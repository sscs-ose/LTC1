* NGSPICE file created from 7b_divider_magic_flat.ext - technology: gf180mcuD

.subckt x7b_divider_magic_flat P2 OUT1 D2_6 D2_2 D2_4 Q5 D2_7 D2_5 Q2 D2_1 Q6 Q3 Q4
+ D2_3 CLK LD Q1 VSS VDD Q7
X0 a_2749_684# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD.t226 VDD.t221 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1 VSS.t103 CLK.t0 a_16065_9774# VSS.t102 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_1209_7469# VDD.t58 VDD.t57 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X3 7b_counter_0.MDFF_6.QB.t0 a_19152_6440# VDD.t1872 VDD.t1871 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X4 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_15865_3363# VSS.t276 VSS.t275 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X5 VDD.t315 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# VDD.t313 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X6 DFF_magic_0.tg_magic_0.IN CLK.t1 DFF_magic_0.tg_magic_3.OUT VSS.t101 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X7 7b_counter_0.3_inp_AND_magic_0.C Q3.t3 a_23207_5885# VDD.t1670 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t11 VSS.t1229 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X9 a_1559_n1526# D2_4.t0 p2_gen_magic_0.xnor_magic_3.OUT VDD.t546 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X10 a_30365_3514# P2.t6 a_30365_4922# VDD.t1473 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X11 VDD.t466 a_14556_n8142# p3_gen_magic_0.3_inp_AND_magic_0.B VDD.t465 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X12 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t472 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X13 VDD.t1672 Q3.t4 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t1671 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X14 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_684# VDD.t661 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X15 VDD.t2029 p3_gen_magic_0.xnor_magic_1.B.t0 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD.t2028 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X16 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_684# VDD.t223 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X17 a_16065_2253# D2_3.t0 VSS.t1183 VSS.t66 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X18 VDD.t810 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_17405_10149# VDD.t806 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X19 7b_counter_0.MDFF_0.QB.t1 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t3 a_5515_3947# VSS.t1171 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X20 p2_gen_magic_0.xnor_magic_1.OUT.t0 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n4081# VDD.t406 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X21 VDD.t665 a_23258_1769# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B VDD.t664 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X22 a_21381_3524# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B VSS.t1279 VSS.t273 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X23 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_19841_9774# VDD.t2176 VDD.t2175 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X24 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t421 VDD.t420 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X25 p3_gen_magic_0.xnor_magic_4.OUT Q2.t3 a_5054_n6471# VSS.t1059 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X26 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t0 VDD.t1814 VDD.t1813 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X27 a_1541_n3597# D2_1.t0 p2_gen_magic_0.xnor_magic_1.OUT VDD.t405 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X28 VDD.t744 p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# VDD.t742 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X29 7b_counter_0.MDFF_5.LD.t5 a_29512_8496.t6 VDD.t1410 VDD.t1409 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X30 a_12174_n8579# p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.AND2_magic_1.A VDD.t549 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X31 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_15865_4557# VSS.t119 VSS.t118 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X32 a_11279_8697# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11191_10149# VDD.t45 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X33 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_5185_2253# VDD.t1553 VDD.t1552 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X34 VDD.t2174 a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD.t2173 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X35 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t9 VDD.t1705 VDD.t1704 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X36 a_12931_7470# D2_2.t0 VSS.t778 VSS.t60 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X37 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_1209_2253# VDD.t2161 VDD.t2160 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X38 a_18891_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_5956# VDD.t2163 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X39 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t9 VSS.t741 VSS.t740 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X40 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_8741# VDD.t371 VDD.t369 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X41 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n1042# VDD.t373 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X42 a_26038_4932# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# VDD.t130 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X43 a_1209_8579# D2_7.t0 VDD.t1950 VDD.t1949 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X44 VSS.t1117 mux_magic_0.IN2.t3 divide_by_2_0.tg_magic_2.IN VSS.t1116 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X45 a_24059_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.D VSS.t362 VSS.t361 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X46 7b_counter_0.MDFF_1.tspc2_magic_0.D a_17405_2092# VDD.t537 VDD.t536 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X47 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK.t2 VSS.t100 VSS.t99 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X48 VDD.t1260 7b_counter_0.NAND_magic_0.A.t6 DFF_magic_0.D.t9 VDD.t1259 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X49 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t3 VDD.t1226 VDD.t1225 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X50 mux_magic_0.AND2_magic_0.A D2_1.t1 VDD.t1777 VDD.t1776 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X51 VDD.t1200 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t3 a_23560_3728# VDD.t531 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X52 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t3 VDD.t1895 VDD.t1894 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X53 VSS.t843 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.P3.t5 VSS.t842 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X54 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT CLK.t4 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VSS.t98 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X55 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t5 VDD.t1910 VDD.t1909 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X56 VDD.t1027 7b_counter_0.MDFF_4.LD.t6 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1026 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X57 a_19307_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK VSS.t1276 VSS.t1275 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X58 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t7 VSS.t592 VSS.t591 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X59 a_7215_10149# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# VDD.t1597 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X60 a_4496_10093# 7b_counter_0.MDFF_3.tspc2_magic_0.D VDD.t1605 VDD.t1603 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X61 a_4651_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t3 VSS.t678 VSS.t677 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X62 a_23985_7877# 7b_counter_0.3_inp_AND_magic_0.B VDD.t1639 VDD.t1637 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X63 VSS.t594 7b_counter_0.MDFF_4.LD.t8 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VSS.t593 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X64 VSS.t97 CLK.t6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS.t96 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X65 VSS.t596 7b_counter_0.MDFF_4.LD.t9 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VSS.t595 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X66 p3_gen_magic_0.3_inp_AND_magic_0.C a_16186_n8142# VSS.t923 VSS.t922 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X67 VSS.t660 D2_5.t0 a_1409_3363# VSS.t31 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X68 VSS.t1093 divide_by_2_1.tg_magic_3.CLK.t0 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VSS.t1092 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X69 VSS.t924 a_11279_1124# 7b_counter_0.MDFF_4.tspc2_magic_0.D VSS.t148 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X70 VDD.t1170 D2_5.t1 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD.t1169 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X71 p2_gen_magic_0.AND2_magic_1.A D2_5.t2 a_12174_n3597# VDD.t407 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X72 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t5 VSS.t958 VSS.t957 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X73 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t10 VSS.t598 VSS.t597 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X74 VDD.t1029 7b_counter_0.MDFF_4.LD.t11 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1028 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X75 a_15865_1059# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VDD.t518 VDD.t517 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X76 VDD.t1031 7b_counter_0.MDFF_4.LD.t12 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t1030 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X77 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t3 VDD.t1428 VDD.t1427 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X78 a_9059_n1973# p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_0.OUT VSS.t250 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X79 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t13 VDD.t1033 VDD.t1032 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X80 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t318 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X81 a_1209_3363# D2_5.t3 VDD.t1172 VDD.t1171 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X82 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t4 VDD.t1838 VDD.t1837 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X83 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t14 VDD.t1035 VDD.t1034 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X84 VDD.t1037 7b_counter_0.MDFF_4.LD.t15 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1036 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X85 a_22991_5885# Q1.t4 VDD.t1228 VDD.t1227 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X86 VDD.t1505 divide_by_2_0.tg_magic_3.CLK.t2 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VDD.t1504 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X87 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.OUT VDD.t1207 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X88 VDD.t1219 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VDD.t1218 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X89 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t3 CLK.t7 VDD.t1912 VDD.t1911 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X90 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_684# VDD.t775 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X91 a_4235_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t4 a_4496_4877# VDD.t2023 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X92 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t6 VSS.t845 VSS.t844 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X93 a_6725_684# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_2092# VDD.t311 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X94 VDD.t716 a_5185_1059# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD.t715 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X95 VSS.t1080 7b_counter_0.MDFF_0.QB.t2 a_1409_4557# VSS.t1079 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X96 a_5185_7469# D2_7.t1 VDD.t1952 VDD.t1951 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X97 VDD.t728 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1209_6275# VDD.t266 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X98 VSS.t588 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT P2.t5 VSS.t587 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X99 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t10 VSS.t743 VSS.t742 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X100 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.VOUT VDD.t501 pfet_03v3 ad=0.4928p pd=3.12u as=1.9712p ps=12.48u w=1.12u l=0.56u
X101 a_15865_3363# 7b_counter_0.MDFF_4.LD.t16 a_16065_3363# VSS.t599 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X102 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t502 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X103 VSS.t980 7b_counter_0.MDFF_5.LD.t10 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VSS.t979 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X104 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t3 VDD.t1507 VDD.t1506 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X105 a_8643_n1526# D2_2.t1 p2_gen_magic_0.xnor_magic_0.OUT VDD.t654 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X106 a_12387_8536# 7b_counter_0.MDFF_5.LD.t11 a_12931_8580# VSS.t981 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X107 p2_gen_magic_0.xnor_magic_3.OUT.t0 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n1042# VDD.t547 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X108 p2_gen_magic_0.xnor_magic_1.OUT.t1 Q7.t3 a_1541_n3150# VSS.t1253 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X109 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t5 CLK.t8 VSS.t95 VSS.t94 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X110 a_8825_1669# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t3 7b_counter_0.MDFF_4.QB.t0 VSS.t1247 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X111 VSS.t93 CLK.t9 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t5 VSS.t92 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X112 a_2749_8740# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B VSS.t112 VSS.t111 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X113 VDD.t25 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n5540# VDD.t24 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X114 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t12 VSS.t983 VSS.t982 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X115 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t6 VDD.t972 VDD.t971 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X116 a_16065_2253# 7b_counter_0.MDFF_4.LD.t17 a_15865_2253# VSS.t600 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X117 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_15865_3363# VDD.t364 VDD.t363 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X118 a_8411_3319# 7b_counter_0.MDFF_4.LD.t18 VDD.t1039 VDD.t1038 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X119 VDD.t649 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11191_684# VDD.t648 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X120 a_1409_1059# Q4.t3 VSS.t873 VSS.t872 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X121 VDD.t1594 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12387_4513# VDD.t1593 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X122 a_11279_3480# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11191_4932# VDD.t77 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X123 VDD.t85 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_5901# VDD.t84 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X124 VDD.t1458 OR_magic_2.A.t6 a_30365_4922# VDD.t1457 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X125 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.NAND_magic_0.VOUT VDD.t733 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X126 a_21381_3524# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_4932# VDD.t2167 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X127 VSS.t1125 D2_7.t2 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS.t1124 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X128 VSS.t91 CLK.t10 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS.t90 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X129 p2_gen_magic_0.3_inp_AND_magic_0.A a_11292_n2115# VSS.t474 VSS.t252 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X130 VDD.t1430 Q6.t4 a_21504_5904# VDD.t1429 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X131 a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_16065_4557# VSS.t911 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X132 VDD.t116 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_26038_684# VDD.t113 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X133 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12931_9774# VSS.t171 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X134 VDD.t1478 p2_gen_magic_0.3_inp_AND_magic_0.C.t1 a_13353_n2115# VDD.t1477 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X135 a_5185_2253# D2_5.t4 VDD.t1174 VDD.t1173 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X136 a_13769_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B a_13553_n2115# VSS.t173 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X137 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t5 VSS.t697 VSS.t696 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X138 VSS.t329 a_26126_1124# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t2 VSS.t178 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X139 VDD.t1041 7b_counter_0.MDFF_4.LD.t19 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1040 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X140 VSS.t331 a_22150_1124# Q4.t2 VSS.t330 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X141 a_9212_739# 7b_counter_0.MDFF_4.tspc2_magic_0.D VSS.t929 VSS.t928 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X142 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t6 a_13353_n6613# VDD.t480 VDD.t478 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X143 VSS.t1231 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t7 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS.t1230 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X144 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t7 7b_counter_0.NAND_magic_0.VOUT VSS.t553 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X145 VDD.t1559 OR_magic_1.VOUT.t2 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VDD.t1558 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X146 a_24536_3947# a_24059_4877# a_23560_3728# VSS.t364 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X147 VSS.t291 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_0.IN VSS.t290 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X148 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t471 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X149 VDD.t2113 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t12 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VDD.t2112 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X150 VDD.t435 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n4081# VDD.t434 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X151 VSS.t1208 p2_gen_magic_0.xnor_magic_3.OUT.t2 a_11708_n2115# VSS.t1207 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X152 VSS.t312 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4235_3947# VSS.t311 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X153 mux_magic_0.IN2.t0 divide_by_2_0.tg_magic_3.IN.t18 VDD.t1983 VDD.t1982 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X154 mux_magic_0.AND2_magic_0.A D2_1.t2 VDD.t1779 VDD.t1778 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X155 VSS.t313 a_11279_6341# 7b_counter_0.MDFF_5.tspc2_magic_0.D VSS.t124 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X156 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t617 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X157 p3_gen_magic_0.3_inp_AND_magic_0.C.t0 a_16186_n8142# VDD.t1609 VDD.t1608 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X158 a_14756_n8142# p3_gen_magic_0.AND2_magic_1.A a_14556_n8142# VSS.t374 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X159 divide_by_2_0.tg_magic_3.IN.t17 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.OUT VDD.t2018 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X160 LD.t0 a_27567_8496.t9 VSS.t576 VSS.t575 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X161 LD.t1 a_27567_8496.t10 VDD.t995 VDD.t994 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X162 a_11492_n6613# p3_gen_magic_0.xnor_magic_4.OUT a_11708_n6613# VSS.t802 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X163 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_19841_8580# VDD.t346 VDD.t345 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X164 VSS.t1184 D2_3.t1 a_16065_2253# VSS.t57 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X165 a_15865_7470# D2_1.t3 VDD.t1781 VDD.t1780 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X166 VDD.t1229 Q1.t6 a_8643_n1526# VDD.t302 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X167 7b_counter_0.MDFF_4.LD.t0 a_31440_8496.t9 VDD.t1924 VDD.t1923 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X168 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_23258_1769# VDD.t663 VDD.t662 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X169 VSS.t274 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_21381_3524# VSS.t273 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X170 7b_counter_0.3_inp_AND_magic_0.C Q3.t6 a_23207_5885# VDD.t1673 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X171 VSS.t1042 D2_6.t1 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS.t1041 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X172 a_17405_10149# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_8741# VDD.t369 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X173 a_5452_n7648# p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.OUT.t1 VSS.t249 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X174 a_5185_1059# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VDD.t368 VDD.t367 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X175 VDD.t431 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_22062_684# VDD.t426 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X176 a_20041_8580# D2_1.t4 VSS.t1018 VSS.t1017 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X177 VDD.t1043 7b_counter_0.MDFF_4.LD.t20 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1042 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X178 VDD.t1412 a_29512_8496.t7 7b_counter_0.MDFF_5.LD.t4 VDD.t1411 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X179 VDD.t1521 Q4.t4 a_1209_1059# VDD.t1520 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X180 VDD.t1162 divide_by_2_1.tg_magic_3.IN.t18 mux_magic_0.IN1.t3 VDD.t1161 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X181 VSS.t803 p3_gen_magic_0.xnor_magic_3.OUT.t2 a_11708_n6613# VSS.t802 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X182 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_3.OUT VDD.t255 VDD.t254 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X183 VDD.t1307 LD.t11 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VDD.t1306 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X184 VDD.t1783 D2_1.t5 p3_gen_magic_0.inverter_magic_0.VOUT VDD.t1782 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X185 VDD.t430 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_22062_684# VDD.t429 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X186 VDD.t1918 CLK.t11 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t1917 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X187 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_15865_6276# VDD.t93 VDD.t35 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X188 divide_by_2_0.tg_magic_3.IN.t9 divide_by_2_0.tg_magic_3.CLK.t4 divide_by_2_0.tg_magic_2.IN VSS.t858 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X189 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_684# VDD.t102 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X190 VSS.t779 D2_2.t2 a_12931_7470# VSS.t55 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X191 p3_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n8579# VDD.t1621 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X192 VSS.t1186 D2_3.t2 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS.t1185 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X193 VSS.t1020 D2_1.t6 mux_magic_0.AND2_magic_0.A VSS.t1019 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X194 DFF_magic_0.D.t2 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.OUT VDD.t229 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X195 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_5901# VDD.t232 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X196 VDD.t1523 Q4.t5 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t1522 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X197 VDD.t1309 LD.t12 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VDD.t1308 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X198 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t13 VDD.t1311 VDD.t1310 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X199 VDD.t988 7b_counter_0.MDFF_4.QB.t2 a_12387_575# VDD.t987 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X200 a_19841_4557# 7b_counter_0.MDFF_1.tspc2_magic_0.Q VDD.t275 VDD.t274 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X201 VDD.t1641 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27234_4513# VDD.t280 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X202 VSS.t1178 p3_gen_magic_0.xnor_magic_1.B.t1 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS.t1177 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X203 a_26126_3480# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26038_4932# VDD.t129 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X204 VDD.t442 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4496_4877# VDD.t441 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X205 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK.t12 VDD.t1905 VDD.t1904 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X206 VSS.t1233 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS.t1232 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X207 VSS.t89 CLK.t13 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS.t88 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X208 DFF_magic_0.tg_magic_2.IN OR_magic_2.A.t7 VDD.t1460 VDD.t1459 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X209 VDD.t1785 D2_1.t7 mux_magic_0.AND2_magic_0.A VDD.t1784 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X210 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t5 VSS.t812 VSS.t811 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X211 VSS.t1153 Q5.t3 7b_counter_0.3_inp_AND_magic_0.A VSS.t1152 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X212 a_20041_9774# 7b_counter_0.MDFF_6.tspc2_magic_0.Q VSS.t198 VSS.t197 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X213 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_3.CLK.t6 DFF_magic_0.D.t5 VSS.t1106 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X214 VSS.t985 7b_counter_0.MDFF_5.LD.t13 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VSS.t984 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X215 VDD.t652 p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# VDD.t650 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X216 a_23793_5904# Q5.t4 7b_counter_0.3_inp_AND_magic_0.A VDD.t1990 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X217 OR_magic_2.A.t3 DFF_magic_0.tg_magic_2.OUT VDD.t1215 VDD.t1214 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X218 VSS.t226 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.IN VSS.t225 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X219 VSS.t781 D2_2.t3 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS.t780 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X220 a_8825_1669# a_8713_1625# VSS.t433 VSS.t432 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X221 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t21 VSS.t602 VSS.t601 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X222 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t22 VSS.t603 VSS.t591 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X223 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.OUT VDD.t738 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X224 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t1 VSS.t1095 VSS.t1094 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X225 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t23 VSS.t605 VSS.t604 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X226 VDD.t637 a_15865_2253# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B VDD.t636 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X227 a_8411_3319# D2_6.t2 VDD.t1816 VDD.t1815 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X228 VSS.t606 7b_counter_0.MDFF_4.LD.t24 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VSS.t593 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X229 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t317 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X230 a_7215_10149# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# VDD.t1596 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X231 a_2749_8740# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_10148# VDD.t18 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X232 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t25 VDD.t1045 VDD.t1044 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X233 VDD.t253 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.IN VDD.t252 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X234 VDD.t500 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.NAND_magic_0.VOUT VDD.t499 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X235 a_11191_10149# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# VDD.t44 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X236 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t1934 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X237 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_8411_8536# VDD.t330 VDD.t329 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X238 VDD.t2073 D2_4.t1 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD.t2072 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X239 mux_magic_0.AND2_magic_0.A D2_1.t8 VDD.t1786 VDD.t1776 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X240 VDD.t1047 7b_counter_0.MDFF_4.LD.t26 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VDD.t1046 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X241 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# VDD.t334 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X242 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT OR_magic_1.VOUT.t3 VDD.t1561 VDD.t1560 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X243 a_11292_n2115# p2_gen_magic_0.xnor_magic_0.OUT a_11492_n2115# VSS.t252 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X244 VDD.t1840 Q2.t5 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t1839 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X245 a_5036_n8579# p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT VDD.t735 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X246 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t5 VSS.t662 VSS.t661 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X247 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VSS.t584 VSS.t583 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X248 a_13769_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B a_13553_n2115# VSS.t173 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X249 a_24401_7877# 7b_counter_0.3_inp_AND_magic_0.B a_24185_7877# VSS.t934 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X250 a_29512_8496.t0 DFF_magic_0.D.t12 VSS.t713 VSS.t712 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X251 a_29512_8496.t1 DFF_magic_0.D.t13 VDD.t1266 VDD.t1265 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X252 VDD.t916 a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD.t915 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X253 a_32616_n2458# mux_magic_0.IN2.t4 VDD.t1938 VDD.t1937 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X254 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.QB.t2 VDD.t1697 VDD.t1696 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X255 VSS.t1212 D2_4.t2 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS.t1211 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X256 a_2749_4932# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD.t931 VDD.t930 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X257 a_22991_5885# Q1.t7 VDD.t1231 VDD.t1230 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X258 a_5470_n1973# p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_4.OUT VSS.t259 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X259 VDD.t1313 LD.t14 a_1209_7469# VDD.t1312 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X260 a_14556_n3644# p2_gen_magic_0.AND2_magic_1.A a_14756_n3644# VSS.t931 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X261 VDD.t342 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.IN VDD.t341 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X262 VSS.t1209 p2_gen_magic_0.xnor_magic_3.OUT.t3 a_11708_n2115# VSS.t1207 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X263 a_9412_739# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t4 a_9212_739# VDD.t2120 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X264 a_23207_5885# Q2.t6 a_22991_5885# VDD.t1841 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X265 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t32 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X266 VDD.t1897 CLK.t14 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t1896 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X267 VDD.t974 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t8 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t973 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X268 VSS.t987 7b_counter_0.MDFF_5.LD.t14 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VSS.t986 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X269 VDD.t1818 D2_6.t3 a_8411_3319# VDD.t1817 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X270 a_15865_7470# 7b_counter_0.MDFF_5.LD.t15 VDD.t1707 VDD.t1706 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X271 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t6 VDD.t1432 VDD.t1431 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X272 a_19152_5956# 7b_counter_0.MDFF_6.tspc2_magic_0.D VDD.t158 VDD.t156 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X273 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t732 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X274 VDD.t162 p2_gen_magic_0.xnor_magic_5.OUT a_16186_n3644# VDD.t161 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X275 a_21381_4932# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD.t360 VDD.t358 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X276 a_20171_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_6.QB.t1 VSS.t1274 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X277 divide_by_2_0.tg_magic_2.IN mux_magic_0.IN2.t5 VDD.t1940 VDD.t1939 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X278 p3_gen_magic_0.AND2_magic_1.A Q4.t6 a_12174_n7648# VSS.t874 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X279 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VDD.t115 VDD.t113 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X280 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# VDD.t111 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X281 a_23672_3947# a_23560_3728# VSS.t461 VSS.t460 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X282 a_12387_3319# 7b_counter_0.MDFF_4.LD.t27 VDD.t1049 VDD.t1048 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X283 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# VDD.t429 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X284 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS.t304 VSS.t303 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X285 VDD.t1315 LD.t15 a_1209_2253# VDD.t1314 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X286 P2.t3 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t1018 VDD.t1017 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X287 VDD.t2075 D2_4.t3 a_27234_3319# VDD.t2074 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X288 a_2749_10148# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD.t922 VDD.t18 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X289 VDD.t1316 LD.t16 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VDD.t1308 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X290 VSS.t377 a_12387_5792# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VSS.t376 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X291 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t4 VSS.t1214 VSS.t1213 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X292 mux_magic_0.IN2.t1 divide_by_2_0.tg_magic_3.IN.t19 VDD.t1985 VDD.t1984 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X293 VSS.t1249 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t5 a_9689_1669# VSS.t1248 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X294 a_12387_1769# 7b_counter_0.MDFF_4.LD.t28 a_12931_2253# VSS.t607 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X295 VDD.t1675 Q3.t7 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t1674 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X296 7b_counter_0.MDFF_7.QB.t1 a_23560_3728# VDD.t709 VDD.t708 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X297 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_1.IN VDD.t793 VDD.t792 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X298 a_17405_10149# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD.t809 VDD.t424 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X299 VDD.t658 a_8713_1625# 7b_counter_0.MDFF_4.QB.t1 VDD.t657 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X300 a_24059_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t4 a_24259_4877# VDD.t1201 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X301 7b_counter_0.3_inp_AND_magic_0.A Q5.t5 a_23793_5904# VDD.t1991 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X302 a_1541_n8579# p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT.t2 VDD.t774 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X303 a_27567_8496.t8 DFF_magic_0.D.t14 VSS.t715 VSS.t714 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X304 a_27567_8496.t5 DFF_magic_0.D.t15 VDD.t1268 VDD.t1267 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X305 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.QB.t2 VDD.t933 VDD.t932 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X306 VDD.t1788 D2_1.t9 a_19841_8580# VDD.t1787 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X307 VSS.t692 DFF_magic_0.tg_magic_2.OUT OR_magic_2.A.t5 VSS.t691 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X308 VDD.t1709 7b_counter_0.MDFF_5.LD.t16 a_15865_7470# VDD.t1708 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X309 a_32616_n1264# mux_magic_0.AND2_magic_0.A a_32816_n1264# VSS.t457 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X310 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t7 VSS.t1061 VSS.t1060 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X311 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t1 a_2749_7308# VDD.t593 VDD.t404 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X312 a_12931_1059# 7b_counter_0.MDFF_4.QB.t3 VSS.t568 VSS.t567 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X313 VDD.t2037 D2_3.t3 a_15865_2253# VDD.t2036 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X314 VSS.t1022 D2_1.t10 a_20041_8580# VSS.t1021 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X315 p3_gen_magic_0.xnor_magic_4.OUT D2_3.t4 a_5054_n6024# VDD.t110 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X316 DFF_magic_0.tg_magic_3.OUT CLK.t15 DFF_magic_0.tg_magic_0.IN VSS.t87 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X317 a_9412_739# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t6 a_9212_739# VDD.t2121 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X318 mux_magic_0.IN1.t2 divide_by_2_1.tg_magic_3.IN.t19 VDD.t1164 VDD.t1163 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X319 VSS.t783 D2_2.t4 a_9059_n6471# VSS.t782 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X320 VSS.t960 Q3.t8 a_27778_1059# VSS.t959 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X321 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t29 VDD.t1051 VDD.t1050 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X322 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t17 VDD.t1318 VDD.t1317 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X323 a_8523_n7648# p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS.t927 VSS.t926 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X324 VSS.t1097 divide_by_2_1.tg_magic_3.CLK.t2 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VSS.t1096 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X325 Q7.t2 a_6725_7308# VSS.t499 VSS.t498 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X326 VDD.t1842 Q2.t8 a_5054_n1526# VDD.t323 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X327 a_27234_3319# 7b_counter_0.MDFF_4.LD.t30 VDD.t1053 VDD.t1052 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X328 a_19152_1223# a_18891_1669# a_19307_1669# VSS.t398 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X329 VDD.t1648 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_19841_4557# VDD.t1647 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X330 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VSS.t1234 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X331 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t3 VDD.t1954 VDD.t1953 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X332 p3_gen_magic_0.xnor_magic_5.OUT.t0 D2_7.t4 a_5036_n8095# VDD.t734 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X333 a_32616_n2458# D2_1.t11 a_32816_n2458# VSS.t1023 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X334 VDD.t707 a_23560_3728# 7b_counter_0.MDFF_7.QB.t1 VDD.t706 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X335 a_24401_7877# 7b_counter_0.3_inp_AND_magic_0.B a_24185_7877# VSS.t934 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X336 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t4 VSS.t1044 VSS.t1043 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X337 VDD.t1901 CLK.t16 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t1900 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X338 VSS.t348 7b_counter_0.3_inp_AND_magic_0.VOUT a_24003_10051# VSS.t347 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X339 a_12387_5792# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t2015 VDD.t1591 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X340 p3_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n8579# VDD.t548 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X341 VSS.t196 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_20041_9774# VSS.t195 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X342 a_17405_5901# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_7309# VDD.t231 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X343 a_16186_n3644# p2_gen_magic_0.xnor_magic_5.OUT a_16386_n3644# VSS.t189 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X344 VSS.t426 a_8411_3319# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B VSS.t425 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X345 VDD.t1993 Q5.t6 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t1992 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X346 VDD.t1433 Q6.t7 a_5036_n3597# VDD.t173 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X347 a_12931_8580# 7b_counter_0.MDFF_5.LD.t17 a_12387_8536# VSS.t988 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X348 VDD.t1213 DFF_magic_0.tg_magic_2.OUT OR_magic_2.A.t2 VDD.t1212 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X349 p3_gen_magic_0.xnor_magic_3.OUT.t1 Q3.t9 a_1559_n6471# VSS.t961 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X350 VDD.t10 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_15865_9774# VDD.t9 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X351 a_7215_10149# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VDD.t289 VDD.t287 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X352 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t5 VDD.t1820 VDD.t1819 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X353 VDD.t293 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11191_4932# VDD.t80 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X354 divide_by_2_0.tg_magic_2.IN mux_magic_0.IN2.t6 VSS.t1119 VSS.t1118 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X355 DFF_magic_0.tg_magic_1.IN CLK.t17 DFF_magic_0.tg_magic_2.OUT VSS.t86 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X356 a_27234_1769# 7b_counter_0.MDFF_4.LD.t31 a_27778_2253# VSS.t608 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X357 VDD.t1877 divide_by_2_1.tg_magic_3.CLK.t3 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VDD.t1876 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X358 VDD.t641 a_8411_3319# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B VDD.t640 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X359 a_12387_575# 7b_counter_0.MDFF_4.QB.t4 VDD.t990 VDD.t989 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X360 a_12387_4513# Q5.t7 VDD.t1994 VDD.t52 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X361 a_27778_1059# Q3.t10 VSS.t963 VSS.t962 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X362 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t32 VSS.t609 VSS.t604 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X363 Q5.t1 a_6725_2092# VDD.t312 VDD.t311 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X364 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_12387_8536# VDD.t2022 VDD.t2021 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X365 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t2 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t172 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X366 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT OR_magic_2.VOUT.t3 VSS.t808 VSS.t807 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X367 a_11279_8697# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VSS.t695 VSS.t150 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X368 a_18891_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_739# VDD.t575 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X369 VSS.t391 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VSS.t390 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X370 p3_gen_magic_0.xnor_magic_3.OUT D2_4.t5 a_1559_n6024# VDD.t561 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X371 a_12931_9774# 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12387_9730# VSS.t170 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X372 p3_gen_magic_0.xnor_magic_6.OUT Q5.t8 a_8523_n7648# VSS.t1154 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X373 VDD.t553 p3_gen_magic_0.AND2_magic_1.A a_14556_n8142# VDD.t552 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X374 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT CLK.t18 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VSS.t85 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X375 VDD.t956 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.NAND_magic_0.A.t3 VDD.t955 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X376 VDD.t1563 OR_magic_1.VOUT.t4 divide_by_2_1.inverter_magic_5.VOUT VDD.t1562 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X377 a_5054_n1973# p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS.t281 VSS.t280 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X378 7b_counter_0.3_inp_AND_magic_0.B Q6.t8 VSS.t814 VSS.t813 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X379 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN P2.t7 VDD.t2061 VDD.t2060 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X380 VDD.t1055 7b_counter_0.MDFF_4.LD.t33 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1054 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X381 VDD.t1386 D2_2.t5 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD.t1385 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X382 VDD.t1487 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.P3.t3 VDD.t1486 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X383 VDD.t1435 Q6.t9 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t1434 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X384 VSS.t1255 Q7.t4 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VSS.t1254 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X385 a_23258_575# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1587 VDD.t1586 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X386 VSS.t1156 Q5.t9 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VSS.t1155 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X387 VDD.t992 7b_counter_0.MDFF_4.QB.t5 7b_counter_0.MDFF_4.tspc2_magic_0.Q VDD.t991 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X388 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t5 VDD.t1509 VDD.t1508 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X389 VDD.t2157 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.IN VDD.t2156 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X390 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t2 CLK.t19 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS.t84 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X391 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.IN VDD.t31 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X392 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t11 VDD.t1677 VDD.t1676 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X393 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12387_9730# VDD.t1217 VDD.t1216 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X394 VDD.t1557 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_19841_9774# VDD.t1556 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X395 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.A VDD.t217 pfet_03v3 ad=0.4928p pd=3.12u as=1.9712p ps=12.48u w=1.12u l=0.56u
X396 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t18 VDD.t1711 VDD.t1710 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X397 VDD.t510 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN VDD.t509 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X398 a_5385_6275# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5185_6275# VSS.t220 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X399 a_23352_n6798# p3_gen_magic_0.P3.t6 VSS.t1143 VSS.t1142 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X400 VDD.t698 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_17405_684# VDD.t697 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X401 a_15865_1059# 7b_counter_0.MDFF_1.QB.t3 VDD.t935 VDD.t934 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X402 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n5540# VDD.t563 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X403 VDD.t1790 D2_1.t12 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD.t1789 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X404 VSS.t368 7b_counter_0.MDFF_1.tspc2_magic_0.D a_18891_1669# VSS.t367 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X405 VDD.t2166 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_6440# VDD.t154 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X406 VDD.t1150 mux_magic_0.IN1.t6 a_32616_n1264# VDD.t1149 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X407 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t9 VDD.t976 VDD.t975 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X408 a_11292_n2115# p2_gen_magic_0.xnor_magic_4.OUT VDD.t126 VDD.t124 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X409 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT CLK.t20 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t1 VSS.t83 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X410 7b_counter_0.MDFF_6.QB.t1 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_20171_6886# VSS.t1273 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X411 VDD.t1437 Q6.t10 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t1436 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X412 a_8713_6842# a_9212_5956# a_9689_6886# VSS.t574 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X413 divide_by_2_0.tg_magic_3.CLK.t0 OR_magic_2.VOUT.t4 VDD.t1422 VDD.t1421 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X414 a_17405_3524# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_4932# VDD.t40 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X415 VSS.t529 7b_counter_0.MDFF_7.QB.t2 7b_counter_0.MDFF_7.tspc2_magic_0.Q VSS.t528 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X416 7b_counter_0.MDFF_5.LD.t8 a_29512_8496.t8 VSS.t797 VSS.t796 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X417 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1209_6275# VSS.t471 VSS.t470 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X418 VDD.t1916 CLK.t21 a_12387_3319# VDD.t1915 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X419 7b_counter_0.MDFF_5.LD.t3 a_29512_8496.t9 VDD.t1414 VDD.t1413 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X420 a_19841_3363# 7b_counter_0.MDFF_4.LD.t34 a_20041_3363# VSS.t610 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X421 divide_by_2_1.tg_magic_3.IN.t2 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT divide_by_2_1.tg_magic_1.IN VDD.t380 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X422 a_27234_3319# D2_4.t6 VDD.t2077 VDD.t2076 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X423 OUT1.t1 a_34156_n2297# VDD.t383 VDD.t381 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X424 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t13 VDD.t2115 VDD.t2114 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X425 a_23352_n6798# p3_gen_magic_0.P3.t7 a_23352_n5390# VDD.t1468 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X426 a_9689_1669# a_9212_739# a_8713_1625# VSS.t333 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X427 VDD.t387 a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD.t386 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X428 VSS.t121 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_17405_3524# VSS.t120 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X429 VDD.t1713 7b_counter_0.MDFF_5.LD.t19 a_12387_6986# VDD.t1712 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X430 VSS.t512 p3_gen_magic_0.xnor_magic_1.OUT.t3 a_16386_n8142# VSS.t511 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X431 VSS.t82 CLK.t22 DFF_magic_0.tg_magic_3.CLK.t5 VSS.t81 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X432 a_17405_8741# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B VSS.t307 VSS.t214 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X433 a_5385_7469# LD.t18 a_5185_7469# VSS.t744 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X434 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t2 a_2749_2092# VSS.t211 VSS.t210 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X435 a_29512_8496.t2 DFF_magic_0.D.t16 VDD.t1270 VDD.t1269 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X436 VDD.t1320 LD.t19 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VDD.t1319 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X437 7b_counter_0.MDFF_4.QB.t1 a_8713_1625# VDD.t656 VDD.t655 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X438 a_24259_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t5 a_24059_4877# VDD.t1202 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X439 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.QB VSS.t139 VSS.t138 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X440 a_12174_n8095# Q4.t7 VDD.t1524 VDD.t238 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X441 VDD.t1636 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n5540# VDD.t1635 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X442 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT divide_by_2_0.tg_magic_0.IN VDD.t196 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X443 a_1559_n1973# p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS.t370 VSS.t369 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X444 divide_by_2_1.tg_magic_3.IN.t5 OR_magic_1.VOUT.t5 divide_by_2_1.tg_magic_1.IN VSS.t892 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X445 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t7 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS.t846 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X446 a_11191_10149# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VDD.t1224 VDD.t1220 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X447 VSS.t80 CLK.t23 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t5 VSS.t79 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X448 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_1209_7469# VSS.t133 VSS.t132 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X449 a_14556_n3644# p2_gen_magic_0.xnor_magic_6.OUT VDD.t759 VDD.t758 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X450 a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_20041_4557# VSS.t938 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X451 VSS.t570 7b_counter_0.MDFF_4.QB.t6 a_12931_1059# VSS.t569 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X452 VDD.t1321 LD.t20 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VDD.t1306 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X453 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t8 p2_gen_magic_0.3_inp_AND_magic_0.VOUT VSS.t847 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X454 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_3.OUT VDD.t2155 VDD.t2154 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X455 a_27778_1059# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27234_575# VSS.t354 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X456 VDD.t1419 p3_gen_magic_0.xnor_magic_3.OUT.t3 a_11292_n6613# VDD.t1418 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X457 a_21381_8741# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_10149# VDD.t348 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X458 divide_by_2_1.tg_magic_3.IN.t14 divide_by_2_1.tg_magic_3.CLK.t4 divide_by_2_1.tg_magic_2.IN VSS.t1098 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X459 a_23802_1059# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23258_575# VSS.t913 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X460 VDD.t1893 DFF_magic_0.tg_magic_3.CLK.t7 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t1892 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X461 a_11708_n6613# p3_gen_magic_0.xnor_magic_4.OUT a_11492_n6613# VSS.t925 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X462 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t7 VDD.t2079 VDD.t2078 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X463 7b_counter_0.3_inp_AND_magic_0.C Q3.t12 a_23207_5885# VDD.t1673 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X464 VDD.t1223 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11191_10149# VDD.t1220 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X465 a_21504_5904# Q6.t11 VDD.t1439 VDD.t1438 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X466 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_5185_1059# VSS.t463 VSS.t462 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X467 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t9 VDD.t1844 VDD.t1843 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X468 a_11708_n6613# p3_gen_magic_0.xnor_magic_4.OUT a_11492_n6613# VSS.t925 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X469 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t9 VDD.t1489 VDD.t1488 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X470 a_2749_4932# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_3524# VDD.t404 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X471 VDD.t49 7b_counter_0.MDFF_5.QB.t2 a_12387_5792# VDD.t48 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X472 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VDD.t1010 VDD.t1009 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X473 VDD.t2039 D2_3.t5 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD.t2038 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X474 VSS.t203 a_12387_3319# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B VSS.t202 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X475 VDD.t514 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27234_575# VDD.t513 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X476 VDD.t1424 OR_magic_2.VOUT.t5 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VDD.t1423 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X477 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.QB.t3 VDD.t1865 VDD.t1864 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X478 a_1957_n7648# p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT.t1 VSS.t492 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X479 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.NAND_magic_0.A.t7 VDD.t1262 VDD.t1261 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X480 divide_by_2_0.tg_magic_1.IN OR_magic_2.VOUT.t6 divide_by_2_0.tg_magic_3.IN.t3 VSS.t809 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X481 VDD.t308 p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# VDD.t306 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X482 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t6 VSS.t860 VSS.t859 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X483 VDD.t377 a_19841_3363# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B VDD.t376 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X484 VDD.t1462 OR_magic_2.A.t8 DFF_magic_0.tg_magic_2.IN VDD.t1461 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X485 a_2749_684# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_2092# VDD.t204 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X486 a_23802_2253# D2_4.t8 VSS.t1216 VSS.t1215 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X487 VDD.t247 a_1209_1059# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD.t246 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X488 VSS.t1127 D2_7.t5 a_5452_n3150# VSS.t1126 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X489 VDD.t1974 p3_gen_magic_0.P3.t8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VDD.t1973 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X490 VDD.t705 mux_magic_0.AND2_magic_0.A a_32616_n1264# VDD.t704 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X491 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t10 VDD.t978 VDD.t977 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X492 VSS.t193 a_7303_3480# Q6.t2 VSS.t192 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X493 VSS.t582 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VSS.t581 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X494 VDD.t1388 D2_2.t6 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD.t1387 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X495 VSS.t145 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VSS.t144 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X496 a_17405_5901# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD.t98 VDD.t37 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X497 a_18891_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_739# VDD.t574 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X498 VDD.t193 a_12387_3319# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B VDD.t192 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X499 7b_counter_0.MDFF_4.LD.t1 a_31440_8496.t10 VSS.t1110 VSS.t1109 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X500 a_1209_6275# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1409_6275# VSS.t469 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X501 a_16186_n8142# p3_gen_magic_0.xnor_magic_5.OUT.t2 VDD.t1920 VDD.t1919 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X502 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t8 VDD.t1526 VDD.t1525 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X503 7b_counter_0.MDFF_4.LD.t2 a_31440_8496.t11 VDD.t1926 VDD.t1925 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X504 divide_by_2_1.inverter_magic_5.VOUT OR_magic_1.VOUT.t6 VDD.t1565 VDD.t1564 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X505 VDD.t83 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_5901# VDD.t76 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X506 VDD.t2097 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t10 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t2096 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X507 VDD.t1426 OR_magic_2.VOUT.t7 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VDD.t1425 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X508 VSS.t185 a_4496_4393# a_5515_3947# VSS.t184 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X509 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_15865_7470# VSS.t272 VSS.t271 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X510 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t13 VDD.t1679 VDD.t1678 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X511 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_3.OUT VSS.t1269 VSS.t1268 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X512 VDD.t1866 7b_counter_0.MDFF_0.QB.t4 a_1209_4557# VDD.t1446 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X513 a_12931_2253# 7b_counter_0.MDFF_4.LD.t35 a_12387_1769# VSS.t611 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X514 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.CLK.t5 divide_by_2_1.tg_magic_3.IN.t11 VSS.t1099 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X515 a_17405_4932# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD.t42 VDD.t37 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X516 a_5515_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t4 7b_counter_0.MDFF_3.QB VSS.t679 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X517 a_8643_n1973# p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS.t429 VSS.t428 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X518 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_3.OUT VDD.t2153 VDD.t2152 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X519 a_17405_8741# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_10149# VDD.t424 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X520 VDD.t1956 D2_7.t6 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD.t1955 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X521 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t30 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X522 mux_magic_0.IN2.t2 divide_by_2_0.tg_magic_3.IN.t20 VSS.t1149 VSS.t1148 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X523 p2_gen_magic_0.xnor_magic_1.OUT D2_1.t13 a_1541_n3597# VDD.t406 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X524 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t24 VSS.t78 VSS.t77 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X525 a_8523_n8095# Q5.t10 VDD.t1995 VDD.t600 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X526 p2_gen_magic_0.xnor_magic_5.OUT p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n4081# VDD.t108 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X527 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t508 VDD.t507 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X528 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t6 VSS.t1188 VSS.t1187 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X529 a_1209_7469# LD.t21 a_1409_7469# VSS.t745 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X530 a_2749_5900# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD.t633 VDD.t631 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X531 a_16186_n3644# p2_gen_magic_0.xnor_magic_1.OUT.t2 VDD.t1861 VDD.t1860 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X532 VDD.t1233 Q1.t8 a_12387_9730# VDD.t1232 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X533 a_8411_8536# 7b_counter_0.MDFF_5.LD.t20 a_8955_8580# VSS.t989 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X534 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK.t25 VDD.t1899 VDD.t1898 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X535 a_32616_n1264# mux_magic_0.IN1.t7 VDD.t1152 VDD.t1151 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X536 VDD.t980 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t11 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t979 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X537 divide_by_2_0.tg_magic_0.IN OR_magic_2.VOUT.t8 divide_by_2_0.tg_magic_3.OUT VSS.t810 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X538 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_1209_8579# VDD.t137 VDD.t136 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X539 a_22991_5885# Q1.t9 VDD.t1234 VDD.t1230 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X540 VSS.t375 a_27234_3319# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B VSS.t247 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X541 a_20171_6886# a_19152_6440# VSS.t1088 VSS.t1087 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X542 a_9689_6886# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t3 VSS.t205 VSS.t204 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X543 VDD.t1322 LD.t22 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VDD.t1306 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X544 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT OR_magic_1.VOUT.t7 VDD.t1567 VDD.t1566 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X545 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_27234_575# VDD.t763 VDD.t762 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X546 VDD.t1569 OR_magic_1.VOUT.t8 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VDD.t1568 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X547 VDD.t526 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8411_4513# VDD.t525 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X548 VSS.t200 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_6725_7308# VSS.t199 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X549 VDD.t627 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23258_575# VDD.t626 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X550 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t1 VDD.t379 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X551 VSS.t649 mux_magic_0.IN1.t8 divide_by_2_1.tg_magic_2.IN VSS.t648 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X552 VDD.t1154 mux_magic_0.IN1.t9 divide_by_2_1.tg_magic_2.IN VDD.t1153 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X553 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t7 VDD.t1390 VDD.t1389 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X554 a_1209_1059# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VDD.t484 VDD.t483 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X555 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t8 VSS.t785 VSS.t784 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X556 a_5185_1059# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5385_1059# VSS.t278 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X557 VDD.t1272 DFF_magic_0.D.t17 a_29512_8496.t3 VDD.t1271 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X558 VDD.t1903 CLK.t26 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t1902 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X559 a_4235_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t5 a_4496_10093# VDD.t1193 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X560 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8955_9774# VSS.t340 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X561 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t5 VDD.t2126 VDD.t2125 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X562 VDD.t559 a_12387_5792# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VDD.t73 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X563 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK.t27 VSS.t76 VSS.t75 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X564 VDD.t492 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VDD.t491 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X565 VSS.t242 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VSS.t241 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X566 a_5385_2253# LD.t23 a_5185_2253# VSS.t746 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X567 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_1209_3363# VDD.t322 VDD.t321 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X568 divide_by_2_1.tg_magic_0.IN OR_magic_1.VOUT.t9 divide_by_2_1.tg_magic_3.OUT VSS.t893 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X569 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n2115# VSS.t477 VSS.t476 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X570 p2_gen_magic_0.xnor_magic_0.OUT Q1.t10 a_8643_n1973# VSS.t698 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X571 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t11 VDD.t1997 VDD.t1996 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X572 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t24 VDD.t1324 VDD.t1323 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X573 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t25 VDD.t1326 VDD.t1325 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X574 a_12387_575# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1025 VDD.t1024 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X575 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_1209_2253# VSS.t1270 VSS.t257 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X576 a_21381_10149# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD.t413 VDD.t410 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X577 p3_gen_magic_0.3_inp_AND_magic_0.A a_11292_n6613# VDD.t766 VDD.t764 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X578 VDD.t1057 7b_counter_0.MDFF_4.LD.t36 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1056 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X579 a_6725_684# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD.t722 VDD.t719 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X580 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B VSS.t319 VSS.t318 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X581 VDD.t2099 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t11 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t2098 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X582 a_13353_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B VDD.t469 VDD.t467 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X583 a_12590_n3150# p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.AND2_magic_1.A VSS.t181 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X584 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B VSS.t294 VSS.t111 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X585 a_14756_n8142# p3_gen_magic_0.xnor_magic_6.OUT VSS.t163 VSS.t162 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X586 VDD.t301 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n8579# VDD.t300 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X587 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t37 VDD.t1059 VDD.t1058 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X588 VDD.t1061 7b_counter_0.MDFF_4.LD.t38 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t1060 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X589 VDD.t169 a_7303_3480# Q6.t1 VDD.t167 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X590 VDD.t1062 7b_counter_0.MDFF_4.LD.t39 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1028 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X591 p2_gen_magic_0.xnor_magic_0.OUT D2_2.t9 a_8643_n1526# VDD.t653 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X592 a_13553_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B a_13769_n6613# VSS.t328 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X593 VDD.t220 VDD.t219 VDD.t220 VDD.t70 pfet_03v3 ad=0.4928p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X594 divide_by_2_1.inverter_magic_5.VOUT OR_magic_1.VOUT.t10 VDD.t1571 VDD.t1570 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X595 VDD.t1063 7b_counter_0.MDFF_4.LD.t40 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t1030 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X596 VDD.t2081 D2_4.t9 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD.t2080 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X597 VDD.t297 a_27234_1769# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B VDD.t296 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X598 a_15865_7470# 7b_counter_0.MDFF_5.LD.t21 a_16065_7470# VSS.t990 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X599 a_2749_3524# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_4932# VDD.t403 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X600 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t41 VDD.t1064 VDD.t1032 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X601 p3_gen_magic_0.P3.t4 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS.t841 VSS.t840 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X602 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t28 VSS.t74 VSS.t73 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X603 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t42 VDD.t1065 VDD.t1034 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X604 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN VDD.t712 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X605 a_16065_6276# 7b_counter_0.MDFF_6.QB.t3 VSS.t974 VSS.t973 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X606 VDD.t1008 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VDD.t1007 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X607 divide_by_2_1.tg_magic_3.OUT OR_magic_1.VOUT.t11 divide_by_2_1.tg_magic_0.IN VSS.t894 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X608 VDD.t148 a_4496_4393# 7b_counter_0.MDFF_0.QB.t0 VDD.t147 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X609 VDD.t1976 p3_gen_magic_0.P3.t9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VDD.t1975 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X610 VDD.t1264 7b_counter_0.NAND_magic_0.A.t8 7b_counter_0.DFF_magic_0.tg_magic_2.IN VDD.t1263 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X611 VSS.t1089 p3_gen_magic_0.3_inp_AND_magic_0.C.t1 a_13769_n6613# VSS.t327 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X612 VSS.t137 7b_counter_0.MDFF_3.QB a_1409_9773# VSS.t136 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X613 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT DFF_magic_0.tg_magic_1.IN VDD.t91 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X614 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t506 VDD.t505 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X615 7b_counter_0.3_inp_AND_magic_0.C Q3.t14 a_23207_5885# VDD.t1670 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X616 a_1409_8579# LD.t26 a_1209_8579# VSS.t747 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X617 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t29 VDD.t1703 VDD.t502 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X618 VDD.t2101 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t12 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t2100 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X619 a_13553_n2115# p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# VSS.t475 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X620 VSS.t991 7b_counter_0.MDFF_5.LD.t22 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VSS.t979 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X621 VDD.t398 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_0.IN VDD.t397 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X622 a_32616_n1264# mux_magic_0.AND2_magic_0.A VDD.t703 VDD.t702 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X623 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_684# VDD.t660 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X624 DFF_magic_0.D.t11 7b_counter_0.NAND_magic_0.A.t9 VSS.t731 VSS.t730 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X625 VDD.t1680 Q3.t15 a_1559_n1526# VDD.t802 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X626 VSS.t993 7b_counter_0.MDFF_5.LD.t23 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VSS.t992 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X627 a_12174_n4081# p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t141 VDD.t140 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X628 VSS.t149 a_11279_3480# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t2 VSS.t148 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X629 VDD.t412 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_21381_10149# VDD.t410 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X630 VSS.t1090 p3_gen_magic_0.3_inp_AND_magic_0.C.t2 a_13769_n6613# VSS.t328 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X631 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_684# VDD.t223 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X632 VSS.t828 OR_magic_2.A.t9 a_30365_3514# VSS.t827 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X633 VDD.t958 DFF_magic_0.tg_magic_3.CLK.t8 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t957 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X634 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t24 VSS.t995 VSS.t994 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X635 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.B.t2 VDD.t2031 VDD.t2030 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X636 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_3.CLK.t9 DFF_magic_0.D.t3 VSS.t540 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X637 Q3.t1 a_21381_3524# VDD.t2172 VDD.t2170 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X638 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t25 VSS.t996 VSS.t982 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X639 VSS.t664 D2_5.t6 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS.t663 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X640 a_31440_8496.t8 DFF_magic_0.D.t18 VSS.t717 VSS.t716 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X641 a_1409_6275# Q6.t12 VSS.t816 VSS.t815 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X642 7b_counter_0.MDFF_3.tspc2_magic_0.D a_2749_8740# VDD.t21 VDD.t20 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X643 a_31440_8496.t5 DFF_magic_0.D.t19 VDD.t1274 VDD.t1273 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X644 VSS.t1112 a_31440_8496.t12 7b_counter_0.MDFF_4.LD.t3 VSS.t1111 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X645 VDD.t1928 a_31440_8496.t13 7b_counter_0.MDFF_4.LD.t4 VDD.t1927 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X646 a_9412_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t4 a_9212_5956# VDD.t197 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X647 VDD.t1958 D2_7.t7 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD.t1957 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X648 VSS.t1091 p3_gen_magic_0.3_inp_AND_magic_0.C.t3 a_13769_n6613# VSS.t327 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X649 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t16 VDD.t2017 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X650 VDD.t2127 Q7.t6 a_1541_n3597# VDD.t434 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X651 divide_by_2_0.tg_magic_3.CLK.t1 OR_magic_2.VOUT.t9 VSS.t944 VSS.t943 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X652 a_1209_4557# 7b_counter_0.MDFF_0.QB.t5 VDD.t1867 VDD.t1449 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X653 Q1.t2 a_21381_8741# VSS.t494 VSS.t493 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X654 P2.t4 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS.t586 VSS.t585 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X655 VDD.t1067 7b_counter_0.MDFF_4.LD.t43 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t1066 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X656 VDD.t366 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5185_1059# VDD.t365 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X657 a_12387_6986# D2_2.t10 VDD.t1392 VDD.t1391 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X658 VSS.t213 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_2749_2092# VSS.t212 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X659 VDD.t1068 7b_counter_0.MDFF_4.LD.t44 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1036 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X660 divide_by_2_1.tg_magic_3.IN.t10 divide_by_2_1.tg_magic_3.CLK.t6 divide_by_2_1.tg_magic_3.OUT VSS.t1100 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X661 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t6 a_5515_9163# VSS.t680 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X662 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VDD.t428 VDD.t426 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X663 VDD.t243 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5185_6275# VDD.t242 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X664 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t45 VDD.t1070 VDD.t1069 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X665 7b_counter_0.MDFF_1.tspc2_magic_0.D a_17405_2092# VDD.t535 VDD.t534 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X666 VDD.t1071 7b_counter_0.MDFF_4.LD.t46 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1040 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X667 a_12174_n7648# p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS.t372 VSS.t371 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X668 a_1409_7469# CLK.t30 VSS.t72 VSS.t71 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X669 7b_counter_0.MDFF_6.tspc2_magic_0.D a_17405_7309# VDD.t235 VDD.t234 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X670 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN CLK.t31 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS.t70 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X671 a_8955_8580# D2_2.t11 VSS.t787 VSS.t786 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X672 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_3.CLK.t7 divide_by_2_0.tg_magic_3.IN.t8 VSS.t861 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X673 VDD.t1822 D2_6.t6 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD.t1821 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X674 a_13353_n2115# p2_gen_magic_0.3_inp_AND_magic_0.A a_13553_n2115# VSS.t476 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X675 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t7 VSS.t1257 VSS.t1256 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X676 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_12387_1769# VDD.t785 VDD.t784 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X677 a_1209_2253# LD.t27 a_1409_2253# VSS.t748 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X678 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t28 VDD.t1328 VDD.t1327 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X679 VDD.t1073 7b_counter_0.MDFF_4.LD.t47 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD.t1072 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X680 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_15865_4557# VDD.t36 VDD.t35 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X681 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT OR_magic_1.VOUT.t12 VDD.t1573 VDD.t1572 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X682 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t524 VDD.t523 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X683 VDD.t1330 LD.t29 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VDD.t1329 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X684 VDD.t1906 CLK.t32 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t502 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X685 a_16386_n8142# p3_gen_magic_0.xnor_magic_1.OUT.t4 VSS.t514 VSS.t513 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X686 a_15865_8580# CLK.t33 VDD.t1908 VDD.t1907 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X687 a_4235_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t7 a_4496_10093# VDD.t1194 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X688 a_8939_n3150# p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.OUT VSS.t106 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X689 VDD.t1074 7b_counter_0.MDFF_4.LD.t48 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1042 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X690 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.QB.t4 VDD.t937 VDD.t936 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X691 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t8 VDD.t778 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X692 a_5385_1059# 7b_counter_0.MDFF_0.tspc2_magic_0.Q VSS.t484 VSS.t483 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X693 VDD.t1332 LD.t30 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VDD.t1331 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X694 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN P2.t8 VSS.t1202 VSS.t1201 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X695 VSS.t179 a_26126_3480# 7b_counter_0.MDFF_7.tspc2_magic_0.D VSS.t178 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X696 a_8955_9774# 7b_counter_0.MDFF_5.tspc2_magic_0.Q VSS.t443 VSS.t442 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X697 7b_counter_0.3_inp_AND_magic_0.VOUT a_23985_7877# VDD.t2149 VDD.t2147 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X698 VDD.t1333 LD.t31 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VDD.t1306 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X699 VDD.t929 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_2749_4932# VDD.t631 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X700 a_22991_5885# Q1.t11 VDD.t1235 VDD.t1227 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X701 a_16065_6276# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_15865_6276# VSS.t117 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X702 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_3.CLK.t10 DFF_magic_0.tg_magic_2.OUT VSS.t541 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X703 a_7303_8697# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7215_10149# VDD.t1595 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X704 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.VOUT VDD.t498 VDD.t497 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X705 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t7 VDD.t2041 VDD.t2040 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X706 a_23207_5885# Q2.t10 a_22991_5885# VDD.t1841 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X707 VDD.t445 a_11279_6341# 7b_counter_0.MDFF_5.tspc2_magic_0.D VDD.t77 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X708 VDD.t533 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24259_4877# VDD.t529 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X709 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t10 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS.t848 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X710 VDD.t1914 CLK.t34 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t2 VDD.t1913 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X711 VDD.t1999 Q5.t12 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t1998 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X712 VSS.t1190 D2_3.t8 a_5470_n6471# VSS.t1189 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X713 VSS.t997 7b_counter_0.MDFF_5.LD.t26 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VSS.t984 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X714 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t14 VSS.t1244 VSS.t1243 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X715 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t32 VSS.t750 VSS.t749 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X716 VSS.t383 a_23258_575# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VSS.t382 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X717 a_13553_n2115# p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# VSS.t475 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X718 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1209_9773# VDD.t914 VDD.t913 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X719 a_8523_n4081# p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t6 VDD.t5 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X720 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t10 VDD.t1644 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X721 VDD.t1076 7b_counter_0.MDFF_4.LD.t49 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1075 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X722 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t4 CLK.t35 VSS.t69 VSS.t68 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X723 a_17405_3524# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_4932# VDD.t230 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X724 VDD.t1078 7b_counter_0.MDFF_4.LD.t50 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VDD.t1077 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X725 VDD.t79 a_11279_3480# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t1 VDD.t77 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X726 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t27 VDD.t1715 VDD.t1714 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X727 p2_gen_magic_0.xnor_magic_4.OUT Q2.t11 a_5054_n1973# VSS.t1062 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X728 a_30365_4922# OR_magic_2.A.t10 VDD.t1463 VDD.t1457 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X729 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t51 VDD.t1079 VDD.t1044 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X730 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_15865_9774# VDD.t14 VDD.t13 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X731 VDD.t362 a_15865_3363# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B VDD.t361 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X732 a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VDD.t1555 VDD.t1554 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X733 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_27234_1769# VDD.t295 VDD.t294 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X734 a_5515_3947# a_4496_4393# VSS.t183 VSS.t182 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X735 a_11292_n6613# p3_gen_magic_0.xnor_magic_4.OUT VDD.t1619 VDD.t1617 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X736 VDD.t812 CLK.t36 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t811 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X737 VDD.t1080 7b_counter_0.MDFF_4.LD.t52 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VDD.t1046 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X738 VSS.t976 7b_counter_0.MDFF_6.QB.t4 a_16065_6276# VSS.t975 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X739 VDD.t114 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_26038_684# VDD.t113 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X740 VSS.t1272 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19307_6886# VSS.t1271 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X741 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t7 VDD.t1176 VDD.t1175 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X742 a_4496_4877# 7b_counter_0.MDFF_0.tspc2_magic_0.D VDD.t440 VDD.t436 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X743 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.NAND_magic_0.A.t10 VDD.t1293 VDD.t1292 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X744 VDD.t820 CLK.t37 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t819 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X745 Q1.t1 a_21381_8741# VDD.t772 VDD.t349 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X746 VDD.t1082 7b_counter_0.MDFF_4.LD.t53 a_23258_1769# VDD.t1081 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X747 VDD.t396 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_0.IN VDD.t395 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X748 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.OUT VDD.t90 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X749 a_19152_5956# 7b_counter_0.MDFF_6.tspc2_magic_0.D VDD.t157 VDD.t156 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X750 a_11279_1124# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VSS.t427 VSS.t245 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X751 a_8955_8580# 7b_counter_0.MDFF_5.LD.t28 a_8411_8536# VSS.t998 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X752 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t29 VSS.t1000 VSS.t999 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X753 VDD.t1335 LD.t33 a_1209_8579# VDD.t1334 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X754 VSS.t684 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t6 a_24536_3947# VSS.t683 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X755 a_1409_3363# LD.t34 a_1209_3363# VSS.t751 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X756 7b_counter_0.MDFF_5.QB.t0 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t5 a_8825_6886# VSS.t206 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X757 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_15865_1059# VSS.t358 VSS.t357 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X758 VDD.t586 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7215_4932# VDD.t580 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X759 a_21381_10149# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_8741# VDD.t349 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X760 p2_gen_magic_0.3_inp_AND_magic_0.C a_16186_n3644# VSS.t191 VSS.t190 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X761 a_23560_3728# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t7 VDD.t1203 VDD.t527 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X762 VSS.t1001 7b_counter_0.MDFF_5.LD.t30 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VSS.t986 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X763 VSS.t719 DFF_magic_0.D.t20 a_31440_8496.t7 VSS.t718 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X764 VDD.t1276 DFF_magic_0.D.t21 a_31440_8496.t4 VDD.t1275 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X765 a_8411_4513# 7b_counter_0.MDFF_4.tspc2_magic_0.Q VDD.t605 VDD.t604 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X766 a_34156_n889# mux_magic_0.OR_magic_0.A VDD.t614 VDD.t610 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X767 a_19841_8580# 7b_counter_0.MDFF_5.LD.t31 VDD.t1717 VDD.t1716 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X768 VSS.t1218 D2_4.t10 a_1975_n6471# VSS.t1217 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X769 VDD.t791 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_0.IN VDD.t790 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X770 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t16 VSS.t965 VSS.t964 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X771 p3_gen_magic_0.xnor_magic_1.OUT.t2 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n8579# VDD.t773 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X772 VDD.t1196 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t8 a_4496_9609# VDD.t1195 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X773 VSS.t921 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4235_9163# VSS.t920 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X774 a_15865_8580# 7b_counter_0.MDFF_5.LD.t32 VDD.t1719 VDD.t1718 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X775 VDD.t314 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# VDD.t313 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X776 a_7303_8697# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VSS.t244 VSS.t243 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X777 a_8955_9774# 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8411_9730# VSS.t339 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X778 VDD.t818 CLK.t38 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t1 VDD.t817 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X779 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t54 VDD.t1084 VDD.t1083 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X780 a_9212_739# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t7 a_9412_739# VDD.t2122 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X781 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.CLK.t7 divide_by_2_1.tg_magic_3.IN.t9 VSS.t1101 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X782 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t55 VDD.t1086 VDD.t1085 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X783 VDD.t1088 7b_counter_0.MDFF_4.LD.t56 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VDD.t1087 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X784 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t8 VDD.t1511 VDD.t1510 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X785 VDD.t1090 7b_counter_0.MDFF_4.LD.t57 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1089 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X786 VDD.t133 a_26126_3480# 7b_counter_0.MDFF_7.tspc2_magic_0.D VDD.t129 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X787 a_1409_4557# 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1209_4557# VSS.t232 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X788 VDD.t1337 LD.t35 a_5185_7469# VDD.t1336 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X789 a_1209_6275# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VDD.t727 VDD.t264 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X790 VDD.t92 a_15865_6276# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD.t33 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X791 VDD.t1092 7b_counter_0.MDFF_4.LD.t58 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VDD.t1091 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X792 VDD.t1237 Q1.t12 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t1236 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X793 VDD.t1339 LD.t36 a_1209_3363# VDD.t1338 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X794 a_16065_3363# CLK.t39 VSS.t67 VSS.t66 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X795 VDD.t106 p3_gen_magic_0.xnor_magic_6.OUT a_14556_n8142# VDD.t105 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X796 VSS.t789 D2_2.t12 a_8955_8580# VSS.t788 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X797 VSS.t1046 D2_6.t7 a_8939_n7648# VSS.t1045 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X798 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n5540# VDD.t110 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X799 a_11191_4932# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VDD.t292 VDD.t80 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X800 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t4 CLK.t40 VSS.t65 VSS.t64 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X801 VDD.t816 CLK.t41 DFF_magic_0.tg_magic_3.CLK.t3 VDD.t815 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X802 a_22150_1124# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VSS.t309 VSS.t308 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X803 a_1409_2253# CLK.t42 VSS.t63 VSS.t62 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X804 VDD.t450 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9412_5956# VDD.t448 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X805 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN P2.t9 VDD.t2063 VDD.t2062 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X806 VSS.t543 DFF_magic_0.tg_magic_3.CLK.t11 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS.t542 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X807 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN VDD.t683 VDD.t682 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X808 a_5036_n8095# Q6.t13 VDD.t1440 VDD.t298 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X809 VDD.t603 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8411_4513# VDD.t602 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X810 VDD.t814 CLK.t43 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t3 VDD.t813 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X811 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t8 VDD.t1178 VDD.t1177 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X812 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t37 VDD.t1341 VDD.t1340 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X813 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_0.IN VDD.t502 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X814 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B VSS.t159 VSS.t158 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X815 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t33 VSS.t1003 VSS.t1002 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X816 divide_by_2_0.tg_magic_3.IN.t2 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT divide_by_2_0.tg_magic_1.IN VDD.t144 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X817 VDD.t1721 7b_counter_0.MDFF_5.LD.t34 a_15865_8580# VDD.t1720 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X818 a_12931_8580# CLK.t44 VSS.t61 VSS.t60 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X819 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t12 VDD.t1590 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X820 VDD.t597 a_19152_1223# 7b_counter_0.MDFF_1.QB.t1 VDD.t596 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X821 a_16065_4557# Q2.t12 VSS.t1064 VSS.t1063 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X822 VSS.t1129 D2_7.t8 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS.t1128 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X823 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t38 VDD.t1343 VDD.t1342 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X824 VDD.t948 a_14556_n3644# p2_gen_magic_0.3_inp_AND_magic_0.B VDD.t947 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X825 VDD.t1345 LD.t39 a_5185_2253# VDD.t1344 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X826 VSS.t441 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8955_9774# VSS.t440 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X827 VDD.t1651 7b_counter_0.3_inp_AND_magic_0.C a_23985_7877# VDD.t1649 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X828 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t40 VDD.t1346 VDD.t1325 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X829 OR_magic_2.VOUT.t2 a_23352_n6798# VSS.t452 VSS.t451 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X830 VDD.t1792 D2_1.t14 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD.t1791 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X831 VDD.t828 CLK.t45 a_15865_3363# VDD.t827 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X832 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# VDD.t333 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X833 VSS.t876 Q4.t9 a_1409_1059# VSS.t875 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X834 VSS.t508 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VSS.t507 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X835 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT VDD.t70 pfet_03v3 ad=0.4928p pd=3.12u as=3.0464p ps=18.880001u w=1.12u l=0.56u
X836 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD.t1592 VDD.t1591 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X837 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# VDD.t462 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X838 a_11279_6341# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VSS.t151 VSS.t150 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X839 a_17405_10149# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD.t808 VDD.t806 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X840 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t9 VDD.t2043 VDD.t2042 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X841 VDD.t940 7b_counter_0.MDFF_7.QB.t3 a_27234_4513# VDD.t280 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X842 a_17405_684# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD.t696 VDD.t695 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X843 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.OUT VDD.t737 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X844 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t8 VDD.t1824 VDD.t1823 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X845 VDD.t2083 D2_4.t11 a_23258_1769# VDD.t2082 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X846 a_24259_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t8 a_24059_4877# VDD.t1204 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X847 a_12931_9774# Q1.t13 VSS.t700 VSS.t699 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X848 a_1209_9773# 7b_counter_0.MDFF_3.QB VDD.t65 VDD.t64 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X849 a_1559_n1042# p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t805 VDD.t804 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X850 OR_magic_2.VOUT.t1 a_23352_n6798# VDD.t690 VDD.t688 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X851 VDD.t2129 Q7.t8 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t2128 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X852 a_5036_n7648# p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS.t473 VSS.t472 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X853 a_14756_n3644# p2_gen_magic_0.AND2_magic_1.A a_14556_n3644# VSS.t930 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X854 a_2749_3524# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_4932# VDD.t748 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X855 VDD.t263 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_0.IN VDD.t262 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X856 a_23207_5885# Q2.t13 a_22991_5885# VDD.t1841 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X857 VDD.t1585 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23258_575# VDD.t1584 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X858 a_23560_3728# a_24059_4877# a_24536_3947# VSS.t363 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X859 p3_gen_magic_0.xnor_magic_3.OUT.t0 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n5540# VDD.t561 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X860 divide_by_2_0.tg_magic_3.IN.t6 divide_by_2_0.tg_magic_3.CLK.t9 divide_by_2_0.tg_magic_3.OUT VSS.t862 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X861 VDD.t1794 D2_1.t15 p3_gen_magic_0.inverter_magic_0.VOUT VDD.t1793 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X862 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t13 VDD.t1394 VDD.t1393 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X863 p3_gen_magic_0.P3.t2 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t1485 VDD.t1484 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X864 a_15865_1059# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_16065_1059# VSS.t356 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X865 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t41 VSS.t753 VSS.t752 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X866 a_17405_4932# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD.t41 VDD.t40 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X867 a_12387_5792# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12931_6276# VSS.t1169 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X868 a_2749_10148# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD.t921 VDD.t920 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X869 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t14 VDD.t1239 VDD.t1238 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X870 VSS.t578 a_27567_8496.t11 LD.t2 VSS.t577 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X871 VDD.t1528 Q4.t10 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t1527 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X872 VDD.t997 a_27567_8496.t12 LD.t3 VDD.t996 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X873 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t13 VSS.t1158 VSS.t1157 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X874 VDD.t199 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t6 a_8713_6842# VDD.t198 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X875 VSS.t1210 p2_gen_magic_0.xnor_magic_3.OUT.t4 a_11708_n2115# VSS.t175 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X876 Q7.t1 a_6725_7308# VDD.t781 VDD.t457 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X877 VSS.t830 OR_magic_2.A.t11 DFF_magic_0.tg_magic_2.IN VSS.t829 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X878 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK.t46 VDD.t826 VDD.t825 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X879 VSS.t946 OR_magic_2.VOUT.t10 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VSS.t945 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X880 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# VDD.t111 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X881 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1640 VDD.t280 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X882 a_19307_6886# a_18891_6886# a_19152_6440# VSS.t1278 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X883 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# VDD.t429 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X884 a_4496_4877# 7b_counter_0.MDFF_0.tspc2_magic_0.D VDD.t439 VDD.t438 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X885 VSS.t832 OR_magic_2.A.t12 a_23352_n6798# VSS.t831 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X886 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT divide_by_2_1.tg_magic_0.IN VDD.t390 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X887 VDD.t288 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7215_10149# VDD.t287 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X888 VDD.t1874 p3_gen_magic_0.3_inp_AND_magic_0.C.t4 a_13353_n6613# VDD.t1873 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X889 VDD.t1180 D2_5.t9 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD.t1179 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X890 VSS.t1025 D2_1.t16 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS.t1024 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X891 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t47 VDD.t824 VDD.t823 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X892 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_3524# VDD.t623 VDD.t231 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X893 VDD.t1699 7b_counter_0.MDFF_6.QB.t5 a_15865_6276# VDD.t1698 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X894 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT DFF_magic_0.tg_magic_1.IN VDD.t89 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X895 a_20041_3363# 7b_counter_0.MDFF_4.LD.t59 a_19841_3363# VSS.t612 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X896 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t14 VDD.t1442 VDD.t1441 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X897 7b_counter_0.3_inp_AND_magic_0.A Q4.t11 VSS.t878 VSS.t877 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X898 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t35 VDD.t1723 VDD.t1722 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X899 VDD.t155 7b_counter_0.MDFF_6.tspc2_magic_0.D a_19152_5956# VDD.t154 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X900 a_16065_3363# 7b_counter_0.MDFF_4.LD.t60 a_15865_3363# VSS.t600 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X901 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t12 VDD.t2085 VDD.t2084 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X902 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B VSS.t215 VSS.t214 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X903 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t42 VDD.t1348 VDD.t1347 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X904 VDD.t910 p3_gen_magic_0.xnor_magic_1.OUT.t5 a_16186_n8142# VDD.t909 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X905 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t12 VDD.t960 VDD.t959 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X906 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_3.OUT VSS.t224 VSS.t223 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X907 VDD.t770 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n8579# VDD.t769 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X908 VSS.t572 7b_counter_0.MDFF_4.QB.t7 7b_counter_0.MDFF_4.tspc2_magic_0.Q VSS.t571 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X909 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t1 VDD.t171 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X910 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t11 VDD.t1491 VDD.t1490 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X911 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_8741# VSS.t279 VSS.t216 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X912 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN VDD.t681 VDD.t680 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X913 VDD.t1879 divide_by_2_1.tg_magic_3.CLK.t8 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VDD.t1878 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X914 a_7215_4932# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# VDD.t1 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X915 a_23352_n5390# OR_magic_2.A.t13 VDD.t1465 VDD.t1464 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X916 a_31440_8496.t6 DFF_magic_0.D.t22 VSS.t721 VSS.t720 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X917 a_32816_n1264# mux_magic_0.AND2_magic_0.A a_32616_n1264# VSS.t456 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X918 a_31440_8496.t3 DFF_magic_0.D.t23 VDD.t1278 VDD.t1277 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X919 VDD.t579 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VDD.t578 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X920 a_1541_n7648# p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS.t496 VSS.t495 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X921 VDD.t1600 a_7303_8697# Q2.t1 VDD.t1599 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X922 7b_counter_0.3_inp_AND_magic_0.A Q5.t14 a_23793_5904# VDD.t1991 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X923 VDD.t1529 Q4.t12 a_12174_n8095# VDD.t236 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X924 a_20041_4557# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_19841_4557# VSS.t937 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X925 VSS.t917 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# VSS.t916 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X926 a_16065_4557# 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_15865_4557# VSS.t910 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X927 mux_magic_0.AND2_magic_0.A D2_1.t17 VSS.t1027 VSS.t1026 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X928 VDD.t1222 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11191_10149# VDD.t44 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X929 7b_counter_0.DFF_magic_0.tg_magic_0.IN CLK.t48 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS.t59 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X930 mux_magic_0.OR_magic_0.B a_32616_n2458# VDD.t926 VDD.t925 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X931 a_2749_5900# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_7308# VDD.t404 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X932 VSS.t702 Q1.t15 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VSS.t701 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X933 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.B.t3 VSS.t1180 VSS.t1179 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X934 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_23258_575# VDD.t567 VDD.t566 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X935 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t10 VSS.t666 VSS.t665 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X936 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t61 VDD.t1094 VDD.t1093 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X937 VDD.t761 a_27234_575# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VDD.t760 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X938 VSS.t58 CLK.t49 a_16065_3363# VSS.t57 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X939 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t62 VDD.t1096 VDD.t1095 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X940 a_1209_7469# LD.t43 VDD.t1350 VDD.t1349 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X941 a_32816_n2458# D2_1.t18 a_32616_n2458# VSS.t1028 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X942 VDD.t1531 Q4.t13 a_23793_5904# VDD.t1530 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X943 a_11492_n6613# p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# VSS.t455 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X944 a_8643_n1042# p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t305 VDD.t304 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X945 VDD.t1725 7b_counter_0.MDFF_5.LD.t36 a_12387_8536# VDD.t1724 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X946 a_21504_5904# Q7.t9 7b_counter_0.3_inp_AND_magic_0.B VDD.t2130 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X947 a_24185_7877# 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# VSS.t256 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X948 VDD.t218 VDD.t216 VDD.t218 VDD.t217 pfet_03v3 ad=0.4928p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X949 VDD.t679 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_0.IN VDD.t678 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X950 VDD.t647 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11191_684# VDD.t646 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X951 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD.t502 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X952 VSS.t864 divide_by_2_0.tg_magic_3.CLK.t10 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VSS.t863 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X953 VSS.t668 D2_5.t11 a_12590_n7648# VSS.t667 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X954 VDD.t1846 Q2.t14 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t1845 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X955 VSS.t56 CLK.t50 a_12931_8580# VSS.t55 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X956 a_11492_n6613# p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# VSS.t455 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X957 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t44 VDD.t1352 VDD.t1351 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X958 a_8523_n8095# D2_6.t9 p3_gen_magic_0.xnor_magic_6.OUT VDD.t1620 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X959 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.OUT VDD.t389 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X960 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t45 VSS.t755 VSS.t754 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X961 VSS.t1066 Q2.t15 a_16065_4557# VSS.t1065 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X962 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t46 VSS.t757 VSS.t756 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X963 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t51 VDD.t822 VDD.t821 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X964 7b_counter_0.MDFF_1.QB.t1 a_19152_1223# VDD.t595 VDD.t594 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X965 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t12 VDD.t982 VDD.t981 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X966 a_2749_10148# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_8740# VDD.t17 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X967 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t37 VSS.t1005 VSS.t1004 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X968 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT OR_magic_2.VOUT.t11 VDD.t1653 VDD.t1652 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X969 p2_gen_magic_0.3_inp_AND_magic_0.C.t0 a_16186_n3644# VDD.t166 VDD.t165 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X970 VSS.t317 a_12387_6986# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B VSS.t316 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X971 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK.t52 VDD.t830 VDD.t829 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X972 a_11492_n2115# p2_gen_magic_0.xnor_magic_4.OUT a_11708_n2115# VSS.t175 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X973 a_1209_2253# LD.t47 VDD.t1354 VDD.t1353 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X974 VSS.t504 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_0.IN VSS.t503 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X975 VDD.t675 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26038_4932# VDD.t671 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X976 VDD.t2000 Q5.t15 a_12387_4513# VDD.t48 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X977 a_34156_n2297# mux_magic_0.OR_magic_0.B VSS.t293 VSS.t292 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X978 7b_counter_0.MDFF_0.tspc2_magic_0.D a_2749_3524# VSS.t480 VSS.t210 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X979 a_27234_4513# 7b_counter_0.MDFF_7.QB.t4 VDD.t941 VDD.t280 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X980 DFF_magic_0.tg_magic_2.IN OR_magic_2.A.t14 VDD.t1467 VDD.t1466 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X981 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.NAND_magic_0.VOUT VDD.t731 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X982 VDD.t1796 D2_1.t19 a_32616_n2458# VDD.t1795 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X983 a_5452_n3150# p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT VSS.t194 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X984 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t13 VSS.t1220 VSS.t1219 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X985 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_15865_7470# VDD.t353 VDD.t352 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X986 VDD.t943 7b_counter_0.MDFF_7.QB.t5 7b_counter_0.MDFF_7.tspc2_magic_0.Q VDD.t942 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X987 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_5185_6275# VSS.t450 VSS.t449 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X988 a_23793_5904# Q4.t14 VDD.t1533 VDD.t1532 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X989 VSS.t704 Q1.t16 a_12931_9774# VSS.t703 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X990 p3_gen_magic_0.3_inp_AND_magic_0.B a_14556_n8142# VSS.t326 VSS.t325 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X991 mux_magic_0.OR_magic_0.A a_32616_n1264# VSS.t395 VSS.t394 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X992 VSS.t1246 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VSS.t1245 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X993 VSS.t657 divide_by_2_1.tg_magic_3.IN.t20 mux_magic_0.IN1.t5 VSS.t656 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X994 VSS.t1259 Q7.t10 7b_counter_0.3_inp_AND_magic_0.B VSS.t1258 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X995 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t48 VDD.t1355 VDD.t1347 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X996 VDD.t1535 Q4.t15 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t1534 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X997 VDD.t836 CLK.t53 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t835 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X998 a_12931_2253# D2_6.t10 VSS.t1047 VSS.t17 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X999 Q5.t2 a_6725_2092# VSS.t254 VSS.t253 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1000 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t13 VDD.t2103 VDD.t2102 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1001 a_24536_3947# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t9 VSS.t686 VSS.t685 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1002 a_34156_n2297# mux_magic_0.OR_magic_0.B a_34156_n889# VDD.t399 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1003 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_3.CLK.t13 DFF_magic_0.tg_magic_2.IN VSS.t544 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1004 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_19841_3363# VDD.t375 VDD.t374 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1005 VDD.t670 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8411_9730# VDD.t669 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1006 VSS.t54 CLK.t54 a_27778_2253# VSS.t53 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1007 a_15865_2253# D2_3.t10 VDD.t2045 VDD.t2044 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1008 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_8741# VDD.t370 VDD.t369 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1009 VSS.t723 DFF_magic_0.D.t24 a_27567_8496.t7 VSS.t722 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1010 VDD.t1280 DFF_magic_0.D.t25 a_27567_8496.t4 VDD.t1279 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1011 LD.t4 a_27567_8496.t13 VSS.t580 VSS.t579 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1012 p2_gen_magic_0.xnor_magic_4.OUT D2_3.t11 a_5054_n1526# VDD.t373 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1013 LD.t5 a_27567_8496.t14 VDD.t999 VDD.t998 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1014 a_19841_8580# D2_1.t20 VDD.t1798 VDD.t1797 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1015 a_8713_6842# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t7 VDD.t201 VDD.t200 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1016 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_5185_7469# VSS.t467 VSS.t466 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1017 VSS.t791 D2_2.t14 a_9059_n1973# VSS.t790 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1018 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t9 VDD.t1960 VDD.t1959 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1019 mux_magic_0.OR_magic_0.B a_32616_n2458# VSS.t519 VSS.t518 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1020 VDD.t532 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24259_4877# VDD.t531 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1021 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT CLK.t55 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VSS.t52 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1022 VDD.t2001 Q5.t16 a_8523_n8095# VDD.t598 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1023 a_19307_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK VSS.t389 VSS.t388 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1024 a_5036_n4081# p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t176 VDD.t175 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1025 a_7215_10149# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# VDD.t285 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1026 VDD.t1166 divide_by_2_1.tg_magic_3.IN.t21 mux_magic_0.IN1.t1 VDD.t1165 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1027 p2_gen_magic_0.xnor_magic_5.OUT D2_7.t10 a_5036_n3597# VDD.t108 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1028 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_1.IN VDD.t261 VDD.t260 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1029 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t5 a_13353_n6613# VDD.t479 VDD.t478 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1030 a_23352_n5390# OR_magic_2.A.t15 VDD.t1469 VDD.t1468 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1031 VDD.t834 CLK.t56 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t833 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1032 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t11 VSS.t1049 VSS.t1048 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1033 VSS.t1030 D2_1.t21 p3_gen_magic_0.inverter_magic_0.VOUT VSS.t1029 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1034 divide_by_2_1.tg_magic_2.IN mux_magic_0.IN1.t10 VDD.t1156 VDD.t1155 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1035 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_19841_8580# VSS.t268 VSS.t267 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1036 VDD.t251 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.IN VDD.t250 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1037 VSS.t880 Q4.t16 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VSS.t879 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1038 p2_gen_magic_0.xnor_magic_3.OUT.t1 Q3.t17 a_1559_n1973# VSS.t966 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1039 a_24185_7877# 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# VSS.t256 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1040 a_27778_2253# CLK.t57 VSS.t51 VSS.t50 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1041 VDD.t279 a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD.t278 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1042 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t58 VDD.t832 VDD.t831 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1043 VDD.t47 a_11279_8697# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t1 VDD.t45 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1044 7b_counter_0.DFF_magic_0.tg_magic_1.IN CLK.t59 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS.t49 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1045 OR_magic_2.A.t1 DFF_magic_0.tg_magic_2.OUT VDD.t1211 VDD.t1210 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1046 a_21381_3524# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_4932# VDD.t2169 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1047 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8411_9730# VDD.t490 VDD.t489 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1048 VDD.t1616 a_11279_1124# 7b_counter_0.MDFF_4.tspc2_magic_0.D VDD.t1615 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1049 VSS.t896 OR_magic_1.VOUT.t13 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VSS.t895 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1050 VDD.t1023 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12387_575# VDD.t1022 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1051 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_19841_9774# VSS.t1282 VSS.t1281 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1052 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t12 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VSS.t849 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1053 a_12387_3319# 7b_counter_0.MDFF_4.LD.t63 a_12931_3363# VSS.t607 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1054 a_11191_4932# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# VDD.t76 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1055 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_5900# VDD.t403 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1056 VDD.t2105 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t14 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t2104 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1057 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_8411_3319# VDD.t639 VDD.t638 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1058 7b_counter_0.NAND_magic_0.A.t2 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t954 VDD.t953 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1059 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t10 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS.t1235 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1060 VDD.t74 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VDD.t73 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1061 p2_gen_magic_0.xnor_magic_3.OUT D2_4.t14 a_1559_n1526# VDD.t547 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1062 VDD.t1356 LD.t49 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VDD.t1331 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1063 p3_gen_magic_0.3_inp_AND_magic_0.B a_14556_n8142# VDD.t464 VDD.t463 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1064 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t13 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS.t554 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1065 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.B.t4 VDD.t2033 VDD.t2032 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1066 VSS.t123 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# VSS.t122 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1067 7b_counter_0.MDFF_0.tspc2_magic_0.D a_2749_3524# VDD.t751 VDD.t404 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1068 VDD.t180 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19841_9774# VDD.t179 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1069 a_5185_6275# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5385_6275# VSS.t219 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1070 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t38 VDD.t1727 VDD.t1726 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1071 VDD.t651 p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# VDD.t650 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1072 VDD.t419 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t5 VDD.t418 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1073 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t16 VDD.t2107 VDD.t2106 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1074 VSS.t1160 Q5.t17 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VSS.t1159 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1075 p2_gen_magic_0.AND2_magic_1.A Q4.t17 a_12174_n3150# VSS.t881 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1076 7b_counter_0.3_inp_AND_magic_0.C Q3.t18 a_23207_5885# VDD.t1670 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1077 7b_counter_0.3_inp_AND_magic_0.B Q7.t11 a_21504_5904# VDD.t2131 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1078 a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VDD.t8 VDD.t7 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1079 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.QB.t6 VSS.t978 VSS.t977 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1080 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12931_4557# VSS.t915 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1081 a_21504_5904# Q6.t15 VDD.t1443 VDD.t1438 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1082 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT OR_magic_2.VOUT.t12 VDD.t1655 VDD.t1654 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1083 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t17 VDD.t1241 VDD.t1240 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1084 a_21381_4932# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_3524# VDD.t2168 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1085 a_15865_2253# 7b_counter_0.MDFF_4.LD.t64 VDD.t1098 VDD.t1097 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1086 a_12931_6276# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12387_5792# VSS.t1168 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1087 a_5054_n1042# p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t326 VDD.t325 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1088 VDD.t1728 7b_counter_0.MDFF_5.LD.t39 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t1028 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1089 VDD.t2047 D2_3.t12 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD.t2046 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1090 OR_magic_1.VOUT.t0 a_30365_3514# VDD.t88 VDD.t86 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1091 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.P3.t10 VDD.t1978 VDD.t1977 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1092 a_5185_7469# LD.t50 a_5385_7469# VSS.t758 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1093 a_6725_5900# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD.t187 VDD.t185 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1094 a_1559_n6024# Q3.t19 VDD.t1681 VDD.t1633 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1095 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t51 VSS.t759 VSS.t756 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1096 a_26038_4932# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# VDD.t128 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1097 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN CLK.t60 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS.t48 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1098 a_19152_6440# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK VDD.t2165 VDD.t152 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1099 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t40 VDD.t1729 VDD.t1034 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1100 VDD.t307 p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# VDD.t306 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1101 VDD.t1182 D2_5.t12 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD.t1181 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1102 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t17 VDD.t2109 VDD.t2108 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1103 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT VDD.t151 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1104 VDD.t1099 7b_counter_0.MDFF_4.LD.t65 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD.t1060 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1105 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.NAND_magic_0.A.t11 a_24003_10051# VSS.t732 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1106 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_1.IN VDD.t394 VDD.t393 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1107 divide_by_2_0.tg_magic_3.IN.t11 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_2.IN VDD.t1589 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1108 VDD.t139 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n4081# VDD.t138 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1109 VSS.t1076 p2_gen_magic_0.xnor_magic_1.OUT.t3 a_16386_n3644# VSS.t1075 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1110 VDD.t474 a_26126_1124# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t1 VDD.t189 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1111 VDD.t477 a_22150_1124# Q4.t1 VDD.t475 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1112 a_1541_n8095# Q7.t12 VDD.t2132 VDD.t767 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1113 VDD.t1101 7b_counter_0.MDFF_4.LD.t66 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t1100 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1114 a_20041_3363# D2_3.t13 VSS.t1192 VSS.t1191 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1115 VDD.t97 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_5901# VDD.t37 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1116 a_8523_n3150# p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS.t306 VSS.t305 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1117 a_27234_3319# 7b_counter_0.MDFF_4.LD.t67 a_27778_3363# VSS.t608 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1118 a_12174_n3597# Q4.t18 VDD.t1536 VDD.t140 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1119 DFF_magic_0.D.t4 DFF_magic_0.tg_magic_3.CLK.t14 DFF_magic_0.tg_magic_3.OUT VSS.t545 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1120 VDD.t557 a_27234_3319# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B VDD.t556 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1121 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_12387_575# VDD.t271 VDD.t270 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1122 VDD.t488 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8411_9730# VDD.t487 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1123 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1209_4557# VDD.t385 VDD.t384 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1124 VSS.t1050 D2_6.t12 a_12931_2253# VSS.t2 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1125 VSS.t459 a_23560_3728# a_23672_3947# VSS.t458 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1126 a_12387_6986# 7b_counter_0.MDFF_5.LD.t41 VDD.t1731 VDD.t1730 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1127 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t11 VDD.t1962 VDD.t1961 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1128 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t52 VDD.t1357 VDD.t1351 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1129 VDD.t2049 D2_3.t14 a_19841_3363# VDD.t2048 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1130 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT DFF_magic_0.tg_magic_0.IN VDD.t736 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1131 VDD.t1016 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT P2.t2 VDD.t1015 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1132 a_27778_2253# 7b_counter_0.MDFF_4.LD.t68 a_27234_1769# VSS.t613 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1133 VDD.t1103 7b_counter_0.MDFF_4.LD.t69 a_15865_2253# VDD.t1102 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1134 VSS.t323 a_4496_9609# a_5515_9163# VSS.t322 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1135 a_27567_8496.t6 DFF_magic_0.D.t26 VSS.t725 VSS.t724 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1136 a_23802_2253# 7b_counter_0.MDFF_4.LD.t70 a_23258_1769# VSS.t614 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1137 a_27567_8496.t3 DFF_magic_0.D.t27 VDD.t1282 VDD.t1281 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1138 VSS.t1007 7b_counter_0.MDFF_5.LD.t42 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VSS.t1006 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1139 VDD.t1733 7b_counter_0.MDFF_5.LD.t43 a_19841_8580# VDD.t1732 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1140 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_3.CLK.t9 divide_by_2_1.tg_magic_3.IN.t13 VSS.t1102 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1141 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_5900# VDD.t183 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1142 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_5900# VDD.t402 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1143 a_20041_4557# 7b_counter_0.MDFF_1.tspc2_magic_0.Q VSS.t238 VSS.t237 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1144 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27778_4557# VSS.t936 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1145 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_5185_2253# VSS.t889 VSS.t888 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1146 VDD.t632 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_5900# VDD.t631 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1147 a_23207_5885# Q2.t16 a_22991_5885# VDD.t1841 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1148 a_22991_5885# Q1.t18 VDD.t1242 VDD.t1227 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1149 mux_magic_0.IN1.t0 divide_by_2_1.tg_magic_3.IN.t22 VDD.t1168 VDD.t1167 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1150 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6.t13 VDD.t1826 VDD.t1825 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1151 a_8523_n4081# p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.OUT VDD.t423 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1152 a_11708_n2115# p2_gen_magic_0.xnor_magic_4.OUT a_11492_n2115# VSS.t174 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1153 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t71 VDD.t1105 VDD.t1104 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1154 DFF_magic_0.tg_magic_2.IN OR_magic_2.A.t16 VSS.t834 VSS.t833 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1155 a_4496_10093# 7b_counter_0.MDFF_3.tspc2_magic_0.D VDD.t1604 VDD.t1603 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1156 VSS.t266 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.IN VSS.t265 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1157 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t53 VDD.t1358 VDD.t1340 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1158 a_11191_10149# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# VDD.t44 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1159 a_12387_8536# CLK.t61 VDD.t846 VDD.t845 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1160 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t12 VSS.t1131 VSS.t1130 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1161 VDD.t1632 p2_gen_magic_0.AND2_magic_1.A a_14556_n3644# VDD.t1631 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1162 p2_gen_magic_0.xnor_magic_6.OUT Q5.t18 a_8523_n3150# VSS.t1161 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1163 a_30365_3514# P2.t10 a_30365_4922# VDD.t1473 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1164 p2_gen_magic_0.3_inp_AND_magic_0.A a_11292_n2115# VDD.t741 VDD.t739 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1165 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t72 VDD.t1106 VDD.t1069 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1166 a_9412_739# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t8 a_9212_739# VDD.t2120 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1167 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.P3.t11 VSS.t1145 VSS.t1144 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1168 a_13353_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B VDD.t123 VDD.t121 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1169 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t73 VDD.t1108 VDD.t1107 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1170 7b_counter_0.DFF_magic_0.tg_magic_2.OUT CLK.t62 7b_counter_0.DFF_magic_0.tg_magic_1.IN VSS.t47 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1171 a_34156_n889# mux_magic_0.OR_magic_0.B a_34156_n2297# VDD.t381 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1172 VDD.t1396 D2_2.t15 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD.t1395 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1173 VDD.t1445 Q6.t16 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t1444 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1174 VSS.t898 OR_magic_1.VOUT.t14 divide_by_2_1.inverter_magic_5.VOUT VSS.t897 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1175 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t13 VDD.t1493 VDD.t1492 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1176 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT OR_magic_1.VOUT.t15 VSS.t900 VSS.t899 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1177 LD.t6 a_27567_8496.t15 VDD.t1000 VDD.t994 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1178 VDD.t1734 7b_counter_0.MDFF_5.LD.t44 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t1042 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1179 VDD.t1657 OR_magic_2.VOUT.t13 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VDD.t1656 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1180 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t18 VSS.t1237 VSS.t1236 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1181 VDD.t1735 7b_counter_0.MDFF_5.LD.t45 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t1028 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1182 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VDD.t470 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1183 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_12387_3319# VDD.t191 VDD.t190 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1184 a_8643_n6024# Q1.t19 VDD.t1244 VDD.t1243 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1185 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_1.IN VSS.t289 VSS.t288 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1186 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t20 VDD.t1683 VDD.t1682 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1187 VDD.t1737 7b_counter_0.MDFF_5.LD.t46 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t1736 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1188 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t16 VDD.t2117 VDD.t2116 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1189 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# VDD.t75 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1190 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t14 7b_counter_0.DFF_magic_0.tg_magic_2.IN VSS.t555 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1191 VSS.t520 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_2749_3524# VSS.t212 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1192 7b_counter_0.MDFF_3.QB a_4496_9609# VDD.t461 VDD.t460 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1193 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t47 VDD.t1738 VDD.t1034 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1194 VSS.t557 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t15 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS.t556 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1195 VSS.t230 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_0.IN VSS.t229 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1196 VSS.t539 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.NAND_magic_0.A.t5 VSS.t538 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1197 VDD.t1828 D2_6.t14 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD.t1827 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1198 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_1209_8579# VSS.t180 VSS.t132 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1199 a_5385_6275# 7b_counter_0.MDFF_3.tspc2_magic_0.Q VSS.t143 VSS.t142 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1200 a_19152_739# 7b_counter_0.MDFF_1.tspc2_magic_0.D VDD.t545 VDD.t544 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1201 p3_gen_magic_0.xnor_magic_5.OUT.t1 Q6.t17 a_5036_n7648# VSS.t817 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1202 VDD.t4 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n4081# VDD.t3 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1203 a_20171_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.QB.t0 VSS.t387 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1204 a_11191_10149# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# VDD.t43 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1205 VDD.t120 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12387_9730# VDD.t119 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1206 VDD.t1942 mux_magic_0.IN2.t7 divide_by_2_0.tg_magic_2.IN VDD.t1941 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1207 VDD.t1575 OR_magic_1.VOUT.t16 divide_by_2_1.inverter_magic_5.VOUT VDD.t1574 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1208 VSS.t1086 a_19152_6440# a_20171_6886# VSS.t1085 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1209 VDD.t1740 7b_counter_0.MDFF_5.LD.t48 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VDD.t1739 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1210 divide_by_2_0.tg_magic_0.IN OR_magic_2.VOUT.t14 divide_by_2_0.tg_magic_3.OUT VSS.t947 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1211 a_8523_n3597# Q5.t19 VDD.t2002 VDD.t5 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1212 VSS.t465 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_6725_2092# VSS.t464 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1213 VDD.t844 CLK.t63 a_15865_9774# VDD.t843 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1214 7b_counter_0.MDFF_5.LD.t7 a_29512_8496.t10 VSS.t799 VSS.t798 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1215 7b_counter_0.MDFF_5.LD.t2 a_29512_8496.t11 VDD.t1415 VDD.t1409 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1216 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t15 VSS.t1194 VSS.t1193 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1217 a_5054_n1042# p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_4.OUT VDD.t372 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1218 a_7215_4932# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VDD.t585 VDD.t584 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1219 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26038_684# VDD.t189 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1220 VSS.t234 a_12387_575# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VSS.t233 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1221 VDD.t701 p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# VDD.t699 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1222 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t19 VDD.t1538 VDD.t1537 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1223 VDD.t1246 Q1.t20 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t1245 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1224 a_19152_739# 7b_counter_0.MDFF_1.tspc2_magic_0.D VDD.t543 VDD.t542 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1225 a_5385_7469# D2_7.t13 VSS.t1133 VSS.t1132 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1226 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t3 CLK.t64 VDD.t842 VDD.t841 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1227 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t65 VDD.t840 VDD.t839 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1228 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t66 VSS.t46 VSS.t45 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1229 VDD.t504 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN VDD.t503 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1230 VDD.t1741 7b_counter_0.MDFF_5.LD.t49 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VDD.t1046 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1231 a_5185_2253# LD.t54 a_5385_2253# VSS.t760 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1232 VDD.t1495 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t14 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t1494 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1233 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_1.IN VDD.t259 VDD.t258 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1234 VSS.t416 a_8713_6842# a_8825_6886# VSS.t415 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1235 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t0 a_2749_7308# VDD.t592 VDD.t591 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1236 VSS.t968 Q3.t21 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VSS.t967 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1237 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12387_5792# VDD.t558 VDD.t71 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1238 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t16 VSS.t793 VSS.t792 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1239 divide_by_2_1.tg_magic_3.IN.t0 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT divide_by_2_1.tg_magic_1.IN VDD.t378 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1240 VSS.t1196 D2_3.t16 a_20041_3363# VSS.t1195 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1241 VDD.t1110 7b_counter_0.MDFF_4.LD.t74 a_12387_1769# VDD.t1109 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1242 divide_by_2_1.tg_magic_2.IN mux_magic_0.IN1.t11 VSS.t651 VSS.t650 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1243 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_27234_3319# VDD.t555 VDD.t554 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1244 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VDD.t316 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1245 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t20 VDD.t2004 VDD.t2003 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1246 a_11708_n2115# p2_gen_magic_0.xnor_magic_4.OUT a_11492_n2115# VSS.t174 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1247 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B VSS.t435 VSS.t434 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1248 VDD.t1398 D2_2.t17 a_12387_6986# VDD.t1397 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1249 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B VSS.t497 VSS.t478 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1250 VDD.t1799 D2_1.t22 mux_magic_0.AND2_magic_0.A VDD.t1784 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1251 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t15 VDD.t2087 VDD.t2086 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1252 a_29512_8496.t3 DFF_magic_0.D.t28 VDD.t1283 VDD.t1265 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1253 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t17 VDD.t1848 VDD.t1847 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1254 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n8579# VDD.t734 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1255 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_15865_8580# VSS.t408 VSS.t271 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1256 VDD.t1513 divide_by_2_0.tg_magic_3.CLK.t11 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VDD.t1512 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1257 a_1559_n1042# p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_3.OUT.t0 VDD.t546 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1258 VSS.t236 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_20041_4557# VSS.t235 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1259 VDD.t1743 7b_counter_0.MDFF_5.LD.t50 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1742 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1260 a_1957_n3150# p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT.t1 VSS.t310 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1261 a_21381_3524# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_4932# VDD.t2167 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1262 a_12931_3363# 7b_counter_0.MDFF_4.LD.t75 a_12387_3319# VSS.t611 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1263 VDD.t1744 7b_counter_0.MDFF_5.LD.t51 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD.t1042 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1264 a_14756_n3644# p2_gen_magic_0.xnor_magic_6.OUT VSS.t488 VSS.t487 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1265 VDD.t838 CLK.t67 DFF_magic_0.tg_magic_3.CLK.t2 VDD.t837 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1266 VSS.t490 a_27234_575# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VSS.t489 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1267 a_16065_7470# D2_1.t23 VSS.t1031 VSS.t10 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1268 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t76 VDD.t1112 VDD.t1111 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1269 VDD.t34 a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD.t33 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1270 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t15 VSS.t547 VSS.t546 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1271 7b_counter_0.MDFF_1.tspc2_magic_0.D a_17405_2092# VSS.t366 VSS.t365 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1272 a_21381_8741# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B VSS.t270 VSS.t269 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1273 VDD.t1113 7b_counter_0.MDFF_4.LD.t77 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t1100 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1274 a_2749_4932# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD.t928 VDD.t631 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1275 a_1209_8579# LD.t55 a_1409_8579# VSS.t745 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1276 VDD.t449 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9412_5956# VDD.t448 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1277 a_12174_n8095# D2_5.t13 p3_gen_magic_0.AND2_magic_1.A VDD.t549 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1278 a_23258_575# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23802_1059# VSS.t912 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1279 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t78 VDD.t1114 VDD.t1085 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1280 a_11279_3480# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VSS.t246 VSS.t245 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1281 a_1409_9773# 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1209_9773# VSS.t344 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1282 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_15865_9774# VSS.t110 VSS.t109 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1283 a_16186_n3644# p2_gen_magic_0.xnor_magic_5.OUT VDD.t160 VDD.t159 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1284 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t16 VSS.t549 VSS.t548 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1285 VSS.t835 p2_gen_magic_0.3_inp_AND_magic_0.C.t2 a_13769_n2115# VSS.t172 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1286 VDD.t1115 7b_counter_0.MDFF_4.LD.t79 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD.t1089 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1287 a_2749_4932# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD.t927 VDD.t402 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1288 VDD.t1116 7b_counter_0.MDFF_4.LD.t80 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VDD.t1091 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1289 a_23207_5885# Q2.t18 a_22991_5885# VDD.t1841 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1290 VDD.t2134 Q7.t13 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t2133 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1291 a_12931_4557# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12387_4513# VSS.t914 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1292 a_34156_n2297# mux_magic_0.OR_magic_0.B a_34156_n889# VDD.t400 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1293 VDD.t565 a_23258_575# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VDD.t564 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1294 VDD.t1420 p3_gen_magic_0.xnor_magic_3.OUT.t4 a_11292_n6613# VDD.t1418 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1295 VDD.t1118 7b_counter_0.MDFF_4.LD.t81 a_27234_1769# VDD.t1117 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1296 a_1541_n4081# p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t433 VDD.t432 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1297 a_27567_8496.t2 DFF_magic_0.D.t29 VDD.t1284 VDD.t1267 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1298 VDD.t1987 divide_by_2_0.tg_magic_3.IN.t21 mux_magic_0.IN2.t0 VDD.t1986 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1299 VDD.t1607 a_16186_n8142# p3_gen_magic_0.3_inp_AND_magic_0.C.t0 VDD.t1606 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1300 VSS.t161 p3_gen_magic_0.xnor_magic_6.OUT a_14756_n8142# VSS.t160 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1301 VDD.t1964 D2_7.t14 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD.t1963 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1302 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t15 VDD.t2016 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1303 a_19152_739# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_18891_1669# VDD.t573 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1304 a_11279_6341# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11191_5901# VDD.t77 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1305 VSS.t1068 Q2.t19 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VSS.t1067 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1306 VDD.t496 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1209_9773# VDD.t495 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1307 VSS.t352 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN VSS.t351 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1308 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t52 VSS.t1008 VSS.t1002 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1309 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t16 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS.t558 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1310 VDD.t2119 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t17 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VDD.t2118 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1311 VDD.t1745 7b_counter_0.MDFF_5.LD.t53 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VDD.t1046 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1312 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t14 VDD.t2136 VDD.t2135 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1313 OR_magic_2.A.t4 DFF_magic_0.tg_magic_2.OUT VSS.t690 VSS.t689 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1314 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t17 VSS.t560 VSS.t559 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1315 VSS.t837 p2_gen_magic_0.3_inp_AND_magic_0.C.t3 a_13769_n2115# VSS.t836 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1316 a_32816_n1264# mux_magic_0.IN1.t12 VSS.t653 VSS.t652 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1317 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_1.IN VSS.t228 VSS.t227 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1318 VSS.t1010 7b_counter_0.MDFF_5.LD.t54 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VSS.t1009 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1319 VSS.t734 7b_counter_0.NAND_magic_0.A.t12 7b_counter_0.DFF_magic_0.tg_magic_2.IN VSS.t733 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1320 a_17405_4932# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_3524# VDD.t231 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1321 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t17 VDD.t1612 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1322 VDD.t572 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_1223# VDD.t571 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1323 VSS.t819 Q6.t18 a_1409_6275# VSS.t818 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1324 VDD.t1747 7b_counter_0.MDFF_5.LD.t55 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1746 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1325 7b_counter_0.MDFF_4.LD.t3 a_31440_8496.t14 VSS.t1114 VSS.t1113 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1326 7b_counter_0.MDFF_4.LD.t4 a_31440_8496.t15 VDD.t1929 VDD.t1923 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1327 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.CLK.t12 divide_by_2_0.tg_magic_3.IN.t5 VSS.t865 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1328 7b_counter_0.MDFF_1.QB.t0 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_20171_1669# VSS.t386 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1329 a_8713_1625# a_9212_739# a_9689_1669# VSS.t332 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1330 VDD.t1749 7b_counter_0.MDFF_5.LD.t56 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t1748 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1331 a_5054_n6024# Q2.t20 VDD.t1849 VDD.t22 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1332 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_1209_3363# VSS.t258 VSS.t257 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1333 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t57 VDD.t1750 VDD.t1714 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1334 mux_magic_0.AND2_magic_0.A D2_1.t24 VSS.t1033 VSS.t1032 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1335 VDD.t267 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1209_4557# VDD.t266 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1336 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t58 VDD.t1751 VDD.t1726 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1337 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t18 VDD.t1400 VDD.t1399 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1338 VSS.t801 a_29512_8496.t12 7b_counter_0.MDFF_5.LD.t6 VSS.t800 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1339 VDD.t1416 a_29512_8496.t13 7b_counter_0.MDFF_5.LD.t1 VDD.t1411 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1340 VDD.t454 a_12387_6986# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B VDD.t453 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1341 VDD.t939 7b_counter_0.MDFF_1.QB.t5 a_15865_1059# VDD.t938 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1342 VSS.t902 OR_magic_1.VOUT.t17 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VSS.t901 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1343 VDD.t583 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7215_4932# VDD.t582 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1344 a_4235_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t5 a_4496_4877# VDD.t2023 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1345 VDD.t848 CLK.t68 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t847 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1346 a_5515_9163# a_4496_9609# VSS.t321 VSS.t320 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1347 VDD.t1753 7b_counter_0.MDFF_5.LD.t59 a_8411_8536# VDD.t1752 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1348 VDD.t447 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9412_5956# VDD.t198 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1349 VDD.t1471 OR_magic_2.A.t17 DFF_magic_0.tg_magic_2.IN VDD.t1470 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1350 a_5185_6275# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VDD.t241 VDD.t240 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1351 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t19 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS.t1238 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1352 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t15 VDD.t2138 VDD.t2137 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1353 a_17405_3524# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B VSS.t521 VSS.t158 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1354 a_32816_n2458# mux_magic_0.IN2.t8 VSS.t1121 VSS.t1120 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1355 VSS.t44 CLK.t69 a_1409_7469# VSS.t43 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1356 7b_counter_0.MDFF_6.tspc2_magic_0.D a_17405_7309# VSS.t217 VSS.t216 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1357 a_8643_n1042# p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_0.OUT VDD.t654 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1358 a_15865_8580# 7b_counter_0.MDFF_5.LD.t60 a_16065_8580# VSS.t990 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1359 a_24003_10051# 7b_counter_0.NAND_magic_0.A.t13 7b_counter_0.NAND_magic_0.VOUT VSS.t735 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1360 a_12174_n8579# p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t239 VDD.t238 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1361 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VSS.t169 VSS.t168 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1362 a_5385_2253# D2_5.t14 VSS.t670 VSS.t669 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1363 a_16386_n3644# p2_gen_magic_0.xnor_magic_1.OUT.t4 VSS.t1078 VSS.t1077 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1364 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1209_4557# VSS.t287 VSS.t286 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1365 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t21 VDD.t2006 VDD.t2005 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1366 VDD.t730 a_1209_6275# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD.t386 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1367 a_8825_6886# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t8 7b_counter_0.MDFF_5.QB.t0 VSS.t207 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1368 VSS.t482 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5385_1059# VSS.t481 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1369 a_4651_3947# a_4235_3947# a_4496_4393# VSS.t412 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1370 a_16065_7470# 7b_counter_0.MDFF_5.LD.t61 a_15865_7470# VSS.t1011 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1371 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t70 VSS.t42 VSS.t41 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1372 VDD.t286 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7215_10149# VDD.t285 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1373 VDD.t1850 Q2.t21 a_15865_4557# VDD.t1698 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1374 VDD.t82 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_5901# VDD.t80 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1375 VDD.t1577 OR_magic_1.VOUT.t18 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VDD.t1576 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1376 DFF_magic_0.tg_magic_2.OUT CLK.t71 DFF_magic_0.tg_magic_1.IN VSS.t40 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1377 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t1 a_2749_2092# VDD.t206 VDD.t204 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1378 a_21381_8741# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_10149# VDD.t348 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1379 VSS.t1182 p3_gen_magic_0.xnor_magic_1.B.t5 a_1957_n7648# VSS.t1181 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1380 VSS.t421 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23802_1059# VSS.t420 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1381 a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_16065_9774# VSS.t108 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1382 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t10 VDD.t1881 VDD.t1880 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1383 VDD.t1483 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.P3.t1 VDD.t1482 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1384 a_13553_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B a_13769_n2115# VSS.t172 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1385 VDD.t1479 p2_gen_magic_0.3_inp_AND_magic_0.C.t4 a_13353_n2115# VDD.t1477 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1386 VDD.t2089 D2_4.t16 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD.t2088 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1387 VSS.t437 a_23258_1769# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B VSS.t436 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1388 VDD.t291 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11191_4932# VDD.t80 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1389 VDD.t1944 mux_magic_0.IN2.t9 a_32616_n2458# VDD.t1943 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1390 a_27234_575# Q3.t22 VDD.t1685 VDD.t1684 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1391 VSS.t762 LD.t56 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VSS.t761 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1392 a_14556_n8142# p3_gen_magic_0.AND2_magic_1.A VDD.t551 VDD.t550 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1393 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN CLK.t72 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS.t39 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1394 a_9212_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.D VSS.t315 VSS.t314 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1395 VSS.t1198 D2_3.t17 a_5470_n1973# VSS.t1197 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1396 VDD.t1158 mux_magic_0.IN1.t13 divide_by_2_1.tg_magic_2.IN VDD.t1157 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1397 a_21381_4932# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD.t359 VDD.t358 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1398 VSS.t821 Q6.t19 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VSS.t820 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1399 DFF_magic_0.tg_magic_3.CLK.t1 CLK.t73 VDD.t850 VDD.t849 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1400 a_26038_4932# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VDD.t674 VDD.t671 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1401 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t74 VSS.t38 VSS.t37 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1402 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.QB.t6 VDD.t1868 VDD.t1864 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1403 VDD.t1515 divide_by_2_0.tg_magic_3.CLK.t13 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VDD.t1514 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1404 VDD.t303 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n1042# VDD.t302 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1405 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VDD.t645 VDD.t644 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1406 VSS.t1034 D2_1.t25 a_16065_7470# VSS.t4 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1407 VSS.t1173 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t6 a_4651_3947# VSS.t1172 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1408 VDD.t1295 7b_counter_0.NAND_magic_0.A.t14 DFF_magic_0.D.t8 VDD.t1294 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1409 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT CLK.t75 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t0 VSS.t36 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1410 VDD.t1687 Q3.t23 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t1686 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1411 a_9412_739# 7b_counter_0.MDFF_4.tspc2_magic_0.D VDD.t1628 VDD.t1627 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1412 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t76 VDD.t852 VDD.t851 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1413 VSS.t300 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_21381_8741# VSS.t299 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1414 VDD.t1359 LD.t57 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VDD.t1319 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1415 VSS.t839 p2_gen_magic_0.3_inp_AND_magic_0.C.t5 a_13769_n2115# VSS.t838 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1416 a_1409_8579# D2_7.t15 VSS.t1134 VSS.t71 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1417 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t82 VDD.t1120 VDD.t1119 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1418 7b_counter_0.MDFF_5.LD.t0 a_29512_8496.t14 VDD.t1417 VDD.t1413 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1419 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_1.t26 VDD.t1801 VDD.t1800 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1420 VDD.t1754 7b_counter_0.MDFF_5.LD.t62 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1742 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1421 p3_gen_magic_0.xnor_magic_6.OUT D2_6.t15 a_8523_n8095# VDD.t1621 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1422 a_17405_684# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD.t694 VDD.t693 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1423 a_1209_3363# LD.t58 a_1409_3363# VSS.t748 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1424 VSS.t302 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t7 VSS.t301 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1425 a_17405_684# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD.t692 VDD.t691 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1426 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t83 VDD.t1121 VDD.t1093 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1427 VDD.t1659 OR_magic_2.VOUT.t15 divide_by_2_0.tg_magic_3.CLK.t1 VDD.t1658 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1428 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n2115# VDD.t747 VDD.t745 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1429 a_17405_5901# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD.t96 VDD.t95 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1430 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_5901# VDD.t40 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1431 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t84 VDD.t1122 VDD.t1095 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1432 VDD.t2024 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t7 a_4496_4393# VDD.t441 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1433 a_1209_8579# LD.t59 VDD.t1361 VDD.t1360 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1434 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_1.IN VSS.t502 VSS.t501 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1435 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_15865_2253# VSS.t424 VSS.t275 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1436 a_23352_n5390# p3_gen_magic_0.P3.t12 a_23352_n6798# VDD.t688 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1437 7b_counter_0.3_inp_AND_magic_0.VOUT a_23985_7877# VDD.t2148 VDD.t2147 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1438 a_23258_1769# 7b_counter_0.MDFF_4.LD.t85 VDD.t1124 VDD.t1123 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1439 VDD.t789 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_0.IN VDD.t788 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1440 a_17405_8741# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_10149# VDD.t425 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1441 a_16386_n8142# p3_gen_magic_0.xnor_magic_5.OUT.t3 a_16186_n8142# VSS.t1107 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1442 a_4235_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t8 a_4496_4877# VDD.t2025 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1443 VSS.t262 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# VSS.t146 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1444 a_17405_3524# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_4932# VDD.t40 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1445 a_12174_n3150# p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS.t298 VSS.t297 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1446 a_4496_9609# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t9 VDD.t1198 VDD.t1197 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1447 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.OUT VDD.t195 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1448 p3_gen_magic_0.inverter_magic_0.VOUT D2_1.t27 VDD.t1803 VDD.t1802 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1449 VSS.t1222 D2_4.t17 a_1975_n1973# VSS.t1221 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1450 a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1409_4557# VSS.t231 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1451 a_8523_n8579# p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t601 VDD.t600 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1452 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t15 p2_gen_magic_0.3_inp_AND_magic_0.VOUT VSS.t850 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1453 VDD.t1447 Q6.t20 a_1209_6275# VDD.t1446 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1454 a_8825_6886# a_8713_6842# VSS.t414 VSS.t413 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1455 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t60 VSS.t763 VSS.t754 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1456 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t63 VSS.t1013 VSS.t1012 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1457 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.NAND_magic_0.A.t15 VSS.t737 VSS.t736 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1458 a_23352_n6798# p3_gen_magic_0.P3.t13 a_23352_n5390# VDD.t1468 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1459 a_8411_3319# 7b_counter_0.MDFF_4.LD.t86 a_8955_3363# VSS.t615 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1460 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t64 VSS.t1014 VSS.t1004 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1461 a_5054_n6024# D2_3.t18 p3_gen_magic_0.xnor_magic_4.OUT VDD.t109 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1462 divide_by_2_1.tg_magic_3.IN.t16 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.OUT VDD.t1611 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1463 a_2749_5900# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD.t630 VDD.t629 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1464 a_2749_8740# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_10148# VDD.t16 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1465 a_20171_1669# a_19152_1223# VSS.t402 VSS.t401 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1466 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_3.CLK.t17 DFF_magic_0.tg_magic_2.OUT VSS.t550 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1467 a_9689_1669# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t9 VSS.t1251 VSS.t1250 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1468 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t65 VDD.t1755 VDD.t1722 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1469 a_12387_1769# D2_6.t16 VDD.t1830 VDD.t1829 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1470 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.NAND_magic_0.A.t16 VDD.t1297 VDD.t1296 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1471 7b_counter_0.MDFF_3.tspc2_magic_0.D a_2749_8740# VSS.t114 VSS.t113 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1472 a_1209_3363# LD.t61 VDD.t1363 VDD.t1362 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1473 VDD.t1757 7b_counter_0.MDFF_5.LD.t66 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VDD.t1756 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1474 a_6725_5900# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_7308# VDD.t457 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1475 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t20 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS.t1239 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1476 a_7215_4932# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# VDD.t2 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1477 a_30365_3514# P2.t11 a_30365_4922# VDD.t2064 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1478 a_5036_n8095# D2_7.t16 p3_gen_magic_0.xnor_magic_5.OUT.t0 VDD.t735 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1479 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t22 VDD.t1852 VDD.t1851 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1480 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t0 CLK.t77 VDD.t858 VDD.t857 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1481 7b_counter_0.3_inp_AND_magic_0.C Q3.t24 VSS.t970 VSS.t969 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1482 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_15865_8580# VDD.t609 VDD.t608 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1483 VSS.t35 CLK.t78 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS.t34 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1484 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN CLK.t79 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS.t33 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1485 a_8411_8536# 7b_counter_0.MDFF_5.LD.t67 VDD.t1759 VDD.t1758 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1486 a_9412_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.D VDD.t446 VDD.t200 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1487 divide_by_2_0.tg_magic_3.IN.t1 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT divide_by_2_0.tg_magic_1.IN VDD.t143 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1488 VDD.t1579 OR_magic_1.VOUT.t19 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VDD.t1578 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1489 a_5185_7469# LD.t62 VDD.t1365 VDD.t1364 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1490 VDD.t1125 7b_counter_0.MDFF_4.LD.t87 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD.t1075 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1491 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8955_4557# VSS.t360 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1492 a_12174_n4081# p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.AND2_magic_1.A VDD.t408 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1493 a_21381_8741# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_10149# VDD.t347 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1494 a_5036_n3597# Q6.t21 VDD.t1448 VDD.t175 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1495 VDD.t417 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t4 VDD.t416 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1496 VDD.t1472 OR_magic_2.A.t18 a_23352_n5390# VDD.t1464 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1497 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t88 VDD.t1126 VDD.t1104 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1498 a_1975_n6471# p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT.t1 VSS.t932 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1499 VDD.t290 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11191_4932# VDD.t76 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1500 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t19 VDD.t2051 VDD.t2050 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1501 VSS.t201 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# VSS.t176 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1502 p3_gen_magic_0.inverter_magic_0.VOUT D2_1.t28 VSS.t1036 VSS.t1035 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1503 a_15865_9774# CLK.t80 VDD.t856 VDD.t855 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1504 DFF_magic_0.tg_magic_3.CLK.t0 CLK.t81 VDD.t854 VDD.t853 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1505 VSS.t439 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# VSS.t438 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1506 a_9412_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t9 a_9212_5956# VDD.t202 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1507 VSS.t32 CLK.t82 a_1409_2253# VSS.t31 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1508 VDD.t56 a_1209_7469# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B VDD.t55 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1509 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t18 7b_counter_0.NAND_magic_0.VOUT VSS.t561 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1510 DFF_magic_0.tg_magic_2.OUT CLK.t83 DFF_magic_0.tg_magic_1.IN VSS.t30 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1511 VDD.t482 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1209_1059# VDD.t481 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1512 a_23985_7877# 7b_counter_0.3_inp_AND_magic_0.B VDD.t1638 VDD.t1637 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1513 p3_gen_magic_0.xnor_magic_1.OUT.t1 Q7.t16 a_1541_n7648# VSS.t1260 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1514 a_15865_3363# CLK.t84 VDD.t860 VDD.t859 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1515 divide_by_2_0.tg_magic_3.IN.t13 OR_magic_2.VOUT.t16 divide_by_2_0.tg_magic_1.IN VSS.t948 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1516 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t20 VSS.t883 VSS.t882 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1517 a_1409_1059# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1209_1059# VSS.t336 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1518 a_4496_4393# a_4235_3947# a_4651_3947# VSS.t411 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1519 VDD.t2008 Q5.t22 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t2007 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1520 a_22150_1124# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22062_684# VDD.t475 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1521 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t2 CLK.t85 VDD.t868 VDD.t867 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1522 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT OR_magic_1.VOUT.t20 VDD.t1581 VDD.t1580 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1523 VDD.t866 CLK.t86 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t2 VDD.t865 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1524 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t0 VDD.t170 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1525 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.OUT VDD.t1206 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1526 VSS.t950 OR_magic_2.VOUT.t17 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VSS.t949 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1527 a_21381_10149# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD.t411 VDD.t410 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1528 7b_counter_0.MDFF_4.LD.t5 a_31440_8496.t16 VDD.t1930 VDD.t1925 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1529 VSS.t29 CLK.t87 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS.t28 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1530 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.P3.t14 VDD.t1980 VDD.t1979 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1531 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t616 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1532 a_6725_684# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD.t721 VDD.t660 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1533 a_1559_n6024# D2_4.t18 p3_gen_magic_0.xnor_magic_3.OUT VDD.t560 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1534 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_3.OUT VDD.t340 VDD.t339 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1535 a_5185_2253# LD.t63 VDD.t1367 VDD.t1366 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1536 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN CLK.t88 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS.t27 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1537 a_13353_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B VDD.t122 VDD.t121 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1538 VSS.t324 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# VSS.t122 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1539 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t16 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS.t851 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1540 VSS.t209 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t10 a_9689_6886# VSS.t208 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1541 a_15865_2253# 7b_counter_0.MDFF_4.LD.t89 a_16065_2253# VSS.t599 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1542 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT OR_magic_2.VOUT.t18 VDD.t1661 VDD.t1660 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1543 a_12387_6986# 7b_counter_0.MDFF_5.LD.t68 a_12931_7470# VSS.t981 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1544 VDD.t2159 a_1209_2253# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B VDD.t2158 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1545 a_16065_1059# 7b_counter_0.MDFF_1.QB.t6 VSS.t523 VSS.t522 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1546 VSS.t765 LD.t64 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VSS.t764 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1547 a_1541_n8095# p3_gen_magic_0.xnor_magic_1.B.t6 p3_gen_magic_0.xnor_magic_1.OUT.t0 VDD.t774 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1548 a_30365_4922# P2.t12 a_30365_3514# VDD.t86 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1549 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_19841_4557# VDD.t277 VDD.t276 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1550 VDD.t621 a_8713_6842# 7b_counter_0.MDFF_5.QB.t1 VDD.t620 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1551 VDD.t673 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26038_4932# VDD.t127 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1552 VDD.t1368 LD.t65 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VDD.t1329 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1553 a_19841_9774# 7b_counter_0.MDFF_6.tspc2_magic_0.Q VDD.t178 VDD.t177 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1554 VDD.t1539 Q4.t21 a_23793_5904# VDD.t1530 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1555 DFF_magic_0.D.t7 7b_counter_0.NAND_magic_0.A.t17 VDD.t1299 VDD.t1298 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1556 a_21504_5904# Q7.t17 7b_counter_0.3_inp_AND_magic_0.B VDD.t2130 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1557 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t23 VSS.t1163 VSS.t1162 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1558 VDD.t864 CLK.t89 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t863 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1559 a_19152_5956# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_18891_6886# VDD.t2164 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1560 VSS.t617 7b_counter_0.MDFF_4.LD.t90 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VSS.t616 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1561 VDD.t919 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_2749_10148# VDD.t917 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1562 7b_counter_0.3_inp_AND_magic_0.C Q1.t21 VSS.t706 VSS.t705 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1563 VSS.t552 DFF_magic_0.tg_magic_3.CLK.t18 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS.t551 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1564 a_12931_6276# 7b_counter_0.MDFF_5.QB.t3 VSS.t127 VSS.t126 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1565 VSS.t619 7b_counter_0.MDFF_4.LD.t91 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VSS.t618 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1566 VSS.t853 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t17 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS.t852 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1567 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t92 VSS.t621 VSS.t620 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1568 a_15865_6276# 7b_counter_0.MDFF_6.QB.t7 VDD.t1701 VDD.t1700 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1569 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t4 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t3 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t4 VDD.t208 pfet_03v3 ad=0.4928p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X1570 a_1409_3363# D2_5.t15 VSS.t671 VSS.t62 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1571 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t11 VSS.t1104 VSS.t1103 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1572 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t93 VSS.t623 VSS.t622 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1573 VDD.t324 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n1042# VDD.t323 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1574 7b_counter_0.MDFF_3.tspc2_magic_0.D a_2749_8740# VDD.t19 VDD.t17 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1575 a_19152_6440# a_18891_6886# a_19307_6886# VSS.t1277 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1576 a_8411_8536# D2_2.t19 VDD.t1402 VDD.t1401 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1577 VDD.t1650 7b_counter_0.3_inp_AND_magic_0.C a_23985_7877# VDD.t1649 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1578 VDD.t351 a_15865_7470# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B VDD.t350 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1579 Q3.t2 a_21381_3524# VSS.t1280 VSS.t273 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1580 a_1559_n5540# p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t1634 VDD.t1633 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1581 p3_gen_magic_0.AND2_magic_1.A D2_5.t16 a_12174_n8095# VDD.t548 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1582 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t1 CLK.t90 VDD.t862 VDD.t861 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1583 a_4496_10093# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t10 a_4235_9163# VDD.t1199 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1584 a_19152_5956# 7b_counter_0.MDFF_6.tspc2_magic_0.D VDD.t153 VDD.t152 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1585 DFF_magic_0.tg_magic_0.IN CLK.t91 DFF_magic_0.tg_magic_3.OUT VSS.t26 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1586 a_4496_4877# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t9 a_4235_3947# VDD.t2026 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1587 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t21 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t9 VSS.t1240 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1588 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t1933 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1589 a_23793_5904# Q4.t22 VDD.t1540 VDD.t1532 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1590 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t10 VDD.t1588 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1591 VDD.t1248 Q1.t22 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t1247 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1592 VSS.t261 a_8411_8536# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B VSS.t260 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1593 a_9059_n6471# p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_0.OUT VSS.t1115 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1594 a_29512_8496.t4 DFF_magic_0.D.t30 VSS.t727 VSS.t726 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1595 a_29512_8496.t5 DFF_magic_0.D.t31 VDD.t1285 VDD.t1269 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1596 VDD.t757 p2_gen_magic_0.xnor_magic_6.OUT a_14556_n3644# VDD.t756 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1597 a_1409_4557# 7b_counter_0.MDFF_0.QB.t7 VSS.t1082 VSS.t1081 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1598 VSS.t1052 D2_6.t17 a_8939_n3150# VSS.t1051 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1599 a_1209_6275# Q6.t22 VDD.t1450 VDD.t1449 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1600 VDD.t1541 Q4.t23 a_12174_n3597# VDD.t138 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1601 a_19841_3363# 7b_counter_0.MDFF_4.LD.t94 VDD.t1128 VDD.t1127 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1602 VDD.t720 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_6725_684# VDD.t719 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1603 VDD.t870 CLK.t92 a_1209_7469# VDD.t869 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1604 a_5185_1059# 7b_counter_0.MDFF_0.tspc2_magic_0.Q VDD.t755 VDD.t754 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1605 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t12 VDD.t1883 VDD.t1882 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1606 a_8955_3363# D2_6.t18 VSS.t1054 VSS.t1053 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1607 a_11292_n6613# p3_gen_magic_0.xnor_magic_4.OUT VDD.t1618 VDD.t1617 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1608 VSS.t1204 P2.t13 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VSS.t1203 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1609 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13353_n2115# VDD.t746 VDD.t745 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1610 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t15 VDD.t1610 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1611 a_15865_3363# 7b_counter_0.MDFF_4.LD.t95 VDD.t1130 VDD.t1129 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1612 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# VDD.t188 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1613 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8411_4513# VDD.t577 VDD.t576 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1614 VSS.t708 Q1.t23 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VSS.t707 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1615 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_1.t29 VSS.t1038 VSS.t1037 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1616 a_23985_7877# 7b_counter_0.3_inp_AND_magic_0.A a_24185_7877# VSS.t255 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1617 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t17 VDD.t1184 VDD.t1183 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1618 a_2749_684# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD.t225 VDD.t221 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1619 VDD.t984 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t19 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t983 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1620 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t150 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1621 a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VDD.t494 VDD.t493 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1622 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_5900# VDD.t456 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1623 a_8643_n6024# D2_2.t20 p3_gen_magic_0.xnor_magic_0.OUT VDD.t562 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1624 7b_counter_0.DFF_magic_0.tg_magic_3.OUT CLK.t93 7b_counter_0.DFF_magic_0.tg_magic_0.IN VSS.t25 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1625 VDD.t2091 D2_4.t19 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD.t2090 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1626 a_30365_4922# OR_magic_2.A.t19 VDD.t1474 VDD.t1473 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1627 VSS.t342 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VSS.t341 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1628 VDD.t1404 D2_2.t21 a_8411_8536# VDD.t1403 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1629 a_11292_n6613# p3_gen_magic_0.xnor_magic_0.OUT a_11492_n6613# VSS.t454 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1630 VDD.t1854 Q2.t23 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t1853 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1631 VSS.t625 7b_counter_0.MDFF_4.LD.t96 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VSS.t624 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1632 VDD.t1497 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t18 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t1496 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1633 VDD.t1006 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VDD.t1005 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1634 a_8955_4557# 7b_counter_0.MDFF_4.tspc2_magic_0.Q VSS.t407 VSS.t406 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1635 a_13769_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B a_13553_n6613# VSS.t328 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1636 VSS.t563 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t20 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS.t562 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1637 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3.t20 VDD.t2053 VDD.t2052 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1638 a_23672_3947# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t10 7b_counter_0.MDFF_7.QB.t0 VSS.t687 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1639 VDD.t876 CLK.t94 a_1209_2253# VDD.t875 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1640 p2_gen_magic_0.xnor_magic_6.OUT p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n4081# VDD.t422 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1641 a_16065_1059# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_15865_1059# VSS.t355 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1642 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT CLK.t95 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VSS.t24 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1643 VDD.t51 7b_counter_0.MDFF_5.QB.t4 7b_counter_0.MDFF_5.tspc2_magic_0.Q VDD.t50 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1644 a_11492_n2115# p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# VSS.t251 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1645 a_12387_8536# 7b_counter_0.MDFF_5.LD.t69 VDD.t1761 VDD.t1760 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1646 p3_gen_magic_0.3_inp_AND_magic_0.A a_11292_n6613# VSS.t491 VSS.t454 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1647 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t21 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS.t564 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1648 VSS.t805 p3_gen_magic_0.xnor_magic_3.OUT.t5 a_11708_n6613# VSS.t804 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1649 a_8523_n3597# D2_6.t19 p2_gen_magic_0.xnor_magic_6.OUT VDD.t423 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1650 VDD.t1602 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4496_10093# VDD.t1195 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1651 VDD.t1626 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9412_739# VDD.t1624 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1652 VDD.t1132 7b_counter_0.MDFF_4.LD.t97 a_15865_3363# VDD.t1131 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1653 VDD.t12 a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD.t11 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1654 a_13769_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B a_13553_n6613# VSS.t327 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1655 OUT1.t2 a_34156_n2297# VSS.t285 VSS.t284 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1656 divide_by_2_1.tg_magic_3.IN.t7 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_2.IN VDD.t777 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1657 VDD.t1614 a_11279_1124# 7b_counter_0.MDFF_4.tspc2_magic_0.D VDD.t1613 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1658 a_4651_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t10 VSS.t1175 VSS.t1174 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1659 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_3.OUT VSS.t264 VSS.t263 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1660 DFF_magic_0.D.t6 7b_counter_0.NAND_magic_0.A.t18 VDD.t1301 VDD.t1300 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1661 VDD.t2140 Q7.t18 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t2139 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1662 VDD.t444 a_11279_6341# 7b_counter_0.MDFF_5.tspc2_magic_0.D VDD.t443 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1663 a_5036_n3150# p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS.t165 VSS.t164 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1664 VDD.t530 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24259_4877# VDD.t529 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1665 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t24 VSS.t710 VSS.t709 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1666 VSS.t187 7b_counter_0.MDFF_6.tspc2_magic_0.D a_18891_6886# VSS.t186 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1667 VSS.t627 7b_counter_0.MDFF_4.LD.t98 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VSS.t626 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1668 VDD.t743 p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# VDD.t742 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1669 a_31440_8496.t2 DFF_magic_0.D.t32 VDD.t1286 VDD.t1273 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1670 VDD.t1931 a_31440_8496.t17 7b_counter_0.MDFF_4.LD.t0 VDD.t1927 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1671 VSS.t767 LD.t66 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VSS.t766 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1672 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t23 VDD.t1452 VDD.t1451 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1673 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t96 VDD.t874 VDD.t873 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1674 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2.t22 VDD.t1406 VDD.t1405 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1675 VSS.t769 LD.t67 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VSS.t768 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1676 VSS.t806 p3_gen_magic_0.xnor_magic_3.OUT.t6 a_11708_n6613# VSS.t804 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1677 VDD.t215 VDD.t213 VDD.t215 VDD.t214 pfet_03v3 ad=0.4928p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X1678 a_17405_684# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_2092# VDD.t101 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1679 a_17405_4932# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD.t39 VDD.t37 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1680 VDD.t522 a_15865_1059# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD.t521 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1681 a_15865_6276# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VDD.t29 VDD.t28 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1682 VDD.t1922 p3_gen_magic_0.xnor_magic_5.OUT.t4 a_16186_n8142# VDD.t1921 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1683 VSS.t855 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t19 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS.t854 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1684 VSS.t448 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_0.IN VSS.t447 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1685 VDD.t1543 Q4.t24 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD.t1542 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1686 a_19841_8580# 7b_counter_0.MDFF_5.LD.t70 a_20041_8580# VSS.t1015 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1687 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT OR_magic_2.VOUT.t19 VDD.t1663 VDD.t1662 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1688 p2_gen_magic_0.3_inp_AND_magic_0.B a_14556_n3644# VSS.t535 VSS.t534 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1689 VDD.t338 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.IN VDD.t337 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1690 OUT1.t0 a_34156_n2297# VDD.t382 VDD.t381 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1691 VDD.t1250 Q1.t25 a_8643_n6024# VDD.t1249 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1692 VDD.t282 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VDD.t280 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1693 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t68 VDD.t1370 VDD.t1369 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1694 a_9689_6886# a_9212_5956# a_8713_6842# VSS.t573 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1695 VSS.t510 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_17405_8741# VSS.t156 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1696 VDD.t1805 D2_1.t30 a_15865_7470# VDD.t1804 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1697 VSS.t1056 D2_6.t20 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS.t1055 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1698 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.D.t1 VDD.t228 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1699 a_8643_n5540# p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t1936 VDD.t1243 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1700 VSS.t525 7b_counter_0.MDFF_1.QB.t7 a_16065_1059# VSS.t524 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1701 VDD.t273 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19841_4557# VDD.t272 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1702 VSS.t385 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19307_1669# VSS.t384 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1703 7b_counter_0.MDFF_5.QB.t1 a_8713_6842# VDD.t619 VDD.t618 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1704 VSS.t1151 divide_by_2_0.tg_magic_3.IN.t22 mux_magic_0.IN2.t2 VSS.t1150 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1705 VSS.t23 CLK.t97 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS.t22 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1706 a_4496_4877# 7b_counter_0.MDFF_0.tspc2_magic_0.D VDD.t437 VDD.t436 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1707 VDD.t1689 Q3.t25 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD.t1688 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1708 Q3.t0 a_21381_3524# VDD.t2171 VDD.t2170 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1709 mux_magic_0.IN1.t4 divide_by_2_1.tg_magic_3.IN.t23 VSS.t659 VSS.t658 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1710 a_5036_n4081# p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT VDD.t107 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1711 7b_counter_0.3_inp_AND_magic_0.B Q7.t19 a_21504_5904# VDD.t2131 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1712 VSS.t1200 D2_3.t21 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS.t1199 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1713 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4.t20 VDD.t2093 VDD.t2092 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1714 VDD.t1863 p2_gen_magic_0.xnor_magic_1.OUT.t5 a_16186_n3644# VDD.t1862 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1715 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t118 VDD.t117 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1716 divide_by_2_0.tg_magic_2.IN mux_magic_0.IN2.t10 VDD.t1946 VDD.t1945 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1717 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.QB VDD.t63 VDD.t61 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1718 VDD.t872 CLK.t98 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t871 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1719 divide_by_2_0.tg_magic_3.OUT OR_magic_2.VOUT.t20 divide_by_2_0.tg_magic_0.IN VSS.t951 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1720 a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_20041_9774# VSS.t891 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1721 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t13 VDD.t1885 VDD.t1884 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1722 VDD.t2009 Q5.t24 a_8523_n3597# VDD.t3 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1723 a_23258_575# 7b_counter_0.MDFF_7.tspc2_magic_0.Q VDD.t625 VDD.t624 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1724 a_8955_3363# 7b_counter_0.MDFF_4.LD.t99 a_8411_3319# VSS.t628 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1725 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t69 VDD.t1372 VDD.t1371 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1726 VSS.t129 7b_counter_0.MDFF_5.QB.t5 a_12931_6276# VSS.t128 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1727 VDD.t1209 DFF_magic_0.tg_magic_2.OUT OR_magic_2.A.t0 VDD.t1208 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1728 VDD.t541 7b_counter_0.MDFF_1.tspc2_magic_0.D a_19152_739# VDD.t540 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1729 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t100 VSS.t630 VSS.t629 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1730 DFF_magic_0.tg_magic_3.CLK.t4 CLK.t99 VSS.t21 VSS.t20 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1731 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6.t24 VSS.t823 VSS.t822 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1732 7b_counter_0.MDFF_4.QB.t0 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t10 a_8825_1669# VSS.t1252 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1733 VDD.t27 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_15865_6276# VDD.t26 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1734 VSS.t631 7b_counter_0.MDFF_4.LD.t101 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VSS.t616 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1735 VSS.t517 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_2749_8740# VSS.t422 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1736 a_1541_n3150# p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS.t296 VSS.t295 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1737 VSS.t633 7b_counter_0.MDFF_4.LD.t102 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VSS.t632 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1738 VDD.t1762 7b_counter_0.MDFF_5.LD.t71 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD.t1746 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1739 7b_counter_0.3_inp_AND_magic_0.VOUT a_23985_7877# VSS.t1265 VSS.t255 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1740 a_24259_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.D VDD.t528 VDD.t527 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1741 VDD.t473 a_26126_1124# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t0 VDD.t189 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1742 VDD.t186 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_6725_5900# VDD.t185 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1743 a_27234_575# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t512 VDD.t511 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1744 VDD.t476 a_22150_1124# Q4.t0 VDD.t475 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1745 VDD.t257 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_0.IN VDD.t256 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1746 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t103 VSS.t634 VSS.t622 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1747 VDD.t1221 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11191_10149# VDD.t1220 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1748 VSS.t795 D2_2.t23 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS.t794 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1749 VDD.t328 a_8411_8536# 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B VDD.t327 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1750 VDD.t1453 Q6.t25 a_21504_5904# VDD.t1429 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1751 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t100 VDD.t878 VDD.t877 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1752 VSS.t885 Q4.t25 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VSS.t884 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1753 VDD.t643 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11191_684# VDD.t642 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1754 a_7303_3480# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VSS.t393 VSS.t392 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1755 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK.t101 VDD.t886 VDD.t885 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1756 a_8955_4557# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8411_4513# VSS.t359 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1757 a_8411_9730# 7b_counter_0.MDFF_5.tspc2_magic_0.Q VDD.t668 VDD.t667 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1758 VSS.t1170 a_12387_8536# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B VSS.t316 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1759 a_21381_4932# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD.t357 VDD.t356 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1760 VSS.t729 DFF_magic_0.D.t33 a_29512_8496.t0 VSS.t728 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1761 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_3.OUT VDD.t249 VDD.t248 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1762 VDD.t1287 DFF_magic_0.D.t34 a_29512_8496.t1 VDD.t1271 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1763 VDD.t2011 Q5.t25 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD.t2010 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1764 a_11492_n2115# p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# VSS.t251 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1765 VDD.t1887 divide_by_2_1.tg_magic_3.CLK.t14 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VDD.t1886 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1766 a_1209_7469# CLK.t102 VDD.t884 VDD.t883 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1767 VSS.t1058 D2_6.t21 a_8955_3363# VSS.t1057 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1768 VDD.t168 a_7303_3480# Q6.t0 VDD.t167 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1769 VDD.t1303 7b_counter_0.NAND_magic_0.A.t19 7b_counter_0.NAND_magic_0.VOUT VDD.t1302 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1770 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12387_4513# VDD.t72 VDD.t71 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1771 VDD.t1625 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9412_739# VDD.t1624 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1772 a_1541_n4081# p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT.t0 VDD.t405 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1773 a_24185_7877# 7b_counter_0.3_inp_AND_magic_0.B a_24401_7877# VSS.t933 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1774 VSS.t1224 D2_4.t21 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS.t1223 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1775 VDD.t677 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_0.IN VDD.t676 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1776 VDD.t1875 p3_gen_magic_0.3_inp_AND_magic_0.C.t5 a_13353_n6613# VDD.t1873 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1777 VSS.t673 D2_5.t18 a_12590_n3150# VSS.t672 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1778 VDD.t1856 Q2.t24 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t1855 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1779 a_5470_n6471# p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.OUT VSS.t115 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1780 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT VDD.t149 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1781 VSS.t919 a_7303_8697# Q2.t2 VSS.t918 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1782 a_14556_n8142# p3_gen_magic_0.AND2_magic_1.A a_14756_n8142# VSS.t373 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1783 a_6725_5900# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD.t184 VDD.t183 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1784 a_5036_n8579# p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t299 VDD.t298 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1785 VSS.t694 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VSS.t693 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1786 7b_counter_0.DFF_magic_0.tg_magic_0.IN CLK.t103 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS.t19 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1787 a_12931_3363# CLK.t104 VSS.t18 VSS.t17 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1788 a_2749_5900# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD.t628 VDD.t402 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1789 a_18891_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_5956# VDD.t2163 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1790 VDD.t590 a_32616_n1264# mux_magic_0.OR_magic_0.A VDD.t589 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1791 a_23207_5885# Q2.t25 a_22991_5885# VDD.t1841 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1792 VDD.t952 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.NAND_magic_0.A.t1 VDD.t951 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1793 VSS.t1225 D2_4.t22 a_27778_3363# VSS.t53 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1794 7b_counter_0.3_inp_AND_magic_0.C Q3.t26 a_23207_5885# VDD.t1670 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1795 VSS.t405 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8955_4557# VSS.t404 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1796 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t22 VSS.t566 VSS.t565 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1797 7b_counter_0.MDFF_7.QB.t0 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t11 a_23672_3947# VSS.t688 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1798 VDD.t1134 7b_counter_0.MDFF_4.LD.t104 a_12387_3319# VDD.t1133 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1799 VSS.t635 7b_counter_0.MDFF_4.LD.t105 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VSS.t624 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1800 VDD.t427 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_22062_684# VDD.t426 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1801 a_12931_7470# 7b_counter_0.MDFF_5.LD.t72 a_12387_6986# VSS.t988 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1802 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.D.t0 VDD.t227 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1803 a_1209_2253# CLK.t105 VDD.t882 VDD.t881 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1804 VDD.t1014 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT P2.t1 VDD.t1013 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1805 VSS.t637 7b_counter_0.MDFF_4.LD.t106 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VSS.t636 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1806 a_17405_8741# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_10149# VDD.t424 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1807 a_17405_10149# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD.t807 VDD.t806 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1808 VDD.t880 CLK.t106 a_12387_8536# VDD.t879 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1809 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_684# VDD.t100 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1810 VSS.t16 CLK.t107 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS.t15 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1811 VDD.t1889 divide_by_2_1.tg_magic_3.CLK.t15 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VDD.t1888 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1812 a_12931_4557# Q5.t26 VSS.t1165 VSS.t1164 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1813 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t22 VDD.t2111 VDD.t2110 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1814 a_24259_4877# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t12 a_24059_4877# VDD.t1204 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1815 a_23793_5904# Q5.t27 7b_counter_0.3_inp_AND_magic_0.A VDD.t1990 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1816 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_1.IN VDD.t392 VDD.t391 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1817 VSS.t531 7b_counter_0.MDFF_7.QB.t6 a_27778_4557# VSS.t530 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1818 p2_gen_magic_0.AND2_magic_1.A p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n4081# VDD.t407 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1819 a_1559_n1526# Q3.t27 VDD.t1690 VDD.t804 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1820 divide_by_2_1.tg_magic_2.IN mux_magic_0.IN1.t14 VDD.t1160 VDD.t1159 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1821 a_21381_10149# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD.t409 VDD.t348 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1822 divide_by_2_1.tg_magic_3.IN.t4 OR_magic_1.VOUT.t21 divide_by_2_1.tg_magic_1.IN VSS.t903 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1823 VDD.t1692 Q3.t28 a_27234_575# VDD.t1691 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1824 VDD.t1288 DFF_magic_0.D.t35 a_31440_8496.t1 VDD.t1275 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1825 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t70 VDD.t1373 VDD.t1371 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1826 VDD.t2035 p3_gen_magic_0.xnor_magic_1.B.t7 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD.t2034 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1827 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t71 VSS.t770 VSS.t742 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1828 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t72 VSS.t772 VSS.t771 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1829 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t73 VDD.t1763 VDD.t1085 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1830 a_11279_1124# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11191_684# VDD.t332 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1831 VSS.t638 7b_counter_0.MDFF_4.LD.t107 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VSS.t626 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1832 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_1.IN VSS.t446 VSS.t445 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1833 VDD.t1455 Q6.t26 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD.t1454 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1834 a_12387_575# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12931_1059# VSS.t590 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1835 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_15865_2253# VDD.t635 VDD.t634 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1836 VSS.t773 LD.t73 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VSS.t768 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1837 a_27778_3363# D2_4.t23 VSS.t1226 VSS.t50 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1838 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t17 VDD.t1966 VDD.t1965 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1839 a_2749_10148# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD.t918 VDD.t917 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1840 a_1541_n3597# Q7.t20 VDD.t2141 VDD.t432 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1841 VDD.t2123 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t11 a_8713_1625# VDD.t1622 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1842 a_2749_3524# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B VSS.t479 VSS.t478 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1843 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27234_4513# VDD.t281 VDD.t280 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1844 VSS.t953 OR_magic_2.VOUT.t21 divide_by_2_0.tg_magic_3.CLK.t1 VSS.t952 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1845 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2.t26 VSS.t1070 VSS.t1069 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1846 VDD.t1623 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9412_739# VDD.t1622 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1847 Q7.t0 a_6725_7308# VDD.t780 VDD.t779 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1848 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.IN VDD.t1205 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1849 VDD.t962 DFF_magic_0.tg_magic_3.CLK.t19 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t961 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1850 a_12387_9730# Q1.t26 VDD.t1252 VDD.t1251 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1851 a_19307_1669# a_18891_1669# a_19152_1223# VSS.t397 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1852 VDD.t581 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7215_4932# VDD.t580 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1853 a_2749_684# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD.t224 VDD.t223 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1854 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_684# VDD.t99 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1855 VDD.t2014 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12387_5792# VDD.t1593 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1856 VDD.t1857 Q2.t27 a_5054_n6024# VDD.t24 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1857 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_15865_1059# VDD.t520 VDD.t519 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1858 a_27778_4557# 7b_counter_0.MDFF_7.QB.t7 VSS.t533 VSS.t532 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1859 a_19841_3363# D2_3.t22 VDD.t2055 VDD.t2054 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1860 P2.t0 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t1012 VDD.t1011 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1861 VDD.t1136 7b_counter_0.MDFF_4.LD.t108 a_27234_3319# VDD.t1135 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1862 a_14556_n8142# p3_gen_magic_0.xnor_magic_6.OUT VDD.t104 VDD.t103 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1863 a_5054_n5540# p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD.t23 VDD.t22 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1864 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.OUT VDD.t388 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1865 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_3524# VSS.t417 VSS.t365 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1866 a_22991_5885# Q1.t27 VDD.t1253 VDD.t1227 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1867 VSS.t942 7b_counter_0.3_inp_AND_magic_0.C a_24401_7877# VSS.t933 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1868 a_16186_n8142# p3_gen_magic_0.xnor_magic_5.OUT.t5 a_16386_n8142# VSS.t1108 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1869 VDD.t1456 Q6.t27 a_5036_n8095# VDD.t300 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1870 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.A VDD.t214 pfet_03v3 ad=0.4928p pd=3.12u as=1.9712p ps=12.48u w=1.12u l=0.56u
X1871 VSS.t640 7b_counter_0.MDFF_4.LD.t109 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VSS.t639 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1872 VSS.t641 7b_counter_0.MDFF_4.LD.t110 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VSS.t632 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1873 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n1042# VDD.t653 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1874 VDD.t344 a_19841_8580# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B VDD.t343 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1875 VDD.t1598 a_7303_8697# Q2.t0 VDD.t1595 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1876 VDD.t1764 7b_counter_0.MDFF_5.LD.t74 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t1736 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1877 VDD.t237 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n8579# VDD.t236 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1878 VSS.t105 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# VSS.t104 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1879 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7.t18 VSS.t1136 VSS.t1135 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1880 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t711 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1881 p2_gen_magic_0.3_inp_AND_magic_0.B a_14556_n3644# VDD.t946 VDD.t945 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1882 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_1.t31 VDD.t1807 VDD.t1806 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1883 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS.t506 VSS.t505 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1884 VDD.t355 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_21381_4932# VDD.t354 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1885 a_27234_575# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27778_1059# VSS.t353 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1886 7b_counter_0.MDFF_0.QB.t0 a_4496_4393# VDD.t146 VDD.t145 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1887 VDD.t212 VDD.t210 VDD.t212 VDD.t211 pfet_03v3 ad=0.4928p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X1888 VDD.t2057 D2_3.t23 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD.t2056 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1889 VDD.t2020 a_12387_8536# 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B VDD.t2019 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1890 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VDD.t615 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1891 VDD.t78 a_11279_3480# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t0 VDD.t77 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1892 a_30365_4922# OR_magic_2.A.t20 VDD.t1475 VDD.t1457 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1893 a_5054_n6471# p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS.t167 VSS.t166 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1894 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t801 VDD.t800 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1895 a_8643_n1526# Q1.t28 VDD.t1254 VDD.t304 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1896 p3_gen_magic_0.P3.t0 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD.t1481 VDD.t1480 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1897 VDD.t803 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n1042# VDD.t802 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1898 divide_by_2_1.inverter_magic_5.VOUT OR_magic_1.VOUT.t22 VSS.t905 VSS.t904 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1899 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1209_9773# VSS.t516 VSS.t515 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1900 VDD.t1499 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t20 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t1498 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1901 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1.t29 VDD.t1256 VDD.t1255 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1902 VSS.t125 a_11279_8697# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t2 VSS.t124 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1903 VSS.t1138 D2_7.t19 a_5452_n7648# VSS.t1137 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1904 VSS.t1262 Q7.t21 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VSS.t1261 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1905 VDD.t1001 a_27567_8496.t16 LD.t7 VDD.t996 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1906 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t1643 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1907 VSS.t141 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5385_6275# VSS.t140 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1908 VSS.t3 CLK.t108 a_12931_3363# VSS.t2 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1909 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t75 VDD.t1765 VDD.t1085 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1910 mux_magic_0.OR_magic_0.A a_32616_n1264# VDD.t588 VDD.t587 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1911 7b_counter_0.NAND_magic_0.A.t0 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD.t950 VDD.t949 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1912 p3_gen_magic_0.inverter_magic_0.VOUT D2_1.t32 VDD.t1809 VDD.t1808 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1913 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VDD.t1004 VDD.t1003 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1914 VDD.t1408 D2_2.t24 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD.t1407 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1915 VDD.t2059 D2_3.t24 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD.t2058 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1916 a_27778_3363# 7b_counter_0.MDFF_4.LD.t111 a_27234_3319# VSS.t613 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1917 a_8523_n8579# p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.OUT VDD.t1620 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1918 VDD.t993 7b_counter_0.MDFF_4.QB.t8 7b_counter_0.MDFF_4.tspc2_magic_0.Q VDD.t991 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1919 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t8 VDD.t1642 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1920 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t26 VDD.t1545 VDD.t1544 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1921 OR_magic_2.VOUT.t0 a_23352_n6798# VDD.t689 VDD.t688 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1922 VDD.t2070 p2_gen_magic_0.xnor_magic_3.OUT.t5 a_11292_n2115# VDD.t2069 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1923 VSS.t500 a_12387_1769# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B VSS.t202 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1924 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t112 VDD.t1137 VDD.t1083 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1925 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t14 VDD.t1517 VDD.t1516 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1926 a_18891_1669# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_739# VDD.t570 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1927 7b_counter_0.NAND_magic_0.A.t4 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS.t537 VSS.t536 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1928 VDD.t1186 D2_5.t19 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD.t1185 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1929 a_2749_3524# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_4932# VDD.t402 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1930 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3.t29 VDD.t1694 VDD.t1693 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1931 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t113 VSS.t643 VSS.t642 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1932 VSS.t941 7b_counter_0.3_inp_AND_magic_0.C a_24401_7877# VSS.t939 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1933 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT OR_magic_2.VOUT.t22 VSS.t955 VSS.t954 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1934 VDD.t2071 p2_gen_magic_0.xnor_magic_3.OUT.t6 a_11292_n2115# VDD.t2069 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1935 VDD.t986 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t23 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD.t985 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1936 p3_gen_magic_0.3_inp_AND_magic_0.A a_11292_n6613# VDD.t765 VDD.t764 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1937 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t20 VDD.t964 VDD.t963 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1938 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_684# VDD.t659 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1939 VSS.t1140 D2_7.t20 a_5385_7469# VSS.t1139 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1940 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_5185_1059# VDD.t714 VDD.t713 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1941 VSS.t1167 Q5.t28 a_12931_4557# VSS.t1166 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1942 7b_counter_0.MDFF_6.tspc2_magic_0.D a_17405_7309# VDD.t233 VDD.t231 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1943 a_13353_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B VDD.t468 VDD.t467 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1944 a_26126_3480# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VSS.t444 VSS.t168 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1945 VDD.t944 7b_counter_0.MDFF_7.QB.t8 7b_counter_0.MDFF_7.tspc2_magic_0.Q VDD.t942 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1946 VDD.t799 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VDD.t798 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1947 VDD.t895 CLK.t109 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t894 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1948 a_27778_4557# 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27234_4513# VSS.t935 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1949 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_5901# VDD.t230 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1950 divide_by_2_1.tg_magic_1.IN OR_magic_1.VOUT.t23 divide_by_2_1.tg_magic_3.IN.t3 VSS.t906 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1951 a_31440_8496.t0 DFF_magic_0.D.t36 VDD.t1289 VDD.t1277 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1952 a_18891_6886# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_5956# VDD.t2162 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1953 a_16186_n8142# p3_gen_magic_0.xnor_magic_1.OUT.t6 VDD.t912 VDD.t911 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1954 a_34156_n2297# mux_magic_0.OR_magic_0.B a_34156_n889# VDD.t399 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1955 a_4496_10093# 7b_counter_0.MDFF_3.tspc2_magic_0.D VDD.t1601 VDD.t1197 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1956 a_1559_n6471# p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS.t379 VSS.t378 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1957 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VDD.t1932 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1958 VSS.t972 Q3.t30 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VSS.t971 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1959 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD.t74 VDD.t1374 VDD.t1310 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1960 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t75 VSS.t774 VSS.t771 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1961 VDD.t132 a_26126_3480# 7b_counter_0.MDFF_7.tspc2_magic_0.D VDD.t131 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1962 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t76 VDD.t1376 VDD.t1375 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1963 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_3524# VDD.t622 VDD.t231 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1964 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t76 VDD.t1766 VDD.t1095 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1965 VDD.t2151 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.IN VDD.t2150 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1966 a_8713_1625# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t12 VDD.t2124 VDD.t1627 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1967 VDD.t687 a_5185_6275# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD.t686 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1968 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_3.CLK.t16 divide_by_2_1.tg_magic_3.IN.t12 VSS.t1105 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1969 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t21 VDD.t966 VDD.t965 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1970 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.QB.t8 VDD.t1702 VDD.t1696 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1971 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t2 a_2749_7308# VSS.t396 VSS.t113 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1972 VDD.t599 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n8579# VDD.t598 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1973 p2_gen_magic_0.3_inp_AND_magic_0.A a_11292_n2115# VDD.t740 VDD.t739 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1974 VDD.t1519 divide_by_2_0.tg_magic_3.CLK.t15 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VDD.t1518 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1975 a_7215_4932# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# VDD.t1 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1976 a_23352_n5390# OR_magic_2.A.t21 VDD.t1476 VDD.t1464 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1977 a_12387_1769# 7b_counter_0.MDFF_4.LD.t114 VDD.t1139 VDD.t1138 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1978 Q5.t0 a_6725_2092# VDD.t310 VDD.t309 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1979 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_3.OUT VDD.t336 VDD.t335 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1980 VDD.t893 CLK.t110 a_27234_1769# VDD.t892 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1981 a_5054_n5540# p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.OUT VDD.t109 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1982 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_19841_3363# VSS.t283 VSS.t282 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1983 VDD.t1141 7b_counter_0.MDFF_4.LD.t115 a_19841_3363# VDD.t1140 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1984 VSS.t248 a_27234_1769# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B VSS.t247 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1985 VDD.t2066 P2.t14 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VDD.t2065 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1986 VDD.t1305 7b_counter_0.NAND_magic_0.A.t20 7b_counter_0.DFF_magic_0.tg_magic_2.IN VDD.t1304 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1987 a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1409_9773# VSS.t343 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1988 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN.t0 VDD.t142 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1989 a_23258_1769# 7b_counter_0.MDFF_4.LD.t116 a_23802_2253# VSS.t644 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1990 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.CLK.t16 VSS.t867 VSS.t866 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1991 VDD.t1948 mux_magic_0.IN2.t11 divide_by_2_0.tg_magic_2.IN VDD.t1947 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1992 7b_counter_0.DFF_magic_0.tg_magic_2.OUT CLK.t111 7b_counter_0.DFF_magic_0.tg_magic_1.IN VSS.t14 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1993 VDD.t46 a_11279_8697# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t0 VDD.t45 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1994 a_12590_n7648# p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.AND2_magic_1.A VSS.t218 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1995 VDD.t222 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_2749_684# VDD.t221 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1996 a_1209_1059# Q4.t27 VDD.t1547 VDD.t1546 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X1997 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t0 a_2749_2092# VDD.t205 VDD.t204 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1998 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t23 VSS.t1242 VSS.t1241 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X1999 a_12174_n3597# D2_5.t20 p2_gen_magic_0.AND2_magic_1.A VDD.t408 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2000 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# VDD.t666 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2001 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_19841_4557# VSS.t240 VSS.t239 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2002 mux_magic_0.AND2_magic_0.A D2_1.t33 VDD.t1810 VDD.t1778 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2003 VDD.t753 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5185_1059# VDD.t752 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2004 VDD.t1665 OR_magic_2.VOUT.t23 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VDD.t1664 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2005 a_2749_8740# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_10148# VDD.t15 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2006 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN VDD.t710 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2007 VDD.t1142 7b_counter_0.MDFF_4.LD.t117 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD.t1066 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2008 a_12387_3319# CLK.t112 VDD.t891 VDD.t890 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2009 VDD.t1989 divide_by_2_0.tg_magic_3.IN.t23 mux_magic_0.IN2.t1 VDD.t1988 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2010 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VDD.t1021 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2011 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VDD.t81 VDD.t80 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2012 a_9412_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t11 a_9212_5956# VDD.t202 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2013 a_27234_1769# 7b_counter_0.MDFF_4.LD.t118 VDD.t1144 VDD.t1143 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2014 a_4651_9163# a_4235_9163# a_4496_9609# VSS.t338 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2015 Q1.t0 a_21381_8741# VDD.t771 VDD.t349 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2016 VDD.t1832 D2_6.t22 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD.t1831 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2017 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.QB.t8 VSS.t1084 VSS.t1083 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2018 VSS.t940 7b_counter_0.3_inp_AND_magic_0.C a_24401_7877# VSS.t939 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2019 a_23802_1059# 7b_counter_0.MDFF_7.tspc2_magic_0.Q VSS.t419 VSS.t418 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2020 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.QB VDD.t62 VDD.t61 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2021 VSS.t410 mux_magic_0.OR_magic_0.A a_34156_n2297# VSS.t409 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2022 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t1 CLK.t113 VDD.t889 VDD.t888 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2023 a_32616_n2458# D2_1.t34 VDD.t1812 VDD.t1811 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2024 VSS.t147 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# VSS.t146 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2025 VDD.t60 7b_counter_0.MDFF_3.QB a_1209_9773# VDD.t59 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2026 p2_gen_magic_0.xnor_magic_5.OUT Q6.t28 a_5036_n3150# VSS.t824 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2027 VSS.t486 p2_gen_magic_0.xnor_magic_6.OUT a_14756_n3644# VSS.t485 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2028 VDD.t797 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VDD.t796 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2029 a_34156_n889# mux_magic_0.OR_magic_0.A VDD.t613 VDD.t399 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2030 VSS.t1072 Q2.t28 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VSS.t1071 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2031 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.QB.t8 VSS.t527 VSS.t526 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2032 VDD.t672 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26038_4932# VDD.t671 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2033 a_1559_n5540# p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT.t0 VDD.t560 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2034 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t21 VDD.t1501 VDD.t1500 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2035 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.CLK.t17 divide_by_2_0.tg_magic_3.IN.t4 VSS.t868 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2036 VDD.t1290 DFF_magic_0.D.t37 a_27567_8496.t1 VDD.t1279 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2037 LD.t8 a_27567_8496.t17 VDD.t1002 VDD.t998 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2038 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t28 VDD.t1549 VDD.t1548 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2039 VSS.t13 CLK.t114 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t4 VSS.t12 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2040 a_1409_6275# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1209_6275# VSS.t468 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2041 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_15865_6276# VSS.t155 VSS.t154 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2042 VDD.t1258 Q1.t30 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD.t1257 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2043 a_8643_n6471# p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS.t381 VSS.t380 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2044 a_34156_n889# mux_magic_0.OR_magic_0.A VDD.t612 VDD.t610 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2045 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t77 VDD.t1378 VDD.t1377 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2046 a_12931_1059# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12387_575# VSS.t589 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2047 VDD.t135 a_1209_8579# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B VDD.t134 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2048 p3_gen_magic_0.xnor_magic_1.OUT.t0 p3_gen_magic_0.xnor_magic_1.B.t8 a_1541_n8095# VDD.t773 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2049 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD.t78 VDD.t1380 VDD.t1379 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2050 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS.t350 VSS.t349 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2051 VDD.t69 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5185_6275# VDD.t68 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2052 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t77 VDD.t1767 VDD.t1095 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2053 a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VDD.t265 VDD.t264 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2054 a_5054_n1526# Q2.t29 VDD.t1858 VDD.t325 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2055 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_12387_6986# VDD.t452 VDD.t451 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2056 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.CLK.t22 VDD.t968 VDD.t967 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2057 a_6725_5900# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD.t182 VDD.t181 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2058 VDD.t1968 D2_7.t21 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD.t1967 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2059 VDD.t887 CLK.t115 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD.t502 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2060 a_19152_1223# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK VDD.t569 VDD.t568 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2061 VSS.t682 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t11 a_4651_9163# VSS.t681 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2062 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t78 VDD.t1769 VDD.t1768 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2063 VDD.t174 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n4081# VDD.t173 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2064 OR_magic_1.VOUT.t1 a_30365_3514# VSS.t153 VSS.t152 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2065 a_24003_10051# 7b_counter_0.3_inp_AND_magic_0.VOUT VSS.t346 VSS.t345 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2066 VDD.t1770 7b_counter_0.MDFF_5.LD.t79 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t1748 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2067 VDD.t1771 7b_counter_0.MDFF_5.LD.t80 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VDD.t1739 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2068 VSS.t177 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# VSS.t176 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2069 a_1409_7469# LD.t79 a_1209_7469# VSS.t747 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2070 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5.t29 VDD.t2013 VDD.t2012 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2071 VDD.t970 DFF_magic_0.tg_magic_3.CLK.t23 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t969 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2072 a_16065_8580# CLK.t116 VSS.t11 VSS.t10 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2073 a_12387_5792# 7b_counter_0.MDFF_5.QB.t6 VDD.t53 VDD.t52 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2074 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT OR_magic_1.VOUT.t24 VSS.t908 VSS.t907 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2075 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_1.IN VDD.t787 VDD.t786 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2076 VSS.t675 D2_5.t21 a_5385_2253# VSS.t674 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2077 a_17405_5901# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD.t94 VDD.t40 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2078 a_1541_n8579# p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t768 VDD.t767 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2079 VDD.t1503 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t22 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t1502 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2080 VDD.t320 a_1209_3363# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B VDD.t319 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2081 a_13353_n6613# p3_gen_magic_0.3_inp_AND_magic_0.A a_13553_n6613# VSS.t328 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2082 VDD.t1834 D2_6.t23 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD.t1833 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2083 VSS.t655 mux_magic_0.IN1.t15 a_32816_n1264# VSS.t654 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2084 a_15865_4557# Q2.t30 VDD.t1859 VDD.t1700 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2085 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VDD.t1020 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2086 VSS.t453 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_17405_2092# VSS.t120 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2087 VSS.t1228 D2_4.t24 a_23802_2253# VSS.t1227 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2088 VSS.t646 7b_counter_0.MDFF_4.LD.t119 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VSS.t645 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2089 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_5185_6275# VDD.t685 VDD.t684 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2090 VDD.t269 a_12387_575# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VDD.t268 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2091 a_4235_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t12 a_4496_10093# VDD.t1194 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2092 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 a_13353_n6613# VSS.t334 VSS.t327 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2093 VDD.t726 a_5185_7469# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B VDD.t725 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2094 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1209_6275# VDD.t729 VDD.t384 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2095 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_5900# VDD.t455 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2096 p3_gen_magic_0.xnor_magic_0.OUT Q1.t31 a_8643_n6471# VSS.t711 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2097 VDD.t924 a_32616_n2458# mux_magic_0.OR_magic_0.B VDD.t923 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2098 a_5385_1059# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5185_1059# VSS.t277 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2099 a_16065_9774# CLK.t117 VSS.t9 VSS.t8 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2100 VDD.t1870 a_19152_6440# 7b_counter_0.MDFF_6.QB.t0 VDD.t1869 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2101 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_5900# VDD.t401 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2102 a_8939_n7648# p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_6.OUT VSS.t403 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2103 VDD.t112 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_26038_684# VDD.t111 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2104 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# VDD.t76 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2105 a_19152_739# 7b_counter_0.MDFF_1.tspc2_magic_0.D VDD.t539 VDD.t538 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2106 VDD.t1836 D2_6.t24 a_12387_1769# VDD.t1835 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2107 VDD.t700 p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# VDD.t699 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2108 VSS.t1147 p3_gen_magic_0.P3.t15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VSS.t1146 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2109 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_3.CLK.t18 divide_by_2_0.tg_magic_3.IN.t7 VSS.t869 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2110 VDD.t2068 P2.t15 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VDD.t2067 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2111 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t80 VDD.t1381 VDD.t1342 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2112 VSS.t1123 mux_magic_0.IN2.t12 a_32816_n2458# VSS.t1122 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2113 a_27234_1769# CLK.t118 VDD.t904 VDD.t903 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2114 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_1209_1059# VSS.t222 VSS.t221 nfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2115 a_5515_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t11 7b_counter_0.MDFF_0.QB.t1 VSS.t1176 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2116 a_23258_1769# D2_4.t25 VDD.t2095 VDD.t2094 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2117 VSS.t7 CLK.t119 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS.t6 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2118 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t120 VDD.t1146 VDD.t1145 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2119 VDD.t607 a_15865_8580# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B VDD.t606 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2120 p3_gen_magic_0.xnor_magic_0.OUT D2_2.t25 a_8643_n6024# VDD.t563 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2121 VSS.t826 Q6.t29 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VSS.t825 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2122 a_11191_4932# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# VDD.t76 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2123 VDD.t1772 7b_counter_0.MDFF_5.LD.t81 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VDD.t1756 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2124 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD.t415 VDD.t414 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2125 VDD.t2143 Q7.t22 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD.t2142 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2126 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD.t81 VSS.t776 VSS.t775 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2127 a_8643_n5540# p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.OUT VDD.t562 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2128 a_1409_9773# 7b_counter_0.MDFF_3.QB VSS.t135 VSS.t134 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2129 VDD.t1551 a_5185_2253# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B VDD.t1550 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2130 VDD.t38 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_17405_4932# VDD.t37 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2131 a_13553_n6613# p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# VSS.t328 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2132 a_15865_6276# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_16065_6276# VSS.t116 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2133 VDD.t1667 OR_magic_2.VOUT.t24 divide_by_2_0.tg_magic_3.CLK.t0 VDD.t1666 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2134 VSS.t739 7b_counter_0.NAND_magic_0.A.t21 DFF_magic_0.D.t10 VSS.t738 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2135 VDD.t209 VDD.t207 VDD.t209 VDD.t208 pfet_03v3 ad=0.4928p pd=3.12u as=0 ps=0 w=1.12u l=0.56u
X2136 VDD.t1970 D2_7.t22 a_1209_8579# VDD.t1969 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2137 VDD.t164 a_16186_n3644# p2_gen_magic_0.3_inp_AND_magic_0.C.t0 VDD.t163 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2138 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN.t6 VDD.t776 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2139 divide_by_2_1.tg_magic_0.IN OR_magic_1.VOUT.t25 divide_by_2_1.tg_magic_3.OUT VSS.t909 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2140 a_30365_3514# P2.t16 VSS.t1206 VSS.t1205 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2141 VDD.t902 CLK.t120 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD.t901 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2142 VDD.t900 CLK.t121 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD.t899 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2143 p2_gen_magic_0.xnor_magic_6.OUT D2_6.t25 a_8523_n3597# VDD.t422 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2144 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD.t1019 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2145 a_13553_n6613# p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# VSS.t327 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2146 VDD.t54 7b_counter_0.MDFF_5.QB.t7 7b_counter_0.MDFF_5.tspc2_magic_0.Q VDD.t50 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2147 a_4496_4393# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t12 VDD.t2027 VDD.t438 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2148 VSS.t1141 D2_7.t23 a_1409_8579# VSS.t43 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2149 VDD.t1695 Q3.t31 a_1559_n6024# VDD.t1635 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2150 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t23 VDD.t2145 VDD.t2144 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2151 VDD.t284 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7215_10149# VDD.t283 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2152 a_9212_5956# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t12 a_9412_5956# VDD.t203 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2153 a_4496_9609# a_4235_9163# a_4651_9163# VSS.t337 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2154 VDD.t459 a_4496_9609# 7b_counter_0.MDFF_3.QB VDD.t458 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2155 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.LD.t121 VSS.t647 VSS.t597 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2156 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5.t22 VDD.t1188 VDD.t1187 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2157 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.OUT VDD.t194 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2158 VSS.t676 D2_5.t23 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS.t661 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2159 a_20041_8580# 7b_counter_0.MDFF_5.LD.t82 a_19841_8580# VSS.t1016 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2160 VDD.t898 CLK.t122 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t0 VDD.t897 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2161 VSS.t157 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_7309# VSS.t156 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2162 a_16386_n3644# p2_gen_magic_0.xnor_magic_5.OUT a_16186_n3644# VSS.t188 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2163 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD.t795 VDD.t794 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2164 OR_magic_1.VOUT a_30365_3514# VDD.t87 VDD.t86 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2165 a_16065_8580# 7b_counter_0.MDFF_5.LD.t83 a_15865_8580# VSS.t1011 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2166 VDD.t611 mux_magic_0.OR_magic_0.A a_34156_n889# VDD.t610 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2167 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t23 VSS.t857 VSS.t856 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2168 VSS.t400 a_19152_1223# a_20171_1669# VSS.t399 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2169 VDD.t2146 Q7.t24 a_1541_n8095# VDD.t769 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2170 a_26038_4932# 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# VDD.t127 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2171 VSS.t131 7b_counter_0.MDFF_5.QB.t8 7b_counter_0.MDFF_5.tspc2_magic_0.Q VSS.t130 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2172 a_27567_8496.t0 DFF_magic_0.D.t38 VDD.t1291 VDD.t1281 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2173 VDD.t1190 D2_5.t24 a_1209_3363# VDD.t1189 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2174 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD.t486 VDD.t485 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2175 a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VDD.t1646 VDD.t1645 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2176 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.CLK.t17 VDD.t1891 VDD.t1890 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2177 a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VDD.t1583 VDD.t28 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2178 a_5054_n1526# D2_3.t25 p2_gen_magic_0.xnor_magic_4.OUT VDD.t372 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2179 VDD.t1935 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n5540# VDD.t1249 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2180 a_5185_6275# 7b_counter_0.MDFF_3.tspc2_magic_0.Q VDD.t67 VDD.t66 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2181 VSS.t1267 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.IN VSS.t1266 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2182 a_20041_9774# 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_19841_9774# VSS.t890 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2183 VDD.t1972 D2_7.t24 a_5185_7469# VDD.t1971 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2184 divide_by_2_0.tg_magic_3.CLK.t1 OR_magic_2.VOUT.t25 VDD.t1669 VDD.t1668 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2185 VSS.t777 LD.t82 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VSS.t766 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2186 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD.t83 VDD.t1382 VDD.t1377 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2187 a_16065_9774# 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_15865_9774# VSS.t107 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2188 VSS.t1074 Q2.t31 7b_counter_0.3_inp_AND_magic_0.C VSS.t1073 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2189 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t123 VDD.t896 VDD.t502 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2190 VSS.t423 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_7308# VSS.t422 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2191 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7.t25 VSS.t1264 VSS.t1263 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2192 a_5036_n3597# D2_7.t25 p2_gen_magic_0.xnor_magic_5.OUT VDD.t107 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2193 a_23352_n6798# p3_gen_magic_0.P3.t16 a_23352_n5390# VDD.t1981 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2194 VSS.t431 a_8713_1625# a_8825_1669# VSS.t430 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2195 a_6725_684# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD.t718 VDD.t717 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2196 VDD.t783 a_12387_1769# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B VDD.t782 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2197 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD.t84 VDD.t1383 VDD.t1323 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2198 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t84 VDD.t1773 VDD.t1704 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2199 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# VDD.t331 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2200 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD.t85 VDD.t1384 VDD.t1375 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2201 a_1209_1059# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1409_1059# VSS.t335 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2202 VDD.t1148 7b_counter_0.MDFF_4.LD.t122 a_8411_3319# VDD.t1147 pfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2203 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t85 VDD.t1774 VDD.t1710 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2204 VSS.t5 CLK.t124 a_16065_8580# VSS.t4 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2205 a_11191_4932# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# VDD.t75 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2206 a_7303_3480# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7215_4932# VDD.t0 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2207 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.LD.t86 VDD.t1775 VDD.t1768 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2208 VSS.t1040 D2_1.t35 a_1957_n3150# VSS.t1039 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2209 divide_by_2_0.tg_magic_3.IN.t14 OR_magic_2.VOUT.t26 divide_by_2_0.tg_magic_1.IN VSS.t956 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2210 a_11292_n2115# p2_gen_magic_0.xnor_magic_4.OUT VDD.t125 VDD.t124 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2211 VSS.t871 divide_by_2_0.tg_magic_3.CLK.t19 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VSS.t870 nfet_03v3 ad=0.4928p pd=3.12u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2212 VDD.t908 CLK.t125 a_15865_8580# VDD.t907 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2213 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK.t126 VSS.t1 VSS.t0 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2214 a_1409_2253# LD.t86 a_1209_2253# VSS.t751 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2215 a_1975_n1973# p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_3.OUT.t1 VSS.t509 nfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2216 VDD.t1582 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_15865_4557# VDD.t26 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2217 VDD.t906 CLK.t127 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t0 VDD.t905 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2218 VDD.t1192 D2_5.t25 a_5185_2253# VDD.t1191 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2219 a_14556_n3644# p2_gen_magic_0.AND2_magic_1.A VDD.t1630 VDD.t1629 pfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2220 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4.t29 VSS.t887 VSS.t886 nfet_03v3 ad=0.2912p pd=1.64u as=0.4928p ps=3.12u w=1.12u l=0.56u
X2221 VDD.t516 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_15865_1059# VDD.t515 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2222 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_1209_1059# VDD.t245 VDD.t244 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2223 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_5185_7469# VDD.t724 VDD.t723 pfet_03v3 ad=0.2912p pd=1.64u as=0.2912p ps=1.64u w=1.12u l=0.56u
X2224 7b_counter_0.MDFF_0.tspc2_magic_0.D a_2749_3524# VDD.t750 VDD.t749 pfet_03v3 ad=0.4928p pd=3.12u as=0.4928p ps=3.12u w=1.12u l=0.56u
R0 VDD.t1015 VDD.t853 2420.69
R1 VDD.t568 VDD.t534 1683.52
R2 VDD.t542 VDD.t101 1646.52
R3 VDD.t1548 VDD.t1821 1275.86
R4 VDD.t1833 VDD.t1537 1275.86
R5 VDD.t991 VDD.t311 1199.13
R6 VDD.t61 VDD.t1595 1198.41
R7 VDD.t629 VDD.t55 1194.81
R8 VDD.t84 VDD.t451 1194.81
R9 VDD.t181 VDD.t725 1194.81
R10 VDD.t1255 VDD.t2058 1168.97
R11 VDD.t2046 VDD.t1240 1168.97
R12 VDD.t1179 VDD.t1629 1105.34
R13 VDD.t550 VDD.t1169 1105.34
R14 VDD.t211 VDD.t1300 1065.08
R15 VDD.t1802 VDD.t1606 1061.39
R16 VDD.t214 VDD.t742 1049.07
R17 VDD.t650 VDD.t217 1049.07
R18 VDD.t509 VDD.t1894 1046.14
R19 VDD.t337 VDD.t1660 1046.14
R20 VDD.t2106 VDD.t416 1046.14
R21 VDD.t798 VDD.t821 1046.14
R22 VDD.t885 VDD.t2150 1046.14
R23 VDD.t250 VDD.t1580 1046.14
R24 VDD.t332 VDD.n1008 1034.06
R25 VDD.t947 VDD.t159 1007.33
R26 VDD.t1919 VDD.t465 1007.33
R27 VDD.n1008 VDD.t1613 1007.16
R28 VDD.t2088 VDD.t1837 1006.9
R29 VDD.t1431 VDD.t1791 1006.9
R30 VDD.t1851 VDD.t2080 1006.9
R31 VDD.t2028 VDD.t1451 1006.9
R32 VDD.t1963 VDD.t2005 993.104
R33 VDD.t1996 VDD.t1955 993.104
R34 VDD.t283 VDD.t329 958.63
R35 VDD.t695 VDD.t636 957.376
R36 VDD.t930 VDD.t319 957.376
R37 VDD.t717 VDD.t1550 957.376
R38 VDD.t642 VDD.t784 957.376
R39 VDD.t920 VDD.t134 957.376
R40 VDD.t95 VDD.t350 957.376
R41 VDD.n1027 VDD.t1119 921.26
R42 VDD.n1027 VDD.t1056 921.26
R43 VDD.t1351 VDD.t204 864.109
R44 VDD.t45 VDD.t1748 864.109
R45 VDD.t369 VDD.t1704 864.109
R46 VDD.t189 VDD.t1036 864.109
R47 VDD.t574 VDD.t594 861.423
R48 VDD.t570 VDD.t932 842.491
R49 VDD.t521 VDD.t697 842.491
R50 VDD.t1107 VDD.t517 842.491
R51 VDD.t1022 VDD.t1026 842.491
R52 VDD.t644 VDD.t270 842.491
R53 VDD.n1527 VDD.t591 841.558
R54 VDD.n897 VDD.t443 841.558
R55 VDD.t1197 VDD.t17 806.37
R56 VDD.t531 VDD.t129 806.37
R57 VDD.t1159 VDD.t1888 787.708
R58 VDD.t1466 VDD.t969 787.708
R59 VDD.t949 VDD.t712 787.708
R60 VDD.t1292 VDD.t983 787.708
R61 VDD.t1939 VDD.t1504 787.708
R62 VDD.t1982 VDD.t143 787.708
R63 VDD.t1977 VDD.t901 787.708
R64 VDD.t1480 VDD.t170 787.708
R65 VDD.t2060 VDD.t1502 787.708
R66 VDD.t1017 VDD.t1021 787.708
R67 VDD.t1210 VDD.t91 787.708
R68 VDD.t1167 VDD.t380 787.708
R69 VDD.t1560 VDD.t388 782.313
R70 VDD.t776 VDD.t1890 782.313
R71 VDD.t839 VDD.t737 782.313
R72 VDD.t1206 VDD.t963 782.313
R73 VDD.t731 VDD.t985 782.313
R74 VDD.t710 VDD.t811 782.313
R75 VDD.t1654 VDD.t194 782.313
R76 VDD.t1590 VDD.t1516 782.313
R77 VDD.t2017 VDD.t1518 782.313
R78 VDD.t144 VDD.t1656 782.313
R79 VDD.t1933 VDD.t1898 782.313
R80 VDD.t2108 VDD.t317 782.313
R81 VDD.t1900 VDD.t1644 782.313
R82 VDD.t171 VDD.t2096 782.313
R83 VDD.t831 VDD.t471 782.313
R84 VDD.t616 VDD.t1488 782.313
R85 VDD.t149 VDD.t1494 782.313
R86 VDD.t1020 VDD.t863 782.313
R87 VDD.t961 VDD.t227 782.313
R88 VDD.t89 VDD.t1917 782.313
R89 VDD.t1610 VDD.t1878 782.313
R90 VDD.t378 VDD.t1568 782.313
R91 VDD.t80 VDD.t190 774.006
R92 VDD.t37 VDD.t361 774.006
R93 VDD.t1710 VDD.t1746 757.283
R94 VDD.n1471 VDD.t1599 757.01
R95 VDD.n977 VDD.t536 755.245
R96 VDD.n1526 VDD.t749 755.245
R97 VDD.n1604 VDD.t309 755.245
R98 VDD.n1007 VDD.t1615 755.245
R99 VDD.n1506 VDD.t20 755.245
R100 VDD.n950 VDD.t234 755.245
R101 VDD.t813 VDD.t977 746.33
R102 VDD.t1904 VDD.t897 746.33
R103 VDD.t1913 VDD.t1500 746.33
R104 VDD.t967 VDD.t837 746.33
R105 VDD.t1666 VDD.t1506 741.497
R106 VDD.t1562 VDD.t1884 741.497
R107 VDD.n146 VDD.n144 721.963
R108 VDD.t1578 VDD.t260 713.571
R109 VDD.t894 VDD.t786 713.571
R110 VDD.t1423 VDD.t393 713.571
R111 VDD.t2104 VDD.t2116 713.571
R112 VDD.t835 VDD.t1009 713.571
R113 VDD.t505 VDD.t733 699.505
R114 VDD.t339 VDD.t2016 699.505
R115 VDD.t1642 VDD.t414 699.505
R116 VDD.t794 VDD.t151 699.505
R117 VDD.t228 VDD.t2152 699.505
R118 VDD.t254 VDD.t1612 699.505
R119 VDD.t1377 VDD.t483 669.359
R120 VDD.t1310 VDD.t367 669.359
R121 VDD.t1323 VDD.t493 669.359
R122 VDD.t487 VDD.t1736 669.359
R123 VDD.t119 VDD.t1742 669.359
R124 VDD.t7 VDD.t1726 669.359
R125 VDD.t1554 VDD.t1714 669.359
R126 VDD.t1584 VDD.t1075 669.359
R127 VDD.t513 VDD.t1100 669.359
R128 VDD.t1776 VDD.t702 669.359
R129 VDD.t580 VDD.t638 643.899
R130 VDD.t358 VDD.t376 643.899
R131 VDD.t1050 VDD.n1027 642.857
R132 VDD.n1027 VDD.t1054 642.857
R133 VDD.t2086 VDD.t546 634.721
R134 VDD.t372 VDD.t2050 634.721
R135 VDD.t1399 VDD.t654 634.721
R136 VDD.t405 VDD.t1800 634.721
R137 VDD.t1961 VDD.t107 634.721
R138 VDD.t423 VDD.t1823 634.721
R139 VDD.t1175 VDD.t408 634.721
R140 VDD.t560 VDD.t2078 634.721
R141 VDD.t2040 VDD.t109 634.721
R142 VDD.t562 VDD.t1389 634.721
R143 VDD.t2030 VDD.t774 634.721
R144 VDD.t735 VDD.t1953 634.721
R145 VDD.t1813 VDD.t1620 634.721
R146 VDD.t549 VDD.t1187 634.721
R147 VDD.t715 VDD.t719 621.245
R148 VDD.t915 VDD.t917 621.245
R149 VDD.t287 VDD.t489 621.072
R150 VDD.n1184 VDD 608.955
R151 VDD.t534 VDD.n978 606.742
R152 VDD.t1277 VDD.t1409 572.513
R153 VDD.t1077 VDD.t1058 566.929
R154 VDD.t1119 VDD.t1077 566.929
R155 VDD.t1056 VDD.t1111 566.929
R156 VDD.t1111 VDD.t1072 566.929
R157 VDD.t1306 VDD.t1379 566.929
R158 VDD.t1306 VDD.t1327 566.929
R159 VDD.t1306 VDD.t1369 566.929
R160 VDD.t1306 VDD.t1317 566.929
R161 VDD.t401 VDD.t629 561.039
R162 VDD.t462 VDD.t84 561.039
R163 VDD.n1212 VDD.t778 549.321
R164 VDD.n1300 VDD.t1207 549.321
R165 VDD.n313 VDD.t1588 549.321
R166 VDD.n367 VDD.t1934 549.321
R167 VDD.n578 VDD.t617 549.321
R168 VDD.t1230 VDD.t2130 541.585
R169 VDD.n1009 VDD.t1613 534.769
R170 VDD.n703 VDD.t128 522.145
R171 VDD.t455 VDD.n145 522.078
R172 VDD.t1530 VDD.t1673 519.126
R173 VDD.n761 VDD.t501 517.442
R174 VDD.t185 VDD.t686 506.267
R175 VDD.t1597 VDD.t283 504.673
R176 VDD.t100 VDD.t695 503.497
R177 VDD.t748 VDD.t930 503.497
R178 VDD.t661 VDD.t717 503.497
R179 VDD.t334 VDD.t642 503.497
R180 VDD.t16 VDD.t920 503.497
R181 VDD.t232 VDD.t95 503.497
R182 VDD.t671 VDD.t128 503.497
R183 VDD.n899 VDD.t77 496.933
R184 VDD.n1212 VDD.t256 491.791
R185 VDD.n1300 VDD.t788 491.791
R186 VDD.n313 VDD.t395 491.791
R187 VDD.n367 VDD.t2118 491.791
R188 VDD.n578 VDD.t1007 491.791
R189 VDD.n703 VDD.t131 484.849
R190 VDD.t1095 VDD.t1028 429.604
R191 VDD.n1685 VDD.t994 423.697
R192 VDD.n56 VDD.t2021 421.245
R193 VDD.n110 VDD.t2158 421.245
R194 VDD.t246 VDD.n110 421.245
R195 VDD.n56 VDD.t1216 421.245
R196 VDD.n1661 VDD.t11 421.245
R197 VDD.n1661 VDD.t606 421.245
R198 VDD.n1668 VDD.t2173 421.245
R199 VDD.n1668 VDD.t343 421.245
R200 VDD.n677 VDD.t294 421.245
R201 VDD.n688 VDD.t662 421.245
R202 VDD.n688 VDD.t566 421.245
R203 VDD.n677 VDD.t762 421.245
R204 VDD.t502 VDD.t554 421.245
R205 VDD.t589 VDD.n1262 421.245
R206 VDD.n1262 VDD.t923 421.245
R207 VDD.n761 VDD.t211 416.668
R208 VDD.t596 VDD.t936 404.495
R209 VDD.t594 VDD.t596 404.495
R210 VDD.t544 VDD.t574 404.495
R211 VDD.t571 VDD.t544 404.495
R212 VDD.t102 VDD.t693 404.495
R213 VDD.t404 VDD.t1347 397.445
R214 VDD.t77 VDD.t1030 397.269
R215 VDD.t1093 VDD.t231 397.269
R216 VDD.n1184 VDD.t676 396.553
R217 VDD.t165 VDD.t163 395.604
R218 VDD.t1862 VDD.t165 395.604
R219 VDD.t1860 VDD.t1862 395.604
R220 VDD.t161 VDD.t1860 395.604
R221 VDD.t159 VDD.t161 395.604
R222 VDD.t945 VDD.t947 395.604
R223 VDD.t756 VDD.t945 395.604
R224 VDD.t758 VDD.t756 395.604
R225 VDD.t1631 VDD.t758 395.604
R226 VDD.t1629 VDD.t1631 395.604
R227 VDD.t1760 VDD.t1724 395.604
R228 VDD.t879 VDD.t1760 395.604
R229 VDD.t845 VDD.t879 395.604
R230 VDD.t2019 VDD.t845 395.604
R231 VDD.t2021 VDD.t2019 395.604
R232 VDD.t636 VDD.t634 395.604
R233 VDD.t634 VDD.t2036 395.604
R234 VDD.t2036 VDD.t2044 395.604
R235 VDD.t2044 VDD.t1102 395.604
R236 VDD.t1102 VDD.t1097 395.604
R237 VDD.t55 VDD.t57 395.604
R238 VDD.t57 VDD.t869 395.604
R239 VDD.t869 VDD.t883 395.604
R240 VDD.t883 VDD.t1312 395.604
R241 VDD.t1312 VDD.t1349 395.604
R242 VDD.t319 VDD.t321 395.604
R243 VDD.t321 VDD.t1189 395.604
R244 VDD.t1189 VDD.t1171 395.604
R245 VDD.t1171 VDD.t1338 395.604
R246 VDD.t1338 VDD.t1362 395.604
R247 VDD.t2158 VDD.t2160 395.604
R248 VDD.t2160 VDD.t875 395.604
R249 VDD.t875 VDD.t881 395.604
R250 VDD.t881 VDD.t1314 395.604
R251 VDD.t1314 VDD.t1353 395.604
R252 VDD.t244 VDD.t246 395.604
R253 VDD.t1520 VDD.t244 395.604
R254 VDD.t1546 VDD.t1520 395.604
R255 VDD.t481 VDD.t1546 395.604
R256 VDD.t483 VDD.t481 395.604
R257 VDD.t713 VDD.t715 395.604
R258 VDD.t752 VDD.t713 395.604
R259 VDD.t754 VDD.t752 395.604
R260 VDD.t365 VDD.t754 395.604
R261 VDD.t367 VDD.t365 395.604
R262 VDD.t1550 VDD.t1552 395.604
R263 VDD.t1552 VDD.t1191 395.604
R264 VDD.t1191 VDD.t1173 395.604
R265 VDD.t1173 VDD.t1344 395.604
R266 VDD.t1344 VDD.t1366 395.604
R267 VDD.t1138 VDD.t1109 395.604
R268 VDD.t1835 VDD.t1138 395.604
R269 VDD.t1829 VDD.t1835 395.604
R270 VDD.t782 VDD.t1829 395.604
R271 VDD.t784 VDD.t782 395.604
R272 VDD.t573 VDD.t570 395.604
R273 VDD.t575 VDD.t538 395.604
R274 VDD.t538 VDD.t540 395.604
R275 VDD.t101 VDD.t99 395.604
R276 VDD.t697 VDD.t691 395.604
R277 VDD.t519 VDD.t521 395.604
R278 VDD.t938 VDD.t519 395.604
R279 VDD.t934 VDD.t938 395.604
R280 VDD.t515 VDD.t934 395.604
R281 VDD.t517 VDD.t515 395.604
R282 VDD.t1024 VDD.t1022 395.604
R283 VDD.t987 VDD.t1024 395.604
R284 VDD.t989 VDD.t987 395.604
R285 VDD.t268 VDD.t989 395.604
R286 VDD.t270 VDD.t268 395.604
R287 VDD.t646 VDD.t644 395.604
R288 VDD.t331 VDD.t332 395.604
R289 VDD.t1730 VDD.t1712 395.604
R290 VDD.t1397 VDD.t1730 395.604
R291 VDD.t1391 VDD.t1397 395.604
R292 VDD.t453 VDD.t1391 395.604
R293 VDD.t451 VDD.t453 395.604
R294 VDD.t1048 VDD.t1133 395.604
R295 VDD.t1915 VDD.t1048 395.604
R296 VDD.t890 VDD.t1915 395.604
R297 VDD.t192 VDD.t890 395.604
R298 VDD.t190 VDD.t192 395.604
R299 VDD.t1038 VDD.t1147 395.604
R300 VDD.t1817 VDD.t1038 395.604
R301 VDD.t1815 VDD.t1817 395.604
R302 VDD.t640 VDD.t1815 395.604
R303 VDD.t638 VDD.t640 395.604
R304 VDD.t725 VDD.t723 395.604
R305 VDD.t723 VDD.t1971 395.604
R306 VDD.t1971 VDD.t1951 395.604
R307 VDD.t1951 VDD.t1336 395.604
R308 VDD.t1336 VDD.t1364 395.604
R309 VDD.t913 VDD.t915 395.604
R310 VDD.t59 VDD.t913 395.604
R311 VDD.t64 VDD.t59 395.604
R312 VDD.t495 VDD.t64 395.604
R313 VDD.t493 VDD.t495 395.604
R314 VDD.t134 VDD.t136 395.604
R315 VDD.t136 VDD.t1969 395.604
R316 VDD.t1969 VDD.t1949 395.604
R317 VDD.t1949 VDD.t1334 395.604
R318 VDD.t1334 VDD.t1360 395.604
R319 VDD.t1758 VDD.t1752 395.604
R320 VDD.t1403 VDD.t1758 395.604
R321 VDD.t1401 VDD.t1403 395.604
R322 VDD.t327 VDD.t1401 395.604
R323 VDD.t329 VDD.t327 395.604
R324 VDD.t485 VDD.t487 395.604
R325 VDD.t669 VDD.t485 395.604
R326 VDD.t667 VDD.t669 395.604
R327 VDD.t491 VDD.t667 395.604
R328 VDD.t489 VDD.t491 395.604
R329 VDD.t117 VDD.t119 395.604
R330 VDD.t1232 VDD.t117 395.604
R331 VDD.t1251 VDD.t1232 395.604
R332 VDD.t1218 VDD.t1251 395.604
R333 VDD.t1216 VDD.t1218 395.604
R334 VDD.t11 VDD.t13 395.604
R335 VDD.t13 VDD.t843 395.604
R336 VDD.t843 VDD.t855 395.604
R337 VDD.t855 VDD.t9 395.604
R338 VDD.t9 VDD.t7 395.604
R339 VDD.t606 VDD.t608 395.604
R340 VDD.t608 VDD.t907 395.604
R341 VDD.t907 VDD.t1907 395.604
R342 VDD.t1907 VDD.t1720 395.604
R343 VDD.t1720 VDD.t1718 395.604
R344 VDD.t2173 VDD.t2175 395.604
R345 VDD.t2175 VDD.t179 395.604
R346 VDD.t179 VDD.t177 395.604
R347 VDD.t177 VDD.t1556 395.604
R348 VDD.t1556 VDD.t1554 395.604
R349 VDD.t343 VDD.t345 395.604
R350 VDD.t345 VDD.t1787 395.604
R351 VDD.t1787 VDD.t1797 395.604
R352 VDD.t1797 VDD.t1732 395.604
R353 VDD.t1732 VDD.t1716 395.604
R354 VDD.t1143 VDD.t1117 395.604
R355 VDD.t892 VDD.t1143 395.604
R356 VDD.t903 VDD.t892 395.604
R357 VDD.t296 VDD.t903 395.604
R358 VDD.t294 VDD.t296 395.604
R359 VDD.t1123 VDD.t1081 395.604
R360 VDD.t2082 VDD.t1123 395.604
R361 VDD.t2094 VDD.t2082 395.604
R362 VDD.t664 VDD.t2094 395.604
R363 VDD.t662 VDD.t664 395.604
R364 VDD.t1586 VDD.t1584 395.604
R365 VDD.t626 VDD.t1586 395.604
R366 VDD.t624 VDD.t626 395.604
R367 VDD.t564 VDD.t624 395.604
R368 VDD.t566 VDD.t564 395.604
R369 VDD.t511 VDD.t513 395.604
R370 VDD.t1691 VDD.t511 395.604
R371 VDD.t1684 VDD.t1691 395.604
R372 VDD.t760 VDD.t1684 395.604
R373 VDD.t762 VDD.t760 395.604
R374 VDD.t1052 VDD.t1135 395.604
R375 VDD.t2074 VDD.t1052 395.604
R376 VDD.t2076 VDD.t2074 395.604
R377 VDD.t556 VDD.t2076 395.604
R378 VDD.t554 VDD.t556 395.604
R379 VDD.t376 VDD.t374 395.604
R380 VDD.t374 VDD.t2048 395.604
R381 VDD.t2048 VDD.t2054 395.604
R382 VDD.t2054 VDD.t1140 395.604
R383 VDD.t1140 VDD.t1127 395.604
R384 VDD.t361 VDD.t363 395.604
R385 VDD.t363 VDD.t827 395.604
R386 VDD.t827 VDD.t859 395.604
R387 VDD.t859 VDD.t1131 395.604
R388 VDD.t1131 VDD.t1129 395.604
R389 VDD.t350 VDD.t352 395.604
R390 VDD.t352 VDD.t1804 395.604
R391 VDD.t1804 VDD.t1780 395.604
R392 VDD.t1780 VDD.t1708 395.604
R393 VDD.t1708 VDD.t1706 395.604
R394 VDD.t1606 VDD.t1608 395.604
R395 VDD.t1608 VDD.t909 395.604
R396 VDD.t909 VDD.t911 395.604
R397 VDD.t911 VDD.t1921 395.604
R398 VDD.t1921 VDD.t1919 395.604
R399 VDD.t465 VDD.t463 395.604
R400 VDD.t463 VDD.t105 395.604
R401 VDD.t105 VDD.t103 395.604
R402 VDD.t103 VDD.t552 395.604
R403 VDD.t552 VDD.t550 395.604
R404 VDD.t587 VDD.t589 395.604
R405 VDD.t1149 VDD.t587 395.604
R406 VDD.t1151 VDD.t1149 395.604
R407 VDD.t704 VDD.t1151 395.604
R408 VDD.t702 VDD.t704 395.604
R409 VDD.t923 VDD.t925 395.604
R410 VDD.t925 VDD.t1943 395.604
R411 VDD.t1943 VDD.t1937 395.604
R412 VDD.t1937 VDD.t1795 395.604
R413 VDD.t1795 VDD.t1811 395.604
R414 VDD.n1045 VDD.t575 390.111
R415 VDD.n1029 VDD.t1087 380.952
R416 VDD.n1006 VDD.t1145 380.952
R417 VDD.t1674 VDD.n1369 377.587
R418 VDD.n1361 VDD.t1839 377.587
R419 VDD.t1257 VDD.n1356 377.587
R420 VDD.n1376 VDD.t2142 377.587
R421 VDD.n1387 VDD.t1436 377.587
R422 VDD.n1395 VDD.t2007 377.587
R423 VDD.n1406 VDD.t1542 377.587
R424 VDD.n522 VDD.t1688 377.587
R425 VDD.n530 VDD.t1853 377.587
R426 VDD.n535 VDD.t1245 377.587
R427 VDD.t2133 VDD.n515 377.587
R428 VDD.n501 VDD.t1454 377.587
R429 VDD.t1998 VDD.n492 377.587
R430 VDD.n478 VDD.t1527 377.587
R431 VDD.t256 VDD.t258 372.414
R432 VDD.t260 VDD.t262 372.414
R433 VDD.t1155 VDD.t1157 372.414
R434 VDD.t1153 VDD.t1159 372.414
R435 VDD.t788 VDD.t792 372.414
R436 VDD.t786 VDD.t790 372.414
R437 VDD.t1459 VDD.t1470 372.414
R438 VDD.t1461 VDD.t1466 372.414
R439 VDD.t1682 VDD.t1674 372.414
R440 VDD.t1671 VDD.t1678 372.414
R441 VDD.t1839 VDD.t1847 372.414
R442 VDD.t1837 VDD.t1855 372.414
R443 VDD.t2092 VDD.t2088 372.414
R444 VDD.t2072 VDD.t2086 372.414
R445 VDD.t1238 VDD.t1257 372.414
R446 VDD.t1247 VDD.t1255 372.414
R447 VDD.t2058 VDD.t2052 372.414
R448 VDD.t2050 VDD.t2038 372.414
R449 VDD.t1405 VDD.t1395 372.414
R450 VDD.t1387 VDD.t1399 372.414
R451 VDD.t2142 VDD.t2137 372.414
R452 VDD.t2139 VDD.t2144 372.414
R453 VDD.t1441 VDD.t1436 372.414
R454 VDD.t1444 VDD.t1431 372.414
R455 VDD.t1791 VDD.t1806 372.414
R456 VDD.t1800 VDD.t1789 372.414
R457 VDD.t2007 VDD.t2012 372.414
R458 VDD.t2005 VDD.t1992 372.414
R459 VDD.t1965 VDD.t1963 372.414
R460 VDD.t1957 VDD.t1961 372.414
R461 VDD.t1525 VDD.t1542 372.414
R462 VDD.t1534 VDD.t1548 372.414
R463 VDD.t1821 VDD.t1825 372.414
R464 VDD.t1823 VDD.t1831 372.414
R465 VDD.t1183 VDD.t1179 372.414
R466 VDD.t1185 VDD.t1175 372.414
R467 VDD.t867 VDD.t813 372.414
R468 VDD.t905 VDD.t861 372.414
R469 VDD.t953 VDD.t955 372.414
R470 VDD.t951 VDD.t949 372.414
R471 VDD.t1298 VDD.t1294 372.414
R472 VDD.t1300 VDD.t1259 372.414
R473 VDD.t1261 VDD.t1304 372.414
R474 VDD.t1263 VDD.t1292 372.414
R475 VDD.t395 VDD.t391 372.414
R476 VDD.t393 VDD.t397 372.414
R477 VDD.t1945 VDD.t1941 372.414
R478 VDD.t1947 VDD.t1939 372.414
R479 VDD.t1984 VDD.t1988 372.414
R480 VDD.t1986 VDD.t1982 372.414
R481 VDD.t1979 VDD.t1973 372.414
R482 VDD.t1975 VDD.t1977 372.414
R483 VDD.t2118 VDD.t2114 372.414
R484 VDD.t2116 VDD.t2112 372.414
R485 VDD.t897 VDD.t841 372.414
R486 VDD.t865 VDD.t888 372.414
R487 VDD.t1484 VDD.t1486 372.414
R488 VDD.t1482 VDD.t1480 372.414
R489 VDD.t1688 VDD.t1676 372.414
R490 VDD.t1686 VDD.t1693 372.414
R491 VDD.t1843 VDD.t1853 372.414
R492 VDD.t1845 VDD.t1851 372.414
R493 VDD.t2080 VDD.t2084 372.414
R494 VDD.t2078 VDD.t2090 372.414
R495 VDD.t1245 VDD.t1225 372.414
R496 VDD.t1240 VDD.t1236 372.414
R497 VDD.t2042 VDD.t2046 372.414
R498 VDD.t2056 VDD.t2040 372.414
R499 VDD.t1393 VDD.t1385 372.414
R500 VDD.t1389 VDD.t1407 372.414
R501 VDD.t2125 VDD.t2133 372.414
R502 VDD.t2128 VDD.t2135 372.414
R503 VDD.t1454 VDD.t1427 372.414
R504 VDD.t1451 VDD.t1434 372.414
R505 VDD.t2032 VDD.t2028 372.414
R506 VDD.t2034 VDD.t2030 372.414
R507 VDD.t2003 VDD.t1998 372.414
R508 VDD.t2010 VDD.t1996 372.414
R509 VDD.t1955 VDD.t1959 372.414
R510 VDD.t1953 VDD.t1967 372.414
R511 VDD.t1527 VDD.t1544 372.414
R512 VDD.t1537 VDD.t1522 372.414
R513 VDD.t1819 VDD.t1833 372.414
R514 VDD.t1827 VDD.t1813 372.414
R515 VDD.t1169 VDD.t1177 372.414
R516 VDD.t1187 VDD.t1181 372.414
R517 VDD.t1808 VDD.t1793 372.414
R518 VDD.t1782 VDD.t1802 372.414
R519 VDD.t1007 VDD.t1003 372.414
R520 VDD.t1009 VDD.t1005 372.414
R521 VDD.t2062 VDD.t2065 372.414
R522 VDD.t2067 VDD.t2060 372.414
R523 VDD.t1911 VDD.t1913 372.414
R524 VDD.t817 VDD.t857 372.414
R525 VDD.t837 VDD.t849 372.414
R526 VDD.t853 VDD.t815 372.414
R527 VDD.t1011 VDD.t1015 372.414
R528 VDD.t1013 VDD.t1017 372.414
R529 VDD.t1214 VDD.t1208 372.414
R530 VDD.t1212 VDD.t1210 372.414
R531 VDD.t1163 VDD.t1161 372.414
R532 VDD.t1165 VDD.t1167 372.414
R533 VDD.t507 VDD.t509 367.974
R534 VDD.t503 VDD.t505 367.974
R535 VDD.t335 VDD.t337 367.974
R536 VDD.t341 VDD.t339 367.974
R537 VDD.t416 VDD.t420 367.974
R538 VDD.t414 VDD.t418 367.974
R539 VDD.t800 VDD.t798 367.974
R540 VDD.t796 VDD.t794 367.974
R541 VDD.t2150 VDD.t2154 367.974
R542 VDD.t2152 VDD.t2156 367.974
R543 VDD.t248 VDD.t250 367.974
R544 VDD.t252 VDD.t254 367.974
R545 VDD.t1566 VDD.t1578 367.348
R546 VDD.t1558 VDD.t1560 367.348
R547 VDD.t388 VDD.t390 367.348
R548 VDD.t390 VDD.t389 367.348
R549 VDD.t1888 VDD.t1880 367.348
R550 VDD.t1890 VDD.t1876 367.348
R551 VDD.t777 VDD.t776 367.348
R552 VDD.t778 VDD.t777 367.348
R553 VDD.t873 VDD.t894 367.348
R554 VDD.t819 VDD.t839 367.348
R555 VDD.t737 VDD.t736 367.348
R556 VDD.t736 VDD.t738 367.348
R557 VDD.t969 VDD.t959 367.348
R558 VDD.t963 VDD.t957 367.348
R559 VDD.t1205 VDD.t1206 367.348
R560 VDD.t1207 VDD.t1205 367.348
R561 VDD.t733 VDD.t732 367.348
R562 VDD.t732 VDD.t731 367.348
R563 VDD.t985 VDD.t975 367.348
R564 VDD.t977 VDD.t979 367.348
R565 VDD.t712 VDD.t711 367.348
R566 VDD.t711 VDD.t710 367.348
R567 VDD.t811 VDD.t851 367.348
R568 VDD.t1894 VDD.t899 367.348
R569 VDD.t983 VDD.t971 367.348
R570 VDD.t1652 VDD.t1423 367.348
R571 VDD.t1664 VDD.t1654 367.348
R572 VDD.t194 VDD.t196 367.348
R573 VDD.t196 VDD.t195 367.348
R574 VDD.t1504 VDD.t1508 367.348
R575 VDD.t1516 VDD.t1514 367.348
R576 VDD.t1589 VDD.t1590 367.348
R577 VDD.t1588 VDD.t1589 367.348
R578 VDD.t2016 VDD.t2018 367.348
R579 VDD.t2018 VDD.t2017 367.348
R580 VDD.t1518 VDD.t1510 367.348
R581 VDD.t1506 VDD.t1512 367.348
R582 VDD.t1421 VDD.t1666 367.348
R583 VDD.t1658 VDD.t1668 367.348
R584 VDD.t143 VDD.t142 367.348
R585 VDD.t142 VDD.t144 367.348
R586 VDD.t1656 VDD.t1662 367.348
R587 VDD.t1660 VDD.t1425 367.348
R588 VDD.t901 VDD.t829 367.348
R589 VDD.t1898 VDD.t871 367.348
R590 VDD.t1932 VDD.t1933 367.348
R591 VDD.t1934 VDD.t1932 367.348
R592 VDD.t2110 VDD.t2104 367.348
R593 VDD.t2100 VDD.t2108 367.348
R594 VDD.t317 VDD.t316 367.348
R595 VDD.t316 VDD.t318 367.348
R596 VDD.t1643 VDD.t1642 367.348
R597 VDD.t1644 VDD.t1643 367.348
R598 VDD.t825 VDD.t1900 367.348
R599 VDD.t847 VDD.t1904 367.348
R600 VDD.t170 VDD.t172 367.348
R601 VDD.t172 VDD.t171 367.348
R602 VDD.t2096 VDD.t2102 367.348
R603 VDD.t2098 VDD.t2106 367.348
R604 VDD.t877 VDD.t835 367.348
R605 VDD.t1902 VDD.t831 367.348
R606 VDD.t471 VDD.t470 367.348
R607 VDD.t470 VDD.t472 367.348
R608 VDD.t1502 VDD.t1490 367.348
R609 VDD.t1488 VDD.t1496 367.348
R610 VDD.t615 VDD.t616 367.348
R611 VDD.t617 VDD.t615 367.348
R612 VDD.t151 VDD.t150 367.348
R613 VDD.t150 VDD.t149 367.348
R614 VDD.t1494 VDD.t1492 367.348
R615 VDD.t1500 VDD.t1498 367.348
R616 VDD.t1021 VDD.t1019 367.348
R617 VDD.t1019 VDD.t1020 367.348
R618 VDD.t863 VDD.t1909 367.348
R619 VDD.t821 VDD.t1896 367.348
R620 VDD.t229 VDD.t228 367.348
R621 VDD.t227 VDD.t229 367.348
R622 VDD.t965 VDD.t961 367.348
R623 VDD.t1892 VDD.t967 367.348
R624 VDD.t91 VDD.t90 367.348
R625 VDD.t90 VDD.t89 367.348
R626 VDD.t1917 VDD.t823 367.348
R627 VDD.t833 VDD.t885 367.348
R628 VDD.t1612 VDD.t1611 367.348
R629 VDD.t1611 VDD.t1610 367.348
R630 VDD.t1878 VDD.t1882 367.348
R631 VDD.t1884 VDD.t1886 367.348
R632 VDD.t1564 VDD.t1562 367.348
R633 VDD.t1574 VDD.t1570 367.348
R634 VDD.t380 VDD.t379 367.348
R635 VDD.t379 VDD.t378 367.348
R636 VDD.t1568 VDD.t1572 367.348
R637 VDD.t1580 VDD.t1576 367.348
R638 VDD.n1690 VDD.t1923 364.93
R639 VDD.t1413 VDD.n1689 364.93
R640 VDD.t998 VDD.n1684 364.93
R641 VDD.t1302 VDD.t1296 363.637
R642 VDD.t333 VDD.t648 357.616
R643 VDD.t99 VDD.n1043 353.481
R644 VDD.t1375 VDD.t264 347.959
R645 VDD.t745 VDD.t70 337.587
R646 VDD.t739 VDD.t214 337.587
R647 VDD.t478 VDD.t208 337.587
R648 VDD.t217 VDD.t764 337.587
R649 VDD.n1028 VDD.t1050 318.682
R650 VDD.t1054 VDD.n1026 318.682
R651 VDD.t676 VDD.t682 316.827
R652 VDD.n68 VDD.t167 313.651
R653 VDD.n961 VDD.t2170 313.651
R654 VDD.n1369 VDD.t802 307.135
R655 VDD.n1361 VDD.t323 307.135
R656 VDD.n1356 VDD.t302 307.135
R657 VDD.n1376 VDD.t434 307.135
R658 VDD.t173 VDD.n1387 307.135
R659 VDD.n1395 VDD.t3 307.135
R660 VDD.t138 VDD.n1406 307.135
R661 VDD.n522 VDD.t1635 307.135
R662 VDD.t24 VDD.n530 307.135
R663 VDD.n535 VDD.t1249 307.135
R664 VDD.n515 VDD.t769 307.135
R665 VDD.n501 VDD.t300 307.135
R666 VDD.n492 VDD.t598 307.135
R667 VDD.n478 VDD.t236 307.135
R668 VDD.t1593 VDD.t1042 284.159
R669 VDD.t28 VDD.t1034 284.159
R670 VDD.n1527 VDD.t401 280.519
R671 VDD.n897 VDD.t462 280.519
R672 VDD.t386 VDD.t631 276.796
R673 VDD.t80 VDD.t71 276.618
R674 VDD.t37 VDD.t33 276.618
R675 VDD.n1044 VDD.t568 256.555
R676 VDD.n1677 VDD.n1676 254.209
R677 VDD.n1471 VDD.t1597 252.337
R678 VDD.n977 VDD.t100 251.749
R679 VDD.n1526 VDD.t748 251.749
R680 VDD.n1604 VDD.t661 251.749
R681 VDD.n1007 VDD.t334 251.749
R682 VDD.n1506 VDD.t16 251.749
R683 VDD.n950 VDD.t232 251.749
R684 VDD.n1044 VDD.t542 250.917
R685 VDD.t354 VDD.t278 244.154
R686 VDD.t576 VDD.t584 238.714
R687 VDD.t1329 VDD.t1377 233.011
R688 VDD.t1319 VDD.t1310 233.011
R689 VDD.t1736 VDD.t1722 233.011
R690 VDD.t1726 VDD.t1756 233.011
R691 VDD.t1742 VDD.t1768 233.011
R692 VDD.t1714 VDD.t1739 233.011
R693 VDD.t1075 VDD.t1083 233.011
R694 VDD.t1100 VDD.t1104 233.011
R695 VDD.t1784 VDD.t1776 233.011
R696 VDD.t497 VDD.n1675 230.641
R697 VDD.n1493 VDD.t1331 224.381
R698 VDD.n1211 VDD.t262 215.518
R699 VDD.n1217 VDD.t1153 215.518
R700 VDD.t790 VDD.n1307 215.518
R701 VDD.n1291 VDD.t1461 215.518
R702 VDD.n1370 VDD.t1682 215.518
R703 VDD.n1364 VDD.t1847 215.518
R704 VDD.n1365 VDD.t2092 215.518
R705 VDD.n1357 VDD.t1238 215.518
R706 VDD.n1360 VDD.t2052 215.518
R707 VDD.n249 VDD.t1405 215.518
R708 VDD.t2137 VDD.n1375 215.518
R709 VDD.n1382 VDD.t1441 215.518
R710 VDD.t1806 VDD.n1381 215.518
R711 VDD.t2012 VDD.n1394 215.518
R712 VDD.n1388 VDD.t1965 215.518
R713 VDD.n1401 VDD.t1525 215.518
R714 VDD.t1825 VDD.n1400 215.518
R715 VDD.n1407 VDD.t1183 215.518
R716 VDD.n744 VDD.t867 215.518
R717 VDD.n728 VDD.t953 215.518
R718 VDD.n760 VDD.t1298 215.518
R719 VDD.n723 VDD.t1263 215.518
R720 VDD.n312 VDD.t397 215.518
R721 VDD.n318 VDD.t1947 215.518
R722 VDD.n323 VDD.t1984 215.518
R723 VDD.n358 VDD.t1975 215.518
R724 VDD.t2112 VDD.n374 215.518
R725 VDD.t841 VDD.n550 215.518
R726 VDD.n285 VDD.t1484 215.518
R727 VDD.t1676 VDD.n521 215.518
R728 VDD.n527 VDD.t1843 215.518
R729 VDD.t2084 VDD.n526 215.518
R730 VDD.t1225 VDD.n534 215.518
R731 VDD.n531 VDD.t2042 215.518
R732 VDD.n404 VDD.t1393 215.518
R733 VDD.n516 VDD.t2125 215.518
R734 VDD.n508 VDD.t1427 215.518
R735 VDD.n509 VDD.t2032 215.518
R736 VDD.n493 VDD.t2003 215.518
R737 VDD.n500 VDD.t1959 215.518
R738 VDD.n485 VDD.t1544 215.518
R739 VDD.n486 VDD.t1819 215.518
R740 VDD.n477 VDD.t1177 215.518
R741 VDD.n462 VDD.t1808 215.518
R742 VDD.n577 VDD.t1005 215.518
R743 VDD.n583 VDD.t2067 215.518
R744 VDD.n1330 VDD.t1911 215.518
R745 VDD.n1314 VDD.t849 215.518
R746 VDD.n1315 VDD.t1011 215.518
R747 VDD.n1286 VDD.t1214 215.518
R748 VDD.n1222 VDD.t1163 215.518
R749 VDD.n735 VDD.t507 212.947
R750 VDD.n330 VDD.t335 212.947
R751 VDD.t420 VDD.n557 212.947
R752 VDD.n1321 VDD.t800 212.947
R753 VDD.t2154 VDD.n1280 212.947
R754 VDD.n1234 VDD.t248 212.947
R755 VDD.n1205 VDD.t1558 212.585
R756 VDD.n1216 VDD.t1876 212.585
R757 VDD.n1308 VDD.t819 212.585
R758 VDD.t957 VDD.n1299 212.585
R759 VDD.n743 VDD.t975 212.585
R760 VDD.n734 VDD.t851 212.585
R761 VDD.n306 VDD.t1664 212.585
R762 VDD.n317 VDD.t1514 212.585
R763 VDD.n338 VDD.t1510 212.585
R764 VDD.n339 VDD.t1421 212.585
R765 VDD.n329 VDD.t1662 212.585
R766 VDD.t871 VDD.n366 212.585
R767 VDD.n375 VDD.t2100 212.585
R768 VDD.n551 VDD.t825 212.585
R769 VDD.n558 VDD.t2102 212.585
R770 VDD.n571 VDD.t1902 212.585
R771 VDD.n582 VDD.t1496 212.585
R772 VDD.n1329 VDD.t1492 212.585
R773 VDD.n1320 VDD.t1909 212.585
R774 VDD.n1274 VDD.t965 212.585
R775 VDD.t823 VDD.n1285 212.585
R776 VDD.n1242 VDD.t1882 212.585
R777 VDD.n1243 VDD.t1564 212.585
R778 VDD.n1233 VDD.t1572 212.585
R779 VDD.t1477 VDD.t745 211.974
R780 VDD.t742 VDD.t121 211.974
R781 VDD.t2069 VDD.t739 211.974
R782 VDD.t124 VDD.t306 211.974
R783 VDD.t1649 VDD.t2147 211.974
R784 VDD.t1637 VDD.t313 211.974
R785 VDD.t1873 VDD.t478 211.974
R786 VDD.t467 VDD.t650 211.974
R787 VDD.t764 VDD.t1418 211.974
R788 VDD.t1617 VDD.t699 211.974
R789 VDD.t546 VDD.t547 209.101
R790 VDD.t547 VDD.t804 209.101
R791 VDD.t804 VDD.t802 209.101
R792 VDD.t373 VDD.t372 209.101
R793 VDD.t325 VDD.t373 209.101
R794 VDD.t323 VDD.t325 209.101
R795 VDD.t654 VDD.t653 209.101
R796 VDD.t653 VDD.t304 209.101
R797 VDD.t304 VDD.t302 209.101
R798 VDD.t406 VDD.t405 209.101
R799 VDD.t432 VDD.t406 209.101
R800 VDD.t434 VDD.t432 209.101
R801 VDD.t107 VDD.t108 209.101
R802 VDD.t108 VDD.t175 209.101
R803 VDD.t175 VDD.t173 209.101
R804 VDD.t422 VDD.t423 209.101
R805 VDD.t5 VDD.t422 209.101
R806 VDD.t3 VDD.t5 209.101
R807 VDD.t408 VDD.t407 209.101
R808 VDD.t407 VDD.t140 209.101
R809 VDD.t140 VDD.t138 209.101
R810 VDD.t1 VDD.t580 209.101
R811 VDD.t2167 VDD.t358 209.101
R812 VDD.t561 VDD.t560 209.101
R813 VDD.t1633 VDD.t561 209.101
R814 VDD.t1635 VDD.t1633 209.101
R815 VDD.t109 VDD.t110 209.101
R816 VDD.t110 VDD.t22 209.101
R817 VDD.t22 VDD.t24 209.101
R818 VDD.t563 VDD.t562 209.101
R819 VDD.t1243 VDD.t563 209.101
R820 VDD.t1249 VDD.t1243 209.101
R821 VDD.t774 VDD.t773 209.101
R822 VDD.t773 VDD.t767 209.101
R823 VDD.t767 VDD.t769 209.101
R824 VDD.t734 VDD.t735 209.101
R825 VDD.t298 VDD.t734 209.101
R826 VDD.t300 VDD.t298 209.101
R827 VDD.t1620 VDD.t1621 209.101
R828 VDD.t1621 VDD.t600 209.101
R829 VDD.t600 VDD.t598 209.101
R830 VDD.t548 VDD.t549 209.101
R831 VDD.t238 VDD.t548 209.101
R832 VDD.t236 VDD.t238 209.101
R833 VDD.n722 VDD.t973 205.751
R834 VDD.t1927 VDD.t1925 204.739
R835 VDD.t1923 VDD.t1927 204.739
R836 VDD.t1273 VDD.t1275 204.739
R837 VDD.t1275 VDD.t1277 204.739
R838 VDD.t1409 VDD.t1411 204.739
R839 VDD.t1411 VDD.t1413 204.739
R840 VDD.t1271 VDD.t1269 204.739
R841 VDD.t1265 VDD.t1271 204.739
R842 VDD.t994 VDD.t996 204.739
R843 VDD.t996 VDD.t998 204.739
R844 VDD.t1267 VDD.t1279 204.739
R845 VDD.t1279 VDD.t1281 204.739
R846 VDD.n978 VDD.t102 202.248
R847 VDD.n1008 VDD.t1622 200.87
R848 VDD.t1991 VDD.t1990 196.721
R849 VDD.n1009 VDD.t331 195.971
R850 VDD.t1622 VDD.t1627 187.827
R851 VDD.t1627 VDD.t1624 187.827
R852 VDD.t1624 VDD.t2120 187.827
R853 VDD.t2122 VDD.t2121 187.827
R854 VDD.t657 VDD.t655 187.827
R855 VDD.t655 VDD.t991 187.827
R856 VDD.t311 VDD.t659 187.827
R857 VDD.t719 VDD.t660 187.827
R858 VDD.t17 VDD.t15 187.827
R859 VDD.t917 VDD.t18 187.827
R860 VDD.t458 VDD.t61 187.827
R861 VDD.t460 VDD.t458 187.827
R862 VDD.t1199 VDD.t1193 187.827
R863 VDD.t1194 VDD.t1603 187.827
R864 VDD.t1603 VDD.t1195 187.827
R865 VDD.t1195 VDD.t1197 187.827
R866 VDD.t527 VDD.t531 187.827
R867 VDD.t529 VDD.t527 187.827
R868 VDD.t671 VDD.t127 187.827
R869 VDD.n111 VDD.t1340 187.702
R870 VDD.n127 VDD.t1351 187.702
R871 VDD.n1492 VDD.t1342 187.702
R872 VDD.t1748 VDD.n1628 187.702
R873 VDD.n1660 VDD.t1710 187.702
R874 VDD.t1746 VDD.n1642 187.702
R875 VDD.n1667 VDD.t1704 187.702
R876 VDD.n687 VDD.t1036 187.702
R877 VDD.n676 VDD.t1066 187.702
R878 VDD.n1263 VDD.t1778 187.702
R879 VDD.t285 VDD.t287 187.663
R880 VDD.t1595 VDD.t1596 187.663
R881 VDD.n1605 VDD.t2120 185.218
R882 VDD.n1507 VDD.t1194 185.218
R883 VDD.n144 VDD.t779 184.579
R884 VDD.t129 VDD.n703 180.87
R885 VDD.n1007 VDD.t333 178.809
R886 VDD.n145 VDD.t183 168.343
R887 VDD.n1176 VDD.t130 167.827
R888 VDD.n1685 VDD.t1265 164.929
R889 VDD.t384 VDD.t386 163.389
R890 VDD.t1446 VDD.t384 163.389
R891 VDD.t1449 VDD.t1446 163.389
R892 VDD.t266 VDD.t1449 163.389
R893 VDD.t264 VDD.t266 163.389
R894 VDD.t1591 VDD.t1593 163.266
R895 VDD.t48 VDD.t1591 163.266
R896 VDD.t52 VDD.t48 163.266
R897 VDD.t73 VDD.t52 163.266
R898 VDD.t71 VDD.t73 163.266
R899 VDD.t33 VDD.t35 163.266
R900 VDD.t35 VDD.t1698 163.266
R901 VDD.t1698 VDD.t1700 163.266
R902 VDD.t1700 VDD.t26 163.266
R903 VDD.t26 VDD.t28 163.266
R904 VDD.n1010 VDD.n1009 157.51
R905 VDD.n1570 VDD.t1306 157.338
R906 VDD.t258 VDD.n1211 156.898
R907 VDD.n1217 VDD.t1155 156.898
R908 VDD.n1307 VDD.t792 156.898
R909 VDD.n1291 VDD.t1459 156.898
R910 VDD.n1370 VDD.t1671 156.898
R911 VDD.t1855 VDD.n1364 156.898
R912 VDD.n1365 VDD.t2072 156.898
R913 VDD.n1357 VDD.t1247 156.898
R914 VDD.t2038 VDD.n1360 156.898
R915 VDD.n249 VDD.t1387 156.898
R916 VDD.n1375 VDD.t2139 156.898
R917 VDD.n1382 VDD.t1444 156.898
R918 VDD.n1381 VDD.t1789 156.898
R919 VDD.n1394 VDD.t1992 156.898
R920 VDD.n1388 VDD.t1957 156.898
R921 VDD.n1401 VDD.t1534 156.898
R922 VDD.n1400 VDD.t1831 156.898
R923 VDD.n1407 VDD.t1185 156.898
R924 VDD.n744 VDD.t905 156.898
R925 VDD.n728 VDD.t951 156.898
R926 VDD.t1259 VDD.n760 156.898
R927 VDD.n723 VDD.t1261 156.898
R928 VDD.t391 VDD.n312 156.898
R929 VDD.n318 VDD.t1945 156.898
R930 VDD.n323 VDD.t1986 156.898
R931 VDD.n358 VDD.t1979 156.898
R932 VDD.n374 VDD.t2114 156.898
R933 VDD.n550 VDD.t865 156.898
R934 VDD.n285 VDD.t1482 156.898
R935 VDD.n521 VDD.t1686 156.898
R936 VDD.n527 VDD.t1845 156.898
R937 VDD.n526 VDD.t2090 156.898
R938 VDD.n534 VDD.t1236 156.898
R939 VDD.n531 VDD.t2056 156.898
R940 VDD.t1407 VDD.n404 156.898
R941 VDD.n516 VDD.t2128 156.898
R942 VDD.t1434 VDD.n508 156.898
R943 VDD.n509 VDD.t2034 156.898
R944 VDD.n493 VDD.t2010 156.898
R945 VDD.t1967 VDD.n500 156.898
R946 VDD.t1522 VDD.n485 156.898
R947 VDD.n486 VDD.t1827 156.898
R948 VDD.t1181 VDD.n477 156.898
R949 VDD.n462 VDD.t1782 156.898
R950 VDD.t1003 VDD.n577 156.898
R951 VDD.n583 VDD.t2062 156.898
R952 VDD.n1330 VDD.t817 156.898
R953 VDD.t815 VDD.n1314 156.898
R954 VDD.n1315 VDD.t1013 156.898
R955 VDD.n1286 VDD.t1212 156.898
R956 VDD.n1222 VDD.t1165 156.898
R957 VDD.t1201 VDD.t1202 156.409
R958 VDD.t708 VDD.t942 156.409
R959 VDD.n735 VDD.t503 155.026
R960 VDD.n330 VDD.t341 155.026
R961 VDD.n557 VDD.t418 155.026
R962 VDD.n1321 VDD.t796 155.026
R963 VDD.n1280 VDD.t2156 155.026
R964 VDD.n1234 VDD.t252 155.026
R965 VDD.n1205 VDD.t1566 154.762
R966 VDD.t1880 VDD.n1216 154.762
R967 VDD.n1308 VDD.t873 154.762
R968 VDD.n1299 VDD.t959 154.762
R969 VDD.t979 VDD.n743 154.762
R970 VDD.t899 VDD.n734 154.762
R971 VDD.t971 VDD.n722 154.762
R972 VDD.n306 VDD.t1652 154.762
R973 VDD.t1508 VDD.n317 154.762
R974 VDD.t1512 VDD.n338 154.762
R975 VDD.n339 VDD.t1658 154.762
R976 VDD.t1425 VDD.n329 154.762
R977 VDD.n366 VDD.t829 154.762
R978 VDD.n375 VDD.t2110 154.762
R979 VDD.n551 VDD.t847 154.762
R980 VDD.n558 VDD.t2098 154.762
R981 VDD.n571 VDD.t877 154.762
R982 VDD.t1490 VDD.n582 154.762
R983 VDD.t1498 VDD.n1329 154.762
R984 VDD.t1896 VDD.n1320 154.762
R985 VDD.n1274 VDD.t1892 154.762
R986 VDD.n1285 VDD.t833 154.762
R987 VDD.t1886 VDD.n1242 154.762
R988 VDD.n1243 VDD.t1574 154.762
R989 VDD.t1576 VDD.n1233 154.762
R990 VDD.n1171 VDD.t1204 154.237
R991 VDD.n1044 VDD.t571 147.94
R992 VDD.n110 VDD.t221 145.662
R993 VDD.t1220 VDD.n56 145.662
R994 VDD.t806 VDD.n1661 145.662
R995 VDD.t410 VDD.n1668 145.662
R996 VDD.t426 VDD.n688 145.662
R997 VDD.t113 VDD.n677 145.662
R998 VDD.n1262 VDD.t610 145.662
R999 VDD.t540 VDD.n1044 144.69
R1000 VDD.t1204 VDD.t529 144.565
R1001 VDD.n1165 VDD.t1230 137.524
R1002 VDD.t204 VDD.t775 136.796
R1003 VDD.t221 VDD.t223 136.796
R1004 VDD.t44 VDD.t1220 136.796
R1005 VDD.t43 VDD.t45 136.796
R1006 VDD.t425 VDD.t369 136.796
R1007 VDD.t424 VDD.t806 136.796
R1008 VDD.t347 VDD.t349 136.796
R1009 VDD.t348 VDD.t410 136.796
R1010 VDD.t429 VDD.t426 136.796
R1011 VDD.t666 VDD.t475 136.796
R1012 VDD.t111 VDD.t113 136.796
R1013 VDD.t188 VDD.t189 136.796
R1014 VDD.t1981 VDD.t688 136.796
R1015 VDD.t1468 VDD.t1464 136.796
R1016 VDD.t400 VDD.t381 136.796
R1017 VDD.t610 VDD.t399 136.796
R1018 VDD.n772 VDD.t1991 133.881
R1019 VDD.n1675 VDD.t1302 132.998
R1020 VDD.n1569 VDD.t1325 131.619
R1021 VDD.t775 VDD.n126 122.23
R1022 VDD.n1629 VDD.t43 122.23
R1023 VDD.n1662 VDD.t425 122.23
R1024 VDD.n1669 VDD.t347 122.23
R1025 VDD.n689 VDD.t666 122.23
R1026 VDD.n678 VDD.t188 122.23
R1027 VDD.n344 VDD.t1981 122.23
R1028 VDD.n1261 VDD.t400 122.23
R1029 VDD.n1170 VDD.t1532 118.397
R1030 VDD.t1841 VDD.t1670 116.947
R1031 VDD.t1841 VDD.t1227 116.947
R1032 VDD.t121 VDD.n1350 115.8
R1033 VDD.n1351 VDD.t124 115.8
R1034 VDD.n762 VDD.t1637 115.8
R1035 VDD.n541 VDD.t467 115.8
R1036 VDD.n540 VDD.t1617 115.8
R1037 VDD.t686 VDD.t684 112.15
R1038 VDD.t578 VDD.t576 112.091
R1039 VDD.t584 VDD.t582 112.091
R1040 VDD.t278 VDD.t276 112.091
R1041 VDD.t684 VDD.t1864 110.593
R1042 VDD.t68 VDD.t147 110.593
R1043 VDD.t66 VDD.t145 110.593
R1044 VDD.t620 VDD.t602 110.535
R1045 VDD.t618 VDD.t604 110.535
R1046 VDD.t50 VDD.t578 110.535
R1047 VDD.t276 VDD.t1696 110.535
R1048 VDD.t272 VDD.t1869 110.535
R1049 VDD.t274 VDD.t1871 110.535
R1050 VDD.t706 VDD.n1170 110.066
R1051 VDD.n1588 VDD.t2023 107.48
R1052 VDD.n1616 VDD.t202 107.424
R1053 VDD.n1063 VDD.t2163 107.424
R1054 VDD.n68 VDD.t1 104.55
R1055 VDD.n961 VDD.t2167 104.55
R1056 VDD.n623 VDD.t680 102.993
R1057 VDD.n898 VDD.n897 102.832
R1058 VDD.n885 VDD.t1085 99.7607
R1059 VDD.n1099 VDD.t1046 99.7607
R1060 VDD.t2025 VDD.t240 99.1698
R1061 VDD.t525 VDD.t197 99.1183
R1062 VDD.t2162 VDD.t1645 99.1183
R1063 VDD.t75 VDD.t77 96.5152
R1064 VDD.n1350 VDD.t1477 96.1732
R1065 VDD.n1351 VDD.t2069 96.1732
R1066 VDD.n762 VDD.t1649 96.1732
R1067 VDD.n541 VDD.t1873 96.1732
R1068 VDD.t1418 VDD.n540 96.1732
R1069 VDD.n1676 VDD.t497 95.9601
R1070 VDD.t502 VDD.t671 95.9138
R1071 VDD.n1169 VDD.n773 94.7182
R1072 VDD.t659 VDD.n1604 93.9135
R1073 VDD.t15 VDD.n1506 93.9135
R1074 VDD.t1596 VDD.n1471 93.832
R1075 VDD.t2023 VDD.t436 93.6286
R1076 VDD.t448 VDD.t202 93.588
R1077 VDD.t2163 VDD.t156 93.588
R1078 VDD.t1371 VDD.t441 92.3282
R1079 VDD.t200 VDD.t1060 92.2882
R1080 VDD.t1032 VDD.t154 92.2882
R1081 VDD.t973 VDD.t981 89.7015
R1082 VDD.t86 VDD.t2064 89.7015
R1083 VDD.n146 VDD.t456 89.2584
R1084 VDD.t31 VDD.n1185 87.6251
R1085 VDD.n1525 VDD.t404 86.263
R1086 VDD.t631 VDD.t402 86.2625
R1087 VDD.t1028 VDD.n917 83.4537
R1088 VDD.n1098 VDD.t1095 83.4537
R1089 VDD.n622 VDD.t678 83.4297
R1090 VDD.t32 VDD.t1457 81.8111
R1091 VDD.n1186 VDD.t2064 80.15
R1092 VDD.n1170 VDD.t1530 78.3247
R1093 VDD.t1087 VDD.n1028 76.9236
R1094 VDD.n1026 VDD.t1145 76.9236
R1095 VDD.t231 VDD.n952 74.7415
R1096 VDD.t76 VDD.t80 74.741
R1097 VDD.t40 VDD.t37 74.741
R1098 VDD.n1587 VDD.t438 74.1227
R1099 VDD.t198 VDD.n896 74.0906
R1100 VDD.n1062 VDD.t152 74.0906
R1101 VDD.n1604 VDD.n1603 73.9135
R1102 VDD.n1506 VDD.n1505 73.9135
R1103 VDD.n1471 VDD.n1470 73.8493
R1104 VDD.n1177 VDD.t502 73.3638
R1105 VDD.n1690 VDD.t1273 71.0905
R1106 VDD.n1689 VDD.t1269 71.0905
R1107 VDD.n1684 VDD.t1267 71.0905
R1108 VDD.t2130 VDD.t2168 65.6005
R1109 VDD.t2131 VDD.t2169 65.6005
R1110 VDD.t1429 VDD.t354 65.6005
R1111 VDD.t1673 VDD.n1169 63.7528
R1112 VDD.n978 VDD.n977 63.1204
R1113 VDD.n1527 VDD.n1526 63.1204
R1114 VDD.n951 VDD.n950 63.1204
R1115 VDD.t1532 VDD.n772 62.842
R1116 VDD.n1165 VDD.t1841 59.199
R1117 VDD.t2147 VDD.n761 56.919
R1118 VDD.t2 VDD.n68 56.0462
R1119 VDD.n1183 VDD.t1040 55.2364
R1120 VDD.n146 VDD.t455 54.121
R1121 VDD.t682 VDD.n1183 52.3595
R1122 VDD.t2168 VDD.t2131 49.6005
R1123 VDD.t356 VDD.t1429 49.6005
R1124 VDD.n898 VDD.t75 47.811
R1125 VDD.n1170 VDD.t708 46.3437
R1126 VDD.n962 VDD.n961 45.3338
R1127 VDD.n111 VDD.t1329 45.3079
R1128 VDD.n127 VDD.t1319 45.3079
R1129 VDD.t1331 VDD.n1492 45.3079
R1130 VDD.n1628 VDD.t1722 45.3079
R1131 VDD.t1756 VDD.n1660 45.3079
R1132 VDD.n1642 VDD.t1768 45.3079
R1133 VDD.t1739 VDD.n1667 45.3079
R1134 VDD.t1083 VDD.n687 45.3079
R1135 VDD.t1104 VDD.n676 45.3079
R1136 VDD.n1263 VDD.t1784 45.3079
R1137 VDD.n1353 VDD 44.41
R1138 VDD VDD.n538 44.41
R1139 VDD.n1615 VDD.n68 44.1105
R1140 VDD.n1527 VDD.n1525 43.132
R1141 VDD.n1043 VDD.t691 42.125
R1142 VDD.n1010 VDD.t646 42.125
R1143 VDD.n144 VDD.t457 40.9969
R1144 VDD.n144 VDD.t0 40.9969
R1145 VDD.n145 VDD.t181 38.9615
R1146 VDD.t1841 VDD.n773 38.2519
R1147 VDD.n952 VDD.n951 37.3712
R1148 VDD.n1164 VDD.t1438 36.8005
R1149 VDD.n1528 VDD.n1527 33.9467
R1150 VDD.t1306 VDD.n1569 31.7705
R1151 VDD.t457 VDD.t2 30.0991
R1152 VDD.t0 VDD.t456 30.0991
R1153 VDD.n900 VDD.n899 29.4128
R1154 VDD.n951 VDD.n926 29.4128
R1155 VDD.t2121 VDD.t657 24.3483
R1156 VDD.t1193 VDD.t460 24.3483
R1157 VDD.t1069 VDD.n622 24.1662
R1158 VDD.n1494 VDD.n1491 20.3263
R1159 VDD.n1347 VDD.t213 20.2823
R1160 VDD.n1334 VDD.t219 20.2823
R1161 VDD.n394 VDD.t216 20.2823
R1162 VDD.n545 VDD.t207 20.2823
R1163 VDD.n749 VDD.t210 20.2775
R1164 VDD.t1202 VDD.t706 20.2757
R1165 VDD.n917 VDD.t1085 20.1444
R1166 VDD.t1046 VDD.n1098 20.1444
R1167 VDD.n1603 VDD.t660 20.0005
R1168 VDD.n1505 VDD.t18 20.0005
R1169 VDD.t127 VDD.n1176 20.0005
R1170 VDD.n1470 VDD.t285 19.9831
R1171 VDD.n1100 VDD.n845 19.8305
R1172 VDD.n916 VDD.n848 19.8305
R1173 VDD.n1030 VDD.n993 19.8305
R1174 VDD.n1025 VDD.n994 19.8305
R1175 VDD.n624 VDD.n621 19.8305
R1176 VDD.n1571 VDD.n1542 19.5344
R1177 VDD.n148 VDD.n147 18.2775
R1178 VDD.t1308 VDD.n1587 18.206
R1179 VDD.n896 VDD.t1044 18.1981
R1180 VDD.t1091 VDD.n1062 18.1981
R1181 VDD.t678 VDD.t1040 16.6863
R1182 VDD.t680 VDD.t1069 16.6863
R1183 VDD.n220 VDD.t1675 15.8102
R1184 VDD.n429 VDD.t1689 15.8102
R1185 VDD.n1681 VDD.n1680 15.6843
R1186 VDD.n1674 VDD.n29 15.4714
R1187 VDD.n1312 VDD.n1311 15.2273
R1188 VDD.n1029 VDD.t1107 14.6525
R1189 VDD.t1026 VDD.n1006 14.6525
R1190 VDD.n126 VDD.t223 14.5667
R1191 VDD.n1629 VDD.t44 14.5667
R1192 VDD.n1662 VDD.t424 14.5667
R1193 VDD.n1669 VDD.t348 14.5667
R1194 VDD.n689 VDD.t429 14.5667
R1195 VDD.n678 VDD.t111 14.5667
R1196 VDD.n344 VDD.t1468 14.5667
R1197 VDD.t399 VDD.n1261 14.5667
R1198 VDD.n747 VDD.n746 13.9985
R1199 VDD.n969 VDD.t595 13.8991
R1200 VDD.n132 VDD.t146 13.8991
R1201 VDD.n80 VDD.t658 13.8991
R1202 VDD.n65 VDD.t621 13.8991
R1203 VDD.n154 VDD.t461 13.8991
R1204 VDD.n934 VDD.t1872 13.8991
R1205 VDD.n643 VDD.t707 13.8991
R1206 VDD.n1456 VDD.n157 13.6237
R1207 VDD.n1457 VDD.n134 13.5005
R1208 VDD.n1459 VDD.n1458 13.5005
R1209 VDD.n991 VDD.n175 13.5005
R1210 VDD.n1102 VDD.n1101 13.5005
R1211 VDD.n1415 VDD.n1414 13.5005
R1212 VDD.n1677 VDD.t499 13.4685
R1213 VDD.t242 VDD.t2025 12.9808
R1214 VDD.t240 VDD.t2026 12.9808
R1215 VDD.t203 VDD.t525 12.974
R1216 VDD.t197 VDD.t523 12.974
R1217 VDD.t1647 VDD.t2162 12.974
R1218 VDD.t1645 VDD.t2164 12.974
R1219 VDD.t2169 VDD.n1164 12.8005
R1220 VDD.n1218 VDD.n1217 12.6005
R1221 VDD.n1216 VDD.n1215 12.6005
R1222 VDD VDD.n1212 12.6005
R1223 VDD.n1211 VDD.n1210 12.6005
R1224 VDD.n1206 VDD.n1205 12.6005
R1225 VDD.n1292 VDD.n1291 12.6005
R1226 VDD.n1299 VDD.n1298 12.6005
R1227 VDD VDD.n1300 12.6005
R1228 VDD.n1307 VDD.n1306 12.6005
R1229 VDD.n1309 VDD.n1308 12.6005
R1230 VDD.n1583 VDD.n1582 12.6005
R1231 VDD.n1582 VDD.n1581 12.6005
R1232 VDD.n126 VDD.n125 12.6005
R1233 VDD.n1603 VDD.n1602 12.6005
R1234 VDD.n1043 VDD.n1042 12.6005
R1235 VDD.n1011 VDD.n1010 12.6005
R1236 VDD.n901 VDD.n884 12.6005
R1237 VDD.n902 VDD.n901 12.6005
R1238 VDD.n1615 VDD.n1614 12.6005
R1239 VDD.n1505 VDD.n1504 12.6005
R1240 VDD.n1470 VDD.n1469 12.6005
R1241 VDD.n1630 VDD.n1629 12.6005
R1242 VDD.n1663 VDD.n1662 12.6005
R1243 VDD VDD.n1685 12.6005
R1244 VDD.n1684 VDD.n1683 12.6005
R1245 VDD.n1670 VDD.n1669 12.6005
R1246 VDD.n729 VDD.n728 12.6005
R1247 VDD.n734 VDD.n733 12.6005
R1248 VDD.n736 VDD.n735 12.6005
R1249 VDD.n743 VDD.n742 12.6005
R1250 VDD.n745 VDD.n744 12.6005
R1251 VDD.n760 VDD.n759 12.6005
R1252 VDD.n690 VDD.n689 12.6005
R1253 VDD.n679 VDD.n678 12.6005
R1254 VDD.n724 VDD.n723 12.6005
R1255 VDD.n722 VDD.n721 12.6005
R1256 VDD.n1187 VDD.n1186 12.6005
R1257 VDD.n1183 VDD.n1182 12.6005
R1258 VDD.n1176 VDD.n1175 12.6005
R1259 VDD.n772 VDD.n771 12.6005
R1260 VDD.n1083 VDD.n1082 12.6005
R1261 VDD.n1084 VDD.n1083 12.6005
R1262 VDD.n963 VDD.n962 12.6005
R1263 VDD.n1164 VDD 12.6005
R1264 VDD.n1408 VDD.n1407 12.6005
R1265 VDD.n1402 VDD.n1401 12.6005
R1266 VDD.n1400 VDD.n1399 12.6005
R1267 VDD.n1394 VDD.n1393 12.6005
R1268 VDD.n1389 VDD.n1388 12.6005
R1269 VDD.n1383 VDD.n1382 12.6005
R1270 VDD.n1381 VDD.n1380 12.6005
R1271 VDD.n1375 VDD.n1374 12.6005
R1272 VDD.n250 VDD.n249 12.6005
R1273 VDD.n1358 VDD.n1357 12.6005
R1274 VDD.n1360 VDD.n1359 12.6005
R1275 VDD.n1364 VDD.n1363 12.6005
R1276 VDD.n1366 VDD.n1365 12.6005
R1277 VDD.n1371 VDD.n1370 12.6005
R1278 VDD.n338 VDD.n337 12.6005
R1279 VDD.n340 VDD.n339 12.6005
R1280 VDD.n331 VDD.n330 12.6005
R1281 VDD.n329 VDD.n328 12.6005
R1282 VDD.n324 VDD.n323 12.6005
R1283 VDD.n319 VDD.n318 12.6005
R1284 VDD.n317 VDD.n316 12.6005
R1285 VDD VDD.n313 12.6005
R1286 VDD.n312 VDD.n311 12.6005
R1287 VDD.n307 VDD.n306 12.6005
R1288 VDD.n345 VDD.n344 12.6005
R1289 VDD.n559 VDD.n558 12.6005
R1290 VDD.n557 VDD.n556 12.6005
R1291 VDD.n552 VDD.n551 12.6005
R1292 VDD.n550 VDD.n549 12.6005
R1293 VDD.n463 VDD.n462 12.6005
R1294 VDD.n477 VDD.n476 12.6005
R1295 VDD.n485 VDD.n484 12.6005
R1296 VDD.n487 VDD.n486 12.6005
R1297 VDD.n494 VDD.n493 12.6005
R1298 VDD.n500 VDD.n499 12.6005
R1299 VDD.n508 VDD.n507 12.6005
R1300 VDD.n510 VDD.n509 12.6005
R1301 VDD.n517 VDD.n516 12.6005
R1302 VDD.n404 VDD.n403 12.6005
R1303 VDD.n534 VDD.n533 12.6005
R1304 VDD.n532 VDD.n531 12.6005
R1305 VDD.n528 VDD.n527 12.6005
R1306 VDD.n526 VDD.n525 12.6005
R1307 VDD.n521 VDD.n520 12.6005
R1308 VDD.n376 VDD.n375 12.6005
R1309 VDD.n374 VDD.n373 12.6005
R1310 VDD VDD.n367 12.6005
R1311 VDD.n366 VDD.n365 12.6005
R1312 VDD.n359 VDD.n358 12.6005
R1313 VDD.n286 VDD.n285 12.6005
R1314 VDD.n584 VDD.n583 12.6005
R1315 VDD.n582 VDD.n581 12.6005
R1316 VDD VDD.n578 12.6005
R1317 VDD.n577 VDD.n576 12.6005
R1318 VDD.n572 VDD.n571 12.6005
R1319 VDD.n1331 VDD.n1330 12.6005
R1320 VDD.n1329 VDD.n1328 12.6005
R1321 VDD.n1322 VDD.n1321 12.6005
R1322 VDD.n1320 VDD.n1319 12.6005
R1323 VDD.n1314 VDD.n1313 12.6005
R1324 VDD.n1316 VDD.n1315 12.6005
R1325 VDD.n1275 VDD.n1274 12.6005
R1326 VDD.n1280 VDD.n1279 12.6005
R1327 VDD.n1285 VDD.n1284 12.6005
R1328 VDD.n1287 VDD.n1286 12.6005
R1329 VDD.n1261 VDD.n1260 12.6005
R1330 VDD.n1242 VDD.n1241 12.6005
R1331 VDD.n1244 VDD.n1243 12.6005
R1332 VDD.n1235 VDD.n1234 12.6005
R1333 VDD.n1233 VDD.n1232 12.6005
R1334 VDD.n1223 VDD.n1222 12.6005
R1335 VDD.n1691 VDD.n1690 12.6005
R1336 VDD.n1689 VDD.n1688 12.6005
R1337 VDD.n145 VDD.t185 12.5633
R1338 VDD.n1228 VDD 12.4951
R1339 VDD.n586 VDD.n585 12.4925
R1340 VDD.n563 VDD.n562 12.4772
R1341 VDD.n219 VDD.t1679 12.4261
R1342 VDD.n428 VDD.t1694 12.4261
R1343 VDD.n1290 VDD.n1289 12.2886
R1344 VDD.n962 VDD.t356 12.2672
R1345 VDD.n752 VDD.n750 12.1927
R1346 VDD.n1340 VDD.n1338 12.1927
R1347 VDD.n253 VDD.n251 12.1927
R1348 VDD.n389 VDD.n387 12.1927
R1349 VDD.n381 VDD.n379 12.1927
R1350 VDD.n754 VDD.n753 12.1904
R1351 VDD.n1342 VDD.n1341 12.1904
R1352 VDD.n255 VDD.n254 12.1904
R1353 VDD.n391 VDD.n390 12.1904
R1354 VDD.n383 VDD.n382 12.1904
R1355 VDD.n1678 VDD.n29 12.0423
R1356 VDD.n726 VDD.n725 12.0317
R1357 VDD.n321 VDD.n320 12.0317
R1358 VDD.n1220 VDD.n1219 12.0317
R1359 VDD.t582 VDD.n1615 11.9362
R1360 VDD.n1672 VDD.n1671 11.814
R1361 VDD.n767 VDD.n766 11.5663
R1362 VDD.t1089 VDD.t280 11.3197
R1363 VDD.n226 VDD.t1258 11.2371
R1364 VDD.n407 VDD.t1246 11.2371
R1365 VDD.n342 VDD.n289 10.6839
R1366 VDD.n1333 VDD.n258 10.6839
R1367 VDD.n1093 VDD.n1092 10.5186
R1368 VDD.n1655 VDD.n1654 10.5186
R1369 VDD.n1500 VDD.n1499 10.5186
R1370 VDD.n880 VDD.n879 10.5186
R1371 VDD.n1021 VDD.n1020 10.5186
R1372 VDD.n1037 VDD.n1036 10.5186
R1373 VDD.n120 VDD.n119 10.5186
R1374 VDD.n1577 VDD.n1576 10.5186
R1375 VDD.n1556 VDD.n1555 10.5186
R1376 VDD.n1638 VDD.n1637 10.5186
R1377 VDD.n912 VDD.n911 10.5186
R1378 VDD.n1077 VDD.n1076 10.5186
R1379 VDD.n631 VDD.n630 10.5186
R1380 VDD.n672 VDD.n671 10.5186
R1381 VDD.n1255 VDD.n1254 10.5186
R1382 VDD.n1185 VDD.n1184 10.4172
R1383 VDD.n1053 VDD.n1047 10.3508
R1384 VDD.n1608 VDD.n1607 10.3508
R1385 VDD.n1623 VDD.n1618 10.3508
R1386 VDD.n949 VDD.n948 10.3508
R1387 VDD.n1596 VDD.n1590 10.3503
R1388 VDD.n1515 VDD.n1509 10.3503
R1389 VDD.n702 VDD.n701 10.3503
R1390 VDD.n1289 VDD.n1266 10.1306
R1391 VDD.n45 VDD.n43 10.0135
R1392 VDD.n983 VDD.n981 10.0135
R1393 VDD.n1523 VDD.n1521 10.0135
R1394 VDD.n1539 VDD.n1537 10.0135
R1395 VDD.n91 VDD.n89 10.0135
R1396 VDD.n103 VDD.n101 10.0135
R1397 VDD.n1003 VDD.n1001 10.0135
R1398 VDD.n71 VDD.n69 10.0135
R1399 VDD.n1462 VDD.n1460 10.0135
R1400 VDD.n55 VDD.n53 10.0135
R1401 VDD.n857 VDD.n855 10.0135
R1402 VDD.n868 VDD.n866 10.0135
R1403 VDD.n142 VDD.n140 10.0135
R1404 VDD.n1482 VDD.n1480 10.0135
R1405 VDD.n35 VDD.n33 10.0135
R1406 VDD.n1069 VDD.n1067 10.0135
R1407 VDD.n606 VDD.n604 10.0135
R1408 VDD.n650 VDD.n648 10.0135
R1409 VDD.n656 VDD.n654 10.0135
R1410 VDD.n613 VDD.n611 10.0135
R1411 VDD.n925 VDD.n923 10.0135
R1412 VDD.n960 VDD.n958 10.0135
R1413 VDD.n348 VDD.n346 10.0135
R1414 VDD.n599 VDD.n597 10.0135
R1415 VDD.n1247 VDD.n1246 9.88805
R1416 VDD.n1186 VDD.t1473 9.552
R1417 VDD.n1566 VDD.n1565 9.49544
R1418 VDD.t402 VDD.n1528 9.1863
R1419 VDD.n1163 VDD.n1162 9.0005
R1420 VDD.n1169 VDD.n1168 8.85441
R1421 VDD.n1166 VDD.n774 8.64281
R1422 VDD.n1493 VDD.t1323 8.63049
R1423 VDD.n1373 VDD.n1372 8.42496
R1424 VDD.n519 VDD.n518 8.42496
R1425 VDD.n240 VDD.t1840 8.3042
R1426 VDD.n421 VDD.t1854 8.3042
R1427 VDD.n961 VDD.t1438 8.0005
R1428 VDD.n900 VDD.t76 7.95948
R1429 VDD.n926 VDD.t40 7.95948
R1430 VDD.t1473 VDD.t32 7.89087
R1431 VDD.t1457 VDD.t31 7.89087
R1432 VDD.n266 VDD.t1018 7.64083
R1433 VDD.n1268 VDD.t1211 7.64083
R1434 VDD.n586 VDD.t1016 7.5993
R1435 VDD.n1288 VDD.t1209 7.5993
R1436 VDD.n147 VDD.t183 7.37043
R1437 VDD.n952 VDD.t230 7.25909
R1438 VDD.n547 VDD.n378 7.20693
R1439 VDD.n703 VDD.t130 6.95702
R1440 VDD.n236 VDD.t2087 6.93712
R1441 VDD.n247 VDD.t1400 6.93712
R1442 VDD.n417 VDD.t2079 6.93712
R1443 VDD.n401 VDD.t1390 6.93712
R1444 VDD.n248 VDD.t1396 6.90536
R1445 VDD.n402 VDD.t1386 6.90536
R1446 VDD.n147 VDD.n146 6.72961
R1447 VDD.n1587 VDD.n1586 6.3005
R1448 VDD.n1569 VDD.n1568 6.3005
R1449 VDD VDD.n1571 6.3005
R1450 VDD.n1571 VDD.n1570 6.3005
R1451 VDD.n112 VDD.n111 6.3005
R1452 VDD.n128 VDD.n127 6.3005
R1453 VDD VDD.n1030 6.3005
R1454 VDD.n1030 VDD.n1029 6.3005
R1455 VDD VDD.n994 6.3005
R1456 VDD.n1006 VDD.n994 6.3005
R1457 VDD.n917 VDD.n847 6.3005
R1458 VDD VDD.n848 6.3005
R1459 VDD.n885 VDD.n848 6.3005
R1460 VDD.n896 VDD.n895 6.3005
R1461 VDD VDD.n1494 6.3005
R1462 VDD.n1494 VDD.n1493 6.3005
R1463 VDD.n1628 VDD.n1627 6.3005
R1464 VDD.n1660 VDD.n1659 6.3005
R1465 VDD.n1642 VDD.n1641 6.3005
R1466 VDD.n1667 VDD.n1666 6.3005
R1467 VDD.n29 VDD.n28 6.3005
R1468 VDD.n1676 VDD.n29 6.3005
R1469 VDD.n1679 VDD.n1678 6.3005
R1470 VDD.n1678 VDD.n1677 6.3005
R1471 VDD.n1674 VDD.n1673 6.3005
R1472 VDD.n1675 VDD.n1674 6.3005
R1473 VDD.n676 VDD.n675 6.3005
R1474 VDD.n687 VDD.n686 6.3005
R1475 VDD VDD.n624 6.3005
R1476 VDD.n624 VDD.n623 6.3005
R1477 VDD.n1167 VDD.n1166 6.3005
R1478 VDD.n1166 VDD.n1165 6.3005
R1479 VDD.n774 VDD.n773 6.3005
R1480 VDD VDD.n1100 6.3005
R1481 VDD.n1100 VDD.n1099 6.3005
R1482 VDD.n1098 VDD.n1097 6.3005
R1483 VDD.n1062 VDD.n1061 6.3005
R1484 VDD.n1406 VDD.n1405 6.3005
R1485 VDD.n1396 VDD.n1395 6.3005
R1486 VDD.n1387 VDD.n1386 6.3005
R1487 VDD.n1377 VDD.n1376 6.3005
R1488 VDD.n1356 VDD.n1355 6.3005
R1489 VDD.n1362 VDD.n1361 6.3005
R1490 VDD.n1369 VDD.n1368 6.3005
R1491 VDD.n479 VDD.n478 6.3005
R1492 VDD.n492 VDD.n491 6.3005
R1493 VDD.n502 VDD.n501 6.3005
R1494 VDD.n515 VDD.n514 6.3005
R1495 VDD.n536 VDD.n535 6.3005
R1496 VDD.n530 VDD.n529 6.3005
R1497 VDD.n523 VDD.n522 6.3005
R1498 VDD.n1264 VDD.n1263 6.3005
R1499 VDD.n350 VDD.n349 6.13942
R1500 VDD.n1570 VDD.t1375 6.05194
R1501 VDD.n1349 VDD.n1348 6.03954
R1502 VDD.n542 VDD.n386 6.03954
R1503 VDD.n948 VDD.n947 6.0205
R1504 VDD.n1054 VDD.n1053 6.0205
R1505 VDD.n1609 VDD.n1608 6.0205
R1506 VDD.n1624 VDD.n1623 6.0205
R1507 VDD.n1597 VDD.n1596 6.02
R1508 VDD.n1516 VDD.n1515 6.02
R1509 VDD.n701 VDD.n695 6.02
R1510 VDD.n1246 VDD.n1188 5.7697
R1511 VDD.n1091 VDD.n1090 5.75329
R1512 VDD.n1091 VDD.n1089 5.75329
R1513 VDD.n1653 VDD.n1652 5.75329
R1514 VDD.n1653 VDD.n1651 5.75329
R1515 VDD.n1498 VDD.n1497 5.75329
R1516 VDD.n1498 VDD.n1496 5.75329
R1517 VDD.n878 VDD.n877 5.75329
R1518 VDD.n878 VDD.n876 5.75329
R1519 VDD.n77 VDD.n76 5.75329
R1520 VDD.n77 VDD.n75 5.75329
R1521 VDD.n1575 VDD.n1574 5.75329
R1522 VDD.n1575 VDD.n1573 5.75329
R1523 VDD.n1578 VDD.n1541 5.75329
R1524 VDD.n1578 VDD.n1540 5.75329
R1525 VDD.n1610 VDD.n73 5.75329
R1526 VDD.n1610 VDD.n72 5.75329
R1527 VDD.n1621 VDD.n1620 5.75329
R1528 VDD.n1621 VDD.n1619 5.75329
R1529 VDD.n1636 VDD.n1635 5.75329
R1530 VDD.n1636 VDD.n1634 5.75329
R1531 VDD.n1633 VDD.n52 5.75329
R1532 VDD.n1633 VDD.n51 5.75329
R1533 VDD.n1465 VDD.n1464 5.75329
R1534 VDD.n1465 VDD.n1463 5.75329
R1535 VDD.n881 VDD.n870 5.75329
R1536 VDD.n881 VDD.n869 5.75329
R1537 VDD.n1501 VDD.n1484 5.75329
R1538 VDD.n1501 VDD.n1483 5.75329
R1539 VDD VDD.n1163 5.68269
R1540 VDD.n6 VDD.t1414 5.62158
R1541 VDD.n0 VDD.t1929 5.62158
R1542 VDD.n22 VDD.t999 5.62158
R1543 VDD.n10 VDD.t1278 5.56425
R1544 VDD.n17 VDD.t1266 5.56425
R1545 VDD.n27 VDD.t1282 5.56425
R1546 VDD.n1045 VDD.t573 5.49501
R1547 VDD.n1091 VDD.t362 5.35308
R1548 VDD.n1653 VDD.t607 5.35308
R1549 VDD.n1498 VDD.t135 5.35308
R1550 VDD.n878 VDD.t191 5.35308
R1551 VDD.n77 VDD.t639 5.35308
R1552 VDD.n1575 VDD.t320 5.35308
R1553 VDD.n1621 VDD.t330 5.35308
R1554 VDD.n1636 VDD.t2022 5.35308
R1555 VDD.n357 VDD.n356 5.19063
R1556 VDD.n784 VDD.t2172 5.17246
R1557 VDD.n43 VDD.t808 5.17246
R1558 VDD.n42 VDD.t371 5.17246
R1559 VDD.n979 VDD.t537 5.17246
R1560 VDD.n981 VDD.t696 5.17246
R1561 VDD.n1520 VDD.t592 5.17246
R1562 VDD.n1521 VDD.t630 5.17246
R1563 VDD.n1537 VDD.t931 5.17246
R1564 VDD.n1529 VDD.t750 5.17246
R1565 VDD.n88 VDD.t310 5.17246
R1566 VDD.n89 VDD.t718 5.17246
R1567 VDD.n99 VDD.t206 5.17246
R1568 VDD.n101 VDD.t225 5.17246
R1569 VDD.n1001 VDD.t643 5.17246
R1570 VDD.n1004 VDD.t1616 5.17246
R1571 VDD.n1613 VDD.t168 5.17246
R1572 VDD.n69 VDD.t586 5.17246
R1573 VDD.n1468 VDD.t1600 5.17246
R1574 VDD.n1460 VDD.t284 5.17246
R1575 VDD.n58 VDD.t47 5.17246
R1576 VDD.n53 VDD.t1221 5.17246
R1577 VDD.n855 VDD.t85 5.17246
R1578 VDD.n858 VDD.t444 5.17246
R1579 VDD.n887 VDD.t78 5.17246
R1580 VDD.n866 VDD.t293 5.17246
R1581 VDD.n143 VDD.t780 5.17246
R1582 VDD.n140 VDD.t182 5.17246
R1583 VDD.n1480 VDD.t921 5.17246
R1584 VDD.n1472 VDD.t21 5.17246
R1585 VDD.n33 VDD.t413 5.17246
R1586 VDD.n32 VDD.t771 5.17246
R1587 VDD.n927 VDD.t235 5.17246
R1588 VDD.n1067 VDD.t96 5.17246
R1589 VDD.n775 VDD.t1242 5.17246
R1590 VDD.n604 VDD.t1475 5.17246
R1591 VDD.n603 VDD.t88 5.17246
R1592 VDD.n648 VDD.t427 5.17246
R1593 VDD.n651 VDD.t477 5.17246
R1594 VDD.n654 VDD.t116 5.17246
R1595 VDD.n653 VDD.t474 5.17246
R1596 VDD.n636 VDD.t132 5.17246
R1597 VDD.n611 VDD.t675 5.17246
R1598 VDD.n923 VDD.t39 5.17246
R1599 VDD.n1058 VDD.t623 5.17246
R1600 VDD.n958 VDD.t359 5.17246
R1601 VDD.n288 VDD.t689 5.17246
R1602 VDD.n346 VDD.t1476 5.17246
R1603 VDD.n597 VDD.t614 5.17246
R1604 VDD.n596 VDD.t383 5.17246
R1605 VDD.n766 VDD.n748 5.16309
R1606 VDD.n758 VDD.t1295 5.155
R1607 VDD.n461 VDD.t1794 5.155
R1608 VDD.n938 VDD.t344 5.10487
R1609 VDD.n1512 VDD.t726 5.10487
R1610 VDD.n1018 VDD.t785 5.10487
R1611 VDD.n1034 VDD.t637 5.10487
R1612 VDD.n1050 VDD.t377 5.10487
R1613 VDD.n117 VDD.t2159 5.10487
R1614 VDD.n1593 VDD.t1551 5.10487
R1615 VDD.n1553 VDD.t56 5.10487
R1616 VDD.n909 VDD.t452 5.10487
R1617 VDD.n1074 VDD.t351 5.10487
R1618 VDD.n628 VDD.t555 5.10487
R1619 VDD.n698 VDD.t663 5.10487
R1620 VDD.n669 VDD.t295 5.10487
R1621 VDD.n178 VDD.t164 5.10487
R1622 VDD.n1252 VDD.t924 5.10487
R1623 VDD.n766 VDD.n765 5.07929
R1624 VDD.n1270 VDD.t2151 5.01686
R1625 VDD.n711 VDD.t510 5.01686
R1626 VDD.n294 VDD.t338 5.01686
R1627 VDD.n263 VDD.t799 5.01686
R1628 VDD.n1193 VDD.t251 5.01686
R1629 VDD VDD.t1895 5.00492
R1630 VDD VDD.t1661 5.00492
R1631 VDD VDD.t822 5.00492
R1632 VDD VDD.t886 5.00492
R1633 VDD VDD.t1581 5.00492
R1634 VDD.n272 VDD.t417 4.97139
R1635 VDD VDD.t2107 4.94116
R1636 VDD.n41 VDD.t1773 4.92985
R1637 VDD.n1658 VDD.t1774 4.92985
R1638 VDD.n1489 VDD.t1343 4.92985
R1639 VDD.n990 VDD.t1120 4.92985
R1640 VDD.n1519 VDD.t1355 4.92985
R1641 VDD.n1567 VDD.t1328 4.92985
R1642 VDD.n1563 VDD.t1318 4.92985
R1643 VDD.n97 VDD.t1357 4.92985
R1644 VDD.n109 VDD.t1341 4.92985
R1645 VDD.n995 VDD.t1057 4.92985
R1646 VDD.n47 VDD.t1747 4.92985
R1647 VDD.n57 VDD.t1749 4.92985
R1648 VDD.n849 VDD.t1735 4.92985
R1649 VDD.n886 VDD.t1031 4.92985
R1650 VDD.n846 VDD.t1029 4.92985
R1651 VDD.n843 VDD.t1767 4.92985
R1652 VDD.n658 VDD.t1067 4.92985
R1653 VDD.n652 VDD.t1068 4.92985
R1654 VDD.n609 VDD.t1041 4.92985
R1655 VDD.n1096 VDD.t1096 4.92985
R1656 VDD.n1057 VDD.t1094 4.92985
R1657 VDD.n1265 VDD.t1810 4.92985
R1658 VDD.n1680 VDD.t500 4.83406
R1659 VDD.n1672 VDD.t1297 4.82952
R1660 VDD.n1562 VDD.n1561 4.75289
R1661 VDD.n748 VDD.t1301 4.75175
R1662 VDD.n357 VDD.t1974 4.73491
R1663 VDD.n351 VDD.n350 4.69305
R1664 VDD.n1219 VDD.t1158 4.6676
R1665 VDD.n1290 VDD.t1471 4.6676
R1666 VDD.n725 VDD.t1305 4.6676
R1667 VDD.n320 VDD.t1942 4.6676
R1668 VDD.n585 VDD.t2066 4.6676
R1669 VDD.n1312 VDD.t854 4.65357
R1670 VDD.n746 VDD.t862 4.65357
R1671 VDD.n341 VDD.t1669 4.65357
R1672 VDD.n1332 VDD.t858 4.65357
R1673 VDD.n1245 VDD.t1571 4.65357
R1674 VDD.n548 VDD.t889 4.65233
R1675 VDD.n1199 VDD.t1889 4.65007
R1676 VDD.n1213 VDD.t1891 4.65007
R1677 VDD.n1201 VDD.t257 4.65007
R1678 VDD.n1208 VDD.t261 4.65007
R1679 VDD.n1207 VDD.t1579 4.65007
R1680 VDD.n602 VDD.t1561 4.65007
R1681 VDD.n1295 VDD.t970 4.65007
R1682 VDD.n590 VDD.t964 4.65007
R1683 VDD.n1301 VDD.t789 4.65007
R1684 VDD.n1304 VDD.t787 4.65007
R1685 VDD.n1303 VDD.t895 4.65007
R1686 VDD.n1311 VDD.t840 4.65007
R1687 VDD.n1278 VDD.t2153 4.65007
R1688 VDD.n1273 VDD.t968 4.65007
R1689 VDD.n1277 VDD.t962 4.65007
R1690 VDD.n1272 VDD.t838 4.65007
R1691 VDD.n731 VDD.t812 4.65007
R1692 VDD.n730 VDD.t950 4.65007
R1693 VDD.n726 VDD.t956 4.65007
R1694 VDD.n737 VDD.t506 4.65007
R1695 VDD.n741 VDD.t978 4.65007
R1696 VDD.n738 VDD.t986 4.65007
R1697 VDD.n740 VDD.t814 4.65007
R1698 VDD.n1178 VDD.t887 4.65007
R1699 VDD.n706 VDD.t1703 4.65007
R1700 VDD.n607 VDD.t677 4.65007
R1701 VDD.n1179 VDD.t681 4.65007
R1702 VDD.n717 VDD.t984 4.65007
R1703 VDD.n719 VDD.t982 4.65007
R1704 VDD.n1410 VDD.t1180 4.65007
R1705 VDD.n188 VDD.t1176 4.65007
R1706 VDD.n192 VDD.t1549 4.65007
R1707 VDD.n193 VDD.t1822 4.65007
R1708 VDD.n1398 VDD.t1824 4.65007
R1709 VDD.n1392 VDD.t2006 4.65007
R1710 VDD.n1391 VDD.t1964 4.65007
R1711 VDD.n202 VDD.t1962 4.65007
R1712 VDD.n209 VDD.t1432 4.65007
R1713 VDD.n210 VDD.t1792 4.65007
R1714 VDD.n1379 VDD.t1801 4.65007
R1715 VDD.n1373 VDD.t2145 4.65007
R1716 VDD.n237 VDD.t2089 4.65007
R1717 VDD.n238 VDD.t1838 4.65007
R1718 VDD.n230 VDD.t2051 4.65007
R1719 VDD.n228 VDD.t2059 4.65007
R1720 VDD.n227 VDD.t1256 4.65007
R1721 VDD.n269 VDD.t1481 4.65007
R1722 VDD.n335 VDD.t1667 4.65007
R1723 VDD.n332 VDD.t340 4.65007
R1724 VDD.n336 VDD.t1507 4.65007
R1725 VDD.n333 VDD.t1519 4.65007
R1726 VDD.n326 VDD.t1657 4.65007
R1727 VDD.n325 VDD.t1983 4.65007
R1728 VDD.n321 VDD.t1989 4.65007
R1729 VDD.n300 VDD.t1505 4.65007
R1730 VDD.n314 VDD.t1517 4.65007
R1731 VDD.n302 VDD.t396 4.65007
R1732 VDD.n309 VDD.t394 4.65007
R1733 VDD.n308 VDD.t1424 4.65007
R1734 VDD.n289 VDD.t1655 4.65007
R1735 VDD.n561 VDD.t2097 4.65007
R1736 VDD.n555 VDD.t415 4.65007
R1737 VDD.n276 VDD.t898 4.65007
R1738 VDD.n275 VDD.t1905 4.65007
R1739 VDD.n554 VDD.t1901 4.65007
R1740 VDD.n464 VDD.t1803 4.65007
R1741 VDD.n473 VDD.t1170 4.65007
R1742 VDD.n475 VDD.t1188 4.65007
R1743 VDD.n483 VDD.t1538 4.65007
R1744 VDD.n482 VDD.t1834 4.65007
R1745 VDD.n488 VDD.t1814 4.65007
R1746 VDD.n495 VDD.t1997 4.65007
R1747 VDD.n496 VDD.t1956 4.65007
R1748 VDD.n498 VDD.t1954 4.65007
R1749 VDD.n506 VDD.t1452 4.65007
R1750 VDD.n505 VDD.t2029 4.65007
R1751 VDD.n511 VDD.t2031 4.65007
R1752 VDD.n518 VDD.t2136 4.65007
R1753 VDD.n418 VDD.t2081 4.65007
R1754 VDD.n419 VDD.t1852 4.65007
R1755 VDD.n411 VDD.t2041 4.65007
R1756 VDD.n409 VDD.t2047 4.65007
R1757 VDD.n408 VDD.t1241 4.65007
R1758 VDD.n370 VDD.t2105 4.65007
R1759 VDD.n378 VDD.t2109 4.65007
R1760 VDD.n368 VDD.t2119 4.65007
R1761 VDD.n371 VDD.t2117 4.65007
R1762 VDD.n362 VDD.t902 4.65007
R1763 VDD.n279 VDD.t1899 4.65007
R1764 VDD.n355 VDD.t1487 4.65007
R1765 VDD.n1317 VDD.t864 4.65007
R1766 VDD.n565 VDD.t1503 4.65007
R1767 VDD.n579 VDD.t1489 4.65007
R1768 VDD.n567 VDD.t1008 4.65007
R1769 VDD.n574 VDD.t1010 4.65007
R1770 VDD.n573 VDD.t836 4.65007
R1771 VDD.n258 VDD.t832 4.65007
R1772 VDD.n1323 VDD.t795 4.65007
R1773 VDD.n1327 VDD.t1501 4.65007
R1774 VDD.n1324 VDD.t1495 4.65007
R1775 VDD.n1326 VDD.t1914 4.65007
R1776 VDD.n1282 VDD.t1918 4.65007
R1777 VDD.n1239 VDD.t1563 4.65007
R1778 VDD.n1236 VDD.t255 4.65007
R1779 VDD.n1240 VDD.t1885 4.65007
R1780 VDD.n1237 VDD.t1879 4.65007
R1781 VDD.n1230 VDD.t1569 4.65007
R1782 VDD.n1229 VDD.t1168 4.65007
R1783 VDD.n1220 VDD.t1162 4.65007
R1784 VDD.n1198 VDD.t1160 4.64811
R1785 VDD.n1294 VDD.t1467 4.64811
R1786 VDD.n716 VDD.t1293 4.64811
R1787 VDD.n299 VDD.t1940 4.64811
R1788 VDD.n361 VDD.t1978 4.64811
R1789 VDD.n564 VDD.t2061 4.64811
R1790 VDD.n1092 VDD.t1130 4.64447
R1791 VDD.n940 VDD.t1717 4.64447
R1792 VDD.n1654 VDD.t1719 4.64447
R1793 VDD.n1499 VDD.t1361 4.64447
R1794 VDD.n1514 VDD.t1365 4.64447
R1795 VDD.n879 VDD.t1134 4.64447
R1796 VDD.n78 VDD.t1148 4.64447
R1797 VDD.n1020 VDD.t1110 4.64447
R1798 VDD.n1036 VDD.t1098 4.64447
R1799 VDD.n1052 VDD.t1128 4.64447
R1800 VDD.n119 VDD.t1354 4.64447
R1801 VDD.n1595 VDD.t1367 4.64447
R1802 VDD.n1576 VDD.t1363 4.64447
R1803 VDD.n1555 VDD.t1350 4.64447
R1804 VDD.n1622 VDD.t1753 4.64447
R1805 VDD.n1637 VDD.t1725 4.64447
R1806 VDD.n911 VDD.t1713 4.64447
R1807 VDD.n1076 VDD.t1707 4.64447
R1808 VDD.n630 VDD.t1136 4.64447
R1809 VDD.n700 VDD.t1082 4.64447
R1810 VDD.n671 VDD.t1118 4.64447
R1811 VDD.n1254 VDD.t1812 4.64447
R1812 VDD.n1404 VDD.t1543 4.6442
R1813 VDD.n199 VDD.t2008 4.6442
R1814 VDD.n1385 VDD.t1437 4.6442
R1815 VDD.n216 VDD.t2143 4.6442
R1816 VDD.n480 VDD.t1528 4.6442
R1817 VDD.n490 VDD.t1999 4.6442
R1818 VDD.n503 VDD.t1455 4.6442
R1819 VDD.n513 VDD.t2134 4.6442
R1820 VDD.n1031 VDD.t518 4.64384
R1821 VDD.n838 VDD.t29 4.64384
R1822 VDD.n1022 VDD.t1023 4.64368
R1823 VDD.n913 VDD.t2014 4.64368
R1824 VDD.n625 VDD.t1641 4.64299
R1825 VDD.n1572 VDD.t265 4.63363
R1826 VDD.n1495 VDD.t494 4.63363
R1827 VDD.n1118 VDD.n1117 4.61621
R1828 VDD.n1648 VDD.t12 4.61485
R1829 VDD.n1656 VDD.t8 4.61485
R1830 VDD.n1040 VDD.t522 4.61485
R1831 VDD.n1548 VDD.t730 4.61485
R1832 VDD.n1557 VDD.t727 4.61485
R1833 VDD.n1579 VDD.t387 4.61485
R1834 VDD.n1600 VDD.t716 4.61485
R1835 VDD.n130 VDD.t368 4.61485
R1836 VDD.n123 VDD.t247 4.61485
R1837 VDD.n114 VDD.t484 4.61485
R1838 VDD.n1013 VDD.t271 4.61485
R1839 VDD.n1611 VDD.t577 4.61485
R1840 VDD.n74 VDD.t526 4.61485
R1841 VDD.n1632 VDD.t1217 4.61485
R1842 VDD.n1639 VDD.t120 4.61485
R1843 VDD.n1466 VDD.t490 4.61485
R1844 VDD.n1625 VDD.t488 4.61485
R1845 VDD.n904 VDD.t558 4.61485
R1846 VDD.n882 VDD.t72 4.61485
R1847 VDD.n875 VDD.t1594 4.61485
R1848 VDD.n150 VDD.t687 4.61485
R1849 VDD.n1517 VDD.t241 4.61485
R1850 VDD.n1502 VDD.t916 4.61485
R1851 VDD.n943 VDD.t2174 4.61485
R1852 VDD.n946 VDD.t1555 4.61485
R1853 VDD.n1080 VDD.t92 4.61485
R1854 VDD.n692 VDD.t567 4.61485
R1855 VDD.n673 VDD.t514 4.61485
R1856 VDD.n664 VDD.t763 4.61485
R1857 VDD.n645 VDD.t1585 4.61485
R1858 VDD.n634 VDD.t281 4.61485
R1859 VDD.n1094 VDD.t1583 4.61485
R1860 VDD.n1086 VDD.t34 4.61485
R1861 VDD.n1055 VDD.t1646 4.61485
R1862 VDD.n965 VDD.t279 4.61485
R1863 VDD.n180 VDD.t160 4.61485
R1864 VDD.n181 VDD.t948 4.61485
R1865 VDD.n1411 VDD.t1630 4.61485
R1866 VDD.n465 VDD.t1607 4.61485
R1867 VDD.n468 VDD.t1920 4.61485
R1868 VDD.n469 VDD.t466 4.61485
R1869 VDD.n472 VDD.t551 4.61485
R1870 VDD.n1258 VDD.t590 4.61485
R1871 VDD.n1249 VDD.t703 4.61485
R1872 VDD.n623 VDD.t1089 4.60349
R1873 VDD.n764 VDD.t212 4.58941
R1874 VDD.t215 VDD.n1346 4.58941
R1875 VDD.n1336 VDD.t220 4.58941
R1876 VDD.n395 VDD.t218 4.58941
R1877 VDD.t209 VDD.n544 4.58941
R1878 VDD.n1155 VDD.n1142 4.56745
R1879 VDD.n1154 VDD.n168 4.55648
R1880 VDD.n1135 VDD.n786 4.53191
R1881 VDD.n548 VDD.n547 4.53105
R1882 VDD.n972 VDD.t569 4.53072
R1883 VDD.n1531 VDD.t2027 4.53072
R1884 VDD.n83 VDD.t2123 4.53072
R1885 VDD.n860 VDD.t199 4.53072
R1886 VDD.n1474 VDD.t1198 4.53072
R1887 VDD.n929 VDD.t2165 4.53072
R1888 VDD.n638 VDD.t1200 4.53072
R1889 VDD.n356 VDD.n355 4.523
R1890 VDD.n831 VDD.n829 4.50213
R1891 VDD.n1431 VDD.n1417 4.50213
R1892 VDD.n1119 VDD.n1118 4.50213
R1893 VDD.n804 VDD.n802 4.50213
R1894 VDD.n1439 VDD.n1438 4.50213
R1895 VDD.n1147 VDD.n1145 4.50213
R1896 VDD.n1104 VDD.n837 4.50176
R1897 VDD.n1428 VDD.n1427 4.50176
R1898 VDD.n1128 VDD.n1127 4.50176
R1899 VDD.n811 VDD.n810 4.50176
R1900 VDD.n1450 VDD.n1449 4.50176
R1901 VDD.n1154 VDD.n1153 4.50176
R1902 VDD.n342 VDD.n341 4.50151
R1903 VDD.n1333 VDD.n1332 4.5015
R1904 VDD.n1451 VDD.n1450 4.50144
R1905 VDD.n1429 VDD.n1428 4.50107
R1906 VDD.n1053 VDD.n1052 4.50102
R1907 VDD.n1608 VDD.n78 4.50102
R1908 VDD.n1623 VDD.n1622 4.50102
R1909 VDD.n948 VDD.n940 4.50102
R1910 VDD.n1157 VDD.n1137 4.50088
R1911 VDD.n832 VDD.n821 4.5005
R1912 VDD.n835 VDD.n834 4.5005
R1913 VDD.n833 VDD.n822 4.5005
R1914 VDD.n836 VDD.n827 4.5005
R1915 VDD.n1109 VDD.n822 4.5005
R1916 VDD.n1105 VDD.n828 4.5005
R1917 VDD.n1110 VDD.n821 4.5005
R1918 VDD.n834 VDD.n823 4.5005
R1919 VDD.n830 VDD.n820 4.5005
R1920 VDD.n1106 VDD.n827 4.5005
R1921 VDD.n1422 VDD.n1421 4.5005
R1922 VDD.n1424 VDD.n173 4.5005
R1923 VDD.n1423 VDD.n172 4.5005
R1924 VDD.n1426 VDD.n1425 4.5005
R1925 VDD.n1435 VDD.n172 4.5005
R1926 VDD.n1420 VDD.n1419 4.5005
R1927 VDD.n1421 VDD.n171 4.5005
R1928 VDD.n1434 VDD.n173 4.5005
R1929 VDD.n1430 VDD.n1418 4.5005
R1930 VDD.n1425 VDD.n174 4.5005
R1931 VDD.n1122 VDD.n1121 4.5005
R1932 VDD.n1124 VDD.n790 4.5005
R1933 VDD.n1123 VDD.n789 4.5005
R1934 VDD.n1126 VDD.n1125 4.5005
R1935 VDD.n1133 VDD.n789 4.5005
R1936 VDD.n1129 VDD.n1116 4.5005
R1937 VDD.n1121 VDD.n788 4.5005
R1938 VDD.n1132 VDD.n790 4.5005
R1939 VDD.n1120 VDD.n786 4.5005
R1940 VDD.n1125 VDD.n791 4.5005
R1941 VDD.n805 VDD.n794 4.5005
R1942 VDD.n808 VDD.n807 4.5005
R1943 VDD.n806 VDD.n795 4.5005
R1944 VDD.n809 VDD.n800 4.5005
R1945 VDD.n816 VDD.n795 4.5005
R1946 VDD.n812 VDD.n801 4.5005
R1947 VDD.n817 VDD.n794 4.5005
R1948 VDD.n807 VDD.n796 4.5005
R1949 VDD.n803 VDD.n793 4.5005
R1950 VDD.n813 VDD.n800 4.5005
R1951 VDD.n1444 VDD.n165 4.5005
R1952 VDD.n1447 VDD.n161 4.5005
R1953 VDD.n1446 VDD.n1445 4.5005
R1954 VDD.n1448 VDD.n162 4.5005
R1955 VDD.n1445 VDD.n160 4.5005
R1956 VDD.n164 VDD.n163 4.5005
R1957 VDD.n1444 VDD.n1443 4.5005
R1958 VDD.n1453 VDD.n161 4.5005
R1959 VDD.n167 VDD.n166 4.5005
R1960 VDD.n1452 VDD.n162 4.5005
R1961 VDD.n160 VDD.n158 4.5005
R1962 VDD.n1443 VDD.n1442 4.5005
R1963 VDD.n1440 VDD.n1439 4.5005
R1964 VDD.n1441 VDD.n167 4.5005
R1965 VDD.n163 VDD.n159 4.5005
R1966 VDD.n1454 VDD.n1453 4.5005
R1967 VDD.n1452 VDD.n1451 4.5005
R1968 VDD.n816 VDD.n815 4.5005
R1969 VDD.n812 VDD.n798 4.5005
R1970 VDD.n818 VDD.n817 4.5005
R1971 VDD.n802 VDD.n792 4.5005
R1972 VDD.n797 VDD.n796 4.5005
R1973 VDD.n811 VDD.n156 4.5005
R1974 VDD.n799 VDD.n793 4.5005
R1975 VDD.n814 VDD.n813 4.5005
R1976 VDD.n1596 VDD.n1595 4.5005
R1977 VDD.n1515 VDD.n1514 4.5005
R1978 VDD.n701 VDD.n700 4.5005
R1979 VDD.n1163 VDD.n780 4.5005
R1980 VDD.n1148 VDD.n1138 4.5005
R1981 VDD.n1151 VDD.n1150 4.5005
R1982 VDD.n1149 VDD.n1139 4.5005
R1983 VDD.n1152 VDD.n1143 4.5005
R1984 VDD.n1159 VDD.n1139 4.5005
R1985 VDD.n1155 VDD.n1144 4.5005
R1986 VDD.n1160 VDD.n1138 4.5005
R1987 VDD.n1150 VDD.n1140 4.5005
R1988 VDD.n1146 VDD.n1137 4.5005
R1989 VDD.n1156 VDD.n1143 4.5005
R1990 VDD.n1159 VDD.n1158 4.5005
R1991 VDD.n1161 VDD.n1160 4.5005
R1992 VDD.n1145 VDD.n1136 4.5005
R1993 VDD.n1141 VDD.n1140 4.5005
R1994 VDD.n1157 VDD.n1156 4.5005
R1995 VDD.n1134 VDD.n1133 4.5005
R1996 VDD.n1128 VDD.n1115 4.5005
R1997 VDD.n1114 VDD.n791 4.5005
R1998 VDD.n1130 VDD.n1129 4.5005
R1999 VDD.n1117 VDD.n788 4.5005
R2000 VDD.n1132 VDD.n1131 4.5005
R2001 VDD.n1436 VDD.n1435 4.5005
R2002 VDD.n1419 VDD.n169 4.5005
R2003 VDD.n1416 VDD.n171 4.5005
R2004 VDD.n1432 VDD.n1431 4.5005
R2005 VDD.n1434 VDD.n1433 4.5005
R2006 VDD.n1430 VDD.n1429 4.5005
R2007 VDD.n174 VDD.n170 4.5005
R2008 VDD.n1109 VDD.n1108 4.5005
R2009 VDD.n1105 VDD.n825 4.5005
R2010 VDD.n1111 VDD.n1110 4.5005
R2011 VDD.n829 VDD.n819 4.5005
R2012 VDD.n824 VDD.n823 4.5005
R2013 VDD.n1104 VDD.n1103 4.5005
R2014 VDD.n826 VDD.n820 4.5005
R2015 VDD.n1107 VDD.n1106 4.5005
R2016 VDD.n350 VDD.n284 4.5005
R2017 VDD.n353 VDD.n352 4.5005
R2018 VDD.n354 VDD.n281 4.5005
R2019 VDD.n1246 VDD.n1245 4.5005
R2020 VDD.n6 VDD.t1417 4.2255
R2021 VDD.n10 VDD.t1289 4.2255
R2022 VDD.n0 VDD.t1924 4.2255
R2023 VDD.n784 VDD.t2171 4.2255
R2024 VDD.n41 VDD.t1705 4.2255
R2025 VDD.n43 VDD.t807 4.2255
R2026 VDD.n42 VDD.t370 4.2255
R2027 VDD.n1658 VDD.t1711 4.2255
R2028 VDD.n1489 VDD.t1381 4.2255
R2029 VDD.n990 VDD.t1051 4.2255
R2030 VDD.n970 VDD.t933 4.2255
R2031 VDD.n973 VDD.t543 4.2255
R2032 VDD.n979 VDD.t535 4.2255
R2033 VDD.n981 VDD.t694 4.2255
R2034 VDD.n1519 VDD.t1348 4.2255
R2035 VDD.n1520 VDD.t593 4.2255
R2036 VDD.n1521 VDD.t633 4.2255
R2037 VDD.n1567 VDD.t1326 4.2255
R2038 VDD.n1563 VDD.t1346 4.2255
R2039 VDD.n1537 VDD.t928 4.2255
R2040 VDD.n1529 VDD.t751 4.2255
R2041 VDD.n1532 VDD.t439 4.2255
R2042 VDD.n133 VDD.t1868 4.2255
R2043 VDD.n88 VDD.t312 4.2255
R2044 VDD.n89 VDD.t722 4.2255
R2045 VDD.n97 VDD.t1352 4.2255
R2046 VDD.n99 VDD.t205 4.2255
R2047 VDD.n101 VDD.t226 4.2255
R2048 VDD.n109 VDD.t1358 4.2255
R2049 VDD.n995 VDD.t1055 4.2255
R2050 VDD.n1001 VDD.t649 4.2255
R2051 VDD.n1004 VDD.t1614 4.2255
R2052 VDD.n84 VDD.t1623 4.2255
R2053 VDD.n81 VDD.t993 4.2255
R2054 VDD.n1613 VDD.t169 4.2255
R2055 VDD.n69 VDD.t581 4.2255
R2056 VDD.n1468 VDD.t1598 4.2255
R2057 VDD.n1460 VDD.t288 4.2255
R2058 VDD.n47 VDD.t1762 4.2255
R2059 VDD.n58 VDD.t46 4.2255
R2060 VDD.n53 VDD.t1223 4.2255
R2061 VDD.n57 VDD.t1770 4.2255
R2062 VDD.n849 VDD.t1728 4.2255
R2063 VDD.n855 VDD.t82 4.2255
R2064 VDD.n858 VDD.t445 4.2255
R2065 VDD.n861 VDD.t447 4.2255
R2066 VDD.n66 VDD.t54 4.2255
R2067 VDD.n886 VDD.t1063 4.2255
R2068 VDD.n887 VDD.t79 4.2255
R2069 VDD.n866 VDD.t291 4.2255
R2070 VDD.n846 VDD.t1062 4.2255
R2071 VDD.n143 VDD.t781 4.2255
R2072 VDD.n140 VDD.t187 4.2255
R2073 VDD.n1475 VDD.t1601 4.2255
R2074 VDD.n155 VDD.t63 4.2255
R2075 VDD.n1480 VDD.t918 4.2255
R2076 VDD.n1472 VDD.t19 4.2255
R2077 VDD.n17 VDD.t1283 4.2255
R2078 VDD.n27 VDD.t1291 4.2255
R2079 VDD.n22 VDD.t1002 4.2255
R2080 VDD.n33 VDD.t411 4.2255
R2081 VDD.n32 VDD.t772 4.2255
R2082 VDD.n843 VDD.t1766 4.2255
R2083 VDD.n927 VDD.t233 4.2255
R2084 VDD.n1067 VDD.t98 4.2255
R2085 VDD.n935 VDD.t1697 4.2255
R2086 VDD.n930 VDD.t153 4.2255
R2087 VDD.n775 VDD.t1228 4.2255
R2088 VDD.n776 VDD.t1235 4.2255
R2089 VDD.n777 VDD.t1253 4.2255
R2090 VDD.n778 VDD.t1231 4.2255
R2091 VDD.n779 VDD.t1234 4.2255
R2092 VDD.n604 VDD.t1463 4.2255
R2093 VDD.n603 VDD.t87 4.2255
R2094 VDD.t212 VDD.n749 4.2255
R2095 VDD.n648 VDD.t431 4.2255
R2096 VDD.n651 VDD.t476 4.2255
R2097 VDD.n658 VDD.t1142 4.2255
R2098 VDD.n654 VDD.t114 4.2255
R2099 VDD.n653 VDD.t473 4.2255
R2100 VDD.n652 VDD.t1037 4.2255
R2101 VDD.n644 VDD.t944 4.2255
R2102 VDD.n639 VDD.t532 4.2255
R2103 VDD.n636 VDD.t133 4.2255
R2104 VDD.n611 VDD.t672 4.2255
R2105 VDD.n609 VDD.t1071 4.2255
R2106 VDD.n1096 VDD.t1122 4.2255
R2107 VDD.n923 VDD.t42 4.2255
R2108 VDD.n1058 VDD.t622 4.2255
R2109 VDD.n1057 VDD.t1121 4.2255
R2110 VDD.n958 VDD.t360 4.2255
R2111 VDD.n1347 VDD.t215 4.2255
R2112 VDD.n1334 VDD.t220 4.2255
R2113 VDD.n288 VDD.t690 4.2255
R2114 VDD.n346 VDD.t1465 4.2255
R2115 VDD.t218 VDD.n394 4.2255
R2116 VDD.n545 VDD.t209 4.2255
R2117 VDD.n597 VDD.t612 4.2255
R2118 VDD.n596 VDD.t382 4.2255
R2119 VDD.n1265 VDD.t1779 4.2255
R2120 VDD.t1042 VDD.n885 3.83743
R2121 VDD.n1099 VDD.t1034 3.83743
R2122 VDD.n972 VDD.n971 3.75093
R2123 VDD.n975 VDD.n974 3.75093
R2124 VDD.n1531 VDD.n1530 3.75093
R2125 VDD.n1534 VDD.n1533 3.75093
R2126 VDD.n83 VDD.n82 3.75093
R2127 VDD.n86 VDD.n85 3.75093
R2128 VDD.n860 VDD.n859 3.75093
R2129 VDD.n863 VDD.n862 3.75093
R2130 VDD.n1474 VDD.n1473 3.75093
R2131 VDD.n1477 VDD.n1476 3.75093
R2132 VDD.n929 VDD.n928 3.75093
R2133 VDD.n932 VDD.n931 3.75093
R2134 VDD.n638 VDD.n637 3.75093
R2135 VDD.n641 VDD.n640 3.75093
R2136 VDD.t981 VDD.t86 3.73804
R2137 VDD.n767 VDD.n747 3.70515
R2138 VDD.n770 VDD.n768 3.54746
R2139 VDD.n783 VDD.n781 3.54746
R2140 VDD.n187 VDD.n185 3.54746
R2141 VDD.n197 VDD.n195 3.54746
R2142 VDD.n205 VDD.n203 3.54746
R2143 VDD.n214 VDD.n212 3.54746
R2144 VDD.n223 VDD.n221 3.54746
R2145 VDD.n233 VDD.n231 3.54746
R2146 VDD.n245 VDD.n243 3.54746
R2147 VDD.n453 VDD.n451 3.54746
R2148 VDD.n447 VDD.n445 3.54746
R2149 VDD.n440 VDD.n438 3.54746
R2150 VDD.n434 VDD.n432 3.54746
R2151 VDD.n426 VDD.n424 3.54746
R2152 VDD.n414 VDD.n412 3.54746
R2153 VDD.n399 VDD.n397 3.54746
R2154 VDD.n16 VDD.n14 3.5318
R2155 VDD.n9 VDD.n7 3.5318
R2156 VDD.n4 VDD.n2 3.5318
R2157 VDD.n1226 VDD.n1224 3.5318
R2158 VDD.n26 VDD.n24 3.5318
R2159 VDD.n20 VDD.n18 3.5318
R2160 VDD.n1525 VDD.t403 3.43297
R2161 VDD.n39 VDD.n37 3.30485
R2162 VDD.n1645 VDD.n1643 3.30485
R2163 VDD.n1487 VDD.n1485 3.30485
R2164 VDD.n988 VDD.n986 3.30485
R2165 VDD.n137 VDD.n135 3.30485
R2166 VDD.n1545 VDD.n1543 3.30485
R2167 VDD.n1561 VDD.n1559 3.30485
R2168 VDD.n96 VDD.n94 3.30485
R2169 VDD.n108 VDD.n106 3.30485
R2170 VDD.n998 VDD.n996 3.30485
R2171 VDD.n50 VDD.n48 3.30485
R2172 VDD.n63 VDD.n61 3.30485
R2173 VDD.n852 VDD.n850 3.30485
R2174 VDD.n892 VDD.n890 3.30485
R2175 VDD.n873 VDD.n871 3.30485
R2176 VDD.n841 VDD.n839 3.30485
R2177 VDD.n618 VDD.n616 3.30485
R2178 VDD.n661 VDD.n659 3.30485
R2179 VDD.n684 VDD.n682 3.30485
R2180 VDD.n920 VDD.n918 3.30485
R2181 VDD.n955 VDD.n953 3.30485
R2182 VDD.n594 VDD.n592 3.30485
R2183 VDD.n1335 VDD.n1333 3.2789
R2184 VDD.n547 VDD.n546 3.25303
R2185 VDD.n1440 VDD.n1437 3.17341
R2186 VDD.n1564 VDD.n1542 3.1505
R2187 VDD.n1569 VDD.n1542 3.1505
R2188 VDD.n993 VDD.n992 3.1505
R2189 VDD.n1028 VDD.n993 3.1505
R2190 VDD.n1025 VDD.n1024 3.1505
R2191 VDD.n1026 VDD.n1025 3.1505
R2192 VDD.n916 VDD.n915 3.1505
R2193 VDD.n917 VDD.n916 3.1505
R2194 VDD.n1491 VDD.n1490 3.1505
R2195 VDD.n1492 VDD.n1491 3.1505
R2196 VDD.n621 VDD.n620 3.1505
R2197 VDD.n622 VDD.n621 3.1505
R2198 VDD.n845 VDD.n844 3.1505
R2199 VDD.n1098 VDD.n845 3.1505
R2200 VDD.n31 VDD.n30 3.07058
R2201 VDD.n343 VDD.n342 3.04391
R2202 VDD.n1197 VDD.n1196 3.02507
R2203 VDD.n1214 VDD.n1200 3.02507
R2204 VDD.n1209 VDD.n1202 3.02507
R2205 VDD.n1204 VDD.n1203 3.02507
R2206 VDD.n1293 VDD.n591 3.02507
R2207 VDD.n1297 VDD.n1296 3.02507
R2208 VDD.n1305 VDD.n1302 3.02507
R2209 VDD.n1310 VDD.n589 3.02507
R2210 VDD.n1270 VDD.n1269 3.02507
R2211 VDD.n1276 VDD.n1271 3.02507
R2212 VDD.n588 VDD.n587 3.02507
R2213 VDD.n732 VDD.n712 3.02507
R2214 VDD.n727 VDD.n713 3.02507
R2215 VDD.n711 VDD.n710 3.02507
R2216 VDD.n739 VDD.n709 3.02507
R2217 VDD.n708 VDD.n707 3.02507
R2218 VDD.n758 VDD.n757 3.02507
R2219 VDD.n705 VDD.n704 3.02507
R2220 VDD.n1181 VDD.n608 3.02507
R2221 VDD.n720 VDD.n718 3.02507
R2222 VDD.n715 VDD.n714 3.02507
R2223 VDD.n1409 VDD.n184 3.02507
R2224 VDD.n1403 VDD.n190 3.02507
R2225 VDD.n194 VDD.n191 3.02507
R2226 VDD.n200 VDD.n198 3.02507
R2227 VDD.n1390 VDD.n201 3.02507
R2228 VDD.n1384 VDD.n207 3.02507
R2229 VDD.n211 VDD.n208 3.02507
R2230 VDD.n217 VDD.n215 3.02507
R2231 VDD.n219 VDD.n218 3.02507
R2232 VDD.n236 VDD.n235 3.02507
R2233 VDD.n239 VDD.n234 3.02507
R2234 VDD.n229 VDD.n224 3.02507
R2235 VDD.n226 VDD.n225 3.02507
R2236 VDD.n247 VDD.n246 3.02507
R2237 VDD.n291 VDD.n290 3.02507
R2238 VDD.n294 VDD.n293 3.02507
R2239 VDD.n334 VDD.n292 3.02507
R2240 VDD.n327 VDD.n295 3.02507
R2241 VDD.n322 VDD.n296 3.02507
R2242 VDD.n298 VDD.n297 3.02507
R2243 VDD.n315 VDD.n301 3.02507
R2244 VDD.n310 VDD.n303 3.02507
R2245 VDD.n305 VDD.n304 3.02507
R2246 VDD.n560 VDD.n270 3.02507
R2247 VDD.n272 VDD.n271 3.02507
R2248 VDD.n277 VDD.n274 3.02507
R2249 VDD.n553 VDD.n273 3.02507
R2250 VDD.n461 VDD.n460 3.02507
R2251 VDD.n474 VDD.n455 3.02507
R2252 VDD.n481 VDD.n450 3.02507
R2253 VDD.n449 VDD.n448 3.02507
R2254 VDD.n444 VDD.n443 3.02507
R2255 VDD.n497 VDD.n442 3.02507
R2256 VDD.n504 VDD.n437 3.02507
R2257 VDD.n436 VDD.n435 3.02507
R2258 VDD.n431 VDD.n430 3.02507
R2259 VDD.n428 VDD.n427 3.02507
R2260 VDD.n417 VDD.n416 3.02507
R2261 VDD.n420 VDD.n415 3.02507
R2262 VDD.n410 VDD.n405 3.02507
R2263 VDD.n407 VDD.n406 3.02507
R2264 VDD.n401 VDD.n400 3.02507
R2265 VDD.n377 VDD.n278 3.02507
R2266 VDD.n372 VDD.n369 3.02507
R2267 VDD.n364 VDD.n363 3.02507
R2268 VDD.n360 VDD.n280 3.02507
R2269 VDD.n283 VDD.n282 3.02507
R2270 VDD.n1318 VDD.n264 3.02507
R2271 VDD.n266 VDD.n265 3.02507
R2272 VDD.n268 VDD.n267 3.02507
R2273 VDD.n580 VDD.n566 3.02507
R2274 VDD.n575 VDD.n568 3.02507
R2275 VDD.n570 VDD.n569 3.02507
R2276 VDD.n263 VDD.n262 3.02507
R2277 VDD.n1325 VDD.n261 3.02507
R2278 VDD.n260 VDD.n259 3.02507
R2279 VDD.n1283 VDD.n1281 3.02507
R2280 VDD.n1268 VDD.n1267 3.02507
R2281 VDD.n1190 VDD.n1189 3.02507
R2282 VDD.n1193 VDD.n1192 3.02507
R2283 VDD.n1238 VDD.n1191 3.02507
R2284 VDD.n1231 VDD.n1194 3.02507
R2285 VDD.n1221 VDD.n1195 3.02507
R2286 VDD.n1413 VDD.n182 2.97615
R2287 VDD.n1412 VDD.n183 2.97615
R2288 VDD.n939 VDD.n936 2.97615
R2289 VDD.n938 VDD.n937 2.97615
R2290 VDD.n1650 VDD.n1646 2.97615
R2291 VDD.n1649 VDD.n1647 2.97615
R2292 VDD.n1512 VDD.n1511 2.97615
R2293 VDD.n1513 VDD.n1510 2.97615
R2294 VDD.n1019 VDD.n1016 2.97615
R2295 VDD.n1018 VDD.n1017 2.97615
R2296 VDD.n1034 VDD.n1033 2.97615
R2297 VDD.n1035 VDD.n1032 2.97615
R2298 VDD.n1039 VDD.n984 2.97615
R2299 VDD.n1038 VDD.n985 2.97615
R2300 VDD.n1051 VDD.n1048 2.97615
R2301 VDD.n1050 VDD.n1049 2.97615
R2302 VDD.n117 VDD.n116 2.97615
R2303 VDD.n118 VDD.n115 2.97615
R2304 VDD.n1593 VDD.n1592 2.97615
R2305 VDD.n1594 VDD.n1591 2.97615
R2306 VDD.n1553 VDD.n1552 2.97615
R2307 VDD.n1554 VDD.n1551 2.97615
R2308 VDD.n1549 VDD.n1547 2.97615
R2309 VDD.n1550 VDD.n1546 2.97615
R2310 VDD.n1599 VDD.n92 2.97615
R2311 VDD.n1598 VDD.n93 2.97615
R2312 VDD.n122 VDD.n104 2.97615
R2313 VDD.n121 VDD.n105 2.97615
R2314 VDD.n1015 VDD.n999 2.97615
R2315 VDD.n1014 VDD.n1000 2.97615
R2316 VDD.n910 VDD.n907 2.97615
R2317 VDD.n909 VDD.n908 2.97615
R2318 VDD.n906 VDD.n853 2.97615
R2319 VDD.n905 VDD.n854 2.97615
R2320 VDD.n151 VDD.n139 2.97615
R2321 VDD.n152 VDD.n138 2.97615
R2322 VDD.n945 VDD.n941 2.97615
R2323 VDD.n944 VDD.n942 2.97615
R2324 VDD.n1074 VDD.n1073 2.97615
R2325 VDD.n1075 VDD.n1072 2.97615
R2326 VDD.n1079 VDD.n1070 2.97615
R2327 VDD.n1078 VDD.n1071 2.97615
R2328 VDD.n628 VDD.n627 2.97615
R2329 VDD.n629 VDD.n626 2.97615
R2330 VDD.n699 VDD.n696 2.97615
R2331 VDD.n698 VDD.n697 2.97615
R2332 VDD.n670 VDD.n667 2.97615
R2333 VDD.n669 VDD.n668 2.97615
R2334 VDD.n694 VDD.n646 2.97615
R2335 VDD.n693 VDD.n647 2.97615
R2336 VDD.n666 VDD.n662 2.97615
R2337 VDD.n665 VDD.n663 2.97615
R2338 VDD.n633 VDD.n614 2.97615
R2339 VDD.n632 VDD.n615 2.97615
R2340 VDD.n1088 VDD.n921 2.97615
R2341 VDD.n1087 VDD.n922 2.97615
R2342 VDD.n967 VDD.n956 2.97615
R2343 VDD.n966 VDD.n957 2.97615
R2344 VDD.n178 VDD.n177 2.97615
R2345 VDD.n179 VDD.n176 2.97615
R2346 VDD.n466 VDD.n459 2.97615
R2347 VDD.n467 VDD.n458 2.97615
R2348 VDD.n470 VDD.n457 2.97615
R2349 VDD.n471 VDD.n456 2.97615
R2350 VDD.n1253 VDD.n1250 2.97615
R2351 VDD.n1252 VDD.n1251 2.97615
R2352 VDD.n1256 VDD.n601 2.97615
R2353 VDD.n1257 VDD.n600 2.97615
R2354 VDD.n1162 VDD.n1161 2.94069
R2355 VDD.n240 VDD.n239 2.93344
R2356 VDD.n421 VDD.n420 2.93344
R2357 VDD.n242 VDD.n230 2.73226
R2358 VDD.n423 VDD.n411 2.73226
R2359 VDD VDD.n88 2.61227
R2360 VDD VDD.n1613 2.61227
R2361 VDD VDD.n1468 2.61227
R2362 VDD VDD.n143 2.61227
R2363 VDD VDD.n651 2.61227
R2364 VDD VDD.n596 2.61227
R2365 VDD.n1605 VDD.t2122 2.6092
R2366 VDD.n1507 VDD.t1199 2.6092
R2367 VDD.n16 VDD.n15 2.6005
R2368 VDD.n9 VDD.n8 2.6005
R2369 VDD.n4 VDD.n3 2.6005
R2370 VDD.n1226 VDD.n1225 2.6005
R2371 VDD.n39 VDD.n38 2.6005
R2372 VDD.n45 VDD.n44 2.6005
R2373 VDD.n1645 VDD.n1644 2.6005
R2374 VDD.n1487 VDD.n1486 2.6005
R2375 VDD.n988 VDD.n987 2.6005
R2376 VDD.n969 VDD.n968 2.6005
R2377 VDD.n983 VDD.n982 2.6005
R2378 VDD.n137 VDD.n136 2.6005
R2379 VDD.n1523 VDD.n1522 2.6005
R2380 VDD.n1545 VDD.n1544 2.6005
R2381 VDD.n1561 VDD.n1560 2.6005
R2382 VDD.n1539 VDD.n1538 2.6005
R2383 VDD.n132 VDD.n131 2.6005
R2384 VDD.n91 VDD.n90 2.6005
R2385 VDD.n96 VDD.n95 2.6005
R2386 VDD.n103 VDD.n102 2.6005
R2387 VDD.n108 VDD.n107 2.6005
R2388 VDD.n998 VDD.n997 2.6005
R2389 VDD.n1003 VDD.n1002 2.6005
R2390 VDD.n80 VDD.n79 2.6005
R2391 VDD.n71 VDD.n70 2.6005
R2392 VDD.n1462 VDD.n1461 2.6005
R2393 VDD.n50 VDD.n49 2.6005
R2394 VDD.n55 VDD.n54 2.6005
R2395 VDD.n63 VDD.n62 2.6005
R2396 VDD.n852 VDD.n851 2.6005
R2397 VDD.n857 VDD.n856 2.6005
R2398 VDD.n65 VDD.n64 2.6005
R2399 VDD.n892 VDD.n891 2.6005
R2400 VDD.n868 VDD.n867 2.6005
R2401 VDD.n873 VDD.n872 2.6005
R2402 VDD.n142 VDD.n141 2.6005
R2403 VDD.n154 VDD.n153 2.6005
R2404 VDD.n1482 VDD.n1481 2.6005
R2405 VDD.n26 VDD.n25 2.6005
R2406 VDD.n20 VDD.n19 2.6005
R2407 VDD.n35 VDD.n34 2.6005
R2408 VDD.n841 VDD.n840 2.6005
R2409 VDD.n1069 VDD.n1068 2.6005
R2410 VDD.n934 VDD.n933 2.6005
R2411 VDD.n606 VDD.n605 2.6005
R2412 VDD.n752 VDD.n751 2.6005
R2413 VDD.n756 VDD.n755 2.6005
R2414 VDD.n770 VDD.n769 2.6005
R2415 VDD.n618 VDD.n617 2.6005
R2416 VDD.n650 VDD.n649 2.6005
R2417 VDD.n661 VDD.n660 2.6005
R2418 VDD.n656 VDD.n655 2.6005
R2419 VDD.n684 VDD.n683 2.6005
R2420 VDD.n643 VDD.n642 2.6005
R2421 VDD.n613 VDD.n612 2.6005
R2422 VDD.n920 VDD.n919 2.6005
R2423 VDD.n925 VDD.n924 2.6005
R2424 VDD.n955 VDD.n954 2.6005
R2425 VDD.n960 VDD.n959 2.6005
R2426 VDD.n783 VDD.n782 2.6005
R2427 VDD.n187 VDD.n186 2.6005
R2428 VDD.n197 VDD.n196 2.6005
R2429 VDD.n205 VDD.n204 2.6005
R2430 VDD.n214 VDD.n213 2.6005
R2431 VDD.n223 VDD.n222 2.6005
R2432 VDD.n233 VDD.n232 2.6005
R2433 VDD.n245 VDD.n244 2.6005
R2434 VDD.n1340 VDD.n1339 2.6005
R2435 VDD.n1344 VDD.n1343 2.6005
R2436 VDD.n253 VDD.n252 2.6005
R2437 VDD.n257 VDD.n256 2.6005
R2438 VDD.n348 VDD.n347 2.6005
R2439 VDD.n453 VDD.n452 2.6005
R2440 VDD.n447 VDD.n446 2.6005
R2441 VDD.n440 VDD.n439 2.6005
R2442 VDD.n434 VDD.n433 2.6005
R2443 VDD.n426 VDD.n425 2.6005
R2444 VDD.n414 VDD.n413 2.6005
R2445 VDD.n399 VDD.n398 2.6005
R2446 VDD.n389 VDD.n388 2.6005
R2447 VDD.n393 VDD.n392 2.6005
R2448 VDD.n381 VDD.n380 2.6005
R2449 VDD.n385 VDD.n384 2.6005
R2450 VDD.n599 VDD.n598 2.6005
R2451 VDD.n594 VDD.n593 2.6005
R2452 VDD.n1168 VDD.n774 2.50668
R2453 VDD.n220 VDD.n219 2.4665
R2454 VDD.n429 VDD.n428 2.4665
R2455 VDD.n228 VDD.n227 2.44638
R2456 VDD.n409 VDD.n408 2.44638
R2457 VDD.n1437 VDD.n168 2.36511
R2458 VDD.n785 VDD.n784 2.32427
R2459 VDD.n832 VDD.n831 2.30085
R2460 VDD.n1422 VDD.n1417 2.30085
R2461 VDD.n1122 VDD.n1119 2.30085
R2462 VDD.n805 VDD.n804 2.30085
R2463 VDD.n1438 VDD.n165 2.30085
R2464 VDD.n1148 VDD.n1147 2.30085
R2465 VDD.n837 VDD.n836 2.29544
R2466 VDD.n1427 VDD.n1426 2.29544
R2467 VDD.n1127 VDD.n1126 2.29544
R2468 VDD.n810 VDD.n809 2.29544
R2469 VDD.n1449 VDD.n1448 2.29544
R2470 VDD.n1153 VDD.n1152 2.29544
R2471 VDD.n227 VDD.n226 2.28756
R2472 VDD.n229 VDD.n228 2.28756
R2473 VDD.n230 VDD.n229 2.28756
R2474 VDD.n239 VDD.n238 2.28756
R2475 VDD.n237 VDD.n236 2.28756
R2476 VDD.n408 VDD.n407 2.28756
R2477 VDD.n410 VDD.n409 2.28756
R2478 VDD.n411 VDD.n410 2.28756
R2479 VDD.n420 VDD.n419 2.28756
R2480 VDD.n418 VDD.n417 2.28756
R2481 VDD.t502 VDD.t1089 2.26039
R2482 VDD.n1188 VDD.n603 2.21779
R2483 VDD VDD.n762 2.20189
R2484 VDD.n1171 VDD.t1201 2.17284
R2485 VDD.n1317 VDD 2.13233
R2486 VDD.n1282 VDD 2.13233
R2487 VDD.n1352 VDD.n1351 2.1005
R2488 VDD.n1350 VDD.n1349 2.1005
R2489 VDD.n540 VDD.n539 2.1005
R2490 VDD.n542 VDD.n541 2.1005
R2491 VDD.n1185 VDD.t30 2.04555
R2492 VDD.n343 VDD.n288 2.04357
R2493 VDD.n242 VDD.n241 2.03874
R2494 VDD.n423 VDD.n422 2.03874
R2495 VDD.n1168 VDD 2.03836
R2496 VDD.n241 VDD.n240 1.99109
R2497 VDD.n422 VDD.n421 1.99109
R2498 VDD.n1112 VDD.n818 1.96654
R2499 VDD.n238 VDD.n237 1.94874
R2500 VDD.n419 VDD.n418 1.94874
R2501 VDD.n1664 VDD.n42 1.88267
R2502 VDD.n980 VDD.n979 1.88267
R2503 VDD.n1584 VDD.n1520 1.88267
R2504 VDD.n1536 VDD.n1529 1.88267
R2505 VDD.n100 VDD.n99 1.88267
R2506 VDD.n1005 VDD.n1004 1.88267
R2507 VDD.n59 VDD.n58 1.88267
R2508 VDD.n865 VDD.n858 1.88267
R2509 VDD.n888 VDD.n887 1.88267
R2510 VDD.n1479 VDD.n1472 1.88267
R2511 VDD.n1671 VDD.n32 1.88267
R2512 VDD.n1066 VDD.n927 1.88267
R2513 VDD.n680 VDD.n653 1.88267
R2514 VDD.n1174 VDD.n636 1.88267
R2515 VDD.n1059 VDD.n1058 1.88267
R2516 VDD.n901 VDD.n900 1.82579
R2517 VDD.n1083 VDD.n926 1.82579
R2518 VDD.n1457 VDD.n1456 1.80258
R2519 VDD.n1589 VDD.n1588 1.8005
R2520 VDD.n1046 VDD.n1045 1.8005
R2521 VDD.n1606 VDD.n1605 1.8005
R2522 VDD.n1617 VDD.n1616 1.8005
R2523 VDD.n1508 VDD.n1507 1.8005
R2524 VDD.n1172 VDD.n1171 1.8005
R2525 VDD.n1064 VDD.n1063 1.8005
R2526 VDD.n1113 VDD.n1112 1.79408
R2527 VDD.n731 VDD.n730 1.68244
R2528 VDD.n326 VDD.n325 1.68244
R2529 VDD.n1230 VDD.n1229 1.68244
R2530 VDD.n1009 VDD.n1007 1.65613
R2531 VDD.n1213 VDD 1.63504
R2532 VDD VDD.n590 1.63504
R2533 VDD.n719 VDD 1.63504
R2534 VDD.n314 VDD 1.63504
R2535 VDD VDD.n279 1.63504
R2536 VDD.n579 VDD 1.63504
R2537 VDD.n15 VDD.t1270 1.6255
R2538 VDD.n15 VDD.t1272 1.6255
R2539 VDD.n14 VDD.t1285 1.6255
R2540 VDD.n14 VDD.t1287 1.6255
R2541 VDD.n8 VDD.t1410 1.6255
R2542 VDD.n8 VDD.t1412 1.6255
R2543 VDD.n7 VDD.t1415 1.6255
R2544 VDD.n7 VDD.t1416 1.6255
R2545 VDD.n3 VDD.t1286 1.6255
R2546 VDD.n3 VDD.t1288 1.6255
R2547 VDD.n2 VDD.t1274 1.6255
R2548 VDD.n2 VDD.t1276 1.6255
R2549 VDD.n1225 VDD.t1930 1.6255
R2550 VDD.n1225 VDD.t1931 1.6255
R2551 VDD.n1224 VDD.t1926 1.6255
R2552 VDD.n1224 VDD.t1928 1.6255
R2553 VDD.n1196 VDD.t1156 1.6255
R2554 VDD.n1196 VDD.t1154 1.6255
R2555 VDD.n1200 VDD.t1881 1.6255
R2556 VDD.n1200 VDD.t1877 1.6255
R2557 VDD.n1202 VDD.t259 1.6255
R2558 VDD.n1202 VDD.t263 1.6255
R2559 VDD.n1203 VDD.t1567 1.6255
R2560 VDD.n1203 VDD.t1559 1.6255
R2561 VDD.n591 VDD.t1460 1.6255
R2562 VDD.n591 VDD.t1462 1.6255
R2563 VDD.n1296 VDD.t960 1.6255
R2564 VDD.n1296 VDD.t958 1.6255
R2565 VDD.n1302 VDD.t793 1.6255
R2566 VDD.n1302 VDD.t791 1.6255
R2567 VDD.n589 VDD.t874 1.6255
R2568 VDD.n589 VDD.t820 1.6255
R2569 VDD.n1269 VDD.t2155 1.6255
R2570 VDD.n1269 VDD.t2157 1.6255
R2571 VDD.n1271 VDD.t966 1.6255
R2572 VDD.n1271 VDD.t1893 1.6255
R2573 VDD.n587 VDD.t850 1.6255
R2574 VDD.n587 VDD.t816 1.6255
R2575 VDD.n182 VDD.t946 1.6255
R2576 VDD.n182 VDD.t757 1.6255
R2577 VDD.n183 VDD.t759 1.6255
R2578 VDD.n183 VDD.t1632 1.6255
R2579 VDD.n1090 VDD.t860 1.6255
R2580 VDD.n1090 VDD.t1132 1.6255
R2581 VDD.n1089 VDD.t364 1.6255
R2582 VDD.n1089 VDD.t828 1.6255
R2583 VDD.n936 VDD.t1798 1.6255
R2584 VDD.n936 VDD.t1733 1.6255
R2585 VDD.n937 VDD.t346 1.6255
R2586 VDD.n937 VDD.t1788 1.6255
R2587 VDD.n1652 VDD.t1908 1.6255
R2588 VDD.n1652 VDD.t1721 1.6255
R2589 VDD.n1651 VDD.t609 1.6255
R2590 VDD.n1651 VDD.t908 1.6255
R2591 VDD.n38 VDD.t1715 1.6255
R2592 VDD.n38 VDD.t1740 1.6255
R2593 VDD.n37 VDD.t1750 1.6255
R2594 VDD.n37 VDD.t1771 1.6255
R2595 VDD.n44 VDD.t809 1.6255
R2596 VDD.n44 VDD.t810 1.6255
R2597 VDD.n1646 VDD.t856 1.6255
R2598 VDD.n1646 VDD.t10 1.6255
R2599 VDD.n1647 VDD.t14 1.6255
R2600 VDD.n1647 VDD.t844 1.6255
R2601 VDD.n1644 VDD.t1727 1.6255
R2602 VDD.n1644 VDD.t1772 1.6255
R2603 VDD.n1643 VDD.t1751 1.6255
R2604 VDD.n1643 VDD.t1757 1.6255
R2605 VDD.n1486 VDD.t1324 1.6255
R2606 VDD.n1486 VDD.t1356 1.6255
R2607 VDD.n1485 VDD.t1383 1.6255
R2608 VDD.n1485 VDD.t1332 1.6255
R2609 VDD.n1497 VDD.t1950 1.6255
R2610 VDD.n1497 VDD.t1335 1.6255
R2611 VDD.n1496 VDD.t137 1.6255
R2612 VDD.n1496 VDD.t1970 1.6255
R2613 VDD.n1511 VDD.t724 1.6255
R2614 VDD.n1511 VDD.t1972 1.6255
R2615 VDD.n1510 VDD.t1952 1.6255
R2616 VDD.n1510 VDD.t1337 1.6255
R2617 VDD.n877 VDD.t891 1.6255
R2618 VDD.n877 VDD.t193 1.6255
R2619 VDD.n876 VDD.t1049 1.6255
R2620 VDD.n876 VDD.t1916 1.6255
R2621 VDD.n76 VDD.t1816 1.6255
R2622 VDD.n76 VDD.t641 1.6255
R2623 VDD.n75 VDD.t1039 1.6255
R2624 VDD.n75 VDD.t1818 1.6255
R2625 VDD.n1016 VDD.t1139 1.6255
R2626 VDD.n1016 VDD.t1836 1.6255
R2627 VDD.n1017 VDD.t1830 1.6255
R2628 VDD.n1017 VDD.t783 1.6255
R2629 VDD.n1033 VDD.t635 1.6255
R2630 VDD.n1033 VDD.t2037 1.6255
R2631 VDD.n1032 VDD.t2045 1.6255
R2632 VDD.n1032 VDD.t1103 1.6255
R2633 VDD.n986 VDD.t1059 1.6255
R2634 VDD.n986 VDD.t1078 1.6255
R2635 VDD.n987 VDD.t1108 1.6255
R2636 VDD.n987 VDD.t1088 1.6255
R2637 VDD.n984 VDD.t520 1.6255
R2638 VDD.n984 VDD.t939 1.6255
R2639 VDD.n985 VDD.t935 1.6255
R2640 VDD.n985 VDD.t516 1.6255
R2641 VDD.n1048 VDD.t2055 1.6255
R2642 VDD.n1048 VDD.t1141 1.6255
R2643 VDD.n1049 VDD.t375 1.6255
R2644 VDD.n1049 VDD.t2049 1.6255
R2645 VDD.n968 VDD.t937 1.6255
R2646 VDD.n968 VDD.t597 1.6255
R2647 VDD.n971 VDD.t545 1.6255
R2648 VDD.n971 VDD.t572 1.6255
R2649 VDD.n974 VDD.t539 1.6255
R2650 VDD.n974 VDD.t541 1.6255
R2651 VDD.n982 VDD.t692 1.6255
R2652 VDD.n982 VDD.t698 1.6255
R2653 VDD.n116 VDD.t2161 1.6255
R2654 VDD.n116 VDD.t876 1.6255
R2655 VDD.n115 VDD.t882 1.6255
R2656 VDD.n115 VDD.t1315 1.6255
R2657 VDD.n1592 VDD.t1553 1.6255
R2658 VDD.n1592 VDD.t1192 1.6255
R2659 VDD.n1591 VDD.t1174 1.6255
R2660 VDD.n1591 VDD.t1345 1.6255
R2661 VDD.n1574 VDD.t1172 1.6255
R2662 VDD.n1574 VDD.t1339 1.6255
R2663 VDD.n1573 VDD.t322 1.6255
R2664 VDD.n1573 VDD.t1190 1.6255
R2665 VDD.n1552 VDD.t58 1.6255
R2666 VDD.n1552 VDD.t870 1.6255
R2667 VDD.n1551 VDD.t884 1.6255
R2668 VDD.n1551 VDD.t1313 1.6255
R2669 VDD.n135 VDD.t1373 1.6255
R2670 VDD.n135 VDD.t1316 1.6255
R2671 VDD.n136 VDD.t1372 1.6255
R2672 VDD.n136 VDD.t1309 1.6255
R2673 VDD.n1522 VDD.t628 1.6255
R2674 VDD.n1522 VDD.t632 1.6255
R2675 VDD.n1547 VDD.t729 1.6255
R2676 VDD.n1547 VDD.t1447 1.6255
R2677 VDD.n1546 VDD.t1450 1.6255
R2678 VDD.n1546 VDD.t728 1.6255
R2679 VDD.n1543 VDD.t1380 1.6255
R2680 VDD.n1543 VDD.t1322 1.6255
R2681 VDD.n1544 VDD.t1376 1.6255
R2682 VDD.n1544 VDD.t1321 1.6255
R2683 VDD.n1560 VDD.t1384 1.6255
R2684 VDD.n1560 VDD.t1333 1.6255
R2685 VDD.n1559 VDD.t1370 1.6255
R2686 VDD.n1559 VDD.t1307 1.6255
R2687 VDD.n1541 VDD.t1867 1.6255
R2688 VDD.n1541 VDD.t267 1.6255
R2689 VDD.n1540 VDD.t385 1.6255
R2690 VDD.n1540 VDD.t1866 1.6255
R2691 VDD.n1538 VDD.t927 1.6255
R2692 VDD.n1538 VDD.t929 1.6255
R2693 VDD.n1530 VDD.t440 1.6255
R2694 VDD.n1530 VDD.t2024 1.6255
R2695 VDD.n1533 VDD.t437 1.6255
R2696 VDD.n1533 VDD.t442 1.6255
R2697 VDD.n131 VDD.t1865 1.6255
R2698 VDD.n131 VDD.t148 1.6255
R2699 VDD.n90 VDD.t721 1.6255
R2700 VDD.n90 VDD.t720 1.6255
R2701 VDD.n92 VDD.t714 1.6255
R2702 VDD.n92 VDD.t753 1.6255
R2703 VDD.n93 VDD.t755 1.6255
R2704 VDD.n93 VDD.t366 1.6255
R2705 VDD.n94 VDD.t1374 1.6255
R2706 VDD.n94 VDD.t1320 1.6255
R2707 VDD.n95 VDD.t1311 1.6255
R2708 VDD.n95 VDD.t1359 1.6255
R2709 VDD.n102 VDD.t224 1.6255
R2710 VDD.n102 VDD.t222 1.6255
R2711 VDD.n104 VDD.t245 1.6255
R2712 VDD.n104 VDD.t1521 1.6255
R2713 VDD.n105 VDD.t1547 1.6255
R2714 VDD.n105 VDD.t482 1.6255
R2715 VDD.n106 VDD.t1382 1.6255
R2716 VDD.n106 VDD.t1330 1.6255
R2717 VDD.n107 VDD.t1378 1.6255
R2718 VDD.n107 VDD.t1368 1.6255
R2719 VDD.n996 VDD.t1112 1.6255
R2720 VDD.n996 VDD.t1073 1.6255
R2721 VDD.n997 VDD.t1146 1.6255
R2722 VDD.n997 VDD.t1027 1.6255
R2723 VDD.n999 VDD.t1025 1.6255
R2724 VDD.n999 VDD.t988 1.6255
R2725 VDD.n1000 VDD.t990 1.6255
R2726 VDD.n1000 VDD.t269 1.6255
R2727 VDD.n1002 VDD.t645 1.6255
R2728 VDD.n1002 VDD.t647 1.6255
R2729 VDD.n82 VDD.t2124 1.6255
R2730 VDD.n82 VDD.t1625 1.6255
R2731 VDD.n85 VDD.t1628 1.6255
R2732 VDD.n85 VDD.t1626 1.6255
R2733 VDD.n79 VDD.t656 1.6255
R2734 VDD.n79 VDD.t992 1.6255
R2735 VDD.n70 VDD.t585 1.6255
R2736 VDD.n70 VDD.t583 1.6255
R2737 VDD.n73 VDD.t605 1.6255
R2738 VDD.n73 VDD.t579 1.6255
R2739 VDD.n72 VDD.t524 1.6255
R2740 VDD.n72 VDD.t603 1.6255
R2741 VDD.n1620 VDD.t1402 1.6255
R2742 VDD.n1620 VDD.t328 1.6255
R2743 VDD.n1619 VDD.t1759 1.6255
R2744 VDD.n1619 VDD.t1404 1.6255
R2745 VDD.n1461 VDD.t289 1.6255
R2746 VDD.n1461 VDD.t286 1.6255
R2747 VDD.n1635 VDD.t846 1.6255
R2748 VDD.n1635 VDD.t2020 1.6255
R2749 VDD.n1634 VDD.t1761 1.6255
R2750 VDD.n1634 VDD.t880 1.6255
R2751 VDD.n49 VDD.t1775 1.6255
R2752 VDD.n49 VDD.t1743 1.6255
R2753 VDD.n48 VDD.t1769 1.6255
R2754 VDD.n48 VDD.t1754 1.6255
R2755 VDD.n52 VDD.t1252 1.6255
R2756 VDD.n52 VDD.t1219 1.6255
R2757 VDD.n51 VDD.t118 1.6255
R2758 VDD.n51 VDD.t1233 1.6255
R2759 VDD.n54 VDD.t1224 1.6255
R2760 VDD.n54 VDD.t1222 1.6255
R2761 VDD.n62 VDD.t1723 1.6255
R2762 VDD.n62 VDD.t1737 1.6255
R2763 VDD.n61 VDD.t1755 1.6255
R2764 VDD.n61 VDD.t1764 1.6255
R2765 VDD.n1464 VDD.t668 1.6255
R2766 VDD.n1464 VDD.t492 1.6255
R2767 VDD.n1463 VDD.t486 1.6255
R2768 VDD.n1463 VDD.t670 1.6255
R2769 VDD.n907 VDD.t1731 1.6255
R2770 VDD.n907 VDD.t1398 1.6255
R2771 VDD.n908 VDD.t1392 1.6255
R2772 VDD.n908 VDD.t454 1.6255
R2773 VDD.n850 VDD.t1765 1.6255
R2774 VDD.n850 VDD.t1744 1.6255
R2775 VDD.n851 VDD.t1763 1.6255
R2776 VDD.n851 VDD.t1734 1.6255
R2777 VDD.n853 VDD.t2015 1.6255
R2778 VDD.n853 VDD.t49 1.6255
R2779 VDD.n854 VDD.t53 1.6255
R2780 VDD.n854 VDD.t559 1.6255
R2781 VDD.n856 VDD.t81 1.6255
R2782 VDD.n856 VDD.t83 1.6255
R2783 VDD.n859 VDD.t201 1.6255
R2784 VDD.n859 VDD.t450 1.6255
R2785 VDD.n862 VDD.t446 1.6255
R2786 VDD.n862 VDD.t449 1.6255
R2787 VDD.n64 VDD.t619 1.6255
R2788 VDD.n64 VDD.t51 1.6255
R2789 VDD.n891 VDD.t1079 1.6255
R2790 VDD.n891 VDD.t1099 1.6255
R2791 VDD.n890 VDD.t1045 1.6255
R2792 VDD.n890 VDD.t1061 1.6255
R2793 VDD.n867 VDD.t292 1.6255
R2794 VDD.n867 VDD.t290 1.6255
R2795 VDD.n870 VDD.t1994 1.6255
R2796 VDD.n870 VDD.t74 1.6255
R2797 VDD.n869 VDD.t1592 1.6255
R2798 VDD.n869 VDD.t2000 1.6255
R2799 VDD.n872 VDD.t1114 1.6255
R2800 VDD.n872 VDD.t1074 1.6255
R2801 VDD.n871 VDD.t1086 1.6255
R2802 VDD.n871 VDD.t1043 1.6255
R2803 VDD.n141 VDD.t184 1.6255
R2804 VDD.n141 VDD.t186 1.6255
R2805 VDD.n139 VDD.t685 1.6255
R2806 VDD.n139 VDD.t69 1.6255
R2807 VDD.n138 VDD.t67 1.6255
R2808 VDD.n138 VDD.t243 1.6255
R2809 VDD.n1473 VDD.t1605 1.6255
R2810 VDD.n1473 VDD.t1196 1.6255
R2811 VDD.n1476 VDD.t1604 1.6255
R2812 VDD.n1476 VDD.t1602 1.6255
R2813 VDD.n153 VDD.t62 1.6255
R2814 VDD.n153 VDD.t459 1.6255
R2815 VDD.n1481 VDD.t922 1.6255
R2816 VDD.n1481 VDD.t919 1.6255
R2817 VDD.n1484 VDD.t65 1.6255
R2818 VDD.n1484 VDD.t496 1.6255
R2819 VDD.n1483 VDD.t914 1.6255
R2820 VDD.n1483 VDD.t60 1.6255
R2821 VDD.n25 VDD.t1284 1.6255
R2822 VDD.n25 VDD.t1290 1.6255
R2823 VDD.n24 VDD.t1268 1.6255
R2824 VDD.n24 VDD.t1280 1.6255
R2825 VDD.n19 VDD.t1000 1.6255
R2826 VDD.n19 VDD.t1001 1.6255
R2827 VDD.n18 VDD.t995 1.6255
R2828 VDD.n18 VDD.t997 1.6255
R2829 VDD.n30 VDD.t498 1.6255
R2830 VDD.n30 VDD.t1303 1.6255
R2831 VDD.n34 VDD.t409 1.6255
R2832 VDD.n34 VDD.t412 1.6255
R2833 VDD.n941 VDD.t178 1.6255
R2834 VDD.n941 VDD.t1557 1.6255
R2835 VDD.n942 VDD.t2176 1.6255
R2836 VDD.n942 VDD.t180 1.6255
R2837 VDD.n1073 VDD.t353 1.6255
R2838 VDD.n1073 VDD.t1805 1.6255
R2839 VDD.n1072 VDD.t1781 1.6255
R2840 VDD.n1072 VDD.t1709 1.6255
R2841 VDD.n839 VDD.t1738 1.6255
R2842 VDD.n839 VDD.t1745 1.6255
R2843 VDD.n840 VDD.t1729 1.6255
R2844 VDD.n840 VDD.t1741 1.6255
R2845 VDD.n1070 VDD.t93 1.6255
R2846 VDD.n1070 VDD.t1699 1.6255
R2847 VDD.n1071 VDD.t1701 1.6255
R2848 VDD.n1071 VDD.t27 1.6255
R2849 VDD.n1068 VDD.t94 1.6255
R2850 VDD.n1068 VDD.t97 1.6255
R2851 VDD.n933 VDD.t1702 1.6255
R2852 VDD.n933 VDD.t1870 1.6255
R2853 VDD.n928 VDD.t158 1.6255
R2854 VDD.n928 VDD.t2166 1.6255
R2855 VDD.n931 VDD.t157 1.6255
R2856 VDD.n931 VDD.t155 1.6255
R2857 VDD.n605 VDD.t1474 1.6255
R2858 VDD.n605 VDD.t1458 1.6255
R2859 VDD.n712 VDD.t852 1.6255
R2860 VDD.n712 VDD.t900 1.6255
R2861 VDD.n713 VDD.t954 1.6255
R2862 VDD.n713 VDD.t952 1.6255
R2863 VDD.n710 VDD.t508 1.6255
R2864 VDD.n710 VDD.t504 1.6255
R2865 VDD.n709 VDD.t976 1.6255
R2866 VDD.n709 VDD.t980 1.6255
R2867 VDD.n707 VDD.t868 1.6255
R2868 VDD.n707 VDD.t906 1.6255
R2869 VDD.n755 VDD.t2149 1.6255
R2870 VDD.n755 VDD.t1651 1.6255
R2871 VDD.n753 VDD.t1638 1.6255
R2872 VDD.n753 VDD.t315 1.6255
R2873 VDD.n751 VDD.t2148 1.6255
R2874 VDD.n751 VDD.t1650 1.6255
R2875 VDD.n750 VDD.t1639 1.6255
R2876 VDD.n750 VDD.t314 1.6255
R2877 VDD.n757 VDD.t1299 1.6255
R2878 VDD.n757 VDD.t1260 1.6255
R2879 VDD.n768 VDD.t1533 1.6255
R2880 VDD.n768 VDD.t1531 1.6255
R2881 VDD.n769 VDD.t1540 1.6255
R2882 VDD.n769 VDD.t1539 1.6255
R2883 VDD.n704 VDD.t896 1.6255
R2884 VDD.n704 VDD.t1906 1.6255
R2885 VDD.n608 VDD.t683 1.6255
R2886 VDD.n608 VDD.t679 1.6255
R2887 VDD.n617 VDD.t1106 1.6255
R2888 VDD.n617 VDD.t1115 1.6255
R2889 VDD.n616 VDD.t1070 1.6255
R2890 VDD.n616 VDD.t1090 1.6255
R2891 VDD.n627 VDD.t2077 1.6255
R2892 VDD.n627 VDD.t557 1.6255
R2893 VDD.n626 VDD.t1053 1.6255
R2894 VDD.n626 VDD.t2075 1.6255
R2895 VDD.n696 VDD.t1124 1.6255
R2896 VDD.n696 VDD.t2083 1.6255
R2897 VDD.n697 VDD.t2095 1.6255
R2898 VDD.n697 VDD.t665 1.6255
R2899 VDD.n667 VDD.t1144 1.6255
R2900 VDD.n667 VDD.t893 1.6255
R2901 VDD.n668 VDD.t904 1.6255
R2902 VDD.n668 VDD.t297 1.6255
R2903 VDD.n646 VDD.t1587 1.6255
R2904 VDD.n646 VDD.t627 1.6255
R2905 VDD.n647 VDD.t625 1.6255
R2906 VDD.n647 VDD.t565 1.6255
R2907 VDD.n649 VDD.t428 1.6255
R2908 VDD.n649 VDD.t430 1.6255
R2909 VDD.n659 VDD.t1105 1.6255
R2910 VDD.n659 VDD.t1113 1.6255
R2911 VDD.n660 VDD.t1126 1.6255
R2912 VDD.n660 VDD.t1101 1.6255
R2913 VDD.n662 VDD.t512 1.6255
R2914 VDD.n662 VDD.t1692 1.6255
R2915 VDD.n663 VDD.t1685 1.6255
R2916 VDD.n663 VDD.t761 1.6255
R2917 VDD.n655 VDD.t115 1.6255
R2918 VDD.n655 VDD.t112 1.6255
R2919 VDD.n682 VDD.t1084 1.6255
R2920 VDD.n682 VDD.t1076 1.6255
R2921 VDD.n683 VDD.t1137 1.6255
R2922 VDD.n683 VDD.t1125 1.6255
R2923 VDD.n642 VDD.t709 1.6255
R2924 VDD.n642 VDD.t943 1.6255
R2925 VDD.n637 VDD.t1203 1.6255
R2926 VDD.n637 VDD.t533 1.6255
R2927 VDD.n640 VDD.t528 1.6255
R2928 VDD.n640 VDD.t530 1.6255
R2929 VDD.n612 VDD.t674 1.6255
R2930 VDD.n612 VDD.t673 1.6255
R2931 VDD.n614 VDD.t941 1.6255
R2932 VDD.n614 VDD.t282 1.6255
R2933 VDD.n615 VDD.t1640 1.6255
R2934 VDD.n615 VDD.t940 1.6255
R2935 VDD.n718 VDD.t972 1.6255
R2936 VDD.n718 VDD.t974 1.6255
R2937 VDD.n714 VDD.t1262 1.6255
R2938 VDD.n714 VDD.t1264 1.6255
R2939 VDD.n919 VDD.t1065 1.6255
R2940 VDD.n919 VDD.t1080 1.6255
R2941 VDD.n918 VDD.t1035 1.6255
R2942 VDD.n918 VDD.t1047 1.6255
R2943 VDD.n921 VDD.t1859 1.6255
R2944 VDD.n921 VDD.t1582 1.6255
R2945 VDD.n922 VDD.t36 1.6255
R2946 VDD.n922 VDD.t1850 1.6255
R2947 VDD.n924 VDD.t41 1.6255
R2948 VDD.n924 VDD.t38 1.6255
R2949 VDD.n954 VDD.t1064 1.6255
R2950 VDD.n954 VDD.t1116 1.6255
R2951 VDD.n953 VDD.t1033 1.6255
R2952 VDD.n953 VDD.t1092 1.6255
R2953 VDD.n956 VDD.t275 1.6255
R2954 VDD.n956 VDD.t1648 1.6255
R2955 VDD.n957 VDD.t277 1.6255
R2956 VDD.n957 VDD.t273 1.6255
R2957 VDD.n959 VDD.t357 1.6255
R2958 VDD.n959 VDD.t355 1.6255
R2959 VDD.n781 VDD.t1439 1.6255
R2960 VDD.n781 VDD.t1453 1.6255
R2961 VDD.n782 VDD.t1443 1.6255
R2962 VDD.n782 VDD.t1430 1.6255
R2963 VDD.n177 VDD.t166 1.6255
R2964 VDD.n177 VDD.t1863 1.6255
R2965 VDD.n176 VDD.t1861 1.6255
R2966 VDD.n176 VDD.t162 1.6255
R2967 VDD.n184 VDD.t1184 1.6255
R2968 VDD.n184 VDD.t1186 1.6255
R2969 VDD.n185 VDD.t1536 1.6255
R2970 VDD.n185 VDD.t1541 1.6255
R2971 VDD.n186 VDD.t141 1.6255
R2972 VDD.n186 VDD.t139 1.6255
R2973 VDD.n190 VDD.t1526 1.6255
R2974 VDD.n190 VDD.t1535 1.6255
R2975 VDD.n191 VDD.t1826 1.6255
R2976 VDD.n191 VDD.t1832 1.6255
R2977 VDD.n195 VDD.t2002 1.6255
R2978 VDD.n195 VDD.t2009 1.6255
R2979 VDD.n196 VDD.t6 1.6255
R2980 VDD.n196 VDD.t4 1.6255
R2981 VDD.n198 VDD.t2013 1.6255
R2982 VDD.n198 VDD.t1993 1.6255
R2983 VDD.n201 VDD.t1966 1.6255
R2984 VDD.n201 VDD.t1958 1.6255
R2985 VDD.n203 VDD.t1448 1.6255
R2986 VDD.n203 VDD.t1433 1.6255
R2987 VDD.n204 VDD.t176 1.6255
R2988 VDD.n204 VDD.t174 1.6255
R2989 VDD.n207 VDD.t1442 1.6255
R2990 VDD.n207 VDD.t1445 1.6255
R2991 VDD.n208 VDD.t1807 1.6255
R2992 VDD.n208 VDD.t1790 1.6255
R2993 VDD.n212 VDD.t2141 1.6255
R2994 VDD.n212 VDD.t2127 1.6255
R2995 VDD.n213 VDD.t433 1.6255
R2996 VDD.n213 VDD.t435 1.6255
R2997 VDD.n215 VDD.t2138 1.6255
R2998 VDD.n215 VDD.t2140 1.6255
R2999 VDD.n218 VDD.t1683 1.6255
R3000 VDD.n218 VDD.t1672 1.6255
R3001 VDD.n222 VDD.t805 1.6255
R3002 VDD.n222 VDD.t803 1.6255
R3003 VDD.n221 VDD.t1690 1.6255
R3004 VDD.n221 VDD.t1680 1.6255
R3005 VDD.n235 VDD.t2093 1.6255
R3006 VDD.n235 VDD.t2073 1.6255
R3007 VDD.n234 VDD.t1848 1.6255
R3008 VDD.n234 VDD.t1856 1.6255
R3009 VDD.n232 VDD.t326 1.6255
R3010 VDD.n232 VDD.t324 1.6255
R3011 VDD.n231 VDD.t1858 1.6255
R3012 VDD.n231 VDD.t1842 1.6255
R3013 VDD.n224 VDD.t2053 1.6255
R3014 VDD.n224 VDD.t2039 1.6255
R3015 VDD.n225 VDD.t1239 1.6255
R3016 VDD.n225 VDD.t1248 1.6255
R3017 VDD.n244 VDD.t305 1.6255
R3018 VDD.n244 VDD.t303 1.6255
R3019 VDD.n243 VDD.t1254 1.6255
R3020 VDD.n243 VDD.t1229 1.6255
R3021 VDD.n246 VDD.t1406 1.6255
R3022 VDD.n246 VDD.t1388 1.6255
R3023 VDD.n1343 VDD.t740 1.6255
R3024 VDD.n1343 VDD.t2071 1.6255
R3025 VDD.n1341 VDD.t126 1.6255
R3026 VDD.n1341 VDD.t307 1.6255
R3027 VDD.n1339 VDD.t741 1.6255
R3028 VDD.n1339 VDD.t2070 1.6255
R3029 VDD.n1338 VDD.t125 1.6255
R3030 VDD.n1338 VDD.t308 1.6255
R3031 VDD.n256 VDD.t747 1.6255
R3032 VDD.n256 VDD.t1479 1.6255
R3033 VDD.n254 VDD.t122 1.6255
R3034 VDD.n254 VDD.t744 1.6255
R3035 VDD.n252 VDD.t746 1.6255
R3036 VDD.n252 VDD.t1478 1.6255
R3037 VDD.n251 VDD.t123 1.6255
R3038 VDD.n251 VDD.t743 1.6255
R3039 VDD.n290 VDD.t1422 1.6255
R3040 VDD.n290 VDD.t1659 1.6255
R3041 VDD.n293 VDD.t336 1.6255
R3042 VDD.n293 VDD.t342 1.6255
R3043 VDD.n292 VDD.t1511 1.6255
R3044 VDD.n292 VDD.t1513 1.6255
R3045 VDD.n295 VDD.t1663 1.6255
R3046 VDD.n295 VDD.t1426 1.6255
R3047 VDD.n296 VDD.t1985 1.6255
R3048 VDD.n296 VDD.t1987 1.6255
R3049 VDD.n297 VDD.t1946 1.6255
R3050 VDD.n297 VDD.t1948 1.6255
R3051 VDD.n301 VDD.t1509 1.6255
R3052 VDD.n301 VDD.t1515 1.6255
R3053 VDD.n303 VDD.t392 1.6255
R3054 VDD.n303 VDD.t398 1.6255
R3055 VDD.n304 VDD.t1653 1.6255
R3056 VDD.n304 VDD.t1665 1.6255
R3057 VDD.n347 VDD.t1469 1.6255
R3058 VDD.n347 VDD.t1472 1.6255
R3059 VDD.n270 VDD.t2103 1.6255
R3060 VDD.n270 VDD.t2099 1.6255
R3061 VDD.n271 VDD.t421 1.6255
R3062 VDD.n271 VDD.t419 1.6255
R3063 VDD.n274 VDD.t842 1.6255
R3064 VDD.n274 VDD.t866 1.6255
R3065 VDD.n273 VDD.t826 1.6255
R3066 VDD.n273 VDD.t848 1.6255
R3067 VDD.n460 VDD.t1809 1.6255
R3068 VDD.n460 VDD.t1783 1.6255
R3069 VDD.n459 VDD.t1609 1.6255
R3070 VDD.n459 VDD.t910 1.6255
R3071 VDD.n458 VDD.t912 1.6255
R3072 VDD.n458 VDD.t1922 1.6255
R3073 VDD.n457 VDD.t464 1.6255
R3074 VDD.n457 VDD.t106 1.6255
R3075 VDD.n456 VDD.t104 1.6255
R3076 VDD.n456 VDD.t553 1.6255
R3077 VDD.n455 VDD.t1178 1.6255
R3078 VDD.n455 VDD.t1182 1.6255
R3079 VDD.n451 VDD.t1524 1.6255
R3080 VDD.n451 VDD.t1529 1.6255
R3081 VDD.n452 VDD.t239 1.6255
R3082 VDD.n452 VDD.t237 1.6255
R3083 VDD.n450 VDD.t1545 1.6255
R3084 VDD.n450 VDD.t1523 1.6255
R3085 VDD.n448 VDD.t1820 1.6255
R3086 VDD.n448 VDD.t1828 1.6255
R3087 VDD.n445 VDD.t1995 1.6255
R3088 VDD.n445 VDD.t2001 1.6255
R3089 VDD.n446 VDD.t601 1.6255
R3090 VDD.n446 VDD.t599 1.6255
R3091 VDD.n443 VDD.t2004 1.6255
R3092 VDD.n443 VDD.t2011 1.6255
R3093 VDD.n442 VDD.t1960 1.6255
R3094 VDD.n442 VDD.t1968 1.6255
R3095 VDD.n438 VDD.t1440 1.6255
R3096 VDD.n438 VDD.t1456 1.6255
R3097 VDD.n439 VDD.t299 1.6255
R3098 VDD.n439 VDD.t301 1.6255
R3099 VDD.n437 VDD.t1428 1.6255
R3100 VDD.n437 VDD.t1435 1.6255
R3101 VDD.n435 VDD.t2033 1.6255
R3102 VDD.n435 VDD.t2035 1.6255
R3103 VDD.n432 VDD.t2132 1.6255
R3104 VDD.n432 VDD.t2146 1.6255
R3105 VDD.n433 VDD.t768 1.6255
R3106 VDD.n433 VDD.t770 1.6255
R3107 VDD.n430 VDD.t2126 1.6255
R3108 VDD.n430 VDD.t2129 1.6255
R3109 VDD.n427 VDD.t1677 1.6255
R3110 VDD.n427 VDD.t1687 1.6255
R3111 VDD.n425 VDD.t1634 1.6255
R3112 VDD.n425 VDD.t1636 1.6255
R3113 VDD.n424 VDD.t1681 1.6255
R3114 VDD.n424 VDD.t1695 1.6255
R3115 VDD.n416 VDD.t2085 1.6255
R3116 VDD.n416 VDD.t2091 1.6255
R3117 VDD.n415 VDD.t1844 1.6255
R3118 VDD.n415 VDD.t1846 1.6255
R3119 VDD.n413 VDD.t23 1.6255
R3120 VDD.n413 VDD.t25 1.6255
R3121 VDD.n412 VDD.t1849 1.6255
R3122 VDD.n412 VDD.t1857 1.6255
R3123 VDD.n405 VDD.t2043 1.6255
R3124 VDD.n405 VDD.t2057 1.6255
R3125 VDD.n406 VDD.t1226 1.6255
R3126 VDD.n406 VDD.t1237 1.6255
R3127 VDD.n398 VDD.t1936 1.6255
R3128 VDD.n398 VDD.t1935 1.6255
R3129 VDD.n397 VDD.t1244 1.6255
R3130 VDD.n397 VDD.t1250 1.6255
R3131 VDD.n400 VDD.t1394 1.6255
R3132 VDD.n400 VDD.t1408 1.6255
R3133 VDD.n392 VDD.t766 1.6255
R3134 VDD.n392 VDD.t1420 1.6255
R3135 VDD.n390 VDD.t1618 1.6255
R3136 VDD.n390 VDD.t700 1.6255
R3137 VDD.n388 VDD.t765 1.6255
R3138 VDD.n388 VDD.t1419 1.6255
R3139 VDD.n387 VDD.t1619 1.6255
R3140 VDD.n387 VDD.t701 1.6255
R3141 VDD.n384 VDD.t479 1.6255
R3142 VDD.n384 VDD.t1875 1.6255
R3143 VDD.n382 VDD.t469 1.6255
R3144 VDD.n382 VDD.t651 1.6255
R3145 VDD.n380 VDD.t480 1.6255
R3146 VDD.n380 VDD.t1874 1.6255
R3147 VDD.n379 VDD.t468 1.6255
R3148 VDD.n379 VDD.t652 1.6255
R3149 VDD.n278 VDD.t2111 1.6255
R3150 VDD.n278 VDD.t2101 1.6255
R3151 VDD.n369 VDD.t2115 1.6255
R3152 VDD.n369 VDD.t2113 1.6255
R3153 VDD.n363 VDD.t830 1.6255
R3154 VDD.n363 VDD.t872 1.6255
R3155 VDD.n280 VDD.t1980 1.6255
R3156 VDD.n280 VDD.t1976 1.6255
R3157 VDD.n282 VDD.t1485 1.6255
R3158 VDD.n282 VDD.t1483 1.6255
R3159 VDD.n264 VDD.t1910 1.6255
R3160 VDD.n264 VDD.t1897 1.6255
R3161 VDD.n265 VDD.t1012 1.6255
R3162 VDD.n265 VDD.t1014 1.6255
R3163 VDD.n267 VDD.t2063 1.6255
R3164 VDD.n267 VDD.t2068 1.6255
R3165 VDD.n566 VDD.t1491 1.6255
R3166 VDD.n566 VDD.t1497 1.6255
R3167 VDD.n568 VDD.t1004 1.6255
R3168 VDD.n568 VDD.t1006 1.6255
R3169 VDD.n569 VDD.t878 1.6255
R3170 VDD.n569 VDD.t1903 1.6255
R3171 VDD.n262 VDD.t801 1.6255
R3172 VDD.n262 VDD.t797 1.6255
R3173 VDD.n261 VDD.t1493 1.6255
R3174 VDD.n261 VDD.t1499 1.6255
R3175 VDD.n259 VDD.t1912 1.6255
R3176 VDD.n259 VDD.t818 1.6255
R3177 VDD.n1281 VDD.t824 1.6255
R3178 VDD.n1281 VDD.t834 1.6255
R3179 VDD.n1267 VDD.t1215 1.6255
R3180 VDD.n1267 VDD.t1213 1.6255
R3181 VDD.n1250 VDD.t1938 1.6255
R3182 VDD.n1250 VDD.t1796 1.6255
R3183 VDD.n1251 VDD.t926 1.6255
R3184 VDD.n1251 VDD.t1944 1.6255
R3185 VDD.n598 VDD.t613 1.6255
R3186 VDD.n598 VDD.t611 1.6255
R3187 VDD.n601 VDD.t1152 1.6255
R3188 VDD.n601 VDD.t705 1.6255
R3189 VDD.n600 VDD.t588 1.6255
R3190 VDD.n600 VDD.t1150 1.6255
R3191 VDD.n593 VDD.t1777 1.6255
R3192 VDD.n593 VDD.t1785 1.6255
R3193 VDD.n592 VDD.t1786 1.6255
R3194 VDD.n592 VDD.t1799 1.6255
R3195 VDD.n1189 VDD.t1565 1.6255
R3196 VDD.n1189 VDD.t1575 1.6255
R3197 VDD.n1192 VDD.t249 1.6255
R3198 VDD.n1192 VDD.t253 1.6255
R3199 VDD.n1191 VDD.t1883 1.6255
R3200 VDD.n1191 VDD.t1887 1.6255
R3201 VDD.n1194 VDD.t1573 1.6255
R3202 VDD.n1194 VDD.t1577 1.6255
R3203 VDD.n1195 VDD.t1164 1.6255
R3204 VDD.n1195 VDD.t1166 1.6255
R3205 VDD.n1278 VDD.n1277 1.61677
R3206 VDD.n738 VDD.n737 1.61677
R3207 VDD.n333 VDD.n332 1.61677
R3208 VDD.n1324 VDD.n1323 1.61677
R3209 VDD.n1237 VDD.n1236 1.61677
R3210 VDD.t1864 VDD.t68 1.55813
R3211 VDD.t147 VDD.t66 1.55813
R3212 VDD.t145 VDD.t242 1.55813
R3213 VDD.n1588 VDD.t2026 1.55813
R3214 VDD.n1616 VDD.t203 1.55732
R3215 VDD.t523 VDD.t620 1.55732
R3216 VDD.t602 VDD.t618 1.55732
R3217 VDD.t604 VDD.t50 1.55732
R3218 VDD.t1696 VDD.t272 1.55732
R3219 VDD.t1869 VDD.t274 1.55732
R3220 VDD.t1871 VDD.t1647 1.55732
R3221 VDD.n1063 VDD.t2164 1.55732
R3222 VDD.n351 VDD.n287 1.5398
R3223 VDD.n1248 VDD.n1247 1.47379
R3224 VDD.n1372 VDD.n220 1.3355
R3225 VDD.n519 VDD.n429 1.3355
R3226 VDD.t436 VDD.t1371 1.30089
R3227 VDD.t441 VDD.t1308 1.30089
R3228 VDD.t1347 VDD.t438 1.30089
R3229 VDD.t1030 VDD.t198 1.30033
R3230 VDD.t1044 VDD.t200 1.30033
R3231 VDD.t1060 VDD.t448 1.30033
R3232 VDD.t156 VDD.t1032 1.30033
R3233 VDD.t154 VDD.t1091 1.30033
R3234 VDD.t152 VDD.t1093 1.30033
R3235 VDD.n747 VDD.n706 1.22931
R3236 VDD.n1359 VDD 1.21734
R3237 VDD VDD.n532 1.21734
R3238 VDD.n1367 VDD 1.20815
R3239 VDD VDD.n524 1.20815
R3240 VDD.n1354 VDD.n1353 1.16958
R3241 VDD.n538 VDD.n537 1.16958
R3242 VDD.n1103 VDD.n1102 1.15088
R3243 VDD.n1366 VDD 1.13101
R3244 VDD.n525 VDD 1.13101
R3245 VDD.n1162 VDD.n1135 1.11767
R3246 VDD.n555 VDD.n554 1.10294
R3247 VDD.n1456 VDD.n1455 1.08484
R3248 VDD.n1416 VDD.n1415 1.07484
R3249 VDD.n1458 VDD.n1457 0.985783
R3250 VDD.n1102 VDD.n175 0.98484
R3251 VDD.n1665 VDD.n1664 0.969146
R3252 VDD.n1585 VDD.n1584 0.969146
R3253 VDD.n100 VDD.n98 0.969146
R3254 VDD.n60 VDD.n59 0.969146
R3255 VDD.n889 VDD.n888 0.969146
R3256 VDD.n681 VDD.n680 0.969146
R3257 VDD.n1060 VDD.n1059 0.969146
R3258 VDD.n970 VDD.n969 0.947457
R3259 VDD.n133 VDD.n132 0.947457
R3260 VDD.n81 VDD.n80 0.947457
R3261 VDD.n66 VDD.n65 0.947457
R3262 VDD.n155 VDD.n154 0.947457
R3263 VDD.n935 VDD.n934 0.947457
R3264 VDD.n776 VDD.n775 0.947457
R3265 VDD.n777 VDD.n776 0.947457
R3266 VDD.n778 VDD.n777 0.947457
R3267 VDD.n644 VDD.n643 0.947457
R3268 VDD VDD.n1227 0.894579
R3269 VDD.n1415 VDD.n175 0.888236
R3270 VDD.n1488 VDD.n1487 0.882891
R3271 VDD.n1582 VDD.n1528 0.863847
R3272 VDD VDD.n242 0.854582
R3273 VDD.n423 VDD 0.854582
R3274 VDD.n1398 VDD.n1397 0.820445
R3275 VDD.n1379 VDD.n1378 0.820445
R3276 VDD.n489 VDD.n488 0.820445
R3277 VDD.n498 VDD.n441 0.820445
R3278 VDD.n512 VDD.n511 0.820445
R3279 VDD.n980 VDD.n976 0.817542
R3280 VDD.n1536 VDD.n1535 0.817542
R3281 VDD.n1005 VDD.n87 0.817542
R3282 VDD.n865 VDD.n864 0.817542
R3283 VDD.n1479 VDD.n1478 0.817542
R3284 VDD.n1066 VDD.n1065 0.817542
R3285 VDD.n1174 VDD.n1173 0.817542
R3286 VDD.n189 VDD.n188 0.81252
R3287 VDD.n475 VDD.n454 0.81252
R3288 VDD.n779 VDD.n778 0.8105
R3289 VDD.n754 VDD.n752 0.778681
R3290 VDD.n1342 VDD.n1340 0.778681
R3291 VDD.n255 VDD.n253 0.778681
R3292 VDD.n391 VDD.n389 0.778681
R3293 VDD.n383 VDD.n381 0.778681
R3294 VDD.n771 VDD.n770 0.763264
R3295 VDD.n1659 VDD.n1658 0.752098
R3296 VDD.n1490 VDD.n1489 0.752098
R3297 VDD.n1568 VDD.n1567 0.752098
R3298 VDD.n1564 VDD.n1563 0.752098
R3299 VDD.n112 VDD.n109 0.752098
R3300 VDD.n1024 VDD.n995 0.752098
R3301 VDD.n1641 VDD.n47 0.752098
R3302 VDD.n915 VDD.n849 0.752098
R3303 VDD.n847 VDD.n846 0.752098
R3304 VDD.n844 VDD.n843 0.752098
R3305 VDD.n675 VDD.n658 0.752098
R3306 VDD.n1097 VDD.n1096 0.752098
R3307 VDD VDD.n783 0.750764
R3308 VDD.n1046 VDD.n976 0.739568
R3309 VDD.n1606 VDD.n87 0.739568
R3310 VDD.n1065 VDD.n1064 0.739568
R3311 VDD.n1173 VDD.n1172 0.739568
R3312 VDD.n1579 VDD.n1578 0.738728
R3313 VDD.n1611 VDD.n1610 0.738728
R3314 VDD.n1633 VDD.n1632 0.738728
R3315 VDD.n1466 VDD.n1465 0.738728
R3316 VDD.n882 VDD.n881 0.738728
R3317 VDD.n1502 VDD.n1501 0.738728
R3318 VDD.n1664 VDD 0.7301
R3319 VDD VDD.n980 0.7301
R3320 VDD.n1584 VDD 0.7301
R3321 VDD VDD.n1536 0.7301
R3322 VDD VDD.n100 0.7301
R3323 VDD VDD.n1005 0.7301
R3324 VDD.n59 VDD 0.7301
R3325 VDD VDD.n865 0.7301
R3326 VDD.n888 VDD 0.7301
R3327 VDD VDD.n1479 0.7301
R3328 VDD.n1671 VDD 0.7301
R3329 VDD VDD.n1066 0.7301
R3330 VDD.n680 VDD 0.7301
R3331 VDD VDD.n1174 0.7301
R3332 VDD.n1059 VDD 0.7301
R3333 VDD.n1247 VDD.n602 0.718056
R3334 VDD.n12 VDD.n11 0.715763
R3335 VDD.n1362 VDD.n242 0.70948
R3336 VDD.n529 VDD.n423 0.70948
R3337 VDD VDD.n1352 0.703633
R3338 VDD.n539 VDD 0.703633
R3339 VDD.n991 VDD.n990 0.694644
R3340 VDD.n610 VDD.n609 0.658723
R3341 VDD.n1648 VDD.n46 0.652313
R3342 VDD.n1041 VDD.n1040 0.652313
R3343 VDD.n1548 VDD.n1524 0.652313
R3344 VDD.n1580 VDD.n1579 0.652313
R3345 VDD.n1601 VDD.n1600 0.652313
R3346 VDD.n124 VDD.n123 0.652313
R3347 VDD.n1013 VDD.n1012 0.652313
R3348 VDD.n1612 VDD.n1611 0.652313
R3349 VDD.n1467 VDD.n1466 0.652313
R3350 VDD.n1632 VDD.n1631 0.652313
R3351 VDD.n904 VDD.n903 0.652313
R3352 VDD.n883 VDD.n882 0.652313
R3353 VDD.n150 VDD.n149 0.652313
R3354 VDD.n1503 VDD.n1502 0.652313
R3355 VDD.n943 VDD.n36 0.652313
R3356 VDD.n1081 VDD.n1080 0.652313
R3357 VDD.n692 VDD.n691 0.652313
R3358 VDD.n664 VDD.n657 0.652313
R3359 VDD.n635 VDD.n634 0.652313
R3360 VDD.n1086 VDD.n1085 0.652313
R3361 VDD.n965 VDD.n964 0.652313
R3362 VDD.n1259 VDD.n1258 0.652313
R3363 VDD.n1187 VDD.n606 0.651457
R3364 VDD.n1478 VDD.n1459 0.650331
R3365 VDD.n562 VDD.n561 0.649202
R3366 VDD.n1535 VDD.n134 0.646517
R3367 VDD VDD.n21 0.639914
R3368 VDD.n780 VDD.n779 0.590391
R3369 VDD.n1266 VDD.n1265 0.582689
R3370 VDD.n1681 VDD.n27 0.569616
R3371 VDD VDD.n767 0.566011
R3372 VDD VDD.n343 0.565631
R3373 VDD.n193 VDD.n192 0.561058
R3374 VDD.n483 VDD.n482 0.561058
R3375 VDD.n1180 VDD.n610 0.55925
R3376 VDD.n1047 VDD.n970 0.552239
R3377 VDD.n973 VDD.n972 0.552239
R3378 VDD.n1532 VDD.n1531 0.552239
R3379 VDD.n1590 VDD.n133 0.552239
R3380 VDD.n84 VDD.n83 0.552239
R3381 VDD.n1607 VDD.n81 0.552239
R3382 VDD.n861 VDD.n860 0.552239
R3383 VDD.n1618 VDD.n66 0.552239
R3384 VDD.n1475 VDD.n1474 0.552239
R3385 VDD.n1509 VDD.n155 0.552239
R3386 VDD.n949 VDD.n935 0.552239
R3387 VDD.n930 VDD.n929 0.552239
R3388 VDD.n702 VDD.n644 0.552239
R3389 VDD.n639 VDD.n638 0.552239
R3390 VDD.n202 VDD.n157 0.530241
R3391 VDD.n946 VDD 0.528114
R3392 VDD VDD.n1656 0.528114
R3393 VDD VDD.n1517 0.528114
R3394 VDD VDD.n1557 0.528114
R3395 VDD.n130 VDD 0.528114
R3396 VDD.n114 VDD 0.528114
R3397 VDD VDD.n1639 0.528114
R3398 VDD VDD.n1625 0.528114
R3399 VDD.n875 VDD 0.528114
R3400 VDD VDD.n673 0.528114
R3401 VDD VDD.n645 0.528114
R3402 VDD VDD.n1094 0.528114
R3403 VDD VDD.n1055 0.528114
R3404 VDD.n1358 VDD 0.513867
R3405 VDD.n1363 VDD 0.513867
R3406 VDD.n1371 VDD 0.513867
R3407 VDD.n533 VDD 0.513867
R3408 VDD VDD.n528 0.513867
R3409 VDD.n520 VDD 0.513867
R3410 VDD.n23 VDD.n21 0.512079
R3411 VDD.n1227 VDD.n1 0.512079
R3412 VDD.n11 VDD.n5 0.512079
R3413 VDD.n13 VDD.n12 0.512079
R3414 VDD.n349 VDD.n348 0.509717
R3415 VDD.n1687 VDD.n1686 0.509533
R3416 VDD.n1209 VDD.n1208 0.505435
R3417 VDD.n1305 VDD.n1304 0.505435
R3418 VDD.n1272 VDD.n588 0.505435
R3419 VDD.n740 VDD.n708 0.505435
R3420 VDD.n335 VDD.n291 0.505435
R3421 VDD.n310 VDD.n309 0.505435
R3422 VDD.n372 VDD.n371 0.505435
R3423 VDD.n575 VDD.n574 0.505435
R3424 VDD.n1326 VDD.n260 0.505435
R3425 VDD.n1239 VDD.n1190 0.505435
R3426 VDD.n1198 VDD.n1197 0.50509
R3427 VDD.n1294 VDD.n1293 0.50509
R3428 VDD.n716 VDD.n715 0.50509
R3429 VDD.n299 VDD.n298 0.50509
R3430 VDD.n361 VDD.n360 0.50509
R3431 VDD.n46 VDD.n45 0.494257
R3432 VDD.n1041 VDD.n983 0.494257
R3433 VDD.n1524 VDD.n1523 0.494257
R3434 VDD.n1580 VDD.n1539 0.494257
R3435 VDD.n1601 VDD.n91 0.494257
R3436 VDD.n124 VDD.n103 0.494257
R3437 VDD.n1012 VDD.n1003 0.494257
R3438 VDD.n1612 VDD.n71 0.494257
R3439 VDD.n1467 VDD.n1462 0.494257
R3440 VDD.n1631 VDD.n55 0.494257
R3441 VDD.n903 VDD.n857 0.494257
R3442 VDD.n883 VDD.n868 0.494257
R3443 VDD.n149 VDD.n142 0.494257
R3444 VDD.n1503 VDD.n1482 0.494257
R3445 VDD.n36 VDD.n35 0.494257
R3446 VDD.n1081 VDD.n1069 0.494257
R3447 VDD.n691 VDD.n650 0.494257
R3448 VDD.n657 VDD.n656 0.494257
R3449 VDD.n635 VDD.n613 0.494257
R3450 VDD.n1085 VDD.n925 0.494257
R3451 VDD.n964 VDD.n960 0.494257
R3452 VDD.n1259 VDD.n599 0.494257
R3453 VDD.n1649 VDD.n1648 0.490519
R3454 VDD.n1040 VDD.n1039 0.490519
R3455 VDD.n1549 VDD.n1548 0.490519
R3456 VDD.n1600 VDD.n1599 0.490519
R3457 VDD.n123 VDD.n122 0.490519
R3458 VDD.n1014 VDD.n1013 0.490519
R3459 VDD.n905 VDD.n904 0.490519
R3460 VDD.n151 VDD.n150 0.490519
R3461 VDD.n944 VDD.n943 0.490519
R3462 VDD.n1080 VDD.n1079 0.490519
R3463 VDD.n693 VDD.n692 0.490519
R3464 VDD.n665 VDD.n664 0.490519
R3465 VDD.n634 VDD.n633 0.490519
R3466 VDD.n1087 VDD.n1086 0.490519
R3467 VDD.n966 VDD.n965 0.490519
R3468 VDD.n180 VDD.n179 0.490519
R3469 VDD.n1412 VDD.n1411 0.490519
R3470 VDD.n466 VDD.n465 0.490519
R3471 VDD.n468 VDD.n467 0.490519
R3472 VDD.n470 VDD.n469 0.490519
R3473 VDD.n472 VDD.n471 0.490519
R3474 VDD.n1258 VDD.n1257 0.490519
R3475 VDD.n1249 VDD.n1248 0.487614
R3476 VDD.n765 VDD.n749 0.485854
R3477 VDD VDD.n1201 0.484396
R3478 VDD VDD.n1301 0.484396
R3479 VDD VDD.n607 0.484396
R3480 VDD VDD.n302 0.484396
R3481 VDD VDD.n368 0.484396
R3482 VDD VDD.n567 0.484396
R3483 VDD VDD.n1312 0.48089
R3484 VDD.n746 VDD 0.48089
R3485 VDD.n341 VDD 0.48089
R3486 VDD.n1332 VDD 0.48089
R3487 VDD.n1245 VDD 0.48089
R3488 VDD.n1219 VDD 0.466864
R3489 VDD VDD.n1290 0.466864
R3490 VDD.n725 VDD 0.466864
R3491 VDD.n320 VDD 0.466864
R3492 VDD.n585 VDD 0.466864
R3493 VDD.n464 VDD 0.465572
R3494 VDD.n1092 VDD 0.46531
R3495 VDD.n1654 VDD 0.46531
R3496 VDD.n1499 VDD 0.46531
R3497 VDD.n879 VDD 0.46531
R3498 VDD.n78 VDD 0.46531
R3499 VDD.n1576 VDD 0.46531
R3500 VDD VDD.n1577 0.46531
R3501 VDD VDD.n1609 0.46531
R3502 VDD.n1622 VDD 0.46531
R3503 VDD.n1637 VDD 0.46531
R3504 VDD.n1638 VDD 0.46531
R3505 VDD.n1624 VDD 0.46531
R3506 VDD VDD.n880 0.46531
R3507 VDD VDD.n1500 0.46531
R3508 VDD.n940 VDD.n939 0.460899
R3509 VDD.n1655 VDD.n1650 0.460899
R3510 VDD.n1514 VDD.n1513 0.460899
R3511 VDD.n1020 VDD.n1019 0.460899
R3512 VDD.n1036 VDD.n1035 0.460899
R3513 VDD.n1038 VDD.n1037 0.460899
R3514 VDD.n1052 VDD.n1051 0.460899
R3515 VDD.n119 VDD.n118 0.460899
R3516 VDD.n1595 VDD.n1594 0.460899
R3517 VDD.n1555 VDD.n1554 0.460899
R3518 VDD.n1556 VDD.n1550 0.460899
R3519 VDD.n1598 VDD.n1597 0.460899
R3520 VDD.n121 VDD.n120 0.460899
R3521 VDD.n1021 VDD.n1015 0.460899
R3522 VDD.n911 VDD.n910 0.460899
R3523 VDD.n912 VDD.n906 0.460899
R3524 VDD.n1516 VDD.n152 0.460899
R3525 VDD.n947 VDD.n945 0.460899
R3526 VDD.n1076 VDD.n1075 0.460899
R3527 VDD.n1078 VDD.n1077 0.460899
R3528 VDD.n630 VDD.n629 0.460899
R3529 VDD.n700 VDD.n699 0.460899
R3530 VDD.n671 VDD.n670 0.460899
R3531 VDD.n695 VDD.n694 0.460899
R3532 VDD.n672 VDD.n666 0.460899
R3533 VDD.n632 VDD.n631 0.460899
R3534 VDD.n1093 VDD.n1088 0.460899
R3535 VDD.n1054 VDD.n967 0.460899
R3536 VDD.n1254 VDD.n1253 0.460899
R3537 VDD.n1256 VDD.n1255 0.460899
R3538 VDD.n1348 VDD.n1347 0.458609
R3539 VDD.n394 VDD.n386 0.458609
R3540 VDD.n1687 VDD.n16 0.458326
R3541 VDD.n12 VDD.n9 0.458326
R3542 VDD.n5 VDD.n4 0.458326
R3543 VDD.n1227 VDD.n1226 0.458326
R3544 VDD.n1682 VDD.n26 0.458326
R3545 VDD.n21 VDD.n20 0.458326
R3546 VDD.n864 VDD.n67 0.456602
R3547 VDD.n13 VDD.n6 0.45408
R3548 VDD.n1 VDD.n0 0.45408
R3549 VDD.n23 VDD.n22 0.45408
R3550 VDD VDD.n938 0.4505
R3551 VDD VDD.n1649 0.4505
R3552 VDD VDD.n1512 0.4505
R3553 VDD VDD.n1018 0.4505
R3554 VDD VDD.n1034 0.4505
R3555 VDD.n1039 VDD 0.4505
R3556 VDD VDD.n1050 0.4505
R3557 VDD VDD.n117 0.4505
R3558 VDD VDD.n1593 0.4505
R3559 VDD VDD.n1553 0.4505
R3560 VDD VDD.n1549 0.4505
R3561 VDD.n1599 VDD 0.4505
R3562 VDD.n122 VDD 0.4505
R3563 VDD VDD.n1014 0.4505
R3564 VDD VDD.n909 0.4505
R3565 VDD VDD.n905 0.4505
R3566 VDD VDD.n151 0.4505
R3567 VDD VDD.n944 0.4505
R3568 VDD VDD.n1074 0.4505
R3569 VDD.n1079 VDD 0.4505
R3570 VDD VDD.n628 0.4505
R3571 VDD VDD.n698 0.4505
R3572 VDD VDD.n669 0.4505
R3573 VDD VDD.n693 0.4505
R3574 VDD VDD.n665 0.4505
R3575 VDD.n633 VDD 0.4505
R3576 VDD VDD.n1087 0.4505
R3577 VDD VDD.n966 0.4505
R3578 VDD VDD.n178 0.4505
R3579 VDD.n1413 VDD 0.4505
R3580 VDD VDD.n466 0.4505
R3581 VDD VDD.n470 0.4505
R3582 VDD VDD.n1252 0.4505
R3583 VDD.n1257 VDD 0.4505
R3584 VDD.n11 VDD.n10 0.450011
R3585 VDD.n899 VDD.n898 0.447328
R3586 VDD.n1414 VDD.n181 0.444278
R3587 VDD.n1686 VDD.n17 0.442185
R3588 VDD.n763 VDD.n756 0.441438
R3589 VDD.n1345 VDD.n1344 0.441438
R3590 VDD.n1337 VDD.n257 0.441438
R3591 VDD.n396 VDD.n393 0.441438
R3592 VDD.n543 VDD.n385 0.441438
R3593 VDD.n1411 VDD.n1410 0.436623
R3594 VDD.n473 VDD.n472 0.436623
R3595 VDD.n1665 VDD.n41 0.434848
R3596 VDD.n40 VDD.n39 0.434848
R3597 VDD.n1657 VDD.n1645 0.434848
R3598 VDD.n1518 VDD.n137 0.434848
R3599 VDD.n1585 VDD.n1519 0.434848
R3600 VDD.n1558 VDD.n1545 0.434848
R3601 VDD.n129 VDD.n96 0.434848
R3602 VDD.n98 VDD.n97 0.434848
R3603 VDD.n113 VDD.n108 0.434848
R3604 VDD.n1640 VDD.n50 0.434848
R3605 VDD.n1626 VDD.n63 0.434848
R3606 VDD.n60 VDD.n57 0.434848
R3607 VDD.n894 VDD.n892 0.434848
R3608 VDD.n889 VDD.n886 0.434848
R3609 VDD.n874 VDD.n873 0.434848
R3610 VDD.n674 VDD.n661 0.434848
R3611 VDD.n681 VDD.n652 0.434848
R3612 VDD.n685 VDD.n684 0.434848
R3613 VDD.n1095 VDD.n920 0.434848
R3614 VDD.n1060 VDD.n1057 0.434848
R3615 VDD.n1056 VDD.n955 0.434848
R3616 VDD.n595 VDD.n594 0.434848
R3617 VDD.n1047 VDD 0.434483
R3618 VDD.n1590 VDD 0.434483
R3619 VDD.n1607 VDD 0.434483
R3620 VDD.n1618 VDD 0.434483
R3621 VDD.n1509 VDD 0.434483
R3622 VDD VDD.n949 0.434483
R3623 VDD VDD.n702 0.434483
R3624 VDD.n989 VDD.n988 0.432891
R3625 VDD.n1023 VDD.n998 0.432891
R3626 VDD.n914 VDD.n852 0.432891
R3627 VDD.n619 VDD.n618 0.432891
R3628 VDD.n465 VDD.n464 0.421551
R3629 VDD.n1335 VDD.n1334 0.421429
R3630 VDD.n546 VDD.n545 0.421429
R3631 VDD.n625 VDD 0.417045
R3632 VDD VDD.n1022 0.40956
R3633 VDD VDD.n913 0.40956
R3634 VDD.n1031 VDD 0.408631
R3635 VDD.n1572 VDD 0.406221
R3636 VDD.n1495 VDD 0.406221
R3637 VDD.n842 VDD.n841 0.4055
R3638 VDD.n727 VDD.n726 0.401325
R3639 VDD.n322 VDD.n321 0.401325
R3640 VDD.n1221 VDD.n1220 0.401325
R3641 VDD VDD.n357 0.398508
R3642 VDD.n1397 VDD.n197 0.397674
R3643 VDD.n206 VDD.n205 0.397674
R3644 VDD.n1378 VDD.n214 0.397674
R3645 VDD.n1367 VDD.n223 0.397674
R3646 VDD.n1354 VDD.n245 0.397674
R3647 VDD.n489 VDD.n447 0.397674
R3648 VDD.n441 VDD.n440 0.397674
R3649 VDD.n512 VDD.n434 0.397674
R3650 VDD.n524 VDD.n426 0.397674
R3651 VDD.n537 VDD.n399 0.397674
R3652 VDD VDD.n785 0.39672
R3653 VDD.n189 VDD.n187 0.395717
R3654 VDD.n454 VDD.n453 0.395717
R3655 VDD.n1682 VDD.n1681 0.392474
R3656 VDD.n764 VDD.n763 0.392399
R3657 VDD.n1346 VDD.n1345 0.392399
R3658 VDD.n1337 VDD.n1336 0.392399
R3659 VDD.n396 VDD.n395 0.392399
R3660 VDD.n544 VDD.n543 0.392399
R3661 VDD.n562 VDD.n269 0.392136
R3662 VDD.n1188 VDD 0.390595
R3663 VDD.n1101 VDD.n838 0.389939
R3664 VDD.n730 VDD 0.384624
R3665 VDD.n325 VDD 0.384624
R3666 VDD VDD.n748 0.382708
R3667 VDD.n181 VDD.n180 0.381006
R3668 VDD.n469 VDD.n468 0.381006
R3669 VDD.n1214 VDD.n1213 0.370786
R3670 VDD.n1204 VDD.n602 0.370786
R3671 VDD.n1297 VDD.n590 0.370786
R3672 VDD.n1311 VDD.n1310 0.370786
R3673 VDD.n1277 VDD.n1276 0.370786
R3674 VDD.n732 VDD.n731 0.370786
R3675 VDD.n739 VDD.n738 0.370786
R3676 VDD.n706 VDD.n705 0.370786
R3677 VDD.n720 VDD.n719 0.370786
R3678 VDD.n334 VDD.n333 0.370786
R3679 VDD.n327 VDD.n326 0.370786
R3680 VDD.n315 VDD.n314 0.370786
R3681 VDD.n305 VDD.n289 0.370786
R3682 VDD.n378 VDD.n377 0.370786
R3683 VDD.n364 VDD.n279 0.370786
R3684 VDD.n1318 VDD.n1317 0.370786
R3685 VDD.n580 VDD.n579 0.370786
R3686 VDD.n570 VDD.n258 0.370786
R3687 VDD.n1325 VDD.n1324 0.370786
R3688 VDD.n1283 VDD.n1282 0.370786
R3689 VDD.n1238 VDD.n1237 0.370786
R3690 VDD.n1231 VDD.n1230 0.370786
R3691 VDD.n241 VDD.n233 0.364413
R3692 VDD.n422 VDD.n414 0.364413
R3693 VDD.n1355 VDD.n1354 0.355908
R3694 VDD.n1368 VDD.n1367 0.355908
R3695 VDD.n537 VDD.n536 0.355908
R3696 VDD.n524 VDD.n523 0.355908
R3697 VDD VDD.n1199 0.355357
R3698 VDD.n1207 VDD 0.355357
R3699 VDD VDD.n1295 0.355357
R3700 VDD.n1303 VDD 0.355357
R3701 VDD VDD.n1273 0.355357
R3702 VDD VDD.n741 0.355357
R3703 VDD.n1178 VDD 0.355357
R3704 VDD VDD.n717 0.355357
R3705 VDD VDD.n336 0.355357
R3706 VDD VDD.n300 0.355357
R3707 VDD.n308 VDD 0.355357
R3708 VDD.n370 VDD 0.355357
R3709 VDD VDD.n362 0.355357
R3710 VDD VDD.n565 0.355357
R3711 VDD.n573 VDD 0.355357
R3712 VDD VDD.n1327 0.355357
R3713 VDD VDD.n1240 0.355357
R3714 VDD VDD.n1278 0.352009
R3715 VDD.n737 VDD 0.352009
R3716 VDD.n332 VDD 0.352009
R3717 VDD.n1323 VDD 0.352009
R3718 VDD.n1236 VDD 0.352009
R3719 VDD VDD.n1201 0.348937
R3720 VDD.n1301 VDD 0.348937
R3721 VDD.n607 VDD 0.348937
R3722 VDD VDD.n302 0.348937
R3723 VDD.n368 VDD 0.348937
R3724 VDD VDD.n567 0.348937
R3725 VDD.n893 VDD.n74 0.345864
R3726 VDD.n1673 VDD.n1672 0.338854
R3727 VDD.n893 VDD.n67 0.337206
R3728 VDD.n1404 VDD.n1403 0.337134
R3729 VDD.n200 VDD.n199 0.337134
R3730 VDD.n1385 VDD.n1384 0.337134
R3731 VDD.n217 VDD.n216 0.337134
R3732 VDD.n481 VDD.n480 0.337134
R3733 VDD.n490 VDD.n444 0.337134
R3734 VDD.n504 VDD.n503 0.337134
R3735 VDD.n513 VDD.n431 0.337134
R3736 VDD.n1410 VDD.n1409 0.335672
R3737 VDD.n194 VDD.n193 0.335672
R3738 VDD.n1391 VDD.n1390 0.335672
R3739 VDD.n211 VDD.n210 0.335672
R3740 VDD.n474 VDD.n473 0.335672
R3741 VDD.n482 VDD.n449 0.335672
R3742 VDD.n497 VDD.n496 0.335672
R3743 VDD.n505 VDD.n436 0.335672
R3744 VDD.n554 VDD.n553 0.327223
R3745 VDD.n277 VDD.n276 0.327223
R3746 VDD VDD.n23 0.326158
R3747 VDD VDD.n1 0.326158
R3748 VDD VDD.n13 0.326158
R3749 VDD.n192 VDD 0.3245
R3750 VDD VDD.n1392 0.3245
R3751 VDD.n209 VDD 0.3245
R3752 VDD VDD.n1373 0.3245
R3753 VDD VDD.n483 0.3245
R3754 VDD.n495 VDD 0.3245
R3755 VDD VDD.n506 0.3245
R3756 VDD.n518 VDD 0.3245
R3757 VDD.n1397 VDD.n1396 0.323688
R3758 VDD.n1386 VDD.n206 0.323688
R3759 VDD.n1378 VDD.n1377 0.323688
R3760 VDD.n491 VDD.n489 0.323688
R3761 VDD.n502 VDD.n441 0.323688
R3762 VDD.n514 VDD.n512 0.323688
R3763 VDD.n1405 VDD.n189 0.322018
R3764 VDD.n479 VDD.n454 0.322018
R3765 VDD.n188 VDD 0.321707
R3766 VDD VDD.n1398 0.321707
R3767 VDD VDD.n202 0.321707
R3768 VDD VDD.n1379 0.321707
R3769 VDD VDD.n475 0.321707
R3770 VDD.n488 VDD 0.321707
R3771 VDD VDD.n498 0.321707
R3772 VDD.n511 VDD 0.321707
R3773 VDD.n1666 VDD.n1665 0.31775
R3774 VDD.n1586 VDD.n1585 0.31775
R3775 VDD.n128 VDD.n98 0.31775
R3776 VDD.n1627 VDD.n60 0.31775
R3777 VDD.n895 VDD.n889 0.31775
R3778 VDD.n686 VDD.n681 0.31775
R3779 VDD.n1061 VDD.n1060 0.31775
R3780 VDD.n275 VDD 0.313609
R3781 VDD VDD.n548 0.31134
R3782 VDD VDD.n555 0.308434
R3783 VDD.n1180 VDD.n1179 0.306734
R3784 VDD.n975 VDD.n973 0.305717
R3785 VDD.n1534 VDD.n1532 0.305717
R3786 VDD.n86 VDD.n84 0.305717
R3787 VDD.n863 VDD.n861 0.305717
R3788 VDD.n1477 VDD.n1475 0.305717
R3789 VDD.n932 VDD.n930 0.305717
R3790 VDD.n641 VDD.n639 0.305717
R3791 VDD.n561 VDD.n560 0.30425
R3792 VDD.n284 VDD.n281 0.291221
R3793 VDD.n206 VDD.n157 0.290704
R3794 VDD.n210 VDD.n209 0.288115
R3795 VDD.n506 VDD.n505 0.288115
R3796 VDD.n1199 VDD.n1198 0.287841
R3797 VDD.n1295 VDD.n1294 0.287841
R3798 VDD.n717 VDD.n716 0.287841
R3799 VDD.n300 VDD.n299 0.287841
R3800 VDD.n362 VDD.n361 0.287841
R3801 VDD.n565 VDD.n564 0.287841
R3802 VDD.n1617 VDD.n67 0.283466
R3803 VDD.n1392 VDD.n1391 0.281855
R3804 VDD.n496 VDD.n495 0.281855
R3805 VDD.n1208 VDD.n1207 0.281308
R3806 VDD.n1304 VDD.n1303 0.281308
R3807 VDD.n1179 VDD.n1178 0.281308
R3808 VDD.n309 VDD.n308 0.281308
R3809 VDD.n371 VDD.n370 0.281308
R3810 VDD.n574 VDD.n573 0.281308
R3811 VDD.n356 VDD.n281 0.261539
R3812 VDD.n563 VDD.n268 0.248462
R3813 VDD.n1130 VDD.n1115 0.244844
R3814 VDD VDD.n1091 0.244297
R3815 VDD VDD.n1653 0.244297
R3816 VDD VDD.n1498 0.244297
R3817 VDD VDD.n878 0.244297
R3818 VDD VDD.n77 0.244297
R3819 VDD VDD.n1575 0.244297
R3820 VDD.n1578 VDD 0.244297
R3821 VDD.n1610 VDD 0.244297
R3822 VDD VDD.n1621 0.244297
R3823 VDD VDD.n1636 0.244297
R3824 VDD VDD.n1633 0.244297
R3825 VDD.n1465 VDD 0.244297
R3826 VDD.n881 VDD 0.244297
R3827 VDD.n1501 VDD 0.244297
R3828 VDD.n1273 VDD.n1272 0.243929
R3829 VDD.n741 VDD.n740 0.243929
R3830 VDD.n336 VDD.n335 0.243929
R3831 VDD.n1327 VDD.n1326 0.243929
R3832 VDD.n1240 VDD.n1239 0.243929
R3833 VDD.n1458 VDD.n156 0.240311
R3834 VDD.n564 VDD.n563 0.228271
R3835 VDD.n1683 VDD.n1682 0.217211
R3836 VDD.n1691 VDD.n5 0.217211
R3837 VDD.n1688 VDD.n1687 0.217211
R3838 VDD.n352 VDD.n351 0.211088
R3839 VDD.n1228 VDD 0.204624
R3840 VDD.n1289 VDD.n1288 0.202923
R3841 VDD.n1181 VDD.n1180 0.199201
R3842 VDD.n31 VDD 0.190753
R3843 VDD VDD.n785 0.1901
R3844 VDD.n1336 VDD.n1335 0.189761
R3845 VDD.n546 VDD.n544 0.189761
R3846 VDD.n287 VDD 0.18149
R3847 VDD.n1229 VDD.n1228 0.1805
R3848 VDD.n1167 VDD.n780 0.174566
R3849 VDD.n1679 VDD.n28 0.172525
R3850 VDD.n1666 VDD.n40 0.16925
R3851 VDD.n1659 VDD.n1657 0.16925
R3852 VDD.n1586 VDD.n1518 0.16925
R3853 VDD.n129 VDD.n128 0.16925
R3854 VDD.n113 VDD.n112 0.16925
R3855 VDD.n1641 VDD.n1640 0.16925
R3856 VDD.n1627 VDD.n1626 0.16925
R3857 VDD.n895 VDD.n894 0.16925
R3858 VDD.n874 VDD.n847 0.16925
R3859 VDD.n675 VDD.n674 0.16925
R3860 VDD.n686 VDD.n685 0.16925
R3861 VDD.n1097 VDD.n1095 0.16925
R3862 VDD.n1061 VDD.n1056 0.16925
R3863 VDD.n1264 VDD.n595 0.16925
R3864 VDD.n1266 VDD.n1264 0.168529
R3865 VDD.n992 VDD.n989 0.168444
R3866 VDD.n1024 VDD.n1023 0.168444
R3867 VDD.n915 VDD.n914 0.168444
R3868 VDD.n620 VDD.n619 0.168444
R3869 VDD.n354 VDD.n353 0.167
R3870 VDD.n276 VDD.n275 0.166887
R3871 VDD.n844 VDD.n842 0.164678
R3872 VDD.n1565 VDD.n1564 0.163625
R3873 VDD.n1490 VDD.n1488 0.163625
R3874 VDD.n1568 VDD.n1566 0.1625
R3875 VDD.n1663 VDD.n46 0.1577
R3876 VDD.n1042 VDD.n1041 0.1577
R3877 VDD.n1583 VDD.n1524 0.1577
R3878 VDD.n1581 VDD.n1580 0.1577
R3879 VDD.n1602 VDD.n1601 0.1577
R3880 VDD.n125 VDD.n124 0.1577
R3881 VDD.n1012 VDD.n1011 0.1577
R3882 VDD.n1614 VDD.n1612 0.1577
R3883 VDD.n1469 VDD.n1467 0.1577
R3884 VDD.n1631 VDD.n1630 0.1577
R3885 VDD.n903 VDD.n902 0.1577
R3886 VDD.n884 VDD.n883 0.1577
R3887 VDD.n149 VDD.n148 0.1577
R3888 VDD.n1504 VDD.n1503 0.1577
R3889 VDD.n1670 VDD.n36 0.1577
R3890 VDD.n1082 VDD.n1081 0.1577
R3891 VDD.n691 VDD.n690 0.1577
R3892 VDD.n679 VDD.n657 0.1577
R3893 VDD.n1175 VDD.n635 0.1577
R3894 VDD.n1085 VDD.n1084 0.1577
R3895 VDD.n964 VDD.n963 0.1577
R3896 VDD.n1260 VDD.n1259 0.1577
R3897 VDD.n976 VDD.n975 0.157022
R3898 VDD.n1535 VDD.n1534 0.157022
R3899 VDD.n87 VDD.n86 0.157022
R3900 VDD.n864 VDD.n863 0.157022
R3901 VDD.n1478 VDD.n1477 0.157022
R3902 VDD.n1065 VDD.n932 0.157022
R3903 VDD.n1173 VDD.n641 0.157022
R3904 VDD.n1348 VDD.n1346 0.149943
R3905 VDD.n395 VDD.n386 0.149943
R3906 VDD.n349 VDD.n345 0.143192
R3907 VDD.n763 VDD 0.133791
R3908 VDD.n1345 VDD 0.133791
R3909 VDD VDD.n1337 0.133791
R3910 VDD VDD.n396 0.133791
R3911 VDD.n543 VDD 0.133791
R3912 VDD.n355 VDD.n354 0.128
R3913 VDD.n287 VDD.n269 0.126502
R3914 VDD.n765 VDD.n764 0.125816
R3915 VDD.n1352 VDD 0.101892
R3916 VDD.n1349 VDD 0.101892
R3917 VDD.n539 VDD 0.101892
R3918 VDD VDD.n542 0.101892
R3919 VDD.n1131 VDD.n1130 0.100143
R3920 VDD.n1131 VDD.n1113 0.0985357
R3921 VDD.n620 VDD.n610 0.093875
R3922 VDD.n1589 VDD.n134 0.0935509
R3923 VDD.n1508 VDD.n1459 0.0897373
R3924 VDD VDD.n893 0.087125
R3925 VDD VDD.n1404 0.0843983
R3926 VDD.n199 VDD 0.0843983
R3927 VDD VDD.n1385 0.0843983
R3928 VDD.n216 VDD 0.0843983
R3929 VDD.n480 VDD 0.0843983
R3930 VDD VDD.n490 0.0843983
R3931 VDD.n503 VDD 0.0843983
R3932 VDD VDD.n513 0.0843983
R3933 VDD.n1686 VDD 0.07475
R3934 VDD.n1488 VDD 0.06125
R3935 VDD.n1565 VDD.n1562 0.060125
R3936 VDD VDD.n40 0.055625
R3937 VDD.n1657 VDD 0.055625
R3938 VDD.n1518 VDD 0.055625
R3939 VDD.n1558 VDD 0.055625
R3940 VDD VDD.n129 0.055625
R3941 VDD VDD.n113 0.055625
R3942 VDD.n1640 VDD 0.055625
R3943 VDD.n1626 VDD 0.055625
R3944 VDD.n894 VDD 0.055625
R3945 VDD VDD.n874 0.055625
R3946 VDD.n674 VDD 0.055625
R3947 VDD.n685 VDD 0.055625
R3948 VDD.n1095 VDD 0.055625
R3949 VDD.n1056 VDD 0.055625
R3950 VDD VDD.n595 0.055625
R3951 VDD.n989 VDD 0.0549444
R3952 VDD.n1023 VDD 0.0549444
R3953 VDD.n914 VDD 0.0549444
R3954 VDD.n619 VDD 0.0549444
R3955 VDD.n834 VDD.n822 0.053063
R3956 VDD.n1109 VDD.n823 0.053063
R3957 VDD.n173 VDD.n172 0.053063
R3958 VDD.n1435 VDD.n1434 0.053063
R3959 VDD.n790 VDD.n789 0.053063
R3960 VDD.n1133 VDD.n1132 0.053063
R3961 VDD.n807 VDD.n795 0.053063
R3962 VDD.n816 VDD.n796 0.053063
R3963 VDD.n1445 VDD.n161 0.053063
R3964 VDD.n1453 VDD.n160 0.053063
R3965 VDD.n1150 VDD.n1139 0.053063
R3966 VDD.n1159 VDD.n1140 0.053063
R3967 VDD.n830 VDD.n821 0.0526849
R3968 VDD.n1110 VDD.n820 0.0526849
R3969 VDD.n1421 VDD.n1418 0.0526849
R3970 VDD.n1430 VDD.n171 0.0526849
R3971 VDD.n1121 VDD.n1120 0.0526849
R3972 VDD.n788 VDD.n786 0.0526849
R3973 VDD.n803 VDD.n794 0.0526849
R3974 VDD.n817 VDD.n793 0.0526849
R3975 VDD.n1444 VDD.n166 0.0526849
R3976 VDD.n1443 VDD.n167 0.0526849
R3977 VDD.n1146 VDD.n1138 0.0526849
R3978 VDD.n1160 VDD.n1137 0.0526849
R3979 VDD.n992 VDD.n991 0.0513605
R3980 VDD.n835 VDD.n833 0.050741
R3981 VDD.n1424 VDD.n1423 0.050741
R3982 VDD.n1124 VDD.n1123 0.050741
R3983 VDD.n808 VDD.n806 0.050741
R3984 VDD.n1447 VDD.n1446 0.050741
R3985 VDD.n1151 VDD.n1149 0.050741
R3986 VDD.n1112 VDD.n1111 0.0506887
R3987 VDD.n828 VDD.n827 0.0470126
R3988 VDD.n1106 VDD.n1105 0.0470126
R3989 VDD.n1425 VDD.n1420 0.0470126
R3990 VDD.n1419 VDD.n174 0.0470126
R3991 VDD.n1125 VDD.n1116 0.0470126
R3992 VDD.n1129 VDD.n791 0.0470126
R3993 VDD.n801 VDD.n800 0.0470126
R3994 VDD.n813 VDD.n812 0.0470126
R3995 VDD.n164 VDD.n162 0.0470126
R3996 VDD.n1452 VDD.n163 0.0470126
R3997 VDD.n1144 VDD.n1143 0.0470126
R3998 VDD.n1156 VDD.n1155 0.0470126
R3999 VDD.n842 VDD 0.0469211
R4000 VDD.n586 VDD.n266 0.0420385
R4001 VDD.n1288 VDD.n1268 0.0420385
R4002 VDD.n1248 VDD 0.041
R4003 VDD.n1353 VDD 0.0390714
R4004 VDD.n538 VDD 0.0390714
R4005 VDD.n1414 VDD.n1413 0.0349922
R4006 VDD.n248 VDD.n247 0.0322647
R4007 VDD.n402 VDD.n401 0.0322647
R4008 VDD.n1577 VDD.n1572 0.0310814
R4009 VDD.n1500 VDD.n1495 0.0310814
R4010 VDD.n353 VDD.n283 0.0305
R4011 VDD.n1115 VDD.n1114 0.0302656
R4012 VDD.n1656 VDD.n1655 0.0301203
R4013 VDD.n1557 VDD.n1556 0.0301203
R4014 VDD.n1597 VDD.n130 0.0301203
R4015 VDD.n120 VDD.n114 0.0301203
R4016 VDD.n1609 VDD.n74 0.0301203
R4017 VDD.n1639 VDD.n1638 0.0301203
R4018 VDD.n1625 VDD.n1624 0.0301203
R4019 VDD.n880 VDD.n875 0.0301203
R4020 VDD.n1517 VDD.n1516 0.0301203
R4021 VDD.n1673 VDD.n31 0.0301203
R4022 VDD.n947 VDD.n946 0.0301203
R4023 VDD.n673 VDD.n672 0.0301203
R4024 VDD.n695 VDD.n645 0.0301203
R4025 VDD.n1094 VDD.n1093 0.0301203
R4026 VDD.n1055 VDD.n1054 0.0301203
R4027 VDD.n1255 VDD.n1249 0.0301203
R4028 VDD.n1114 VDD.n787 0.0297969
R4029 VDD.n1037 VDD.n1031 0.0295001
R4030 VDD.n1077 VDD.n838 0.0295001
R4031 VDD.n631 VDD.n625 0.0285654
R4032 VDD.n1022 VDD.n1021 0.0285499
R4033 VDD.n913 VDD.n912 0.0285499
R4034 VDD.n1442 VDD.n1441 0.0265377
R4035 VDD.n1316 VDD.n586 0.0251429
R4036 VDD.n1288 VDD.n1287 0.0251429
R4037 VDD.n250 VDD.n248 0.0216225
R4038 VDD.n1372 VDD 0.0216225
R4039 VDD.n403 VDD.n402 0.0216225
R4040 VDD VDD.n519 0.0216225
R4041 VDD.n1451 VDD.n159 0.0212547
R4042 VDD.n815 VDD.n798 0.0208774
R4043 VDD.n1108 VDD.n825 0.0208774
R4044 VDD.n1218 VDD.n1197 0.0203701
R4045 VDD.n1210 VDD.n1209 0.0203701
R4046 VDD.n1293 VDD.n1292 0.0203701
R4047 VDD.n1306 VDD.n1305 0.0203701
R4048 VDD.n1313 VDD.n588 0.0203701
R4049 VDD.n745 VDD.n708 0.0203701
R4050 VDD.n759 VDD.n758 0.0203701
R4051 VDD.n1182 VDD.n1181 0.0203701
R4052 VDD.n724 VDD.n715 0.0203701
R4053 VDD.n340 VDD.n291 0.0203701
R4054 VDD.n319 VDD.n298 0.0203701
R4055 VDD.n311 VDD.n310 0.0203701
R4056 VDD.n463 VDD.n461 0.0203701
R4057 VDD.n373 VDD.n372 0.0203701
R4058 VDD.n360 VDD.n359 0.0203701
R4059 VDD.n584 VDD.n268 0.0203701
R4060 VDD.n576 VDD.n575 0.0203701
R4061 VDD.n1331 VDD.n260 0.0203701
R4062 VDD.n1244 VDD.n1190 0.0203701
R4063 VDD.n729 VDD.n727 0.0162732
R4064 VDD.n324 VDD.n322 0.0162732
R4065 VDD.n1223 VDD.n1221 0.0162732
R4066 VDD.n1455 VDD.n158 0.0161604
R4067 VDD.n1117 VDD.n787 0.0149643
R4068 VDD.n1279 VDD.n1270 0.014934
R4069 VDD.n736 VDD.n711 0.014934
R4070 VDD.n331 VDD.n294 0.014934
R4071 VDD.n1322 VDD.n263 0.014934
R4072 VDD.n1235 VDD.n1193 0.014934
R4073 VDD.n1437 VDD.n1436 0.0144623
R4074 VDD.n1403 VDD.n1402 0.0138043
R4075 VDD.n1393 VDD.n200 0.0138043
R4076 VDD.n1384 VDD.n1383 0.0138043
R4077 VDD.n1374 VDD.n217 0.0138043
R4078 VDD.n484 VDD.n481 0.0138043
R4079 VDD.n494 VDD.n444 0.0138043
R4080 VDD.n507 VDD.n504 0.0138043
R4081 VDD.n517 VDD.n431 0.0138043
R4082 VDD.n1409 VDD.n1408 0.0136897
R4083 VDD.n1399 VDD.n194 0.0136897
R4084 VDD.n1390 VDD.n1389 0.0136897
R4085 VDD.n1380 VDD.n211 0.0136897
R4086 VDD.n476 VDD.n474 0.0136897
R4087 VDD.n487 VDD.n449 0.0136897
R4088 VDD.n499 VDD.n497 0.0136897
R4089 VDD.n510 VDD.n436 0.0136897
R4090 VDD.n549 VDD.n277 0.0133571
R4091 VDD.n286 VDD.n283 0.01325
R4092 VDD.n556 VDD.n272 0.0131446
R4093 VDD.n1142 VDD.n1141 0.0125755
R4094 VDD VDD.n1214 0.0125
R4095 VDD VDD.n1204 0.0125
R4096 VDD VDD.n1297 0.0125
R4097 VDD.n1310 VDD 0.0125
R4098 VDD.n1276 VDD 0.0125
R4099 VDD VDD.n732 0.0125
R4100 VDD VDD.n739 0.0125
R4101 VDD.n705 VDD 0.0125
R4102 VDD VDD.n720 0.0125
R4103 VDD VDD.n334 0.0125
R4104 VDD VDD.n327 0.0125
R4105 VDD VDD.n315 0.0125
R4106 VDD VDD.n305 0.0125
R4107 VDD.n377 VDD 0.0125
R4108 VDD VDD.n364 0.0125
R4109 VDD VDD.n1318 0.0125
R4110 VDD VDD.n580 0.0125
R4111 VDD VDD.n570 0.0125
R4112 VDD VDD.n1325 0.0125
R4113 VDD VDD.n1283 0.0125
R4114 VDD VDD.n1238 0.0125
R4115 VDD VDD.n1231 0.0125
R4116 VDD.n553 VDD 0.0110882
R4117 VDD.n560 VDD 0.0103438
R4118 VDD.n1158 VDD.n1142 0.00936793
R4119 VDD.n756 VDD.n754 0.00878947
R4120 VDD.n1344 VDD.n1342 0.00878947
R4121 VDD.n257 VDD.n255 0.00878947
R4122 VDD.n393 VDD.n391 0.00878947
R4123 VDD.n385 VDD.n383 0.00878947
R4124 VDD.n1566 VDD.n1558 0.00725
R4125 VDD.n1437 VDD.n169 0.00691509
R4126 VDD.n1101 VDD 0.00569231
R4127 VDD.n1455 VDD.n1454 0.00427358
R4128 VDD.n1134 VDD.n787 0.00401562
R4129 VDD.n1680 VDD.n1679 0.00391772
R4130 VDD.n1142 VDD.n168 0.00379268
R4131 VDD.n1215 VDD 0.00307143
R4132 VDD.n1206 VDD 0.00307143
R4133 VDD.n1298 VDD 0.00307143
R4134 VDD VDD.n1309 0.00307143
R4135 VDD VDD.n1275 0.00307143
R4136 VDD.n733 VDD 0.00307143
R4137 VDD.n742 VDD 0.00307143
R4138 VDD.n1177 VDD 0.00307143
R4139 VDD.n721 VDD 0.00307143
R4140 VDD.n337 VDD 0.00307143
R4141 VDD.n328 VDD 0.00307143
R4142 VDD.n316 VDD 0.00307143
R4143 VDD.n307 VDD 0.00307143
R4144 VDD VDD.n376 0.00307143
R4145 VDD.n365 VDD 0.00307143
R4146 VDD.n1319 VDD 0.00307143
R4147 VDD.n581 VDD 0.00307143
R4148 VDD.n572 VDD 0.00307143
R4149 VDD.n1328 VDD 0.00307143
R4150 VDD.n1284 VDD 0.00307143
R4151 VDD.n1241 VDD 0.00307143
R4152 VDD.n1232 VDD 0.00307143
R4153 VDD.n1683 VDD 0.00286842
R4154 VDD VDD.n1691 0.00286842
R4155 VDD.n1688 VDD 0.00286842
R4156 VDD.n829 VDD.n820 0.00276891
R4157 VDD.n1431 VDD.n1430 0.00276891
R4158 VDD.n1118 VDD.n786 0.00276891
R4159 VDD.n802 VDD.n793 0.00276891
R4160 VDD.n1439 VDD.n167 0.00276891
R4161 VDD.n1145 VDD.n1137 0.00276891
R4162 VDD VDD.n552 0.00276891
R4163 VDD VDD.n559 0.00260938
R4164 VDD.n939 VDD 0.00259302
R4165 VDD.n1650 VDD 0.00259302
R4166 VDD.n1513 VDD 0.00259302
R4167 VDD.n1019 VDD 0.00259302
R4168 VDD.n1035 VDD 0.00259302
R4169 VDD VDD.n1038 0.00259302
R4170 VDD.n1051 VDD 0.00259302
R4171 VDD.n118 VDD 0.00259302
R4172 VDD.n1594 VDD 0.00259302
R4173 VDD.n1554 VDD 0.00259302
R4174 VDD.n1550 VDD 0.00259302
R4175 VDD VDD.n1598 0.00259302
R4176 VDD VDD.n121 0.00259302
R4177 VDD.n1015 VDD 0.00259302
R4178 VDD.n910 VDD 0.00259302
R4179 VDD.n906 VDD 0.00259302
R4180 VDD.n152 VDD 0.00259302
R4181 VDD.n945 VDD 0.00259302
R4182 VDD.n1075 VDD 0.00259302
R4183 VDD VDD.n1078 0.00259302
R4184 VDD.n629 VDD 0.00259302
R4185 VDD.n699 VDD 0.00259302
R4186 VDD.n670 VDD 0.00259302
R4187 VDD.n694 VDD 0.00259302
R4188 VDD.n666 VDD 0.00259302
R4189 VDD VDD.n632 0.00259302
R4190 VDD.n1088 VDD 0.00259302
R4191 VDD.n967 VDD 0.00259302
R4192 VDD.n179 VDD 0.00259302
R4193 VDD VDD.n1412 0.00259302
R4194 VDD.n467 VDD 0.00259302
R4195 VDD.n471 VDD 0.00259302
R4196 VDD.n1253 VDD 0.00259302
R4197 VDD VDD.n1256 0.00259302
R4198 VDD.n1135 VDD.n1134 0.00214062
R4199 VDD.n831 VDD.n830 0.00213389
R4200 VDD.n1418 VDD.n1417 0.00213389
R4201 VDD.n1120 VDD.n1119 0.00213389
R4202 VDD.n804 VDD.n803 0.00213389
R4203 VDD.n1438 VDD.n166 0.00213389
R4204 VDD.n1147 VDD.n1146 0.00213389
R4205 VDD.n1113 VDD.n787 0.00210714
R4206 VDD VDD.n1046 0.00202542
R4207 VDD VDD.n1589 0.00202542
R4208 VDD VDD.n1606 0.00202542
R4209 VDD VDD.n1617 0.00202542
R4210 VDD VDD.n1508 0.00202542
R4211 VDD.n1064 VDD 0.00202542
R4212 VDD.n1172 VDD 0.00202542
R4213 VDD.n1105 VDD.n1104 0.00201261
R4214 VDD.n1428 VDD.n1419 0.00201261
R4215 VDD.n1129 VDD.n1128 0.00201261
R4216 VDD.n812 VDD.n811 0.00201261
R4217 VDD.n1450 VDD.n163 0.00201261
R4218 VDD.n1155 VDD.n1154 0.00201261
R4219 VDD.n837 VDD.n828 0.00175605
R4220 VDD.n1427 VDD.n1420 0.00175605
R4221 VDD.n1127 VDD.n1116 0.00175605
R4222 VDD.n810 VDD.n801 0.00175605
R4223 VDD.n1449 VDD.n164 0.00175605
R4224 VDD.n1153 VDD.n1144 0.00175605
R4225 VDD.n771 VDD 0.00175
R4226 VDD VDD.n1663 0.0017
R4227 VDD.n1042 VDD 0.0017
R4228 VDD VDD.n1583 0.0017
R4229 VDD.n1581 VDD 0.0017
R4230 VDD.n1602 VDD 0.0017
R4231 VDD.n125 VDD 0.0017
R4232 VDD.n1011 VDD 0.0017
R4233 VDD.n1614 VDD 0.0017
R4234 VDD.n1469 VDD 0.0017
R4235 VDD.n1630 VDD 0.0017
R4236 VDD.n902 VDD 0.0017
R4237 VDD VDD.n884 0.0017
R4238 VDD.n148 VDD 0.0017
R4239 VDD.n1504 VDD 0.0017
R4240 VDD VDD.n1670 0.0017
R4241 VDD.n1082 VDD 0.0017
R4242 VDD VDD.n1187 0.0017
R4243 VDD.n690 VDD 0.0017
R4244 VDD VDD.n679 0.0017
R4245 VDD.n1175 VDD 0.0017
R4246 VDD.n1084 VDD 0.0017
R4247 VDD.n963 VDD 0.0017
R4248 VDD.n345 VDD 0.0017
R4249 VDD.n1260 VDD 0.0017
R4250 VDD VDD.n1218 0.00166883
R4251 VDD.n1210 VDD 0.00166883
R4252 VDD.n1292 VDD 0.00166883
R4253 VDD.n1306 VDD 0.00166883
R4254 VDD.n1313 VDD 0.00166883
R4255 VDD VDD.n745 0.00166883
R4256 VDD.n759 VDD 0.00166883
R4257 VDD.n1182 VDD 0.00166883
R4258 VDD VDD.n724 0.00166883
R4259 VDD VDD.n340 0.00166883
R4260 VDD VDD.n319 0.00166883
R4261 VDD.n311 VDD 0.00166883
R4262 VDD VDD.n463 0.00166883
R4263 VDD.n373 VDD 0.00166883
R4264 VDD.n359 VDD 0.00166883
R4265 VDD VDD.n584 0.00166883
R4266 VDD.n576 VDD 0.00166883
R4267 VDD VDD.n1331 0.00166883
R4268 VDD VDD.n1244 0.00166883
R4269 VDD VDD.n1167 0.00165385
R4270 VDD VDD.n28 0.00163924
R4271 VDD.n822 VDD.n821 0.00163445
R4272 VDD.n1110 VDD.n1109 0.00163445
R4273 VDD.n1421 VDD.n172 0.00163445
R4274 VDD.n1435 VDD.n171 0.00163445
R4275 VDD.n1121 VDD.n789 0.00163445
R4276 VDD.n1133 VDD.n788 0.00163445
R4277 VDD.n795 VDD.n794 0.00163445
R4278 VDD.n817 VDD.n816 0.00163445
R4279 VDD.n1445 VDD.n1444 0.00163445
R4280 VDD.n1443 VDD.n160 0.00163445
R4281 VDD.n1139 VDD.n1138 0.00163445
R4282 VDD.n1160 VDD.n1159 0.00163445
R4283 VDD.n1441 VDD.n1440 0.00163208
R4284 VDD.n1562 VDD 0.001625
R4285 VDD.n352 VDD.n284 0.00159756
R4286 VDD.n833 VDD.n832 0.00158434
R4287 VDD.n1423 VDD.n1422 0.00158434
R4288 VDD.n1123 VDD.n1122 0.00158434
R4289 VDD.n806 VDD.n805 0.00158434
R4290 VDD.n1446 VDD.n165 0.00158434
R4291 VDD.n1149 VDD.n1148 0.00158434
R4292 VDD VDD.n1316 0.00157143
R4293 VDD.n1287 VDD 0.00157143
R4294 VDD VDD.n729 0.00142783
R4295 VDD VDD.n324 0.00142783
R4296 VDD VDD.n1223 0.00142783
R4297 VDD VDD.n250 0.00141837
R4298 VDD.n1355 VDD 0.00141837
R4299 VDD VDD.n1358 0.00141837
R4300 VDD.n1359 VDD 0.00141837
R4301 VDD VDD.n1362 0.00141837
R4302 VDD.n1363 VDD 0.00141837
R4303 VDD VDD.n1366 0.00141837
R4304 VDD.n1368 VDD 0.00141837
R4305 VDD VDD.n1371 0.00141837
R4306 VDD.n403 VDD 0.00141837
R4307 VDD.n536 VDD 0.00141837
R4308 VDD.n533 VDD 0.00141837
R4309 VDD.n532 VDD 0.00141837
R4310 VDD.n529 VDD 0.00141837
R4311 VDD.n528 VDD 0.00141837
R4312 VDD.n525 VDD 0.00141837
R4313 VDD.n523 VDD 0.00141837
R4314 VDD.n520 VDD 0.00141837
R4315 VDD.n1215 VDD 0.00135714
R4316 VDD VDD.n1206 0.00135714
R4317 VDD.n1298 VDD 0.00135714
R4318 VDD.n1309 VDD 0.00135714
R4319 VDD.n1275 VDD 0.00135714
R4320 VDD.n733 VDD 0.00135714
R4321 VDD.n742 VDD 0.00135714
R4322 VDD VDD.n1177 0.00135714
R4323 VDD.n721 VDD 0.00135714
R4324 VDD.n337 VDD 0.00135714
R4325 VDD.n328 VDD 0.00135714
R4326 VDD.n316 VDD 0.00135714
R4327 VDD VDD.n307 0.00135714
R4328 VDD.n376 VDD 0.00135714
R4329 VDD.n365 VDD 0.00135714
R4330 VDD.n1319 VDD 0.00135714
R4331 VDD.n581 VDD 0.00135714
R4332 VDD VDD.n572 0.00135714
R4333 VDD.n1328 VDD 0.00135714
R4334 VDD.n1284 VDD 0.00135714
R4335 VDD.n1241 VDD 0.00135714
R4336 VDD.n1232 VDD 0.00135714
R4337 VDD.n1279 VDD 0.00134906
R4338 VDD VDD.n736 0.00134906
R4339 VDD VDD.n331 0.00134906
R4340 VDD VDD.n1322 0.00134906
R4341 VDD VDD.n1235 0.00134906
R4342 VDD.n1402 VDD 0.00128261
R4343 VDD.n1393 VDD 0.00128261
R4344 VDD.n1383 VDD 0.00128261
R4345 VDD.n1374 VDD 0.00128261
R4346 VDD.n484 VDD 0.00128261
R4347 VDD VDD.n494 0.00128261
R4348 VDD.n507 VDD 0.00128261
R4349 VDD VDD.n517 0.00128261
R4350 VDD.n1408 VDD 0.00127586
R4351 VDD.n1399 VDD 0.00127586
R4352 VDD.n1389 VDD 0.00127586
R4353 VDD.n1380 VDD 0.00127586
R4354 VDD.n476 VDD 0.00127586
R4355 VDD VDD.n487 0.00127586
R4356 VDD.n499 VDD 0.00127586
R4357 VDD VDD.n510 0.00127586
R4358 VDD.n1405 VDD 0.00126271
R4359 VDD.n1396 VDD 0.00126271
R4360 VDD.n1386 VDD 0.00126271
R4361 VDD.n1377 VDD 0.00126271
R4362 VDD VDD.n479 0.00126271
R4363 VDD.n491 VDD 0.00126271
R4364 VDD VDD.n502 0.00126271
R4365 VDD.n514 VDD 0.00126271
R4366 VDD.n552 VDD 0.0012563
R4367 VDD.n549 VDD 0.0012563
R4368 VDD.n797 VDD.n792 0.00125472
R4369 VDD.n1141 VDD.n1136 0.00125472
R4370 VDD.n824 VDD.n819 0.00125472
R4371 VDD.n1433 VDD.n1432 0.00125472
R4372 VDD VDD.n286 0.00125
R4373 VDD.n556 VDD 0.0012438
R4374 VDD.n559 VDD 0.00120312
R4375 VDD.n1442 VDD.n158 0.00106604
R4376 VDD.n798 VDD.n797 0.00106604
R4377 VDD.n799 VDD.n156 0.00106604
R4378 VDD.n1454 VDD.n159 0.00106604
R4379 VDD.n825 VDD.n824 0.00106604
R4380 VDD.n1103 VDD.n826 0.00106604
R4381 VDD.n1433 VDD.n169 0.00106604
R4382 VDD.n834 VDD.n827 0.000878151
R4383 VDD.n1106 VDD.n823 0.000878151
R4384 VDD.n1425 VDD.n173 0.000878151
R4385 VDD.n1434 VDD.n174 0.000878151
R4386 VDD.n1125 VDD.n790 0.000878151
R4387 VDD.n1132 VDD.n791 0.000878151
R4388 VDD.n807 VDD.n800 0.000878151
R4389 VDD.n813 VDD.n796 0.000878151
R4390 VDD.n162 VDD.n161 0.000878151
R4391 VDD.n1453 VDD.n1452 0.000878151
R4392 VDD.n1150 VDD.n1143 0.000878151
R4393 VDD.n1156 VDD.n1140 0.000878151
R4394 VDD.n818 VDD.n792 0.000877358
R4395 VDD.n815 VDD.n814 0.000877358
R4396 VDD.n814 VDD.n799 0.000877358
R4397 VDD.n1161 VDD.n1136 0.000877358
R4398 VDD.n1158 VDD.n1157 0.000877358
R4399 VDD.n1111 VDD.n819 0.000877358
R4400 VDD.n1108 VDD.n1107 0.000877358
R4401 VDD.n1107 VDD.n826 0.000877358
R4402 VDD.n1432 VDD.n1416 0.000877358
R4403 VDD.n1436 VDD.n170 0.000877358
R4404 VDD.n1429 VDD.n170 0.000877358
R4405 VDD.n836 VDD.n835 0.000861446
R4406 VDD.n1426 VDD.n1424 0.000861446
R4407 VDD.n1126 VDD.n1124 0.000861446
R4408 VDD.n809 VDD.n808 0.000861446
R4409 VDD.n1448 VDD.n1447 0.000861446
R4410 VDD.n1152 VDD.n1151 0.000861446
R4411 CLK.n29 CLK.t108 52.9255
R4412 CLK.n36 CLK.t50 52.9255
R4413 CLK.t40 CLK.t9 47.8944
R4414 CLK.t28 CLK.t119 47.8944
R4415 CLK.t78 CLK.t126 47.8944
R4416 CLK.t13 CLK.t66 47.8944
R4417 CLK.t70 CLK.t107 47.8944
R4418 CLK.t8 CLK.t114 47.8944
R4419 CLK.t99 CLK.t22 47.8944
R4420 CLK.t27 CLK.t6 47.8944
R4421 CLK.t35 CLK.t23 47.8944
R4422 CLK.t87 CLK.t2 47.8944
R4423 CLK.t10 CLK.t74 47.8944
R4424 CLK.t24 CLK.t97 47.8944
R4425 CLK.n15 CLK.t59 47.3388
R4426 CLK.n53 CLK.t60 47.3388
R4427 CLK.n4 CLK.t17 47.3388
R4428 CLK.n73 CLK.t55 47.2524
R4429 CLK.n33 CLK.t116 38.8649
R4430 CLK.n31 CLK.t117 38.8649
R4431 CLK.n39 CLK.t30 38.8649
R4432 CLK.n42 CLK.t42 38.8649
R4433 CLK.n26 CLK.t39 38.8649
R4434 CLK.n6 CLK.t54 38.8649
R4435 CLK.n9 CLK.t90 38.7949
R4436 CLK.n8 CLK.t43 38.7949
R4437 CLK.n13 CLK.t3 38.7949
R4438 CLK.n12 CLK.t36 38.7949
R4439 CLK.n18 CLK.t29 38.7949
R4440 CLK.n19 CLK.t115 38.7949
R4441 CLK.n55 CLK.t58 38.7949
R4442 CLK.n56 CLK.t53 38.7949
R4443 CLK.n51 CLK.t51 38.7949
R4444 CLK.n50 CLK.t89 38.7949
R4445 CLK.n62 CLK.t77 38.7949
R4446 CLK.n61 CLK.t34 38.7949
R4447 CLK.n67 CLK.t81 38.7949
R4448 CLK.n66 CLK.t67 38.7949
R4449 CLK.n79 CLK.t12 38.7949
R4450 CLK.n78 CLK.t16 38.7949
R4451 CLK.n75 CLK.t113 38.7949
R4452 CLK.n74 CLK.t122 38.7949
R4453 CLK.n70 CLK.t25 38.7949
R4454 CLK.n71 CLK.t120 38.7949
R4455 CLK.n87 CLK.t65 38.7949
R4456 CLK.n88 CLK.t109 38.7949
R4457 CLK.n2 CLK.t101 38.7949
R4458 CLK.n1 CLK.t11 38.7949
R4459 CLK.n9 CLK.n8 31.4949
R4460 CLK.n13 CLK.n12 31.4949
R4461 CLK.n19 CLK.n18 31.4949
R4462 CLK.n56 CLK.n55 31.4949
R4463 CLK.n51 CLK.n50 31.4949
R4464 CLK.n62 CLK.n61 31.4949
R4465 CLK.n67 CLK.n66 31.4949
R4466 CLK.n79 CLK.n78 31.4949
R4467 CLK.n75 CLK.n74 31.4949
R4468 CLK.n71 CLK.n70 31.4949
R4469 CLK.n88 CLK.n87 31.4949
R4470 CLK.n2 CLK.n1 31.4949
R4471 CLK.n21 CLK.t93 31.3561
R4472 CLK.n58 CLK.t18 31.3561
R4473 CLK.n90 CLK.t15 31.3561
R4474 CLK.n81 CLK.t19 31.3542
R4475 CLK.n28 CLK.t112 28.8568
R4476 CLK.n35 CLK.t61 28.8568
R4477 CLK.n32 CLK.t125 28.8568
R4478 CLK.n30 CLK.t63 28.8568
R4479 CLK.n38 CLK.t92 28.8568
R4480 CLK.n41 CLK.t94 28.8568
R4481 CLK.n25 CLK.t45 28.8568
R4482 CLK.n5 CLK.t118 28.8568
R4483 CLK.n11 CLK.t62 26.9781
R4484 CLK.n11 CLK.t111 26.9781
R4485 CLK.n17 CLK.t103 26.9781
R4486 CLK.n17 CLK.t48 26.9781
R4487 CLK.n54 CLK.t72 26.9781
R4488 CLK.n54 CLK.t88 26.9781
R4489 CLK.n49 CLK.t95 26.9781
R4490 CLK.n49 CLK.t4 26.9781
R4491 CLK.n77 CLK.t75 26.9781
R4492 CLK.n77 CLK.t20 26.9781
R4493 CLK.n69 CLK.t79 26.9781
R4494 CLK.n69 CLK.t31 26.9781
R4495 CLK.n86 CLK.t91 26.9781
R4496 CLK.n86 CLK.t1 26.9781
R4497 CLK.n0 CLK.t71 26.9781
R4498 CLK.n0 CLK.t83 26.9781
R4499 CLK.n83 CLK 19.7538
R4500 CLK.n44 CLK.n43 19.2225
R4501 CLK.n10 CLK.t127 17.9416
R4502 CLK.n14 CLK.t121 17.9416
R4503 CLK.n20 CLK.t123 17.9416
R4504 CLK.n57 CLK.t100 17.9416
R4505 CLK.n52 CLK.t14 17.9416
R4506 CLK.n63 CLK.t38 17.9416
R4507 CLK.n68 CLK.t41 17.9416
R4508 CLK.n80 CLK.t68 17.9416
R4509 CLK.n72 CLK.t52 17.9416
R4510 CLK.n89 CLK.t96 17.9416
R4511 CLK.n3 CLK.t56 17.9416
R4512 CLK.n76 CLK.t86 17.6937
R4513 CLK.n45 CLK.n44 17.1932
R4514 CLK.t108 CLK.n28 17.0773
R4515 CLK.t50 CLK.n35 17.0773
R4516 CLK.t116 CLK.n32 17.0773
R4517 CLK.t117 CLK.n30 17.0773
R4518 CLK.t30 CLK.n38 17.0773
R4519 CLK.t42 CLK.n41 17.0773
R4520 CLK.t39 CLK.n25 17.0773
R4521 CLK.t54 CLK.n5 17.0773
R4522 CLK.n65 CLK.n64 15.7794
R4523 CLK.n48 CLK 15.7041
R4524 CLK.n84 CLK.n83 14.5859
R4525 CLK.n24 CLK.n23 14.0672
R4526 CLK.n60 CLK.n59 12.5623
R4527 CLK.n92 CLK.n91 12.5623
R4528 CLK.n10 CLK.t40 11.957
R4529 CLK.n14 CLK.t28 11.957
R4530 CLK.n20 CLK.t78 11.957
R4531 CLK.n57 CLK.t13 11.957
R4532 CLK.n52 CLK.t70 11.957
R4533 CLK.n63 CLK.t8 11.957
R4534 CLK.n68 CLK.t99 11.957
R4535 CLK.n80 CLK.t27 11.957
R4536 CLK.n72 CLK.t87 11.957
R4537 CLK.n89 CLK.t10 11.957
R4538 CLK.n3 CLK.t24 11.957
R4539 CLK CLK.n47 11.7171
R4540 CLK.n28 CLK.t21 11.6023
R4541 CLK.n35 CLK.t106 11.6023
R4542 CLK.n32 CLK.t33 11.6023
R4543 CLK.n30 CLK.t80 11.6023
R4544 CLK.n38 CLK.t102 11.6023
R4545 CLK.n41 CLK.t105 11.6023
R4546 CLK.n25 CLK.t84 11.6023
R4547 CLK.n5 CLK.t110 11.6023
R4548 CLK.n46 CLK.n45 10.9637
R4549 CLK.n16 CLK 10.8825
R4550 CLK CLK.n29 10.5737
R4551 CLK CLK.n36 10.5737
R4552 CLK.n64 CLK 10.1333
R4553 CLK CLK.n10 9.96162
R4554 CLK CLK.n63 9.96162
R4555 CLK CLK.n68 9.96162
R4556 CLK.n15 CLK.n14 9.77618
R4557 CLK.n21 CLK.n20 9.77618
R4558 CLK.n58 CLK.n57 9.77618
R4559 CLK.n53 CLK.n52 9.77618
R4560 CLK.n81 CLK.n80 9.77618
R4561 CLK.n73 CLK.n72 9.77618
R4562 CLK.n90 CLK.n89 9.77618
R4563 CLK.n4 CLK.n3 9.77618
R4564 CLK.n44 CLK.n40 9.49711
R4565 CLK.n24 CLK.n7 9.40928
R4566 CLK CLK.n33 9.27587
R4567 CLK CLK.n31 9.27587
R4568 CLK CLK.n39 9.27587
R4569 CLK CLK.n42 9.27587
R4570 CLK CLK.n26 9.27587
R4571 CLK CLK.n6 9.27587
R4572 CLK.n76 CLK.t35 9.20812
R4573 CLK.n29 CLK.t104 9.1255
R4574 CLK.n36 CLK.t44 9.1255
R4575 CLK.n48 CLK.n24 8.87892
R4576 CLK CLK.n76 8.68152
R4577 CLK.n82 CLK 8.10194
R4578 CLK.n23 CLK.n22 8.05322
R4579 CLK.n92 CLK 7.82643
R4580 CLK.n33 CLK.t124 7.3005
R4581 CLK.n31 CLK.t0 7.3005
R4582 CLK.n39 CLK.t69 7.3005
R4583 CLK.n42 CLK.t82 7.3005
R4584 CLK.n26 CLK.t49 7.3005
R4585 CLK.n8 CLK.t85 7.3005
R4586 CLK.t127 CLK.n9 7.3005
R4587 CLK.n12 CLK.t76 7.3005
R4588 CLK.t121 CLK.n13 7.3005
R4589 CLK.t59 CLK.n11 7.3005
R4590 CLK.n18 CLK.t32 7.3005
R4591 CLK.t123 CLK.n19 7.3005
R4592 CLK.t93 CLK.n17 7.3005
R4593 CLK.n6 CLK.t57 7.3005
R4594 CLK.n55 CLK.t26 7.3005
R4595 CLK.t100 CLK.n56 7.3005
R4596 CLK.t18 CLK.n54 7.3005
R4597 CLK.n50 CLK.t5 7.3005
R4598 CLK.t14 CLK.n51 7.3005
R4599 CLK.t60 CLK.n49 7.3005
R4600 CLK.n61 CLK.t7 7.3005
R4601 CLK.t38 CLK.n62 7.3005
R4602 CLK.n66 CLK.t73 7.3005
R4603 CLK.t41 CLK.n67 7.3005
R4604 CLK.n78 CLK.t46 7.3005
R4605 CLK.t68 CLK.n79 7.3005
R4606 CLK.t19 CLK.n77 7.3005
R4607 CLK.n74 CLK.t64 7.3005
R4608 CLK.t86 CLK.n75 7.3005
R4609 CLK.n70 CLK.t98 7.3005
R4610 CLK.t52 CLK.n71 7.3005
R4611 CLK.t55 CLK.n69 7.3005
R4612 CLK.n87 CLK.t37 7.3005
R4613 CLK.t96 CLK.n88 7.3005
R4614 CLK.t15 CLK.n86 7.3005
R4615 CLK.n1 CLK.t47 7.3005
R4616 CLK.t56 CLK.n2 7.3005
R4617 CLK.t17 CLK.n0 7.3005
R4618 CLK.n34 CLK 6.38571
R4619 CLK.n83 CLK.n82 6.20465
R4620 CLK.n47 CLK.n27 4.88121
R4621 CLK.n45 CLK.n37 4.83739
R4622 CLK.n46 CLK 4.8335
R4623 CLK.n85 CLK.n65 4.81202
R4624 CLK.n37 CLK 4.53484
R4625 CLK.n34 CLK 4.51896
R4626 CLK.n23 CLK.n16 4.50961
R4627 CLK.n65 CLK.n48 4.17208
R4628 CLK.n82 CLK 3.83185
R4629 CLK.n37 CLK.n34 3.08408
R4630 CLK.n47 CLK.n46 2.40407
R4631 CLK CLK.n85 1.33289
R4632 CLK.n85 CLK.n84 1.08658
R4633 CLK.n16 CLK 0.81937
R4634 CLK.n60 CLK 0.81937
R4635 CLK CLK.n92 0.81937
R4636 CLK.n64 CLK.n60 0.749691
R4637 CLK.n84 CLK 0.473978
R4638 CLK CLK.n15 0.185948
R4639 CLK CLK.n53 0.185948
R4640 CLK CLK.n73 0.185948
R4641 CLK CLK.n4 0.185948
R4642 CLK CLK.n81 0.183616
R4643 CLK.n40 CLK 0.183172
R4644 CLK CLK.n21 0.181221
R4645 CLK CLK.n58 0.181221
R4646 CLK CLK.n90 0.181221
R4647 CLK.n43 CLK 0.141537
R4648 CLK.n22 CLK 0.0449156
R4649 CLK.n59 CLK 0.0449156
R4650 CLK.n91 CLK 0.0449156
R4651 CLK.n22 CLK 0.0332273
R4652 CLK.n59 CLK 0.0332273
R4653 CLK.n91 CLK 0.0332273
R4654 CLK.n43 CLK 0.0329
R4655 CLK.n27 CLK 0.0123421
R4656 CLK.n7 CLK 0.01175
R4657 CLK.n27 CLK 0.0111579
R4658 CLK.n7 CLK 0.010625
R4659 CLK.n40 CLK 0.00517532
R4660 VSS.n1952 VSS.n1066 7.02563e+06
R4661 VSS.n1989 VSS.t19 952901
R4662 VSS.n1130 VSS.n1129 216125
R4663 VSS.n1969 VSS.n1039 216125
R4664 VSS.n142 VSS.n114 216125
R4665 VSS.n2879 VSS.n2878 216125
R4666 VSS.n1889 VSS.n1428 216125
R4667 VSS.n1840 VSS.n1821 216125
R4668 VSS.t733 VSS.n1953 170380
R4669 VSS.t1116 VSS.n2 133419
R4670 VSS.n2906 VSS.n2 57096.1
R4671 VSS.n1953 VSS.n1064 57034.3
R4672 VSS.n65 VSS.n22 42762.3
R4673 VSS.n2777 VSS.n2776 42503.8
R4674 VSS.t1071 VSS.t824 42027.8
R4675 VSS.t1067 VSS.t817 42027.8
R4676 VSS.t1037 VSS.t369 41809.4
R4677 VSS.t1135 VSS.t280 41809.4
R4678 VSS.t1130 VSS.t166 41809.4
R4679 VSS.t1179 VSS.t378 41809.4
R4680 VSS.n1064 VSS.t1109 40174.8
R4681 VSS.n2779 VSS.n64 34205.5
R4682 VSS.n1186 VSS.n1067 33626.6
R4683 VSS.n1422 VSS.n1067 31810.9
R4684 VSS.n1186 VSS.n1185 25310.9
R4685 VSS.n2776 VSS.n67 19756
R4686 VSS.n1596 VSS.n1064 18483.1
R4687 VSS.n1104 VSS.n67 17380.9
R4688 VSS.n1993 VSS.t730 15929
R4689 VSS.n2435 VSS.n63 15509.4
R4690 VSS.n1185 VSS.n64 15026.9
R4691 VSS.n2905 VSS.n2904 13611.1
R4692 VSS.n1910 VSS.n1424 12835.5
R4693 VSS.n2829 VSS.n21 12239.9
R4694 VSS.n1320 VSS.t756 12172.3
R4695 VSS.t284 VSS.n1424 12050.7
R4696 VSS.n2542 VSS.n64 12047.2
R4697 VSS.n2776 VSS.n2775 12047.2
R4698 VSS.n2037 VSS.n2036 8490.89
R4699 VSS.n2027 VSS.n565 8044.55
R4700 VSS.n2905 VSS.n3 8008.43
R4701 VSS.n1104 VSS.n5 7098.75
R4702 VSS.n1829 VSS.n2 7002.9
R4703 VSS.t1161 VSS.t707 6847.71
R4704 VSS.t1154 VSS.t701 6847.71
R4705 VSS.t428 VSS.t1048 6829.13
R4706 VSS.t1043 VSS.t380 6829.13
R4707 VSS.n2778 VSS.n2777 6658.88
R4708 VSS.n66 VSS.n65 6624.26
R4709 VSS.n1993 VSS.t64 6019.86
R4710 VSS.n2037 VSS.n561 5714.4
R4711 VSS.n1423 VSS.n23 5530.63
R4712 VSS.n21 VSS.n5 5241.73
R4713 VSS.n2904 VSS.n4 5123.32
R4714 VSS.n2829 VSS.n2828 5035.12
R4715 VSS.n1392 VSS.n1186 4922.24
R4716 VSS.n1087 VSS.t438 4869.56
R4717 VSS VSS.n1320 4818.45
R4718 VSS.n1182 VSS.t838 4530.79
R4719 VSS.n2435 VSS.n2434 4483.26
R4720 VSS.n1947 VSS.n1067 4291.67
R4721 VSS.n1185 VSS.n1184 3845.48
R4722 VSS.n200 VSS.n67 3818.95
R4723 VSS.t190 VSS.n1104 3722.48
R4724 VSS.n1422 VSS.n3 3720.83
R4725 VSS.t231 VSS.t286 3685.04
R4726 VSS.n2037 VSS.n560 3443.07
R4727 VSS.n2779 VSS.n2778 3352.96
R4728 VSS.n2777 VSS.n66 3352.96
R4729 VSS.n1952 VSS.t152 3250.86
R4730 VSS.n2780 VSS.n2779 3142.25
R4731 VSS.n2903 VSS.t1203 3046.22
R4732 VSS.t780 VSS.t792 2937.24
R4733 VSS.t794 VSS.t784 2937.24
R4734 VSS.t838 VSS.t836 2881.77
R4735 VSS.t1035 VSS.t922 2827.3
R4736 VSS.n2827 VSS.n23 2515.11
R4737 VSS.t798 VSS.t720 2456.82
R4738 VSS.t256 VSS.t969 2368.09
R4739 VSS.n1953 VSS.n1952 2355.86
R4740 VSS.t220 VSS.t749 2072.98
R4741 VSS.t277 VSS.t752 2072.98
R4742 VSS.n2780 VSS.n63 1995.52
R4743 VSS.n2027 VSS.n2026 1892.95
R4744 VSS.t1081 VSS.t1079 1842.52
R4745 VSS.t1079 VSS.t232 1842.52
R4746 VSS.n2827 VSS.n24 1827
R4747 VSS.t98 VSS.t585 1824.89
R4748 VSS.t536 VSS.t14 1824.89
R4749 VSS.t658 VSS.t903 1824.89
R4750 VSS.t840 VSS.t1229 1824.89
R4751 VSS.t30 VSS.t689 1824.89
R4752 VSS.t956 VSS.t1148 1824.89
R4753 VSS.n2778 VSS.t1256 1779.25
R4754 VSS.n66 VSS.t1263 1779.25
R4755 VSS.n1424 VSS.n1423 1769.44
R4756 VSS.t505 VSS.t847 1705.23
R4757 VSS.t349 VSS.t561 1705.23
R4758 VSS.t303 VSS.t83 1705.23
R4759 VSS.t1268 VSS.t540 1705.23
R4760 VSS.t223 VSS.t1099 1705.23
R4761 VSS.t263 VSS.t868 1705.23
R4762 VSS.t24 VSS.t848 1701.21
R4763 VSS.t47 VSS.t554 1701.21
R4764 VSS.t1240 VSS.t70 1701.21
R4765 VSS.t40 VSS.t541 1701.21
R4766 VSS.t892 VSS.t1105 1701.21
R4767 VSS.t948 VSS.t869 1701.21
R4768 VSS.t850 VSS.t27 1699.79
R4769 VSS.t553 VSS.t59 1699.79
R4770 VSS.t36 VSS.t1239 1699.79
R4771 VSS.t1106 VSS.t101 1699.79
R4772 VSS.t1101 VSS.t909 1699.79
R4773 VSS.t947 VSS.t865 1699.79
R4774 VSS.t1029 VSS.n22 1584.15
R4775 VSS.t1256 VSS.t1254 1549.67
R4776 VSS.t1263 VSS.t1261 1549.67
R4777 VSS.n1912 VSS.n1422 1515.27
R4778 VSS.t724 VSS.n565 1506.44
R4779 VSS.n1757 VSS.n1596 1496.69
R4780 VSS.t152 VSS.n1951 1475.68
R4781 VSS.n2121 VSS.t170 1439.43
R4782 VSS.n2094 VSS.t1168 1439.43
R4783 VSS.n2197 VSS.t339 1439.43
R4784 VSS.n2186 VSS.t219 1439.43
R4785 VSS.t335 VSS.n1318 1439.43
R4786 VSS.n1361 VSS.t914 1439.43
R4787 VSS.n1342 VSS.t359 1439.43
R4788 VSS.n1330 VSS.t278 1439.43
R4789 VSS.n1257 VSS.t589 1439.43
R4790 VSS.n1401 VSS.t913 1439.43
R4791 VSS.n1927 VSS.t354 1439.43
R4792 VSS.n1939 VSS.t935 1439.43
R4793 VSS.n1387 VSS.t938 1439.43
R4794 VSS.n1374 VSS.t911 1439.43
R4795 VSS.n1227 VSS.t356 1439.43
R4796 VSS.n2104 VSS.t108 1439.43
R4797 VSS.n2080 VSS.t116 1439.43
R4798 VSS.t343 VSS.n2163 1439.43
R4799 VSS.t469 VSS.n2178 1439.43
R4800 VSS.t891 VSS.n2057 1439.43
R4801 VSS.n1872 VSS.t457 1439.43
R4802 VSS.t712 VSS.n1057 1374.84
R4803 VSS.t886 VSS.n2542 1374.11
R4804 VSS.n2775 VSS.t882 1374.11
R4805 VSS.n2904 VSS.n2903 1342.09
R4806 VSS.n1129 VSS.t851 1317.42
R4807 VSS.t558 VSS.n1969 1317.42
R4808 VSS.t33 VSS.n142 1317.42
R4809 VSS.n2878 VSS.t550 1317.42
R4810 VSS.t1102 VSS.n1889 1317.42
R4811 VSS.n1821 VSS.t861 1317.42
R4812 VSS.n2828 VSS.n22 1301.11
R4813 VSS.t811 VSS.t1211 1301.04
R4814 VSS.t822 VSS.t1223 1301.04
R4815 VSS.t1185 VSS.t1162 1290.61
R4816 VSS.t1199 VSS.t1157 1290.61
R4817 VSS.n202 VSS.n201 1273.97
R4818 VSS.t738 VSS.n565 1272.89
R4819 VSS.t971 VSS.t1253 1205.23
R4820 VSS.t967 VSS.t1260 1205.23
R4821 VSS.t829 VSS.n3 1183.66
R4822 VSS.t1146 VSS.n21 1183.26
R4823 VSS.t171 VSS.n2120 1153.55
R4824 VSS.n2120 VSS.t1169 1153.55
R4825 VSS.n2206 VSS.t340 1153.55
R4826 VSS.n1319 VSS.t336 1153.55
R4827 VSS.n1366 VSS.t915 1153.55
R4828 VSS.t360 VSS.n1341 1153.55
R4829 VSS.n1366 VSS.t590 1153.55
R4830 VSS.t912 VSS.n1400 1153.55
R4831 VSS.n1938 VSS.t353 1153.55
R4832 VSS.t936 VSS.n1938 1153.55
R4833 VSS.t937 VSS.n1386 1153.55
R4834 VSS.t910 VSS.n1373 1153.55
R4835 VSS.n1373 VSS.t355 1153.55
R4836 VSS.t107 VSS.n2103 1153.55
R4837 VSS.n2103 VSS.t117 1153.55
R4838 VSS.n2179 VSS.t344 1153.55
R4839 VSS.n2179 VSS.t468 1153.55
R4840 VSS.n2058 VSS.t890 1153.55
R4841 VSS.t456 VSS.n1871 1153.55
R4842 VSS.n1057 VSS.t575 1151.13
R4843 VSS.n2039 VSS.n2038 1136.96
R4844 VSS.n2903 VSS.n5 1126.94
R4845 VSS.t210 VSS.n1296 1088.19
R4846 VSS.t113 VSS.n2161 1088.19
R4847 VSS.t365 VSS.t367 1088.19
R4848 VSS.t148 VSS.t928 1088.19
R4849 VSS.t314 VSS.t124 1088.19
R4850 VSS.t216 VSS.t186 1088.19
R4851 VSS.t178 VSS.t361 1088.19
R4852 VSS.t699 VSS.t171 1083.33
R4853 VSS.t703 VSS.t699 1083.33
R4854 VSS.t170 VSS.t703 1083.33
R4855 VSS.t126 VSS.t1169 1083.33
R4856 VSS.t128 VSS.t126 1083.33
R4857 VSS.t1168 VSS.t128 1083.33
R4858 VSS.t442 VSS.t340 1083.33
R4859 VSS.t440 VSS.t442 1083.33
R4860 VSS.t339 VSS.t440 1083.33
R4861 VSS.t219 VSS.t142 1083.33
R4862 VSS.t142 VSS.t140 1083.33
R4863 VSS.t140 VSS.t220 1083.33
R4864 VSS.t872 VSS.t335 1083.33
R4865 VSS.t875 VSS.t872 1083.33
R4866 VSS.t336 VSS.t875 1083.33
R4867 VSS.t1164 VSS.t915 1083.33
R4868 VSS.t1166 VSS.t1164 1083.33
R4869 VSS.t914 VSS.t1166 1083.33
R4870 VSS.t406 VSS.t360 1083.33
R4871 VSS.t404 VSS.t406 1083.33
R4872 VSS.t359 VSS.t404 1083.33
R4873 VSS.t278 VSS.t483 1083.33
R4874 VSS.t483 VSS.t481 1083.33
R4875 VSS.t481 VSS.t277 1083.33
R4876 VSS.t567 VSS.t590 1083.33
R4877 VSS.t569 VSS.t567 1083.33
R4878 VSS.t589 VSS.t569 1083.33
R4879 VSS.t418 VSS.t912 1083.33
R4880 VSS.t420 VSS.t418 1083.33
R4881 VSS.t913 VSS.t420 1083.33
R4882 VSS.t962 VSS.t353 1083.33
R4883 VSS.t959 VSS.t962 1083.33
R4884 VSS.t354 VSS.t959 1083.33
R4885 VSS.t532 VSS.t936 1083.33
R4886 VSS.t530 VSS.t532 1083.33
R4887 VSS.t935 VSS.t530 1083.33
R4888 VSS.t938 VSS.t237 1083.33
R4889 VSS.t237 VSS.t235 1083.33
R4890 VSS.t235 VSS.t937 1083.33
R4891 VSS.t911 VSS.t1063 1083.33
R4892 VSS.t1063 VSS.t1065 1083.33
R4893 VSS.t1065 VSS.t910 1083.33
R4894 VSS.t356 VSS.t522 1083.33
R4895 VSS.t522 VSS.t524 1083.33
R4896 VSS.t524 VSS.t355 1083.33
R4897 VSS.t108 VSS.t8 1083.33
R4898 VSS.t8 VSS.t102 1083.33
R4899 VSS.t102 VSS.t107 1083.33
R4900 VSS.t116 VSS.t973 1083.33
R4901 VSS.t973 VSS.t975 1083.33
R4902 VSS.t975 VSS.t117 1083.33
R4903 VSS.t134 VSS.t343 1083.33
R4904 VSS.t136 VSS.t134 1083.33
R4905 VSS.t344 VSS.t136 1083.33
R4906 VSS.t815 VSS.t469 1083.33
R4907 VSS.t818 VSS.t815 1083.33
R4908 VSS.t468 VSS.t818 1083.33
R4909 VSS.t197 VSS.t891 1083.33
R4910 VSS.t195 VSS.t197 1083.33
R4911 VSS.t890 VSS.t195 1083.33
R4912 VSS.t457 VSS.t652 1083.33
R4913 VSS.t652 VSS.t654 1083.33
R4914 VSS.t654 VSS.t456 1083.33
R4915 VSS.n1394 VSS.n1086 1067.69
R4916 VSS.t648 VSS.n1066 1060.95
R4917 VSS.n1147 VSS.t189 987.038
R4918 VSS.n185 VSS.t1108 982.878
R4919 VSS.n1054 VSS.t579 977.444
R4920 VSS.t1113 VSS.n1063 976.221
R4921 VSS.n1058 VSS.t796 976.221
R4922 VSS.n998 VSS.n566 931.149
R4923 VSS.n1129 VSS.t581 927.644
R4924 VSS.n1969 VSS.t447 927.644
R4925 VSS.n142 VSS.t1245 927.644
R4926 VSS.n2878 VSS.t503 927.644
R4927 VSS.n1889 VSS.t229 927.644
R4928 VSS.n1821 VSS.t290 927.644
R4929 VSS.n1320 VSS.t231 921.26
R4930 VSS.n1320 VSS.t1081 921.26
R4931 VSS.n1423 VSS.n1066 914.535
R4932 VSS.t212 VSS.t257 905.265
R4933 VSS.t275 VSS.t120 905.265
R4934 VSS.t245 VSS.t202 905.265
R4935 VSS.t156 VSS.t271 905.265
R4936 VSS.t316 VSS.t150 905.265
R4937 VSS.t422 VSS.t132 905.265
R4938 VSS.t247 VSS.t168 905.265
R4939 VSS.n1054 VSS.t714 895.99
R4940 VSS.n1063 VSS.t716 894.87
R4941 VSS.n1058 VSS.t726 894.87
R4942 VSS.n2038 VSS.t732 880.448
R4943 VSS.t579 VSS.t577 879.699
R4944 VSS.t714 VSS.t722 879.699
R4945 VSS.t722 VSS.t724 879.699
R4946 VSS.t577 VSS.t575 879.414
R4947 VSS.t1109 VSS.t1111 878.598
R4948 VSS.t1111 VSS.t1113 878.598
R4949 VSS.t718 VSS.t716 878.598
R4950 VSS.t720 VSS.t718 878.598
R4951 VSS.t800 VSS.t798 878.598
R4952 VSS.t796 VSS.t800 878.598
R4953 VSS.t726 VSS.t728 878.598
R4954 VSS.t728 VSS.t712 878.598
R4955 VSS.n1953 VSS.n1065 872.524
R4956 VSS.t740 VSS.t764 863.47
R4957 VSS.t775 VSS.t761 863.47
R4958 VSS.t752 VSS.n1329 859.471
R4959 VSS.t749 VSS.n2185 859.471
R4960 VSS.t297 VSS.t475 849.053
R4961 VSS.t81 VSS.n2894 831.183
R4962 VSS.t347 VSS.t345 826.856
R4963 VSS.t735 VSS.t732 826.856
R4964 VSS.n981 VSS.n560 820.544
R4965 VSS.n1086 VSS.t273 797.835
R4966 VSS.t328 VSS.t327 768.221
R4967 VSS.n2036 VSS.t705 762.755
R4968 VSS.t189 VSS.t1077 742.857
R4969 VSS.t1077 VSS.t1075 742.857
R4970 VSS.t1108 VSS.t513 739.726
R4971 VSS.t513 VSS.t511 739.726
R4972 VSS.n1989 VSS.t92 735.85
R4973 VSS.n2036 VSS.t493 733.75
R4974 VSS.n2781 VSS.n62 729.693
R4975 VSS.n2781 VSS.n24 729.611
R4976 VSS.t616 VSS.t604 728.448
R4977 VSS.t1004 VSS.t979 728.448
R4978 VSS.n1948 VSS.n1947 727.861
R4979 VSS.n2121 VSS.t693 727.239
R4980 VSS.n2094 VSS.t376 727.239
R4981 VSS.n2197 VSS.t341 727.239
R4982 VSS.n2186 VSS.t449 727.239
R4983 VSS.n1318 VSS.t221 727.239
R4984 VSS.n1361 VSS.t144 727.239
R4985 VSS.n1342 VSS.t390 727.239
R4986 VSS.n1330 VSS.t462 727.239
R4987 VSS.n1257 VSS.t233 727.239
R4988 VSS.n1401 VSS.t382 727.239
R4989 VSS.n1927 VSS.t489 727.239
R4990 VSS.n1939 VSS.t241 727.239
R4991 VSS.n1387 VSS.t239 727.239
R4992 VSS.n1374 VSS.t118 727.239
R4993 VSS.n1227 VSS.t357 727.239
R4994 VSS.n2104 VSS.t109 727.239
R4995 VSS.n2080 VSS.t154 727.239
R4996 VSS.n2163 VSS.t515 727.239
R4997 VSS.n2178 VSS.t470 727.239
R4998 VSS.n2057 VSS.t1281 727.239
R4999 VSS.n1872 VSS.t394 727.239
R5000 VSS.n107 VSS.t328 725.543
R5001 VSS.n1629 VSS.n23 720.585
R5002 VSS.t308 VSS.t436 713.264
R5003 VSS.t1075 VSS.n1146 694.71
R5004 VSS.t511 VSS.n184 691.782
R5005 VSS.t392 VSS.t425 687.824
R5006 VSS.t243 VSS.t260 687.824
R5007 VSS.t466 VSS.t199 687.824
R5008 VSS.t267 VSS.t299 677.587
R5009 VSS.n1393 VSS.n1087 676.828
R5010 VSS.n202 VSS.t661 672.193
R5011 VSS.n2894 VSS.t26 656.51
R5012 VSS.n1146 VSS.t39 625.524
R5013 VSS.n184 VSS.t1238 625.524
R5014 VSS.n1910 VSS.t893 625.524
R5015 VSS.n1829 VSS.t810 625.524
R5016 VSS.n1324 VSS.t748 619.356
R5017 VSS.n1231 VSS.t599 619.356
R5018 VSS.t611 VSS.n1365 619.356
R5019 VSS.n2068 VSS.t990 619.356
R5020 VSS.t988 VSS.n2119 619.356
R5021 VSS.n2180 VSS.t745 619.356
R5022 VSS.t613 VSS.n1937 619.356
R5023 VSS.n982 VSS.n981 618.819
R5024 VSS.n1381 VSS.t365 597.375
R5025 VSS.n1355 VSS.t148 597.375
R5026 VSS.n1325 VSS.t210 597.375
R5027 VSS.t124 VSS.n2131 597.375
R5028 VSS.n2181 VSS.t113 597.375
R5029 VSS.n2070 VSS.t216 597.375
R5030 VSS.n1936 VSS.t178 597.375
R5031 VSS.n2903 VSS.t20 592.4
R5032 VSS.t742 VSS.n2435 587.324
R5033 VSS.t888 VSS.t464 561.297
R5034 VSS.t1205 VSS.n1948 554.497
R5035 VSS.n2034 VSS.n562 543.879
R5036 VSS.n1145 VSS.t12 543.255
R5037 VSS.n180 VSS.t79 542.461
R5038 VSS.n65 VSS.n24 534.372
R5039 VSS.n2028 VSS.t735 524.441
R5040 VSS.n1912 VSS.n1911 506.974
R5041 VSS.n1147 VSS.t190 498.678
R5042 VSS.n185 VSS.t922 496.575
R5043 VSS.n1319 VSS.t751 496.349
R5044 VSS.n1373 VSS.t600 496.349
R5045 VSS.n1366 VSS.t607 496.349
R5046 VSS.n2103 VSS.t1011 496.349
R5047 VSS.n2120 VSS.t981 496.349
R5048 VSS.t747 VSS.n2179 496.349
R5049 VSS.n1938 VSS.t608 496.349
R5050 VSS.n1394 VSS.n1393 472.248
R5051 VSS.t62 VSS.t748 466.135
R5052 VSS.t31 VSS.t62 466.135
R5053 VSS.t751 VSS.t31 466.135
R5054 VSS.t599 VSS.t66 466.135
R5055 VSS.t66 VSS.t57 466.135
R5056 VSS.t57 VSS.t600 466.135
R5057 VSS.t607 VSS.t17 466.135
R5058 VSS.t17 VSS.t2 466.135
R5059 VSS.t2 VSS.t611 466.135
R5060 VSS.t990 VSS.t10 466.135
R5061 VSS.t10 VSS.t4 466.135
R5062 VSS.t4 VSS.t1011 466.135
R5063 VSS.t981 VSS.t60 466.135
R5064 VSS.t60 VSS.t55 466.135
R5065 VSS.t55 VSS.t988 466.135
R5066 VSS.t745 VSS.t71 466.135
R5067 VSS.t71 VSS.t43 466.135
R5068 VSS.t43 VSS.t747 466.135
R5069 VSS.t608 VSS.t50 466.135
R5070 VSS.t50 VSS.t53 466.135
R5071 VSS.t53 VSS.t613 466.135
R5072 VSS.t852 VSS.t98 449.122
R5073 VSS.t851 VSS.t41 449.122
R5074 VSS.t14 VSS.t562 449.122
R5075 VSS.t73 VSS.t558 449.122
R5076 VSS.t1229 VSS.t28 449.122
R5077 VSS.t1241 VSS.t33 449.122
R5078 VSS.t551 VSS.t30 449.122
R5079 VSS.t550 VSS.t77 449.122
R5080 VSS.t903 VSS.t1096 449.122
R5081 VSS.t907 VSS.t1102 449.122
R5082 VSS.t863 VSS.t956 449.122
R5083 VSS.t861 VSS.t954 449.122
R5084 VSS.t847 VSS.t88 448.745
R5085 VSS.t856 VSS.t39 448.745
R5086 VSS.t561 VSS.t34 448.745
R5087 VSS.t19 VSS.t559 448.745
R5088 VSS.t83 VSS.t1230 448.745
R5089 VSS.t1238 VSS.t75 448.745
R5090 VSS.t540 VSS.t90 448.745
R5091 VSS.t546 VSS.t26 448.745
R5092 VSS.t1099 VSS.t895 448.745
R5093 VSS.t893 VSS.t1094 448.745
R5094 VSS.t868 VSS.t949 448.745
R5095 VSS.t810 VSS.t859 448.745
R5096 VSS.t943 VSS.n4 436.135
R5097 VSS.n2778 VSS.t964 423.776
R5098 VSS.t957 VSS.n66 423.776
R5099 VSS.n1951 VSS.t1205 421.623
R5100 VSS.t874 VSS.t454 418.253
R5101 VSS.t252 VSS.t881 418.253
R5102 VSS.n107 VSS.t371 415.048
R5103 VSS.t966 VSS.t310 405.483
R5104 VSS.t1062 VSS.t194 405.483
R5105 VSS.t1059 VSS.t249 405.483
R5106 VSS.t961 VSS.t492 405.483
R5107 VSS.n171 VSS.t1029 397.815
R5108 VSS.t933 VSS.t255 388.274
R5109 VSS.t120 VSS.t158 384.026
R5110 VSS.t146 VSS.t245 384.026
R5111 VSS.t478 VSS.t212 384.026
R5112 VSS.t150 VSS.t122 384.026
R5113 VSS.t111 VSS.t422 384.026
R5114 VSS.t214 VSS.t156 384.026
R5115 VSS.t168 VSS.t176 384.026
R5116 VSS.t1073 VSS.n559 371.43
R5117 VSS.n1034 VSS.t738 370.296
R5118 VSS.n171 VSS.t1035 369.399
R5119 VSS.t730 VSS.n1034 343.846
R5120 VSS.t255 VSS.t939 343.034
R5121 VSS.n1155 VSS.t931 341.918
R5122 VSS.t373 VSS.n199 341.418
R5123 VSS.t412 VSS.t1172 334.925
R5124 VSS.t411 VSS.t412 334.925
R5125 VSS.t1174 VSS.t411 334.925
R5126 VSS.t338 VSS.t681 334.925
R5127 VSS.t337 VSS.t338 334.925
R5128 VSS.t677 VSS.t337 334.925
R5129 VSS.n1392 VSS.t282 329.661
R5130 VSS.t451 VSS.n4 328.772
R5131 VSS.n1336 VSS.t253 316.466
R5132 VSS.t192 VSS.n1335 316.466
R5133 VSS.n2192 VSS.t498 316.293
R5134 VSS.t918 VSS.n2191 316.293
R5135 VSS.n1832 VSS.t952 314.183
R5136 VSS.t257 VSS.n1324 312.916
R5137 VSS.n1231 VSS.t275 312.916
R5138 VSS.n1365 VSS.t202 312.916
R5139 VSS.t271 VSS.n2068 312.916
R5140 VSS.n2119 VSS.t316 312.916
R5141 VSS.t132 VSS.n2180 312.916
R5142 VSS.n1937 VSS.t247 312.916
R5143 VSS.t476 VSS.t172 311.447
R5144 VSS.t175 VSS.t252 311.447
R5145 VSS.t454 VSS.t802 311.447
R5146 VSS.t438 VSS.t308 311.034
R5147 VSS.t104 VSS.t392 311.033
R5148 VSS.t916 VSS.t243 311.033
R5149 VSS.t199 VSS.t318 311.033
R5150 VSS.t299 VSS.t269 304.029
R5151 VSS.n2028 VSS.t347 302.416
R5152 VSS.n2830 VSS.t451 293.077
R5153 VSS.n1117 VSS.t844 291.248
R5154 VSS.t15 VSS.n1107 291.248
R5155 VSS.n1963 VSS.t565 291.248
R5156 VSS.n1968 VSS.t6 291.248
R5157 VSS.n136 VSS.t99 291.248
R5158 VSS.n141 VSS.t1232 291.248
R5159 VSS.n2866 VSS.t548 291.248
R5160 VSS.t22 VSS.n2852 291.248
R5161 VSS.n1883 VSS.t1103 291.248
R5162 VSS.n1888 VSS.t901 291.248
R5163 VSS.n1853 VSS.t866 291.248
R5164 VSS.t945 VSS.n1852 291.248
R5165 VSS.n1136 VSS.t45 291.005
R5166 VSS.n1140 VSS.t854 291.005
R5167 VSS.n1984 VSS.t0 291.005
R5168 VSS.t556 VSS.n1036 291.005
R5169 VSS.n158 VSS.t1236 291.005
R5170 VSS.t96 VSS.n111 291.005
R5171 VSS.n2885 VSS.t37 291.005
R5172 VSS.n2889 VSS.t542 291.005
R5173 VSS.n1904 VSS.t899 291.005
R5174 VSS.t1092 VSS.n1425 291.005
R5175 VSS.t807 VSS.n1823 291.005
R5176 VSS.n1836 VSS.t870 291.005
R5177 VSS.n2038 VSS.n2037 284.241
R5178 VSS.t253 VSS.t192 280.909
R5179 VSS.t498 VSS.t918 280.755
R5180 VSS.n108 VSS.n107 275.279
R5181 VSS.t756 VSS.n1319 260.909
R5182 VSS.t931 VSS.t487 257.332
R5183 VSS.t162 VSS.t373 256.955
R5184 VSS.n1295 VSS.t1174 248.093
R5185 VSS.n2160 VSS.t677 248.093
R5186 VSS.t305 VSS.t428 245.748
R5187 VSS.t698 VSS.t1161 245.748
R5188 VSS.t380 VSS.t926 245.748
R5189 VSS.t711 VSS.t1154 245.748
R5190 VSS.t432 VSS.n1346 243.44
R5191 VSS.n1286 VSS.t184 243.44
R5192 VSS.n2140 VSS.t413 243.44
R5193 VSS.n2151 VSS.t322 243.44
R5194 VSS.n2052 VSS.t1085 243.44
R5195 VSS.t460 VSS.n1405 243.44
R5196 VSS.n1391 VSS.t399 243.44
R5197 VSS.n1182 VSS.t476 242.237
R5198 VSS.n1373 VSS.t622 238.666
R5199 VSS.t626 VSS.n1366 238.666
R5200 VSS.n2103 VSS.t982 238.666
R5201 VSS.n2120 VSS.t984 238.666
R5202 VSS.n2179 VSS.t754 238.666
R5203 VSS.n1947 VSS.t624 238.666
R5204 VSS.n1938 VSS.t593 238.666
R5205 VSS.t939 VSS.n1993 237.25
R5206 VSS.t485 VSS.n1183 234.696
R5207 VSS.n201 VSS.t160 234.352
R5208 VSS.n2040 VSS.t877 228.292
R5209 VSS.t604 VSS.t632 224.138
R5210 VSS.t591 VSS.t616 224.138
R5211 VSS.t986 VSS.t1004 224.138
R5212 VSS.t979 VSS.t1002 224.138
R5213 VSS.t766 VSS.t742 224.138
R5214 VSS.t624 VSS.t597 224.138
R5215 VSS.t768 VSS.t771 224.138
R5216 VSS.t371 VSS.n103 223.766
R5217 VSS.n1166 VSS.t297 223.766
R5218 VSS.n1341 VSS.t1250 223.282
R5219 VSS.n2206 VSS.t204 223.282
R5220 VSS.t1271 VSS.n2058 223.282
R5221 VSS.n1400 VSS.t685 223.282
R5222 VSS.n1386 VSS.t384 223.282
R5223 VSS.t756 VSS.n384 223.101
R5224 VSS.t622 VSS.n1372 223.101
R5225 VSS.n1367 VSS.t626 223.101
R5226 VSS.t982 VSS.n2102 223.101
R5227 VSS.n2101 VSS.t984 223.101
R5228 VSS.n2436 VSS.t754 223.101
R5229 VSS.n1946 VSS.t593 223.101
R5230 VSS.t475 VSS.t665 222.05
R5231 VSS.n998 VSS.n997 218.912
R5232 VSS.n997 VSS.n996 218.912
R5233 VSS.n996 VSS.n601 218.912
R5234 VSS.n990 VSS.n601 218.912
R5235 VSS.n990 VSS.n989 218.912
R5236 VSS.n989 VSS.n988 218.912
R5237 VSS.n988 VSS.n606 218.912
R5238 VSS.n982 VSS.n606 218.912
R5239 VSS.t295 VSS.n2475 217.077
R5240 VSS.t164 VSS.n2493 217.077
R5241 VSS.t472 VSS.n2735 217.077
R5242 VSS.t495 VSS.n2717 217.077
R5243 VSS.t969 VSS.n2039 215.561
R5244 VSS.n1395 VSS.n1394 215.53
R5245 VSS.n258 VSS.t106 210.934
R5246 VSS.n2589 VSS.t403 210.934
R5247 VSS.t1026 VSS.n2905 209.091
R5248 VSS.n201 VSS.n108 206.994
R5249 VSS.n2895 VSS.t81 204.15
R5250 VSS.t615 VSS.t430 201.575
R5251 VSS.t1053 VSS.t1247 201.575
R5252 VSS.t1057 VSS.t1252 201.575
R5253 VSS.t628 VSS.t432 201.575
R5254 VSS.t184 VSS.t760 201.575
R5255 VSS.t1176 VSS.t669 201.575
R5256 VSS.t1171 VSS.t674 201.575
R5257 VSS.t182 VSS.t746 201.575
R5258 VSS.t415 VSS.t989 201.575
R5259 VSS.t207 VSS.t786 201.575
R5260 VSS.t206 VSS.t788 201.575
R5261 VSS.t413 VSS.t998 201.575
R5262 VSS.t322 VSS.t758 201.575
R5263 VSS.t679 VSS.t1132 201.575
R5264 VSS.t680 VSS.t1139 201.575
R5265 VSS.t320 VSS.t744 201.575
R5266 VSS.t1085 VSS.t1015 201.575
R5267 VSS.t1274 VSS.t1017 201.575
R5268 VSS.t1273 VSS.t1021 201.575
R5269 VSS.t1087 VSS.t1016 201.575
R5270 VSS.t644 VSS.t458 201.575
R5271 VSS.t1215 VSS.t687 201.575
R5272 VSS.t1227 VSS.t688 201.575
R5273 VSS.t614 VSS.t460 201.575
R5274 VSS.t610 VSS.t399 201.575
R5275 VSS.t1191 VSS.t387 201.575
R5276 VSS.t1195 VSS.t386 201.575
R5277 VSS.t612 VSS.t401 201.575
R5278 VSS.t831 VSS.n2829 200.618
R5279 VSS.t804 VSS.t874 200.305
R5280 VSS.t881 VSS.t1207 200.305
R5281 VSS.n1184 VSS.t487 200.148
R5282 VSS.n200 VSS.t162 199.855
R5283 VSS.t106 VSS.t698 196.597
R5284 VSS.t403 VSS.t711 196.597
R5285 VSS.t1019 VSS.t1026 196.364
R5286 VSS.t464 VSS.t434 193.017
R5287 VSS.n2895 VSS.t20 189.569
R5288 VSS.t218 VSS.t804 189.478
R5289 VSS.t1207 VSS.t181 189.478
R5290 VSS.t1142 VSS.t831 188.406
R5291 VSS.n212 VSS.n211 187.674
R5292 VSS.n1176 VSS.n1096 187.674
R5293 VSS.n212 VSS.t218 185.869
R5294 VSS.t181 VSS.n1176 185.869
R5295 VSS.n1087 VSS.t330 185.817
R5296 VSS.t518 VSS.t409 185.346
R5297 VSS.n1992 VSS.t92 180.736
R5298 VSS.n980 VSS.n610 179.448
R5299 VSS.n974 VSS.n973 179.448
R5300 VSS.n973 VSS.n972 179.448
R5301 VSS.n972 VSS.n637 179.448
R5302 VSS.n966 VSS.n637 179.448
R5303 VSS.n966 VSS.n965 179.448
R5304 VSS.n965 VSS.n964 179.448
R5305 VSS.n964 VSS.n641 179.448
R5306 VSS.n958 VSS.n641 179.448
R5307 VSS.n958 VSS.n957 179.448
R5308 VSS.n957 VSS.n956 179.448
R5309 VSS.n956 VSS.n645 179.448
R5310 VSS.n950 VSS.n645 179.448
R5311 VSS.n950 VSS.n949 179.448
R5312 VSS.n949 VSS.n948 179.448
R5313 VSS.n948 VSS.n649 179.448
R5314 VSS.n942 VSS.n649 179.448
R5315 VSS.n942 VSS.n941 179.448
R5316 VSS.n941 VSS.n940 179.448
R5317 VSS.n940 VSS.n653 179.448
R5318 VSS.n934 VSS.n653 179.448
R5319 VSS.n934 VSS.n933 179.448
R5320 VSS.n933 VSS.n932 179.448
R5321 VSS.n932 VSS.n657 179.448
R5322 VSS.n926 VSS.n657 179.448
R5323 VSS.n926 VSS.n925 179.448
R5324 VSS.n925 VSS.n924 179.448
R5325 VSS.n924 VSS.n661 179.448
R5326 VSS.n913 VSS.n661 179.448
R5327 VSS.n913 VSS.n912 179.448
R5328 VSS.n912 VSS.n911 179.448
R5329 VSS.n911 VSS.n691 179.448
R5330 VSS.n905 VSS.n691 179.448
R5331 VSS.n905 VSS.n904 179.448
R5332 VSS.n904 VSS.n903 179.448
R5333 VSS.n903 VSS.n695 179.448
R5334 VSS.n897 VSS.n695 179.448
R5335 VSS.n897 VSS.n896 179.448
R5336 VSS.n896 VSS.n895 179.448
R5337 VSS.n895 VSS.n699 179.448
R5338 VSS.n889 VSS.n699 179.448
R5339 VSS.n889 VSS.n888 179.448
R5340 VSS.n888 VSS.n887 179.448
R5341 VSS.n887 VSS.n703 179.448
R5342 VSS.n881 VSS.n703 179.448
R5343 VSS.n881 VSS.n880 179.448
R5344 VSS.n880 VSS.n879 179.448
R5345 VSS.n879 VSS.n707 179.448
R5346 VSS.n873 VSS.n707 179.448
R5347 VSS.n873 VSS.n872 179.448
R5348 VSS.n872 VSS.n871 179.448
R5349 VSS.n871 VSS.n711 179.448
R5350 VSS.n865 VSS.n711 179.448
R5351 VSS.n865 VSS.n864 179.448
R5352 VSS.n864 VSS.n863 179.448
R5353 VSS.n863 VSS.n715 179.448
R5354 VSS.n857 VSS.n715 179.448
R5355 VSS.n857 VSS.n856 179.448
R5356 VSS.n856 VSS.n855 179.448
R5357 VSS.n855 VSS.n719 179.448
R5358 VSS.n849 VSS.n719 179.448
R5359 VSS.n849 VSS.n848 179.448
R5360 VSS.n848 VSS.n847 179.448
R5361 VSS.n847 VSS.n723 179.448
R5362 VSS.n841 VSS.n723 179.448
R5363 VSS.n841 VSS.n840 179.448
R5364 VSS.n840 VSS.n839 179.448
R5365 VSS.n839 VSS.n727 179.448
R5366 VSS.n833 VSS.n727 179.448
R5367 VSS.n833 VSS.n832 179.448
R5368 VSS.n832 VSS.n831 179.448
R5369 VSS.n831 VSS.n731 179.448
R5370 VSS.n825 VSS.n731 179.448
R5371 VSS.n825 VSS.n824 179.448
R5372 VSS.n824 VSS.n823 179.448
R5373 VSS.n823 VSS.n735 179.448
R5374 VSS.n817 VSS.n735 179.448
R5375 VSS.n817 VSS.n816 179.448
R5376 VSS.n816 VSS.n815 179.448
R5377 VSS.n815 VSS.n739 179.448
R5378 VSS.n809 VSS.n739 179.448
R5379 VSS.n809 VSS.n808 179.448
R5380 VSS.n808 VSS.n807 179.448
R5381 VSS.n807 VSS.n743 179.448
R5382 VSS.n801 VSS.n743 179.448
R5383 VSS.n801 VSS.n800 179.448
R5384 VSS.n800 VSS.n799 179.448
R5385 VSS.n799 VSS.n747 179.448
R5386 VSS.n793 VSS.n747 179.448
R5387 VSS.n793 VSS.n792 179.448
R5388 VSS.n792 VSS.n791 179.448
R5389 VSS.n791 VSS.n751 179.448
R5390 VSS.n762 VSS.n751 179.448
R5391 VSS.n779 VSS.n762 179.448
R5392 VSS.n779 VSS.n778 179.448
R5393 VSS.n778 VSS.n777 179.448
R5394 VSS.n777 VSS.n500 179.448
R5395 VSS.n2220 VSS.n500 179.448
R5396 VSS.n2221 VSS.n2220 179.448
R5397 VSS.n2222 VSS.n2221 179.448
R5398 VSS.n2222 VSS.n496 179.448
R5399 VSS.n2228 VSS.n496 179.448
R5400 VSS.n2229 VSS.n2228 179.448
R5401 VSS.n2230 VSS.n2229 179.448
R5402 VSS.n2230 VSS.n492 179.448
R5403 VSS.n2236 VSS.n492 179.448
R5404 VSS.n2237 VSS.n2236 179.448
R5405 VSS.n2238 VSS.n2237 179.448
R5406 VSS.n2238 VSS.n488 179.448
R5407 VSS.n2244 VSS.n488 179.448
R5408 VSS.n2245 VSS.n2244 179.448
R5409 VSS.n2246 VSS.n2245 179.448
R5410 VSS.n2246 VSS.n484 179.448
R5411 VSS.n2252 VSS.n484 179.448
R5412 VSS.n2253 VSS.n2252 179.448
R5413 VSS.n2254 VSS.n2253 179.448
R5414 VSS.n2254 VSS.n480 179.448
R5415 VSS.n2260 VSS.n480 179.448
R5416 VSS.n2261 VSS.n2260 179.448
R5417 VSS.n2262 VSS.n2261 179.448
R5418 VSS.n2262 VSS.n476 179.448
R5419 VSS.n2268 VSS.n476 179.448
R5420 VSS.n2269 VSS.n2268 179.448
R5421 VSS.n2270 VSS.n2269 179.448
R5422 VSS.n2270 VSS.n472 179.448
R5423 VSS.n2276 VSS.n472 179.448
R5424 VSS.n2277 VSS.n2276 179.448
R5425 VSS.n2278 VSS.n2277 179.448
R5426 VSS.n2278 VSS.n468 179.448
R5427 VSS.n2284 VSS.n468 179.448
R5428 VSS.n2285 VSS.n2284 179.448
R5429 VSS.n2286 VSS.n2285 179.448
R5430 VSS.n2286 VSS.n464 179.448
R5431 VSS.n2292 VSS.n464 179.448
R5432 VSS.n2293 VSS.n2292 179.448
R5433 VSS.n2294 VSS.n2293 179.448
R5434 VSS.n2294 VSS.n460 179.448
R5435 VSS.n2300 VSS.n460 179.448
R5436 VSS.n2301 VSS.n2300 179.381
R5437 VSS.n2302 VSS.n2301 179.363
R5438 VSS.n2302 VSS.n456 179.363
R5439 VSS.n2308 VSS.n456 179.363
R5440 VSS.n2309 VSS.n2308 179.363
R5441 VSS.n2310 VSS.n2309 179.363
R5442 VSS.n2310 VSS.n452 179.363
R5443 VSS.n2316 VSS.n452 179.363
R5444 VSS.n2317 VSS.n2316 179.363
R5445 VSS.n2318 VSS.n2317 179.363
R5446 VSS.n2318 VSS.n448 179.363
R5447 VSS.n2324 VSS.n448 179.363
R5448 VSS.n2325 VSS.n2324 179.363
R5449 VSS.n2326 VSS.n2325 179.363
R5450 VSS.n2326 VSS.n444 179.363
R5451 VSS.n2332 VSS.n444 179.363
R5452 VSS.n2333 VSS.n2332 179.363
R5453 VSS.n2334 VSS.n2333 179.363
R5454 VSS.n2334 VSS.n440 179.363
R5455 VSS.n2340 VSS.n440 179.363
R5456 VSS.n2341 VSS.n2340 179.363
R5457 VSS.n2342 VSS.n2341 179.363
R5458 VSS.n2342 VSS.n436 179.363
R5459 VSS.n2348 VSS.n436 179.363
R5460 VSS.n2349 VSS.n2348 179.363
R5461 VSS.n2350 VSS.n2349 179.363
R5462 VSS.n2350 VSS.n432 179.363
R5463 VSS.n2356 VSS.n432 179.363
R5464 VSS.n2357 VSS.n2356 179.363
R5465 VSS.n2358 VSS.n2357 179.363
R5466 VSS.n2358 VSS.n428 179.363
R5467 VSS.n2364 VSS.n428 179.363
R5468 VSS.n2365 VSS.n2364 179.363
R5469 VSS.n2366 VSS.n2365 179.363
R5470 VSS.n2366 VSS.n424 179.363
R5471 VSS.n2375 VSS.n424 179.363
R5472 VSS.n2376 VSS.n2375 179.363
R5473 VSS.n2377 VSS.n2376 179.363
R5474 VSS.n2377 VSS.n409 179.363
R5475 VSS.n2401 VSS.n409 179.363
R5476 VSS.n2402 VSS.n2401 179.363
R5477 VSS.n2403 VSS.n2402 179.363
R5478 VSS.n2403 VSS.n405 179.363
R5479 VSS.n2409 VSS.n405 179.363
R5480 VSS.n2410 VSS.n2409 179.363
R5481 VSS.n2411 VSS.n2410 179.363
R5482 VSS.n2411 VSS.n401 179.363
R5483 VSS.n2417 VSS.n401 179.363
R5484 VSS.n2418 VSS.n2417 179.363
R5485 VSS.n2419 VSS.n2418 179.363
R5486 VSS.n2419 VSS.n397 179.363
R5487 VSS.n2425 VSS.n397 179.363
R5488 VSS.n2426 VSS.n2425 179.363
R5489 VSS.n2427 VSS.n2426 179.363
R5490 VSS.n2427 VSS.n393 179.363
R5491 VSS.n2035 VSS.t813 178.757
R5492 VSS.n371 VSS.t971 178.431
R5493 VSS.n2699 VSS.t967 178.431
R5494 VSS.t250 VSS.n257 178.167
R5495 VSS.t1115 VSS.n2588 178.167
R5496 VSS.n1131 VSS.n1106 176.779
R5497 VSS.n1977 VSS.n1976 176.779
R5498 VSS.n151 VSS.n150 176.779
R5499 VSS.n2880 VSS.n2851 176.779
R5500 VSS.n1897 VSS.n1896 176.779
R5501 VSS.n1841 VSS.n1820 176.779
R5502 VSS.t397 VSS.t620 176.522
R5503 VSS.t601 VSS.t388 176.522
R5504 VSS.t618 VSS.t1248 176.522
R5505 VSS.t332 VSS.t645 176.522
R5506 VSS.t208 VSS.t992 176.522
R5507 VSS.t1006 VSS.t574 176.522
R5508 VSS.t1278 VSS.t994 176.522
R5509 VSS.t1012 VSS.t1275 176.522
R5510 VSS.t636 VSS.t683 176.522
R5511 VSS.t363 VSS.t639 176.522
R5512 VSS.n1994 VSS.t1152 176.161
R5513 VSS.n2468 VSS.n336 176.119
R5514 VSS.n2486 VSS.n279 176.119
R5515 VSS.n2728 VSS.n2610 176.119
R5516 VSS.n2710 VSS.n2664 176.119
R5517 VSS.n1177 VSS.t174 175.911
R5518 VSS.n2568 VSS.t925 175.911
R5519 VSS.t398 VSS.n1385 175.405
R5520 VSS.n1354 VSS.t333 175.405
R5521 VSS.n2207 VSS.t573 175.405
R5522 VSS.n2067 VSS.t1277 175.405
R5523 VSS.n1413 VSS.t364 175.405
R5524 VSS.t509 VSS.n354 174.071
R5525 VSS.t259 VSS.n311 174.071
R5526 VSS.t115 VSS.n2639 174.071
R5527 VSS.t932 VSS.n2682 174.071
R5528 VSS.n1381 VSS.t158 170.679
R5529 VSS.n1355 VSS.t146 170.679
R5530 VSS.n1325 VSS.t478 170.679
R5531 VSS.n2131 VSS.t122 170.679
R5532 VSS.n2181 VSS.t111 170.679
R5533 VSS.n2070 VSS.t214 170.679
R5534 VSS.t176 VSS.n1936 170.679
R5535 VSS.n1994 VSS.t933 168.971
R5536 VSS.t64 VSS.n1992 167.826
R5537 VSS.n2543 VSS.t884 161.492
R5538 VSS.t780 VSS.n226 161.492
R5539 VSS.t879 VSS.n2567 161.492
R5540 VSS.t794 VSS.n2774 161.492
R5541 VSS.n2902 VSS.n6 158.471
R5542 VSS.n1958 VSS.n1957 158.471
R5543 VSS.n1878 VSS.n1877 158.471
R5544 VSS.n128 VSS.n127 158.471
R5545 VSS.n2861 VSS.n2855 158.471
R5546 VSS.n1859 VSS.n1858 158.471
R5547 VSS.t581 VSS.t507 155.022
R5548 VSS.t583 VSS.t505 155.022
R5549 VSS.t447 VSS.t351 155.022
R5550 VSS.t445 VSS.t349 155.022
R5551 VSS.t1245 VSS.t301 155.022
R5552 VSS.t1243 VSS.t303 155.022
R5553 VSS.t503 VSS.t1266 155.022
R5554 VSS.t501 VSS.t1268 155.022
R5555 VSS.t229 VSS.t225 155.022
R5556 VSS.t227 VSS.t223 155.022
R5557 VSS.t290 VSS.t265 155.022
R5558 VSS.t288 VSS.t263 155.022
R5559 VSS.n974 VSS.n561 154.909
R5560 VSS.n2541 VSS.t1048 149.957
R5561 VSS.n2576 VSS.t1043 149.957
R5562 VSS.n1395 VSS.t438 148.856
R5563 VSS.n2508 VSS.t707 146.01
R5564 VSS.n2753 VSS.t701 146.01
R5565 VSS.t705 VSS.n2034 145.918
R5566 VSS.t345 VSS.n2027 145.419
R5567 VSS.n1948 VSS.t827 144.732
R5568 VSS.n1116 VSS.t48 144.263
R5569 VSS.t849 VSS.n1128 144.263
R5570 VSS.n1964 VSS.t49 144.263
R5571 VSS.n1970 VSS.t555 144.263
R5572 VSS.n137 VSS.t1235 144.263
R5573 VSS.n143 VSS.t52 144.263
R5574 VSS.n2865 VSS.t86 144.263
R5575 VSS.t544 VSS.n2877 144.263
R5576 VSS.n1884 VSS.t906 144.263
R5577 VSS.n1890 VSS.t1098 144.263
R5578 VSS.n1816 VSS.t809 144.263
R5579 VSS.t858 VSS.n1817 144.263
R5580 VSS.n1137 VSS.t846 144.143
R5581 VSS.n1141 VSS.t85 144.143
R5582 VSS.n1983 VSS.t564 144.143
R5583 VSS.t25 VSS.n1988 144.143
R5584 VSS.n157 VSS.t84 144.143
R5585 VSS.t1234 VSS.n183 144.143
R5586 VSS.n2886 VSS.t545 144.143
R5587 VSS.n2890 VSS.t87 144.143
R5588 VSS.n1903 VSS.t1100 144.143
R5589 VSS.t894 VSS.n1909 144.143
R5590 VSS.t862 VSS.n1839 144.143
R5591 VSS.n1835 VSS.t951 144.143
R5592 VSS.n2434 VSS.n393 144.105
R5593 VSS.t587 VSS.n2902 142.356
R5594 VSS.t1201 VSS.n6 142.356
R5595 VSS.n1957 VSS.t538 142.356
R5596 VSS.n1958 VSS.t736 142.356
R5597 VSS.n1877 VSS.t656 142.356
R5598 VSS.n1878 VSS.t650 142.356
R5599 VSS.n128 VSS.t842 142.356
R5600 VSS.n127 VSS.t1144 142.356
R5601 VSS.n2855 VSS.t691 142.356
R5602 VSS.t833 VSS.n2861 142.356
R5603 VSS.n1859 VSS.t1150 142.356
R5604 VSS.n1858 VSS.t1118 142.356
R5605 VSS.t48 VSS.t852 138.82
R5606 VSS.t844 VSS.t24 138.82
R5607 VSS.t848 VSS.t15 138.82
R5608 VSS.t41 VSS.t849 138.82
R5609 VSS.t562 VSS.t49 138.82
R5610 VSS.t565 VSS.t47 138.82
R5611 VSS.t554 VSS.t6 138.82
R5612 VSS.t555 VSS.t73 138.82
R5613 VSS.t28 VSS.t1235 138.82
R5614 VSS.t99 VSS.t1240 138.82
R5615 VSS.t70 VSS.t1232 138.82
R5616 VSS.t52 VSS.t1241 138.82
R5617 VSS.t86 VSS.t551 138.82
R5618 VSS.t548 VSS.t40 138.82
R5619 VSS.t541 VSS.t22 138.82
R5620 VSS.t77 VSS.t544 138.82
R5621 VSS.t1096 VSS.t906 138.82
R5622 VSS.t1103 VSS.t892 138.82
R5623 VSS.t1105 VSS.t901 138.82
R5624 VSS.t1098 VSS.t907 138.82
R5625 VSS.t809 VSS.t863 138.82
R5626 VSS.t866 VSS.t948 138.82
R5627 VSS.t869 VSS.t945 138.82
R5628 VSS.t954 VSS.t858 138.82
R5629 VSS.t88 VSS.t846 138.703
R5630 VSS.t45 VSS.t850 138.703
R5631 VSS.t27 VSS.t854 138.703
R5632 VSS.t85 VSS.t856 138.703
R5633 VSS.t34 VSS.t564 138.703
R5634 VSS.t0 VSS.t553 138.703
R5635 VSS.t59 VSS.t556 138.703
R5636 VSS.t559 VSS.t25 138.703
R5637 VSS.t1230 VSS.t84 138.703
R5638 VSS.t1236 VSS.t36 138.703
R5639 VSS.t1239 VSS.t96 138.703
R5640 VSS.t75 VSS.t1234 138.703
R5641 VSS.t90 VSS.t545 138.703
R5642 VSS.t37 VSS.t1106 138.703
R5643 VSS.t101 VSS.t542 138.703
R5644 VSS.t87 VSS.t546 138.703
R5645 VSS.t895 VSS.t1100 138.703
R5646 VSS.t899 VSS.t1101 138.703
R5647 VSS.t909 VSS.t1092 138.703
R5648 VSS.t1094 VSS.t894 138.703
R5649 VSS.t949 VSS.t862 138.703
R5650 VSS.t865 VSS.t807 138.703
R5651 VSS.t870 VSS.t947 138.703
R5652 VSS.t859 VSS.t951 138.703
R5653 VSS.t792 VSS.t1041 138.422
R5654 VSS.t1055 VSS.t784 138.422
R5655 VSS.n372 VSS.t964 137.011
R5656 VSS.n2700 VSS.t957 137.011
R5657 VSS.t1203 VSS.t587 136.983
R5658 VSS.t585 VSS.t1201 136.983
R5659 VSS.t538 VSS.t733 136.983
R5660 VSS.t736 VSS.t536 136.983
R5661 VSS.t656 VSS.t648 136.983
R5662 VSS.t650 VSS.t658 136.983
R5663 VSS.t842 VSS.t1146 136.983
R5664 VSS.t1144 VSS.t840 136.983
R5665 VSS.t691 VSS.t829 136.983
R5666 VSS.t689 VSS.t833 136.983
R5667 VSS.t1150 VSS.t1116 136.983
R5668 VSS.t1148 VSS.t1118 136.983
R5669 VSS.n1183 VSS.n1182 136.084
R5670 VSS.n2507 VSS.t1162 135.581
R5671 VSS.n2752 VSS.t1157 135.581
R5672 VSS.n1177 VSS.t175 135.537
R5673 VSS.n2568 VSS.t802 135.537
R5674 VSS.t269 VSS.n2051 135.124
R5675 VSS.t430 VSS.t1053 133.35
R5676 VSS.t1247 VSS.t1057 133.35
R5677 VSS.t1252 VSS.t628 133.35
R5678 VSS.t425 VSS.t571 133.35
R5679 VSS.t1083 VSS.t888 133.35
R5680 VSS.t760 VSS.t1176 133.35
R5681 VSS.t669 VSS.t1171 133.35
R5682 VSS.t674 VSS.t182 133.35
R5683 VSS.t786 VSS.t415 133.35
R5684 VSS.t788 VSS.t207 133.35
R5685 VSS.t998 VSS.t206 133.35
R5686 VSS.t260 VSS.t130 133.35
R5687 VSS.t138 VSS.t466 133.35
R5688 VSS.t758 VSS.t679 133.35
R5689 VSS.t1132 VSS.t680 133.35
R5690 VSS.t1139 VSS.t320 133.35
R5691 VSS.t977 VSS.t267 133.35
R5692 VSS.t1015 VSS.t1274 133.35
R5693 VSS.t1017 VSS.t1273 133.35
R5694 VSS.t1021 VSS.t1087 133.35
R5695 VSS.t458 VSS.t1215 133.35
R5696 VSS.t687 VSS.t1227 133.35
R5697 VSS.t688 VSS.t614 133.35
R5698 VSS.t436 VSS.t528 133.35
R5699 VSS.t282 VSS.t526 133.35
R5700 VSS.t387 VSS.t610 133.35
R5701 VSS.t386 VSS.t1191 133.35
R5702 VSS.t401 VSS.t1195 133.35
R5703 VSS.n1809 VSS.t284 132.734
R5704 VSS.n1595 VSS.n1594 131.986
R5705 VSS.n1594 VSS.n1460 131.986
R5706 VSS.n1588 VSS.n1460 131.986
R5707 VSS.n1588 VSS.n1587 131.986
R5708 VSS.n1587 VSS.n1586 131.986
R5709 VSS.n1586 VSS.n1464 131.986
R5710 VSS.n1580 VSS.n1464 131.986
R5711 VSS.n1580 VSS.n1579 131.986
R5712 VSS.n1579 VSS.n1578 131.986
R5713 VSS.n1578 VSS.n1468 131.986
R5714 VSS.n1572 VSS.n1468 131.986
R5715 VSS.n1572 VSS.n1571 131.986
R5716 VSS.n1571 VSS.n1570 131.986
R5717 VSS.n1570 VSS.n1472 131.986
R5718 VSS.n1564 VSS.n1472 131.986
R5719 VSS.n1564 VSS.n1563 131.986
R5720 VSS.n1563 VSS.n1562 131.986
R5721 VSS.n1562 VSS.n1476 131.986
R5722 VSS.n1556 VSS.n1476 131.986
R5723 VSS.n1556 VSS.n1555 131.986
R5724 VSS.n1555 VSS.n1554 131.986
R5725 VSS.n1554 VSS.n1480 131.986
R5726 VSS.n1548 VSS.n1480 131.986
R5727 VSS.n1548 VSS.n1547 131.986
R5728 VSS.n1547 VSS.n1546 131.986
R5729 VSS.n1546 VSS.n1484 131.986
R5730 VSS.n1540 VSS.n1484 131.986
R5731 VSS.n1540 VSS.n1539 131.986
R5732 VSS.n1539 VSS.n1538 131.986
R5733 VSS.n1538 VSS.n1488 131.986
R5734 VSS.n1532 VSS.n1488 131.986
R5735 VSS.n1532 VSS.n1531 131.986
R5736 VSS.n1531 VSS.n1530 131.986
R5737 VSS.n1530 VSS.n1492 131.986
R5738 VSS.n1524 VSS.n1492 131.986
R5739 VSS.n1524 VSS.n1523 131.986
R5740 VSS.n1523 VSS.n1522 131.986
R5741 VSS.n1522 VSS.n1496 131.986
R5742 VSS.n1516 VSS.n1496 131.986
R5743 VSS.n1516 VSS.n1515 131.986
R5744 VSS.n1515 VSS.n1514 131.986
R5745 VSS.n1514 VSS.n1500 131.986
R5746 VSS.n1508 VSS.n1500 131.986
R5747 VSS.n1508 VSS.n1507 131.986
R5748 VSS.n1507 VSS.n1506 131.986
R5749 VSS.n1506 VSS.n567 131.986
R5750 VSS.n2025 VSS.n567 131.986
R5751 VSS.t493 VSS.t1258 130.901
R5752 VSS.n2039 VSS.n559 129.338
R5753 VSS.n2542 VSS.t780 129.061
R5754 VSS.n2775 VSS.t794 129.061
R5755 VSS.t507 VSS.n1106 127.825
R5756 VSS.n1977 VSS.t351 127.825
R5757 VSS.n151 VSS.t301 127.825
R5758 VSS.t1266 VSS.n2851 127.825
R5759 VSS.n1897 VSS.t225 127.825
R5760 VSS.t265 VSS.n1820 127.825
R5761 VSS.n1336 VSS.t104 127.457
R5762 VSS.n2192 VSS.t916 127.398
R5763 VSS.n2191 VSS.t318 127.398
R5764 VSS.n1913 VSS.t897 125.344
R5765 VSS.t1258 VSS.n2035 125.272
R5766 VSS.t1159 VSS.t696 125.15
R5767 VSS.t1155 VSS.t709 125.15
R5768 VSS.t771 VSS.n63 124.522
R5769 VSS.t94 VSS.n1154 123.9
R5770 VSS.n179 VSS.t68 123.719
R5771 VSS.n320 VSS.t825 122.543
R5772 VSS.t1024 VSS.n296 122.543
R5773 VSS.n266 VSS.t1128 122.543
R5774 VSS.n2597 VSS.t1124 122.543
R5775 VSS.n2648 VSS.t820 122.543
R5776 VSS.t1177 VSS.n2624 122.543
R5777 VSS.n1335 VSS.t434 118.618
R5778 VSS.n2040 VSS.t934 116.843
R5779 VSS.n1913 VSS.t904 116.391
R5780 VSS.t1023 VSS.n1870 115.641
R5781 VSS.n1181 VSS.n1088 115.35
R5782 VSS.n319 VSS.t1060 112.115
R5783 VSS.n2476 VSS.t1219 112.115
R5784 VSS.n2494 VSS.t1193 112.115
R5785 VSS.n2736 VSS.t1187 112.115
R5786 VSS.n2647 VSS.t1069 112.115
R5787 VSS.n2718 VSS.t1213 112.115
R5788 VSS.t661 VSS.t374 108.832
R5789 VSS.t12 VSS.t534 108.413
R5790 VSS.t79 VSS.t325 108.254
R5791 VSS.n2026 VSS.n566 108.046
R5792 VSS.n2522 VSS.n2521 104.442
R5793 VSS.n255 VSS.n233 104.442
R5794 VSS.n2767 VSS.n2766 104.442
R5795 VSS.n2586 VSS.n72 104.442
R5796 VSS.t904 VSS.n1067 102.962
R5797 VSS.n2026 VSS.n2025 97.0154
R5798 VSS.n1871 VSS.t1028 92.6735
R5799 VSS.n210 VSS.n103 92.0327
R5800 VSS.n1167 VSS.n1166 92.0327
R5801 VSS.n1346 VSS.t571 91.4843
R5802 VSS.n1286 VSS.t1083 91.4843
R5803 VSS.t130 VSS.n2140 91.4843
R5804 VSS.n2151 VSS.t138 91.4843
R5805 VSS.n2052 VSS.t977 91.4843
R5806 VSS.n1405 VSS.t528 91.4843
R5807 VSS.t526 VSS.n1391 91.4843
R5808 VSS.t172 VSS.t663 89.3971
R5809 VSS.t665 VSS.t173 89.3971
R5810 VSS.t1120 VSS.t1023 87.0325
R5811 VSS.t1122 VSS.t1120 87.0325
R5812 VSS.t1028 VSS.t1122 87.0325
R5813 VSS.t409 VSS.t292 85.3293
R5814 VSS.n1871 VSS.t1032 84.1879
R5815 VSS.n2521 VSS.t790 83.964
R5816 VSS.n2766 VSS.t782 83.964
R5817 VSS.n2830 VSS.t1142 83.7364
R5818 VSS.n1596 VSS.n1595 81.2223
R5819 VSS.n2543 VSS.t251 80.7458
R5820 VSS.n2567 VSS.t455 80.7458
R5821 VSS.n1386 VSS.t397 80.4405
R5822 VSS.n1341 VSS.t332 80.4405
R5823 VSS.t574 VSS.n2206 80.4405
R5824 VSS.n2058 VSS.t1278 80.4405
R5825 VSS.n1400 VSS.t363 80.4405
R5826 VSS.t952 VSS.n1831 77.1682
R5827 VSS.t667 VSS.n210 73.9872
R5828 VSS.n1167 VSS.t672 73.9872
R5829 VSS.n1831 VSS.t943 71.6562
R5830 VSS.n1347 VSS.t1250 71.3268
R5831 VSS.t1172 VSS.n1294 71.3268
R5832 VSS.t204 VSS.n2205 71.3268
R5833 VSS.t681 VSS.n2159 71.3268
R5834 VSS.n2059 VSS.t1271 71.3268
R5835 VSS.n1406 VSS.t685 71.3268
R5836 VSS.n1200 VSS.t384 71.3268
R5837 VSS.n256 VSS.n255 69.6287
R5838 VSS.n2587 VSS.n2586 69.6287
R5839 VSS.t174 VSS.t884 69.2108
R5840 VSS.t251 VSS.t886 69.2108
R5841 VSS.t925 VSS.t879 69.2108
R5842 VSS.t455 VSS.t882 69.2108
R5843 VSS.n1130 VSS.t583 67.9921
R5844 VSS.n1039 VSS.t445 67.9921
R5845 VSS.n114 VSS.t1243 67.9921
R5846 VSS.n2879 VSS.t501 67.9921
R5847 VSS.n1428 VSS.t227 67.9921
R5848 VSS.n1840 VSS.t288 67.9921
R5849 VSS.n337 VSS.n297 67.5808
R5850 VSS.n280 VSS.n267 67.5808
R5851 VSS.n2611 VSS.n2598 67.5808
R5852 VSS.n2665 VSS.n2625 67.5808
R5853 VSS.t620 VSS.t398 64.7994
R5854 VSS.t388 VSS.t595 64.7994
R5855 VSS.t367 VSS.t601 64.7994
R5856 VSS.t928 VSS.t618 64.7994
R5857 VSS.t1248 VSS.t629 64.7994
R5858 VSS.t645 VSS.t333 64.7994
R5859 VSS.t992 VSS.t314 64.7994
R5860 VSS.t999 VSS.t208 64.7994
R5861 VSS.t573 VSS.t1006 64.7994
R5862 VSS.t994 VSS.t1277 64.7994
R5863 VSS.t1275 VSS.t1009 64.7994
R5864 VSS.t186 VSS.t1012 64.7994
R5865 VSS.t361 VSS.t636 64.7994
R5866 VSS.t683 VSS.t642 64.7994
R5867 VSS.t639 VSS.t364 64.7994
R5868 VSS.n1296 VSS.n1295 62.5655
R5869 VSS.n2161 VSS.n2160 62.5655
R5870 VSS.n1347 VSS.t615 62.0234
R5871 VSS.n1294 VSS.t746 62.0234
R5872 VSS.n2205 VSS.t989 62.0234
R5873 VSS.n2159 VSS.t744 62.0234
R5874 VSS.n2059 VSS.t1016 62.0234
R5875 VSS.n1406 VSS.t644 62.0234
R5876 VSS.n1200 VSS.t612 62.0234
R5877 VSS.t173 VSS.n1088 60.5595
R5878 VSS.n1131 VSS.n1130 59.8331
R5879 VSS.n1976 VSS.n1039 59.8331
R5880 VSS.n150 VSS.n114 59.8331
R5881 VSS.n2880 VSS.n2879 59.8331
R5882 VSS.n1896 VSS.n1428 59.8331
R5883 VSS.n1841 VSS.n1840 59.8331
R5884 VSS.n1870 VSS.t518 58.4247
R5885 VSS.n1184 VSS.t485 57.1852
R5886 VSS.t160 VSS.n200 57.1015
R5887 VSS.n338 VSS.t1221 47.1019
R5888 VSS.n281 VSS.t1197 47.1019
R5889 VSS.n2612 VSS.t1189 47.1019
R5890 VSS.n2666 VSS.t1217 47.1019
R5891 VSS.t663 VSS.n1181 46.1407
R5892 VSS.t1152 VSS.t934 43.1421
R5893 VSS.t877 VSS.t256 43.1421
R5894 VSS.n2434 VSS.n2433 40.075
R5895 VSS.n2520 VSS.n233 38.9104
R5896 VSS.n2765 VSS.n72 38.9104
R5897 VSS.n2051 VSS.t813 38.004
R5898 VSS.t292 VSS.n1809 37.9249
R5899 VSS.t369 VSS.t295 36.8625
R5900 VSS.n2475 VSS.n297 36.8625
R5901 VSS.n338 VSS.n337 36.8625
R5902 VSS.n354 VSS.n336 36.8625
R5903 VSS.t310 VSS.t509 36.8625
R5904 VSS.t1253 VSS.t966 36.8625
R5905 VSS.t280 VSS.t164 36.8625
R5906 VSS.n2493 VSS.n267 36.8625
R5907 VSS.n281 VSS.n280 36.8625
R5908 VSS.n311 VSS.n279 36.8625
R5909 VSS.t194 VSS.t259 36.8625
R5910 VSS.t824 VSS.t1062 36.8625
R5911 VSS.t166 VSS.t472 36.8625
R5912 VSS.n2735 VSS.n2598 36.8625
R5913 VSS.n2612 VSS.n2611 36.8625
R5914 VSS.n2639 VSS.n2610 36.8625
R5915 VSS.t249 VSS.t115 36.8625
R5916 VSS.t817 VSS.t1059 36.8625
R5917 VSS.t378 VSS.t495 36.8625
R5918 VSS.n2717 VSS.n2625 36.8625
R5919 VSS.n2666 VSS.n2665 36.8625
R5920 VSS.n2682 VSS.n2664 36.8625
R5921 VSS.t492 VSS.t932 36.8625
R5922 VSS.t1260 VSS.t961 36.8625
R5923 VSS.t1032 VSS.n2 35.1396
R5924 VSS.n258 VSS.t250 34.8146
R5925 VSS.n2589 VSS.t1115 34.8146
R5926 VSS.n372 VSS.n371 28.677
R5927 VSS.n2700 VSS.n2699 28.677
R5928 VSS.n981 VSS.n980 27.6079
R5929 VSS.n562 VSS.t1073 26.5311
R5930 VSS.n1393 VSS.n1392 26.1752
R5931 VSS.n1154 VSS.t534 25.0188
R5932 VSS.t325 VSS.n179 24.9822
R5933 VSS.n610 VSS.n561 24.5404
R5934 VSS.n1155 VSS.t94 23.8275
R5935 VSS.n199 VSS.t68 23.7926
R5936 VSS.t825 VSS.t1071 23.4662
R5937 VSS.n320 VSS.n319 23.4662
R5938 VSS.t1060 VSS.t811 23.4662
R5939 VSS.t1211 VSS.t1024 23.4662
R5940 VSS.n2476 VSS.n296 23.4662
R5941 VSS.t1219 VSS.t1037 23.4662
R5942 VSS.t1128 VSS.t1185 23.4662
R5943 VSS.n2494 VSS.n266 23.4662
R5944 VSS.t1193 VSS.t1135 23.4662
R5945 VSS.t1124 VSS.t1199 23.4662
R5946 VSS.n2736 VSS.n2597 23.4662
R5947 VSS.t1187 VSS.t1130 23.4662
R5948 VSS.t820 VSS.t1067 23.4662
R5949 VSS.n2648 VSS.n2647 23.4662
R5950 VSS.t1069 VSS.t822 23.4662
R5951 VSS.t1223 VSS.t1177 23.4662
R5952 VSS.n2718 VSS.n2624 23.4662
R5953 VSS.t1213 VSS.t1179 23.4662
R5954 VSS.t792 VSS.n2541 23.0706
R5955 VSS.n2576 VSS.t784 23.0706
R5956 VSS.t374 VSS.n201 22.5772
R5957 VSS.n1183 VSS.t930 22.5687
R5958 VSS.n1296 VSS.t311 22.2219
R5959 VSS.n2161 VSS.t920 22.2219
R5960 VSS.t696 VSS.n2507 20.8589
R5961 VSS.t709 VSS.n2752 20.8589
R5962 VSS.n1911 VSS.n1910 19.026
R5963 VSS.n2469 VSS.t1221 18.4315
R5964 VSS.n2469 VSS.t1039 18.4315
R5965 VSS.t1039 VSS.n2468 18.4315
R5966 VSS.n2487 VSS.t1197 18.4315
R5967 VSS.n2487 VSS.t1126 18.4315
R5968 VSS.t1126 VSS.n2486 18.4315
R5969 VSS.t790 VSS.n2520 18.4315
R5970 VSS.n257 VSS.t1051 18.4315
R5971 VSS.t782 VSS.n2765 18.4315
R5972 VSS.n2588 VSS.t1045 18.4315
R5973 VSS.n2729 VSS.t1189 18.4315
R5974 VSS.n2729 VSS.t1137 18.4315
R5975 VSS.t1137 VSS.n2728 18.4315
R5976 VSS.n2711 VSS.t1217 18.4315
R5977 VSS.n2711 VSS.t1181 18.4315
R5978 VSS.t1181 VSS.n2710 18.4315
R5979 VSS.n1759 VSS.n1458 16.7834
R5980 VSS.n211 VSS.t667 16.2415
R5981 VSS.t672 VSS.n1096 16.2415
R5982 VSS.n2464 VSS.n2459 14.4905
R5983 VSS.n2453 VSS.n2452 14.384
R5984 VSS.t1051 VSS.n256 14.3357
R5985 VSS.t1045 VSS.n2587 14.3357
R5986 VSS.n915 VSS.n689 14.3087
R5987 VSS.n2446 VSS.n2445 13.7962
R5988 VSS.n2062 VSS.n2061 13.6668
R5989 VSS.n2129 VSS.n507 13.6367
R5990 VSS.n1265 VSS.n221 13.6318
R5991 VSS.n1920 VSS.n1916 13.6285
R5992 VSS.n1117 VSS.n1116 13.6102
R5993 VSS.n1128 VSS.n1107 13.6102
R5994 VSS.n1964 VSS.n1963 13.6102
R5995 VSS.n1970 VSS.n1968 13.6102
R5996 VSS.n137 VSS.n136 13.6102
R5997 VSS.n143 VSS.n141 13.6102
R5998 VSS.n2866 VSS.n2865 13.6102
R5999 VSS.n2877 VSS.n2852 13.6102
R6000 VSS.n1884 VSS.n1883 13.6102
R6001 VSS.n1890 VSS.n1888 13.6102
R6002 VSS.n1853 VSS.n1816 13.6102
R6003 VSS.n1852 VSS.n1817 13.6102
R6004 VSS.n1137 VSS.n1136 13.5988
R6005 VSS.n1141 VSS.n1140 13.5988
R6006 VSS.n1984 VSS.n1983 13.5988
R6007 VSS.n1988 VSS.n1036 13.5988
R6008 VSS.n158 VSS.n157 13.5988
R6009 VSS.n183 VSS.n111 13.5988
R6010 VSS.n2886 VSS.n2885 13.5988
R6011 VSS.n2890 VSS.n2889 13.5988
R6012 VSS.n1904 VSS.n1903 13.5988
R6013 VSS.n1909 VSS.n1425 13.5988
R6014 VSS.n1839 VSS.n1823 13.5988
R6015 VSS.n1836 VSS.n1835 13.5988
R6016 VSS.n2211 VSS.n2210 13.5448
R6017 VSS.n1205 VSS.n547 13.5005
R6018 VSS.n2445 VSS.n2444 13.5005
R6019 VSS.n2064 VSS.n2063 13.5005
R6020 VSS.n1019 VSS.n1018 13.4554
R6021 VSS.n2033 VSS.n563 13.3493
R6022 VSS.n2217 VSS.n2216 13.0165
R6023 VSS.n1804 VSS.n1803 12.9534
R6024 VSS.n191 VSS.n190 12.8678
R6025 VSS.n94 VSS.n93 12.8678
R6026 VSS.n1090 VSS.n1089 12.8678
R6027 VSS.n1094 VSS.n1093 12.8678
R6028 VSS.n1030 VSS.n1029 12.8678
R6029 VSS.n2031 VSS.n2029 12.7598
R6030 VSS.n1146 VSS.t188 12.3882
R6031 VSS.n184 VSS.t1107 12.3613
R6032 VSS.n2045 VSS.n558 12.282
R6033 VSS.n2433 VSS.n62 12.0492
R6034 VSS.n2802 VSS.n2801 11.8868
R6035 VSS.n1832 VSS.n1829 11.7135
R6036 VSS.t1041 VSS.n226 11.5355
R6037 VSS.n2774 VSS.t1055 11.5355
R6038 VSS.n2814 VSS.n2813 11.3796
R6039 VSS.n1197 VSS.n1085 11.3589
R6040 VSS.n2209 VSS.n2208 11.2341
R6041 VSS.n1267 VSS.n1262 11.2341
R6042 VSS.n1384 VSS.n1383 11.2325
R6043 VSS.n1328 VSS.n1327 11.2325
R6044 VSS.n2184 VSS.n2183 11.2325
R6045 VSS.n2066 VSS.n533 11.2325
R6046 VSS.n1875 VSS.n1874 11.079
R6047 VSS.n1809 VSS.n1808 10.9898
R6048 VSS.n2405 VSS.n407 10.8241
R6049 VSS.n2079 VSS.n2078 10.7317
R6050 VSS.n2196 VSS.n2195 10.7317
R6051 VSS.n2188 VSS.n2187 10.7317
R6052 VSS.n1308 VSS.n1305 10.7317
R6053 VSS.n1344 VSS.n1343 10.7317
R6054 VSS.n1332 VSS.n1331 10.7317
R6055 VSS.n1194 VSS.n1193 10.7317
R6056 VSS.n1376 VSS.n1375 10.7317
R6057 VSS.n2074 VSS.n525 10.7317
R6058 VSS.n2168 VSS.n2167 10.7317
R6059 VSS.n2175 VSS.n2174 10.7317
R6060 VSS.n2123 VSS.n2122 10.7317
R6061 VSS.n2093 VSS.n512 10.7317
R6062 VSS.n1315 VSS.n1314 10.7317
R6063 VSS.n1363 VSS.n1362 10.7317
R6064 VSS.n1259 VSS.n1258 10.7317
R6065 VSS.n1226 VSS.n1208 10.7317
R6066 VSS.n1403 VSS.n1402 10.7317
R6067 VSS.n1929 VSS.n1928 10.7317
R6068 VSS.n1416 VSS.n1073 10.7317
R6069 VSS.n2048 VSS.n553 10.7317
R6070 VSS.n2177 VSS.n387 10.5272
R6071 VSS.n2442 VSS.n2441 10.5272
R6072 VSS.n2083 VSS.n2082 10.5272
R6073 VSS.n2107 VSS.n2106 10.5272
R6074 VSS.n2118 VSS.n515 10.5272
R6075 VSS.n2096 VSS.n2095 10.5272
R6076 VSS.n1323 VSS.n1322 10.5272
R6077 VSS.n1232 VSS.n1213 10.5272
R6078 VSS.n1360 VSS.n1244 10.5272
R6079 VSS.n1256 VSS.n1255 10.5272
R6080 VSS.n1230 VSS.n1229 10.5272
R6081 VSS.n1390 VSS.n1389 10.5272
R6082 VSS.n1399 VSS.n1083 10.5272
R6083 VSS.n1926 VSS.n1925 10.5272
R6084 VSS.n1941 VSS.n1940 10.5272
R6085 VSS.n2199 VSS.n2198 10.5272
R6086 VSS.n2152 VSS.n2145 10.5272
R6087 VSS.n1317 VSS.n380 10.5272
R6088 VSS.n1340 VSS.n1273 10.5272
R6089 VSS.n1287 VSS.n1280 10.5272
R6090 VSS.n2056 VSS.n2055 10.5272
R6091 VSS.n1633 VSS.n1627 10.5005
R6092 VSS.n1637 VSS.n1635 10.5005
R6093 VSS.n1641 VSS.n1625 10.5005
R6094 VSS.n1645 VSS.n1643 10.5005
R6095 VSS.n1649 VSS.n1623 10.5005
R6096 VSS.n1653 VSS.n1651 10.5005
R6097 VSS.n1657 VSS.n1621 10.5005
R6098 VSS.n1661 VSS.n1659 10.5005
R6099 VSS.n1665 VSS.n1619 10.5005
R6100 VSS.n1669 VSS.n1667 10.5005
R6101 VSS.n1673 VSS.n1617 10.5005
R6102 VSS.n1677 VSS.n1675 10.5005
R6103 VSS.n1681 VSS.n1615 10.5005
R6104 VSS.n1685 VSS.n1683 10.5005
R6105 VSS.n1689 VSS.n1613 10.5005
R6106 VSS.n1693 VSS.n1691 10.5005
R6107 VSS.n1697 VSS.n1611 10.5005
R6108 VSS.n1701 VSS.n1699 10.5005
R6109 VSS.n1705 VSS.n1609 10.5005
R6110 VSS.n1709 VSS.n1707 10.5005
R6111 VSS.n1713 VSS.n1607 10.5005
R6112 VSS.n1717 VSS.n1715 10.5005
R6113 VSS.n1721 VSS.n1605 10.5005
R6114 VSS.n1725 VSS.n1723 10.5005
R6115 VSS.n1729 VSS.n1603 10.5005
R6116 VSS.n1733 VSS.n1731 10.5005
R6117 VSS.n1737 VSS.n1601 10.5005
R6118 VSS.n1740 VSS.n1739 10.5005
R6119 VSS.n1747 VSS.n1745 10.5005
R6120 VSS.n1756 VSS.n1597 10.5005
R6121 VSS.n1758 VSS.n1459 10.5005
R6122 VSS.n1593 VSS.n1459 10.5005
R6123 VSS.n1593 VSS.n1461 10.5005
R6124 VSS.n1589 VSS.n1461 10.5005
R6125 VSS.n1589 VSS.n1463 10.5005
R6126 VSS.n1585 VSS.n1463 10.5005
R6127 VSS.n1585 VSS.n1465 10.5005
R6128 VSS.n1581 VSS.n1465 10.5005
R6129 VSS.n1581 VSS.n1467 10.5005
R6130 VSS.n1577 VSS.n1467 10.5005
R6131 VSS.n1577 VSS.n1469 10.5005
R6132 VSS.n1573 VSS.n1469 10.5005
R6133 VSS.n1573 VSS.n1471 10.5005
R6134 VSS.n1569 VSS.n1471 10.5005
R6135 VSS.n1569 VSS.n1473 10.5005
R6136 VSS.n1565 VSS.n1473 10.5005
R6137 VSS.n1565 VSS.n1475 10.5005
R6138 VSS.n1561 VSS.n1475 10.5005
R6139 VSS.n1561 VSS.n1477 10.5005
R6140 VSS.n1557 VSS.n1477 10.5005
R6141 VSS.n1557 VSS.n1479 10.5005
R6142 VSS.n1553 VSS.n1479 10.5005
R6143 VSS.n1553 VSS.n1481 10.5005
R6144 VSS.n1549 VSS.n1481 10.5005
R6145 VSS.n1549 VSS.n1483 10.5005
R6146 VSS.n1545 VSS.n1483 10.5005
R6147 VSS.n1545 VSS.n1485 10.5005
R6148 VSS.n1541 VSS.n1485 10.5005
R6149 VSS.n1541 VSS.n1487 10.5005
R6150 VSS.n1537 VSS.n1487 10.5005
R6151 VSS.n1537 VSS.n1489 10.5005
R6152 VSS.n1533 VSS.n1489 10.5005
R6153 VSS.n1533 VSS.n1491 10.5005
R6154 VSS.n1529 VSS.n1491 10.5005
R6155 VSS.n1529 VSS.n1493 10.5005
R6156 VSS.n1525 VSS.n1493 10.5005
R6157 VSS.n1525 VSS.n1495 10.5005
R6158 VSS.n1521 VSS.n1495 10.5005
R6159 VSS.n1521 VSS.n1497 10.5005
R6160 VSS.n1517 VSS.n1497 10.5005
R6161 VSS.n1517 VSS.n1499 10.5005
R6162 VSS.n1513 VSS.n1499 10.5005
R6163 VSS.n1513 VSS.n1501 10.5005
R6164 VSS.n1509 VSS.n1501 10.5005
R6165 VSS.n1509 VSS.n1503 10.5005
R6166 VSS.n1505 VSS.n1503 10.5005
R6167 VSS.n1505 VSS.n568 10.5005
R6168 VSS.n2024 VSS.n568 10.5005
R6169 VSS.n2024 VSS.n569 10.5005
R6170 VSS.n2020 VSS.n2018 10.5005
R6171 VSS.n2016 VSS.n572 10.5005
R6172 VSS.n2012 VSS.n2011 10.5005
R6173 VSS.n592 VSS.n588 10.5005
R6174 VSS.n593 VSS.n592 10.5005
R6175 VSS.n1017 VSS.n1016 10.5005
R6176 VSS.n1014 VSS.n595 10.5005
R6177 VSS.n1010 VSS.n1008 10.5005
R6178 VSS.n1006 VSS.n597 10.5005
R6179 VSS.n1002 VSS.n1000 10.5005
R6180 VSS.n1000 VSS.n999 10.5005
R6181 VSS.n999 VSS.n599 10.5005
R6182 VSS.n995 VSS.n599 10.5005
R6183 VSS.n995 VSS.n602 10.5005
R6184 VSS.n991 VSS.n602 10.5005
R6185 VSS.n991 VSS.n605 10.5005
R6186 VSS.n987 VSS.n605 10.5005
R6187 VSS.n987 VSS.n607 10.5005
R6188 VSS.n983 VSS.n607 10.5005
R6189 VSS.n983 VSS.n609 10.5005
R6190 VSS.n620 VSS.n617 10.5005
R6191 VSS.n624 VSS.n622 10.5005
R6192 VSS.n628 VSS.n614 10.5005
R6193 VSS.n632 VSS.n630 10.5005
R6194 VSS.n979 VSS.n611 10.5005
R6195 VSS.n979 VSS.n612 10.5005
R6196 VSS.n975 VSS.n612 10.5005
R6197 VSS.n975 VSS.n636 10.5005
R6198 VSS.n971 VSS.n636 10.5005
R6199 VSS.n971 VSS.n638 10.5005
R6200 VSS.n967 VSS.n638 10.5005
R6201 VSS.n967 VSS.n640 10.5005
R6202 VSS.n963 VSS.n640 10.5005
R6203 VSS.n963 VSS.n642 10.5005
R6204 VSS.n959 VSS.n642 10.5005
R6205 VSS.n959 VSS.n644 10.5005
R6206 VSS.n955 VSS.n644 10.5005
R6207 VSS.n955 VSS.n646 10.5005
R6208 VSS.n951 VSS.n646 10.5005
R6209 VSS.n951 VSS.n648 10.5005
R6210 VSS.n947 VSS.n648 10.5005
R6211 VSS.n947 VSS.n650 10.5005
R6212 VSS.n943 VSS.n650 10.5005
R6213 VSS.n943 VSS.n652 10.5005
R6214 VSS.n939 VSS.n652 10.5005
R6215 VSS.n939 VSS.n654 10.5005
R6216 VSS.n935 VSS.n654 10.5005
R6217 VSS.n935 VSS.n656 10.5005
R6218 VSS.n931 VSS.n656 10.5005
R6219 VSS.n931 VSS.n658 10.5005
R6220 VSS.n927 VSS.n658 10.5005
R6221 VSS.n927 VSS.n660 10.5005
R6222 VSS.n923 VSS.n660 10.5005
R6223 VSS.n923 VSS.n662 10.5005
R6224 VSS.n914 VSS.n662 10.5005
R6225 VSS.n914 VSS.n690 10.5005
R6226 VSS.n910 VSS.n690 10.5005
R6227 VSS.n910 VSS.n692 10.5005
R6228 VSS.n906 VSS.n692 10.5005
R6229 VSS.n906 VSS.n694 10.5005
R6230 VSS.n902 VSS.n694 10.5005
R6231 VSS.n902 VSS.n696 10.5005
R6232 VSS.n898 VSS.n696 10.5005
R6233 VSS.n898 VSS.n698 10.5005
R6234 VSS.n894 VSS.n698 10.5005
R6235 VSS.n894 VSS.n700 10.5005
R6236 VSS.n890 VSS.n700 10.5005
R6237 VSS.n890 VSS.n702 10.5005
R6238 VSS.n886 VSS.n702 10.5005
R6239 VSS.n886 VSS.n704 10.5005
R6240 VSS.n882 VSS.n704 10.5005
R6241 VSS.n882 VSS.n706 10.5005
R6242 VSS.n878 VSS.n706 10.5005
R6243 VSS.n878 VSS.n708 10.5005
R6244 VSS.n874 VSS.n708 10.5005
R6245 VSS.n874 VSS.n710 10.5005
R6246 VSS.n870 VSS.n710 10.5005
R6247 VSS.n870 VSS.n712 10.5005
R6248 VSS.n866 VSS.n712 10.5005
R6249 VSS.n866 VSS.n714 10.5005
R6250 VSS.n862 VSS.n714 10.5005
R6251 VSS.n862 VSS.n716 10.5005
R6252 VSS.n858 VSS.n716 10.5005
R6253 VSS.n858 VSS.n718 10.5005
R6254 VSS.n854 VSS.n718 10.5005
R6255 VSS.n854 VSS.n720 10.5005
R6256 VSS.n850 VSS.n720 10.5005
R6257 VSS.n850 VSS.n722 10.5005
R6258 VSS.n846 VSS.n722 10.5005
R6259 VSS.n846 VSS.n724 10.5005
R6260 VSS.n842 VSS.n724 10.5005
R6261 VSS.n842 VSS.n726 10.5005
R6262 VSS.n838 VSS.n726 10.5005
R6263 VSS.n838 VSS.n728 10.5005
R6264 VSS.n834 VSS.n728 10.5005
R6265 VSS.n834 VSS.n730 10.5005
R6266 VSS.n830 VSS.n730 10.5005
R6267 VSS.n830 VSS.n732 10.5005
R6268 VSS.n826 VSS.n732 10.5005
R6269 VSS.n826 VSS.n734 10.5005
R6270 VSS.n822 VSS.n734 10.5005
R6271 VSS.n822 VSS.n736 10.5005
R6272 VSS.n818 VSS.n736 10.5005
R6273 VSS.n818 VSS.n738 10.5005
R6274 VSS.n814 VSS.n738 10.5005
R6275 VSS.n814 VSS.n740 10.5005
R6276 VSS.n810 VSS.n740 10.5005
R6277 VSS.n810 VSS.n742 10.5005
R6278 VSS.n806 VSS.n742 10.5005
R6279 VSS.n806 VSS.n744 10.5005
R6280 VSS.n802 VSS.n744 10.5005
R6281 VSS.n802 VSS.n746 10.5005
R6282 VSS.n798 VSS.n746 10.5005
R6283 VSS.n798 VSS.n748 10.5005
R6284 VSS.n794 VSS.n748 10.5005
R6285 VSS.n794 VSS.n750 10.5005
R6286 VSS.n790 VSS.n750 10.5005
R6287 VSS.n790 VSS.n752 10.5005
R6288 VSS.n760 VSS.n752 10.5005
R6289 VSS.n780 VSS.n760 10.5005
R6290 VSS.n780 VSS.n761 10.5005
R6291 VSS.n776 VSS.n761 10.5005
R6292 VSS.n776 VSS.n501 10.5005
R6293 VSS.n2219 VSS.n501 10.5005
R6294 VSS.n2219 VSS.n499 10.5005
R6295 VSS.n2223 VSS.n499 10.5005
R6296 VSS.n2223 VSS.n497 10.5005
R6297 VSS.n2227 VSS.n497 10.5005
R6298 VSS.n2227 VSS.n495 10.5005
R6299 VSS.n2231 VSS.n495 10.5005
R6300 VSS.n2231 VSS.n493 10.5005
R6301 VSS.n2235 VSS.n493 10.5005
R6302 VSS.n2235 VSS.n491 10.5005
R6303 VSS.n2239 VSS.n491 10.5005
R6304 VSS.n2239 VSS.n489 10.5005
R6305 VSS.n2243 VSS.n489 10.5005
R6306 VSS.n2243 VSS.n487 10.5005
R6307 VSS.n2247 VSS.n487 10.5005
R6308 VSS.n2247 VSS.n485 10.5005
R6309 VSS.n2251 VSS.n485 10.5005
R6310 VSS.n2251 VSS.n483 10.5005
R6311 VSS.n2255 VSS.n483 10.5005
R6312 VSS.n2255 VSS.n481 10.5005
R6313 VSS.n2259 VSS.n481 10.5005
R6314 VSS.n2259 VSS.n479 10.5005
R6315 VSS.n2263 VSS.n479 10.5005
R6316 VSS.n2263 VSS.n477 10.5005
R6317 VSS.n2267 VSS.n477 10.5005
R6318 VSS.n2267 VSS.n475 10.5005
R6319 VSS.n2271 VSS.n475 10.5005
R6320 VSS.n2271 VSS.n473 10.5005
R6321 VSS.n2275 VSS.n473 10.5005
R6322 VSS.n2275 VSS.n471 10.5005
R6323 VSS.n2279 VSS.n471 10.5005
R6324 VSS.n2279 VSS.n469 10.5005
R6325 VSS.n2283 VSS.n469 10.5005
R6326 VSS.n2283 VSS.n467 10.5005
R6327 VSS.n2287 VSS.n467 10.5005
R6328 VSS.n2287 VSS.n465 10.5005
R6329 VSS.n2291 VSS.n465 10.5005
R6330 VSS.n2291 VSS.n463 10.5005
R6331 VSS.n2295 VSS.n463 10.5005
R6332 VSS.n2295 VSS.n461 10.5005
R6333 VSS.n2299 VSS.n461 10.5005
R6334 VSS.n2299 VSS.n459 10.5005
R6335 VSS.n2303 VSS.n459 10.5005
R6336 VSS.n2303 VSS.n457 10.5005
R6337 VSS.n2307 VSS.n457 10.5005
R6338 VSS.n2307 VSS.n455 10.5005
R6339 VSS.n2311 VSS.n455 10.5005
R6340 VSS.n2311 VSS.n453 10.5005
R6341 VSS.n2315 VSS.n453 10.5005
R6342 VSS.n2315 VSS.n451 10.5005
R6343 VSS.n2319 VSS.n451 10.5005
R6344 VSS.n2319 VSS.n449 10.5005
R6345 VSS.n2323 VSS.n449 10.5005
R6346 VSS.n2323 VSS.n447 10.5005
R6347 VSS.n2327 VSS.n447 10.5005
R6348 VSS.n2327 VSS.n445 10.5005
R6349 VSS.n2331 VSS.n445 10.5005
R6350 VSS.n2331 VSS.n443 10.5005
R6351 VSS.n2335 VSS.n443 10.5005
R6352 VSS.n2335 VSS.n441 10.5005
R6353 VSS.n2339 VSS.n441 10.5005
R6354 VSS.n2339 VSS.n439 10.5005
R6355 VSS.n2343 VSS.n439 10.5005
R6356 VSS.n2343 VSS.n437 10.5005
R6357 VSS.n2347 VSS.n437 10.5005
R6358 VSS.n2347 VSS.n435 10.5005
R6359 VSS.n2351 VSS.n435 10.5005
R6360 VSS.n2351 VSS.n433 10.5005
R6361 VSS.n2355 VSS.n433 10.5005
R6362 VSS.n2355 VSS.n431 10.5005
R6363 VSS.n2359 VSS.n431 10.5005
R6364 VSS.n2359 VSS.n429 10.5005
R6365 VSS.n2363 VSS.n429 10.5005
R6366 VSS.n2363 VSS.n427 10.5005
R6367 VSS.n2367 VSS.n427 10.5005
R6368 VSS.n2367 VSS.n425 10.5005
R6369 VSS.n2374 VSS.n425 10.5005
R6370 VSS.n2374 VSS.n423 10.5005
R6371 VSS.n2378 VSS.n423 10.5005
R6372 VSS.n2378 VSS.n410 10.5005
R6373 VSS.n2400 VSS.n410 10.5005
R6374 VSS.n2400 VSS.n408 10.5005
R6375 VSS.n2404 VSS.n408 10.5005
R6376 VSS.n2404 VSS.n406 10.5005
R6377 VSS.n2408 VSS.n406 10.5005
R6378 VSS.n2408 VSS.n404 10.5005
R6379 VSS.n2412 VSS.n404 10.5005
R6380 VSS.n2412 VSS.n402 10.5005
R6381 VSS.n2416 VSS.n402 10.5005
R6382 VSS.n2416 VSS.n400 10.5005
R6383 VSS.n2420 VSS.n400 10.5005
R6384 VSS.n2420 VSS.n398 10.5005
R6385 VSS.n2424 VSS.n398 10.5005
R6386 VSS.n2424 VSS.n396 10.5005
R6387 VSS.n2428 VSS.n396 10.5005
R6388 VSS.n2428 VSS.n394 10.5005
R6389 VSS.n2432 VSS.n394 10.5005
R6390 VSS.n2508 VSS.t1159 10.4297
R6391 VSS.n2753 VSS.t1155 10.4297
R6392 VSS.n1852 VSS 10.4038
R6393 VSS VSS.n2852 10.4038
R6394 VSS.n2889 VSS 10.4038
R6395 VSS VSS.n1107 10.4038
R6396 VSS.n1140 VSS 10.4038
R6397 VSS VSS.n1425 10.4038
R6398 VSS.n141 VSS 10.4038
R6399 VSS VSS.n111 10.4038
R6400 VSS VSS.n1036 10.4038
R6401 VSS.n1968 VSS 10.4038
R6402 VSS.n1888 VSS 10.4038
R6403 VSS VSS.n1836 10.4038
R6404 VSS VSS.n2121 10.4005
R6405 VSS VSS.n2094 10.4005
R6406 VSS VSS.n2197 10.4005
R6407 VSS VSS.n2186 10.4005
R6408 VSS.n2902 VSS.n2901 10.4005
R6409 VSS.n1110 VSS.n6 10.4005
R6410 VSS.n1116 VSS.n1115 10.4005
R6411 VSS.n1118 VSS.n1117 10.4005
R6412 VSS.n1128 VSS.n1127 10.4005
R6413 VSS.n1138 VSS.n1137 10.4005
R6414 VSS.n1122 VSS.n1106 10.4005
R6415 VSS.n1132 VSS.n1131 10.4005
R6416 VSS.n1136 VSS.n1135 10.4005
R6417 VSS.n1142 VSS.n1141 10.4005
R6418 VSS.n1318 VSS 10.4005
R6419 VSS VSS.n2455 10.4005
R6420 VSS.n2455 VSS 10.4005
R6421 VSS.n1324 VSS 10.4005
R6422 VSS VSS.n1361 10.4005
R6423 VSS VSS.n1342 10.4005
R6424 VSS VSS.n1330 10.4005
R6425 VSS VSS.n1257 10.4005
R6426 VSS VSS.n1401 10.4005
R6427 VSS VSS.n1927 10.4005
R6428 VSS VSS.n1939 10.4005
R6429 VSS VSS.n1387 10.4005
R6430 VSS.n1385 VSS 10.4005
R6431 VSS.n1382 VSS.n1381 10.4005
R6432 VSS.n1381 VSS.n1380 10.4005
R6433 VSS VSS.n1374 10.4005
R6434 VSS VSS.n1227 10.4005
R6435 VSS.n1231 VSS 10.4005
R6436 VSS VSS.n1231 10.4005
R6437 VSS.n1372 VSS 10.4005
R6438 VSS.n1367 VSS 10.4005
R6439 VSS.n1372 VSS 10.4005
R6440 VSS VSS.n1367 10.4005
R6441 VSS.n1365 VSS 10.4005
R6442 VSS.n1365 VSS 10.4005
R6443 VSS.n1355 VSS.n1266 10.4005
R6444 VSS.n1356 VSS.n1355 10.4005
R6445 VSS.n1354 VSS 10.4005
R6446 VSS.n1346 VSS 10.4005
R6447 VSS.n1335 VSS.n1334 10.4005
R6448 VSS.n1337 VSS.n1336 10.4005
R6449 VSS VSS.n1286 10.4005
R6450 VSS.n1329 VSS 10.4005
R6451 VSS.n1325 VSS.n1297 10.4005
R6452 VSS.n1326 VSS.n1325 10.4005
R6453 VSS.n1324 VSS 10.4005
R6454 VSS.n319 VSS.n318 10.4005
R6455 VSS.n2477 VSS.n2476 10.4005
R6456 VSS.n321 VSS.n320 10.4005
R6457 VSS.n329 VSS.n296 10.4005
R6458 VSS.n2495 VSS.n2494 10.4005
R6459 VSS.n2509 VSS.n2508 10.4005
R6460 VSS.n272 VSS.n266 10.4005
R6461 VSS.n2507 VSS.n2506 10.4005
R6462 VSS.n1159 VSS.n1088 10.4005
R6463 VSS.n1181 VSS.n1180 10.4005
R6464 VSS.n2544 VSS.n2543 10.4005
R6465 VSS.n2541 VSS.n2540 10.4005
R6466 VSS.n1178 VSS.n1177 10.4005
R6467 VSS.n2528 VSS.n226 10.4005
R6468 VSS.n373 VSS.n372 10.4005
R6469 VSS.n371 VSS.n370 10.4005
R6470 VSS.n2752 VSS.n2751 10.4005
R6471 VSS.n2737 VSS.n2736 10.4005
R6472 VSS.n2754 VSS.n2753 10.4005
R6473 VSS.n2603 VSS.n2597 10.4005
R6474 VSS.n2647 VSS.n2646 10.4005
R6475 VSS.n2719 VSS.n2718 10.4005
R6476 VSS.n2649 VSS.n2648 10.4005
R6477 VSS.n2657 VSS.n2624 10.4005
R6478 VSS VSS.n185 10.4005
R6479 VSS.n172 VSS.n171 10.4005
R6480 VSS.n2701 VSS.n2700 10.4005
R6481 VSS.n2699 VSS.n2698 10.4005
R6482 VSS.n2567 VSS.n2566 10.4005
R6483 VSS.n2774 VSS.n2773 10.4005
R6484 VSS.n2577 VSS.n2576 10.4005
R6485 VSS.n2569 VSS.n2568 10.4005
R6486 VSS.n189 VSS.n108 10.4005
R6487 VSS.n203 VSS.n202 10.4005
R6488 VSS VSS.n2104 10.4005
R6489 VSS VSS.n2080 10.4005
R6490 VSS.n2068 VSS 10.4005
R6491 VSS.n2068 VSS 10.4005
R6492 VSS.n2102 VSS 10.4005
R6493 VSS.n2101 VSS 10.4005
R6494 VSS.n2102 VSS 10.4005
R6495 VSS.n2101 VSS 10.4005
R6496 VSS.n2119 VSS 10.4005
R6497 VSS.n2119 VSS 10.4005
R6498 VSS.n2131 VSS.n2130 10.4005
R6499 VSS.n2131 VSS.n508 10.4005
R6500 VSS VSS.n2207 10.4005
R6501 VSS.n2140 VSS 10.4005
R6502 VSS.n2191 VSS.n2190 10.4005
R6503 VSS.n2193 VSS.n2192 10.4005
R6504 VSS VSS.n2151 10.4005
R6505 VSS.n2185 VSS 10.4005
R6506 VSS.n2181 VSS.n2162 10.4005
R6507 VSS.n2182 VSS.n2181 10.4005
R6508 VSS.n2163 VSS 10.4005
R6509 VSS.n2178 VSS 10.4005
R6510 VSS.n2180 VSS 10.4005
R6511 VSS.n2180 VSS 10.4005
R6512 VSS.n2436 VSS 10.4005
R6513 VSS VSS.n2436 10.4005
R6514 VSS VSS.n2028 10.4005
R6515 VSS.n1034 VSS.n1033 10.4005
R6516 VSS.n1957 VSS.n1956 10.4005
R6517 VSS.n1959 VSS.n1958 10.4005
R6518 VSS.n1965 VSS.n1964 10.4005
R6519 VSS.n1963 VSS.n1962 10.4005
R6520 VSS.n1971 VSS.n1970 10.4005
R6521 VSS.n1978 VSS.n1977 10.4005
R6522 VSS.n1983 VSS.n1982 10.4005
R6523 VSS.n1976 VSS.n1975 10.4005
R6524 VSS.n1985 VSS.n1984 10.4005
R6525 VSS.n1988 VSS.n1987 10.4005
R6526 VSS VSS.n1989 10.4005
R6527 VSS.n1992 VSS.n1991 10.4005
R6528 VSS VSS.n2040 10.4005
R6529 VSS.n2057 VSS 10.4005
R6530 VSS.n2070 VSS.n2069 10.4005
R6531 VSS.n2071 VSS.n2070 10.4005
R6532 VSS.n2067 VSS 10.4005
R6533 VSS VSS.n2052 10.4005
R6534 VSS.n2051 VSS.n2050 10.4005
R6535 VSS.n2035 VSS 10.4005
R6536 VSS.n1995 VSS.n1994 10.4005
R6537 VSS.n1063 VSS 10.4005
R6538 VSS VSS.n1058 10.4005
R6539 VSS.n1057 VSS 10.4005
R6540 VSS VSS.n1054 10.4005
R6541 VSS.n1951 VSS.n1950 10.4005
R6542 VSS.n1946 VSS 10.4005
R6543 VSS.n1946 VSS 10.4005
R6544 VSS.n1937 VSS 10.4005
R6545 VSS.n1937 VSS 10.4005
R6546 VSS.n1936 VSS.n1074 10.4005
R6547 VSS.n1936 VSS.n1935 10.4005
R6548 VSS.n1413 VSS 10.4005
R6549 VSS.n1396 VSS.n1395 10.4005
R6550 VSS.n1405 VSS 10.4005
R6551 VSS.n1191 VSS.n1086 10.4005
R6552 VSS.n1391 VSS 10.4005
R6553 VSS VSS.n1155 10.4005
R6554 VSS.n1145 VSS 10.4005
R6555 VSS.n1154 VSS.n1153 10.4005
R6556 VSS VSS.n1147 10.4005
R6557 VSS.n199 VSS 10.4005
R6558 VSS VSS.n180 10.4005
R6559 VSS.n179 VSS.n178 10.4005
R6560 VSS.n152 VSS.n151 10.4005
R6561 VSS.n157 VSS.n156 10.4005
R6562 VSS.n150 VSS.n149 10.4005
R6563 VSS.n159 VSS.n158 10.4005
R6564 VSS.n183 VSS.n182 10.4005
R6565 VSS.n138 VSS.n137 10.4005
R6566 VSS.n136 VSS.n135 10.4005
R6567 VSS.n144 VSS.n143 10.4005
R6568 VSS.n129 VSS.n128 10.4005
R6569 VSS.n127 VSS.n126 10.4005
R6570 VSS.n2894 VSS 10.4005
R6571 VSS.n2896 VSS.n2895 10.4005
R6572 VSS.n2871 VSS.n2851 10.4005
R6573 VSS.n2887 VSS.n2886 10.4005
R6574 VSS.n2881 VSS.n2880 10.4005
R6575 VSS.n2885 VSS.n2884 10.4005
R6576 VSS.n2891 VSS.n2890 10.4005
R6577 VSS.n2865 VSS.n2864 10.4005
R6578 VSS.n2867 VSS.n2866 10.4005
R6579 VSS.n2877 VSS.n2876 10.4005
R6580 VSS.n2856 VSS.n2855 10.4005
R6581 VSS.n2861 VSS.n2860 10.4005
R6582 VSS.n1911 VSS 10.4005
R6583 VSS.n1914 VSS.n1913 10.4005
R6584 VSS.n1898 VSS.n1897 10.4005
R6585 VSS.n1903 VSS.n1902 10.4005
R6586 VSS.n1896 VSS.n1895 10.4005
R6587 VSS.n1905 VSS.n1904 10.4005
R6588 VSS.n1909 VSS.n1908 10.4005
R6589 VSS.n1885 VSS.n1884 10.4005
R6590 VSS.n1883 VSS.n1882 10.4005
R6591 VSS.n1891 VSS.n1890 10.4005
R6592 VSS.n1879 VSS.n1878 10.4005
R6593 VSS.n1877 VSS.n1876 10.4005
R6594 VSS VSS.n1872 10.4005
R6595 VSS.n1860 VSS.n1859 10.4005
R6596 VSS.n1858 VSS.n1857 10.4005
R6597 VSS.n1849 VSS.n1816 10.4005
R6598 VSS.n1854 VSS.n1853 10.4005
R6599 VSS.n1846 VSS.n1817 10.4005
R6600 VSS.n1839 VSS.n1838 10.4005
R6601 VSS.n1824 VSS.n1820 10.4005
R6602 VSS.n1842 VSS.n1841 10.4005
R6603 VSS.n1823 VSS.n1822 10.4005
R6604 VSS.n1835 VSS.n1834 10.4005
R6605 VSS VSS.n1832 10.4005
R6606 VSS.n1831 VSS.n1830 10.4005
R6607 VSS.n2831 VSS.n2830 10.4005
R6608 VSS.n1870 VSS 10.4005
R6609 VSS VSS.n2906 10.4005
R6610 VSS.n1076 VSS.n10 10.295
R6611 VSS.n2202 VSS.n2201 10.1984
R6612 VSS.n2155 VSS.n2154 10.1984
R6613 VSS.n1352 VSS.n1351 10.1984
R6614 VSS.n1290 VSS.n1289 10.1984
R6615 VSS.n1411 VSS.n1410 10.1984
R6616 VSS.n1204 VSS.n1203 10.1984
R6617 VSS.n551 VSS.n535 10.1984
R6618 VSS.n2113 VSS.n2112 9.91668
R6619 VSS.n1370 VSS.n1369 9.82067
R6620 VSS.n1845 VSS.n1844 9.80927
R6621 VSS.n2875 VSS.n2874 9.80927
R6622 VSS.n1126 VSS.n1125 9.80927
R6623 VSS.n1973 VSS.n1972 9.80927
R6624 VSS.n1893 VSS.n1892 9.80927
R6625 VSS.n2030 VSS.n563 9.76794
R6626 VSS.n1856 VSS.n1855 9.65366
R6627 VSS.n2859 VSS.n2854 9.65366
R6628 VSS.n1112 VSS.n1111 9.65366
R6629 VSS.n1961 VSS.n1960 9.65366
R6630 VSS.n1881 VSS.n1880 9.65366
R6631 VSS.n2782 VSS.n61 9.38226
R6632 VSS.n2783 VSS.n2782 9.3812
R6633 VSS.n2465 VSS.n2464 9.36934
R6634 VSS.n1630 VSS.n1438 9.26515
R6635 VSS.n2561 VSS.n2560 9.0005
R6636 VSS.n2551 VSS.n2550 9.0005
R6637 VSS.n1999 VSS.n1998 9.0005
R6638 VSS.n2043 VSS.n2042 8.85306
R6639 VSS.n2898 VSS.n2849 8.84039
R6640 VSS.n2522 VSS.t305 8.19206
R6641 VSS.n2767 VSS.t926 8.19206
R6642 VSS.n1295 VSS.t740 7.99558
R6643 VSS.n2160 VSS.t775 7.99558
R6644 VSS.n213 VSS.n102 7.74518
R6645 VSS.n1175 VSS.n1097 7.74518
R6646 VSS.n259 VSS.n250 7.74518
R6647 VSS.n2488 VSS.n278 7.74518
R6648 VSS.n2485 VSS.n283 7.74518
R6649 VSS.n2470 VSS.n335 7.74518
R6650 VSS.n2467 VSS.n340 7.74518
R6651 VSS.n2519 VSS.n234 7.74518
R6652 VSS.n2712 VSS.n2663 7.74518
R6653 VSS.n2709 VSS.n2668 7.74518
R6654 VSS.n2730 VSS.n2609 7.74518
R6655 VSS.n2727 VSS.n2614 7.74518
R6656 VSS.n2764 VSS.n73 7.74518
R6657 VSS.n2590 VSS.n89 7.74518
R6658 VSS.n1998 VSS.n1997 7.49868
R6659 VSS.n2849 VSS.n9 7.29194
R6660 VSS.n1792 VSS.n1791 7.23784
R6661 VSS.n1152 VSS.n1151 7.12494
R6662 VSS.n2898 VSS.n2897 6.52095
R6663 VSS.n1874 VSS.n1873 6.2086
R6664 VSS.n1077 VSS.n1076 6.04619
R6665 VSS.n1437 VSS.n1435 6.00324
R6666 VSS.n177 VSS.n176 5.992
R6667 VSS.n1052 VSS.n1027 5.70095
R6668 VSS.n187 VSS.n186 5.43653
R6669 VSS VSS.t1027 5.43302
R6670 VSS VSS.t1119 5.39046
R6671 VSS VSS.t834 5.39046
R6672 VSS VSS.t737 5.39046
R6673 VSS.n1914 VSS.t905 5.38269
R6674 VSS.n1033 VSS.t731 5.38269
R6675 VSS VSS.t814 5.36235
R6676 VSS.n1950 VSS.t153 5.3339
R6677 VSS.n2162 VSS.t114 5.3339
R6678 VSS.n1297 VSS.t480 5.3339
R6679 VSS.n1935 VSS.t179 5.3339
R6680 VSS.n1191 VSS.t1280 5.3339
R6681 VSS.n1380 VSS.t366 5.3339
R6682 VSS.n2069 VSS.t217 5.3339
R6683 VSS VSS.t1153 5.31891
R6684 VSS.n146 VSS.n115 5.29395
R6685 VSS VSS.t191 5.2709
R6686 VSS.n2456 VSS.t774 5.247
R6687 VSS.n187 VSS.t326 5.24136
R6688 VSS.n2175 VSS.t471 5.23126
R6689 VSS.n2166 VSS.t180 5.23126
R6690 VSS.n2077 VSS.t272 5.23126
R6691 VSS.n2079 VSS.t155 5.23126
R6692 VSS.n2122 VSS.t694 5.23126
R6693 VSS.n2093 VSS.t377 5.23126
R6694 VSS.n516 VSS.t317 5.23126
R6695 VSS.n2196 VSS.t342 5.23126
R6696 VSS.n2187 VSS.t450 5.23126
R6697 VSS.n2143 VSS.t467 5.23126
R6698 VSS.n2137 VSS.t261 5.23126
R6699 VSS.n1149 VSS.t535 5.23126
R6700 VSS.n1315 VSS.t222 5.23126
R6701 VSS.n1298 VSS.t258 5.23126
R6702 VSS.n1305 VSS.t287 5.23126
R6703 VSS.n1362 VSS.t145 5.23126
R6704 VSS.n1343 VSS.t391 5.23126
R6705 VSS.n1331 VSS.t463 5.23126
R6706 VSS.n1278 VSS.t889 5.23126
R6707 VSS.n1345 VSS.t426 5.23126
R6708 VSS.n1258 VSS.t234 5.23126
R6709 VSS.n1245 VSS.t500 5.23126
R6710 VSS.n1364 VSS.t203 5.23126
R6711 VSS.n1226 VSS.t358 5.23126
R6712 VSS.n1217 VSS.t424 5.23126
R6713 VSS.n1402 VSS.t383 5.23126
R6714 VSS.n1928 VSS.t490 5.23126
R6715 VSS.n1417 VSS.t248 5.23126
R6716 VSS.n1073 VSS.t242 5.23126
R6717 VSS.n1415 VSS.t375 5.23126
R6718 VSS.n1404 VSS.t437 5.23126
R6719 VSS.n1187 VSS.t283 5.23126
R6720 VSS.n1194 VSS.t240 5.23126
R6721 VSS.n1211 VSS.t276 5.23126
R6722 VSS.n1375 VSS.t119 5.23126
R6723 VSS.n1313 VSS.t1270 5.23126
R6724 VSS.n174 VSS.t923 5.23126
R6725 VSS.n513 VSS.t1170 5.23126
R6726 VSS.n2073 VSS.t408 5.23126
R6727 VSS.n525 VSS.t110 5.23126
R6728 VSS.n2173 VSS.t133 5.23126
R6729 VSS.n2167 VSS.t516 5.23126
R6730 VSS.n553 VSS.t1282 5.23126
R6731 VSS.n555 VSS.t268 5.23126
R6732 VSS.n1873 VSS.t395 5.23126
R6733 VSS.n1810 VSS.t519 5.23126
R6734 VSS.n2042 VSS 5.21831
R6735 VSS.n2088 VSS.t980 5.21498
R6736 VSS.n1248 VSS.t631 5.21498
R6737 VSS.n1068 VSS.t625 5.21498
R6738 VSS.n2437 VSS.t743 5.21406
R6739 VSS.n2087 VSS.t1005 5.21406
R6740 VSS.n1219 VSS.t609 5.21406
R6741 VSS.n300 VSS.t1220 5.20602
R6742 VSS.n270 VSS.t1194 5.20602
R6743 VSS.n265 VSS.t1136 5.20602
R6744 VSS.n295 VSS.t1038 5.20602
R6745 VSS.n2527 VSS.t793 5.20602
R6746 VSS.n2539 VSS.t1049 5.20602
R6747 VSS.n1099 VSS.t666 5.20602
R6748 VSS.n2772 VSS.t785 5.20602
R6749 VSS.n2628 VSS.t1214 5.20602
R6750 VSS.n2601 VSS.t1188 5.20602
R6751 VSS.n2623 VSS.t1180 5.20602
R6752 VSS.n2738 VSS.t1131 5.20602
R6753 VSS.n92 VSS.t1044 5.20602
R6754 VSS.n204 VSS.t662 5.20602
R6755 VSS VSS.n340 5.2005
R6756 VSS.n354 VSS.n340 5.2005
R6757 VSS.n345 VSS.n344 5.2005
R6758 VSS.n344 VSS.n297 5.2005
R6759 VSS.n346 VSS.n339 5.2005
R6760 VSS.n339 VSS.n338 5.2005
R6761 VSS.n2467 VSS.n2466 5.2005
R6762 VSS.n2468 VSS.n2467 5.2005
R6763 VSS.n2471 VSS.n2470 5.2005
R6764 VSS.n2470 VSS.n2469 5.2005
R6765 VSS.n2472 VSS.n298 5.2005
R6766 VSS.n337 VSS.n298 5.2005
R6767 VSS.n2474 VSS.n2473 5.2005
R6768 VSS.n2475 VSS.n2474 5.2005
R6769 VSS.n335 VSS 5.2005
R6770 VSS.n336 VSS.n335 5.2005
R6771 VSS VSS.n283 5.2005
R6772 VSS.n311 VSS.n283 5.2005
R6773 VSS.n288 VSS.n287 5.2005
R6774 VSS.n287 VSS.n267 5.2005
R6775 VSS.n289 VSS.n282 5.2005
R6776 VSS.n282 VSS.n281 5.2005
R6777 VSS.n2485 VSS.n2484 5.2005
R6778 VSS.n2486 VSS.n2485 5.2005
R6779 VSS.n2489 VSS.n2488 5.2005
R6780 VSS.n2488 VSS.n2487 5.2005
R6781 VSS.n2490 VSS.n268 5.2005
R6782 VSS.n280 VSS.n268 5.2005
R6783 VSS.n2492 VSS.n2491 5.2005
R6784 VSS.n2493 VSS.n2492 5.2005
R6785 VSS.n278 VSS 5.2005
R6786 VSS.n279 VSS.n278 5.2005
R6787 VSS.n2519 VSS.n2518 5.2005
R6788 VSS.n2520 VSS.n2519 5.2005
R6789 VSS.n232 VSS.n231 5.2005
R6790 VSS.n2521 VSS.n232 5.2005
R6791 VSS.n2524 VSS.n2523 5.2005
R6792 VSS.n2523 VSS.n2522 5.2005
R6793 VSS VSS.n234 5.2005
R6794 VSS.n256 VSS.n234 5.2005
R6795 VSS VSS.n259 5.2005
R6796 VSS.n259 VSS.n258 5.2005
R6797 VSS.n252 VSS.n251 5.2005
R6798 VSS.n251 VSS.n233 5.2005
R6799 VSS.n254 VSS.n253 5.2005
R6800 VSS.n255 VSS.n254 5.2005
R6801 VSS.n250 VSS.n249 5.2005
R6802 VSS.n257 VSS.n250 5.2005
R6803 VSS.n1175 VSS 5.2005
R6804 VSS.n1176 VSS.n1175 5.2005
R6805 VSS.n1165 VSS.n1164 5.2005
R6806 VSS.n1166 VSS.n1165 5.2005
R6807 VSS.n1169 VSS.n1168 5.2005
R6808 VSS.n1168 VSS.n1167 5.2005
R6809 VSS.n1170 VSS.n1097 5.2005
R6810 VSS.n1097 VSS.n1096 5.2005
R6811 VSS VSS.n2590 5.2005
R6812 VSS.n2590 VSS.n2589 5.2005
R6813 VSS.n2583 VSS.n90 5.2005
R6814 VSS.n90 VSS.n72 5.2005
R6815 VSS.n2585 VSS.n2584 5.2005
R6816 VSS.n2586 VSS.n2585 5.2005
R6817 VSS.n89 VSS.n88 5.2005
R6818 VSS.n2588 VSS.n89 5.2005
R6819 VSS.n2764 VSS.n2763 5.2005
R6820 VSS.n2765 VSS.n2764 5.2005
R6821 VSS.n71 VSS.n70 5.2005
R6822 VSS.n2766 VSS.n71 5.2005
R6823 VSS.n2769 VSS.n2768 5.2005
R6824 VSS.n2768 VSS.n2767 5.2005
R6825 VSS VSS.n73 5.2005
R6826 VSS.n2587 VSS.n73 5.2005
R6827 VSS VSS.n2614 5.2005
R6828 VSS.n2639 VSS.n2614 5.2005
R6829 VSS.n2616 VSS.n2615 5.2005
R6830 VSS.n2615 VSS.n2598 5.2005
R6831 VSS.n2617 VSS.n2613 5.2005
R6832 VSS.n2613 VSS.n2612 5.2005
R6833 VSS.n2727 VSS.n2726 5.2005
R6834 VSS.n2728 VSS.n2727 5.2005
R6835 VSS.n2731 VSS.n2730 5.2005
R6836 VSS.n2730 VSS.n2729 5.2005
R6837 VSS.n2732 VSS.n2599 5.2005
R6838 VSS.n2611 VSS.n2599 5.2005
R6839 VSS.n2734 VSS.n2733 5.2005
R6840 VSS.n2735 VSS.n2734 5.2005
R6841 VSS.n2609 VSS 5.2005
R6842 VSS.n2610 VSS.n2609 5.2005
R6843 VSS VSS.n2668 5.2005
R6844 VSS.n2682 VSS.n2668 5.2005
R6845 VSS.n2673 VSS.n2672 5.2005
R6846 VSS.n2672 VSS.n2625 5.2005
R6847 VSS.n2674 VSS.n2667 5.2005
R6848 VSS.n2667 VSS.n2666 5.2005
R6849 VSS.n2709 VSS.n2708 5.2005
R6850 VSS.n2710 VSS.n2709 5.2005
R6851 VSS.n2713 VSS.n2712 5.2005
R6852 VSS.n2712 VSS.n2711 5.2005
R6853 VSS.n2714 VSS.n2626 5.2005
R6854 VSS.n2665 VSS.n2626 5.2005
R6855 VSS.n2716 VSS.n2715 5.2005
R6856 VSS.n2717 VSS.n2716 5.2005
R6857 VSS.n2663 VSS 5.2005
R6858 VSS.n2664 VSS.n2663 5.2005
R6859 VSS VSS.n213 5.2005
R6860 VSS.n213 VSS.n212 5.2005
R6861 VSS.n207 VSS.n104 5.2005
R6862 VSS.n104 VSS.n103 5.2005
R6863 VSS.n209 VSS.n208 5.2005
R6864 VSS.n210 VSS.n209 5.2005
R6865 VSS.n102 VSS.n101 5.2005
R6866 VSS.n211 VSS.n102 5.2005
R6867 VSS.n2033 VSS.n2032 5.2005
R6868 VSS.n2034 VSS.n2033 5.2005
R6869 VSS.n2031 VSS.n2030 5.2005
R6870 VSS.n2030 VSS.n559 5.2005
R6871 VSS VSS.n563 5.2005
R6872 VSS.n563 VSS.n562 5.2005
R6873 VSS.n2405 VSS.n2404 5.2005
R6874 VSS.n2404 VSS.n2403 5.2005
R6875 VSS.n2406 VSS.n406 5.2005
R6876 VSS.n406 VSS.n405 5.2005
R6877 VSS.n2408 VSS.n2407 5.2005
R6878 VSS.n2409 VSS.n2408 5.2005
R6879 VSS.n404 VSS.n403 5.2005
R6880 VSS.n2410 VSS.n404 5.2005
R6881 VSS.n2413 VSS.n2412 5.2005
R6882 VSS.n2412 VSS.n2411 5.2005
R6883 VSS.n2414 VSS.n402 5.2005
R6884 VSS.n402 VSS.n401 5.2005
R6885 VSS.n2416 VSS.n2415 5.2005
R6886 VSS.n2417 VSS.n2416 5.2005
R6887 VSS.n400 VSS.n399 5.2005
R6888 VSS.n2418 VSS.n400 5.2005
R6889 VSS.n2421 VSS.n2420 5.2005
R6890 VSS.n2420 VSS.n2419 5.2005
R6891 VSS.n2422 VSS.n398 5.2005
R6892 VSS.n398 VSS.n397 5.2005
R6893 VSS.n2424 VSS.n2423 5.2005
R6894 VSS.n2425 VSS.n2424 5.2005
R6895 VSS.n396 VSS.n395 5.2005
R6896 VSS.n2426 VSS.n396 5.2005
R6897 VSS.n2429 VSS.n2428 5.2005
R6898 VSS.n2428 VSS.n2427 5.2005
R6899 VSS.n2430 VSS.n394 5.2005
R6900 VSS.n394 VSS.n393 5.2005
R6901 VSS.n2432 VSS.n2431 5.2005
R6902 VSS.n62 VSS.n61 5.2005
R6903 VSS.n2372 VSS.n423 5.2005
R6904 VSS.n2376 VSS.n423 5.2005
R6905 VSS.n2379 VSS.n2378 5.2005
R6906 VSS.n2378 VSS.n2377 5.2005
R6907 VSS.n2382 VSS.n410 5.2005
R6908 VSS.n410 VSS.n409 5.2005
R6909 VSS.n2400 VSS.n2399 5.2005
R6910 VSS.n2401 VSS.n2400 5.2005
R6911 VSS.n408 VSS.n407 5.2005
R6912 VSS.n2402 VSS.n408 5.2005
R6913 VSS.n2217 VSS.n501 5.2005
R6914 VSS.n501 VSS.n500 5.2005
R6915 VSS.n2219 VSS.n2218 5.2005
R6916 VSS.n2220 VSS.n2219 5.2005
R6917 VSS.n499 VSS.n498 5.2005
R6918 VSS.n2221 VSS.n499 5.2005
R6919 VSS.n2224 VSS.n2223 5.2005
R6920 VSS.n2223 VSS.n2222 5.2005
R6921 VSS.n2225 VSS.n497 5.2005
R6922 VSS.n497 VSS.n496 5.2005
R6923 VSS.n2227 VSS.n2226 5.2005
R6924 VSS.n2228 VSS.n2227 5.2005
R6925 VSS.n495 VSS.n494 5.2005
R6926 VSS.n2229 VSS.n495 5.2005
R6927 VSS.n2232 VSS.n2231 5.2005
R6928 VSS.n2231 VSS.n2230 5.2005
R6929 VSS.n2233 VSS.n493 5.2005
R6930 VSS.n493 VSS.n492 5.2005
R6931 VSS.n2235 VSS.n2234 5.2005
R6932 VSS.n2236 VSS.n2235 5.2005
R6933 VSS.n491 VSS.n490 5.2005
R6934 VSS.n2237 VSS.n491 5.2005
R6935 VSS.n2240 VSS.n2239 5.2005
R6936 VSS.n2239 VSS.n2238 5.2005
R6937 VSS.n2241 VSS.n489 5.2005
R6938 VSS.n489 VSS.n488 5.2005
R6939 VSS.n2243 VSS.n2242 5.2005
R6940 VSS.n2244 VSS.n2243 5.2005
R6941 VSS.n487 VSS.n486 5.2005
R6942 VSS.n2245 VSS.n487 5.2005
R6943 VSS.n2248 VSS.n2247 5.2005
R6944 VSS.n2247 VSS.n2246 5.2005
R6945 VSS.n2249 VSS.n485 5.2005
R6946 VSS.n485 VSS.n484 5.2005
R6947 VSS.n2251 VSS.n2250 5.2005
R6948 VSS.n2252 VSS.n2251 5.2005
R6949 VSS.n483 VSS.n482 5.2005
R6950 VSS.n2253 VSS.n483 5.2005
R6951 VSS.n2256 VSS.n2255 5.2005
R6952 VSS.n2255 VSS.n2254 5.2005
R6953 VSS.n2257 VSS.n481 5.2005
R6954 VSS.n481 VSS.n480 5.2005
R6955 VSS.n2259 VSS.n2258 5.2005
R6956 VSS.n2260 VSS.n2259 5.2005
R6957 VSS.n479 VSS.n478 5.2005
R6958 VSS.n2261 VSS.n479 5.2005
R6959 VSS.n2264 VSS.n2263 5.2005
R6960 VSS.n2263 VSS.n2262 5.2005
R6961 VSS.n2265 VSS.n477 5.2005
R6962 VSS.n477 VSS.n476 5.2005
R6963 VSS.n2267 VSS.n2266 5.2005
R6964 VSS.n2268 VSS.n2267 5.2005
R6965 VSS.n475 VSS.n474 5.2005
R6966 VSS.n2269 VSS.n475 5.2005
R6967 VSS.n2272 VSS.n2271 5.2005
R6968 VSS.n2271 VSS.n2270 5.2005
R6969 VSS.n2273 VSS.n473 5.2005
R6970 VSS.n473 VSS.n472 5.2005
R6971 VSS.n2275 VSS.n2274 5.2005
R6972 VSS.n2276 VSS.n2275 5.2005
R6973 VSS.n471 VSS.n470 5.2005
R6974 VSS.n2277 VSS.n471 5.2005
R6975 VSS.n2280 VSS.n2279 5.2005
R6976 VSS.n2279 VSS.n2278 5.2005
R6977 VSS.n2281 VSS.n469 5.2005
R6978 VSS.n469 VSS.n468 5.2005
R6979 VSS.n2283 VSS.n2282 5.2005
R6980 VSS.n2284 VSS.n2283 5.2005
R6981 VSS.n467 VSS.n466 5.2005
R6982 VSS.n2285 VSS.n467 5.2005
R6983 VSS.n2288 VSS.n2287 5.2005
R6984 VSS.n2287 VSS.n2286 5.2005
R6985 VSS.n2289 VSS.n465 5.2005
R6986 VSS.n465 VSS.n464 5.2005
R6987 VSS.n2291 VSS.n2290 5.2005
R6988 VSS.n2292 VSS.n2291 5.2005
R6989 VSS.n463 VSS.n462 5.2005
R6990 VSS.n2293 VSS.n463 5.2005
R6991 VSS.n2296 VSS.n2295 5.2005
R6992 VSS.n2295 VSS.n2294 5.2005
R6993 VSS.n2297 VSS.n461 5.2005
R6994 VSS.n461 VSS.n460 5.2005
R6995 VSS.n2299 VSS.n2298 5.2005
R6996 VSS.n2300 VSS.n2299 5.2005
R6997 VSS.n459 VSS.n458 5.2005
R6998 VSS.n2301 VSS.n459 5.2005
R6999 VSS.n2304 VSS.n2303 5.2005
R7000 VSS.n2303 VSS.n2302 5.2005
R7001 VSS.n2305 VSS.n457 5.2005
R7002 VSS.n457 VSS.n456 5.2005
R7003 VSS.n2307 VSS.n2306 5.2005
R7004 VSS.n2308 VSS.n2307 5.2005
R7005 VSS.n455 VSS.n454 5.2005
R7006 VSS.n2309 VSS.n455 5.2005
R7007 VSS.n2312 VSS.n2311 5.2005
R7008 VSS.n2311 VSS.n2310 5.2005
R7009 VSS.n2313 VSS.n453 5.2005
R7010 VSS.n453 VSS.n452 5.2005
R7011 VSS.n2315 VSS.n2314 5.2005
R7012 VSS.n2316 VSS.n2315 5.2005
R7013 VSS.n451 VSS.n450 5.2005
R7014 VSS.n2317 VSS.n451 5.2005
R7015 VSS.n2320 VSS.n2319 5.2005
R7016 VSS.n2319 VSS.n2318 5.2005
R7017 VSS.n2321 VSS.n449 5.2005
R7018 VSS.n449 VSS.n448 5.2005
R7019 VSS.n2323 VSS.n2322 5.2005
R7020 VSS.n2324 VSS.n2323 5.2005
R7021 VSS.n447 VSS.n446 5.2005
R7022 VSS.n2325 VSS.n447 5.2005
R7023 VSS.n2328 VSS.n2327 5.2005
R7024 VSS.n2327 VSS.n2326 5.2005
R7025 VSS.n2329 VSS.n445 5.2005
R7026 VSS.n445 VSS.n444 5.2005
R7027 VSS.n2331 VSS.n2330 5.2005
R7028 VSS.n2332 VSS.n2331 5.2005
R7029 VSS.n443 VSS.n442 5.2005
R7030 VSS.n2333 VSS.n443 5.2005
R7031 VSS.n2336 VSS.n2335 5.2005
R7032 VSS.n2335 VSS.n2334 5.2005
R7033 VSS.n2337 VSS.n441 5.2005
R7034 VSS.n441 VSS.n440 5.2005
R7035 VSS.n2339 VSS.n2338 5.2005
R7036 VSS.n2340 VSS.n2339 5.2005
R7037 VSS.n439 VSS.n438 5.2005
R7038 VSS.n2341 VSS.n439 5.2005
R7039 VSS.n2344 VSS.n2343 5.2005
R7040 VSS.n2343 VSS.n2342 5.2005
R7041 VSS.n2345 VSS.n437 5.2005
R7042 VSS.n437 VSS.n436 5.2005
R7043 VSS.n2347 VSS.n2346 5.2005
R7044 VSS.n2348 VSS.n2347 5.2005
R7045 VSS.n435 VSS.n434 5.2005
R7046 VSS.n2349 VSS.n435 5.2005
R7047 VSS.n2352 VSS.n2351 5.2005
R7048 VSS.n2351 VSS.n2350 5.2005
R7049 VSS.n2353 VSS.n433 5.2005
R7050 VSS.n433 VSS.n432 5.2005
R7051 VSS.n2355 VSS.n2354 5.2005
R7052 VSS.n2356 VSS.n2355 5.2005
R7053 VSS.n431 VSS.n430 5.2005
R7054 VSS.n2357 VSS.n431 5.2005
R7055 VSS.n2360 VSS.n2359 5.2005
R7056 VSS.n2359 VSS.n2358 5.2005
R7057 VSS.n2361 VSS.n429 5.2005
R7058 VSS.n429 VSS.n428 5.2005
R7059 VSS.n2363 VSS.n2362 5.2005
R7060 VSS.n2364 VSS.n2363 5.2005
R7061 VSS.n427 VSS.n426 5.2005
R7062 VSS.n2365 VSS.n427 5.2005
R7063 VSS.n2368 VSS.n2367 5.2005
R7064 VSS.n2367 VSS.n2366 5.2005
R7065 VSS.n2369 VSS.n425 5.2005
R7066 VSS.n425 VSS.n424 5.2005
R7067 VSS.n2374 VSS.n2373 5.2005
R7068 VSS.n2375 VSS.n2374 5.2005
R7069 VSS.n788 VSS.n752 5.2005
R7070 VSS.n752 VSS.n751 5.2005
R7071 VSS.n760 VSS.n758 5.2005
R7072 VSS.n762 VSS.n760 5.2005
R7073 VSS.n781 VSS.n780 5.2005
R7074 VSS.n780 VSS.n779 5.2005
R7075 VSS.n761 VSS.n759 5.2005
R7076 VSS.n778 VSS.n761 5.2005
R7077 VSS.n776 VSS.n775 5.2005
R7078 VSS.n777 VSS.n776 5.2005
R7079 VSS.n690 VSS.n689 5.2005
R7080 VSS.n912 VSS.n690 5.2005
R7081 VSS.n910 VSS.n909 5.2005
R7082 VSS.n911 VSS.n910 5.2005
R7083 VSS.n908 VSS.n692 5.2005
R7084 VSS.n692 VSS.n691 5.2005
R7085 VSS.n907 VSS.n906 5.2005
R7086 VSS.n906 VSS.n905 5.2005
R7087 VSS.n694 VSS.n693 5.2005
R7088 VSS.n904 VSS.n694 5.2005
R7089 VSS.n902 VSS.n901 5.2005
R7090 VSS.n903 VSS.n902 5.2005
R7091 VSS.n900 VSS.n696 5.2005
R7092 VSS.n696 VSS.n695 5.2005
R7093 VSS.n899 VSS.n898 5.2005
R7094 VSS.n898 VSS.n897 5.2005
R7095 VSS.n698 VSS.n697 5.2005
R7096 VSS.n896 VSS.n698 5.2005
R7097 VSS.n894 VSS.n893 5.2005
R7098 VSS.n895 VSS.n894 5.2005
R7099 VSS.n892 VSS.n700 5.2005
R7100 VSS.n700 VSS.n699 5.2005
R7101 VSS.n891 VSS.n890 5.2005
R7102 VSS.n890 VSS.n889 5.2005
R7103 VSS.n702 VSS.n701 5.2005
R7104 VSS.n888 VSS.n702 5.2005
R7105 VSS.n886 VSS.n885 5.2005
R7106 VSS.n887 VSS.n886 5.2005
R7107 VSS.n884 VSS.n704 5.2005
R7108 VSS.n704 VSS.n703 5.2005
R7109 VSS.n883 VSS.n882 5.2005
R7110 VSS.n882 VSS.n881 5.2005
R7111 VSS.n706 VSS.n705 5.2005
R7112 VSS.n880 VSS.n706 5.2005
R7113 VSS.n878 VSS.n877 5.2005
R7114 VSS.n879 VSS.n878 5.2005
R7115 VSS.n876 VSS.n708 5.2005
R7116 VSS.n708 VSS.n707 5.2005
R7117 VSS.n875 VSS.n874 5.2005
R7118 VSS.n874 VSS.n873 5.2005
R7119 VSS.n710 VSS.n709 5.2005
R7120 VSS.n872 VSS.n710 5.2005
R7121 VSS.n870 VSS.n869 5.2005
R7122 VSS.n871 VSS.n870 5.2005
R7123 VSS.n868 VSS.n712 5.2005
R7124 VSS.n712 VSS.n711 5.2005
R7125 VSS.n867 VSS.n866 5.2005
R7126 VSS.n866 VSS.n865 5.2005
R7127 VSS.n714 VSS.n713 5.2005
R7128 VSS.n864 VSS.n714 5.2005
R7129 VSS.n862 VSS.n861 5.2005
R7130 VSS.n863 VSS.n862 5.2005
R7131 VSS.n860 VSS.n716 5.2005
R7132 VSS.n716 VSS.n715 5.2005
R7133 VSS.n859 VSS.n858 5.2005
R7134 VSS.n858 VSS.n857 5.2005
R7135 VSS.n718 VSS.n717 5.2005
R7136 VSS.n856 VSS.n718 5.2005
R7137 VSS.n854 VSS.n853 5.2005
R7138 VSS.n855 VSS.n854 5.2005
R7139 VSS.n852 VSS.n720 5.2005
R7140 VSS.n720 VSS.n719 5.2005
R7141 VSS.n851 VSS.n850 5.2005
R7142 VSS.n850 VSS.n849 5.2005
R7143 VSS.n722 VSS.n721 5.2005
R7144 VSS.n848 VSS.n722 5.2005
R7145 VSS.n846 VSS.n845 5.2005
R7146 VSS.n847 VSS.n846 5.2005
R7147 VSS.n844 VSS.n724 5.2005
R7148 VSS.n724 VSS.n723 5.2005
R7149 VSS.n843 VSS.n842 5.2005
R7150 VSS.n842 VSS.n841 5.2005
R7151 VSS.n726 VSS.n725 5.2005
R7152 VSS.n840 VSS.n726 5.2005
R7153 VSS.n838 VSS.n837 5.2005
R7154 VSS.n839 VSS.n838 5.2005
R7155 VSS.n836 VSS.n728 5.2005
R7156 VSS.n728 VSS.n727 5.2005
R7157 VSS.n835 VSS.n834 5.2005
R7158 VSS.n834 VSS.n833 5.2005
R7159 VSS.n730 VSS.n729 5.2005
R7160 VSS.n832 VSS.n730 5.2005
R7161 VSS.n830 VSS.n829 5.2005
R7162 VSS.n831 VSS.n830 5.2005
R7163 VSS.n828 VSS.n732 5.2005
R7164 VSS.n732 VSS.n731 5.2005
R7165 VSS.n827 VSS.n826 5.2005
R7166 VSS.n826 VSS.n825 5.2005
R7167 VSS.n734 VSS.n733 5.2005
R7168 VSS.n824 VSS.n734 5.2005
R7169 VSS.n822 VSS.n821 5.2005
R7170 VSS.n823 VSS.n822 5.2005
R7171 VSS.n820 VSS.n736 5.2005
R7172 VSS.n736 VSS.n735 5.2005
R7173 VSS.n819 VSS.n818 5.2005
R7174 VSS.n818 VSS.n817 5.2005
R7175 VSS.n738 VSS.n737 5.2005
R7176 VSS.n816 VSS.n738 5.2005
R7177 VSS.n814 VSS.n813 5.2005
R7178 VSS.n815 VSS.n814 5.2005
R7179 VSS.n812 VSS.n740 5.2005
R7180 VSS.n740 VSS.n739 5.2005
R7181 VSS.n811 VSS.n810 5.2005
R7182 VSS.n810 VSS.n809 5.2005
R7183 VSS.n742 VSS.n741 5.2005
R7184 VSS.n808 VSS.n742 5.2005
R7185 VSS.n806 VSS.n805 5.2005
R7186 VSS.n807 VSS.n806 5.2005
R7187 VSS.n804 VSS.n744 5.2005
R7188 VSS.n744 VSS.n743 5.2005
R7189 VSS.n803 VSS.n802 5.2005
R7190 VSS.n802 VSS.n801 5.2005
R7191 VSS.n746 VSS.n745 5.2005
R7192 VSS.n800 VSS.n746 5.2005
R7193 VSS.n798 VSS.n797 5.2005
R7194 VSS.n799 VSS.n798 5.2005
R7195 VSS.n796 VSS.n748 5.2005
R7196 VSS.n748 VSS.n747 5.2005
R7197 VSS.n795 VSS.n794 5.2005
R7198 VSS.n794 VSS.n793 5.2005
R7199 VSS.n750 VSS.n749 5.2005
R7200 VSS.n792 VSS.n750 5.2005
R7201 VSS.n790 VSS.n789 5.2005
R7202 VSS.n791 VSS.n790 5.2005
R7203 VSS.n928 VSS.n927 5.2005
R7204 VSS.n927 VSS.n926 5.2005
R7205 VSS.n677 VSS.n660 5.2005
R7206 VSS.n925 VSS.n660 5.2005
R7207 VSS.n923 VSS.n922 5.2005
R7208 VSS.n924 VSS.n923 5.2005
R7209 VSS.n688 VSS.n662 5.2005
R7210 VSS.n662 VSS.n661 5.2005
R7211 VSS.n915 VSS.n914 5.2005
R7212 VSS.n914 VSS.n913 5.2005
R7213 VSS.n1018 VSS.n1017 5.2005
R7214 VSS.n1016 VSS.n587 5.2005
R7215 VSS.n1014 VSS.n1013 5.2005
R7216 VSS.n1012 VSS.n595 5.2005
R7217 VSS.n1011 VSS.n1010 5.2005
R7218 VSS.n1008 VSS.n596 5.2005
R7219 VSS.n1006 VSS.n1005 5.2005
R7220 VSS.n1004 VSS.n597 5.2005
R7221 VSS.n1003 VSS.n1002 5.2005
R7222 VSS.n1000 VSS.n598 5.2005
R7223 VSS.n1000 VSS.n566 5.2005
R7224 VSS.n999 VSS.n600 5.2005
R7225 VSS.n999 VSS.n998 5.2005
R7226 VSS.n603 VSS.n599 5.2005
R7227 VSS.n997 VSS.n599 5.2005
R7228 VSS.n995 VSS.n994 5.2005
R7229 VSS.n996 VSS.n995 5.2005
R7230 VSS.n993 VSS.n602 5.2005
R7231 VSS.n602 VSS.n601 5.2005
R7232 VSS.n992 VSS.n991 5.2005
R7233 VSS.n991 VSS.n990 5.2005
R7234 VSS.n605 VSS.n604 5.2005
R7235 VSS.n989 VSS.n605 5.2005
R7236 VSS.n987 VSS.n986 5.2005
R7237 VSS.n988 VSS.n987 5.2005
R7238 VSS.n985 VSS.n607 5.2005
R7239 VSS.n607 VSS.n606 5.2005
R7240 VSS.n984 VSS.n983 5.2005
R7241 VSS.n983 VSS.n982 5.2005
R7242 VSS.n609 VSS.n608 5.2005
R7243 VSS.n618 VSS.n617 5.2005
R7244 VSS.n620 VSS.n619 5.2005
R7245 VSS.n622 VSS.n615 5.2005
R7246 VSS.n625 VSS.n624 5.2005
R7247 VSS.n626 VSS.n614 5.2005
R7248 VSS.n628 VSS.n627 5.2005
R7249 VSS.n630 VSS.n613 5.2005
R7250 VSS.n633 VSS.n632 5.2005
R7251 VSS.n634 VSS.n611 5.2005
R7252 VSS.n979 VSS.n978 5.2005
R7253 VSS.n980 VSS.n979 5.2005
R7254 VSS.n977 VSS.n612 5.2005
R7255 VSS.n612 VSS.n610 5.2005
R7256 VSS.n976 VSS.n975 5.2005
R7257 VSS.n975 VSS.n974 5.2005
R7258 VSS.n636 VSS.n635 5.2005
R7259 VSS.n973 VSS.n636 5.2005
R7260 VSS.n971 VSS.n970 5.2005
R7261 VSS.n972 VSS.n971 5.2005
R7262 VSS.n969 VSS.n638 5.2005
R7263 VSS.n638 VSS.n637 5.2005
R7264 VSS.n968 VSS.n967 5.2005
R7265 VSS.n967 VSS.n966 5.2005
R7266 VSS.n640 VSS.n639 5.2005
R7267 VSS.n965 VSS.n640 5.2005
R7268 VSS.n963 VSS.n962 5.2005
R7269 VSS.n964 VSS.n963 5.2005
R7270 VSS.n961 VSS.n642 5.2005
R7271 VSS.n642 VSS.n641 5.2005
R7272 VSS.n960 VSS.n959 5.2005
R7273 VSS.n959 VSS.n958 5.2005
R7274 VSS.n644 VSS.n643 5.2005
R7275 VSS.n957 VSS.n644 5.2005
R7276 VSS.n955 VSS.n954 5.2005
R7277 VSS.n956 VSS.n955 5.2005
R7278 VSS.n953 VSS.n646 5.2005
R7279 VSS.n646 VSS.n645 5.2005
R7280 VSS.n952 VSS.n951 5.2005
R7281 VSS.n951 VSS.n950 5.2005
R7282 VSS.n648 VSS.n647 5.2005
R7283 VSS.n949 VSS.n648 5.2005
R7284 VSS.n947 VSS.n946 5.2005
R7285 VSS.n948 VSS.n947 5.2005
R7286 VSS.n945 VSS.n650 5.2005
R7287 VSS.n650 VSS.n649 5.2005
R7288 VSS.n944 VSS.n943 5.2005
R7289 VSS.n943 VSS.n942 5.2005
R7290 VSS.n652 VSS.n651 5.2005
R7291 VSS.n941 VSS.n652 5.2005
R7292 VSS.n939 VSS.n938 5.2005
R7293 VSS.n940 VSS.n939 5.2005
R7294 VSS.n937 VSS.n654 5.2005
R7295 VSS.n654 VSS.n653 5.2005
R7296 VSS.n936 VSS.n935 5.2005
R7297 VSS.n935 VSS.n934 5.2005
R7298 VSS.n656 VSS.n655 5.2005
R7299 VSS.n933 VSS.n656 5.2005
R7300 VSS.n931 VSS.n930 5.2005
R7301 VSS.n932 VSS.n931 5.2005
R7302 VSS.n929 VSS.n658 5.2005
R7303 VSS.n658 VSS.n657 5.2005
R7304 VSS.n2013 VSS.n2012 5.2005
R7305 VSS.n2011 VSS.n2010 5.2005
R7306 VSS.n588 VSS.n577 5.2005
R7307 VSS.n592 VSS.n591 5.2005
R7308 VSS.n592 VSS.n566 5.2005
R7309 VSS.n593 VSS.n586 5.2005
R7310 VSS.n1459 VSS.n1458 5.2005
R7311 VSS.n1595 VSS.n1459 5.2005
R7312 VSS.n1593 VSS.n1592 5.2005
R7313 VSS.n1594 VSS.n1593 5.2005
R7314 VSS.n1591 VSS.n1461 5.2005
R7315 VSS.n1461 VSS.n1460 5.2005
R7316 VSS.n1590 VSS.n1589 5.2005
R7317 VSS.n1589 VSS.n1588 5.2005
R7318 VSS.n1463 VSS.n1462 5.2005
R7319 VSS.n1587 VSS.n1463 5.2005
R7320 VSS.n1585 VSS.n1584 5.2005
R7321 VSS.n1586 VSS.n1585 5.2005
R7322 VSS.n1583 VSS.n1465 5.2005
R7323 VSS.n1465 VSS.n1464 5.2005
R7324 VSS.n1582 VSS.n1581 5.2005
R7325 VSS.n1581 VSS.n1580 5.2005
R7326 VSS.n1467 VSS.n1466 5.2005
R7327 VSS.n1579 VSS.n1467 5.2005
R7328 VSS.n1577 VSS.n1576 5.2005
R7329 VSS.n1578 VSS.n1577 5.2005
R7330 VSS.n1575 VSS.n1469 5.2005
R7331 VSS.n1469 VSS.n1468 5.2005
R7332 VSS.n1574 VSS.n1573 5.2005
R7333 VSS.n1573 VSS.n1572 5.2005
R7334 VSS.n1471 VSS.n1470 5.2005
R7335 VSS.n1571 VSS.n1471 5.2005
R7336 VSS.n1569 VSS.n1568 5.2005
R7337 VSS.n1570 VSS.n1569 5.2005
R7338 VSS.n1567 VSS.n1473 5.2005
R7339 VSS.n1473 VSS.n1472 5.2005
R7340 VSS.n1566 VSS.n1565 5.2005
R7341 VSS.n1565 VSS.n1564 5.2005
R7342 VSS.n1475 VSS.n1474 5.2005
R7343 VSS.n1563 VSS.n1475 5.2005
R7344 VSS.n1561 VSS.n1560 5.2005
R7345 VSS.n1562 VSS.n1561 5.2005
R7346 VSS.n1559 VSS.n1477 5.2005
R7347 VSS.n1477 VSS.n1476 5.2005
R7348 VSS.n1558 VSS.n1557 5.2005
R7349 VSS.n1557 VSS.n1556 5.2005
R7350 VSS.n1479 VSS.n1478 5.2005
R7351 VSS.n1555 VSS.n1479 5.2005
R7352 VSS.n1553 VSS.n1552 5.2005
R7353 VSS.n1554 VSS.n1553 5.2005
R7354 VSS.n1551 VSS.n1481 5.2005
R7355 VSS.n1481 VSS.n1480 5.2005
R7356 VSS.n1550 VSS.n1549 5.2005
R7357 VSS.n1549 VSS.n1548 5.2005
R7358 VSS.n1483 VSS.n1482 5.2005
R7359 VSS.n1547 VSS.n1483 5.2005
R7360 VSS.n1545 VSS.n1544 5.2005
R7361 VSS.n1546 VSS.n1545 5.2005
R7362 VSS.n1543 VSS.n1485 5.2005
R7363 VSS.n1485 VSS.n1484 5.2005
R7364 VSS.n1542 VSS.n1541 5.2005
R7365 VSS.n1541 VSS.n1540 5.2005
R7366 VSS.n1487 VSS.n1486 5.2005
R7367 VSS.n1539 VSS.n1487 5.2005
R7368 VSS.n1537 VSS.n1536 5.2005
R7369 VSS.n1538 VSS.n1537 5.2005
R7370 VSS.n1535 VSS.n1489 5.2005
R7371 VSS.n1489 VSS.n1488 5.2005
R7372 VSS.n1534 VSS.n1533 5.2005
R7373 VSS.n1533 VSS.n1532 5.2005
R7374 VSS.n1491 VSS.n1490 5.2005
R7375 VSS.n1531 VSS.n1491 5.2005
R7376 VSS.n1529 VSS.n1528 5.2005
R7377 VSS.n1530 VSS.n1529 5.2005
R7378 VSS.n1527 VSS.n1493 5.2005
R7379 VSS.n1493 VSS.n1492 5.2005
R7380 VSS.n1526 VSS.n1525 5.2005
R7381 VSS.n1525 VSS.n1524 5.2005
R7382 VSS.n1495 VSS.n1494 5.2005
R7383 VSS.n1523 VSS.n1495 5.2005
R7384 VSS.n1521 VSS.n1520 5.2005
R7385 VSS.n1522 VSS.n1521 5.2005
R7386 VSS.n1519 VSS.n1497 5.2005
R7387 VSS.n1497 VSS.n1496 5.2005
R7388 VSS.n1518 VSS.n1517 5.2005
R7389 VSS.n1517 VSS.n1516 5.2005
R7390 VSS.n1499 VSS.n1498 5.2005
R7391 VSS.n1515 VSS.n1499 5.2005
R7392 VSS.n1513 VSS.n1512 5.2005
R7393 VSS.n1514 VSS.n1513 5.2005
R7394 VSS.n1511 VSS.n1501 5.2005
R7395 VSS.n1501 VSS.n1500 5.2005
R7396 VSS.n1510 VSS.n1509 5.2005
R7397 VSS.n1509 VSS.n1508 5.2005
R7398 VSS.n1503 VSS.n1502 5.2005
R7399 VSS.n1507 VSS.n1503 5.2005
R7400 VSS.n1505 VSS.n1504 5.2005
R7401 VSS.n1506 VSS.n1505 5.2005
R7402 VSS.n570 VSS.n568 5.2005
R7403 VSS.n568 VSS.n567 5.2005
R7404 VSS.n2024 VSS.n2023 5.2005
R7405 VSS.n2025 VSS.n2024 5.2005
R7406 VSS.n2022 VSS.n569 5.2005
R7407 VSS.n2021 VSS.n2020 5.2005
R7408 VSS.n2018 VSS.n571 5.2005
R7409 VSS.n2016 VSS.n2015 5.2005
R7410 VSS.n2014 VSS.n572 5.2005
R7411 VSS.n1745 VSS.n1744 5.2005
R7412 VSS.n1748 VSS.n1747 5.2005
R7413 VSS.n1752 VSS.n1597 5.2005
R7414 VSS.n1756 VSS.n1755 5.2005
R7415 VSS.n1759 VSS.n1758 5.2005
R7416 VSS.n1631 VSS.n1627 5.2005
R7417 VSS.n1633 VSS.n1632 5.2005
R7418 VSS.n1635 VSS.n1626 5.2005
R7419 VSS.n1638 VSS.n1637 5.2005
R7420 VSS.n1639 VSS.n1625 5.2005
R7421 VSS.n1641 VSS.n1640 5.2005
R7422 VSS.n1643 VSS.n1624 5.2005
R7423 VSS.n1646 VSS.n1645 5.2005
R7424 VSS.n1647 VSS.n1623 5.2005
R7425 VSS.n1649 VSS.n1648 5.2005
R7426 VSS.n1651 VSS.n1622 5.2005
R7427 VSS.n1654 VSS.n1653 5.2005
R7428 VSS.n1655 VSS.n1621 5.2005
R7429 VSS.n1657 VSS.n1656 5.2005
R7430 VSS.n1659 VSS.n1620 5.2005
R7431 VSS.n1662 VSS.n1661 5.2005
R7432 VSS.n1663 VSS.n1619 5.2005
R7433 VSS.n1665 VSS.n1664 5.2005
R7434 VSS.n1667 VSS.n1618 5.2005
R7435 VSS.n1670 VSS.n1669 5.2005
R7436 VSS.n1671 VSS.n1617 5.2005
R7437 VSS.n1673 VSS.n1672 5.2005
R7438 VSS.n1675 VSS.n1616 5.2005
R7439 VSS.n1678 VSS.n1677 5.2005
R7440 VSS.n1679 VSS.n1615 5.2005
R7441 VSS.n1681 VSS.n1680 5.2005
R7442 VSS.n1683 VSS.n1614 5.2005
R7443 VSS.n1686 VSS.n1685 5.2005
R7444 VSS.n1687 VSS.n1613 5.2005
R7445 VSS.n1689 VSS.n1688 5.2005
R7446 VSS.n1691 VSS.n1612 5.2005
R7447 VSS.n1694 VSS.n1693 5.2005
R7448 VSS.n1695 VSS.n1611 5.2005
R7449 VSS.n1697 VSS.n1696 5.2005
R7450 VSS.n1699 VSS.n1610 5.2005
R7451 VSS.n1702 VSS.n1701 5.2005
R7452 VSS.n1703 VSS.n1609 5.2005
R7453 VSS.n1705 VSS.n1704 5.2005
R7454 VSS.n1707 VSS.n1608 5.2005
R7455 VSS.n1710 VSS.n1709 5.2005
R7456 VSS.n1711 VSS.n1607 5.2005
R7457 VSS.n1713 VSS.n1712 5.2005
R7458 VSS.n1715 VSS.n1606 5.2005
R7459 VSS.n1718 VSS.n1717 5.2005
R7460 VSS.n1719 VSS.n1605 5.2005
R7461 VSS.n1721 VSS.n1720 5.2005
R7462 VSS.n1723 VSS.n1604 5.2005
R7463 VSS.n1726 VSS.n1725 5.2005
R7464 VSS.n1727 VSS.n1603 5.2005
R7465 VSS.n1729 VSS.n1728 5.2005
R7466 VSS.n1731 VSS.n1602 5.2005
R7467 VSS.n1734 VSS.n1733 5.2005
R7468 VSS.n1735 VSS.n1601 5.2005
R7469 VSS.n1737 VSS.n1736 5.2005
R7470 VSS.n1739 VSS.n1600 5.2005
R7471 VSS.n1741 VSS.n1740 5.2005
R7472 VSS.n1630 VSS.n1629 5.2005
R7473 VSS.n1076 VSS.n1075 5.18836
R7474 VSS.n1276 VSS.t254 5.18736
R7475 VSS.n147 VSS.n146 5.17894
R7476 VSS.n1052 VSS.t725 5.17491
R7477 VSS.n1875 VSS.t651 5.1725
R7478 VSS.n2900 VSS.t1202 5.16935
R7479 VSS.n2208 VSS.t993 5.1621
R7480 VSS.n2184 VSS.t776 5.1621
R7481 VSS.n1267 VSS.t619 5.1621
R7482 VSS.n1328 VSS.t741 5.1621
R7483 VSS.n1077 VSS.t637 5.1621
R7484 VSS.n1384 VSS.t602 5.1621
R7485 VSS.n2066 VSS.t1013 5.1621
R7486 VSS.n1265 VSS.t924 5.1539
R7487 VSS.n1843 VSS.t266 5.14713
R7488 VSS.n1819 VSS.t264 5.14713
R7489 VSS.n1827 VSS.t871 5.14713
R7490 VSS.n1833 VSS.t860 5.14713
R7491 VSS.n1828 VSS.t953 5.14713
R7492 VSS.n20 VSS.t944 5.14713
R7493 VSS.n1847 VSS.t946 5.14713
R7494 VSS.n1845 VSS.t955 5.14713
R7495 VSS.n1850 VSS.t867 5.14713
R7496 VSS.n1815 VSS.t864 5.14713
R7497 VSS.n1862 VSS.t1151 5.14713
R7498 VSS.n1856 VSS.t1149 5.14713
R7499 VSS.n1861 VSS.t1117 5.14713
R7500 VSS.n1429 VSS.t902 5.14713
R7501 VSS.n1892 VSS.t908 5.14713
R7502 VSS.n196 VSS.t676 5.14713
R7503 VSS.n97 VSS.t883 5.14713
R7504 VSS.n216 VSS.t880 5.14713
R7505 VSS.n1124 VSS.t508 5.14713
R7506 VSS.n1133 VSS.t506 5.14713
R7507 VSS.n1134 VSS.t855 5.14713
R7508 VSS.n1143 VSS.t857 5.14713
R7509 VSS.n1144 VSS.t13 5.14713
R7510 VSS.n1152 VSS.t95 5.14713
R7511 VSS.n2858 VSS.t692 5.14713
R7512 VSS.n2859 VSS.t690 5.14713
R7513 VSS.n2857 VSS.t830 5.14713
R7514 VSS.n2869 VSS.t23 5.14713
R7515 VSS.n2875 VSS.t78 5.14713
R7516 VSS.n2863 VSS.t549 5.14713
R7517 VSS.n2862 VSS.t552 5.14713
R7518 VSS.n2873 VSS.t1267 5.14713
R7519 VSS.n2882 VSS.t1269 5.14713
R7520 VSS.n2883 VSS.t543 5.14713
R7521 VSS.n2892 VSS.t547 5.14713
R7522 VSS.n2893 VSS.t82 5.14713
R7523 VSS.n2897 VSS.t21 5.14713
R7524 VSS.n2888 VSS.t38 5.14713
R7525 VSS.n2850 VSS.t91 5.14713
R7526 VSS.n2870 VSS.t502 5.14713
R7527 VSS.n2872 VSS.t504 5.14713
R7528 VSS.n1120 VSS.t16 5.14713
R7529 VSS.n1126 VSS.t42 5.14713
R7530 VSS.n1114 VSS.t845 5.14713
R7531 VSS.n1113 VSS.t853 5.14713
R7532 VSS.n1109 VSS.t588 5.14713
R7533 VSS.n1111 VSS.t586 5.14713
R7534 VSS.n7 VSS.t1204 5.14713
R7535 VSS.n1139 VSS.t46 5.14713
R7536 VSS.n1105 VSS.t89 5.14713
R7537 VSS.n1121 VSS.t584 5.14713
R7538 VSS.n1123 VSS.t582 5.14713
R7539 VSS.n1158 VSS.t664 5.14713
R7540 VSS.n1915 VSS.t898 5.14713
R7541 VSS.n1894 VSS.t226 5.14713
R7542 VSS.n1426 VSS.t224 5.14713
R7543 VSS.n1906 VSS.t1093 5.14713
R7544 VSS.n1907 VSS.t1095 5.14713
R7545 VSS.n1901 VSS.t900 5.14713
R7546 VSS.n1900 VSS.t896 5.14713
R7547 VSS.n1899 VSS.t228 5.14713
R7548 VSS.n1427 VSS.t230 5.14713
R7549 VSS.n375 VSS.t1257 5.14713
R7550 VSS.n351 VSS.t1255 5.14713
R7551 VSS.n307 VSS.t1072 5.14713
R7552 VSS.n308 VSS.t1061 5.14713
R7553 VSS.n361 VSS.t972 5.14713
R7554 VSS.n355 VSS.t965 5.14713
R7555 VSS.n330 VSS.t1212 5.14713
R7556 VSS.n273 VSS.t1186 5.14713
R7557 VSS.n2497 VSS.t1129 5.14713
R7558 VSS.n315 VSS.t812 5.14713
R7559 VSS.n312 VSS.t826 5.14713
R7560 VSS.n2479 VSS.t1025 5.14713
R7561 VSS.n240 VSS.t708 5.14713
R7562 VSS.n2510 VSS.t697 5.14713
R7563 VSS.n2530 VSS.t781 5.14713
R7564 VSS.n242 VSS.t1163 5.14713
R7565 VSS.n245 VSS.t1160 5.14713
R7566 VSS.n2535 VSS.t1042 5.14713
R7567 VSS.n2545 VSS.t887 5.14713
R7568 VSS.n1172 VSS.t885 5.14713
R7569 VSS.n79 VSS.t702 5.14713
R7570 VSS.n2755 VSS.t710 5.14713
R7571 VSS.n2571 VSS.t795 5.14713
R7572 VSS.n2635 VSS.t1068 5.14713
R7573 VSS.n2636 VSS.t1070 5.14713
R7574 VSS.n2689 VSS.t968 5.14713
R7575 VSS.n2683 VSS.t958 5.14713
R7576 VSS.n2658 VSS.t1224 5.14713
R7577 VSS.n2604 VSS.t1200 5.14713
R7578 VSS.n2721 VSS.t1178 5.14713
R7579 VSS.n2703 VSS.t1264 5.14713
R7580 VSS.n2679 VSS.t1262 5.14713
R7581 VSS.n2643 VSS.t823 5.14713
R7582 VSS.n2640 VSS.t821 5.14713
R7583 VSS.n2742 VSS.t1125 5.14713
R7584 VSS.n81 VSS.t1158 5.14713
R7585 VSS.n84 VSS.t1156 5.14713
R7586 VSS.n173 VSS.t1036 5.14713
R7587 VSS.n170 VSS.t1030 5.14713
R7588 VSS.n124 VSS.t843 5.14713
R7589 VSS.n121 VSS.t841 5.14713
R7590 VSS.n131 VSS.t1145 5.14713
R7591 VSS.n123 VSS.t1147 5.14713
R7592 VSS.n116 VSS.t1233 5.14713
R7593 VSS.n145 VSS.t1242 5.14713
R7594 VSS.n139 VSS.t100 5.14713
R7595 VSS.n118 VSS.t29 5.14713
R7596 VSS.n148 VSS.t302 5.14713
R7597 VSS.n112 VSS.t304 5.14713
R7598 VSS.n160 VSS.t97 5.14713
R7599 VSS.n181 VSS.t76 5.14713
R7600 VSS.n161 VSS.t80 5.14713
R7601 VSS.n177 VSS.t69 5.14713
R7602 VSS.n155 VSS.t1237 5.14713
R7603 VSS.n154 VSS.t1231 5.14713
R7604 VSS.n153 VSS.t1244 5.14713
R7605 VSS.n113 VSS.t1246 5.14713
R7606 VSS.n2578 VSS.t1056 5.14713
R7607 VSS.n1032 VSS.t739 5.14713
R7608 VSS.n1974 VSS.t352 5.14713
R7609 VSS.n1037 VSS.t350 5.14713
R7610 VSS.n1986 VSS.t557 5.14713
R7611 VSS.n1035 VSS.t560 5.14713
R7612 VSS.n1990 VSS.t93 5.14713
R7613 VSS.n1028 VSS.t65 5.14713
R7614 VSS.n1981 VSS.t1 5.14713
R7615 VSS.n1980 VSS.t35 5.14713
R7616 VSS.n1979 VSS.t446 5.14713
R7617 VSS.n1038 VSS.t448 5.14713
R7618 VSS.n1040 VSS.t7 5.14713
R7619 VSS.n1972 VSS.t74 5.14713
R7620 VSS.n1966 VSS.t566 5.14713
R7621 VSS.n1042 VSS.t563 5.14713
R7622 VSS.n1954 VSS.t539 5.14713
R7623 VSS.n1960 VSS.t537 5.14713
R7624 VSS.n1955 VSS.t734 5.14713
R7625 VSS.n1886 VSS.t1104 5.14713
R7626 VSS.n1431 VSS.t1097 5.14713
R7627 VSS.n1432 VSS.t657 5.14713
R7628 VSS.n1880 VSS.t659 5.14713
R7629 VSS.n1433 VSS.t649 5.14713
R7630 VSS.n1837 VSS.t808 5.14713
R7631 VSS.n1826 VSS.t950 5.14713
R7632 VSS.n1825 VSS.t289 5.14713
R7633 VSS.n1818 VSS.t291 5.14713
R7634 VSS.n2114 VSS.t991 5.1454
R7635 VSS.n1237 VSS.t617 5.1454
R7636 VSS.n1917 VSS.t635 5.1454
R7637 VSS.n1236 VSS.t605 5.14447
R7638 VSS.n2111 VSS.t1014 5.14447
R7639 VSS.n2041 VSS.t878 5.13735
R7640 VSS.n2044 VSS.t1259 5.13413
R7641 VSS.n2452 VSS.t770 5.13148
R7642 VSS.n2453 VSS.t772 5.12074
R7643 VSS.n2129 VSS.t313 5.08183
R7644 VSS.n2139 VSS.t919 5.07198
R7645 VSS.n2832 VSS.t452 5.07083
R7646 VSS.n2046 VSS.t494 5.07083
R7647 VSS.n533 VSS.t279 5.07083
R7648 VSS.n2141 VSS.t499 5.07083
R7649 VSS.n2209 VSS.t125 5.07083
R7650 VSS.n1275 VSS.t193 5.07083
R7651 VSS.n1262 VSS.t149 5.07083
R7652 VSS.n1075 VSS.t329 5.07083
R7653 VSS.n1085 VSS.t331 5.07083
R7654 VSS.n1383 VSS.t417 5.07083
R7655 VSS.n1327 VSS.t211 5.07083
R7656 VSS.n2183 VSS.t396 5.07083
R7657 VSS.n1805 VSS.t285 5.07083
R7658 VSS.n1044 VSS.t1114 5.05713
R7659 VSS.n1061 VSS.t721 5.05713
R7660 VSS.n1059 VSS.t797 5.05713
R7661 VSS.n1049 VSS.t713 5.05713
R7662 VSS.n1055 VSS.t580 5.05713
R7663 VSS.n125 VSS.n119 5.00971
R7664 VSS.n134 VSS.n133 4.9259
R7665 VSS.n557 VSS.t706 4.92017
R7666 VSS.n2900 VSS.n2899 4.7456
R7667 VSS.n2899 VSS.n8 4.71732
R7668 VSS.n2575 VSS.n2574 4.70151
R7669 VSS.n175 VSS.n174 4.66121
R7670 VSS.n1864 VSS.n1814 4.64694
R7671 VSS VSS.n2132 4.63333
R7672 VSS VSS.n2157 4.63333
R7673 VSS VSS.n1272 4.63333
R7674 VSS VSS.n1292 4.63333
R7675 VSS VSS.n1082 4.63333
R7676 VSS VSS.n1199 4.63333
R7677 VSS.n1921 VSS.n1920 4.63083
R7678 VSS.n1150 VSS.n1149 4.62479
R7679 VSS.n1920 VSS.n1919 4.62145
R7680 VSS.n2563 VSS.n97 4.61606
R7681 VSS.n376 VSS.n375 4.61606
R7682 VSS.n308 VSS.n301 4.61606
R7683 VSS.n367 VSS.n355 4.61606
R7684 VSS.n315 VSS.n293 4.61606
R7685 VSS.n2510 VSS.n239 4.61606
R7686 VSS.n2503 VSS.n242 4.61606
R7687 VSS.n2545 VSS.n225 4.61606
R7688 VSS.n2755 VSS.n78 4.61606
R7689 VSS.n2636 VSS.n2629 4.61606
R7690 VSS.n2695 VSS.n2683 4.61606
R7691 VSS.n2704 VSS.n2703 4.61606
R7692 VSS.n2643 VSS.n2621 4.61606
R7693 VSS.n2748 VSS.n81 4.61606
R7694 VSS.n192 VSS.t1090 4.613
R7695 VSS.n191 VSS.t1091 4.613
R7696 VSS.n95 VSS.t805 4.613
R7697 VSS.n94 VSS.t806 4.613
R7698 VSS.n1091 VSS.t839 4.613
R7699 VSS.n1090 VSS.t837 4.613
R7700 VSS.n1095 VSS.t1209 4.613
R7701 VSS.n1094 VSS.t1208 4.613
R7702 VSS.n1031 VSS.t941 4.613
R7703 VSS.n1030 VSS.t940 4.613
R7704 VSS.n2042 VSS.n2041 4.61061
R7705 VSS.n2534 VSS.n2533 4.60595
R7706 VSS.n673 VSS.n670 4.58492
R7707 VSS.n2387 VSS.n414 4.5725
R7708 VSS.n770 VSS.n504 4.56576
R7709 VSS.n133 VSS.n132 4.56421
R7710 VSS.n1768 VSS.n1449 4.55603
R7711 VSS.n2202 VSS.n2134 4.54133
R7712 VSS.n2155 VSS.n2149 4.54133
R7713 VSS.n1351 VSS.n1350 4.54133
R7714 VSS.n1290 VSS.n1284 4.54133
R7715 VSS.n1410 VSS.n1409 4.54133
R7716 VSS.n551 VSS.n550 4.54133
R7717 VSS.n1784 VSS.n1783 4.53674
R7718 VSS.n1769 VSS.n1768 4.52628
R7719 VSS.n538 VSS.n28 4.52406
R7720 VSS.n766 VSS.n754 4.51151
R7721 VSS.n1865 VSS.n1864 4.50944
R7722 VSS.n686 VSS.n685 4.50899
R7723 VSS.n420 VSS.n416 4.50877
R7724 VSS.n2800 VSS.n47 4.50386
R7725 VSS.n58 VSS.n56 4.50345
R7726 VSS.n1780 VSS.n1779 4.50176
R7727 VSS.n2552 VSS.n45 4.50176
R7728 VSS.n542 VSS.n35 4.50176
R7729 VSS.n585 VSS.n583 4.50176
R7730 VSS.n2838 VSS.n2837 4.50176
R7731 VSS.n1762 VSS.n1761 4.50176
R7732 VSS.n2001 VSS.n579 4.50139
R7733 VSS.n2002 VSS.n2001 4.50103
R7734 VSS.n2553 VSS.n38 4.50092
R7735 VSS.n1775 VSS.n1441 4.50089
R7736 VSS.n1864 VSS.n1863 4.5005
R7737 VSS.n1151 VSS.n1102 4.5005
R7738 VSS.n683 VSS.n665 4.5005
R7739 VSS.n918 VSS.n668 4.5005
R7740 VSS.n682 VSS.n679 4.5005
R7741 VSS.n674 VSS.n673 4.5005
R7742 VSS.n920 VSS.n666 4.5005
R7743 VSS.n687 VSS.n686 4.5005
R7744 VSS.n675 VSS.n672 4.5005
R7745 VSS.n919 VSS.n667 4.5005
R7746 VSS.n669 VSS.n668 4.5005
R7747 VSS.n682 VSS.n681 4.5005
R7748 VSS.n680 VSS.n666 4.5005
R7749 VSS.n540 VSS.n30 4.5005
R7750 VSS.n2816 VSS.n34 4.5005
R7751 VSS.n2822 VSS.n29 4.5005
R7752 VSS.n2824 VSS.n27 4.5005
R7753 VSS.n2818 VSS.n32 4.5005
R7754 VSS.n2823 VSS.n28 4.5005
R7755 VSS.n2817 VSS.n33 4.5005
R7756 VSS.n537 VSS.n27 4.5005
R7757 VSS.n541 VSS.n540 4.5005
R7758 VSS.n539 VSS.n29 4.5005
R7759 VSS.n544 VSS.n32 4.5005
R7760 VSS.n543 VSS.n33 4.5005
R7761 VSS.n684 VSS.n683 4.5005
R7762 VSS.n672 VSS.n536 4.5005
R7763 VSS.n671 VSS.n667 4.5005
R7764 VSS.n2793 VSS.n2792 4.5005
R7765 VSS.n2788 VSS.n57 4.5005
R7766 VSS.n54 VSS.n53 4.5005
R7767 VSS.n2794 VSS.n52 4.5005
R7768 VSS.n2798 VSS.n49 4.5005
R7769 VSS.n2787 VSS.n2786 4.5005
R7770 VSS.n2799 VSS.n48 4.5005
R7771 VSS.n2461 VSS.n50 4.5005
R7772 VSS.n2792 VSS.n2791 4.5005
R7773 VSS.n2789 VSS.n2788 4.5005
R7774 VSS.n2790 VSS.n54 4.5005
R7775 VSS.n55 VSS.n52 4.5005
R7776 VSS.n2460 VSS.n49 4.5005
R7777 VSS.n2462 VSS.n2461 4.5005
R7778 VSS.n374 VSS.n350 4.5005
R7779 VSS.n353 VSS.n352 4.5005
R7780 VSS.n369 VSS.n368 4.5005
R7781 VSS.n363 VSS.n362 4.5005
R7782 VSS.n310 VSS.n309 4.5005
R7783 VSS.n323 VSS.n322 4.5005
R7784 VSS.n317 VSS.n316 4.5005
R7785 VSS.n314 VSS.n313 4.5005
R7786 VSS.n2512 VSS.n2511 4.5005
R7787 VSS.n241 VSS.n238 4.5005
R7788 VSS.n2505 VSS.n2504 4.5005
R7789 VSS.n247 VSS.n246 4.5005
R7790 VSS.n2501 VSS.n2500 4.5005
R7791 VSS.n2547 VSS.n2546 4.5005
R7792 VSS.n1171 VSS.n223 4.5005
R7793 VSS.n2757 VSS.n2756 4.5005
R7794 VSS.n80 VSS.n77 4.5005
R7795 VSS.n2697 VSS.n2696 4.5005
R7796 VSS.n2691 VSS.n2690 4.5005
R7797 VSS.n2638 VSS.n2637 4.5005
R7798 VSS.n2651 VSS.n2650 4.5005
R7799 VSS.n2702 VSS.n2678 4.5005
R7800 VSS.n2681 VSS.n2680 4.5005
R7801 VSS.n2645 VSS.n2644 4.5005
R7802 VSS.n2642 VSS.n2641 4.5005
R7803 VSS.n2750 VSS.n2749 4.5005
R7804 VSS.n86 VSS.n85 4.5005
R7805 VSS.n2746 VSS.n2745 4.5005
R7806 VSS.n120 VSS.n119 4.5005
R7807 VSS.n176 VSS.n110 4.5005
R7808 VSS.n2565 VSS.n2564 4.5005
R7809 VSS.n218 VSS.n217 4.5005
R7810 VSS.n2554 VSS.n40 4.5005
R7811 VSS.n2804 VSS.n44 4.5005
R7812 VSS.n2810 VSS.n39 4.5005
R7813 VSS.n2812 VSS.n37 4.5005
R7814 VSS.n2806 VSS.n42 4.5005
R7815 VSS.n2811 VSS.n38 4.5005
R7816 VSS.n2805 VSS.n43 4.5005
R7817 VSS.n765 VSS.n757 4.5005
R7818 VSS.n504 VSS.n503 4.5005
R7819 VSS.n784 VSS.n756 4.5005
R7820 VSS.n786 VSS.n754 4.5005
R7821 VSS.n771 VSS.n764 4.5005
R7822 VSS.n2215 VSS.n2214 4.5005
R7823 VSS.n785 VSS.n755 4.5005
R7824 VSS.n773 VSS.n772 4.5005
R7825 VSS.n755 VSS.n506 4.5005
R7826 VSS.n767 VSS.n756 4.5005
R7827 VSS.n771 VSS.n770 4.5005
R7828 VSS.n768 VSS.n765 4.5005
R7829 VSS.n2214 VSS.n2213 4.5005
R7830 VSS.n772 VSS.n505 4.5005
R7831 VSS.n2555 VSS.n2554 4.5005
R7832 VSS.n2559 VSS.n39 4.5005
R7833 VSS.n2558 VSS.n37 4.5005
R7834 VSS.n2557 VSS.n42 4.5005
R7835 VSS.n2553 VSS.n43 4.5005
R7836 VSS.n421 VSS.n419 4.5005
R7837 VSS.n2397 VSS.n414 4.5005
R7838 VSS.n2391 VSS.n418 4.5005
R7839 VSS.n2370 VSS.n416 4.5005
R7840 VSS.n2386 VSS.n2384 4.5005
R7841 VSS.n2396 VSS.n2395 4.5005
R7842 VSS.n2392 VSS.n417 4.5005
R7843 VSS.n2385 VSS.n413 4.5005
R7844 VSS.n2391 VSS.n2390 4.5005
R7845 VSS.n2387 VSS.n2386 4.5005
R7846 VSS.n2388 VSS.n419 4.5005
R7847 VSS.n2395 VSS.n2394 4.5005
R7848 VSS.n2393 VSS.n2392 4.5005
R7849 VSS.n2385 VSS.n415 4.5005
R7850 VSS.n2007 VSS.n2006 4.5005
R7851 VSS.n1022 VSS.n1021 4.5005
R7852 VSS.n2008 VSS.n579 4.5005
R7853 VSS.n2002 VSS.n2000 4.5005
R7854 VSS.n582 VSS.n581 4.5005
R7855 VSS.n2003 VSS.n578 4.5005
R7856 VSS.n1023 VSS.n584 4.5005
R7857 VSS.n1025 VSS.n582 4.5005
R7858 VSS.n1024 VSS.n1023 4.5005
R7859 VSS.n2849 VSS.n2848 4.5005
R7860 VSS.n2006 VSS.n2005 4.5005
R7861 VSS.n2004 VSS.n2003 4.5005
R7862 VSS.n14 VSS.n12 4.5005
R7863 VSS.n1786 VSS.n1785 4.5005
R7864 VSS.n1782 VSS.n11 4.5005
R7865 VSS.n2845 VSS.n2844 4.5005
R7866 VSS.n15 VSS.n13 4.5005
R7867 VSS.n16 VSS.n14 4.5005
R7868 VSS.n2839 VSS.n2836 4.5005
R7869 VSS.n1788 VSS.n1786 4.5005
R7870 VSS.n1790 VSS.n1782 4.5005
R7871 VSS.n2844 VSS.n2843 4.5005
R7872 VSS.n1789 VSS.n1783 4.5005
R7873 VSS.n17 VSS.n15 4.5005
R7874 VSS.n1750 VSS.n1452 4.5005
R7875 VSS.n1763 VSS.n1456 4.5005
R7876 VSS.n1769 VSS.n1451 4.5005
R7877 VSS.n1742 VSS.n1449 4.5005
R7878 VSS.n1765 VSS.n1454 4.5005
R7879 VSS.n1770 VSS.n1450 4.5005
R7880 VSS.n1764 VSS.n1455 4.5005
R7881 VSS.n1766 VSS.n1765 4.5005
R7882 VSS.n1764 VSS.n1453 4.5005
R7883 VSS.n1452 VSS.n1448 4.5005
R7884 VSS.n1771 VSS.n1770 4.5005
R7885 VSS.n1777 VSS.n1776 4.5005
R7886 VSS.n1772 VSS.n1442 4.5005
R7887 VSS.n1773 VSS.n1440 4.5005
R7888 VSS.n1774 VSS.n1445 4.5005
R7889 VSS.n1775 VSS.n1446 4.5005
R7890 VSS.n1776 VSS.n1443 4.5005
R7891 VSS.n1794 VSS.n1447 4.5005
R7892 VSS.n1800 VSS.n1442 4.5005
R7893 VSS.n1802 VSS.n1440 4.5005
R7894 VSS.n1796 VSS.n1445 4.5005
R7895 VSS.n1801 VSS.n1441 4.5005
R7896 VSS.n1795 VSS.n1446 4.5005
R7897 VSS.n1800 VSS.n1799 4.5005
R7898 VSS.n1803 VSS.n1802 4.5005
R7899 VSS.n1797 VSS.n1796 4.5005
R7900 VSS.n1794 VSS.n1793 4.5005
R7901 VSS.n1798 VSS.n1443 4.5005
R7902 VSS.n1801 VSS.n1439 4.5005
R7903 VSS.n1792 VSS.n1780 4.5005
R7904 VSS.n1795 VSS.n1444 4.5005
R7905 VSS.n1788 VSS.n1787 4.5005
R7906 VSS.n1791 VSS.n1790 4.5005
R7907 VSS.n2843 VSS.n2842 4.5005
R7908 VSS.n2840 VSS.n2839 4.5005
R7909 VSS.n18 VSS.n16 4.5005
R7910 VSS.n1789 VSS.n1781 4.5005
R7911 VSS.n2838 VSS.n2835 4.5005
R7912 VSS.n2841 VSS.n17 4.5005
R7913 VSS.n2822 VSS.n2821 4.5005
R7914 VSS.n2825 VSS.n2824 4.5005
R7915 VSS.n2819 VSS.n2818 4.5005
R7916 VSS.n2816 VSS.n2815 4.5005
R7917 VSS.n2820 VSS.n30 4.5005
R7918 VSS.n2823 VSS.n26 4.5005
R7919 VSS.n2814 VSS.n35 4.5005
R7920 VSS.n2817 VSS.n31 4.5005
R7921 VSS.n2810 VSS.n2809 4.5005
R7922 VSS.n2813 VSS.n2812 4.5005
R7923 VSS.n2807 VSS.n2806 4.5005
R7924 VSS.n2804 VSS.n2803 4.5005
R7925 VSS.n2808 VSS.n40 4.5005
R7926 VSS.n2811 VSS.n36 4.5005
R7927 VSS.n2802 VSS.n45 4.5005
R7928 VSS.n2805 VSS.n41 4.5005
R7929 VSS.n2799 VSS.n46 4.5005
R7930 VSS.n59 VSS.n53 4.5005
R7931 VSS.n2795 VSS.n2794 4.5005
R7932 VSS.n2798 VSS.n2797 4.5005
R7933 VSS.n2801 VSS.n2800 4.5005
R7934 VSS.n2786 VSS.n2785 4.5005
R7935 VSS.n2784 VSS.n58 4.5005
R7936 VSS.n60 VSS.n57 4.5005
R7937 VSS.n2793 VSS.n51 4.5005
R7938 VSS.n2796 VSS.n50 4.5005
R7939 VSS.n2396 VSS.n412 4.5005
R7940 VSS.n2381 VSS.n421 4.5005
R7941 VSS.n2398 VSS.n2397 4.5005
R7942 VSS.n2380 VSS.n418 4.5005
R7943 VSS.n2371 VSS.n2370 4.5005
R7944 VSS.n2384 VSS.n2383 4.5005
R7945 VSS.n422 VSS.n417 4.5005
R7946 VSS.n413 VSS.n411 4.5005
R7947 VSS.n2216 VSS.n2215 4.5005
R7948 VSS.n782 VSS.n757 4.5005
R7949 VSS.n503 VSS.n502 4.5005
R7950 VSS.n784 VSS.n783 4.5005
R7951 VSS.n787 VSS.n786 4.5005
R7952 VSS.n764 VSS.n763 4.5005
R7953 VSS.n785 VSS.n753 4.5005
R7954 VSS.n774 VSS.n773 4.5005
R7955 VSS.n916 VSS.n687 4.5005
R7956 VSS.n665 VSS.n663 4.5005
R7957 VSS.n918 VSS.n917 4.5005
R7958 VSS.n679 VSS.n678 4.5005
R7959 VSS.n674 VSS.n659 4.5005
R7960 VSS.n921 VSS.n920 4.5005
R7961 VSS.n676 VSS.n675 4.5005
R7962 VSS.n919 VSS.n664 4.5005
R7963 VSS.n1019 VSS.n585 4.5005
R7964 VSS.n2007 VSS.n580 4.5005
R7965 VSS.n1021 VSS.n1020 4.5005
R7966 VSS.n2009 VSS.n2008 4.5005
R7967 VSS.n2000 VSS.n573 4.5005
R7968 VSS.n590 VSS.n581 4.5005
R7969 VSS.n578 VSS.n576 4.5005
R7970 VSS.n589 VSS.n584 4.5005
R7971 VSS.n1761 VSS.n1760 4.5005
R7972 VSS.n1751 VSS.n1750 4.5005
R7973 VSS.n1457 VSS.n1456 4.5005
R7974 VSS.n1749 VSS.n1451 4.5005
R7975 VSS.n1743 VSS.n1742 4.5005
R7976 VSS.n1753 VSS.n1454 4.5005
R7977 VSS.n1598 VSS.n1450 4.5005
R7978 VSS.n1754 VSS.n1455 4.5005
R7979 VSS.n1867 VSS.n1866 4.5005
R7980 VSS.n1865 VSS.n1813 4.5005
R7981 VSS.n1874 VSS.n1434 4.5005
R7982 VSS.n1869 VSS.n1435 4.5005
R7983 VSS.n2177 VSS.n2176 4.39555
R7984 VSS.n2082 VSS.n2081 4.39555
R7985 VSS.n515 VSS.n514 4.39555
R7986 VSS.n2095 VSS.n2092 4.39555
R7987 VSS.n2198 VSS.n2136 4.39555
R7988 VSS.n2145 VSS.n2144 4.39555
R7989 VSS.n1317 VSS.n1316 4.39555
R7990 VSS.n1322 VSS.n1321 4.39555
R7991 VSS.n1360 VSS.n1359 4.39555
R7992 VSS.n1340 VSS.n1339 4.39555
R7993 VSS.n1280 VSS.n1279 4.39555
R7994 VSS.n1256 VSS.n1246 4.39555
R7995 VSS.n1229 VSS.n1228 4.39555
R7996 VSS.n1399 VSS.n1398 4.39555
R7997 VSS.n1926 VSS.n1418 4.39555
R7998 VSS.n1940 VSS.n1072 4.39555
R7999 VSS.n1389 VSS.n1388 4.39555
R8000 VSS.n1213 VSS.n1212 4.39555
R8001 VSS.n2106 VSS.n2105 4.39555
R8002 VSS.n2056 VSS.n554 4.39555
R8003 VSS.n1437 VSS.n1436 4.39555
R8004 VSS.n557 VSS.n556 4.30289
R8005 VSS.n2061 VSS.n548 4.12333
R8006 VSS.n1772 VSS.n1771 4.09657
R8007 VSS.n1044 VSS.n1043 4.07463
R8008 VSS.n1329 VSS.t764 3.99804
R8009 VSS.n2185 VSS.t761 3.99804
R8010 VSS VSS.n1949 3.8414
R8011 VSS.n2203 VSS.n2133 3.83333
R8012 VSS.n2156 VSS.n2148 3.83333
R8013 VSS.n1349 VSS.n1271 3.83333
R8014 VSS.n1291 VSS.n1283 3.83333
R8015 VSS.n1408 VSS.n1081 3.83333
R8016 VSS.n1202 VSS.n1198 3.83333
R8017 VSS.n1197 VSS.n1196 3.83333
R8018 VSS.n552 VSS.n549 3.83333
R8019 VSS.n209 VSS.n104 3.79837
R8020 VSS.n1168 VSS.n1165 3.79837
R8021 VSS.n254 VSS.n251 3.79837
R8022 VSS.n2492 VSS.n268 3.79837
R8023 VSS.n287 VSS.n282 3.79837
R8024 VSS.n2474 VSS.n298 3.79837
R8025 VSS.n344 VSS.n339 3.79837
R8026 VSS.n2523 VSS.n232 3.79837
R8027 VSS.n2716 VSS.n2626 3.79837
R8028 VSS.n2672 VSS.n2667 3.79837
R8029 VSS.n2734 VSS.n2599 3.79837
R8030 VSS.n2615 VSS.n2613 3.79837
R8031 VSS.n2768 VSS.n71 3.79837
R8032 VSS.n2585 VSS.n90 3.79837
R8033 VSS.n2440 VSS.n389 3.76876
R8034 VSS.n2084 VSS.n529 3.76876
R8035 VSS.n2097 VSS.n2091 3.76876
R8036 VSS.n2153 VSS.n2150 3.76876
R8037 VSS.n2200 VSS.n2135 3.76876
R8038 VSS.n1148 VSS.n1103 3.76876
R8039 VSS.n1156 VSS.n1101 3.76876
R8040 VSS.n1304 VSS.n1299 3.76876
R8041 VSS.n1288 VSS.n1285 3.76876
R8042 VSS.n1270 VSS.n1269 3.76876
R8043 VSS.n1254 VSS.n1247 3.76876
R8044 VSS.n1243 VSS.n1241 3.76876
R8045 VSS.n1225 VSS.n1218 3.76876
R8046 VSS.n1924 VSS.n1419 3.76876
R8047 VSS.n1942 VSS.n1071 3.76876
R8048 VSS.n1080 VSS.n1079 3.76876
R8049 VSS.n1189 VSS.n1188 3.76876
R8050 VSS.n1233 VSS.n1216 3.76876
R8051 VSS.n2458 VSS.n381 3.76876
R8052 VSS.n198 VSS.n188 3.76876
R8053 VSS.n186 VSS.n109 3.76876
R8054 VSS.n2117 VSS.n517 3.76876
R8055 VSS.n2108 VSS.n524 3.76876
R8056 VSS.n2447 VSS.n386 3.76876
R8057 VSS.n2054 VSS.n2053 3.76876
R8058 VSS.n1868 VSS.n1811 3.76876
R8059 VSS.n2029 VSS.n564 3.76485
R8060 VSS.n1805 VSS.n1804 3.7496
R8061 VSS.n209 VSS.n102 3.7239
R8062 VSS.n1168 VSS.n1097 3.7239
R8063 VSS.n254 VSS.n250 3.7239
R8064 VSS.n2488 VSS.n268 3.7239
R8065 VSS.n2485 VSS.n282 3.7239
R8066 VSS.n2470 VSS.n298 3.7239
R8067 VSS.n2467 VSS.n339 3.7239
R8068 VSS.n2519 VSS.n232 3.7239
R8069 VSS.n2712 VSS.n2626 3.7239
R8070 VSS.n2709 VSS.n2667 3.7239
R8071 VSS.n2730 VSS.n2599 3.7239
R8072 VSS.n2727 VSS.n2613 3.7239
R8073 VSS.n2764 VSS.n71 3.7239
R8074 VSS.n2585 VSS.n89 3.7239
R8075 VSS.n2444 VSS.n2443 3.70003
R8076 VSS.n1 VSS.n0 3.66898
R8077 VSS.n391 VSS.n390 3.66898
R8078 VSS.n528 VSS.n527 3.66898
R8079 VSS.n519 VSS.n518 3.66898
R8080 VSS.n2099 VSS.n2090 3.66898
R8081 VSS.n510 VSS.n509 3.66898
R8082 VSS.n2147 VSS.n2146 3.66898
R8083 VSS.n383 VSS.n382 3.66898
R8084 VSS.n2449 VSS.n2448 3.66898
R8085 VSS.n1301 VSS.n1300 3.66898
R8086 VSS.n1240 VSS.n1239 3.66898
R8087 VSS.n1353 VSS.n1268 3.66898
R8088 VSS.n1282 VSS.n1281 3.66898
R8089 VSS.n1252 VSS.n1250 3.66898
R8090 VSS.n1215 VSS.n1214 3.66898
R8091 VSS.n1223 VSS.n1221 3.66898
R8092 VSS.n1922 VSS.n1421 3.66898
R8093 VSS.n1070 VSS.n1069 3.66898
R8094 VSS.n1412 VSS.n1078 3.66898
R8095 VSS.n1206 VSS.n1195 3.66898
R8096 VSS.n523 VSS.n522 3.66898
R8097 VSS.n2065 VSS.n534 3.66898
R8098 VSS.n334 VSS.n299 3.61615
R8099 VSS.n277 VSS.n269 3.61615
R8100 VSS.n286 VSS.n284 3.61615
R8101 VSS.n343 VSS.n341 3.61615
R8102 VSS.n2525 VSS.n230 3.61615
R8103 VSS.n228 VSS.n227 3.61615
R8104 VSS.n1163 VSS.n1098 3.61615
R8105 VSS.n2770 VSS.n69 3.61615
R8106 VSS.n2662 VSS.n2627 3.61615
R8107 VSS.n2608 VSS.n2600 3.61615
R8108 VSS.n2671 VSS.n2669 3.61615
R8109 VSS.n2596 VSS.n2595 3.61615
R8110 VSS.n2582 VSS.n91 3.61615
R8111 VSS.n206 VSS.n105 3.61615
R8112 VSS.n165 VSS.n164 3.60833
R8113 VSS.n2049 VSS.n2047 3.60833
R8114 VSS.n2072 VSS.n532 3.60833
R8115 VSS.n2165 VSS.n2164 3.60833
R8116 VSS.n2194 VSS.n2138 3.60833
R8117 VSS.n2189 VSS.n2142 3.60833
R8118 VSS.n2125 VSS.n2124 3.60833
R8119 VSS.n1307 VSS.n1306 3.60833
R8120 VSS.n1338 VSS.n1274 3.60833
R8121 VSS.n1333 VSS.n1277 3.60833
R8122 VSS.n1357 VSS.n1261 3.60833
R8123 VSS.n1264 VSS.n1263 3.60833
R8124 VSS.n1934 VSS.n1414 3.60833
R8125 VSS.n1931 VSS.n1930 3.60833
R8126 VSS.n1397 VSS.n1084 3.60833
R8127 VSS.n1210 VSS.n1209 3.60833
R8128 VSS.n1192 VSS.n1190 3.60833
R8129 VSS.n1379 VSS.n1207 3.60833
R8130 VSS.n1311 VSS.n1310 3.60833
R8131 VSS.n2128 VSS.n511 3.60833
R8132 VSS.n2171 VSS.n2170 3.60833
R8133 VSS.n531 VSS.n530 3.60833
R8134 VSS.n1807 VSS.n1806 3.60833
R8135 VSS.n1062 VSS.n1045 3.59463
R8136 VSS.n1060 VSS.n1046 3.59463
R8137 VSS.n1048 VSS.n1047 3.59463
R8138 VSS.n1056 VSS.n1050 3.59463
R8139 VSS.n1053 VSS.n1051 3.59463
R8140 VSS.t188 VSS.n1145 3.57455
R8141 VSS.n180 VSS.t1107 3.56931
R8142 VSS.n1804 VSS.n1438 3.45169
R8143 VSS.t897 VSS.n1912 3.35794
R8144 VSS.n1150 VSS.n1148 3.12356
R8145 VSS.n2481 VSS.n293 3.11877
R8146 VSS.n2503 VSS.n2502 3.11877
R8147 VSS.n2723 VSS.n2621 3.11877
R8148 VSS.n2748 VSS.n2747 3.11877
R8149 VSS.n2481 VSS.n292 3.07838
R8150 VSS.n2502 VSS.n243 3.07838
R8151 VSS.n2723 VSS.n2620 3.07838
R8152 VSS.n2747 VSS.n82 3.07838
R8153 VSS.n2899 VSS.n2898 3.01251
R8154 VSS.n175 VSS.n173 2.96041
R8155 VSS.n547 VSS.n546 2.73113
R8156 VSS.n1634 VSS.n1633 2.61344
R8157 VSS.n1637 VSS.n1636 2.61344
R8158 VSS.n1642 VSS.n1641 2.61344
R8159 VSS.n1645 VSS.n1644 2.61344
R8160 VSS.n1650 VSS.n1649 2.61344
R8161 VSS.n1653 VSS.n1652 2.61344
R8162 VSS.n1658 VSS.n1657 2.61344
R8163 VSS.n1661 VSS.n1660 2.61344
R8164 VSS.n1666 VSS.n1665 2.61344
R8165 VSS.n1669 VSS.n1668 2.61344
R8166 VSS.n1674 VSS.n1673 2.61344
R8167 VSS.n1677 VSS.n1676 2.61344
R8168 VSS.n1682 VSS.n1681 2.61344
R8169 VSS.n1685 VSS.n1684 2.61344
R8170 VSS.n1690 VSS.n1689 2.61344
R8171 VSS.n1693 VSS.n1692 2.61344
R8172 VSS.n1698 VSS.n1697 2.61344
R8173 VSS.n1701 VSS.n1700 2.61344
R8174 VSS.n1706 VSS.n1705 2.61344
R8175 VSS.n1709 VSS.n1708 2.61344
R8176 VSS.n1714 VSS.n1713 2.61344
R8177 VSS.n1717 VSS.n1716 2.61344
R8178 VSS.n1722 VSS.n1721 2.61344
R8179 VSS.n1725 VSS.n1724 2.61344
R8180 VSS.n1730 VSS.n1729 2.61344
R8181 VSS.n1733 VSS.n1732 2.61344
R8182 VSS.n1738 VSS.n1737 2.61344
R8183 VSS.n1745 VSS.n1599 2.61344
R8184 VSS.n1747 VSS.n1746 2.61344
R8185 VSS.n1757 VSS.n1756 2.61344
R8186 VSS.n2019 VSS.n569 2.61344
R8187 VSS.n2018 VSS.n2017 2.61344
R8188 VSS.n2012 VSS.n574 2.61344
R8189 VSS.n2011 VSS.n575 2.61344
R8190 VSS.n1017 VSS.n594 2.61344
R8191 VSS.n1016 VSS.n1015 2.61344
R8192 VSS.n1009 VSS.n595 2.61344
R8193 VSS.n1008 VSS.n1007 2.61344
R8194 VSS.n1001 VSS.n597 2.61344
R8195 VSS.n616 VSS.n609 2.61344
R8196 VSS.n621 VSS.n620 2.61344
R8197 VSS.n624 VSS.n623 2.61344
R8198 VSS.n629 VSS.n628 2.61344
R8199 VSS.n632 VSS.n631 2.61344
R8200 VSS.n1015 VSS.n1014 2.61344
R8201 VSS.n1010 VSS.n1009 2.61344
R8202 VSS.n1007 VSS.n1006 2.61344
R8203 VSS.n1002 VSS.n1001 2.61344
R8204 VSS.n617 VSS.n616 2.61344
R8205 VSS.n622 VSS.n621 2.61344
R8206 VSS.n623 VSS.n614 2.61344
R8207 VSS.n630 VSS.n629 2.61344
R8208 VSS.n631 VSS.n611 2.61344
R8209 VSS.n588 VSS.n575 2.61344
R8210 VSS.n594 VSS.n593 2.61344
R8211 VSS.n2020 VSS.n2019 2.61344
R8212 VSS.n2017 VSS.n2016 2.61344
R8213 VSS.n574 VSS.n572 2.61344
R8214 VSS.n1746 VSS.n1597 2.61344
R8215 VSS.n1758 VSS.n1757 2.61344
R8216 VSS.n1635 VSS.n1634 2.61344
R8217 VSS.n1636 VSS.n1625 2.61344
R8218 VSS.n1643 VSS.n1642 2.61344
R8219 VSS.n1644 VSS.n1623 2.61344
R8220 VSS.n1651 VSS.n1650 2.61344
R8221 VSS.n1652 VSS.n1621 2.61344
R8222 VSS.n1659 VSS.n1658 2.61344
R8223 VSS.n1660 VSS.n1619 2.61344
R8224 VSS.n1667 VSS.n1666 2.61344
R8225 VSS.n1668 VSS.n1617 2.61344
R8226 VSS.n1675 VSS.n1674 2.61344
R8227 VSS.n1676 VSS.n1615 2.61344
R8228 VSS.n1683 VSS.n1682 2.61344
R8229 VSS.n1684 VSS.n1613 2.61344
R8230 VSS.n1691 VSS.n1690 2.61344
R8231 VSS.n1692 VSS.n1611 2.61344
R8232 VSS.n1699 VSS.n1698 2.61344
R8233 VSS.n1700 VSS.n1609 2.61344
R8234 VSS.n1707 VSS.n1706 2.61344
R8235 VSS.n1708 VSS.n1607 2.61344
R8236 VSS.n1715 VSS.n1714 2.61344
R8237 VSS.n1716 VSS.n1605 2.61344
R8238 VSS.n1723 VSS.n1722 2.61344
R8239 VSS.n1724 VSS.n1603 2.61344
R8240 VSS.n1731 VSS.n1730 2.61344
R8241 VSS.n1732 VSS.n1601 2.61344
R8242 VSS.n1739 VSS.n1738 2.61344
R8243 VSS.n1740 VSS.n1599 2.61344
R8244 VSS.n1628 VSS.n1627 2.57967
R8245 VSS.n1629 VSS.n1628 2.57967
R8246 VSS.n2835 VSS.n2834 2.53357
R8247 VSS.n2501 VSS.n262 2.45051
R8248 VSS.n2746 VSS.n2593 2.45051
R8249 VSS.n351 VSS.n347 2.39297
R8250 VSS.n312 VSS.n290 2.39297
R8251 VSS.n248 VSS.n245 2.39297
R8252 VSS.n1173 VSS.n1172 2.39297
R8253 VSS.n2679 VSS.n2675 2.39297
R8254 VSS.n2640 VSS.n2618 2.39297
R8255 VSS.n87 VSS.n84 2.39297
R8256 VSS.n1032 VSS.n1027 2.37619
R8257 VSS.n216 VSS.n215 2.34602
R8258 VSS.n307 VSS.n306 2.34602
R8259 VSS.n361 VSS.n360 2.34602
R8260 VSS.n240 VSS.n235 2.34602
R8261 VSS.n79 VSS.n74 2.34602
R8262 VSS.n2635 VSS.n2634 2.34602
R8263 VSS.n2689 VSS.n2688 2.34602
R8264 VSS.n146 VSS.n145 2.31541
R8265 VSS.n543 VSS.n542 2.30642
R8266 VSS.n2837 VSS.n13 2.30135
R8267 VSS.n1024 VSS.n583 2.29751
R8268 VSS.n1762 VSS.n1453 2.29751
R8269 VSS.n2460 VSS.n47 2.296
R8270 VSS.n2789 VSS.n56 2.29314
R8271 VSS.n1779 VSS.n1778 2.29039
R8272 VSS.n2556 VSS.n2552 2.27007
R8273 VSS.n2481 VSS.n2480 2.21254
R8274 VSS.n2723 VSS.n2722 2.21254
R8275 VSS.n2201 VSS.n510 2.17814
R8276 VSS.n1353 VSS.n1352 2.17814
R8277 VSS.n2154 VSS.n2147 2.17664
R8278 VSS.n1289 VSS.n1282 2.17664
R8279 VSS.n1412 VSS.n1411 2.17664
R8280 VSS.n170 VSS.n169 2.10867
R8281 VSS VSS.n2483 2.09372
R8282 VSS.n260 VSS 2.09372
R8283 VSS VSS.n1174 2.09372
R8284 VSS VSS.n2707 2.09372
R8285 VSS VSS.n2725 2.09372
R8286 VSS.n2591 VSS 2.09372
R8287 VSS.n2784 VSS.n2783 2.07629
R8288 VSS.n328 VSS.n327 2.06712
R8289 VSS.n2656 VSS.n2655 2.06712
R8290 VSS.n305 VSS 1.99329
R8291 VSS VSS.n2517 1.99329
R8292 VSS VSS.n2762 1.99329
R8293 VSS.n2633 VSS 1.99329
R8294 VSS.n359 VSS 1.99329
R8295 VSS.n2687 VSS 1.99329
R8296 VSS.n214 VSS 1.9923
R8297 VSS.n2833 VSS.n20 1.91985
R8298 VSS.n1813 VSS.n1812 1.8127
R8299 VSS.n1348 VSS.n1347 1.73383
R8300 VSS.n1294 VSS.n1293 1.73383
R8301 VSS.n2205 VSS.n2204 1.73383
R8302 VSS.n2159 VSS.n2158 1.73383
R8303 VSS.n2060 VSS.n2059 1.73383
R8304 VSS.n1407 VSS.n1406 1.73383
R8305 VSS.n1201 VSS.n1200 1.73383
R8306 VSS.n2783 VSS.n24 1.73383
R8307 VSS.n2045 VSS.n2044 1.64468
R8308 VSS VSS.n2465 1.61221
R8309 VSS.n2141 VSS.n2139 1.58545
R8310 VSS.n1205 VSS.n1204 1.54391
R8311 VSS.n2064 VSS.n535 1.5047
R8312 VSS.n2848 VSS.n10 1.49567
R8313 VSS.n0 VSS.t1033 1.463
R8314 VSS.n0 VSS.t1020 1.463
R8315 VSS.n164 VSS.t1143 1.463
R8316 VSS.n164 VSS.t832 1.463
R8317 VSS.n1949 VSS.t1206 1.463
R8318 VSS.n1949 VSS.t828 1.463
R8319 VSS.n2047 VSS.t270 1.463
R8320 VSS.n2047 VSS.t300 1.463
R8321 VSS.n532 VSS.t307 1.463
R8322 VSS.n532 VSS.t510 1.463
R8323 VSS.n2176 VSS.t816 1.463
R8324 VSS.n2176 VSS.t819 1.463
R8325 VSS.n2164 VSS.t112 1.463
R8326 VSS.n2164 VSS.t517 1.463
R8327 VSS.n390 VSS.t763 1.463
R8328 VSS.n390 VSS.t777 1.463
R8329 VSS.n389 VSS.t1134 1.463
R8330 VSS.n389 VSS.t1141 1.463
R8331 VSS.n527 VSS.t983 1.463
R8332 VSS.n527 VSS.t987 1.463
R8333 VSS.n529 VSS.t1031 1.463
R8334 VSS.n529 VSS.t1034 1.463
R8335 VSS.n2081 VSS.t974 1.463
R8336 VSS.n2081 VSS.t976 1.463
R8337 VSS.n518 VSS.t1008 1.463
R8338 VSS.n518 VSS.t997 1.463
R8339 VSS.n514 VSS.t700 1.463
R8340 VSS.n514 VSS.t704 1.463
R8341 VSS.n2092 VSS.t127 1.463
R8342 VSS.n2092 VSS.t129 1.463
R8343 VSS.n2090 VSS.t1003 1.463
R8344 VSS.n2090 VSS.t985 1.463
R8345 VSS.n2091 VSS.t778 1.463
R8346 VSS.n2091 VSS.t779 1.463
R8347 VSS.n509 VSS.t1000 1.463
R8348 VSS.n509 VSS.t1007 1.463
R8349 VSS.n2134 VSS.t414 1.463
R8350 VSS.n2134 VSS.t131 1.463
R8351 VSS.n2133 VSS.t205 1.463
R8352 VSS.n2133 VSS.t416 1.463
R8353 VSS.n2132 VSS.t315 1.463
R8354 VSS.n2132 VSS.t209 1.463
R8355 VSS.n2136 VSS.t443 1.463
R8356 VSS.n2136 VSS.t441 1.463
R8357 VSS.n2138 VSS.t244 1.463
R8358 VSS.n2138 VSS.t917 1.463
R8359 VSS.n2144 VSS.t143 1.463
R8360 VSS.n2144 VSS.t141 1.463
R8361 VSS.n2149 VSS.t139 1.463
R8362 VSS.n2149 VSS.t323 1.463
R8363 VSS.n2148 VSS.t321 1.463
R8364 VSS.n2148 VSS.t682 1.463
R8365 VSS.n2157 VSS.t678 1.463
R8366 VSS.n2157 VSS.t921 1.463
R8367 VSS.n2146 VSS.t750 1.463
R8368 VSS.n2146 VSS.t762 1.463
R8369 VSS.n2150 VSS.t1133 1.463
R8370 VSS.n2150 VSS.t1140 1.463
R8371 VSS.n2142 VSS.t319 1.463
R8372 VSS.n2142 VSS.t200 1.463
R8373 VSS.n2135 VSS.t787 1.463
R8374 VSS.n2135 VSS.t789 1.463
R8375 VSS.n2124 VSS.t695 1.463
R8376 VSS.n2124 VSS.t123 1.463
R8377 VSS.n190 VSS.t334 1.463
R8378 VSS.n190 VSS.t1089 1.463
R8379 VSS.n93 VSS.t491 1.463
R8380 VSS.n93 VSS.t803 1.463
R8381 VSS.n1103 VSS.t1078 1.463
R8382 VSS.n1103 VSS.t1076 1.463
R8383 VSS.n1101 VSS.t488 1.463
R8384 VSS.n1101 VSS.t486 1.463
R8385 VSS.n1089 VSS.t477 1.463
R8386 VSS.n1089 VSS.t835 1.463
R8387 VSS.n1093 VSS.t474 1.463
R8388 VSS.n1093 VSS.t1210 1.463
R8389 VSS.n1316 VSS.t873 1.463
R8390 VSS.n1316 VSS.t876 1.463
R8391 VSS.n382 VSS.t759 1.463
R8392 VSS.n382 VSS.t773 1.463
R8393 VSS.n2448 VSS.t755 1.463
R8394 VSS.n2448 VSS.t767 1.463
R8395 VSS.n1300 VSS.t757 1.463
R8396 VSS.n1300 VSS.t769 1.463
R8397 VSS.n1306 VSS.t479 1.463
R8398 VSS.n1306 VSS.t520 1.463
R8399 VSS.n1299 VSS.t671 1.463
R8400 VSS.n1299 VSS.t660 1.463
R8401 VSS.n1321 VSS.t1082 1.463
R8402 VSS.n1321 VSS.t1080 1.463
R8403 VSS.n1239 VSS.t592 1.463
R8404 VSS.n1239 VSS.t627 1.463
R8405 VSS.n1359 VSS.t1165 1.463
R8406 VSS.n1359 VSS.t1167 1.463
R8407 VSS.n1268 VSS.t630 1.463
R8408 VSS.n1268 VSS.t646 1.463
R8409 VSS.n1350 VSS.t433 1.463
R8410 VSS.n1350 VSS.t572 1.463
R8411 VSS.n1271 VSS.t1251 1.463
R8412 VSS.n1271 VSS.t431 1.463
R8413 VSS.n1272 VSS.t929 1.463
R8414 VSS.n1272 VSS.t1249 1.463
R8415 VSS.n1339 VSS.t407 1.463
R8416 VSS.n1339 VSS.t405 1.463
R8417 VSS.n1274 VSS.t393 1.463
R8418 VSS.n1274 VSS.t105 1.463
R8419 VSS.n1279 VSS.t484 1.463
R8420 VSS.n1279 VSS.t482 1.463
R8421 VSS.n1284 VSS.t1084 1.463
R8422 VSS.n1284 VSS.t185 1.463
R8423 VSS.n1283 VSS.t183 1.463
R8424 VSS.n1283 VSS.t1173 1.463
R8425 VSS.n1292 VSS.t1175 1.463
R8426 VSS.n1292 VSS.t312 1.463
R8427 VSS.n1281 VSS.t753 1.463
R8428 VSS.n1281 VSS.t765 1.463
R8429 VSS.n1285 VSS.t670 1.463
R8430 VSS.n1285 VSS.t675 1.463
R8431 VSS.n1277 VSS.t435 1.463
R8432 VSS.n1277 VSS.t465 1.463
R8433 VSS.n1269 VSS.t1054 1.463
R8434 VSS.n1269 VSS.t1058 1.463
R8435 VSS.n1261 VSS.t246 1.463
R8436 VSS.n1261 VSS.t147 1.463
R8437 VSS.n1246 VSS.t568 1.463
R8438 VSS.n1246 VSS.t570 1.463
R8439 VSS.n1250 VSS.t603 1.463
R8440 VSS.n1250 VSS.t638 1.463
R8441 VSS.n1247 VSS.t1047 1.463
R8442 VSS.n1247 VSS.t1050 1.463
R8443 VSS.n1263 VSS.t427 1.463
R8444 VSS.n1263 VSS.t262 1.463
R8445 VSS.n1241 VSS.t18 1.463
R8446 VSS.n1241 VSS.t3 1.463
R8447 VSS.n1214 VSS.t623 1.463
R8448 VSS.n1214 VSS.t633 1.463
R8449 VSS.n1228 VSS.t523 1.463
R8450 VSS.n1228 VSS.t525 1.463
R8451 VSS.n1221 VSS.t634 1.463
R8452 VSS.n1221 VSS.t641 1.463
R8453 VSS.n1218 VSS.t1183 1.463
R8454 VSS.n1218 VSS.t1184 1.463
R8455 VSS.n1082 VSS.t362 1.463
R8456 VSS.n1082 VSS.t684 1.463
R8457 VSS.n1081 VSS.t686 1.463
R8458 VSS.n1081 VSS.t459 1.463
R8459 VSS.n1409 VSS.t461 1.463
R8460 VSS.n1409 VSS.t529 1.463
R8461 VSS.n1398 VSS.t419 1.463
R8462 VSS.n1398 VSS.t421 1.463
R8463 VSS.n1418 VSS.t963 1.463
R8464 VSS.n1418 VSS.t960 1.463
R8465 VSS.n1421 VSS.t598 1.463
R8466 VSS.n1421 VSS.t606 1.463
R8467 VSS.n1419 VSS.t51 1.463
R8468 VSS.n1419 VSS.t54 1.463
R8469 VSS.n1072 VSS.t533 1.463
R8470 VSS.n1072 VSS.t531 1.463
R8471 VSS.n1069 VSS.t647 1.463
R8472 VSS.n1069 VSS.t594 1.463
R8473 VSS.n1071 VSS.t1226 1.463
R8474 VSS.n1071 VSS.t1225 1.463
R8475 VSS.n1414 VSS.t444 1.463
R8476 VSS.n1414 VSS.t177 1.463
R8477 VSS.n1930 VSS.t169 1.463
R8478 VSS.n1930 VSS.t201 1.463
R8479 VSS.n1078 VSS.t643 1.463
R8480 VSS.n1078 VSS.t640 1.463
R8481 VSS.n1079 VSS.t1216 1.463
R8482 VSS.n1079 VSS.t1228 1.463
R8483 VSS.n1084 VSS.t309 1.463
R8484 VSS.n1084 VSS.t439 1.463
R8485 VSS.n1199 VSS.t389 1.463
R8486 VSS.n1199 VSS.t368 1.463
R8487 VSS.n1198 VSS.t402 1.463
R8488 VSS.n1198 VSS.t385 1.463
R8489 VSS.n1196 VSS.t527 1.463
R8490 VSS.n1196 VSS.t400 1.463
R8491 VSS.n549 VSS.t1088 1.463
R8492 VSS.n549 VSS.t1272 1.463
R8493 VSS.n550 VSS.t978 1.463
R8494 VSS.n550 VSS.t1086 1.463
R8495 VSS.n548 VSS.t1276 1.463
R8496 VSS.n548 VSS.t187 1.463
R8497 VSS.n1209 VSS.t521 1.463
R8498 VSS.n1209 VSS.t121 1.463
R8499 VSS.n1195 VSS.t621 1.463
R8500 VSS.n1195 VSS.t596 1.463
R8501 VSS.n1190 VSS.t1279 1.463
R8502 VSS.n1190 VSS.t274 1.463
R8503 VSS.n1188 VSS.t1192 1.463
R8504 VSS.n1188 VSS.t1196 1.463
R8505 VSS.n1388 VSS.t238 1.463
R8506 VSS.n1388 VSS.t236 1.463
R8507 VSS.n1207 VSS.t159 1.463
R8508 VSS.n1207 VSS.t453 1.463
R8509 VSS.n1216 VSS.t67 1.463
R8510 VSS.n1216 VSS.t58 1.463
R8511 VSS.n1212 VSS.t1064 1.463
R8512 VSS.n1212 VSS.t1066 1.463
R8513 VSS.n1310 VSS.t497 1.463
R8514 VSS.n1310 VSS.t213 1.463
R8515 VSS.n381 VSS.t63 1.463
R8516 VSS.n381 VSS.t32 1.463
R8517 VSS.n299 VSS.t370 1.463
R8518 VSS.n299 VSS.t1222 1.463
R8519 VSS.n269 VSS.t281 1.463
R8520 VSS.n269 VSS.t1198 1.463
R8521 VSS.n284 VSS.t165 1.463
R8522 VSS.n284 VSS.t1127 1.463
R8523 VSS.n341 VSS.t296 1.463
R8524 VSS.n341 VSS.t1040 1.463
R8525 VSS.n230 VSS.t429 1.463
R8526 VSS.n230 VSS.t791 1.463
R8527 VSS.n227 VSS.t306 1.463
R8528 VSS.n227 VSS.t1052 1.463
R8529 VSS.n1098 VSS.t298 1.463
R8530 VSS.n1098 VSS.t673 1.463
R8531 VSS.n69 VSS.t381 1.463
R8532 VSS.n69 VSS.t783 1.463
R8533 VSS.n2627 VSS.t379 1.463
R8534 VSS.n2627 VSS.t1218 1.463
R8535 VSS.n2600 VSS.t167 1.463
R8536 VSS.n2600 VSS.t1190 1.463
R8537 VSS.n2669 VSS.t496 1.463
R8538 VSS.n2669 VSS.t1182 1.463
R8539 VSS.n2595 VSS.t473 1.463
R8540 VSS.n2595 VSS.t1138 1.463
R8541 VSS.n91 VSS.t927 1.463
R8542 VSS.n91 VSS.t1046 1.463
R8543 VSS.n188 VSS.t163 1.463
R8544 VSS.n188 VSS.t161 1.463
R8545 VSS.n109 VSS.t514 1.463
R8546 VSS.n109 VSS.t512 1.463
R8547 VSS.n105 VSS.t372 1.463
R8548 VSS.n105 VSS.t668 1.463
R8549 VSS.n511 VSS.t151 1.463
R8550 VSS.n511 VSS.t324 1.463
R8551 VSS.n517 VSS.t61 1.463
R8552 VSS.n517 VSS.t56 1.463
R8553 VSS.n522 VSS.t996 1.463
R8554 VSS.n522 VSS.t1001 1.463
R8555 VSS.n524 VSS.t11 1.463
R8556 VSS.n524 VSS.t5 1.463
R8557 VSS.n2105 VSS.t9 1.463
R8558 VSS.n2105 VSS.t103 1.463
R8559 VSS.n2170 VSS.t294 1.463
R8560 VSS.n2170 VSS.t423 1.463
R8561 VSS.n386 VSS.t72 1.463
R8562 VSS.n386 VSS.t44 1.463
R8563 VSS.n2443 VSS.t135 1.463
R8564 VSS.n2443 VSS.t137 1.463
R8565 VSS.n564 VSS.t346 1.463
R8566 VSS.n564 VSS.t348 1.463
R8567 VSS.n556 VSS.t970 1.463
R8568 VSS.n556 VSS.t1074 1.463
R8569 VSS.n554 VSS.t198 1.463
R8570 VSS.n554 VSS.t196 1.463
R8571 VSS.n530 VSS.t215 1.463
R8572 VSS.n530 VSS.t157 1.463
R8573 VSS.n534 VSS.t995 1.463
R8574 VSS.n534 VSS.t1010 1.463
R8575 VSS.n2053 VSS.t1018 1.463
R8576 VSS.n2053 VSS.t1022 1.463
R8577 VSS.n1029 VSS.t1265 1.463
R8578 VSS.n1029 VSS.t942 1.463
R8579 VSS.n1043 VSS.t1110 1.463
R8580 VSS.n1043 VSS.t1112 1.463
R8581 VSS.n1045 VSS.t717 1.463
R8582 VSS.n1045 VSS.t719 1.463
R8583 VSS.n1046 VSS.t799 1.463
R8584 VSS.n1046 VSS.t801 1.463
R8585 VSS.n1047 VSS.t727 1.463
R8586 VSS.n1047 VSS.t729 1.463
R8587 VSS.n1050 VSS.t576 1.463
R8588 VSS.n1050 VSS.t578 1.463
R8589 VSS.n1051 VSS.t715 1.463
R8590 VSS.n1051 VSS.t723 1.463
R8591 VSS.n1436 VSS.t653 1.463
R8592 VSS.n1436 VSS.t655 1.463
R8593 VSS.n1806 VSS.t293 1.463
R8594 VSS.n1806 VSS.t410 1.463
R8595 VSS.n1811 VSS.t1121 1.463
R8596 VSS.n1811 VSS.t1123 1.463
R8597 VSS VSS.n1179 1.4209
R8598 VSS VSS.n96 1.4209
R8599 VSS.n1238 VSS.n1237 1.41164
R8600 VSS.n1236 VSS.n1235 1.41164
R8601 VSS.n2115 VSS.n2114 1.41164
R8602 VSS.n2111 VSS.n2110 1.41164
R8603 VSS.n1917 VSS.n1420 1.41016
R8604 VSS.n1628 VSS.n1065 1.31166
R8605 VSS.n2439 VSS.n391 1.30108
R8606 VSS.n1303 VSS.n1301 1.30108
R8607 VSS.n1242 VSS.n1240 1.30108
R8608 VSS.n1234 VSS.n1215 1.30108
R8609 VSS.n1943 VSS.n1070 1.30108
R8610 VSS.n2116 VSS.n519 1.30108
R8611 VSS.n2109 VSS.n523 1.30108
R8612 VSS.n2085 VSS.n528 1.29958
R8613 VSS.n2099 VSS.n2098 1.29958
R8614 VSS.n2457 VSS.n383 1.29958
R8615 VSS.n2450 VSS.n2449 1.29958
R8616 VSS.n1253 VSS.n1252 1.29958
R8617 VSS.n1224 VSS.n1223 1.29958
R8618 VSS.n1923 VSS.n1922 1.29958
R8619 VSS.n594 VSS.n566 1.29478
R8620 VSS.n1015 VSS.n566 1.29478
R8621 VSS.n1009 VSS.n566 1.29478
R8622 VSS.n1007 VSS.n566 1.29478
R8623 VSS.n1001 VSS.n566 1.29478
R8624 VSS.n616 VSS.n560 1.29478
R8625 VSS.n621 VSS.n560 1.29478
R8626 VSS.n623 VSS.n560 1.29478
R8627 VSS.n629 VSS.n560 1.29478
R8628 VSS.n631 VSS.n560 1.29478
R8629 VSS.n574 VSS.n566 1.29478
R8630 VSS.n575 VSS.n566 1.29478
R8631 VSS.n2019 VSS.n566 1.29478
R8632 VSS.n2017 VSS.n566 1.29478
R8633 VSS.n1599 VSS.n1065 1.29478
R8634 VSS.n1746 VSS.n1065 1.29478
R8635 VSS.n1634 VSS.n1065 1.29478
R8636 VSS.n1636 VSS.n1065 1.29478
R8637 VSS.n1642 VSS.n1065 1.29478
R8638 VSS.n1644 VSS.n1065 1.29478
R8639 VSS.n1650 VSS.n1065 1.29478
R8640 VSS.n1652 VSS.n1065 1.29478
R8641 VSS.n1658 VSS.n1065 1.29478
R8642 VSS.n1660 VSS.n1065 1.29478
R8643 VSS.n1666 VSS.n1065 1.29478
R8644 VSS.n1668 VSS.n1065 1.29478
R8645 VSS.n1674 VSS.n1065 1.29478
R8646 VSS.n1676 VSS.n1065 1.29478
R8647 VSS.n1682 VSS.n1065 1.29478
R8648 VSS.n1684 VSS.n1065 1.29478
R8649 VSS.n1690 VSS.n1065 1.29478
R8650 VSS.n1692 VSS.n1065 1.29478
R8651 VSS.n1698 VSS.n1065 1.29478
R8652 VSS.n1700 VSS.n1065 1.29478
R8653 VSS.n1706 VSS.n1065 1.29478
R8654 VSS.n1708 VSS.n1065 1.29478
R8655 VSS.n1714 VSS.n1065 1.29478
R8656 VSS.n1716 VSS.n1065 1.29478
R8657 VSS.n1722 VSS.n1065 1.29478
R8658 VSS.n1724 VSS.n1065 1.29478
R8659 VSS.n1730 VSS.n1065 1.29478
R8660 VSS.n1732 VSS.n1065 1.29478
R8661 VSS.n1738 VSS.n1065 1.29478
R8662 VSS.n2464 VSS.n2463 1.27516
R8663 VSS.n1997 VSS.n1996 1.26524
R8664 VSS.n1276 VSS.n1275 1.25337
R8665 VSS.n1999 VSS.n10 1.20218
R8666 VSS.n2834 VSS.n2833 1.18807
R8667 VSS.n379 VSS.n347 1.17119
R8668 VSS.n2483 VSS.n290 1.17119
R8669 VSS.n260 VSS.n248 1.17119
R8670 VSS.n1174 VSS.n1173 1.17119
R8671 VSS.n2707 VSS.n2675 1.17119
R8672 VSS.n2725 VSS.n2618 1.17119
R8673 VSS.n2591 VSS.n87 1.17119
R8674 VSS.n2551 VSS.n221 1.15749
R8675 VSS.n193 VSS.n192 1.11939
R8676 VSS.n1092 VSS.n1091 1.11939
R8677 VSS.n1385 VSS.t595 1.11772
R8678 VSS.t629 VSS.n1354 1.11772
R8679 VSS.n2207 VSS.t999 1.11772
R8680 VSS.t1009 VSS.n2067 1.11772
R8681 VSS.t642 VSS.n1413 1.11772
R8682 VSS.n163 VSS.n19 1.11742
R8683 VSS.n507 VSS.n221 1.08721
R8684 VSS.n168 VSS.n162 1.07034
R8685 VSS.n169 VSS.n25 1.07034
R8686 VSS.n384 VSS.t768 1.03868
R8687 VSS.n1372 VSS.t632 1.03818
R8688 VSS.n1367 VSS.t591 1.03818
R8689 VSS.n2102 VSS.t986 1.03818
R8690 VSS.t1002 VSS.n2101 1.03818
R8691 VSS.n2436 VSS.t766 1.03818
R8692 VSS.t597 VSS.n1946 1.03818
R8693 VSS.n2848 VSS.n2847 1.03581
R8694 VSS.n2440 VSS.n2439 1.03184
R8695 VSS.n2085 VSS.n2084 1.03184
R8696 VSS.n2098 VSS.n2097 1.03184
R8697 VSS.n2458 VSS.n2457 1.03184
R8698 VSS.n1304 VSS.n1303 1.03184
R8699 VSS.n1254 VSS.n1253 1.03184
R8700 VSS.n1243 VSS.n1242 1.03184
R8701 VSS.n1234 VSS.n1233 1.03184
R8702 VSS.n1225 VSS.n1224 1.03184
R8703 VSS.n1924 VSS.n1923 1.03184
R8704 VSS.n1943 VSS.n1942 1.03184
R8705 VSS.n2117 VSS.n2116 1.03184
R8706 VSS.n2109 VSS.n2108 1.03184
R8707 VSS.n2450 VSS.n2447 1.0114
R8708 VSS.n163 VSS.n162 0.955147
R8709 VSS.n2500 VSS.n2499 0.939167
R8710 VSS.n2745 VSS.n2744 0.939167
R8711 VSS.n1997 VSS.n1028 0.936031
R8712 VSS.n2560 VSS.n2551 0.932808
R8713 VSS.n2457 VSS.n2456 0.92521
R8714 VSS.n2451 VSS.n2450 0.92521
R8715 VSS.n2906 VSS.t1019 0.909591
R8716 VSS.n2834 VSS.n19 0.899346
R8717 VSS.n2884 VSS.n2882 0.881611
R8718 VSS.n1135 VSS.n1133 0.881611
R8719 VSS.n1905 VSS.n1426 0.881611
R8720 VSS.n159 VSS.n112 0.881611
R8721 VSS.n1985 VSS.n1037 0.881611
R8722 VSS.n1822 VSS.n1819 0.881611
R8723 VSS.n166 VSS.n19 0.880263
R8724 VSS.n1403 VSS.n1397 0.877263
R8725 VSS.n2195 VSS.n2194 0.87647
R8726 VSS.n1344 VSS.n1338 0.87647
R8727 VSS.n2049 VSS.n2048 0.876129
R8728 VSS.n1193 VSS.n1192 0.875129
R8729 VSS.n1807 VSS.n1434 0.875129
R8730 VSS.n2189 VSS.n2188 0.874923
R8731 VSS.n1333 VSS.n1332 0.874923
R8732 VSS.n1157 VSS.n1156 0.874807
R8733 VSS.n198 VSS.n197 0.874807
R8734 VSS.n1866 VSS.n1435 0.845198
R8735 VSS.n2062 VSS.n547 0.839031
R8736 VSS.n167 VSS.n163 0.83553
R8737 VSS VSS.n2437 0.827919
R8738 VSS.n2087 VSS 0.827919
R8739 VSS.n2454 VSS 0.827919
R8740 VSS VSS.n1219 0.827919
R8741 VSS VSS.n2088 0.826952
R8742 VSS VSS.n1248 0.826952
R8743 VSS VSS.n1068 0.826952
R8744 VSS VSS.n2888 0.803833
R8745 VSS VSS.n2883 0.803833
R8746 VSS VSS.n1139 0.803833
R8747 VSS VSS.n1134 0.803833
R8748 VSS.n1901 VSS 0.803833
R8749 VSS.n1906 VSS 0.803833
R8750 VSS.n155 VSS 0.803833
R8751 VSS.n160 VSS 0.803833
R8752 VSS.n1981 VSS 0.803833
R8753 VSS.n1986 VSS 0.803833
R8754 VSS.n1837 VSS 0.803833
R8755 VSS.n1368 VSS.n1238 0.803577
R8756 VSS.n1371 VSS.n1235 0.803577
R8757 VSS.n2115 VSS.n520 0.803577
R8758 VSS.n2110 VSS.n521 0.803577
R8759 VSS.n1918 VSS.n1420 0.802588
R8760 VSS.n96 VSS.n95 0.777239
R8761 VSS.n1179 VSS.n1095 0.777239
R8762 VSS.n1996 VSS.n1031 0.777239
R8763 VSS.n2532 VSS 0.77007
R8764 VSS.n2573 VSS 0.77007
R8765 VSS.n2438 VSS.n392 0.728242
R8766 VSS.n2086 VSS.n526 0.728242
R8767 VSS.n2100 VSS.n2089 0.728242
R8768 VSS.n1302 VSS.n385 0.728242
R8769 VSS.n1251 VSS.n1249 0.728242
R8770 VSS.n1222 VSS.n1220 0.728242
R8771 VSS.n1945 VSS.n1944 0.728242
R8772 VSS.n2870 VSS.n2850 0.71601
R8773 VSS.n1121 VSS.n1105 0.71601
R8774 VSS.n1900 VSS.n1899 0.71601
R8775 VSS.n154 VSS.n153 0.71601
R8776 VSS.n1980 VSS.n1979 0.71601
R8777 VSS.n1826 VSS.n1825 0.71601
R8778 VSS.n1203 VSS.n1197 0.7085
R8779 VSS.n2563 VSS.n2562 0.699191
R8780 VSS.n192 VSS.n191 0.67334
R8781 VSS.n95 VSS.n94 0.67334
R8782 VSS.n1091 VSS.n1090 0.67334
R8783 VSS.n1095 VSS.n1094 0.67334
R8784 VSS.n1031 VSS.n1030 0.67334
R8785 VSS.n1061 VSS.n1060 0.671611
R8786 VSS.n377 VSS.n376 0.670885
R8787 VSS.n367 VSS.n366 0.670885
R8788 VSS.n239 VSS.n237 0.670885
R8789 VSS.n225 VSS.n224 0.670885
R8790 VSS.n78 VSS.n76 0.670885
R8791 VSS.n2695 VSS.n2694 0.670885
R8792 VSS.n2705 VSS.n2704 0.670885
R8793 VSS.n2004 VSS.n1999 0.662178
R8794 VSS.n2212 VSS.n2211 0.656724
R8795 VSS.n1148 VSS 0.655143
R8796 VSS.n1156 VSS 0.655143
R8797 VSS VSS.n198 0.655143
R8798 VSS.n186 VSS 0.655143
R8799 VSS.n2441 VSS.n2440 0.627286
R8800 VSS.n2084 VSS.n2083 0.627286
R8801 VSS.n2097 VSS.n2096 0.627286
R8802 VSS.n2153 VSS.n2152 0.627286
R8803 VSS.n2200 VSS.n2199 0.627286
R8804 VSS.n1323 VSS.n1304 0.627286
R8805 VSS.n1288 VSS.n1287 0.627286
R8806 VSS.n1273 VSS.n1270 0.627286
R8807 VSS.n1255 VSS.n1254 0.627286
R8808 VSS.n1244 VSS.n1243 0.627286
R8809 VSS.n1230 VSS.n1225 0.627286
R8810 VSS.n1925 VSS.n1924 0.627286
R8811 VSS.n1942 VSS.n1941 0.627286
R8812 VSS.n1083 VSS.n1080 0.627286
R8813 VSS.n1390 VSS.n1189 0.627286
R8814 VSS.n1233 VSS.n1232 0.627286
R8815 VSS.n2118 VSS.n2117 0.627286
R8816 VSS.n2108 VSS.n2107 0.627286
R8817 VSS.n2055 VSS.n2054 0.627286
R8818 VSS.n1869 VSS.n1868 0.627286
R8819 VSS.n2502 VSS.n2501 0.597038
R8820 VSS.n2747 VSS.n2746 0.597038
R8821 VSS.n2065 VSS.n2064 0.590319
R8822 VSS.n2063 VSS.n536 0.584346
R8823 VSS.n1848 VSS 0.582722
R8824 VSS.n2868 VSS 0.582722
R8825 VSS.n1119 VSS 0.582722
R8826 VSS VSS.n117 0.582722
R8827 VSS VSS.n1041 0.582722
R8828 VSS VSS.n1430 0.582722
R8829 VSS.n1932 VSS.n1931 0.574328
R8830 VSS.n2126 VSS.n2125 0.573536
R8831 VSS.n1358 VSS.n1357 0.573536
R8832 VSS.n1934 VSS.n1933 0.573536
R8833 VSS.n1264 VSS.n1260 0.573328
R8834 VSS.n2128 VSS.n2127 0.573328
R8835 VSS.n2169 VSS.n2165 0.573195
R8836 VSS.n2075 VSS.n2072 0.573195
R8837 VSS.n1309 VSS.n1307 0.572195
R8838 VSS.n1377 VSS.n1210 0.572195
R8839 VSS.n1379 VSS.n1378 0.571989
R8840 VSS.n1312 VSS.n1311 0.571989
R8841 VSS.n2172 VSS.n2171 0.571989
R8842 VSS.n2076 VSS.n531 0.571989
R8843 VSS.n1179 VSS.n1178 0.568021
R8844 VSS.n2569 VSS.n96 0.568021
R8845 VSS.n1996 VSS.n1995 0.568021
R8846 VSS.n167 VSS.n166 0.561269
R8847 VSS.n1206 VSS.n1205 0.554405
R8848 VSS.n2446 VSS.n387 0.551399
R8849 VSS.n2444 VSS.n2442 0.534241
R8850 VSS.n2459 VSS.n380 0.527643
R8851 VSS.n360 VSS.n359 0.50401
R8852 VSS.n306 VSS.n305 0.50401
R8853 VSS.n2517 VSS.n235 0.50401
R8854 VSS.n2762 VSS.n74 0.50401
R8855 VSS.n2688 VSS.n2687 0.50401
R8856 VSS.n2634 VSS.n2633 0.50401
R8857 VSS.n215 VSS.n214 0.50401
R8858 VSS.n334 VSS.n333 0.50331
R8859 VSS.n277 VSS.n276 0.50331
R8860 VSS.n286 VSS.n285 0.50331
R8861 VSS.n343 VSS.n342 0.50331
R8862 VSS.n2526 VSS.n2525 0.50331
R8863 VSS.n2538 VSS.n228 0.50331
R8864 VSS.n1163 VSS.n1162 0.50331
R8865 VSS.n2771 VSS.n2770 0.50331
R8866 VSS.n2662 VSS.n2661 0.50331
R8867 VSS.n2608 VSS.n2607 0.50331
R8868 VSS.n2671 VSS.n2670 0.50331
R8869 VSS.n2739 VSS.n2596 0.50331
R8870 VSS.n2582 VSS.n2581 0.50331
R8871 VSS.n206 VSS.n205 0.50331
R8872 VSS.n168 VSS.n167 0.499494
R8873 VSS.n2858 VSS.n2857 0.487216
R8874 VSS.n124 VSS.n123 0.487216
R8875 VSS.n1955 VSS.n1954 0.487216
R8876 VSS.n1433 VSS.n1432 0.487216
R8877 VSS.n2465 VSS.n379 0.483016
R8878 VSS.n1062 VSS.n1061 0.4805
R8879 VSS.n1060 VSS.n1059 0.4805
R8880 VSS.n1049 VSS.n1048 0.4805
R8881 VSS.n1056 VSS.n1055 0.4805
R8882 VSS.n162 VSS.n25 0.467417
R8883 VSS.n2560 VSS.n2559 0.465605
R8884 VSS VSS.n1851 0.457167
R8885 VSS.n2853 VSS 0.457167
R8886 VSS.n1108 VSS 0.457167
R8887 VSS VSS.n140 0.457167
R8888 VSS VSS.n1967 0.457167
R8889 VSS VSS.n1887 0.457167
R8890 VSS.n1109 VSS.n8 0.454994
R8891 VSS.n1242 VSS.n1238 0.4505
R8892 VSS.n1235 VSS.n1234 0.4505
R8893 VSS.n1923 VSS.n1420 0.4505
R8894 VSS.n2116 VSS.n2115 0.4505
R8895 VSS.n2110 VSS.n2109 0.4505
R8896 VSS VSS.n9 0.44806
R8897 VSS.n366 VSS.n356 0.445885
R8898 VSS.n2513 VSS.n237 0.445885
R8899 VSS.n2758 VSS.n76 0.445885
R8900 VSS.n2694 VSS.n2684 0.445885
R8901 VSS.n327 VSS.n301 0.441269
R8902 VSS.n2655 VSS.n2629 0.441269
R8903 VSS VSS.n1056 0.434944
R8904 VSS.n166 VSS.n165 0.413044
R8905 VSS.n2061 VSS 0.4125
R8906 VSS.n378 VSS.n348 0.4055
R8907 VSS.n365 VSS.n364 0.4055
R8908 VSS.n325 VSS.n324 0.4055
R8909 VSS.n2482 VSS.n291 0.4055
R8910 VSS.n2515 VSS.n2514 0.4055
R8911 VSS.n261 VSS.n244 0.4055
R8912 VSS.n2760 VSS.n2759 0.4055
R8913 VSS.n2693 VSS.n2692 0.4055
R8914 VSS.n2653 VSS.n2652 0.4055
R8915 VSS.n2706 VSS.n2676 0.4055
R8916 VSS.n2724 VSS.n2619 0.4055
R8917 VSS.n2592 VSS.n83 0.4055
R8918 VSS.n220 VSS.n219 0.4055
R8919 VSS.n377 VSS.n349 0.403192
R8920 VSS.n2548 VSS.n224 0.403192
R8921 VSS.n2705 VSS.n2677 0.403192
R8922 VSS.n358 VSS.n357 0.400885
R8923 VSS.n326 VSS.n302 0.400885
R8924 VSS.n304 VSS.n303 0.400885
R8925 VSS.n2516 VSS.n236 0.400885
R8926 VSS.n2761 VSS.n75 0.400885
R8927 VSS.n2686 VSS.n2685 0.400885
R8928 VSS.n2654 VSS.n2630 0.400885
R8929 VSS.n2632 VSS.n2631 0.400885
R8930 VSS.n100 VSS.n99 0.400885
R8931 VSS.n1863 VSS.n1861 0.398328
R8932 VSS.n2826 VSS.n25 0.393224
R8933 VSS.n2482 VSS.n2481 0.388192
R8934 VSS.n2502 VSS.n261 0.388192
R8935 VSS.n2724 VSS.n2723 0.388192
R8936 VSS.n2747 VSS.n2592 0.388192
R8937 VSS VSS.n2893 0.387167
R8938 VSS VSS.n1144 0.387167
R8939 VSS VSS.n161 0.387167
R8940 VSS.n1990 VSS 0.387167
R8941 VSS VSS.n1828 0.387167
R8942 VSS.n271 VSS.n263 0.37418
R8943 VSS.n2602 VSS.n2594 0.37418
R8944 VSS.n169 VSS.n168 0.367956
R8945 VSS VSS.n1062 0.364944
R8946 VSS VSS.n1048 0.364944
R8947 VSS VSS.n1053 0.364944
R8948 VSS.n2445 VSS.n388 0.362755
R8949 VSS.n1053 VSS.n1052 0.362722
R8950 VSS.n2562 VSS.n98 0.352423
R8951 VSS.n1827 VSS.n9 0.349633
R8952 VSS.n1851 VSS.n1850 0.347167
R8953 VSS.n2863 VSS.n2853 0.347167
R8954 VSS.n1114 VSS.n1108 0.347167
R8955 VSS.n140 VSS.n139 0.347167
R8956 VSS.n1967 VSS.n1966 0.347167
R8957 VSS.n1887 VSS.n1886 0.347167
R8958 VSS VSS.n2892 0.338278
R8959 VSS VSS.n1143 0.338278
R8960 VSS.n181 VSS 0.338278
R8961 VSS VSS.n1035 0.338278
R8962 VSS.n1833 VSS 0.338278
R8963 VSS.n1907 VSS 0.336905
R8964 VSS.n379 VSS.n378 0.3305
R8965 VSS.n2483 VSS.n2482 0.3305
R8966 VSS.n261 VSS.n260 0.3305
R8967 VSS.n2707 VSS.n2706 0.3305
R8968 VSS.n2725 VSS.n2724 0.3305
R8969 VSS.n2592 VSS.n2591 0.3305
R8970 VSS.n2550 VSS.n2549 0.330435
R8971 VSS.n1855 VSS.n1854 0.328278
R8972 VSS.n2867 VSS.n2854 0.328278
R8973 VSS.n1118 VSS.n1112 0.328278
R8974 VSS.n135 VSS.n134 0.328278
R8975 VSS.n1962 VSS.n1961 0.328278
R8976 VSS.n1882 VSS.n1881 0.328278
R8977 VSS.n1916 VSS.n1915 0.32733
R8978 VSS.n2172 VSS.n2169 0.320287
R8979 VSS.n1312 VSS.n1309 0.320287
R8980 VSS.n1358 VSS.n1260 0.320287
R8981 VSS.n1933 VSS.n1932 0.320287
R8982 VSS.n1378 VSS.n1377 0.320287
R8983 VSS.n2127 VSS.n2126 0.320287
R8984 VSS.n2076 VSS.n2075 0.320287
R8985 VSS.n332 VSS.n331 0.30866
R8986 VSS.n275 VSS.n274 0.30866
R8987 VSS.n2496 VSS.n264 0.30866
R8988 VSS.n2478 VSS.n294 0.30866
R8989 VSS.n2529 VSS.n229 0.30866
R8990 VSS.n2537 VSS.n2536 0.30866
R8991 VSS.n1161 VSS.n1160 0.30866
R8992 VSS.n2570 VSS.n68 0.30866
R8993 VSS.n2660 VSS.n2659 0.30866
R8994 VSS.n2606 VSS.n2605 0.30866
R8995 VSS.n2720 VSS.n2622 0.30866
R8996 VSS.n2741 VSS.n2740 0.30866
R8997 VSS.n2580 VSS.n2579 0.30866
R8998 VSS.n195 VSS.n106 0.30866
R8999 VSS.n2480 VSS.n2479 0.304466
R9000 VSS.n2722 VSS.n2721 0.304466
R9001 VSS.n1174 VSS.n222 0.303962
R9002 VSS.n2078 VSS.n2076 0.303434
R9003 VSS.n1309 VSS.n1308 0.303434
R9004 VSS.n1363 VSS.n1358 0.303434
R9005 VSS.n1377 VSS.n1376 0.303434
R9006 VSS.n1314 VSS.n1312 0.303434
R9007 VSS.n2126 VSS.n2123 0.303434
R9008 VSS.n2075 VSS.n2074 0.303434
R9009 VSS.n2174 VSS.n2172 0.303434
R9010 VSS.n2169 VSS.n2168 0.303434
R9011 VSS.n2127 VSS.n512 0.303434
R9012 VSS.n1260 VSS.n1259 0.303434
R9013 VSS.n1378 VSS.n1208 0.303434
R9014 VSS.n1932 VSS.n1929 0.303434
R9015 VSS.n1933 VSS.n1416 0.303434
R9016 VSS.n330 VSS.n328 0.301214
R9017 VSS.n2658 VSS.n2656 0.301214
R9018 VSS.n2874 VSS.n2872 0.293141
R9019 VSS.n1125 VSS.n1123 0.293141
R9020 VSS.n1893 VSS.n1427 0.293141
R9021 VSS.n147 VSS.n113 0.293141
R9022 VSS.n1973 VSS.n1038 0.293141
R9023 VSS.n1844 VSS.n1818 0.293141
R9024 VSS.n132 VSS.n131 0.286056
R9025 VSS.n1874 VSS.n1435 0.284171
R9026 VSS.n333 VSS.n300 0.27986
R9027 VSS.n276 VSS.n270 0.27986
R9028 VSS.n2527 VSS.n2526 0.27986
R9029 VSS.n2772 VSS.n2771 0.27986
R9030 VSS.n2661 VSS.n2628 0.27986
R9031 VSS.n2607 VSS.n2601 0.27986
R9032 VSS.n224 VSS.n222 0.279618
R9033 VSS.n273 VSS.n271 0.279241
R9034 VSS.n2604 VSS.n2602 0.279241
R9035 VSS.n285 VSS.n265 0.27914
R9036 VSS.n342 VSS.n295 0.27914
R9037 VSS.n2539 VSS.n2538 0.27914
R9038 VSS.n1162 VSS.n1099 0.27914
R9039 VSS.n2670 VSS.n2623 0.27914
R9040 VSS.n2739 VSS.n2738 0.27914
R9041 VSS.n2581 VSS.n92 0.27914
R9042 VSS.n205 VSS.n204 0.27914
R9043 VSS.n2433 VSS.n2432 0.276403
R9044 VSS VSS.n2184 0.271428
R9045 VSS.n2208 VSS 0.271428
R9046 VSS VSS.n1328 0.271428
R9047 VSS VSS.n1267 0.271428
R9048 VSS VSS.n1077 0.271428
R9049 VSS VSS.n1384 0.271428
R9050 VSS VSS.n2066 0.271428
R9051 VSS.n2499 VSS.n2498 0.26546
R9052 VSS.n2744 VSS.n2743 0.26546
R9053 VSS.n1866 VSS.n1865 0.265311
R9054 VSS.n2190 VSS.n2141 0.263577
R9055 VSS.n1337 VSS.n1275 0.263577
R9056 VSS.n1356 VSS.n1262 0.263577
R9057 VSS.n1075 VSS.n1074 0.263577
R9058 VSS.n1396 VSS.n1085 0.263577
R9059 VSS.n1383 VSS.n1382 0.263577
R9060 VSS.n1327 VSS.n1326 0.263577
R9061 VSS.n2183 VSS.n2182 0.263577
R9062 VSS.n2071 VSS.n533 0.263577
R9063 VSS.n2050 VSS.n2046 0.263577
R9064 VSS.n1808 VSS.n1805 0.263577
R9065 VSS.n1867 VSS.n1813 0.263
R9066 VSS.n2193 VSS.n2139 0.262423
R9067 VSS.n327 VSS.n326 0.26172
R9068 VSS.n2655 VSS.n2654 0.26172
R9069 VSS VSS.n1049 0.256056
R9070 VSS.n378 VSS.n377 0.25308
R9071 VSS.n2706 VSS.n2705 0.25308
R9072 VSS.n2063 VSS.n2062 0.251199
R9073 VSS.n349 VSS.n348 0.250885
R9074 VSS.n364 VSS.n356 0.250885
R9075 VSS.n324 VSS.n302 0.250885
R9076 VSS.n292 VSS.n291 0.250885
R9077 VSS.n2514 VSS.n2513 0.250885
R9078 VSS.n244 VSS.n243 0.250885
R9079 VSS.n2549 VSS.n2548 0.250885
R9080 VSS.n2759 VSS.n2758 0.250885
R9081 VSS.n2692 VSS.n2684 0.250885
R9082 VSS.n2652 VSS.n2630 0.250885
R9083 VSS.n2677 VSS.n2676 0.250885
R9084 VSS.n2620 VSS.n2619 0.250885
R9085 VSS.n83 VSS.n82 0.250885
R9086 VSS.n219 VSS.n98 0.250885
R9087 VSS.n2874 VSS.n2873 0.249389
R9088 VSS.n1125 VSS.n1124 0.249389
R9089 VSS.n1894 VSS.n1893 0.249389
R9090 VSS.n148 VSS.n147 0.249389
R9091 VSS.n1974 VSS.n1973 0.249389
R9092 VSS.n1844 VSS.n1843 0.249389
R9093 VSS.n326 VSS.n325 0.248689
R9094 VSS.n2654 VSS.n2653 0.248689
R9095 VSS.n1850 VSS 0.243833
R9096 VSS.n1847 VSS 0.243833
R9097 VSS VSS.n2858 0.243833
R9098 VSS VSS.n2863 0.243833
R9099 VSS VSS.n2869 0.243833
R9100 VSS.n2888 VSS 0.243833
R9101 VSS VSS.n2870 0.243833
R9102 VSS.n2873 VSS 0.243833
R9103 VSS.n2883 VSS 0.243833
R9104 VSS.n2893 VSS 0.243833
R9105 VSS VSS.n1114 0.243833
R9106 VSS VSS.n1120 0.243833
R9107 VSS VSS.n1109 0.243833
R9108 VSS.n1139 VSS 0.243833
R9109 VSS VSS.n1121 0.243833
R9110 VSS.n1124 VSS 0.243833
R9111 VSS.n1134 VSS 0.243833
R9112 VSS.n1144 VSS 0.243833
R9113 VSS.n1915 VSS 0.243833
R9114 VSS VSS.n1901 0.243833
R9115 VSS.n1899 VSS 0.243833
R9116 VSS VSS.n1894 0.243833
R9117 VSS VSS.n1906 0.243833
R9118 VSS VSS.n170 0.243833
R9119 VSS.n139 VSS 0.243833
R9120 VSS VSS.n116 0.243833
R9121 VSS VSS.n155 0.243833
R9122 VSS.n153 VSS 0.243833
R9123 VSS VSS.n148 0.243833
R9124 VSS VSS.n160 0.243833
R9125 VSS VSS.n161 0.243833
R9126 VSS VSS.n1032 0.243833
R9127 VSS VSS.n1981 0.243833
R9128 VSS.n1979 VSS 0.243833
R9129 VSS VSS.n1974 0.243833
R9130 VSS VSS.n1986 0.243833
R9131 VSS VSS.n1990 0.243833
R9132 VSS.n1966 VSS 0.243833
R9133 VSS.n1040 VSS 0.243833
R9134 VSS.n1954 VSS 0.243833
R9135 VSS.n1886 VSS 0.243833
R9136 VSS.n1429 VSS 0.243833
R9137 VSS.n1432 VSS 0.243833
R9138 VSS VSS.n1837 0.243833
R9139 VSS.n1825 VSS 0.243833
R9140 VSS.n1843 VSS 0.243833
R9141 VSS VSS.n1827 0.243833
R9142 VSS VSS.n1828 0.243833
R9143 VSS.n2531 VSS.n2530 0.238749
R9144 VSS.n2572 VSS.n2571 0.238749
R9145 VSS.n2086 VSS.n2085 0.237
R9146 VSS.n1224 VSS.n1220 0.237
R9147 VSS.n2533 VSS.n2532 0.236264
R9148 VSS.n1849 VSS.n1815 0.236056
R9149 VSS.n1846 VSS.n1845 0.236056
R9150 VSS.n1861 VSS.n1860 0.236056
R9151 VSS.n1857 VSS.n1856 0.236056
R9152 VSS.n2857 VSS.n2856 0.236056
R9153 VSS.n2860 VSS.n2859 0.236056
R9154 VSS.n2864 VSS.n2862 0.236056
R9155 VSS.n2876 VSS.n2875 0.236056
R9156 VSS.n2887 VSS.n2850 0.236056
R9157 VSS.n2872 VSS.n2871 0.236056
R9158 VSS.n2882 VSS.n2881 0.236056
R9159 VSS.n2892 VSS.n2891 0.236056
R9160 VSS.n2897 VSS.n2896 0.236056
R9161 VSS.n1115 VSS.n1113 0.236056
R9162 VSS.n1127 VSS.n1126 0.236056
R9163 VSS.n1111 VSS.n1110 0.236056
R9164 VSS.n2901 VSS.n7 0.236056
R9165 VSS.n1138 VSS.n1105 0.236056
R9166 VSS.n1123 VSS.n1122 0.236056
R9167 VSS.n1133 VSS.n1132 0.236056
R9168 VSS.n1143 VSS.n1142 0.236056
R9169 VSS.n1153 VSS.n1152 0.236056
R9170 VSS.n1902 VSS.n1900 0.236056
R9171 VSS.n1898 VSS.n1427 0.236056
R9172 VSS.n1895 VSS.n1426 0.236056
R9173 VSS.n1908 VSS.n1907 0.236056
R9174 VSS.n173 VSS.n172 0.236056
R9175 VSS.n129 VSS.n123 0.236056
R9176 VSS.n138 VSS.n118 0.236056
R9177 VSS.n145 VSS.n144 0.236056
R9178 VSS.n156 VSS.n154 0.236056
R9179 VSS.n152 VSS.n113 0.236056
R9180 VSS.n149 VSS.n112 0.236056
R9181 VSS.n182 VSS.n181 0.236056
R9182 VSS.n178 VSS.n177 0.236056
R9183 VSS.n1982 VSS.n1980 0.236056
R9184 VSS.n1978 VSS.n1038 0.236056
R9185 VSS.n1975 VSS.n1037 0.236056
R9186 VSS.n1987 VSS.n1035 0.236056
R9187 VSS.n1991 VSS.n1028 0.236056
R9188 VSS.n1965 VSS.n1042 0.236056
R9189 VSS.n1972 VSS.n1971 0.236056
R9190 VSS.n1960 VSS.n1959 0.236056
R9191 VSS.n1956 VSS.n1955 0.236056
R9192 VSS.n1885 VSS.n1431 0.236056
R9193 VSS.n1892 VSS.n1891 0.236056
R9194 VSS.n1880 VSS.n1879 0.236056
R9195 VSS.n1876 VSS.n1433 0.236056
R9196 VSS.n1838 VSS.n1826 0.236056
R9197 VSS.n1824 VSS.n1818 0.236056
R9198 VSS.n1842 VSS.n1819 0.236056
R9199 VSS.n1834 VSS.n1833 0.236056
R9200 VSS.n1830 VSS.n20 0.236056
R9201 VSS.n2098 VSS.n2089 0.236043
R9202 VSS.n1253 VSS.n1249 0.236043
R9203 VSS.n2439 VSS.n2438 0.2355
R9204 VSS.n1303 VSS.n1302 0.2355
R9205 VSS.n1944 VSS.n1943 0.234543
R9206 VSS.n2165 VSS 0.233577
R9207 VSS VSS.n2189 0.233577
R9208 VSS.n2194 VSS 0.233577
R9209 VSS.n2125 VSS 0.233577
R9210 VSS.n1307 VSS 0.233577
R9211 VSS VSS.n1333 0.233577
R9212 VSS.n1338 VSS 0.233577
R9213 VSS.n1357 VSS 0.233577
R9214 VSS VSS.n1264 0.233577
R9215 VSS VSS.n1934 0.233577
R9216 VSS.n1931 VSS 0.233577
R9217 VSS.n1397 VSS 0.233577
R9218 VSS.n1210 VSS 0.233577
R9219 VSS.n1192 VSS 0.233577
R9220 VSS VSS.n1379 0.233577
R9221 VSS.n1311 VSS 0.233577
R9222 VSS VSS.n2128 0.233577
R9223 VSS.n2171 VSS 0.233577
R9224 VSS VSS.n531 0.233577
R9225 VSS.n2072 VSS 0.233577
R9226 VSS VSS.n2049 0.233577
R9227 VSS VSS.n1807 0.233577
R9228 VSS.n2535 VSS.n2534 0.233545
R9229 VSS.n2578 VSS.n2575 0.233545
R9230 VSS.n130 VSS 0.2305
R9231 VSS.n365 VSS.n357 0.229074
R9232 VSS.n325 VSS.n303 0.229074
R9233 VSS.n2516 VSS.n2515 0.229074
R9234 VSS.n2761 VSS.n2760 0.229074
R9235 VSS.n2693 VSS.n2685 0.229074
R9236 VSS.n2653 VSS.n2631 0.229074
R9237 VSS.n220 VSS.n99 0.229074
R9238 VSS.n2041 VSS 0.2255
R9239 VSS.n1848 VSS.n1847 0.221611
R9240 VSS.n2869 VSS.n2868 0.221611
R9241 VSS.n1120 VSS.n1119 0.221611
R9242 VSS VSS.n2900 0.221611
R9243 VSS.n1041 VSS.n1040 0.221611
R9244 VSS.n1430 VSS.n1429 0.221611
R9245 VSS.n2437 VSS 0.219469
R9246 VSS VSS.n2087 0.219469
R9247 VSS VSS.n2454 0.219469
R9248 VSS.n1219 VSS 0.219469
R9249 VSS VSS.n1875 0.219205
R9250 VSS VSS.n2088 0.218541
R9251 VSS.n1248 VSS 0.218541
R9252 VSS VSS.n1068 0.218541
R9253 VSS VSS.n125 0.217167
R9254 VSS.n2532 VSS.n2531 0.214098
R9255 VSS.n2573 VSS.n2572 0.214098
R9256 VSS.n117 VSS.n115 0.212722
R9257 VSS.n133 VSS.n119 0.21207
R9258 VSS.n366 VSS.n365 0.2105
R9259 VSS.n2515 VSS.n237 0.2105
R9260 VSS.n2760 VSS.n76 0.2105
R9261 VSS.n2694 VSS.n2693 0.2105
R9262 VSS.n352 VSS.n347 0.210483
R9263 VSS.n313 VSS.n290 0.210483
R9264 VSS.n248 VSS.n247 0.210483
R9265 VSS.n1173 VSS.n223 0.210483
R9266 VSS.n2680 VSS.n2675 0.210483
R9267 VSS.n2641 VSS.n2618 0.210483
R9268 VSS.n87 VSS.n86 0.210483
R9269 VSS.n1100 VSS.n1092 0.20138
R9270 VSS.n194 VSS.n193 0.20138
R9271 VSS.n2168 VSS.n2166 0.199786
R9272 VSS.n2078 VSS.n2077 0.199786
R9273 VSS.n516 VSS.n512 0.199786
R9274 VSS.n2188 VSS.n2143 0.199786
R9275 VSS.n2195 VSS.n2137 0.199786
R9276 VSS.n1308 VSS.n1298 0.199786
R9277 VSS.n1332 VSS.n1278 0.199786
R9278 VSS.n1345 VSS.n1344 0.199786
R9279 VSS.n1259 VSS.n1245 0.199786
R9280 VSS.n1364 VSS.n1363 0.199786
R9281 VSS.n1217 VSS.n1208 0.199786
R9282 VSS.n1929 VSS.n1417 0.199786
R9283 VSS.n1416 VSS.n1415 0.199786
R9284 VSS.n1404 VSS.n1403 0.199786
R9285 VSS.n1193 VSS.n1187 0.199786
R9286 VSS.n1376 VSS.n1211 0.199786
R9287 VSS.n1314 VSS.n1313 0.199786
R9288 VSS.n2123 VSS.n513 0.199786
R9289 VSS.n2074 VSS.n2073 0.199786
R9290 VSS.n2174 VSS.n2173 0.199786
R9291 VSS.n2048 VSS.n555 0.199786
R9292 VSS.n1810 VSS.n1434 0.199786
R9293 VSS.n2826 VSS.n2825 0.196456
R9294 VSS.n2566 VSS.n2565 0.189389
R9295 VSS.n374 VSS.n373 0.189389
R9296 VSS.n321 VSS.n310 0.189389
R9297 VSS.n370 VSS.n369 0.189389
R9298 VSS.n318 VSS.n317 0.189389
R9299 VSS.n2511 VSS.n2509 0.189389
R9300 VSS.n2506 VSS.n2505 0.189389
R9301 VSS.n2546 VSS.n2544 0.189389
R9302 VSS.n2756 VSS.n2754 0.189389
R9303 VSS.n2649 VSS.n2638 0.189389
R9304 VSS.n2698 VSS.n2697 0.189389
R9305 VSS.n2702 VSS.n2701 0.189389
R9306 VSS.n2646 VSS.n2645 0.189389
R9307 VSS.n2751 VSS.n2750 0.189389
R9308 VSS.n359 VSS.n357 0.18928
R9309 VSS.n305 VSS.n303 0.18928
R9310 VSS.n2517 VSS.n2516 0.18928
R9311 VSS.n2762 VSS.n2761 0.18928
R9312 VSS.n2687 VSS.n2685 0.18928
R9313 VSS.n2633 VSS.n2631 0.18928
R9314 VSS.n214 VSS.n99 0.18928
R9315 VSS.n1266 VSS.n1265 0.1805
R9316 VSS.n217 VSS 0.178278
R9317 VSS VSS.n353 0.178278
R9318 VSS.n322 VSS 0.178278
R9319 VSS.n362 VSS 0.178278
R9320 VSS VSS.n314 0.178278
R9321 VSS VSS.n241 0.178278
R9322 VSS.n246 VSS 0.178278
R9323 VSS.n1171 VSS 0.178278
R9324 VSS VSS.n80 0.178278
R9325 VSS.n2650 VSS 0.178278
R9326 VSS.n2690 VSS 0.178278
R9327 VSS VSS.n2681 0.178278
R9328 VSS VSS.n2642 0.178278
R9329 VSS.n85 VSS 0.178278
R9330 VSS.n329 VSS.n300 0.177167
R9331 VSS.n272 VSS.n270 0.177167
R9332 VSS.n2495 VSS.n265 0.177167
R9333 VSS.n2477 VSS.n295 0.177167
R9334 VSS.n2528 VSS.n2527 0.177167
R9335 VSS.n2540 VSS.n2539 0.177167
R9336 VSS.n1159 VSS.n1099 0.177167
R9337 VSS.n2773 VSS.n2772 0.177167
R9338 VSS.n2657 VSS.n2628 0.177167
R9339 VSS.n2603 VSS.n2601 0.177167
R9340 VSS.n2719 VSS.n2623 0.177167
R9341 VSS.n2738 VSS.n2737 0.177167
R9342 VSS.n2577 VSS.n92 0.177167
R9343 VSS.n204 VSS.n203 0.177167
R9344 VSS.n176 VSS.n175 0.176722
R9345 VSS.n1868 VSS.n1867 0.175143
R9346 VSS.n2456 VSS 0.175034
R9347 VSS.n2451 VSS 0.175034
R9348 VSS.n558 VSS.n557 0.173341
R9349 VSS.n2032 VSS 0.172842
R9350 VSS.n2112 VSS.n521 0.170294
R9351 VSS.n376 VSS.n350 0.168962
R9352 VSS.n368 VSS.n367 0.168962
R9353 VSS.n309 VSS.n301 0.168962
R9354 VSS.n316 VSS.n293 0.168962
R9355 VSS.n2512 VSS.n239 0.168962
R9356 VSS.n2504 VSS.n2503 0.168962
R9357 VSS.n2547 VSS.n225 0.168962
R9358 VSS.n2757 VSS.n78 0.168962
R9359 VSS.n2696 VSS.n2695 0.168962
R9360 VSS.n2637 VSS.n2629 0.168962
R9361 VSS.n2704 VSS.n2678 0.168962
R9362 VSS.n2644 VSS.n2621 0.168962
R9363 VSS.n2749 VSS.n2748 0.168962
R9364 VSS.n2564 VSS.n2563 0.168962
R9365 VSS.n1369 VSS.n1368 0.168438
R9366 VSS.n2431 VSS.n61 0.167808
R9367 VSS.n197 VSS.n196 0.166424
R9368 VSS.n1158 VSS.n1157 0.166424
R9369 VSS.n126 VSS.n122 0.166056
R9370 VSS.n363 VSS.n358 0.1655
R9371 VSS.n323 VSS.n304 0.1655
R9372 VSS.n238 VSS.n236 0.1655
R9373 VSS.n77 VSS.n75 0.1655
R9374 VSS.n2691 VSS.n2686 0.1655
R9375 VSS.n2651 VSS.n2632 0.1655
R9376 VSS.n218 VSS.n100 0.1655
R9377 VSS.n2203 VSS.n2202 0.1565
R9378 VSS.n2156 VSS.n2155 0.1565
R9379 VSS.n1351 VSS.n1349 0.1565
R9380 VSS.n1291 VSS.n1290 0.1565
R9381 VSS.n1410 VSS.n1408 0.1565
R9382 VSS.n1203 VSS.n1202 0.1565
R9383 VSS.n552 VSS.n551 0.1565
R9384 VSS.n1855 VSS.n1815 0.155275
R9385 VSS.n2862 VSS.n2854 0.155275
R9386 VSS.n1113 VSS.n1112 0.155275
R9387 VSS.n134 VSS.n118 0.155275
R9388 VSS.n1961 VSS.n1042 0.155275
R9389 VSS.n1881 VSS.n1431 0.155275
R9390 VSS.n2154 VSS.n2153 0.154786
R9391 VSS.n2201 VSS.n2200 0.154786
R9392 VSS.n1289 VSS.n1288 0.154786
R9393 VSS.n1352 VSS.n1270 0.154786
R9394 VSS.n1411 VSS.n1080 0.154786
R9395 VSS.n1204 VSS.n1189 0.154786
R9396 VSS.n2054 VSS.n535 0.154786
R9397 VSS.n1371 VSS.n1370 0.152665
R9398 VSS.n2561 VSS.n220 0.151747
R9399 VSS.n2210 VSS.n508 0.1505
R9400 VSS.n1151 VSS.n1150 0.149389
R9401 VSS VSS.n1044 0.147167
R9402 VSS.n1059 VSS 0.147167
R9403 VSS.n1055 VSS 0.147167
R9404 VSS.n1334 VSS.n1276 0.147038
R9405 VSS.n2029 VSS 0.144346
R9406 VSS.n2574 VSS.n2573 0.140703
R9407 VSS.n2537 VSS.n2534 0.138684
R9408 VSS.n2580 VSS.n2575 0.138684
R9409 VSS.n2046 VSS.n2045 0.137808
R9410 VSS.n2406 VSS.n2405 0.1355
R9411 VSS.n2407 VSS.n2406 0.1355
R9412 VSS.n2407 VSS.n403 0.1355
R9413 VSS.n2413 VSS.n403 0.1355
R9414 VSS.n2414 VSS.n2413 0.1355
R9415 VSS.n2415 VSS.n2414 0.1355
R9416 VSS.n2415 VSS.n399 0.1355
R9417 VSS.n2421 VSS.n399 0.1355
R9418 VSS.n2422 VSS.n2421 0.1355
R9419 VSS.n2423 VSS.n2422 0.1355
R9420 VSS.n2423 VSS.n395 0.1355
R9421 VSS.n2429 VSS.n395 0.1355
R9422 VSS.n2430 VSS.n2429 0.1355
R9423 VSS.n2431 VSS.n2430 0.1355
R9424 VSS.n2218 VSS.n2217 0.1355
R9425 VSS.n2218 VSS.n498 0.1355
R9426 VSS.n2224 VSS.n498 0.1355
R9427 VSS.n2225 VSS.n2224 0.1355
R9428 VSS.n2226 VSS.n2225 0.1355
R9429 VSS.n2226 VSS.n494 0.1355
R9430 VSS.n2232 VSS.n494 0.1355
R9431 VSS.n2233 VSS.n2232 0.1355
R9432 VSS.n2234 VSS.n2233 0.1355
R9433 VSS.n2234 VSS.n490 0.1355
R9434 VSS.n2240 VSS.n490 0.1355
R9435 VSS.n2241 VSS.n2240 0.1355
R9436 VSS.n2242 VSS.n2241 0.1355
R9437 VSS.n2242 VSS.n486 0.1355
R9438 VSS.n2248 VSS.n486 0.1355
R9439 VSS.n2249 VSS.n2248 0.1355
R9440 VSS.n2250 VSS.n2249 0.1355
R9441 VSS.n2250 VSS.n482 0.1355
R9442 VSS.n2256 VSS.n482 0.1355
R9443 VSS.n2257 VSS.n2256 0.1355
R9444 VSS.n2258 VSS.n2257 0.1355
R9445 VSS.n2258 VSS.n478 0.1355
R9446 VSS.n2264 VSS.n478 0.1355
R9447 VSS.n2265 VSS.n2264 0.1355
R9448 VSS.n2266 VSS.n2265 0.1355
R9449 VSS.n2266 VSS.n474 0.1355
R9450 VSS.n2272 VSS.n474 0.1355
R9451 VSS.n2273 VSS.n2272 0.1355
R9452 VSS.n2274 VSS.n2273 0.1355
R9453 VSS.n2274 VSS.n470 0.1355
R9454 VSS.n2280 VSS.n470 0.1355
R9455 VSS.n2281 VSS.n2280 0.1355
R9456 VSS.n2282 VSS.n2281 0.1355
R9457 VSS.n2282 VSS.n466 0.1355
R9458 VSS.n2288 VSS.n466 0.1355
R9459 VSS.n2289 VSS.n2288 0.1355
R9460 VSS.n2290 VSS.n2289 0.1355
R9461 VSS.n2290 VSS.n462 0.1355
R9462 VSS.n2296 VSS.n462 0.1355
R9463 VSS.n2297 VSS.n2296 0.1355
R9464 VSS.n2298 VSS.n2297 0.1355
R9465 VSS.n2298 VSS.n458 0.1355
R9466 VSS.n2304 VSS.n458 0.1355
R9467 VSS.n2305 VSS.n2304 0.1355
R9468 VSS.n2306 VSS.n2305 0.1355
R9469 VSS.n2306 VSS.n454 0.1355
R9470 VSS.n2312 VSS.n454 0.1355
R9471 VSS.n2313 VSS.n2312 0.1355
R9472 VSS.n2314 VSS.n2313 0.1355
R9473 VSS.n2314 VSS.n450 0.1355
R9474 VSS.n2320 VSS.n450 0.1355
R9475 VSS.n2321 VSS.n2320 0.1355
R9476 VSS.n2322 VSS.n2321 0.1355
R9477 VSS.n2322 VSS.n446 0.1355
R9478 VSS.n2328 VSS.n446 0.1355
R9479 VSS.n2329 VSS.n2328 0.1355
R9480 VSS.n2330 VSS.n2329 0.1355
R9481 VSS.n2330 VSS.n442 0.1355
R9482 VSS.n2336 VSS.n442 0.1355
R9483 VSS.n2337 VSS.n2336 0.1355
R9484 VSS.n2338 VSS.n2337 0.1355
R9485 VSS.n2338 VSS.n438 0.1355
R9486 VSS.n2344 VSS.n438 0.1355
R9487 VSS.n2345 VSS.n2344 0.1355
R9488 VSS.n2346 VSS.n2345 0.1355
R9489 VSS.n2346 VSS.n434 0.1355
R9490 VSS.n2352 VSS.n434 0.1355
R9491 VSS.n2353 VSS.n2352 0.1355
R9492 VSS.n2354 VSS.n2353 0.1355
R9493 VSS.n2354 VSS.n430 0.1355
R9494 VSS.n2360 VSS.n430 0.1355
R9495 VSS.n2361 VSS.n2360 0.1355
R9496 VSS.n2362 VSS.n2361 0.1355
R9497 VSS.n2362 VSS.n426 0.1355
R9498 VSS.n2368 VSS.n426 0.1355
R9499 VSS.n2369 VSS.n2368 0.1355
R9500 VSS.n2373 VSS.n2369 0.1355
R9501 VSS.n909 VSS.n689 0.1355
R9502 VSS.n909 VSS.n908 0.1355
R9503 VSS.n908 VSS.n907 0.1355
R9504 VSS.n907 VSS.n693 0.1355
R9505 VSS.n901 VSS.n693 0.1355
R9506 VSS.n901 VSS.n900 0.1355
R9507 VSS.n900 VSS.n899 0.1355
R9508 VSS.n899 VSS.n697 0.1355
R9509 VSS.n893 VSS.n697 0.1355
R9510 VSS.n893 VSS.n892 0.1355
R9511 VSS.n892 VSS.n891 0.1355
R9512 VSS.n891 VSS.n701 0.1355
R9513 VSS.n885 VSS.n701 0.1355
R9514 VSS.n885 VSS.n884 0.1355
R9515 VSS.n884 VSS.n883 0.1355
R9516 VSS.n883 VSS.n705 0.1355
R9517 VSS.n877 VSS.n705 0.1355
R9518 VSS.n877 VSS.n876 0.1355
R9519 VSS.n876 VSS.n875 0.1355
R9520 VSS.n875 VSS.n709 0.1355
R9521 VSS.n869 VSS.n709 0.1355
R9522 VSS.n869 VSS.n868 0.1355
R9523 VSS.n868 VSS.n867 0.1355
R9524 VSS.n867 VSS.n713 0.1355
R9525 VSS.n861 VSS.n713 0.1355
R9526 VSS.n861 VSS.n860 0.1355
R9527 VSS.n860 VSS.n859 0.1355
R9528 VSS.n859 VSS.n717 0.1355
R9529 VSS.n853 VSS.n717 0.1355
R9530 VSS.n853 VSS.n852 0.1355
R9531 VSS.n852 VSS.n851 0.1355
R9532 VSS.n851 VSS.n721 0.1355
R9533 VSS.n845 VSS.n721 0.1355
R9534 VSS.n845 VSS.n844 0.1355
R9535 VSS.n844 VSS.n843 0.1355
R9536 VSS.n843 VSS.n725 0.1355
R9537 VSS.n837 VSS.n725 0.1355
R9538 VSS.n837 VSS.n836 0.1355
R9539 VSS.n836 VSS.n835 0.1355
R9540 VSS.n835 VSS.n729 0.1355
R9541 VSS.n829 VSS.n729 0.1355
R9542 VSS.n829 VSS.n828 0.1355
R9543 VSS.n828 VSS.n827 0.1355
R9544 VSS.n827 VSS.n733 0.1355
R9545 VSS.n821 VSS.n733 0.1355
R9546 VSS.n821 VSS.n820 0.1355
R9547 VSS.n820 VSS.n819 0.1355
R9548 VSS.n819 VSS.n737 0.1355
R9549 VSS.n813 VSS.n737 0.1355
R9550 VSS.n813 VSS.n812 0.1355
R9551 VSS.n812 VSS.n811 0.1355
R9552 VSS.n811 VSS.n741 0.1355
R9553 VSS.n805 VSS.n741 0.1355
R9554 VSS.n805 VSS.n804 0.1355
R9555 VSS.n804 VSS.n803 0.1355
R9556 VSS.n803 VSS.n745 0.1355
R9557 VSS.n797 VSS.n745 0.1355
R9558 VSS.n797 VSS.n796 0.1355
R9559 VSS.n796 VSS.n795 0.1355
R9560 VSS.n795 VSS.n749 0.1355
R9561 VSS.n789 VSS.n749 0.1355
R9562 VSS.n1018 VSS.n587 0.1355
R9563 VSS.n1013 VSS.n587 0.1355
R9564 VSS.n1013 VSS.n1012 0.1355
R9565 VSS.n1012 VSS.n1011 0.1355
R9566 VSS.n1011 VSS.n596 0.1355
R9567 VSS.n1005 VSS.n596 0.1355
R9568 VSS.n1005 VSS.n1004 0.1355
R9569 VSS.n1004 VSS.n1003 0.1355
R9570 VSS.n1003 VSS.n598 0.1355
R9571 VSS.n600 VSS.n598 0.1355
R9572 VSS.n603 VSS.n600 0.1355
R9573 VSS.n994 VSS.n603 0.1355
R9574 VSS.n994 VSS.n993 0.1355
R9575 VSS.n993 VSS.n992 0.1355
R9576 VSS.n992 VSS.n604 0.1355
R9577 VSS.n986 VSS.n604 0.1355
R9578 VSS.n986 VSS.n985 0.1355
R9579 VSS.n985 VSS.n984 0.1355
R9580 VSS.n984 VSS.n608 0.1355
R9581 VSS.n618 VSS.n608 0.1355
R9582 VSS.n619 VSS.n618 0.1355
R9583 VSS.n619 VSS.n615 0.1355
R9584 VSS.n625 VSS.n615 0.1355
R9585 VSS.n626 VSS.n625 0.1355
R9586 VSS.n627 VSS.n626 0.1355
R9587 VSS.n627 VSS.n613 0.1355
R9588 VSS.n633 VSS.n613 0.1355
R9589 VSS.n634 VSS.n633 0.1355
R9590 VSS.n978 VSS.n634 0.1355
R9591 VSS.n978 VSS.n977 0.1355
R9592 VSS.n977 VSS.n976 0.1355
R9593 VSS.n976 VSS.n635 0.1355
R9594 VSS.n970 VSS.n635 0.1355
R9595 VSS.n970 VSS.n969 0.1355
R9596 VSS.n969 VSS.n968 0.1355
R9597 VSS.n968 VSS.n639 0.1355
R9598 VSS.n962 VSS.n639 0.1355
R9599 VSS.n962 VSS.n961 0.1355
R9600 VSS.n961 VSS.n960 0.1355
R9601 VSS.n960 VSS.n643 0.1355
R9602 VSS.n954 VSS.n643 0.1355
R9603 VSS.n954 VSS.n953 0.1355
R9604 VSS.n953 VSS.n952 0.1355
R9605 VSS.n952 VSS.n647 0.1355
R9606 VSS.n946 VSS.n647 0.1355
R9607 VSS.n946 VSS.n945 0.1355
R9608 VSS.n945 VSS.n944 0.1355
R9609 VSS.n944 VSS.n651 0.1355
R9610 VSS.n938 VSS.n651 0.1355
R9611 VSS.n938 VSS.n937 0.1355
R9612 VSS.n937 VSS.n936 0.1355
R9613 VSS.n936 VSS.n655 0.1355
R9614 VSS.n930 VSS.n655 0.1355
R9615 VSS.n930 VSS.n929 0.1355
R9616 VSS.n1592 VSS.n1458 0.1355
R9617 VSS.n1592 VSS.n1591 0.1355
R9618 VSS.n1591 VSS.n1590 0.1355
R9619 VSS.n1590 VSS.n1462 0.1355
R9620 VSS.n1584 VSS.n1462 0.1355
R9621 VSS.n1584 VSS.n1583 0.1355
R9622 VSS.n1583 VSS.n1582 0.1355
R9623 VSS.n1582 VSS.n1466 0.1355
R9624 VSS.n1576 VSS.n1466 0.1355
R9625 VSS.n1576 VSS.n1575 0.1355
R9626 VSS.n1575 VSS.n1574 0.1355
R9627 VSS.n1574 VSS.n1470 0.1355
R9628 VSS.n1568 VSS.n1470 0.1355
R9629 VSS.n1568 VSS.n1567 0.1355
R9630 VSS.n1567 VSS.n1566 0.1355
R9631 VSS.n1566 VSS.n1474 0.1355
R9632 VSS.n1560 VSS.n1474 0.1355
R9633 VSS.n1560 VSS.n1559 0.1355
R9634 VSS.n1559 VSS.n1558 0.1355
R9635 VSS.n1558 VSS.n1478 0.1355
R9636 VSS.n1552 VSS.n1478 0.1355
R9637 VSS.n1552 VSS.n1551 0.1355
R9638 VSS.n1551 VSS.n1550 0.1355
R9639 VSS.n1550 VSS.n1482 0.1355
R9640 VSS.n1544 VSS.n1482 0.1355
R9641 VSS.n1544 VSS.n1543 0.1355
R9642 VSS.n1543 VSS.n1542 0.1355
R9643 VSS.n1542 VSS.n1486 0.1355
R9644 VSS.n1536 VSS.n1486 0.1355
R9645 VSS.n1536 VSS.n1535 0.1355
R9646 VSS.n1535 VSS.n1534 0.1355
R9647 VSS.n1534 VSS.n1490 0.1355
R9648 VSS.n1528 VSS.n1490 0.1355
R9649 VSS.n1528 VSS.n1527 0.1355
R9650 VSS.n1527 VSS.n1526 0.1355
R9651 VSS.n1526 VSS.n1494 0.1355
R9652 VSS.n1520 VSS.n1494 0.1355
R9653 VSS.n1520 VSS.n1519 0.1355
R9654 VSS.n1519 VSS.n1518 0.1355
R9655 VSS.n1518 VSS.n1498 0.1355
R9656 VSS.n1512 VSS.n1498 0.1355
R9657 VSS.n1512 VSS.n1511 0.1355
R9658 VSS.n1511 VSS.n1510 0.1355
R9659 VSS.n1510 VSS.n1502 0.1355
R9660 VSS.n1504 VSS.n1502 0.1355
R9661 VSS.n1504 VSS.n570 0.1355
R9662 VSS.n2023 VSS.n570 0.1355
R9663 VSS.n2023 VSS.n2022 0.1355
R9664 VSS.n2022 VSS.n2021 0.1355
R9665 VSS.n2021 VSS.n571 0.1355
R9666 VSS.n2015 VSS.n571 0.1355
R9667 VSS.n2015 VSS.n2014 0.1355
R9668 VSS.n1632 VSS.n1631 0.1355
R9669 VSS.n1632 VSS.n1626 0.1355
R9670 VSS.n1638 VSS.n1626 0.1355
R9671 VSS.n1639 VSS.n1638 0.1355
R9672 VSS.n1640 VSS.n1639 0.1355
R9673 VSS.n1640 VSS.n1624 0.1355
R9674 VSS.n1646 VSS.n1624 0.1355
R9675 VSS.n1647 VSS.n1646 0.1355
R9676 VSS.n1648 VSS.n1647 0.1355
R9677 VSS.n1648 VSS.n1622 0.1355
R9678 VSS.n1654 VSS.n1622 0.1355
R9679 VSS.n1655 VSS.n1654 0.1355
R9680 VSS.n1656 VSS.n1655 0.1355
R9681 VSS.n1656 VSS.n1620 0.1355
R9682 VSS.n1662 VSS.n1620 0.1355
R9683 VSS.n1663 VSS.n1662 0.1355
R9684 VSS.n1664 VSS.n1663 0.1355
R9685 VSS.n1664 VSS.n1618 0.1355
R9686 VSS.n1670 VSS.n1618 0.1355
R9687 VSS.n1671 VSS.n1670 0.1355
R9688 VSS.n1672 VSS.n1671 0.1355
R9689 VSS.n1672 VSS.n1616 0.1355
R9690 VSS.n1678 VSS.n1616 0.1355
R9691 VSS.n1679 VSS.n1678 0.1355
R9692 VSS.n1680 VSS.n1679 0.1355
R9693 VSS.n1680 VSS.n1614 0.1355
R9694 VSS.n1686 VSS.n1614 0.1355
R9695 VSS.n1687 VSS.n1686 0.1355
R9696 VSS.n1688 VSS.n1687 0.1355
R9697 VSS.n1688 VSS.n1612 0.1355
R9698 VSS.n1694 VSS.n1612 0.1355
R9699 VSS.n1695 VSS.n1694 0.1355
R9700 VSS.n1696 VSS.n1695 0.1355
R9701 VSS.n1696 VSS.n1610 0.1355
R9702 VSS.n1702 VSS.n1610 0.1355
R9703 VSS.n1703 VSS.n1702 0.1355
R9704 VSS.n1704 VSS.n1703 0.1355
R9705 VSS.n1704 VSS.n1608 0.1355
R9706 VSS.n1710 VSS.n1608 0.1355
R9707 VSS.n1711 VSS.n1710 0.1355
R9708 VSS.n1712 VSS.n1711 0.1355
R9709 VSS.n1712 VSS.n1606 0.1355
R9710 VSS.n1718 VSS.n1606 0.1355
R9711 VSS.n1719 VSS.n1718 0.1355
R9712 VSS.n1720 VSS.n1719 0.1355
R9713 VSS.n1720 VSS.n1604 0.1355
R9714 VSS.n1726 VSS.n1604 0.1355
R9715 VSS.n1727 VSS.n1726 0.1355
R9716 VSS.n1728 VSS.n1727 0.1355
R9717 VSS.n1728 VSS.n1602 0.1355
R9718 VSS.n1734 VSS.n1602 0.1355
R9719 VSS.n1735 VSS.n1734 0.1355
R9720 VSS.n1736 VSS.n1735 0.1355
R9721 VSS.n1736 VSS.n1600 0.1355
R9722 VSS.n1741 VSS.n1600 0.1355
R9723 VSS.n2089 VSS 0.13409
R9724 VSS.n1249 VSS 0.13409
R9725 VSS.n1944 VSS 0.13409
R9726 VSS.n2438 VSS 0.133132
R9727 VSS VSS.n2086 0.133132
R9728 VSS.n1302 VSS 0.133132
R9729 VSS.n1220 VSS 0.133132
R9730 VSS.n1180 VSS.n1092 0.132897
R9731 VSS.n193 VSS.n189 0.132897
R9732 VSS VSS.n1814 0.132722
R9733 VSS.n1631 VSS.n1630 0.132038
R9734 VSS.n132 VSS.n120 0.129738
R9735 VSS.n2014 VSS.n2013 0.126287
R9736 VSS VSS.n2031 0.126081
R9737 VSS.n2211 VSS.n507 0.122388
R9738 VSS VSS.n1371 0.116479
R9739 VSS VSS.n521 0.116479
R9740 VSS.n2832 VSS.n2831 0.116432
R9741 VSS.n2452 VSS.n2451 0.116021
R9742 VSS.n1368 VSS 0.115552
R9743 VSS.n1918 VSS 0.115552
R9744 VSS VSS.n520 0.115552
R9745 VSS.n2044 VSS.n2043 0.115394
R9746 VSS.n789 VSS.n788 0.113655
R9747 VSS.n681 VSS.n680 0.113597
R9748 VSS.n2210 VSS.n2209 0.113577
R9749 VSS.n2500 VSS.n263 0.112682
R9750 VSS.n2745 VSS.n2594 0.112682
R9751 VSS.n1862 VSS.n1814 0.111611
R9752 VSS.n420 VSS.n388 0.109786
R9753 VSS.n2531 VSS.n229 0.109456
R9754 VSS.n2572 VSS.n68 0.109456
R9755 VSS.n2113 VSS.n520 0.106273
R9756 VSS.n165 VSS 0.103212
R9757 VSS.n1157 VSS.n1100 0.102619
R9758 VSS.n197 VSS.n194 0.102619
R9759 VSS.n2459 VSS.n2458 0.100143
R9760 VSS VSS.n2147 0.0997784
R9761 VSS VSS.n510 0.0997784
R9762 VSS VSS.n383 0.0997784
R9763 VSS.n2449 VSS 0.0997784
R9764 VSS VSS.n1282 0.0997784
R9765 VSS VSS.n1353 0.0997784
R9766 VSS VSS.n1240 0.0997784
R9767 VSS VSS.n1215 0.0997784
R9768 VSS VSS.n1412 0.0997784
R9769 VSS VSS.n1206 0.0997784
R9770 VSS VSS.n519 0.0997784
R9771 VSS VSS.n523 0.0997784
R9772 VSS VSS.n2065 0.0997784
R9773 VSS VSS.n1 0.0997784
R9774 VSS.n2455 VSS.n384 0.0972571
R9775 VSS.n392 VSS.n391 0.0951392
R9776 VSS.n528 VSS.n526 0.0951392
R9777 VSS.n1301 VSS.n385 0.0951392
R9778 VSS.n1223 VSS.n1222 0.0951392
R9779 VSS.n196 VSS.n195 0.0949444
R9780 VSS.n1160 VSS.n1158 0.0949444
R9781 VSS.n331 VSS.n330 0.0949444
R9782 VSS.n274 VSS.n273 0.0949444
R9783 VSS.n2497 VSS.n2496 0.0949444
R9784 VSS.n2479 VSS.n2478 0.0949444
R9785 VSS.n2530 VSS.n2529 0.0949444
R9786 VSS.n2536 VSS.n2535 0.0949444
R9787 VSS.n2571 VSS.n2570 0.0949444
R9788 VSS.n2659 VSS.n2658 0.0949444
R9789 VSS.n2605 VSS.n2604 0.0949444
R9790 VSS.n2721 VSS.n2720 0.0949444
R9791 VSS.n2742 VSS.n2741 0.0949444
R9792 VSS.n2579 VSS.n2578 0.0949444
R9793 VSS.n2100 VSS.n2099 0.0942113
R9794 VSS.n1252 VSS.n1251 0.0942113
R9795 VSS.n1945 VSS.n1070 0.0942113
R9796 VSS.n360 VSS.n358 0.0931962
R9797 VSS.n306 VSS.n304 0.0931962
R9798 VSS.n236 VSS.n235 0.0931962
R9799 VSS.n75 VSS.n74 0.0931962
R9800 VSS.n2688 VSS.n2686 0.0931962
R9801 VSS.n2634 VSS.n2632 0.0931962
R9802 VSS.n215 VSS.n100 0.0931962
R9803 VSS.n1919 VSS.n1917 0.0923557
R9804 VSS.n275 VSS.n271 0.0919876
R9805 VSS.n1161 VSS.n1100 0.0919876
R9806 VSS.n2606 VSS.n2602 0.0919876
R9807 VSS.n194 VSS.n106 0.0919876
R9808 VSS.n2130 VSS.n2129 0.0916538
R9809 VSS.n929 VSS.n928 0.0898504
R9810 VSS.n1863 VSS.n1862 0.0893889
R9811 VSS.n2032 VSS.n558 0.0883824
R9812 VSS.n2390 VSS.n420 0.0841129
R9813 VSS.n1812 VSS.n1 0.0830773
R9814 VSS.n1919 VSS.n1918 0.0812216
R9815 VSS.n130 VSS.n122 0.0805
R9816 VSS.n333 VSS.n332 0.079343
R9817 VSS.n276 VSS.n275 0.079343
R9818 VSS.n285 VSS.n264 0.079343
R9819 VSS.n342 VSS.n294 0.079343
R9820 VSS.n2526 VSS.n229 0.079343
R9821 VSS.n2538 VSS.n2537 0.079343
R9822 VSS.n1162 VSS.n1161 0.079343
R9823 VSS.n2771 VSS.n68 0.079343
R9824 VSS.n2661 VSS.n2660 0.079343
R9825 VSS.n2607 VSS.n2606 0.079343
R9826 VSS.n2670 VSS.n2622 0.079343
R9827 VSS.n2740 VSS.n2739 0.079343
R9828 VSS.n2581 VSS.n2580 0.079343
R9829 VSS.n205 VSS.n106 0.079343
R9830 VSS.n2471 VSS 0.0778554
R9831 VSS.n2489 VSS 0.0778554
R9832 VSS.n2484 VSS 0.0778554
R9833 VSS.n2466 VSS 0.0778554
R9834 VSS.n2518 VSS 0.0778554
R9835 VSS VSS.n249 0.0778554
R9836 VSS VSS.n1170 0.0778554
R9837 VSS.n2763 VSS 0.0778554
R9838 VSS.n2713 VSS 0.0778554
R9839 VSS.n2731 VSS 0.0778554
R9840 VSS.n2708 VSS 0.0778554
R9841 VSS.n2726 VSS 0.0778554
R9842 VSS VSS.n88 0.0778554
R9843 VSS VSS.n101 0.0778554
R9844 VSS.n1851 VSS.n1848 0.0746176
R9845 VSS.n2868 VSS.n2853 0.0746176
R9846 VSS.n1119 VSS.n1108 0.0746176
R9847 VSS.n140 VSS.n117 0.0746176
R9848 VSS.n1967 VSS.n1041 0.0746176
R9849 VSS.n1887 VSS.n1430 0.0746176
R9850 VSS.n2454 VSS.n2453 0.073799
R9851 VSS.n264 VSS.n262 0.072156
R9852 VSS.n2740 VSS.n2593 0.072156
R9853 VSS.n332 VSS.n328 0.0719368
R9854 VSS.n2660 VSS.n2656 0.0719368
R9855 VSS.n122 VSS.n121 0.0705
R9856 VSS.n2043 VSS 0.0703936
R9857 VSS.n2373 VSS.n2372 0.0695408
R9858 VSS.n2480 VSS.n294 0.0683965
R9859 VSS.n2722 VSS.n2622 0.0683965
R9860 VSS.n1921 VSS 0.0673041
R9861 VSS.n2114 VSS.n2113 0.0673041
R9862 VSS.n766 VSS.n506 0.0665432
R9863 VSS.n352 VSS.n348 0.0662692
R9864 VSS.n350 VSS.n349 0.0662692
R9865 VSS.n364 VSS.n363 0.0662692
R9866 VSS.n368 VSS.n356 0.0662692
R9867 VSS.n324 VSS.n323 0.0662692
R9868 VSS.n309 VSS.n302 0.0662692
R9869 VSS.n313 VSS.n291 0.0662692
R9870 VSS.n316 VSS.n292 0.0662692
R9871 VSS.n2514 VSS.n238 0.0662692
R9872 VSS.n2513 VSS.n2512 0.0662692
R9873 VSS.n247 VSS.n244 0.0662692
R9874 VSS.n2504 VSS.n243 0.0662692
R9875 VSS.n2549 VSS.n223 0.0662692
R9876 VSS.n2548 VSS.n2547 0.0662692
R9877 VSS.n2759 VSS.n77 0.0662692
R9878 VSS.n2758 VSS.n2757 0.0662692
R9879 VSS.n2692 VSS.n2691 0.0662692
R9880 VSS.n2696 VSS.n2684 0.0662692
R9881 VSS.n2652 VSS.n2651 0.0662692
R9882 VSS.n2637 VSS.n2630 0.0662692
R9883 VSS.n2680 VSS.n2676 0.0662692
R9884 VSS.n2678 VSS.n2677 0.0662692
R9885 VSS.n2641 VSS.n2619 0.0662692
R9886 VSS.n2644 VSS.n2620 0.0662692
R9887 VSS.n86 VSS.n83 0.0662692
R9888 VSS.n2749 VSS.n82 0.0662692
R9889 VSS.n219 VSS.n218 0.0662692
R9890 VSS.n2564 VSS.n98 0.0662692
R9891 VSS.n217 VSS.n216 0.0660556
R9892 VSS.n353 VSS.n351 0.0660556
R9893 VSS.n322 VSS.n307 0.0660556
R9894 VSS.n362 VSS.n361 0.0660556
R9895 VSS.n314 VSS.n312 0.0660556
R9896 VSS.n241 VSS.n240 0.0660556
R9897 VSS.n246 VSS.n245 0.0660556
R9898 VSS.n1172 VSS.n1171 0.0660556
R9899 VSS.n80 VSS.n79 0.0660556
R9900 VSS.n2650 VSS.n2635 0.0660556
R9901 VSS.n2690 VSS.n2689 0.0660556
R9902 VSS.n2681 VSS.n2679 0.0660556
R9903 VSS.n2642 VSS.n2640 0.0660556
R9904 VSS.n85 VSS.n84 0.0660556
R9905 VSS.n2498 VSS.n262 0.0656521
R9906 VSS.n2743 VSS.n2593 0.0656521
R9907 VSS.n2204 VSS.n2203 0.0625
R9908 VSS.n2158 VSS.n2156 0.0625
R9909 VSS.n1349 VSS.n1348 0.0625
R9910 VSS.n1293 VSS.n1291 0.0625
R9911 VSS.n1408 VSS.n1407 0.0625
R9912 VSS.n1202 VSS.n1201 0.0625
R9913 VSS.n2060 VSS.n552 0.0625
R9914 VSS.n545 VSS.n541 0.0608
R9915 VSS.n769 VSS.n767 0.058921
R9916 VSS.n685 VSS.n669 0.0571038
R9917 VSS.n1998 VSS.n1027 0.0548374
R9918 VSS.n767 VSS.n766 0.0547105
R9919 VSS.n920 VSS.n665 0.053063
R9920 VSS.n683 VSS.n666 0.053063
R9921 VSS.n2818 VSS.n30 0.053063
R9922 VSS.n540 VSS.n32 0.053063
R9923 VSS.n2806 VSS.n40 0.053063
R9924 VSS.n2554 VSS.n42 0.053063
R9925 VSS.n764 VSS.n757 0.053063
R9926 VSS.n771 VSS.n765 0.053063
R9927 VSS.n2384 VSS.n421 0.053063
R9928 VSS.n2386 VSS.n419 0.053063
R9929 VSS.n2007 VSS.n581 0.053063
R9930 VSS.n2006 VSS.n582 0.053063
R9931 VSS.n2844 VSS.n14 0.053063
R9932 VSS.n2843 VSS.n16 0.053063
R9933 VSS.n1750 VSS.n1454 0.053063
R9934 VSS.n1765 VSS.n1452 0.053063
R9935 VSS.n1776 VSS.n1445 0.053063
R9936 VSS.n1796 VSS.n1443 0.053063
R9937 VSS.n2390 VSS.n2389 0.0527581
R9938 VSS.n679 VSS.n675 0.0526849
R9939 VSS.n682 VSS.n672 0.0526849
R9940 VSS.n2823 VSS.n2822 0.0526849
R9941 VSS.n29 VSS.n28 0.0526849
R9942 VSS.n2811 VSS.n2810 0.0526849
R9943 VSS.n39 VSS.n38 0.0526849
R9944 VSS.n785 VSS.n784 0.0526849
R9945 VSS.n756 VSS.n755 0.0526849
R9946 VSS.n418 VSS.n417 0.0526849
R9947 VSS.n2392 VSS.n2391 0.0526849
R9948 VSS.n2008 VSS.n578 0.0526849
R9949 VSS.n2003 VSS.n579 0.0526849
R9950 VSS.n1786 VSS.n1783 0.0526849
R9951 VSS.n1789 VSS.n1788 0.0526849
R9952 VSS.n1451 VSS.n1450 0.0526849
R9953 VSS.n1770 VSS.n1769 0.0526849
R9954 VSS.n1442 VSS.n1441 0.0526849
R9955 VSS.n1801 VSS.n1800 0.0526849
R9956 VSS.n2833 VSS.n2832 0.0503305
R9957 VSS.n2562 VSS.n2561 0.049129
R9958 VSS.n2565 VSS.n97 0.0471667
R9959 VSS.n375 VSS.n374 0.0471667
R9960 VSS.n310 VSS.n308 0.0471667
R9961 VSS.n369 VSS.n355 0.0471667
R9962 VSS.n317 VSS.n315 0.0471667
R9963 VSS.n2511 VSS.n2510 0.0471667
R9964 VSS.n2505 VSS.n242 0.0471667
R9965 VSS.n2546 VSS.n2545 0.0471667
R9966 VSS.n2756 VSS.n2755 0.0471667
R9967 VSS.n2638 VSS.n2636 0.0471667
R9968 VSS.n2697 VSS.n2683 0.0471667
R9969 VSS.n2703 VSS.n2702 0.0471667
R9970 VSS.n2645 VSS.n2643 0.0471667
R9971 VSS.n2750 VSS.n81 0.0471667
R9972 VSS.n919 VSS.n918 0.0470126
R9973 VSS.n668 VSS.n667 0.0470126
R9974 VSS.n2817 VSS.n2816 0.0470126
R9975 VSS.n34 VSS.n33 0.0470126
R9976 VSS.n2805 VSS.n2804 0.0470126
R9977 VSS.n44 VSS.n43 0.0470126
R9978 VSS.n773 VSS.n503 0.0470126
R9979 VSS.n772 VSS.n504 0.0470126
R9980 VSS.n2397 VSS.n413 0.0470126
R9981 VSS.n2385 VSS.n414 0.0470126
R9982 VSS.n1021 VSS.n584 0.0470126
R9983 VSS.n1023 VSS.n1022 0.0470126
R9984 VSS.n2836 VSS.n15 0.0470126
R9985 VSS.n2839 VSS.n17 0.0470126
R9986 VSS.n1456 VSS.n1455 0.0470126
R9987 VSS.n1764 VSS.n1763 0.0470126
R9988 VSS.n1447 VSS.n1446 0.0470126
R9989 VSS.n1795 VSS.n1794 0.0470126
R9990 VSS.n2846 VSS.n12 0.0467273
R9991 VSS.n2799 VSS.n2798 0.0455
R9992 VSS.n49 VSS.n48 0.0455
R9993 VSS.n2797 VSS.n46 0.0455
R9994 VSS.n2793 VSS.n53 0.0434545
R9995 VSS.n2792 VSS.n54 0.0434545
R9996 VSS.n2791 VSS.n2790 0.0434545
R9997 VSS.n59 VSS.n51 0.0434545
R9998 VSS.n2499 VSS.n2497 0.0427222
R9999 VSS.n2744 VSS.n2742 0.0427222
R10000 VSS.n2786 VSS.n57 0.0426364
R10001 VSS.n2788 VSS.n2787 0.0426364
R10002 VSS.n2785 VSS.n60 0.0426364
R10003 VSS.n1744 VSS.n1741 0.0425965
R10004 VSS.n1767 VSS.n1766 0.0417185
R10005 VSS.n2533 VSS 0.040834
R10006 VSS.n1916 VSS 0.0402059
R10007 VSS VSS.n2175 0.0401429
R10008 VSS.n2166 VSS 0.0401429
R10009 VSS.n2077 VSS 0.0401429
R10010 VSS VSS.n2079 0.0401429
R10011 VSS.n2122 VSS 0.0401429
R10012 VSS VSS.n2093 0.0401429
R10013 VSS VSS.n516 0.0401429
R10014 VSS VSS.n2196 0.0401429
R10015 VSS.n2187 VSS 0.0401429
R10016 VSS VSS.n2143 0.0401429
R10017 VSS.n2137 VSS 0.0401429
R10018 VSS VSS.n1315 0.0401429
R10019 VSS VSS.n1298 0.0401429
R10020 VSS VSS.n1305 0.0401429
R10021 VSS.n1362 VSS 0.0401429
R10022 VSS.n1343 VSS 0.0401429
R10023 VSS.n1331 VSS 0.0401429
R10024 VSS VSS.n1278 0.0401429
R10025 VSS VSS.n1345 0.0401429
R10026 VSS.n1258 VSS 0.0401429
R10027 VSS.n1245 VSS 0.0401429
R10028 VSS VSS.n1364 0.0401429
R10029 VSS VSS.n1226 0.0401429
R10030 VSS VSS.n1217 0.0401429
R10031 VSS.n1402 VSS 0.0401429
R10032 VSS.n1928 VSS 0.0401429
R10033 VSS.n1417 VSS 0.0401429
R10034 VSS VSS.n1073 0.0401429
R10035 VSS.n1415 VSS 0.0401429
R10036 VSS VSS.n1404 0.0401429
R10037 VSS VSS.n1187 0.0401429
R10038 VSS VSS.n1194 0.0401429
R10039 VSS VSS.n1211 0.0401429
R10040 VSS.n1375 VSS 0.0401429
R10041 VSS.n1313 VSS 0.0401429
R10042 VSS VSS.n513 0.0401429
R10043 VSS.n2073 VSS 0.0401429
R10044 VSS VSS.n525 0.0401429
R10045 VSS.n2173 VSS 0.0401429
R10046 VSS.n2167 VSS 0.0401429
R10047 VSS VSS.n553 0.0401429
R10048 VSS VSS.n555 0.0401429
R10049 VSS.n1873 VSS 0.0401429
R10050 VSS VSS.n1810 0.0401429
R10051 VSS.n1785 VSS.n1784 0.0385455
R10052 VSS.n2473 VSS.n2472 0.0384339
R10053 VSS.n2491 VSS.n2490 0.0384339
R10054 VSS.n289 VSS.n288 0.0384339
R10055 VSS.n346 VSS.n345 0.0384339
R10056 VSS.n2524 VSS.n231 0.0384339
R10057 VSS.n253 VSS.n252 0.0384339
R10058 VSS.n1169 VSS.n1164 0.0384339
R10059 VSS.n2769 VSS.n70 0.0384339
R10060 VSS.n2715 VSS.n2714 0.0384339
R10061 VSS.n2733 VSS.n2732 0.0384339
R10062 VSS.n2674 VSS.n2673 0.0384339
R10063 VSS.n2617 VSS.n2616 0.0384339
R10064 VSS.n2584 VSS.n2583 0.0384339
R10065 VSS.n208 VSS.n207 0.0384339
R10066 VSS.n1026 VSS.n1025 0.0383151
R10067 VSS.n2472 VSS.n2471 0.0376901
R10068 VSS.n2490 VSS.n2489 0.0376901
R10069 VSS.n2484 VSS.n289 0.0376901
R10070 VSS.n2466 VSS.n346 0.0376901
R10071 VSS.n2518 VSS.n231 0.0376901
R10072 VSS.n253 VSS.n249 0.0376901
R10073 VSS.n1170 VSS.n1169 0.0376901
R10074 VSS.n2763 VSS.n70 0.0376901
R10075 VSS.n2714 VSS.n2713 0.0376901
R10076 VSS.n2732 VSS.n2731 0.0376901
R10077 VSS.n2708 VSS.n2674 0.0376901
R10078 VSS.n2726 VSS.n2617 0.0376901
R10079 VSS.n2584 VSS.n88 0.0376901
R10080 VSS.n208 VSS.n101 0.0376901
R10081 VSS.n2794 VSS.n50 0.0369091
R10082 VSS.n2461 VSS.n52 0.0369091
R10083 VSS.n2796 VSS.n2795 0.0369091
R10084 VSS.n2847 VSS.n11 0.0367416
R10085 VSS.n1798 VSS.n1797 0.0366561
R10086 VSS.n2842 VSS.n18 0.0364483
R10087 VSS.n1799 VSS.n1439 0.036396
R10088 VSS.n1787 VSS.n1781 0.0361897
R10089 VSS.n1784 VSS.n11 0.0361376
R10090 VSS.n2820 VSS.n2819 0.0345872
R10091 VSS.n2821 VSS.n26 0.034342
R10092 VSS.n2808 VSS.n2807 0.0339492
R10093 VSS.n2809 VSS.n36 0.0337086
R10094 VSS.n538 VSS.n537 0.0330131
R10095 VSS.n1922 VSS.n1921 0.0329742
R10096 VSS.n8 VSS.n7 0.0327222
R10097 VSS.n1793 VSS.n1444 0.0324942
R10098 VSS.n2841 VSS.n2840 0.0323103
R10099 VSS.n2550 VSS.n222 0.03218
R10100 VSS VSS.n187 0.0310055
R10101 VSS.n681 VSS.n670 0.0307655
R10102 VSS.n2389 VSS.n2387 0.0306935
R10103 VSS.n2815 VSS.n31 0.0306635
R10104 VSS.n2803 VSS.n41 0.0300989
R10105 VSS.n680 VSS.n669 0.0295733
R10106 VSS VSS.n2177 0.0283571
R10107 VSS.n2441 VSS 0.0283571
R10108 VSS.n2083 VSS 0.0283571
R10109 VSS.n2082 VSS 0.0283571
R10110 VSS VSS.n515 0.0283571
R10111 VSS.n2095 VSS 0.0283571
R10112 VSS.n2096 VSS 0.0283571
R10113 VSS.n2198 VSS 0.0283571
R10114 VSS VSS.n2145 0.0283571
R10115 VSS.n2152 VSS 0.0283571
R10116 VSS.n2199 VSS 0.0283571
R10117 VSS VSS.n1317 0.0283571
R10118 VSS VSS.n1323 0.0283571
R10119 VSS.n1322 VSS 0.0283571
R10120 VSS VSS.n1360 0.0283571
R10121 VSS VSS.n1340 0.0283571
R10122 VSS VSS.n1280 0.0283571
R10123 VSS.n1287 VSS 0.0283571
R10124 VSS VSS.n1273 0.0283571
R10125 VSS VSS.n1256 0.0283571
R10126 VSS.n1255 VSS 0.0283571
R10127 VSS VSS.n1244 0.0283571
R10128 VSS.n1229 VSS 0.0283571
R10129 VSS VSS.n1230 0.0283571
R10130 VSS VSS.n1399 0.0283571
R10131 VSS VSS.n1926 0.0283571
R10132 VSS.n1925 VSS 0.0283571
R10133 VSS.n1940 VSS 0.0283571
R10134 VSS.n1941 VSS 0.0283571
R10135 VSS VSS.n1083 0.0283571
R10136 VSS VSS.n1390 0.0283571
R10137 VSS.n1389 VSS 0.0283571
R10138 VSS.n1232 VSS 0.0283571
R10139 VSS VSS.n1213 0.0283571
R10140 VSS VSS.n380 0.0283571
R10141 VSS VSS.n2118 0.0283571
R10142 VSS.n2107 VSS 0.0283571
R10143 VSS.n2106 VSS 0.0283571
R10144 VSS VSS.n387 0.0283571
R10145 VSS.n2442 VSS 0.0283571
R10146 VSS VSS.n2056 0.0283571
R10147 VSS.n2055 VSS 0.0283571
R10148 VSS VSS.n1437 0.0283571
R10149 VSS VSS.n1869 0.0283571
R10150 VSS.n591 VSS.n580 0.0274767
R10151 VSS.n2010 VSS.n2009 0.0272442
R10152 VSS.n125 VSS.n124 0.0271667
R10153 VSS.n2574 VSS 0.02496
R10154 VSS.n121 VSS.n120 0.0249444
R10155 VSS.n2379 VSS.n422 0.0246463
R10156 VSS.n917 VSS.n688 0.0245
R10157 VSS.n781 VSS.n759 0.0243775
R10158 VSS.n1438 VSS.n23 0.0242443
R10159 VSS.n2782 VSS.n2781 0.0241364
R10160 VSS.n2781 VSS.n2780 0.0241364
R10161 VSS.n546 VSS.n537 0.0240602
R10162 VSS.n539 VSS.n538 0.02345
R10163 VSS.n2463 VSS.n2462 0.023
R10164 VSS.n2399 VSS.n2398 0.023
R10165 VSS.n922 VSS.n921 0.0229444
R10166 VSS.n775 VSS.n774 0.0221327
R10167 VSS.n589 VSS.n586 0.0221279
R10168 VSS.n1748 VSS.n1598 0.0220686
R10169 VSS.n783 VSS.n758 0.0213163
R10170 VSS.n2383 VSS.n2382 0.0210793
R10171 VSS.n2013 VSS.n573 0.0209651
R10172 VSS.n1370 VSS.n1236 0.0209124
R10173 VSS VSS.n1102 0.0208571
R10174 VSS.n174 VSS.n110 0.0208571
R10175 VSS.n2447 VSS.n2446 0.0207649
R10176 VSS.n1149 VSS.n1102 0.0197857
R10177 VSS VSS.n110 0.0197857
R10178 VSS.n2382 VSS.n2381 0.018061
R10179 VSS.n678 VSS.n677 0.0173889
R10180 VSS.n1752 VSS.n1751 0.0173627
R10181 VSS.n2798 VSS.n50 0.0172727
R10182 VSS.n2461 VSS.n49 0.0172727
R10183 VSS.n2462 VSS.n2460 0.0172727
R10184 VSS.n2797 VSS.n2796 0.0172727
R10185 VSS.n1812 VSS 0.017201
R10186 VSS.n770 VSS.n769 0.0168158
R10187 VSS.n2001 VSS.n1026 0.0162531
R10188 VSS.n2794 VSS.n2793 0.0160455
R10189 VSS.n2792 VSS.n52 0.0160455
R10190 VSS.n2791 VSS.n55 0.0160455
R10191 VSS.n2795 VSS.n51 0.0160455
R10192 VSS.n788 VSS.n787 0.0158061
R10193 VSS.n2463 VSS.n55 0.0144091
R10194 VSS.n677 VSS.n676 0.0142778
R10195 VSS.n2380 VSS.n2379 0.0142195
R10196 VSS.n2556 VSS.n2555 0.0141364
R10197 VSS.n2498 VSS.n263 0.0138884
R10198 VSS.n2743 VSS.n2594 0.0138884
R10199 VSS.n131 VSS.n130 0.0138333
R10200 VSS.n685 VSS.n670 0.0137168
R10201 VSS.n1778 VSS.n1777 0.013135
R10202 VSS.n1755 VSS.n1754 0.0128529
R10203 VSS.n2827 VSS.n2826 0.0126495
R10204 VSS.n2828 VSS.n2827 0.0126495
R10205 VSS.n2473 VSS.n334 0.0124008
R10206 VSS.n2491 VSS.n277 0.0124008
R10207 VSS.n288 VSS.n286 0.0124008
R10208 VSS.n345 VSS.n343 0.0124008
R10209 VSS.n2525 VSS.n2524 0.0124008
R10210 VSS.n252 VSS.n228 0.0124008
R10211 VSS.n1164 VSS.n1163 0.0124008
R10212 VSS.n2770 VSS.n2769 0.0124008
R10213 VSS.n2715 VSS.n2662 0.0124008
R10214 VSS.n2733 VSS.n2608 0.0124008
R10215 VSS.n2673 VSS.n2671 0.0124008
R10216 VSS.n2616 VSS.n2596 0.0124008
R10217 VSS.n2583 VSS.n2582 0.0124008
R10218 VSS.n207 VSS.n206 0.0124008
R10219 VSS.n1755 VSS.n1457 0.0122647
R10220 VSS.n2399 VSS.n411 0.01175
R10221 VSS.n2212 VSS.n506 0.0115072
R10222 VSS.n928 VSS.n659 0.0113889
R10223 VSS.n2846 VSS.n2845 0.0111364
R10224 VSS.n1753 VSS.n1752 0.0108922
R10225 VSS.n1760 VSS.n1759 0.0108922
R10226 VSS.n331 VSS 0.0105
R10227 VSS.n274 VSS 0.0105
R10228 VSS.n2496 VSS 0.0105
R10229 VSS.n2478 VSS 0.0105
R10230 VSS.n2529 VSS 0.0105
R10231 VSS.n2536 VSS 0.0105
R10232 VSS.n1160 VSS 0.0105
R10233 VSS.n2570 VSS 0.0105
R10234 VSS.n2659 VSS 0.0105
R10235 VSS.n2605 VSS 0.0105
R10236 VSS.n2720 VSS 0.0105
R10237 VSS.n2741 VSS 0.0105
R10238 VSS.n2579 VSS 0.0105
R10239 VSS.n195 VSS 0.0105
R10240 VSS.n2557 VSS.n2556 0.0101503
R10241 VSS.n1778 VSS.n1774 0.00944168
R10242 VSS.n116 VSS.n115 0.00938889
R10243 VSS.n412 VSS.n407 0.0090061
R10244 VSS.n922 VSS.n663 0.00894444
R10245 VSS.n2005 VSS.n1026 0.00826224
R10246 VSS.n758 VSS.n753 0.00784694
R10247 VSS.n1020 VSS.n586 0.00747674
R10248 VSS.n2372 VSS.n2371 0.00681098
R10249 VSS.n2800 VSS.n2799 0.00622727
R10250 VSS.n2801 VSS.n46 0.00622727
R10251 VSS VSS.n2100 0.00606701
R10252 VSS.n1251 VSS 0.00606701
R10253 VSS VSS.n1945 0.00606701
R10254 VSS.n1749 VSS.n1748 0.0059902
R10255 VSS.n2389 VSS.n2388 0.00594885
R10256 VSS.n2010 VSS.n576 0.00584884
R10257 VSS.n591 VSS.n590 0.00584884
R10258 VSS.n57 VSS.n53 0.00540909
R10259 VSS.n2786 VSS.n58 0.00540909
R10260 VSS.n2788 VSS.n54 0.00540909
R10261 VSS.n2790 VSS.n2789 0.00540909
R10262 VSS.n60 VSS.n59 0.00540909
R10263 VSS.n2785 VSS.n2784 0.00540909
R10264 VSS.n1767 VSS.n1448 0.00516523
R10265 VSS VSS.n392 0.00513918
R10266 VSS VSS.n526 0.00513918
R10267 VSS VSS.n385 0.00513918
R10268 VSS.n1369 VSS.n1237 0.00513918
R10269 VSS.n1222 VSS 0.00513918
R10270 VSS.n546 VSS.n545 0.00448601
R10271 VSS.n1768 VSS.n1767 0.00436002
R10272 VSS.n775 VSS.n502 0.00396939
R10273 VSS.n48 VSS.n47 0.00386
R10274 VSS.n1854 VSS 0.00383333
R10275 VSS VSS.n2867 0.00383333
R10276 VSS.n2884 VSS 0.00383333
R10277 VSS VSS.n1118 0.00383333
R10278 VSS.n1135 VSS 0.00383333
R10279 VSS VSS.n1905 0.00383333
R10280 VSS.n135 VSS 0.00383333
R10281 VSS VSS.n159 0.00383333
R10282 VSS VSS.n1985 0.00383333
R10283 VSS.n1962 VSS 0.00383333
R10284 VSS.n1882 VSS 0.00383333
R10285 VSS.n1822 VSS 0.00383333
R10286 VSS.n688 VSS.n664 0.00383333
R10287 VSS.n2787 VSS.n56 0.00345187
R10288 VSS.n2213 VSS.n2212 0.00343706
R10289 VSS.n2112 VSS.n2111 0.00328351
R10290 VSS.n769 VSS.n768 0.00322727
R10291 VSS.n782 VSS.n781 0.00294898
R10292 VSS.n1950 VSS 0.00280769
R10293 VSS VSS.n2162 0.00280769
R10294 VSS.n2190 VSS 0.00280769
R10295 VSS VSS.n2193 0.00280769
R10296 VSS VSS.n508 0.00280769
R10297 VSS VSS.n1297 0.00280769
R10298 VSS.n1334 VSS 0.00280769
R10299 VSS VSS.n1337 0.00280769
R10300 VSS VSS.n1356 0.00280769
R10301 VSS.n1266 VSS 0.00280769
R10302 VSS.n1935 VSS 0.00280769
R10303 VSS VSS.n1074 0.00280769
R10304 VSS VSS.n1396 0.00280769
R10305 VSS.n1382 VSS 0.00280769
R10306 VSS VSS.n1191 0.00280769
R10307 VSS.n1380 VSS 0.00280769
R10308 VSS.n1326 VSS 0.00280769
R10309 VSS.n2130 VSS 0.00280769
R10310 VSS.n2182 VSS 0.00280769
R10311 VSS.n2069 VSS 0.00280769
R10312 VSS VSS.n2071 0.00280769
R10313 VSS.n2050 VSS 0.00280769
R10314 VSS.n1808 VSS 0.00280769
R10315 VSS.n675 VSS.n674 0.00276891
R10316 VSS.n673 VSS.n672 0.00276891
R10317 VSS.n2824 VSS.n2823 0.00276891
R10318 VSS.n28 VSS.n27 0.00276891
R10319 VSS.n2812 VSS.n2811 0.00276891
R10320 VSS.n38 VSS.n37 0.00276891
R10321 VSS.n786 VSS.n785 0.00276891
R10322 VSS.n755 VSS.n754 0.00276891
R10323 VSS.n2370 VSS.n417 0.00276891
R10324 VSS.n2392 VSS.n416 0.00276891
R10325 VSS.n2000 VSS.n578 0.00276891
R10326 VSS.n2003 VSS.n2002 0.00276891
R10327 VSS.n1783 VSS.n1782 0.00276891
R10328 VSS.n1790 VSS.n1789 0.00276891
R10329 VSS.n1742 VSS.n1450 0.00276891
R10330 VSS.n1770 VSS.n1449 0.00276891
R10331 VSS.n1441 VSS.n1440 0.00276891
R10332 VSS.n1802 VSS.n1801 0.00276891
R10333 VSS.n545 VSS.n544 0.00275
R10334 VSS.n763 VSS.n759 0.00254082
R10335 VSS.n2204 VSS 0.0025
R10336 VSS.n2158 VSS 0.0025
R10337 VSS.n1348 VSS 0.0025
R10338 VSS.n1293 VSS 0.0025
R10339 VSS.n1407 VSS 0.0025
R10340 VSS.n1201 VSS 0.0025
R10341 VSS VSS.n2060 0.0025
R10342 VSS.n2847 VSS.n2846 0.00238811
R10343 VSS.n685 VSS.n684 0.00217832
R10344 VSS.n2371 VSS.n422 0.00214634
R10345 VSS.n1803 VSS.n1439 0.00206069
R10346 VSS.n1791 VSS.n1781 0.00205172
R10347 VSS.n918 VSS.n687 0.00201261
R10348 VSS.n686 VSS.n668 0.00201261
R10349 VSS.n2816 VSS.n35 0.00201261
R10350 VSS.n2804 VSS.n45 0.00201261
R10351 VSS.n2215 VSS.n503 0.00201261
R10352 VSS.n2214 VSS.n504 0.00201261
R10353 VSS.n2397 VSS.n2396 0.00201261
R10354 VSS.n2395 VSS.n414 0.00201261
R10355 VSS.n1021 VSS.n585 0.00201261
R10356 VSS.n2839 VSS.n2838 0.00201261
R10357 VSS.n1761 VSS.n1456 0.00201261
R10358 VSS.n1794 VSS.n1780 0.00201261
R10359 VSS.n2825 VSS.n26 0.00197139
R10360 VSS.n2813 VSS.n36 0.00194385
R10361 VSS.n576 VSS.n573 0.00189535
R10362 VSS.n541 VSS.n539 0.00185
R10363 VSS.n676 VSS.n659 0.00183333
R10364 VSS.n1022 VSS.n583 0.00175605
R10365 VSS.n1763 VSS.n1762 0.00175605
R10366 VSS.n2837 VSS.n2836 0.00175604
R10367 VSS.n542 VSS.n34 0.00175602
R10368 VSS.n2552 VSS.n44 0.00175454
R10369 VSS.n1779 VSS.n1447 0.00175286
R10370 VSS.n1785 VSS.n12 0.00172727
R10371 VSS.n787 VSS.n753 0.00172449
R10372 VSS.n1743 VSS.n1598 0.00167647
R10373 VSS.n679 VSS.n665 0.00163445
R10374 VSS.n683 VSS.n682 0.00163445
R10375 VSS.n2822 VSS.n30 0.00163445
R10376 VSS.n540 VSS.n29 0.00163445
R10377 VSS.n2810 VSS.n40 0.00163445
R10378 VSS.n2554 VSS.n39 0.00163445
R10379 VSS.n784 VSS.n757 0.00163445
R10380 VSS.n765 VSS.n756 0.00163445
R10381 VSS.n421 VSS.n418 0.00163445
R10382 VSS.n2391 VSS.n419 0.00163445
R10383 VSS.n2008 VSS.n2007 0.00163445
R10384 VSS.n2006 VSS.n579 0.00163445
R10385 VSS.n1786 VSS.n14 0.00163445
R10386 VSS.n1788 VSS.n16 0.00163445
R10387 VSS.n1750 VSS.n1451 0.00163445
R10388 VSS.n1769 VSS.n1452 0.00163445
R10389 VSS.n1776 VSS.n1442 0.00163445
R10390 VSS.n1800 VSS.n1443 0.00163445
R10391 VSS.n2394 VSS.n388 0.00162735
R10392 VSS VSS.n1849 0.00161111
R10393 VSS VSS.n1846 0.00161111
R10394 VSS.n1860 VSS 0.00161111
R10395 VSS.n1857 VSS 0.00161111
R10396 VSS.n2566 VSS 0.00161111
R10397 VSS.n2856 VSS 0.00161111
R10398 VSS.n2860 VSS 0.00161111
R10399 VSS.n2864 VSS 0.00161111
R10400 VSS.n2876 VSS 0.00161111
R10401 VSS VSS.n2887 0.00161111
R10402 VSS.n2871 VSS 0.00161111
R10403 VSS.n2881 VSS 0.00161111
R10404 VSS.n2891 VSS 0.00161111
R10405 VSS.n2896 VSS 0.00161111
R10406 VSS.n1115 VSS 0.00161111
R10407 VSS.n1127 VSS 0.00161111
R10408 VSS.n1110 VSS 0.00161111
R10409 VSS.n2901 VSS 0.00161111
R10410 VSS VSS.n1138 0.00161111
R10411 VSS.n1122 VSS 0.00161111
R10412 VSS.n1132 VSS 0.00161111
R10413 VSS.n1142 VSS 0.00161111
R10414 VSS.n1153 VSS 0.00161111
R10415 VSS VSS.n1914 0.00161111
R10416 VSS.n1902 VSS 0.00161111
R10417 VSS VSS.n1898 0.00161111
R10418 VSS.n1895 VSS 0.00161111
R10419 VSS.n1908 VSS 0.00161111
R10420 VSS.n373 VSS 0.00161111
R10421 VSS VSS.n321 0.00161111
R10422 VSS.n370 VSS 0.00161111
R10423 VSS VSS.n329 0.00161111
R10424 VSS VSS.n272 0.00161111
R10425 VSS VSS.n2495 0.00161111
R10426 VSS.n318 VSS 0.00161111
R10427 VSS VSS.n2477 0.00161111
R10428 VSS.n2509 VSS 0.00161111
R10429 VSS VSS.n2528 0.00161111
R10430 VSS.n2506 VSS 0.00161111
R10431 VSS.n2540 VSS 0.00161111
R10432 VSS.n2544 VSS 0.00161111
R10433 VSS VSS.n1159 0.00161111
R10434 VSS.n2754 VSS 0.00161111
R10435 VSS.n2773 VSS 0.00161111
R10436 VSS VSS.n2649 0.00161111
R10437 VSS.n2698 VSS 0.00161111
R10438 VSS VSS.n2657 0.00161111
R10439 VSS VSS.n2603 0.00161111
R10440 VSS.n2701 VSS 0.00161111
R10441 VSS VSS.n2719 0.00161111
R10442 VSS.n2646 VSS 0.00161111
R10443 VSS.n2737 VSS 0.00161111
R10444 VSS.n2751 VSS 0.00161111
R10445 VSS.n172 VSS 0.00161111
R10446 VSS VSS.n129 0.00161111
R10447 VSS.n126 VSS 0.00161111
R10448 VSS VSS.n138 0.00161111
R10449 VSS.n144 VSS 0.00161111
R10450 VSS.n156 VSS 0.00161111
R10451 VSS VSS.n152 0.00161111
R10452 VSS.n149 VSS 0.00161111
R10453 VSS.n182 VSS 0.00161111
R10454 VSS.n178 VSS 0.00161111
R10455 VSS VSS.n2577 0.00161111
R10456 VSS.n203 VSS 0.00161111
R10457 VSS.n1033 VSS 0.00161111
R10458 VSS.n1982 VSS 0.00161111
R10459 VSS VSS.n1978 0.00161111
R10460 VSS.n1975 VSS 0.00161111
R10461 VSS.n1987 VSS 0.00161111
R10462 VSS.n1991 VSS 0.00161111
R10463 VSS VSS.n1965 0.00161111
R10464 VSS.n1971 VSS 0.00161111
R10465 VSS.n1959 VSS 0.00161111
R10466 VSS.n1956 VSS 0.00161111
R10467 VSS VSS.n1885 0.00161111
R10468 VSS.n1891 VSS 0.00161111
R10469 VSS.n1879 VSS 0.00161111
R10470 VSS.n1876 VSS 0.00161111
R10471 VSS.n1838 VSS 0.00161111
R10472 VSS VSS.n1824 0.00161111
R10473 VSS VSS.n1842 0.00161111
R10474 VSS.n1834 VSS 0.00161111
R10475 VSS.n1830 VSS 0.00161111
R10476 VSS.n916 VSS.n915 0.00161111
R10477 VSS.n2398 VSS.n412 0.00159756
R10478 VSS.n2213 VSS.n505 0.00154895
R10479 VSS.n1793 VSS.n1792 0.00154046
R10480 VSS.n2840 VSS.n2835 0.00153448
R10481 VSS.n2831 VSS 0.00151695
R10482 VSS.n2815 VSS.n2814 0.00148093
R10483 VSS.n2803 VSS.n2802 0.00146257
R10484 VSS.n1020 VSS.n1019 0.00143023
R10485 VSS.n917 VSS.n916 0.00138889
R10486 VSS.n2558 VSS.n2557 0.00133916
R10487 VSS.n2005 VSS.n2004 0.00133916
R10488 VSS.n2381 VSS.n2380 0.00132317
R10489 VSS.n2216 VSS.n502 0.00131633
R10490 VSS.n1760 VSS.n1457 0.00128431
R10491 VSS.n1799 VSS.n1798 0.00128035
R10492 VSS.n1771 VSS.n1448 0.00127754
R10493 VSS.n1774 VSS.n1773 0.00127754
R10494 VSS.n1787 VSS.n18 0.00127586
R10495 VSS.n1178 VSS 0.0012438
R10496 VSS.n1180 VSS 0.0012438
R10497 VSS VSS.n2569 0.0012438
R10498 VSS.n189 VSS 0.0012438
R10499 VSS.n1995 VSS 0.0012438
R10500 VSS.n2821 VSS.n2820 0.0012357
R10501 VSS.n2809 VSS.n2808 0.00122193
R10502 VSS.n678 VSS.n663 0.00116667
R10503 VSS.n783 VSS.n782 0.00111224
R10504 VSS.n1751 VSS.n1749 0.00108824
R10505 VSS.n2394 VSS.n2393 0.00106367
R10506 VSS.n2009 VSS.n577 0.000965116
R10507 VSS.n544 VSS.n543 0.00095
R10508 VSS.n684 VSS.n671 0.00091958
R10509 VSS.n671 VSS.n536 0.00091958
R10510 VSS.n768 VSS.n505 0.00091958
R10511 VSS.n2559 VSS.n2558 0.00091958
R10512 VSS.n2555 VSS.n2553 0.00091958
R10513 VSS.n2845 VSS.n13 0.000909091
R10514 VSS.n1773 VSS.n1772 0.000888769
R10515 VSS.n1777 VSS.n1775 0.000888769
R10516 VSS.n920 VSS.n919 0.000878151
R10517 VSS.n667 VSS.n666 0.000878151
R10518 VSS.n2818 VSS.n2817 0.000878151
R10519 VSS.n33 VSS.n32 0.000878151
R10520 VSS.n2806 VSS.n2805 0.000878151
R10521 VSS.n43 VSS.n42 0.000878151
R10522 VSS.n773 VSS.n764 0.000878151
R10523 VSS.n772 VSS.n771 0.000878151
R10524 VSS.n2384 VSS.n413 0.000878151
R10525 VSS.n2386 VSS.n2385 0.000878151
R10526 VSS.n584 VSS.n581 0.000878151
R10527 VSS.n1023 VSS.n582 0.000878151
R10528 VSS.n1025 VSS.n1024 0.000878151
R10529 VSS.n2844 VSS.n15 0.000878151
R10530 VSS.n2843 VSS.n17 0.000878151
R10531 VSS.n1455 VSS.n1454 0.000878151
R10532 VSS.n1765 VSS.n1764 0.000878151
R10533 VSS.n1766 VSS.n1453 0.000878151
R10534 VSS.n1446 VSS.n1445 0.000878151
R10535 VSS.n1796 VSS.n1795 0.000878151
R10536 VSS.n2388 VSS.n415 0.000875783
R10537 VSS.n2393 VSS.n415 0.000875783
R10538 VSS.n2383 VSS.n411 0.00077439
R10539 VSS.n1797 VSS.n1444 0.000760116
R10540 VSS.n2842 VSS.n2841 0.000758621
R10541 VSS.n2819 VSS.n31 0.000745232
R10542 VSS.n2807 VSS.n41 0.000740642
R10543 VSS.n580 VSS.n577 0.000732558
R10544 VSS.n590 VSS.n589 0.000732558
R10545 VSS.n921 VSS.n664 0.000722222
R10546 VSS.n774 VSS.n763 0.000704082
R10547 VSS.n1744 VSS.n1743 0.000696078
R10548 VSS.n1754 VSS.n1753 0.000696078
R10549 7b_counter_0.MDFF_6.QB.n3 7b_counter_0.MDFF_6.QB.t6 53.2954
R10550 7b_counter_0.MDFF_6.QB.n1 7b_counter_0.MDFF_6.QB.t3 38.8649
R10551 7b_counter_0.MDFF_6.QB.n0 7b_counter_0.MDFF_6.QB.t5 28.8568
R10552 7b_counter_0.MDFF_6.tspc2_magic_0.QB 7b_counter_0.MDFF_6.QB.n4 23.3781
R10553 7b_counter_0.MDFF_6.tspc2_magic_0.QB 7b_counter_0.MDFF_6.mux_magic_0.IN1 19.3581
R10554 7b_counter_0.MDFF_6.QB.n4 7b_counter_0.MDFF_6.QB.t2 17.1425
R10555 7b_counter_0.MDFF_6.QB.t3 7b_counter_0.MDFF_6.QB.n0 17.0773
R10556 7b_counter_0.MDFF_6.QB.n4 7b_counter_0.MDFF_6.QB.t8 14.405
R10557 7b_counter_0.MDFF_6.QB.n0 7b_counter_0.MDFF_6.QB.t7 11.6023
R10558 7b_counter_0.MDFF_6.mux_magic_0.IN1 7b_counter_0.MDFF_6.QB.n1 9.42108
R10559 7b_counter_0.MDFF_6.QB.n3 7b_counter_0.MDFF_6.QB.n2 8.51584
R10560 7b_counter_0.MDFF_6.QB.n1 7b_counter_0.MDFF_6.QB.t4 7.3005
R10561 7b_counter_0.MDFF_6.QB.t8 7b_counter_0.MDFF_6.QB.n3 7.3005
R10562 7b_counter_0.MDFF_6.QB.n2 7b_counter_0.MDFF_6.QB.t1 3.62007
R10563 7b_counter_0.MDFF_6.QB.n2 7b_counter_0.MDFF_6.QB.t0 3.15478
R10564 Q3.t16 Q3.t30 47.8944
R10565 Q3.t5 Q3.t21 47.8944
R10566 Q3.t15 Q3.t27 47.5387
R10567 Q3.t31 Q3.t19 47.5387
R10568 Q3.n19 Q3.n18 43.2428
R10569 Q3.n4 Q3.t8 38.8649
R10570 Q3.n13 Q3.t13 38.7949
R10571 Q3.n12 Q3.t7 38.7949
R10572 Q3.n8 Q3.t29 38.7949
R10573 Q3.n7 Q3.t25 38.7949
R10574 Q3.t3 Q3.t18 31.5469
R10575 Q3.t26 Q3.t6 31.5469
R10576 Q3.t14 Q3.t26 31.5469
R10577 Q3.n13 Q3.n12 31.4949
R10578 Q3.n8 Q3.n7 31.4949
R10579 Q3.n3 Q3.t22 28.8568
R10580 Q3.t18 Q3.t24 28.8094
R10581 Q3.t6 Q3.t12 26.9844
R10582 Q3.n20 Q3.n19 24.9435
R10583 Q3.n14 Q3.t4 17.9416
R10584 Q3.n9 Q3.t23 17.9416
R10585 Q3 Q3.n0 17.8451
R10586 Q3.t8 Q3.n3 17.0773
R10587 Q3.n0 Q3.t14 16.4255
R10588 Q3.n15 Q3.t15 15.7085
R10589 Q3.n6 Q3.t31 15.7085
R10590 Q3.n0 Q3.t3 15.1219
R10591 Q3.n15 Q3.t17 13.4273
R10592 Q3.n6 Q3.t9 13.4273
R10593 Q3.n19 Q3.n5 12.0001
R10594 Q3.n14 Q3.t16 11.957
R10595 Q3.n9 Q3.t5 11.957
R10596 Q3.n3 Q3.t28 11.6023
R10597 Q3.n11 Q3.n10 10.1437
R10598 Q3 Q3.n14 9.94647
R10599 Q3 Q3.n9 9.94647
R10600 Q3 Q3.n4 9.27587
R10601 Q3.n16 Q3.n11 9.00165
R10602 Q3.n18 Q3.n17 9.00165
R10603 Q3 Q3.n15 8.08021
R10604 Q3 Q3.n6 8.08021
R10605 Q3.n4 Q3.t10 7.3005
R10606 Q3.n12 Q3.t20 7.3005
R10607 Q3.t4 Q3.n13 7.3005
R10608 Q3.n7 Q3.t11 7.3005
R10609 Q3.t23 Q3.n8 7.3005
R10610 Q3.n1 Q3.t2 5.47387
R10611 Q3.n2 Q3.t0 4.65398
R10612 Q3.n1 Q3.t1 4.2255
R10613 Q3.n10 Q3 2.64076
R10614 Q3.n16 Q3 2.37798
R10615 Q3.n10 Q3 0.477999
R10616 Q3.n17 Q3 0.473682
R10617 Q3.n2 Q3.n1 0.427022
R10618 Q3 Q3.n2 0.257096
R10619 Q3.n17 Q3.n16 0.229175
R10620 Q3.n18 Q3.n11 0.2075
R10621 Q3 Q3.n21 0.184413
R10622 Q3.n20 Q3 0.0260556
R10623 Q3.n21 Q3 0.0238333
R10624 Q3.n5 Q3 0.0130316
R10625 Q3.n5 Q3 0.00733544
R10626 Q3.n21 Q3.n20 0.00383333
R10627 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t7 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t18 47.8944
R10628 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t23 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t8 47.8944
R10629 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n1 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t17 38.7949
R10630 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n2 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t14 38.7949
R10631 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t16 38.7949
R10632 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n5 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t10 38.7949
R10633 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n2 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n1 31.4949
R10634 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n5 31.4949
R10635 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t9 31.3561
R10636 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t15 31.3559
R10637 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n0 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t19 26.9781
R10638 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n0 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t20 26.9781
R10639 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n4 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t21 26.9781
R10640 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n4 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t6 26.9781
R10641 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t22 17.9416
R10642 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n7 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t11 17.9416
R10643 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t7 11.957
R10644 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n7 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t23 11.957
R10645 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 10.0107
R10646 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n3 10.0013
R10647 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n7 9.77618
R10648 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 8.14207
R10649 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n1 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t12 7.3005
R10650 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t22 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n2 7.3005
R10651 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n0 7.3005
R10652 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n5 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t13 7.3005
R10653 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t11 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n6 7.3005
R10654 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n4 7.3005
R10655 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n8 4.9131
R10656 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n9 3.6455
R10657 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n11 3.4888
R10658 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n10 3.31072
R10659 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n10 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t2 1.6255
R10660 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n10 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t1 1.6255
R10661 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n11 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t0 1.6255
R10662 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n11 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t3 1.6255
R10663 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t5 1.463
R10664 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t4 1.463
R10665 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t15 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t14 47.8944
R10666 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n0 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t16 38.7949
R10667 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n1 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t17 38.7949
R10668 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n1 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n0 31.4949
R10669 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n2 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t13 17.9416
R10670 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n2 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t15 11.957
R10671 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n7 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 10.4306
R10672 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n2 9.96162
R10673 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n0 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t12 7.3005
R10674 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t13 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n1 7.3005
R10675 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n4 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t1 5.68115
R10676 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t9 4.92604
R10677 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n8 3.6455
R10678 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n9 3.31072
R10679 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n5 3.1505
R10680 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n10 2.90572
R10681 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n4 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n3 2.6005
R10682 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n7 1.91911
R10683 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n7 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 1.88467
R10684 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t0 1.6255
R10685 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t2 1.6255
R10686 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t5 1.6255
R10687 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n9 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t3 1.6255
R10688 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n10 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t4 1.6255
R10689 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n10 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t6 1.6255
R10690 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n5 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t11 1.463
R10691 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n5 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t10 1.463
R10692 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t7 1.463
R10693 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n8 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t8 1.463
R10694 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n6 1.34968
R10695 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n6 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n4 0.898543
R10696 D2_4.t13 D2_4.t2 47.8944
R10697 D2_4.t4 D2_4.t21 47.8944
R10698 D2_4.t14 D2_4.t0 47.5387
R10699 D2_4.t5 D2_4.t18 47.5387
R10700 D2_4.n14 D2_4.n11 43.5378
R10701 D2_4.n17 D2_4.t22 38.8649
R10702 D2_4.n13 D2_4.t24 38.8649
R10703 D2_4.n7 D2_4.t15 38.7949
R10704 D2_4.n6 D2_4.t16 38.7949
R10705 D2_4.n2 D2_4.t7 38.7949
R10706 D2_4.n1 D2_4.t9 38.7949
R10707 D2_4.n7 D2_4.n6 31.4949
R10708 D2_4.n2 D2_4.n1 31.4949
R10709 D2_4.n16 D2_4.t6 28.8568
R10710 D2_4.n12 D2_4.t25 28.8568
R10711 D2_4.n11 D2_4.n5 20.6621
R10712 D2_4.n8 D2_4.t1 17.9416
R10713 D2_4.n3 D2_4.t19 17.9416
R10714 D2_4.t22 D2_4.n16 17.0773
R10715 D2_4.t24 D2_4.n12 17.0773
R10716 D2_4.n9 D2_4.t14 16.621
R10717 D2_4.n4 D2_4.t5 16.621
R10718 D2_4.n9 D2_4.t17 12.5148
R10719 D2_4.n4 D2_4.t10 12.5148
R10720 D2_4.n8 D2_4.t13 11.957
R10721 D2_4.n3 D2_4.t4 11.957
R10722 D2_4.n16 D2_4.t3 11.6023
R10723 D2_4.n12 D2_4.t11 11.6023
R10724 D2_4.n15 D2_4.n14 10.5535
R10725 D2_4 D2_4.n8 9.95286
R10726 D2_4 D2_4.n3 9.95286
R10727 D2_4 D2_4.n17 9.27587
R10728 D2_4 D2_4.n13 9.27587
R10729 D2_4 D2_4.n9 8.59246
R10730 D2_4 D2_4.n4 8.59246
R10731 D2_4.n17 D2_4.t23 7.3005
R10732 D2_4.n13 D2_4.t8 7.3005
R10733 D2_4.n6 D2_4.t20 7.3005
R10734 D2_4.t1 D2_4.n7 7.3005
R10735 D2_4.n1 D2_4.t12 7.3005
R10736 D2_4.t19 D2_4.n2 7.3005
R10737 D2_4.n14 D2_4 5.5699
R10738 D2_4.n11 D2_4.n10 4.86714
R10739 D2_4.n5 D2_4 1.37202
R10740 D2_4.n10 D2_4 1.30354
R10741 D2_4.n10 D2_4 0.24123
R10742 D2_4.n5 D2_4 0.172752
R10743 D2_4.n15 D2_4.n0 0.0468264
R10744 D2_4 D2_4.n15 0.0339615
R10745 D2_4.n0 D2_4 0.0108108
R10746 D2_4.n0 D2_4 0.00311992
R10747 p2_gen_magic_0.xnor_magic_3.OUT.n0 p2_gen_magic_0.xnor_magic_3.OUT.t3 39.1562
R10748 p2_gen_magic_0.xnor_magic_3.OUT.t5 p2_gen_magic_0.xnor_magic_3.OUT.t4 28.8746
R10749 p2_gen_magic_0.xnor_magic_3.OUT.t3 p2_gen_magic_0.xnor_magic_3.OUT.t2 23.4648
R10750 p2_gen_magic_0.xnor_magic_3.OUT.n2 p2_gen_magic_0.xnor_magic_3.OUT.n0 17.1813
R10751 p2_gen_magic_0.xnor_magic_3.OUT.n1 p2_gen_magic_0.xnor_magic_3.OUT.t6 14.1443
R10752 p2_gen_magic_0.xnor_magic_3.OUT.n1 p2_gen_magic_0.xnor_magic_3.OUT.t5 13.8835
R10753 p2_gen_magic_0.xnor_magic_3.OUT.n0 p2_gen_magic_0.xnor_magic_3.OUT.n1 12.5017
R10754 p2_gen_magic_0.xnor_magic_3.OUT.n2 p2_gen_magic_0.xnor_magic_3.OUT.t1 9.23184
R10755 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_3.OUT.n2 5.86488
R10756 p2_gen_magic_0.xnor_magic_3.OUT.n0 p2_gen_magic_0.xnor_magic_3.OUT 5.43085
R10757 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_3.OUT.t0 3.11311
R10758 P2.t13 P2.t8 47.8944
R10759 P2.t11 P2.t12 44.6331
R10760 P2.t6 P2.t11 43.4094
R10761 P2.n0 P2.t7 38.7949
R10762 P2.n1 P2.t14 38.7949
R10763 P2.t10 P2.t6 31.5469
R10764 P2.n1 P2.n0 31.4949
R10765 P2.n4 P2 27.0879
R10766 P2.n2 P2.t9 17.9416
R10767 P2.n3 P2.t10 15.0567
R10768 P2.n3 P2.t16 13.6228
R10769 P2.n2 P2.t13 11.957
R10770 P2 P2.n2 9.95929
R10771 P2 P2.n3 8.2675
R10772 P2.n0 P2.t15 7.3005
R10773 P2.t9 P2.n1 7.3005
R10774 P2.n8 P2.n6 3.6455
R10775 P2.n8 P2.n7 3.31072
R10776 P2.n9 P2.n5 2.90572
R10777 P2.n5 P2.t2 1.6255
R10778 P2.n5 P2.t0 1.6255
R10779 P2.n7 P2.t1 1.6255
R10780 P2.n7 P2.t3 1.6255
R10781 P2.n6 P2.t5 1.463
R10782 P2.n6 P2.t4 1.463
R10783 P2.n10 P2 0.642239
R10784 P2.n4 P2 0.629125
R10785 P2.n9 P2.n8 0.4055
R10786 P2 P2.n4 0.383157
R10787 P2 P2.n9 0.178625
R10788 P2.n10 P2 0.12963
R10789 P2 P2.n10 0.112022
R10790 p3_gen_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VIN 53.9092
R10791 p3_gen_magic_0.xnor_magic_1.B.t3 p3_gen_magic_0.xnor_magic_1.B.t1 47.8944
R10792 p3_gen_magic_0.xnor_magic_1.B.t8 p3_gen_magic_0.xnor_magic_1.B.t6 47.5387
R10793 p3_gen_magic_0.xnor_magic_1.B.n1 p3_gen_magic_0.xnor_magic_1.B.t2 38.7949
R10794 p3_gen_magic_0.xnor_magic_1.B.n0 p3_gen_magic_0.xnor_magic_1.B.t0 38.7949
R10795 p3_gen_magic_0.xnor_magic_1.B.n1 p3_gen_magic_0.xnor_magic_1.B.n0 31.4949
R10796 p3_gen_magic_0.xnor_magic_1.B.n2 p3_gen_magic_0.xnor_magic_1.B.t7 17.9416
R10797 p3_gen_magic_0.xnor_magic_1.B.n3 p3_gen_magic_0.xnor_magic_1.B.t8 16.621
R10798 p3_gen_magic_0.xnor_magic_1.B.n3 p3_gen_magic_0.xnor_magic_1.B.t5 12.5148
R10799 p3_gen_magic_0.xnor_magic_1.B.n2 p3_gen_magic_0.xnor_magic_1.B.t3 11.957
R10800 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VIN p3_gen_magic_0.xnor_magic_1.B.n3 10.0765
R10801 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VIN p3_gen_magic_0.xnor_magic_1.B.n2 9.95286
R10802 p3_gen_magic_0.xnor_magic_1.B.n0 p3_gen_magic_0.xnor_magic_1.B.t4 7.3005
R10803 p3_gen_magic_0.xnor_magic_1.B.t7 p3_gen_magic_0.xnor_magic_1.B.n1 7.3005
R10804 D2_3.t6 D2_3.t21 47.8944
R10805 D2_3.t15 D2_3.t2 47.8944
R10806 D2_3.t4 D2_3.t18 47.5387
R10807 D2_3.t11 D2_3.t25 47.5387
R10808 D2_3.n4 D2_3.t13 38.8649
R10809 D2_3.n1 D2_3.t0 38.8649
R10810 D2_3.n11 D2_3.t7 38.7949
R10811 D2_3.n10 D2_3.t12 38.7949
R10812 D2_3.n7 D2_3.t19 38.7949
R10813 D2_3.n6 D2_3.t24 38.7949
R10814 D2_3.n15 D2_3.n14 35.6362
R10815 D2_3.n11 D2_3.n10 31.4949
R10816 D2_3.n7 D2_3.n6 31.4949
R10817 D2_3.n3 D2_3.t14 28.8568
R10818 D2_3.n0 D2_3.t3 28.8568
R10819 D2_3.n15 D2_3.n9 22.1721
R10820 D2_3.n12 D2_3.t23 17.9416
R10821 D2_3.n8 D2_3.t5 17.9416
R10822 D2_3.t13 D2_3.n3 17.0773
R10823 D2_3.t0 D2_3.n0 17.0773
R10824 D2_3.n13 D2_3.t4 16.621
R10825 D2_3.n5 D2_3.t11 16.621
R10826 D2_3.n13 D2_3.t8 12.5148
R10827 D2_3.n5 D2_3.t17 12.5148
R10828 D2_3.n12 D2_3.t6 11.957
R10829 D2_3.n8 D2_3.t15 11.957
R10830 D2_3.n16 D2_3 11.8418
R10831 D2_3.n3 D2_3.t22 11.6023
R10832 D2_3.n0 D2_3.t10 11.6023
R10833 D2_3 D2_3.n12 9.95286
R10834 D2_3 D2_3.n8 9.95286
R10835 D2_3 D2_3.n4 9.27587
R10836 D2_3 D2_3.n1 9.27587
R10837 D2_3 D2_3.n13 8.59246
R10838 D2_3 D2_3.n5 8.59246
R10839 D2_3.n10 D2_3.t9 7.3005
R10840 D2_3.t23 D2_3.n11 7.3005
R10841 D2_3.n6 D2_3.t20 7.3005
R10842 D2_3.t5 D2_3.n7 7.3005
R10843 D2_3.n4 D2_3.t16 7.3005
R10844 D2_3.n1 D2_3.t1 7.3005
R10845 D2_3.n16 D2_3.n15 5.5297
R10846 D2_3.n17 D2_3.n16 4.5005
R10847 D2_3.n14 D2_3 1.4092
R10848 D2_3.n9 D2_3 1.25659
R10849 D2_3.n14 D2_3 0.135578
R10850 D2_3.n9 D2_3 0.133622
R10851 D2_3.n17 D2_3.n2 0.0468409
R10852 D2_3 D2_3.n17 0.0339615
R10853 D2_3.n2 D2_3 0.0108063
R10854 D2_3.n2 D2_3 0.00911964
R10855 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t10 130.41
R10856 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n5 36.752
R10857 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t7 35.3186
R10858 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t8 33.5023
R10859 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t4 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n0 33.5023
R10860 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t11 32.2349
R10861 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n2 27.7405
R10862 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t6 26.3857
R10863 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t4 16.3786
R10864 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t6 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n3 13.2317
R10865 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n1 12.5032
R10866 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t5 11.3259
R10867 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t3 11.146
R10868 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t12 7.3005
R10869 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t9 7.3005
R10870 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n4 5.87653
R10871 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t2 5.47387
R10872 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t1 5.28011
R10873 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t0 4.65398
R10874 7b_counter_0.MDFF_0.QB.n3 7b_counter_0.MDFF_0.QB.t8 53.0716
R10875 7b_counter_0.MDFF_0.QB.n1 7b_counter_0.MDFF_0.QB.t7 38.8649
R10876 7b_counter_0.MDFF_0.QB.n0 7b_counter_0.MDFF_0.QB.t4 28.8568
R10877 7b_counter_0.MDFF_0.tspc2_magic_0.QB 7b_counter_0.MDFF_0.QB.n4 23.3781
R10878 7b_counter_0.MDFF_0.tspc2_magic_0.QB 7b_counter_0.MDFF_0.mux_magic_0.IN1 17.999
R10879 7b_counter_0.MDFF_0.QB.n4 7b_counter_0.MDFF_0.QB.t6 17.2076
R10880 7b_counter_0.MDFF_0.QB.t7 7b_counter_0.MDFF_0.QB.n0 17.0773
R10881 7b_counter_0.MDFF_0.QB.n4 7b_counter_0.MDFF_0.QB.t3 14.3398
R10882 7b_counter_0.MDFF_0.QB.n0 7b_counter_0.MDFF_0.QB.t5 11.6023
R10883 7b_counter_0.MDFF_0.mux_magic_0.IN1 7b_counter_0.MDFF_0.QB.n1 9.42008
R10884 7b_counter_0.MDFF_0.QB.n3 7b_counter_0.MDFF_0.QB.n2 8.51584
R10885 7b_counter_0.MDFF_0.QB.n1 7b_counter_0.MDFF_0.QB.t2 7.3005
R10886 7b_counter_0.MDFF_0.QB.t3 7b_counter_0.MDFF_0.QB.n3 7.3005
R10887 7b_counter_0.MDFF_0.QB.n2 7b_counter_0.MDFF_0.QB.t1 3.62007
R10888 7b_counter_0.MDFF_0.QB.n2 7b_counter_0.MDFF_0.QB.t0 3.15478
R10889 p2_gen_magic_0.xnor_magic_1.OUT.n2 p2_gen_magic_0.xnor_magic_1.OUT 49.7902
R10890 p2_gen_magic_0.xnor_magic_1.OUT.n1 p2_gen_magic_0.xnor_magic_1.OUT.t4 38.8649
R10891 p2_gen_magic_0.xnor_magic_1.OUT.n0 p2_gen_magic_0.xnor_magic_1.OUT.t5 28.8568
R10892 p2_gen_magic_0.xnor_magic_1.OUT.t4 p2_gen_magic_0.xnor_magic_1.OUT.n0 17.0773
R10893 p2_gen_magic_0.xnor_magic_1.OUT.n0 p2_gen_magic_0.xnor_magic_1.OUT.t2 11.6023
R10894 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_1.OUT.n1 9.27587
R10895 p2_gen_magic_0.xnor_magic_1.OUT.n2 p2_gen_magic_0.xnor_magic_1.OUT.t1 9.23184
R10896 p2_gen_magic_0.xnor_magic_1.OUT.n1 p2_gen_magic_0.xnor_magic_1.OUT.t3 7.3005
R10897 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_1.OUT.n2 5.86488
R10898 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_1.OUT.t0 3.11311
R10899 Q2.t26 Q2.t19 47.8944
R10900 Q2.t7 Q2.t28 47.8944
R10901 Q2.t27 Q2.t20 47.5387
R10902 Q2.t8 Q2.t29 47.5387
R10903 Q2 Q2.n18 39.7641
R10904 Q2.n17 Q2.t12 38.8649
R10905 Q2.n10 Q2.t22 38.7949
R10906 Q2.n9 Q2.t23 38.7949
R10907 Q2.n5 Q2.t4 38.7949
R10908 Q2.n4 Q2.t5 38.7949
R10909 Q2.n15 Q2.n3 37.8543
R10910 Q2.t6 Q2.t13 31.5469
R10911 Q2.t18 Q2.t6 31.5469
R10912 Q2.t10 Q2.t18 31.5469
R10913 Q2.n10 Q2.n9 31.4949
R10914 Q2.n5 Q2.n4 31.4949
R10915 Q2.n15 Q2.n14 29.8511
R10916 Q2.n16 Q2.t21 28.8568
R10917 Q2.t25 Q2.t31 28.8094
R10918 Q2.n14 Q2.n13 27.0771
R10919 Q2.t13 Q2.t16 26.9844
R10920 Q2.n11 Q2.t14 17.9416
R10921 Q2.n6 Q2.t24 17.9416
R10922 Q2.t12 Q2.n16 17.0773
R10923 Q2.n2 Q2.t10 15.9693
R10924 Q2.n12 Q2.t27 15.7085
R10925 Q2.n7 Q2.t8 15.7085
R10926 Q2.n2 Q2.t25 15.5782
R10927 Q2.n12 Q2.t3 13.4273
R10928 Q2.n7 Q2.t11 13.4273
R10929 Q2.n3 Q2.n2 13.012
R10930 Q2.n14 Q2.n8 12.8746
R10931 Q2.n11 Q2.t26 11.957
R10932 Q2.n6 Q2.t7 11.957
R10933 Q2.n16 Q2.t30 11.6023
R10934 Q2 Q2.n11 9.94647
R10935 Q2 Q2.n6 9.94647
R10936 Q2 Q2.n17 9.27587
R10937 Q2 Q2.n12 8.08021
R10938 Q2 Q2.n7 8.08021
R10939 Q2.n9 Q2.t9 7.3005
R10940 Q2.t14 Q2.n10 7.3005
R10941 Q2.n4 Q2.t17 7.3005
R10942 Q2.t24 Q2.n5 7.3005
R10943 Q2.n17 Q2.t15 7.3005
R10944 Q2.n0 Q2.t2 5.47387
R10945 Q2.n1 Q2.t0 4.65398
R10946 Q2.n3 Q2 4.57782
R10947 Q2.n0 Q2.t1 4.2255
R10948 Q2.n8 Q2 2.60172
R10949 Q2.n13 Q2 2.48458
R10950 Q2 Q2.n15 1.96301
R10951 Q2.n13 Q2 0.550045
R10952 Q2.n8 Q2 0.469045
R10953 Q2.n1 Q2.n0 0.427022
R10954 Q2 Q2.n1 0.257096
R10955 Q2.n18 Q2 0.18746
R10956 Q2.n18 Q2 0.00286842
R10957 D2_6.t11 D2_6.t1 47.8944
R10958 D2_6.t4 D2_6.t20 47.8944
R10959 D2_6.t25 D2_6.t19 47.5387
R10960 D2_6.t15 D2_6.t9 47.5387
R10961 D2_6.n13 D2_6.n4 40.7121
R10962 D2_6.n16 D2_6.t12 38.8649
R10963 D2_6.n11 D2_6.t21 38.8649
R10964 D2_6.n6 D2_6.t8 38.7949
R10965 D2_6.n5 D2_6.t6 38.7949
R10966 D2_6.n1 D2_6.t0 38.7949
R10967 D2_6.n0 D2_6.t23 38.7949
R10968 D2_6.n6 D2_6.n5 31.4949
R10969 D2_6.n1 D2_6.n0 31.4949
R10970 D2_6.n15 D2_6.t16 28.8568
R10971 D2_6.n10 D2_6.t2 28.8568
R10972 D2_6.n7 D2_6.t22 17.9416
R10973 D2_6.n2 D2_6.t14 17.9416
R10974 D2_6.t12 D2_6.n15 17.0773
R10975 D2_6.t21 D2_6.n10 17.0773
R10976 D2_6.n12 D2_6.n9 16.749
R10977 D2_6.n8 D2_6.t25 16.621
R10978 D2_6.n3 D2_6.t15 16.621
R10979 D2_6.n8 D2_6.t17 12.5148
R10980 D2_6.n3 D2_6.t7 12.5148
R10981 D2_6.n7 D2_6.t11 11.957
R10982 D2_6.n2 D2_6.t4 11.957
R10983 D2_6.n15 D2_6.t24 11.6023
R10984 D2_6.n10 D2_6.t3 11.6023
R10985 D2_6 D2_6.n7 9.95286
R10986 D2_6 D2_6.n2 9.95286
R10987 D2_6 D2_6.n16 9.27587
R10988 D2_6 D2_6.n11 9.27587
R10989 D2_6 D2_6.n8 8.59246
R10990 D2_6 D2_6.n3 8.59246
R10991 D2_6.n16 D2_6.t10 7.3005
R10992 D2_6.n5 D2_6.t13 7.3005
R10993 D2_6.t22 D2_6.n6 7.3005
R10994 D2_6.n11 D2_6.t18 7.3005
R10995 D2_6.n0 D2_6.t5 7.3005
R10996 D2_6.t14 D2_6.n1 7.3005
R10997 D2_6.n13 D2_6.n12 5.61914
R10998 D2_6.n14 D2_6.n13 4.95532
R10999 D2_6.n12 D2_6 3.5062
R11000 D2_6.n9 D2_6 1.36028
R11001 D2_6.n4 D2_6 1.34267
R11002 D2_6.n4 D2_6 0.2021
R11003 D2_6.n9 D2_6 0.184491
R11004 D2_6.n14 D2_6 0.0740348
R11005 D2_6 D2_6.n14 0.0339615
R11006 D2_1.t18 D2_1.t11 144.929
R11007 D2_1.n23 D2_1.n22 60.7838
R11008 D2_1.t28 D2_1.t21 47.8944
R11009 D2_1.t29 D2_1.t16 47.8944
R11010 D2_1.t13 D2_1.t0 47.5387
R11011 D2_1.n4 D2_1.t4 38.8649
R11012 D2_1.n1 D2_1.t23 38.8649
R11013 D2_1.n11 D2_1.t27 38.7949
R11014 D2_1.n10 D2_1.t15 38.7949
R11015 D2_1.n6 D2_1.t26 38.7949
R11016 D2_1.n5 D2_1.t14 38.7949
R11017 D2_1.n18 D2_1.t24 32.714
R11018 D2_1.n11 D2_1.n10 31.4949
R11019 D2_1.n6 D2_1.n5 31.4949
R11020 D2_1.n3 D2_1.t9 28.8568
R11021 D2_1.n0 D2_1.t30 28.8568
R11022 D2_1.n22 D2_1.n21 25.7355
R11023 D2_1.n16 D2_1.t19 24.9839
R11024 D2_1.n19 D2_1.n18 21.0471
R11025 D2_1.t24 D2_1 20.2341
R11026 D2_1.n12 D2_1.t5 17.9416
R11027 D2_1.n7 D2_1.t12 17.9416
R11028 D2_1.t4 D2_1.n3 17.0773
R11029 D2_1.t23 D2_1.n0 17.0773
R11030 D2_1.n8 D2_1.t13 16.621
R11031 D2_1.n21 D2_1 16.3186
R11032 D2_1.n14 D2_1.n13 15.8172
R11033 D2_1.n15 D2_1.n14 15.8172
R11034 D2_1.n17 D2_1.t18 14.7032
R11035 D2_1.n20 D2_1.t33 14.5353
R11036 D2_1 D2_1.n17 13.7626
R11037 D2_1.n21 D2_1 12.9567
R11038 D2_1.n8 D2_1.t35 12.5148
R11039 D2_1.n12 D2_1.t28 11.957
R11040 D2_1.n7 D2_1.t29 11.957
R11041 D2_1.n13 D2_1.t1 11.7326
R11042 D2_1.n13 D2_1.t8 11.7326
R11043 D2_1.n14 D2_1.t7 11.7326
R11044 D2_1.n14 D2_1.t22 11.7326
R11045 D2_1.n15 D2_1.t2 11.7326
R11046 D2_1.t33 D2_1.n15 11.7326
R11047 D2_1.n19 D2_1.t17 11.6675
R11048 D2_1.n3 D2_1.t20 11.6023
R11049 D2_1.n0 D2_1.t3 11.6023
R11050 D2_1.n16 D2_1.t34 11.4552
R11051 D2_1 D2_1.n12 9.95286
R11052 D2_1 D2_1.n7 9.95286
R11053 D2_1 D2_1.n4 9.27587
R11054 D2_1 D2_1.n1 9.27587
R11055 D2_1.n24 D2_1.n23 8.99292
R11056 D2_1 D2_1.n8 8.59246
R11057 D2_1 D2_1.n20 8.19616
R11058 D2_1.n23 D2_1 7.33027
R11059 D2_1.n18 D2_1.t6 7.3005
R11060 D2_1.n10 D2_1.t32 7.3005
R11061 D2_1.t5 D2_1.n11 7.3005
R11062 D2_1.n5 D2_1.t31 7.3005
R11063 D2_1.t12 D2_1.n6 7.3005
R11064 D2_1.n4 D2_1.t10 7.3005
R11065 D2_1.n1 D2_1.t25 7.3005
R11066 D2_1.n22 D2_1.n9 3.80981
R11067 D2_1.n20 D2_1.n19 2.47729
R11068 D2_1.n17 D2_1.n16 2.45537
R11069 D2_1.n9 D2_1 1.3505
R11070 D2_1.n9 D2_1 0.194274
R11071 D2_1.n24 D2_1.n2 0.0468336
R11072 D2_1 D2_1.n24 0.0339615
R11073 D2_1.n2 D2_1 0.0115019
R11074 D2_1.n2 D2_1 0.00541341
R11075 a_29512_8496.n2 a_29512_8496.t14 39.6673
R11076 a_29512_8496.t6 a_29512_8496.n2 39.6673
R11077 a_29512_8496.n3 a_29512_8496.t10 39.3349
R11078 a_29512_8496.t8 a_29512_8496.n3 39.3349
R11079 a_29512_8496.t11 a_29512_8496.t6 31.0255
R11080 a_29512_8496.t7 a_29512_8496.t13 31.0255
R11081 a_29512_8496.t10 a_29512_8496.t11 29.1353
R11082 a_29512_8496.t13 a_29512_8496.t12 29.1353
R11083 a_29512_8496.t9 a_29512_8496.t8 29.1353
R11084 a_29512_8496.n4 a_29512_8496.t14 13.6103
R11085 a_29512_8496.n4 a_29512_8496.t9 12.9295
R11086 a_29512_8496.n0 a_29512_8496.n1 4.43082
R11087 a_29512_8496.n1 a_29512_8496.n4 8.42281
R11088 a_29512_8496.n2 a_29512_8496.t7 7.3005
R11089 a_29512_8496.n3 a_29512_8496.t12 7.3005
R11090 a_29512_8496.n1 a_29512_8496.t2 5.86791
R11091 a_29512_8496.n0 a_29512_8496.t0 4.62819
R11092 a_29512_8496.n1 a_29512_8496.t4 4.62001
R11093 a_29512_8496.n0 a_29512_8496.t3 5.02161
R11094 a_29512_8496.t1 a_29512_8496.n0 5.01918
R11095 a_29512_8496.n1 a_29512_8496.t5 4.2255
R11096 7b_counter_0.MDFF_5.LD.t82 7b_counter_0.MDFF_5.LD.t70 144.929
R11097 7b_counter_0.MDFF_5.LD.t61 7b_counter_0.MDFF_5.LD.t21 144.929
R11098 7b_counter_0.MDFF_5.LD.t83 7b_counter_0.MDFF_5.LD.t60 144.929
R11099 7b_counter_0.MDFF_5.LD.t68 7b_counter_0.MDFF_5.LD.t72 144.929
R11100 7b_counter_0.MDFF_5.LD.t11 7b_counter_0.MDFF_5.LD.t17 144.929
R11101 7b_counter_0.MDFF_5.LD.t20 7b_counter_0.MDFF_5.LD.t28 144.929
R11102 7b_counter_0.MDFF_5.LD.n2 7b_counter_0.MDFF_5.LD.n1 45.1331
R11103 7b_counter_0.MDFF_5.LD.n41 7b_counter_0.MDFF_5.LD.t24 32.714
R11104 7b_counter_0.MDFF_5.LD.n22 7b_counter_0.MDFF_5.LD.t12 32.714
R11105 7b_counter_0.MDFF_5.LD.n33 7b_counter_0.MDFF_5.LD.t25 32.714
R11106 7b_counter_0.MDFF_5.LD.n6 7b_counter_0.MDFF_5.LD.t13 32.714
R11107 7b_counter_0.MDFF_5.LD.n17 7b_counter_0.MDFF_5.LD.t26 32.714
R11108 7b_counter_0.MDFF_5.LD.n56 7b_counter_0.MDFF_5.LD.t42 32.714
R11109 7b_counter_0.MDFF_5.LD.n31 7b_counter_0.MDFF_5.LD.t34 25.1498
R11110 7b_counter_0.MDFF_5.LD.n4 7b_counter_0.MDFF_5.LD.t41 25.0633
R11111 7b_counter_0.MDFF_5.LD.n15 7b_counter_0.MDFF_5.LD.t69 25.0633
R11112 7b_counter_0.MDFF_5.LD.n54 7b_counter_0.MDFF_5.LD.t67 25.0633
R11113 7b_counter_0.MDFF_5.LD.n39 7b_counter_0.MDFF_5.LD.t43 24.9839
R11114 7b_counter_0.MDFF_5.LD.n20 7b_counter_0.MDFF_5.LD.t16 24.9839
R11115 7b_counter_0.MDFF_5.LD.n42 7b_counter_0.MDFF_5.LD.n41 21.0471
R11116 7b_counter_0.MDFF_5.LD.n23 7b_counter_0.MDFF_5.LD.n22 21.0471
R11117 7b_counter_0.MDFF_5.LD.n34 7b_counter_0.MDFF_5.LD.n33 21.0471
R11118 7b_counter_0.MDFF_5.LD.n7 7b_counter_0.MDFF_5.LD.n6 21.0471
R11119 7b_counter_0.MDFF_5.LD.n18 7b_counter_0.MDFF_5.LD.n17 21.0471
R11120 7b_counter_0.MDFF_5.LD.n57 7b_counter_0.MDFF_5.LD.n56 21.0471
R11121 7b_counter_0.MDFF_5.LD.t24 7b_counter_0.MDFF_5.LD 20.2341
R11122 7b_counter_0.MDFF_5.LD.t12 7b_counter_0.MDFF_5.LD 20.2341
R11123 7b_counter_0.MDFF_5.LD.t25 7b_counter_0.MDFF_5.LD 20.2341
R11124 7b_counter_0.MDFF_5.LD.t13 7b_counter_0.MDFF_5.LD 20.2328
R11125 7b_counter_0.MDFF_5.LD.t26 7b_counter_0.MDFF_5.LD 20.2328
R11126 7b_counter_0.MDFF_5.LD.t42 7b_counter_0.MDFF_5.LD 20.2328
R11127 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n3 18.9288
R11128 7b_counter_0.MDFF_5.LD.n2 7b_counter_0.MDFF_5.LD 18.294
R11129 7b_counter_0.MDFF_5.LD.n37 7b_counter_0.MDFF_5.LD.n36 15.8172
R11130 7b_counter_0.MDFF_5.LD.n38 7b_counter_0.MDFF_5.LD.n37 15.8172
R11131 7b_counter_0.MDFF_5.LD.n25 7b_counter_0.MDFF_5.LD.n24 15.8172
R11132 7b_counter_0.MDFF_5.LD.n26 7b_counter_0.MDFF_5.LD.n25 15.8172
R11133 7b_counter_0.MDFF_5.LD.n29 7b_counter_0.MDFF_5.LD.n28 15.8172
R11134 7b_counter_0.MDFF_5.LD.n30 7b_counter_0.MDFF_5.LD.n29 15.8172
R11135 7b_counter_0.MDFF_5.LD.n9 7b_counter_0.MDFF_5.LD.n8 15.8172
R11136 7b_counter_0.MDFF_5.LD.n10 7b_counter_0.MDFF_5.LD.n9 15.8172
R11137 7b_counter_0.MDFF_5.LD.n13 7b_counter_0.MDFF_5.LD.n12 15.8172
R11138 7b_counter_0.MDFF_5.LD.n14 7b_counter_0.MDFF_5.LD.n13 15.8172
R11139 7b_counter_0.MDFF_5.LD.n52 7b_counter_0.MDFF_5.LD.n51 15.8172
R11140 7b_counter_0.MDFF_5.LD.n53 7b_counter_0.MDFF_5.LD.n52 15.8172
R11141 7b_counter_0.MDFF_5.LD.n21 7b_counter_0.MDFF_5.LD.t61 14.7678
R11142 7b_counter_0.MDFF_5.LD.n5 7b_counter_0.MDFF_5.LD.t68 14.7678
R11143 7b_counter_0.MDFF_5.LD.n40 7b_counter_0.MDFF_5.LD.t82 14.7032
R11144 7b_counter_0.MDFF_5.LD.n32 7b_counter_0.MDFF_5.LD.t83 14.7032
R11145 7b_counter_0.MDFF_5.LD.n16 7b_counter_0.MDFF_5.LD.t11 14.7032
R11146 7b_counter_0.MDFF_5.LD.n55 7b_counter_0.MDFF_5.LD.t20 14.7032
R11147 7b_counter_0.MDFF_5.LD.n43 7b_counter_0.MDFF_5.LD.t84 14.5353
R11148 7b_counter_0.MDFF_5.LD.n27 7b_counter_0.MDFF_5.LD.t77 14.5353
R11149 7b_counter_0.MDFF_5.LD.n35 7b_counter_0.MDFF_5.LD.t85 14.5353
R11150 7b_counter_0.MDFF_5.LD.n11 7b_counter_0.MDFF_5.LD.t45 14.5353
R11151 7b_counter_0.MDFF_5.LD.n19 7b_counter_0.MDFF_5.LD.t55 14.5353
R11152 7b_counter_0.MDFF_5.LD.n58 7b_counter_0.MDFF_5.LD.t56 14.5353
R11153 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n40 13.7626
R11154 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n21 13.7626
R11155 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n32 13.7626
R11156 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n5 13.7626
R11157 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n16 13.7626
R11158 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n55 13.7626
R11159 7b_counter_0.MDFF_5.LD.n36 7b_counter_0.MDFF_5.LD.t27 11.7326
R11160 7b_counter_0.MDFF_5.LD.n36 7b_counter_0.MDFF_5.LD.t57 11.7326
R11161 7b_counter_0.MDFF_5.LD.n37 7b_counter_0.MDFF_5.LD.t48 11.7326
R11162 7b_counter_0.MDFF_5.LD.n37 7b_counter_0.MDFF_5.LD.t80 11.7326
R11163 7b_counter_0.MDFF_5.LD.n38 7b_counter_0.MDFF_5.LD.t9 11.7326
R11164 7b_counter_0.MDFF_5.LD.t84 7b_counter_0.MDFF_5.LD.n38 11.7326
R11165 7b_counter_0.MDFF_5.LD.n24 7b_counter_0.MDFF_5.LD.t47 11.7326
R11166 7b_counter_0.MDFF_5.LD.n24 7b_counter_0.MDFF_5.LD.t40 11.7326
R11167 7b_counter_0.MDFF_5.LD.n25 7b_counter_0.MDFF_5.LD.t53 11.7326
R11168 7b_counter_0.MDFF_5.LD.n25 7b_counter_0.MDFF_5.LD.t49 11.7326
R11169 7b_counter_0.MDFF_5.LD.n26 7b_counter_0.MDFF_5.LD.t76 11.7326
R11170 7b_counter_0.MDFF_5.LD.t77 7b_counter_0.MDFF_5.LD.n26 11.7326
R11171 7b_counter_0.MDFF_5.LD.n28 7b_counter_0.MDFF_5.LD.t38 11.7326
R11172 7b_counter_0.MDFF_5.LD.n28 7b_counter_0.MDFF_5.LD.t58 11.7326
R11173 7b_counter_0.MDFF_5.LD.n29 7b_counter_0.MDFF_5.LD.t81 11.7326
R11174 7b_counter_0.MDFF_5.LD.n29 7b_counter_0.MDFF_5.LD.t66 11.7326
R11175 7b_counter_0.MDFF_5.LD.n30 7b_counter_0.MDFF_5.LD.t18 11.7326
R11176 7b_counter_0.MDFF_5.LD.t85 7b_counter_0.MDFF_5.LD.n30 11.7326
R11177 7b_counter_0.MDFF_5.LD.n8 7b_counter_0.MDFF_5.LD.t51 11.7326
R11178 7b_counter_0.MDFF_5.LD.n8 7b_counter_0.MDFF_5.LD.t44 11.7326
R11179 7b_counter_0.MDFF_5.LD.n9 7b_counter_0.MDFF_5.LD.t75 11.7326
R11180 7b_counter_0.MDFF_5.LD.n9 7b_counter_0.MDFF_5.LD.t73 11.7326
R11181 7b_counter_0.MDFF_5.LD.n10 7b_counter_0.MDFF_5.LD.t39 11.7326
R11182 7b_counter_0.MDFF_5.LD.t45 7b_counter_0.MDFF_5.LD.n10 11.7326
R11183 7b_counter_0.MDFF_5.LD.n12 7b_counter_0.MDFF_5.LD.t50 11.7326
R11184 7b_counter_0.MDFF_5.LD.n12 7b_counter_0.MDFF_5.LD.t62 11.7326
R11185 7b_counter_0.MDFF_5.LD.n13 7b_counter_0.MDFF_5.LD.t86 11.7326
R11186 7b_counter_0.MDFF_5.LD.n13 7b_counter_0.MDFF_5.LD.t78 11.7326
R11187 7b_counter_0.MDFF_5.LD.n14 7b_counter_0.MDFF_5.LD.t71 11.7326
R11188 7b_counter_0.MDFF_5.LD.t55 7b_counter_0.MDFF_5.LD.n14 11.7326
R11189 7b_counter_0.MDFF_5.LD.n51 7b_counter_0.MDFF_5.LD.t46 11.7326
R11190 7b_counter_0.MDFF_5.LD.n51 7b_counter_0.MDFF_5.LD.t74 11.7326
R11191 7b_counter_0.MDFF_5.LD.n52 7b_counter_0.MDFF_5.LD.t35 11.7326
R11192 7b_counter_0.MDFF_5.LD.n52 7b_counter_0.MDFF_5.LD.t65 11.7326
R11193 7b_counter_0.MDFF_5.LD.n53 7b_counter_0.MDFF_5.LD.t79 11.7326
R11194 7b_counter_0.MDFF_5.LD.t56 7b_counter_0.MDFF_5.LD.n53 11.7326
R11195 7b_counter_0.MDFF_5.LD.n42 7b_counter_0.MDFF_5.LD.t63 11.6675
R11196 7b_counter_0.MDFF_5.LD.n23 7b_counter_0.MDFF_5.LD.t37 11.6675
R11197 7b_counter_0.MDFF_5.LD.n34 7b_counter_0.MDFF_5.LD.t64 11.6675
R11198 7b_counter_0.MDFF_5.LD.n7 7b_counter_0.MDFF_5.LD.t10 11.6675
R11199 7b_counter_0.MDFF_5.LD.n18 7b_counter_0.MDFF_5.LD.t22 11.6675
R11200 7b_counter_0.MDFF_5.LD.n57 7b_counter_0.MDFF_5.LD.t23 11.6675
R11201 7b_counter_0.MDFF_5.LD.n39 7b_counter_0.MDFF_5.LD.t31 11.4552
R11202 7b_counter_0.MDFF_5.LD.n31 7b_counter_0.MDFF_5.LD.t32 11.4552
R11203 7b_counter_0.MDFF_5.LD.n15 7b_counter_0.MDFF_5.LD.t36 11.4552
R11204 7b_counter_0.MDFF_5.LD.n54 7b_counter_0.MDFF_5.LD.t59 11.4552
R11205 7b_counter_0.MDFF_5.LD.n20 7b_counter_0.MDFF_5.LD.t15 11.3906
R11206 7b_counter_0.MDFF_5.LD.n4 7b_counter_0.MDFF_5.LD.t19 11.3906
R11207 7b_counter_0.MDFF_5.LD.n0 7b_counter_0.MDFF_5.LD.n50 9.69373
R11208 7b_counter_0.MDFF_5.LD.n46 7b_counter_0.MDFF_5.LD.n45 9.64291
R11209 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n43 8.19616
R11210 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n27 8.19616
R11211 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n35 8.19616
R11212 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n11 8.19616
R11213 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n19 8.19616
R11214 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.LD.n58 8.19616
R11215 7b_counter_0.MDFF_5.LD.n41 7b_counter_0.MDFF_5.LD.t54 7.3005
R11216 7b_counter_0.MDFF_5.LD.n22 7b_counter_0.MDFF_5.LD.t14 7.3005
R11217 7b_counter_0.MDFF_5.LD.n33 7b_counter_0.MDFF_5.LD.t30 7.3005
R11218 7b_counter_0.MDFF_5.LD.n6 7b_counter_0.MDFF_5.LD.t33 7.3005
R11219 7b_counter_0.MDFF_5.LD.n17 7b_counter_0.MDFF_5.LD.t52 7.3005
R11220 7b_counter_0.MDFF_5.LD.n56 7b_counter_0.MDFF_5.LD.t29 7.3005
R11221 7b_counter_0.MDFF_5.LD.n45 7b_counter_0.MDFF_5.LD.t7 4.63638
R11222 7b_counter_0.MDFF_5.LD.n1 7b_counter_0.MDFF_5.LD.t2 4.2255
R11223 7b_counter_0.MDFF_5.LD.n0 7b_counter_0.MDFF_5.LD.t5 4.2255
R11224 7b_counter_0.MDFF_5.LD.n46 7b_counter_0.MDFF_5.LD.n44 3.17388
R11225 7b_counter_0.MDFF_5.LD.n50 7b_counter_0.MDFF_5.LD.n49 2.6005
R11226 7b_counter_0.MDFF_5.LD.n48 7b_counter_0.MDFF_5.LD.n47 2.6005
R11227 7b_counter_0.MDFF_5.LD.n43 7b_counter_0.MDFF_5.LD.n42 2.47729
R11228 7b_counter_0.MDFF_5.LD.n27 7b_counter_0.MDFF_5.LD.n23 2.47729
R11229 7b_counter_0.MDFF_5.LD.n35 7b_counter_0.MDFF_5.LD.n34 2.47729
R11230 7b_counter_0.MDFF_5.LD.n11 7b_counter_0.MDFF_5.LD.n7 2.47729
R11231 7b_counter_0.MDFF_5.LD.n19 7b_counter_0.MDFF_5.LD.n18 2.47729
R11232 7b_counter_0.MDFF_5.LD.n58 7b_counter_0.MDFF_5.LD.n57 2.47729
R11233 7b_counter_0.MDFF_5.LD.n40 7b_counter_0.MDFF_5.LD.n39 2.45537
R11234 7b_counter_0.MDFF_5.LD.n21 7b_counter_0.MDFF_5.LD.n20 2.45537
R11235 7b_counter_0.MDFF_5.LD.n32 7b_counter_0.MDFF_5.LD.n31 2.45537
R11236 7b_counter_0.MDFF_5.LD.n5 7b_counter_0.MDFF_5.LD.n4 2.45537
R11237 7b_counter_0.MDFF_5.LD.n16 7b_counter_0.MDFF_5.LD.n15 2.45537
R11238 7b_counter_0.MDFF_5.LD.n55 7b_counter_0.MDFF_5.LD.n54 2.45537
R11239 7b_counter_0.MDFF_5.LD.n47 7b_counter_0.MDFF_5.LD.t1 1.6255
R11240 7b_counter_0.MDFF_5.LD.n47 7b_counter_0.MDFF_5.LD.t3 1.6255
R11241 7b_counter_0.MDFF_5.LD.n49 7b_counter_0.MDFF_5.LD.t4 1.6255
R11242 7b_counter_0.MDFF_5.LD.n49 7b_counter_0.MDFF_5.LD.t0 1.6255
R11243 7b_counter_0.MDFF_5.LD.n44 7b_counter_0.MDFF_5.LD.t6 1.463
R11244 7b_counter_0.MDFF_5.LD.n44 7b_counter_0.MDFF_5.LD.t8 1.463
R11245 7b_counter_0.MDFF_5.LD.n3 7b_counter_0.MDFF_5.LD 1.27725
R11246 7b_counter_0.MDFF_5.LD.n3 7b_counter_0.MDFF_5.LD 1.27582
R11247 7b_counter_0.MDFF_5.LD.n50 7b_counter_0.MDFF_5.LD.n48 0.925383
R11248 7b_counter_0.MDFF_5.LD.n3 7b_counter_0.MDFF_5.LD.n2 0.834839
R11249 7b_counter_0.MDFF_5.LD.n1 7b_counter_0.MDFF_5.LD.n0 0.833778
R11250 7b_counter_0.MDFF_5.LD.n48 7b_counter_0.MDFF_5.LD.n46 0.805215
R11251 7b_counter_0.MDFF_5.LD.n45 7b_counter_0.MDFF_5.LD.n1 0.805215
R11252 D2_2.t8 D2_2.t23 47.8944
R11253 D2_2.t16 D2_2.t3 47.8944
R11254 D2_2.t25 D2_2.t20 47.5387
R11255 D2_2.t9 D2_2.t1 47.5387
R11256 D2_2.n16 D2_2.t2 38.8649
R11257 D2_2.n1 D2_2.t12 38.8649
R11258 D2_2.n3 D2_2.t7 38.7949
R11259 D2_2.n2 D2_2.t5 38.7949
R11260 D2_2.n8 D2_2.t18 38.7949
R11261 D2_2.n7 D2_2.t15 38.7949
R11262 D2_2.n3 D2_2.n2 31.4949
R11263 D2_2.n8 D2_2.n7 31.4949
R11264 D2_2.n15 D2_2.t10 28.8568
R11265 D2_2.n0 D2_2.t19 28.8568
R11266 D2_2.n13 D2_2.n12 21.7014
R11267 D2_2.n4 D2_2.t24 17.9416
R11268 D2_2.n9 D2_2.t6 17.9416
R11269 D2_2.t2 D2_2.n15 17.0773
R11270 D2_2.t12 D2_2.n0 17.0773
R11271 D2_2.n5 D2_2.t25 16.621
R11272 D2_2.n10 D2_2.t9 16.621
R11273 D2_2.n12 D2_2.n6 14.1695
R11274 D2_2.n5 D2_2.t4 12.5148
R11275 D2_2.n10 D2_2.t14 12.5148
R11276 D2_2.n4 D2_2.t8 11.957
R11277 D2_2.n9 D2_2.t16 11.957
R11278 D2_2.n12 D2_2.n11 11.825
R11279 D2_2.n15 D2_2.t17 11.6023
R11280 D2_2.n0 D2_2.t21 11.6023
R11281 D2_2 D2_2.n4 9.95286
R11282 D2_2 D2_2.n9 9.95286
R11283 D2_2 D2_2.n16 9.27587
R11284 D2_2 D2_2.n1 9.27587
R11285 D2_2 D2_2.n5 8.59246
R11286 D2_2 D2_2.n10 8.59246
R11287 D2_2.n14 D2_2.n13 7.97639
R11288 D2_2.n16 D2_2.t0 7.3005
R11289 D2_2.n2 D2_2.t13 7.3005
R11290 D2_2.t24 D2_2.n3 7.3005
R11291 D2_2.n7 D2_2.t22 7.3005
R11292 D2_2.t6 D2_2.n8 7.3005
R11293 D2_2.n1 D2_2.t11 7.3005
R11294 D2_2.n13 D2_2 6.09406
R11295 D2_2.n11 D2_2 1.36924
R11296 D2_2.n6 D2_2 1.36028
R11297 D2_2.n6 D2_2 0.184491
R11298 D2_2.n11 D2_2 0.108743
R11299 D2_2.n14 D2_2 0.0738303
R11300 D2_2 D2_2.n14 0.0339615
R11301 LD.t26 LD.t55 144.929
R11302 LD.t23 LD.t54 144.929
R11303 LD.t86 LD.t27 144.929
R11304 LD.t34 LD.t58 144.929
R11305 LD.t18 LD.t50 144.929
R11306 LD.t79 LD.t21 144.929
R11307 LD.n18 LD.n17 55.3638
R11308 LD.n32 LD.n31 32.8505
R11309 LD.n33 LD.n32 32.8505
R11310 LD.n59 LD.n58 32.8505
R11311 LD.n60 LD.n59 32.8505
R11312 LD.n5 LD.t60 32.714
R11313 LD.n21 LD.t41 32.714
R11314 LD.n29 LD.t51 32.714
R11315 LD.n41 LD.t46 32.714
R11316 LD.n47 LD.t32 32.714
R11317 LD.n56 LD.t45 32.714
R11318 LD.n3 LD.t33 24.9839
R11319 LD.n19 LD.t39 24.9839
R11320 LD.n27 LD.t15 24.9839
R11321 LD.n39 LD.t36 24.9839
R11322 LD.n45 LD.t35 24.9839
R11323 LD.n54 LD.t14 24.9839
R11324 LD.n6 LD.n5 21.0471
R11325 LD.n22 LD.n21 21.0471
R11326 LD.n30 LD.n29 21.0471
R11327 LD.n42 LD.n41 21.0471
R11328 LD.n48 LD.n47 21.0471
R11329 LD.n57 LD.n56 21.0471
R11330 LD.t60 LD 20.2341
R11331 LD.t41 LD 20.2341
R11332 LD.t51 LD 20.2341
R11333 LD.t46 LD 20.2341
R11334 LD.t32 LD 20.2341
R11335 LD.t45 LD 20.2341
R11336 LD.n35 LD 20.116
R11337 LD.n53 LD 18.3333
R11338 LD.n1 LD.n0 15.8172
R11339 LD.n2 LD.n1 15.8172
R11340 LD.n24 LD.n23 15.8172
R11341 LD.n25 LD.n24 15.8172
R11342 LD.n37 LD.n36 15.8172
R11343 LD.n38 LD.n37 15.8172
R11344 LD.n50 LD.n49 15.8172
R11345 LD.n51 LD.n50 15.8172
R11346 LD.n20 LD.t23 14.7678
R11347 LD.n28 LD.t86 14.7678
R11348 LD.n46 LD.t18 14.7678
R11349 LD.n55 LD.t79 14.7678
R11350 LD.n4 LD.t26 14.7032
R11351 LD.n40 LD.t34 14.7032
R11352 LD.n7 LD.t38 14.5353
R11353 LD.n26 LD.t52 14.5353
R11354 LD.n34 LD.t37 14.5353
R11355 LD.n43 LD.t17 14.5353
R11356 LD.n52 LD.t48 14.5353
R11357 LD.n61 LD.t28 14.5353
R11358 LD LD.n4 13.7626
R11359 LD LD.n20 13.7626
R11360 LD LD.n28 13.7626
R11361 LD LD.n40 13.7626
R11362 LD LD.n46 13.7626
R11363 LD LD.n55 13.7626
R11364 LD.n0 LD.t24 11.7326
R11365 LD.n0 LD.t84 11.7326
R11366 LD.n1 LD.t49 11.7326
R11367 LD.n1 LD.t30 11.7326
R11368 LD.n2 LD.t80 11.7326
R11369 LD.t38 LD.n2 11.7326
R11370 LD.n23 LD.t74 11.7326
R11371 LD.n23 LD.t13 11.7326
R11372 LD.n24 LD.t19 11.7326
R11373 LD.n24 LD.t57 11.7326
R11374 LD.n25 LD.t44 11.7326
R11375 LD.t52 LD.n25 11.7326
R11376 LD.n36 LD.t85 11.7326
R11377 LD.n36 LD.t68 11.7326
R11378 LD.n37 LD.t31 11.7326
R11379 LD.n37 LD.t11 11.7326
R11380 LD.n38 LD.t40 11.7326
R11381 LD.t17 LD.n38 11.7326
R11382 LD.n49 LD.t70 11.7326
R11383 LD.n49 LD.t69 11.7326
R11384 LD.n50 LD.t16 11.7326
R11385 LD.n50 LD.t12 11.7326
R11386 LD.n51 LD.t42 11.7326
R11387 LD.t48 LD.n51 11.7326
R11388 LD.n6 LD.t10 11.6675
R11389 LD.n22 LD.t9 11.6675
R11390 LD.n30 LD.t75 11.6675
R11391 LD.n42 LD.t72 11.6675
R11392 LD.n48 LD.t81 11.6675
R11393 LD.n57 LD.t71 11.6675
R11394 LD.n3 LD.t59 11.4552
R11395 LD.n39 LD.t61 11.4552
R11396 LD.n19 LD.t63 11.3906
R11397 LD.n27 LD.t47 11.3906
R11398 LD.n45 LD.t62 11.3906
R11399 LD.n54 LD.t43 11.3906
R11400 LD.n33 LD.t53 10.1684
R11401 LD.n31 LD.t77 10.1684
R11402 LD.n31 LD.t83 10.1684
R11403 LD.n32 LD.t65 10.1684
R11404 LD.n32 LD.t29 10.1684
R11405 LD.t37 LD.n33 10.1684
R11406 LD.n60 LD.t25 10.1684
R11407 LD.n58 LD.t76 10.1684
R11408 LD.n58 LD.t78 10.1684
R11409 LD.n59 LD.t20 10.1684
R11410 LD.n59 LD.t22 10.1684
R11411 LD.t28 LD.n60 10.1684
R11412 LD.n10 LD.n8 9.69373
R11413 LD.n15 LD.n14 9.64291
R11414 LD LD.n7 8.19616
R11415 LD LD.n26 8.19616
R11416 LD LD.n34 8.19616
R11417 LD LD.n43 8.19616
R11418 LD LD.n52 8.19616
R11419 LD LD.n61 8.19616
R11420 LD.n5 LD.t82 7.3005
R11421 LD.n21 LD.t64 7.3005
R11422 LD.n29 LD.t73 7.3005
R11423 LD.n41 LD.t67 7.3005
R11424 LD.n47 LD.t56 7.3005
R11425 LD.n56 LD.t66 7.3005
R11426 LD.n15 LD.t0 4.63638
R11427 LD.n16 LD.t1 4.2255
R11428 LD.n8 LD.t6 4.2255
R11429 LD.n44 LD 4.02178
R11430 LD.n14 LD.n13 3.17388
R11431 LD.n12 LD.n11 2.6005
R11432 LD.n10 LD.n9 2.6005
R11433 LD.n7 LD.n6 2.47729
R11434 LD.n26 LD.n22 2.47729
R11435 LD.n34 LD.n30 2.47729
R11436 LD.n43 LD.n42 2.47729
R11437 LD.n52 LD.n48 2.47729
R11438 LD.n61 LD.n57 2.47729
R11439 LD.n4 LD.n3 2.45537
R11440 LD.n20 LD.n19 2.45537
R11441 LD.n28 LD.n27 2.45537
R11442 LD.n40 LD.n39 2.45537
R11443 LD.n46 LD.n45 2.45537
R11444 LD.n55 LD.n54 2.45537
R11445 LD LD.n35 1.93071
R11446 LD LD.n62 1.93071
R11447 LD.n53 LD.n44 1.92305
R11448 LD.n62 LD.n53 1.78327
R11449 LD.n9 LD.t7 1.6255
R11450 LD.n9 LD.t8 1.6255
R11451 LD.n11 LD.t3 1.6255
R11452 LD.n11 LD.t5 1.6255
R11453 LD.n13 LD.t2 1.463
R11454 LD.n13 LD.t4 1.463
R11455 LD.n12 LD.n10 0.925383
R11456 LD.n16 LD.n15 0.805215
R11457 LD.n14 LD.n12 0.805215
R11458 LD LD.n18 0.643813
R11459 LD.n17 LD.n8 0.460082
R11460 LD.n17 LD.n16 0.374196
R11461 LD.n18 LD 0.193357
R11462 LD.n35 LD 0.181929
R11463 LD.n44 LD 0.181929
R11464 LD.n62 LD 0.181929
R11465 D2_7.t12 D2_7.t2 47.8944
R11466 D2_7.t18 D2_7.t8 47.8944
R11467 D2_7.t4 D2_7.t16 47.5387
R11468 D2_7.t10 D2_7.t25 47.5387
R11469 D2_7.n3 D2_7.t13 38.8649
R11470 D2_7.n1 D2_7.t15 38.8649
R11471 D2_7.n6 D2_7.t3 38.7949
R11472 D2_7.n5 D2_7.t6 38.7949
R11473 D2_7.n10 D2_7.t11 38.7949
R11474 D2_7.n9 D2_7.t14 38.7949
R11475 D2_7.n14 D2_7.n8 33.9151
R11476 D2_7.n6 D2_7.n5 31.4949
R11477 D2_7.n10 D2_7.n9 31.4949
R11478 D2_7.n2 D2_7.t24 28.8568
R11479 D2_7.n0 D2_7.t22 28.8568
R11480 D2_7.n15 D2_7.n14 22.2998
R11481 D2_7.n7 D2_7.t21 17.9416
R11482 D2_7.n11 D2_7.t7 17.9416
R11483 D2_7.t13 D2_7.n2 17.0773
R11484 D2_7.t15 D2_7.n0 17.0773
R11485 D2_7.n4 D2_7.t4 16.621
R11486 D2_7.n12 D2_7.t10 16.621
R11487 D2_7.n14 D2_7.n13 16.1008
R11488 D2_7.n4 D2_7.t19 12.5148
R11489 D2_7.n12 D2_7.t5 12.5148
R11490 D2_7.n7 D2_7.t12 11.957
R11491 D2_7.n11 D2_7.t18 11.957
R11492 D2_7.n2 D2_7.t1 11.6023
R11493 D2_7.n0 D2_7.t0 11.6023
R11494 D2_7.n15 D2_7 11.489
R11495 D2_7 D2_7.n7 9.95286
R11496 D2_7 D2_7.n11 9.95286
R11497 D2_7 D2_7.n3 9.27587
R11498 D2_7 D2_7.n1 9.27587
R11499 D2_7 D2_7.n4 8.59246
R11500 D2_7 D2_7.n12 8.59246
R11501 D2_7.n5 D2_7.t9 7.3005
R11502 D2_7.t21 D2_7.n6 7.3005
R11503 D2_7.n9 D2_7.t17 7.3005
R11504 D2_7.t7 D2_7.n10 7.3005
R11505 D2_7.n3 D2_7.t20 7.3005
R11506 D2_7.n1 D2_7.t23 7.3005
R11507 D2_7.n16 D2_7.n15 2.69384
R11508 D2_7.n13 D2_7 1.3818
R11509 D2_7.n8 D2_7 1.31528
R11510 D2_7.n13 D2_7 0.16297
R11511 D2_7.n8 D2_7 0.137535
R11512 D2_7 D2_7.n16 0.113082
R11513 D2_7.n16 D2_7 0.00371263
R11514 mux_magic_0.IN2.t3 mux_magic_0.IN2.t6 47.8944
R11515 mux_magic_0.IN2.n1 mux_magic_0.IN2.t8 38.8649
R11516 mux_magic_0.IN2.n2 mux_magic_0.IN2.t5 38.7949
R11517 mux_magic_0.IN2.n3 mux_magic_0.IN2.t7 38.7949
R11518 mux_magic_0.IN2.n3 mux_magic_0.IN2.n2 31.4949
R11519 mux_magic_0.IN2.n0 mux_magic_0.IN2.t9 28.8568
R11520 mux_magic_0.IN2.n4 mux_magic_0.IN2.t10 17.9416
R11521 mux_magic_0.IN2.t8 mux_magic_0.IN2.n0 17.0773
R11522 mux_magic_0.IN2.t1 mux_magic_0.IN2 12.3547
R11523 mux_magic_0.IN2.n4 mux_magic_0.IN2.t3 11.957
R11524 mux_magic_0.IN2.n0 mux_magic_0.IN2.t4 11.6023
R11525 mux_magic_0.IN2 mux_magic_0.IN2.n4 9.95929
R11526 mux_magic_0.IN2 mux_magic_0.IN2.n1 9.47416
R11527 mux_magic_0.IN2.n2 mux_magic_0.IN2.t11 7.3005
R11528 mux_magic_0.IN2.t10 mux_magic_0.IN2.n3 7.3005
R11529 mux_magic_0.IN2.n1 mux_magic_0.IN2.t12 7.3005
R11530 mux_magic_0.IN2.t1 mux_magic_0.IN2.t0 4.93572
R11531 mux_magic_0.IN2.t1 mux_magic_0.IN2 4.15573
R11532 mux_magic_0.IN2.t1 mux_magic_0.IN2.t2 3.6455
R11533 7b_counter_0.NAND_magic_0.A.t12 7b_counter_0.NAND_magic_0.A.t15 47.8944
R11534 7b_counter_0.NAND_magic_0.A.t9 7b_counter_0.NAND_magic_0.A.t21 47.8944
R11535 7b_counter_0.NAND_magic_0.A.n9 7b_counter_0.NAND_magic_0.A.t10 38.7949
R11536 7b_counter_0.NAND_magic_0.A.n10 7b_counter_0.NAND_magic_0.A.t20 38.7949
R11537 7b_counter_0.NAND_magic_0.A.n3 7b_counter_0.NAND_magic_0.A.t18 38.7949
R11538 7b_counter_0.NAND_magic_0.A.n2 7b_counter_0.NAND_magic_0.A.t14 38.7949
R11539 7b_counter_0.NAND_magic_0.A.n5 7b_counter_0.NAND_magic_0.A.t19 31.9191
R11540 7b_counter_0.NAND_magic_0.A.n10 7b_counter_0.NAND_magic_0.A.n9 31.4949
R11541 7b_counter_0.NAND_magic_0.A.n3 7b_counter_0.NAND_magic_0.A.n2 31.4949
R11542 7b_counter_0.NAND_magic_0.A.n6 7b_counter_0.NAND_magic_0.A.t13 31.1267
R11543 7b_counter_0.NAND_magic_0.A.n0 7b_counter_0.NAND_magic_0.A.n8 19.1157
R11544 7b_counter_0.NAND_magic_0.A.n11 7b_counter_0.NAND_magic_0.A.t7 17.9416
R11545 7b_counter_0.NAND_magic_0.A.n4 7b_counter_0.NAND_magic_0.A.t6 17.9416
R11546 7b_counter_0.NAND_magic_0.A.n11 7b_counter_0.NAND_magic_0.A.t12 11.957
R11547 7b_counter_0.NAND_magic_0.A.n4 7b_counter_0.NAND_magic_0.A.t9 11.957
R11548 7b_counter_0.NAND_magic_0.A.n6 7b_counter_0.NAND_magic_0.A.t11 10.9505
R11549 7b_counter_0.NAND_magic_0.A.n5 7b_counter_0.NAND_magic_0.A.t16 10.3639
R11550 7b_counter_0.NAND_magic_0.A 7b_counter_0.NAND_magic_0.A.n4 9.96162
R11551 7b_counter_0.NAND_magic_0.A 7b_counter_0.NAND_magic_0.A.n11 9.95929
R11552 7b_counter_0.NAND_magic_0.A 7b_counter_0.NAND_magic_0.A.n7 8.22152
R11553 7b_counter_0.NAND_magic_0.A.n8 7b_counter_0.NAND_magic_0.A 7.60603
R11554 7b_counter_0.NAND_magic_0.A.n9 7b_counter_0.NAND_magic_0.A.t8 7.3005
R11555 7b_counter_0.NAND_magic_0.A.t7 7b_counter_0.NAND_magic_0.A.n10 7.3005
R11556 7b_counter_0.NAND_magic_0.A.n2 7b_counter_0.NAND_magic_0.A.t17 7.3005
R11557 7b_counter_0.NAND_magic_0.A.t6 7b_counter_0.NAND_magic_0.A.n3 7.3005
R11558 7b_counter_0.NAND_magic_0.A.n7 7b_counter_0.NAND_magic_0.A.n5 6.32282
R11559 7b_counter_0.NAND_magic_0.A.n7 7b_counter_0.NAND_magic_0.A.n6 4.75854
R11560 7b_counter_0.NAND_magic_0.A.n1 7b_counter_0.NAND_magic_0.A.n12 3.6455
R11561 7b_counter_0.NAND_magic_0.A.n1 7b_counter_0.NAND_magic_0.A.n13 3.31072
R11562 7b_counter_0.NAND_magic_0.A.n1 7b_counter_0.NAND_magic_0.A.n14 2.90572
R11563 7b_counter_0.NAND_magic_0.A.n8 7b_counter_0.NAND_magic_0.A 2.29941
R11564 7b_counter_0.NAND_magic_0.A.n13 7b_counter_0.NAND_magic_0.A.t1 1.6255
R11565 7b_counter_0.NAND_magic_0.A.n13 7b_counter_0.NAND_magic_0.A.t0 1.6255
R11566 7b_counter_0.NAND_magic_0.A.n14 7b_counter_0.NAND_magic_0.A.t3 1.6255
R11567 7b_counter_0.NAND_magic_0.A.n14 7b_counter_0.NAND_magic_0.A.t2 1.6255
R11568 7b_counter_0.NAND_magic_0.A.n12 7b_counter_0.NAND_magic_0.A.t5 1.463
R11569 7b_counter_0.NAND_magic_0.A.n12 7b_counter_0.NAND_magic_0.A.t4 1.463
R11570 7b_counter_0.NAND_magic_0.A.n0 7b_counter_0.NAND_magic_0.A 1.25072
R11571 7b_counter_0.NAND_magic_0.A.n1 7b_counter_0.NAND_magic_0.A.n0 1.22536
R11572 DFF_magic_0.D.n12 DFF_magic_0.D.t38 39.8579
R11573 DFF_magic_0.D.t29 DFF_magic_0.D.n12 39.8579
R11574 DFF_magic_0.D.n8 DFF_magic_0.D.t28 39.8579
R11575 DFF_magic_0.D.t16 DFF_magic_0.D.n8 39.8579
R11576 DFF_magic_0.D.n4 DFF_magic_0.D.t36 39.8579
R11577 DFF_magic_0.D.t32 DFF_magic_0.D.n4 39.8579
R11578 DFF_magic_0.D.n13 DFF_magic_0.D.t14 39.3349
R11579 DFF_magic_0.D.t26 DFF_magic_0.D.n13 39.3349
R11580 DFF_magic_0.D.n9 DFF_magic_0.D.t30 39.3349
R11581 DFF_magic_0.D.t12 DFF_magic_0.D.n9 39.3349
R11582 DFF_magic_0.D.n5 DFF_magic_0.D.t18 39.3349
R11583 DFF_magic_0.D.t22 DFF_magic_0.D.n5 39.3349
R11584 DFF_magic_0.D.t15 DFF_magic_0.D.t29 31.0255
R11585 DFF_magic_0.D.t37 DFF_magic_0.D.t25 31.0255
R11586 DFF_magic_0.D.t31 DFF_magic_0.D.t16 31.0255
R11587 DFF_magic_0.D.t17 DFF_magic_0.D.t34 31.0255
R11588 DFF_magic_0.D.t19 DFF_magic_0.D.t32 31.0255
R11589 DFF_magic_0.D.t35 DFF_magic_0.D.t21 31.0255
R11590 DFF_magic_0.D.t14 DFF_magic_0.D.t15 29.1353
R11591 DFF_magic_0.D.t25 DFF_magic_0.D.t24 29.1353
R11592 DFF_magic_0.D.t27 DFF_magic_0.D.t26 29.1353
R11593 DFF_magic_0.D.t30 DFF_magic_0.D.t31 29.1353
R11594 DFF_magic_0.D.t34 DFF_magic_0.D.t33 29.1353
R11595 DFF_magic_0.D.t13 DFF_magic_0.D.t12 29.1353
R11596 DFF_magic_0.D.t18 DFF_magic_0.D.t19 29.1353
R11597 DFF_magic_0.D.t21 DFF_magic_0.D.t20 29.1353
R11598 DFF_magic_0.D.t23 DFF_magic_0.D.t22 29.1353
R11599 DFF_magic_0.D.n7 DFF_magic_0.D 28.4293
R11600 DFF_magic_0.D.n14 DFF_magic_0.D.t38 13.5376
R11601 DFF_magic_0.D.n10 DFF_magic_0.D.t28 13.5376
R11602 DFF_magic_0.D.n6 DFF_magic_0.D.t36 13.5376
R11603 DFF_magic_0.D.n7 DFF_magic_0.D.n6 13.1086
R11604 DFF_magic_0.D.n11 DFF_magic_0.D.n10 13.0416
R11605 DFF_magic_0.D.n14 DFF_magic_0.D.t27 12.5549
R11606 DFF_magic_0.D.n10 DFF_magic_0.D.t13 12.5549
R11607 DFF_magic_0.D.n6 DFF_magic_0.D.t23 12.5549
R11608 DFF_magic_0.D.n15 DFF_magic_0.D.n14 12.5041
R11609 DFF_magic_0.D.n12 DFF_magic_0.D.t37 7.3005
R11610 DFF_magic_0.D.n13 DFF_magic_0.D.t24 7.3005
R11611 DFF_magic_0.D.n8 DFF_magic_0.D.t17 7.3005
R11612 DFF_magic_0.D.n9 DFF_magic_0.D.t33 7.3005
R11613 DFF_magic_0.D.n4 DFF_magic_0.D.t35 7.3005
R11614 DFF_magic_0.D.n5 DFF_magic_0.D.t20 7.3005
R11615 DFF_magic_0.D DFF_magic_0.D.n15 5.8063
R11616 DFF_magic_0.D.n1 DFF_magic_0.D.t0 5.68115
R11617 DFF_magic_0.D DFF_magic_0.D.t5 4.928
R11618 DFF_magic_0.D DFF_magic_0.D.n17 3.6455
R11619 DFF_magic_0.D DFF_magic_0.D.n18 3.31072
R11620 DFF_magic_0.D DFF_magic_0.D.n16 3.31072
R11621 DFF_magic_0.D.n3 DFF_magic_0.D.n2 3.1505
R11622 DFF_magic_0.D.n1 DFF_magic_0.D.n0 2.6005
R11623 DFF_magic_0.D.n15 DFF_magic_0.D.n11 2.54426
R11624 DFF_magic_0.D.n11 DFF_magic_0.D.n7 2.36537
R11625 DFF_magic_0.D.n0 DFF_magic_0.D.t1 1.6255
R11626 DFF_magic_0.D.n0 DFF_magic_0.D.t2 1.6255
R11627 DFF_magic_0.D.n16 DFF_magic_0.D.t8 1.6255
R11628 DFF_magic_0.D.n16 DFF_magic_0.D.t7 1.6255
R11629 DFF_magic_0.D.n18 DFF_magic_0.D.t9 1.6255
R11630 DFF_magic_0.D.n18 DFF_magic_0.D.t6 1.6255
R11631 DFF_magic_0.D.n2 DFF_magic_0.D.t3 1.463
R11632 DFF_magic_0.D.n2 DFF_magic_0.D.t4 1.463
R11633 DFF_magic_0.D.n17 DFF_magic_0.D.t10 1.463
R11634 DFF_magic_0.D.n17 DFF_magic_0.D.t11 1.463
R11635 DFF_magic_0.D DFF_magic_0.D.n3 1.45209
R11636 DFF_magic_0.D.n3 DFF_magic_0.D.n1 0.898543
R11637 Q1.t5 Q1.t23 47.8944
R11638 Q1.t24 Q1.t15 47.8944
R11639 Q1.t6 Q1.t28 47.5387
R11640 Q1.t25 Q1.t19 47.5387
R11641 Q1.n20 Q1.n6 46.1005
R11642 Q1.n5 Q1.t16 38.8649
R11643 Q1.n14 Q1.t29 38.7949
R11644 Q1.n13 Q1.t30 38.7949
R11645 Q1.n9 Q1.t17 38.7949
R11646 Q1.n8 Q1.t20 38.7949
R11647 Q1.t27 Q1.t7 31.5469
R11648 Q1.t11 Q1.t27 31.5469
R11649 Q1.t4 Q1.t11 31.5469
R11650 Q1.t18 Q1.t4 31.5469
R11651 Q1.n14 Q1.n13 31.4949
R11652 Q1.n9 Q1.n8 31.4949
R11653 Q1.n4 Q1.t26 28.8568
R11654 Q1.t7 Q1.t9 26.9844
R11655 Q1.n20 Q1.n19 24.0695
R11656 Q1.n12 Q1.n11 18.9058
R11657 Q1.n15 Q1.t22 17.9416
R11658 Q1.n10 Q1.t12 17.9416
R11659 Q1.t16 Q1.n4 17.0773
R11660 Q1.n16 Q1.t6 15.7085
R11661 Q1.n7 Q1.t25 15.7085
R11662 Q1.n3 Q1.t18 15.3175
R11663 Q1.n3 Q1.t21 13.4925
R11664 Q1.n16 Q1.t10 13.4273
R11665 Q1.n7 Q1.t31 13.4273
R11666 Q1.n15 Q1.t5 11.957
R11667 Q1.n10 Q1.t24 11.957
R11668 Q1.n4 Q1.t8 11.6023
R11669 Q1 Q1.n15 9.94647
R11670 Q1 Q1.n10 9.94647
R11671 Q1 Q1.n5 9.27587
R11672 Q1.n19 Q1.n18 9.00923
R11673 Q1.n17 Q1.n12 9.00165
R11674 Q1 Q1.n3 8.10124
R11675 Q1 Q1.n16 8.08021
R11676 Q1 Q1.n7 8.08021
R11677 Q1.n5 Q1.t13 7.3005
R11678 Q1.n13 Q1.t14 7.3005
R11679 Q1.t22 Q1.n14 7.3005
R11680 Q1.n8 Q1.t3 7.3005
R11681 Q1.t12 Q1.n9 7.3005
R11682 Q1.n21 Q1.n20 5.71336
R11683 Q1.n0 Q1.t2 5.47387
R11684 Q1.n1 Q1.t1 4.65398
R11685 Q1.n0 Q1.t0 4.2255
R11686 Q1.n17 Q1 2.46385
R11687 Q1.n11 Q1 2.46321
R11688 Q1 Q1.n21 0.8075
R11689 Q1.n11 Q1 0.58743
R11690 Q1.n21 Q1 0.454173
R11691 Q1.n1 Q1.n0 0.427022
R11692 Q1.n18 Q1 0.259591
R11693 Q1 Q1.n1 0.257096
R11694 Q1.n19 Q1.n12 0.232459
R11695 Q1.n18 Q1.n17 0.229763
R11696 Q1.n6 Q1 0.18935
R11697 Q1.n2 Q1 0.186245
R11698 Q1 Q1.n2 0.0995
R11699 Q1.n2 Q1 0.0139043
R11700 Q1.n6 Q1 0.00166883
R11701 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t6 130.41
R11702 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n5 36.752
R11703 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t7 35.3186
R11704 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t5 33.5023
R11705 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t12 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n0 33.5023
R11706 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t11 32.2349
R11707 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n2 27.7405
R11708 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t9 26.3857
R11709 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t12 16.3786
R11710 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t9 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n3 13.2317
R11711 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n1 12.5032
R11712 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t8 11.3259
R11713 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t10 11.146
R11714 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t3 7.3005
R11715 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t4 7.3005
R11716 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n4 5.87653
R11717 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t2 5.47387
R11718 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t1 5.28011
R11719 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t0 4.65398
R11720 p3_gen_magic_0.P3.t15 p3_gen_magic_0.P3.t11 47.8944
R11721 p3_gen_magic_0.P3.t16 p3_gen_magic_0.P3.t12 44.6331
R11722 p3_gen_magic_0.P3.t7 p3_gen_magic_0.P3.t16 43.4094
R11723 p3_gen_magic_0.P3.n1 p3_gen_magic_0.P3.t10 38.7949
R11724 p3_gen_magic_0.P3.n2 p3_gen_magic_0.P3.t8 38.7949
R11725 p3_gen_magic_0.P3.t13 p3_gen_magic_0.P3.t7 31.5469
R11726 p3_gen_magic_0.P3.n2 p3_gen_magic_0.P3.n1 31.4949
R11727 p3_gen_magic_0.P3.n3 p3_gen_magic_0.P3.t14 17.9416
R11728 p3_gen_magic_0.P3.n4 p3_gen_magic_0.P3.t13 15.0567
R11729 p3_gen_magic_0.P3.n4 p3_gen_magic_0.P3.t6 13.6228
R11730 p3_gen_magic_0.P3.n3 p3_gen_magic_0.P3.t15 11.957
R11731 p3_gen_magic_0.P3 p3_gen_magic_0.P3.n3 9.95929
R11732 p3_gen_magic_0.P3 p3_gen_magic_0.P3.n4 8.2675
R11733 p3_gen_magic_0.P3.n1 p3_gen_magic_0.P3.t9 7.3005
R11734 p3_gen_magic_0.P3.t14 p3_gen_magic_0.P3.n2 7.3005
R11735 p3_gen_magic_0.P3.n0 p3_gen_magic_0.P3.n5 3.6455
R11736 p3_gen_magic_0.P3.n0 p3_gen_magic_0.P3.n6 3.31072
R11737 p3_gen_magic_0.P3.n0 p3_gen_magic_0.P3.n7 2.90572
R11738 p3_gen_magic_0.P3.n6 p3_gen_magic_0.P3.t1 1.6255
R11739 p3_gen_magic_0.P3.n6 p3_gen_magic_0.P3.t0 1.6255
R11740 p3_gen_magic_0.P3.n7 p3_gen_magic_0.P3.t3 1.6255
R11741 p3_gen_magic_0.P3.n7 p3_gen_magic_0.P3.t2 1.6255
R11742 p3_gen_magic_0.P3.n5 p3_gen_magic_0.P3.t5 1.463
R11743 p3_gen_magic_0.P3.n5 p3_gen_magic_0.P3.t4 1.463
R11744 p3_gen_magic_0.P3.n0 p3_gen_magic_0.P3 1.34878
R11745 7b_counter_0.MDFF_4.LD.t28 7b_counter_0.MDFF_4.LD.t35 144.929
R11746 7b_counter_0.MDFF_4.LD.t59 7b_counter_0.MDFF_4.LD.t34 144.929
R11747 7b_counter_0.MDFF_4.LD.t60 7b_counter_0.MDFF_4.LD.t16 144.929
R11748 7b_counter_0.MDFF_4.LD.t17 7b_counter_0.MDFF_4.LD.t89 144.929
R11749 7b_counter_0.MDFF_4.LD.t86 7b_counter_0.MDFF_4.LD.t99 144.929
R11750 7b_counter_0.MDFF_4.LD.t63 7b_counter_0.MDFF_4.LD.t75 144.929
R11751 7b_counter_0.MDFF_4.LD.t116 7b_counter_0.MDFF_4.LD.t70 144.929
R11752 7b_counter_0.MDFF_4.LD.t31 7b_counter_0.MDFF_4.LD.t68 144.929
R11753 7b_counter_0.MDFF_4.LD.t67 7b_counter_0.MDFF_4.LD.t111 144.929
R11754 7b_counter_0.MDFF_4.LD.n11 7b_counter_0.MDFF_4.LD.t85 69.1459
R11755 7b_counter_0.MDFF_4.LD.n42 7b_counter_0.MDFF_4.LD.t69 66.03
R11756 7b_counter_0.MDFF_4.LD.n68 7b_counter_0.MDFF_4.LD.t107 32.714
R11757 7b_counter_0.MDFF_4.LD.n31 7b_counter_0.MDFF_4.LD.t92 32.714
R11758 7b_counter_0.MDFF_4.LD.n39 7b_counter_0.MDFF_4.LD.t93 32.714
R11759 7b_counter_0.MDFF_4.LD.n44 7b_counter_0.MDFF_4.LD.t103 32.714
R11760 7b_counter_0.MDFF_4.LD.n55 7b_counter_0.MDFF_4.LD.t119 32.714
R11761 7b_counter_0.MDFF_4.LD.n63 7b_counter_0.MDFF_4.LD.t98 32.714
R11762 7b_counter_0.MDFF_4.LD.n12 7b_counter_0.MDFF_4.LD.t109 32.714
R11763 7b_counter_0.MDFF_4.LD.n20 7b_counter_0.MDFF_4.LD.t24 32.714
R11764 7b_counter_0.MDFF_4.LD.n8 7b_counter_0.MDFF_4.LD.t8 32.714
R11765 7b_counter_0.MDFF_4.LD.n66 7b_counter_0.MDFF_4.LD.t114 27.7917
R11766 7b_counter_0.MDFF_4.LD.n37 7b_counter_0.MDFF_4.LD.t97 25.1498
R11767 7b_counter_0.MDFF_4.LD.n53 7b_counter_0.MDFF_4.LD.t18 25.0633
R11768 7b_counter_0.MDFF_4.LD.n61 7b_counter_0.MDFF_4.LD.t27 25.0633
R11769 7b_counter_0.MDFF_4.LD.n18 7b_counter_0.MDFF_4.LD.t118 25.0633
R11770 7b_counter_0.MDFF_4.LD.n6 7b_counter_0.MDFF_4.LD.t30 25.0633
R11771 7b_counter_0.MDFF_4.LD.n29 7b_counter_0.MDFF_4.LD.t115 24.9839
R11772 7b_counter_0.MDFF_4.LD.n69 7b_counter_0.MDFF_4.LD.n68 21.0471
R11773 7b_counter_0.MDFF_4.LD.n32 7b_counter_0.MDFF_4.LD.n31 21.0471
R11774 7b_counter_0.MDFF_4.LD.n40 7b_counter_0.MDFF_4.LD.n39 21.0471
R11775 7b_counter_0.MDFF_4.LD.n45 7b_counter_0.MDFF_4.LD.n44 21.0471
R11776 7b_counter_0.MDFF_4.LD.n56 7b_counter_0.MDFF_4.LD.n55 21.0471
R11777 7b_counter_0.MDFF_4.LD.n64 7b_counter_0.MDFF_4.LD.n63 21.0471
R11778 7b_counter_0.MDFF_4.LD.n13 7b_counter_0.MDFF_4.LD.n12 21.0471
R11779 7b_counter_0.MDFF_4.LD.n21 7b_counter_0.MDFF_4.LD.n20 21.0471
R11780 7b_counter_0.MDFF_4.LD.n9 7b_counter_0.MDFF_4.LD.n8 21.0471
R11781 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n0 20.2647
R11782 7b_counter_0.MDFF_4.LD.t92 7b_counter_0.MDFF_4.LD 20.2341
R11783 7b_counter_0.MDFF_4.LD.t93 7b_counter_0.MDFF_4.LD 20.2341
R11784 7b_counter_0.MDFF_4.LD.t103 7b_counter_0.MDFF_4.LD 20.2341
R11785 7b_counter_0.MDFF_4.LD.t107 7b_counter_0.MDFF_4.LD 20.2328
R11786 7b_counter_0.MDFF_4.LD.t119 7b_counter_0.MDFF_4.LD 20.2328
R11787 7b_counter_0.MDFF_4.LD.t98 7b_counter_0.MDFF_4.LD 20.2328
R11788 7b_counter_0.MDFF_4.LD.t109 7b_counter_0.MDFF_4.LD 20.2328
R11789 7b_counter_0.MDFF_4.LD.t24 7b_counter_0.MDFF_4.LD 20.2328
R11790 7b_counter_0.MDFF_4.LD.t8 7b_counter_0.MDFF_4.LD 20.2328
R11791 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n11 18.0523
R11792 7b_counter_0.MDFF_4.LD.n71 7b_counter_0.MDFF_4.LD.n70 15.8172
R11793 7b_counter_0.MDFF_4.LD.n72 7b_counter_0.MDFF_4.LD.n71 15.8172
R11794 7b_counter_0.MDFF_4.LD.n27 7b_counter_0.MDFF_4.LD.n26 15.8172
R11795 7b_counter_0.MDFF_4.LD.n28 7b_counter_0.MDFF_4.LD.n27 15.8172
R11796 7b_counter_0.MDFF_4.LD.n35 7b_counter_0.MDFF_4.LD.n34 15.8172
R11797 7b_counter_0.MDFF_4.LD.n36 7b_counter_0.MDFF_4.LD.n35 15.8172
R11798 7b_counter_0.MDFF_4.LD.n47 7b_counter_0.MDFF_4.LD.n46 15.8172
R11799 7b_counter_0.MDFF_4.LD.n48 7b_counter_0.MDFF_4.LD.n47 15.8172
R11800 7b_counter_0.MDFF_4.LD.n51 7b_counter_0.MDFF_4.LD.n50 15.8172
R11801 7b_counter_0.MDFF_4.LD.n52 7b_counter_0.MDFF_4.LD.n51 15.8172
R11802 7b_counter_0.MDFF_4.LD.n59 7b_counter_0.MDFF_4.LD.n58 15.8172
R11803 7b_counter_0.MDFF_4.LD.n60 7b_counter_0.MDFF_4.LD.n59 15.8172
R11804 7b_counter_0.MDFF_4.LD.n15 7b_counter_0.MDFF_4.LD.n14 15.8172
R11805 7b_counter_0.MDFF_4.LD.n16 7b_counter_0.MDFF_4.LD.n15 15.8172
R11806 7b_counter_0.MDFF_4.LD.n23 7b_counter_0.MDFF_4.LD.n22 15.8172
R11807 7b_counter_0.MDFF_4.LD.n24 7b_counter_0.MDFF_4.LD.n23 15.8172
R11808 7b_counter_0.MDFF_4.LD.n4 7b_counter_0.MDFF_4.LD.n3 15.8172
R11809 7b_counter_0.MDFF_4.LD.n5 7b_counter_0.MDFF_4.LD.n4 15.8172
R11810 7b_counter_0.MDFF_4.LD.n67 7b_counter_0.MDFF_4.LD.t28 14.7678
R11811 7b_counter_0.MDFF_4.LD.n43 7b_counter_0.MDFF_4.LD.t17 14.7678
R11812 7b_counter_0.MDFF_4.LD.n19 7b_counter_0.MDFF_4.LD.t31 14.7678
R11813 7b_counter_0.MDFF_4.LD.n30 7b_counter_0.MDFF_4.LD.t59 14.7032
R11814 7b_counter_0.MDFF_4.LD.n38 7b_counter_0.MDFF_4.LD.t60 14.7032
R11815 7b_counter_0.MDFF_4.LD.n54 7b_counter_0.MDFF_4.LD.t86 14.7032
R11816 7b_counter_0.MDFF_4.LD.n62 7b_counter_0.MDFF_4.LD.t63 14.7032
R11817 7b_counter_0.MDFF_4.LD.n7 7b_counter_0.MDFF_4.LD.t67 14.7032
R11818 7b_counter_0.MDFF_4.LD.n73 7b_counter_0.MDFF_4.LD.t36 14.5353
R11819 7b_counter_0.MDFF_4.LD.n33 7b_counter_0.MDFF_4.LD.t61 14.5353
R11820 7b_counter_0.MDFF_4.LD.n41 7b_counter_0.MDFF_4.LD.t62 14.5353
R11821 7b_counter_0.MDFF_4.LD.n49 7b_counter_0.MDFF_4.LD.t82 14.5353
R11822 7b_counter_0.MDFF_4.LD.n57 7b_counter_0.MDFF_4.LD.t12 14.5353
R11823 7b_counter_0.MDFF_4.LD.n65 7b_counter_0.MDFF_4.LD.t11 14.5353
R11824 7b_counter_0.MDFF_4.LD.n17 7b_counter_0.MDFF_4.LD.t44 14.5353
R11825 7b_counter_0.MDFF_4.LD.n25 7b_counter_0.MDFF_4.LD.t43 14.5353
R11826 7b_counter_0.MDFF_4.LD.n10 7b_counter_0.MDFF_4.LD.t19 14.5353
R11827 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n67 13.7626
R11828 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n30 13.7626
R11829 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n38 13.7626
R11830 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n43 13.7626
R11831 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n54 13.7626
R11832 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n62 13.7626
R11833 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n19 13.7626
R11834 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n7 13.7626
R11835 7b_counter_0.MDFF_4.LD.n70 7b_counter_0.MDFF_4.LD.t47 11.7326
R11836 7b_counter_0.MDFF_4.LD.n70 7b_counter_0.MDFF_4.LD.t6 11.7326
R11837 7b_counter_0.MDFF_4.LD.n71 7b_counter_0.MDFF_4.LD.t76 11.7326
R11838 7b_counter_0.MDFF_4.LD.n71 7b_counter_0.MDFF_4.LD.t120 11.7326
R11839 7b_counter_0.MDFF_4.LD.n72 7b_counter_0.MDFF_4.LD.t33 11.7326
R11840 7b_counter_0.MDFF_4.LD.t36 7b_counter_0.MDFF_4.LD.n72 11.7326
R11841 7b_counter_0.MDFF_4.LD.n26 7b_counter_0.MDFF_4.LD.t41 11.7326
R11842 7b_counter_0.MDFF_4.LD.n26 7b_counter_0.MDFF_4.LD.t13 11.7326
R11843 7b_counter_0.MDFF_4.LD.n27 7b_counter_0.MDFF_4.LD.t80 11.7326
R11844 7b_counter_0.MDFF_4.LD.n27 7b_counter_0.MDFF_4.LD.t58 11.7326
R11845 7b_counter_0.MDFF_4.LD.n28 7b_counter_0.MDFF_4.LD.t83 11.7326
R11846 7b_counter_0.MDFF_4.LD.t61 7b_counter_0.MDFF_4.LD.n28 11.7326
R11847 7b_counter_0.MDFF_4.LD.n34 7b_counter_0.MDFF_4.LD.t42 11.7326
R11848 7b_counter_0.MDFF_4.LD.n34 7b_counter_0.MDFF_4.LD.t14 11.7326
R11849 7b_counter_0.MDFF_4.LD.n35 7b_counter_0.MDFF_4.LD.t52 11.7326
R11850 7b_counter_0.MDFF_4.LD.n35 7b_counter_0.MDFF_4.LD.t26 11.7326
R11851 7b_counter_0.MDFF_4.LD.n36 7b_counter_0.MDFF_4.LD.t84 11.7326
R11852 7b_counter_0.MDFF_4.LD.t62 7b_counter_0.MDFF_4.LD.n36 11.7326
R11853 7b_counter_0.MDFF_4.LD.n46 7b_counter_0.MDFF_4.LD.t37 11.7326
R11854 7b_counter_0.MDFF_4.LD.n46 7b_counter_0.MDFF_4.LD.t73 11.7326
R11855 7b_counter_0.MDFF_4.LD.n47 7b_counter_0.MDFF_4.LD.t50 11.7326
R11856 7b_counter_0.MDFF_4.LD.n47 7b_counter_0.MDFF_4.LD.t56 11.7326
R11857 7b_counter_0.MDFF_4.LD.n48 7b_counter_0.MDFF_4.LD.t29 11.7326
R11858 7b_counter_0.MDFF_4.LD.t82 7b_counter_0.MDFF_4.LD.n48 11.7326
R11859 7b_counter_0.MDFF_4.LD.n50 7b_counter_0.MDFF_4.LD.t65 11.7326
R11860 7b_counter_0.MDFF_4.LD.n50 7b_counter_0.MDFF_4.LD.t38 11.7326
R11861 7b_counter_0.MDFF_4.LD.n51 7b_counter_0.MDFF_4.LD.t51 11.7326
R11862 7b_counter_0.MDFF_4.LD.n51 7b_counter_0.MDFF_4.LD.t25 11.7326
R11863 7b_counter_0.MDFF_4.LD.n52 7b_counter_0.MDFF_4.LD.t40 11.7326
R11864 7b_counter_0.MDFF_4.LD.t12 7b_counter_0.MDFF_4.LD.n52 11.7326
R11865 7b_counter_0.MDFF_4.LD.n58 7b_counter_0.MDFF_4.LD.t48 11.7326
R11866 7b_counter_0.MDFF_4.LD.n58 7b_counter_0.MDFF_4.LD.t20 11.7326
R11867 7b_counter_0.MDFF_4.LD.n59 7b_counter_0.MDFF_4.LD.t78 11.7326
R11868 7b_counter_0.MDFF_4.LD.n59 7b_counter_0.MDFF_4.LD.t55 11.7326
R11869 7b_counter_0.MDFF_4.LD.n60 7b_counter_0.MDFF_4.LD.t39 11.7326
R11870 7b_counter_0.MDFF_4.LD.t11 7b_counter_0.MDFF_4.LD.n60 11.7326
R11871 7b_counter_0.MDFF_4.LD.n14 7b_counter_0.MDFF_4.LD.t49 11.7326
R11872 7b_counter_0.MDFF_4.LD.n14 7b_counter_0.MDFF_4.LD.t87 11.7326
R11873 7b_counter_0.MDFF_4.LD.n15 7b_counter_0.MDFF_4.LD.t54 11.7326
R11874 7b_counter_0.MDFF_4.LD.n15 7b_counter_0.MDFF_4.LD.t112 11.7326
R11875 7b_counter_0.MDFF_4.LD.n16 7b_counter_0.MDFF_4.LD.t15 11.7326
R11876 7b_counter_0.MDFF_4.LD.t44 7b_counter_0.MDFF_4.LD.n16 11.7326
R11877 7b_counter_0.MDFF_4.LD.n22 7b_counter_0.MDFF_4.LD.t77 11.7326
R11878 7b_counter_0.MDFF_4.LD.n22 7b_counter_0.MDFF_4.LD.t66 11.7326
R11879 7b_counter_0.MDFF_4.LD.n23 7b_counter_0.MDFF_4.LD.t71 11.7326
R11880 7b_counter_0.MDFF_4.LD.n23 7b_counter_0.MDFF_4.LD.t88 11.7326
R11881 7b_counter_0.MDFF_4.LD.n24 7b_counter_0.MDFF_4.LD.t117 11.7326
R11882 7b_counter_0.MDFF_4.LD.t43 7b_counter_0.MDFF_4.LD.n24 11.7326
R11883 7b_counter_0.MDFF_4.LD.n3 7b_counter_0.MDFF_4.LD.t79 11.7326
R11884 7b_counter_0.MDFF_4.LD.n3 7b_counter_0.MDFF_4.LD.t57 11.7326
R11885 7b_counter_0.MDFF_4.LD.n4 7b_counter_0.MDFF_4.LD.t72 11.7326
R11886 7b_counter_0.MDFF_4.LD.n4 7b_counter_0.MDFF_4.LD.t45 11.7326
R11887 7b_counter_0.MDFF_4.LD.n5 7b_counter_0.MDFF_4.LD.t46 11.7326
R11888 7b_counter_0.MDFF_4.LD.t19 7b_counter_0.MDFF_4.LD.n5 11.7326
R11889 7b_counter_0.MDFF_4.LD.n69 7b_counter_0.MDFF_4.LD.t101 11.6675
R11890 7b_counter_0.MDFF_4.LD.n32 7b_counter_0.MDFF_4.LD.t21 11.6675
R11891 7b_counter_0.MDFF_4.LD.n40 7b_counter_0.MDFF_4.LD.t23 11.6675
R11892 7b_counter_0.MDFF_4.LD.n45 7b_counter_0.MDFF_4.LD.t32 11.6675
R11893 7b_counter_0.MDFF_4.LD.n56 7b_counter_0.MDFF_4.LD.t91 11.6675
R11894 7b_counter_0.MDFF_4.LD.n64 7b_counter_0.MDFF_4.LD.t90 11.6675
R11895 7b_counter_0.MDFF_4.LD.n13 7b_counter_0.MDFF_4.LD.t106 11.6675
R11896 7b_counter_0.MDFF_4.LD.n21 7b_counter_0.MDFF_4.LD.t105 11.6675
R11897 7b_counter_0.MDFF_4.LD.n9 7b_counter_0.MDFF_4.LD.t96 11.6675
R11898 7b_counter_0.MDFF_4.LD.n11 7b_counter_0.MDFF_4.LD.t116 11.6023
R11899 7b_counter_0.MDFF_4.LD.n29 7b_counter_0.MDFF_4.LD.t94 11.4552
R11900 7b_counter_0.MDFF_4.LD.n37 7b_counter_0.MDFF_4.LD.t95 11.4552
R11901 7b_counter_0.MDFF_4.LD.n53 7b_counter_0.MDFF_4.LD.t122 11.4552
R11902 7b_counter_0.MDFF_4.LD.n61 7b_counter_0.MDFF_4.LD.t104 11.4552
R11903 7b_counter_0.MDFF_4.LD.n6 7b_counter_0.MDFF_4.LD.t108 11.4552
R11904 7b_counter_0.MDFF_4.LD.n66 7b_counter_0.MDFF_4.LD.t74 11.3906
R11905 7b_counter_0.MDFF_4.LD.n18 7b_counter_0.MDFF_4.LD.t81 11.3906
R11906 7b_counter_0.MDFF_4.LD.n42 7b_counter_0.MDFF_4.LD.t64 11.3901
R11907 7b_counter_0.MDFF_4.LD.n1 7b_counter_0.MDFF_4.LD.n0 4.43798
R11908 7b_counter_0.MDFF_4.LD.n1 7b_counter_0.MDFF_4.LD.n2 0.792707
R11909 7b_counter_0.MDFF_4.LD.n11 7b_counter_0.MDFF_4.LD.t53 9.58175
R11910 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n73 8.19616
R11911 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n33 8.19616
R11912 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n41 8.19616
R11913 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n49 8.19616
R11914 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n57 8.19616
R11915 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n65 8.19616
R11916 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n17 8.19616
R11917 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n25 8.19616
R11918 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.LD.n10 8.19616
R11919 7b_counter_0.MDFF_4.LD.n68 7b_counter_0.MDFF_4.LD.t22 7.3005
R11920 7b_counter_0.MDFF_4.LD.n31 7b_counter_0.MDFF_4.LD.t9 7.3005
R11921 7b_counter_0.MDFF_4.LD.n39 7b_counter_0.MDFF_4.LD.t102 7.3005
R11922 7b_counter_0.MDFF_4.LD.n44 7b_counter_0.MDFF_4.LD.t110 7.3005
R11923 7b_counter_0.MDFF_4.LD.n55 7b_counter_0.MDFF_4.LD.t100 7.3005
R11924 7b_counter_0.MDFF_4.LD.n63 7b_counter_0.MDFF_4.LD.t7 7.3005
R11925 7b_counter_0.MDFF_4.LD.n12 7b_counter_0.MDFF_4.LD.t113 7.3005
R11926 7b_counter_0.MDFF_4.LD.n20 7b_counter_0.MDFF_4.LD.t10 7.3005
R11927 7b_counter_0.MDFF_4.LD.n8 7b_counter_0.MDFF_4.LD.t121 7.3005
R11928 7b_counter_0.MDFF_4.LD.n0 7b_counter_0.MDFF_4.LD.t2 5.86349
R11929 7b_counter_0.MDFF_4.LD.n2 7b_counter_0.MDFF_4.LD.t3 4.63638
R11930 7b_counter_0.MDFF_4.LD.n0 7b_counter_0.MDFF_4.LD.t1 4.63638
R11931 7b_counter_0.MDFF_4.LD.n2 7b_counter_0.MDFF_4.LD.t4 4.2255
R11932 7b_counter_0.MDFF_4.LD.n0 7b_counter_0.MDFF_4.LD.t5 4.2255
R11933 7b_counter_0.MDFF_4.LD.n73 7b_counter_0.MDFF_4.LD.n69 2.47729
R11934 7b_counter_0.MDFF_4.LD.n33 7b_counter_0.MDFF_4.LD.n32 2.47729
R11935 7b_counter_0.MDFF_4.LD.n41 7b_counter_0.MDFF_4.LD.n40 2.47729
R11936 7b_counter_0.MDFF_4.LD.n49 7b_counter_0.MDFF_4.LD.n45 2.47729
R11937 7b_counter_0.MDFF_4.LD.n57 7b_counter_0.MDFF_4.LD.n56 2.47729
R11938 7b_counter_0.MDFF_4.LD.n65 7b_counter_0.MDFF_4.LD.n64 2.47729
R11939 7b_counter_0.MDFF_4.LD.n17 7b_counter_0.MDFF_4.LD.n13 2.47729
R11940 7b_counter_0.MDFF_4.LD.n25 7b_counter_0.MDFF_4.LD.n21 2.47729
R11941 7b_counter_0.MDFF_4.LD.n10 7b_counter_0.MDFF_4.LD.n9 2.47729
R11942 7b_counter_0.MDFF_4.LD.n67 7b_counter_0.MDFF_4.LD.n66 2.45537
R11943 7b_counter_0.MDFF_4.LD.n30 7b_counter_0.MDFF_4.LD.n29 2.45537
R11944 7b_counter_0.MDFF_4.LD.n38 7b_counter_0.MDFF_4.LD.n37 2.45537
R11945 7b_counter_0.MDFF_4.LD.n54 7b_counter_0.MDFF_4.LD.n53 2.45537
R11946 7b_counter_0.MDFF_4.LD.n62 7b_counter_0.MDFF_4.LD.n61 2.45537
R11947 7b_counter_0.MDFF_4.LD.n19 7b_counter_0.MDFF_4.LD.n18 2.45537
R11948 7b_counter_0.MDFF_4.LD.n7 7b_counter_0.MDFF_4.LD.n6 2.45537
R11949 7b_counter_0.MDFF_4.LD.n43 7b_counter_0.MDFF_4.LD.n42 2.42339
R11950 7b_counter_0.MDFF_4.LD.n1 7b_counter_0.MDFF_4.LD.t0 5.02188
R11951 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t3 130.41
R11952 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n5 36.752
R11953 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t8 35.3186
R11954 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t5 33.5023
R11955 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t12 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n0 33.5023
R11956 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t4 32.2349
R11957 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n2 27.7405
R11958 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t11 26.3857
R11959 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t12 16.3786
R11960 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t11 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n3 13.2317
R11961 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n1 12.5032
R11962 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t7 11.3259
R11963 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t6 11.146
R11964 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t9 7.3005
R11965 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t10 7.3005
R11966 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n4 5.87653
R11967 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t2 5.47387
R11968 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t0 5.28011
R11969 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t1 4.65398
R11970 p3_gen_magic_0.3_inp_AND_magic_0.C.n1 p3_gen_magic_0.3_inp_AND_magic_0.C.t2 39.1562
R11971 p3_gen_magic_0.3_inp_AND_magic_0.C.t4 p3_gen_magic_0.3_inp_AND_magic_0.C.t1 28.8746
R11972 p3_gen_magic_0.3_inp_AND_magic_0.C.t2 p3_gen_magic_0.3_inp_AND_magic_0.C.t3 23.4648
R11973 p3_gen_magic_0.3_inp_AND_magic_0.C.n0 p3_gen_magic_0.3_inp_AND_magic_0.C.t5 14.1443
R11974 p3_gen_magic_0.3_inp_AND_magic_0.C.n0 p3_gen_magic_0.3_inp_AND_magic_0.C.t4 13.8835
R11975 p3_gen_magic_0.3_inp_AND_magic_0.C.n1 p3_gen_magic_0.3_inp_AND_magic_0.C.n0 12.5017
R11976 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.3_inp_AND_magic_0.C.n1 5.35629
R11977 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.3_inp_AND_magic_0.C.t0 3.46108
R11978 D2_5.t5 D2_5.t23 47.8944
R11979 D2_5.t10 D2_5.t6 47.8944
R11980 D2_5.t16 D2_5.t13 47.5387
R11981 D2_5.t2 D2_5.t20 47.5387
R11982 D2_5.n3 D2_5.t14 38.8649
R11983 D2_5.n1 D2_5.t15 38.8649
R11984 D2_5.n5 D2_5.t22 38.7949
R11985 D2_5.n4 D2_5.t1 38.7949
R11986 D2_5.n10 D2_5.t7 38.7949
R11987 D2_5.n9 D2_5.t9 38.7949
R11988 D2_5.n5 D2_5.n4 31.4949
R11989 D2_5.n10 D2_5.n9 31.4949
R11990 D2_5.n2 D2_5.t25 28.8568
R11991 D2_5.n0 D2_5.t24 28.8568
R11992 D2_5.n14 D2_5.n8 18.892
R11993 D2_5.n14 D2_5.n13 18.602
R11994 D2_5.n6 D2_5.t12 17.9416
R11995 D2_5.n11 D2_5.t19 17.9416
R11996 D2_5.t14 D2_5.n2 17.0773
R11997 D2_5.t15 D2_5.n0 17.0773
R11998 D2_5.n7 D2_5.t16 16.621
R11999 D2_5.n12 D2_5.t2 16.621
R12000 D2_5.n15 D2_5.n14 15.3785
R12001 D2_5.n7 D2_5.t11 12.5148
R12002 D2_5.n12 D2_5.t18 12.5148
R12003 D2_5.n6 D2_5.t5 11.957
R12004 D2_5.n11 D2_5.t10 11.957
R12005 D2_5.n2 D2_5.t4 11.6023
R12006 D2_5.n0 D2_5.t3 11.6023
R12007 D2_5 D2_5.n6 9.95286
R12008 D2_5 D2_5.n11 9.95286
R12009 D2_5 D2_5.n3 9.27587
R12010 D2_5 D2_5.n1 9.27587
R12011 D2_5 D2_5.n7 8.59246
R12012 D2_5 D2_5.n12 8.59246
R12013 D2_5.n16 D2_5.n15 8.11394
R12014 D2_5.n15 D2_5 7.97404
R12015 D2_5.n4 D2_5.t8 7.3005
R12016 D2_5.t12 D2_5.n5 7.3005
R12017 D2_5.n9 D2_5.t17 7.3005
R12018 D2_5.t19 D2_5.n10 7.3005
R12019 D2_5.n3 D2_5.t21 7.3005
R12020 D2_5.n1 D2_5.t0 7.3005
R12021 D2_5.n8 D2_5 1.4268
R12022 D2_5.n13 D2_5 1.35441
R12023 D2_5.n13 D2_5 0.190361
R12024 D2_5.n8 D2_5 0.11797
R12025 D2_5.n16 D2_5 0.0740494
R12026 D2_5 D2_5.n16 0.0339615
R12027 divide_by_2_1.tg_magic_3.CLK.t2 divide_by_2_1.tg_magic_3.CLK.t11 47.8944
R12028 divide_by_2_1.tg_magic_3.CLK.t1 divide_by_2_1.tg_magic_3.CLK.t0 47.8944
R12029 divide_by_2_1.inverter_magic_5.VOUT divide_by_2_1.tg_magic_3.CLK.t6 47.3388
R12030 divide_by_2_1.tg_magic_2.CLK divide_by_2_1.tg_magic_3.CLK.t4 47.2524
R12031 divide_by_2_1.tg_magic_3.CLK.n5 divide_by_2_1.tg_magic_3.CLK.t17 38.7949
R12032 divide_by_2_1.tg_magic_3.CLK.n6 divide_by_2_1.tg_magic_3.CLK.t15 38.7949
R12033 divide_by_2_1.tg_magic_3.CLK.n2 divide_by_2_1.tg_magic_3.CLK.t13 38.7949
R12034 divide_by_2_1.tg_magic_3.CLK.n1 divide_by_2_1.tg_magic_3.CLK.t8 38.7949
R12035 divide_by_2_1.tg_magic_3.CLK.n6 divide_by_2_1.tg_magic_3.CLK.n5 31.4949
R12036 divide_by_2_1.tg_magic_3.CLK.n2 divide_by_2_1.tg_magic_3.CLK.n1 31.4949
R12037 divide_by_2_1.tg_magic_3.CLK.n4 divide_by_2_1.tg_magic_3.CLK.t9 26.9781
R12038 divide_by_2_1.tg_magic_3.CLK.n4 divide_by_2_1.tg_magic_3.CLK.t16 26.9781
R12039 divide_by_2_1.tg_magic_3.CLK.n0 divide_by_2_1.tg_magic_3.CLK.t7 26.9781
R12040 divide_by_2_1.tg_magic_3.CLK.n0 divide_by_2_1.tg_magic_3.CLK.t5 26.9781
R12041 divide_by_2_1.inverter_magic_5.VOUT divide_by_2_1.tg_magic_2.CLK 20.617
R12042 divide_by_2_1.tg_magic_3.CLK.n7 divide_by_2_1.tg_magic_3.CLK.t10 17.9416
R12043 divide_by_2_1.tg_magic_3.CLK.n3 divide_by_2_1.tg_magic_3.CLK.t14 17.9416
R12044 divide_by_2_1.tg_magic_3.CLK.n7 divide_by_2_1.tg_magic_3.CLK.t2 11.957
R12045 divide_by_2_1.tg_magic_3.CLK.n3 divide_by_2_1.tg_magic_3.CLK.t1 11.957
R12046 divide_by_2_1.inverter_magic_5.VOUT divide_by_2_1.tg_magic_3.CLK.n3 10.8079
R12047 divide_by_2_1.tg_magic_2.CLK divide_by_2_1.tg_magic_3.CLK.n7 10.0908
R12048 divide_by_2_1.tg_magic_3.CLK.n5 divide_by_2_1.tg_magic_3.CLK.t3 7.3005
R12049 divide_by_2_1.tg_magic_3.CLK.t10 divide_by_2_1.tg_magic_3.CLK.n6 7.3005
R12050 divide_by_2_1.tg_magic_3.CLK.t4 divide_by_2_1.tg_magic_3.CLK.n4 7.3005
R12051 divide_by_2_1.tg_magic_3.CLK.n1 divide_by_2_1.tg_magic_3.CLK.t12 7.3005
R12052 divide_by_2_1.tg_magic_3.CLK.t14 divide_by_2_1.tg_magic_3.CLK.n2 7.3005
R12053 divide_by_2_1.tg_magic_3.CLK.t6 divide_by_2_1.tg_magic_3.CLK.n0 7.3005
R12054 Q6.n6 Q6 52.5285
R12055 Q6.t15 Q6.t4 48.3065
R12056 Q6.t5 Q6.t29 47.8944
R12057 Q6.t24 Q6.t19 47.8944
R12058 Q6.t7 Q6.t21 47.5387
R12059 Q6.t27 Q6.t13 47.5387
R12060 Q6.n4 Q6.t12 38.8649
R12061 Q6.n13 Q6.t6 38.7949
R12062 Q6.n12 Q6.t10 38.7949
R12063 Q6.n8 Q6.t23 38.7949
R12064 Q6.n7 Q6.t26 38.7949
R12065 Q6.t4 Q6.t25 31.5469
R12066 Q6.t11 Q6.t15 31.5469
R12067 Q6.n13 Q6.n12 31.4949
R12068 Q6.n8 Q6.n7 31.4949
R12069 Q6.n3 Q6.t20 28.8568
R12070 Q6.n6 Q6.n5 28.2186
R12071 Q6 Q6.n2 24.7556
R12072 Q6 Q6.n17 19.4925
R12073 Q6.n17 Q6.n11 18.3057
R12074 Q6.n2 Q6.t11 18.2505
R12075 Q6.n14 Q6.t16 17.9416
R12076 Q6.n9 Q6.t9 17.9416
R12077 Q6.t12 Q6.n3 17.0773
R12078 Q6.n15 Q6.t7 15.7085
R12079 Q6.n10 Q6.t27 15.7085
R12080 Q6.n15 Q6.t28 13.4273
R12081 Q6.n10 Q6.t17 13.4273
R12082 Q6.n14 Q6.t5 11.957
R12083 Q6.n9 Q6.t24 11.957
R12084 Q6.n3 Q6.t22 11.6023
R12085 Q6.n2 Q6.t8 11.4067
R12086 Q6 Q6.n14 9.94647
R12087 Q6 Q6.n9 9.94647
R12088 Q6 Q6.n4 9.27587
R12089 Q6 Q6.n15 8.08021
R12090 Q6 Q6.n10 8.08021
R12091 Q6.n4 Q6.t18 7.3005
R12092 Q6.n12 Q6.t14 7.3005
R12093 Q6.t16 Q6.n13 7.3005
R12094 Q6.n7 Q6.t3 7.3005
R12095 Q6.t9 Q6.n8 7.3005
R12096 Q6.n0 Q6.t2 5.47387
R12097 Q6.n17 Q6.n16 4.95531
R12098 Q6.n1 Q6.t1 4.65398
R12099 Q6.n0 Q6.t0 4.2255
R12100 Q6.n11 Q6 2.41882
R12101 Q6.n16 Q6 1.96503
R12102 Q6 Q6.n6 1.88133
R12103 Q6.n16 Q6 1.15959
R12104 Q6.n11 Q6 0.651998
R12105 Q6.n1 Q6.n0 0.427022
R12106 Q6 Q6.n1 0.257096
R12107 Q6.n5 Q6 0.010625
R12108 Q6.n5 Q6 0.0095
R12109 divide_by_2_0.tg_magic_3.CLK.t10 divide_by_2_0.tg_magic_3.CLK.t16 47.8944
R12110 divide_by_2_0.tg_magic_3.CLK.t6 divide_by_2_0.tg_magic_3.CLK.t19 47.8944
R12111 divide_by_2_0.tg_magic_3.CLK.t1 divide_by_2_0.tg_magic_3.CLK.t9 47.3388
R12112 divide_by_2_0.tg_magic_2.CLK divide_by_2_0.tg_magic_3.CLK.t4 47.2524
R12113 divide_by_2_0.tg_magic_3.CLK.n5 divide_by_2_0.tg_magic_3.CLK.t14 38.7949
R12114 divide_by_2_0.tg_magic_3.CLK.n6 divide_by_2_0.tg_magic_3.CLK.t2 38.7949
R12115 divide_by_2_0.tg_magic_3.CLK.n2 divide_by_2_0.tg_magic_3.CLK.t3 38.7949
R12116 divide_by_2_0.tg_magic_3.CLK.n1 divide_by_2_0.tg_magic_3.CLK.t15 38.7949
R12117 divide_by_2_0.tg_magic_3.CLK.n6 divide_by_2_0.tg_magic_3.CLK.n5 31.4949
R12118 divide_by_2_0.tg_magic_3.CLK.n2 divide_by_2_0.tg_magic_3.CLK.n1 31.4949
R12119 divide_by_2_0.tg_magic_3.CLK.n4 divide_by_2_0.tg_magic_3.CLK.t7 26.9781
R12120 divide_by_2_0.tg_magic_3.CLK.n4 divide_by_2_0.tg_magic_3.CLK.t18 26.9781
R12121 divide_by_2_0.tg_magic_3.CLK.n0 divide_by_2_0.tg_magic_3.CLK.t12 26.9781
R12122 divide_by_2_0.tg_magic_3.CLK.n0 divide_by_2_0.tg_magic_3.CLK.t17 26.9781
R12123 divide_by_2_0.tg_magic_3.CLK.t1 divide_by_2_0.tg_magic_2.CLK 20.617
R12124 divide_by_2_0.tg_magic_3.CLK.n7 divide_by_2_0.tg_magic_3.CLK.t5 17.9416
R12125 divide_by_2_0.tg_magic_3.CLK.n3 divide_by_2_0.tg_magic_3.CLK.t11 17.9416
R12126 divide_by_2_0.tg_magic_3.CLK.n7 divide_by_2_0.tg_magic_3.CLK.t10 11.957
R12127 divide_by_2_0.tg_magic_3.CLK.n3 divide_by_2_0.tg_magic_3.CLK.t6 11.957
R12128 divide_by_2_0.tg_magic_2.CLK divide_by_2_0.tg_magic_3.CLK.n7 10.0908
R12129 divide_by_2_0.tg_magic_3.CLK.t1 divide_by_2_0.tg_magic_3.CLK.n3 9.77618
R12130 divide_by_2_0.tg_magic_3.CLK.n5 divide_by_2_0.tg_magic_3.CLK.t13 7.3005
R12131 divide_by_2_0.tg_magic_3.CLK.t5 divide_by_2_0.tg_magic_3.CLK.n6 7.3005
R12132 divide_by_2_0.tg_magic_3.CLK.t4 divide_by_2_0.tg_magic_3.CLK.n4 7.3005
R12133 divide_by_2_0.tg_magic_3.CLK.n1 divide_by_2_0.tg_magic_3.CLK.t8 7.3005
R12134 divide_by_2_0.tg_magic_3.CLK.t11 divide_by_2_0.tg_magic_3.CLK.n2 7.3005
R12135 divide_by_2_0.tg_magic_3.CLK.t9 divide_by_2_0.tg_magic_3.CLK.n0 7.3005
R12136 divide_by_2_0.tg_magic_3.CLK.t1 divide_by_2_0.tg_magic_3.CLK.t0 5.84563
R12137 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t17 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t6 47.8944
R12138 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t23 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t19 47.8944
R12139 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n1 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t7 47.3388
R12140 p2_gen_magic_0.DFF_magic_0.tg_magic_2.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t12 47.2524
R12141 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n10 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t9 38.7949
R12142 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n11 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t22 38.7949
R12143 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n7 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t21 38.7949
R12144 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n6 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t14 38.7949
R12145 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n11 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n10 31.4949
R12146 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n7 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n6 31.4949
R12147 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n9 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t16 26.9781
R12148 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n9 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t10 26.9781
R12149 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n5 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t15 26.9781
R12150 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n5 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t8 26.9781
R12151 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n0 p2_gen_magic_0.DFF_magic_0.tg_magic_2.CLK 20.617
R12152 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n12 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t11 17.9416
R12153 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n8 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t20 17.9416
R12154 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n12 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t17 11.957
R12155 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n8 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t23 11.957
R12156 p2_gen_magic_0.DFF_magic_0.tg_magic_2.CLK p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n12 10.0908
R12157 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n1 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n8 9.77618
R12158 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n10 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t18 7.3005
R12159 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t11 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n11 7.3005
R12160 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t12 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n9 7.3005
R12161 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n6 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t13 7.3005
R12162 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t20 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n7 7.3005
R12163 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t7 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n5 7.3005
R12164 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n0 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n2 3.6455
R12165 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n0 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n3 3.31072
R12166 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n0 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n4 2.90572
R12167 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n0 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n1 1.72041
R12168 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n3 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t1 1.6255
R12169 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n3 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t0 1.6255
R12170 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n4 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t2 1.6255
R12171 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n4 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t3 1.6255
R12172 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n2 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t4 1.463
R12173 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n2 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t5 1.463
R12174 Q7.t17 Q7.t19 48.5227
R12175 Q7.t7 Q7.t4 47.8944
R12176 Q7.t25 Q7.t21 47.8944
R12177 Q7.t6 Q7.t20 47.5387
R12178 Q7.t24 Q7.t12 47.5387
R12179 Q7.n8 Q7.t23 38.7949
R12180 Q7.n7 Q7.t22 38.7949
R12181 Q7.n4 Q7.t14 38.7949
R12182 Q7.n3 Q7.t13 38.7949
R12183 Q7.n13 Q7.n12 38.5887
R12184 Q7.n13 Q7.n1 34.6748
R12185 Q7.t19 Q7.t11 31.5469
R12186 Q7.n8 Q7.n7 31.4949
R12187 Q7.n4 Q7.n3 31.4949
R12188 Q7.t11 Q7.t10 29.6567
R12189 Q7.n12 Q7.n6 21.1404
R12190 Q7.n9 Q7.t18 17.9416
R12191 Q7.n5 Q7.t8 17.9416
R12192 Q7.n0 Q7.t17 16.8166
R12193 Q7.n10 Q7.t6 15.7085
R12194 Q7.n2 Q7.t24 15.7085
R12195 Q7.n0 Q7.t9 14.7309
R12196 Q7.n1 Q7.n0 13.8453
R12197 Q7.n10 Q7.t3 13.4273
R12198 Q7.n2 Q7.t16 13.4273
R12199 Q7.n9 Q7.t7 11.957
R12200 Q7.n5 Q7.t25 11.957
R12201 Q7 Q7.n9 9.94647
R12202 Q7 Q7.n5 9.94647
R12203 Q7 Q7.n10 8.08021
R12204 Q7 Q7.n2 8.08021
R12205 Q7.n7 Q7.t15 7.3005
R12206 Q7.t18 Q7.n8 7.3005
R12207 Q7.n3 Q7.t5 7.3005
R12208 Q7.t8 Q7.n4 7.3005
R12209 Q7.n15 Q7.t2 5.47387
R12210 Q7.n14 Q7.n13 4.91049
R12211 Q7.n16 Q7.t1 4.65398
R12212 Q7.n12 Q7.n11 4.62973
R12213 Q7.n1 Q7 4.6123
R12214 Q7.n15 Q7.t0 4.2255
R12215 Q7.n11 Q7 3.0464
R12216 Q7.n6 Q7 2.87302
R12217 Q7.n16 Q7.n15 0.427022
R12218 Q7 Q7.n16 0.257096
R12219 Q7.n6 Q7 0.170113
R12220 Q7.n11 Q7 0.0782273
R12221 Q7.n14 Q7 0.030875
R12222 Q7 Q7.n14 0.023
R12223 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t5 130.41
R12224 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n5 36.752
R12225 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t12 35.3186
R12226 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t6 33.5023
R12227 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t8 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n2 33.5023
R12228 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t10 32.2349
R12229 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n0 27.7405
R12230 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t9 26.3866
R12231 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t8 16.3786
R12232 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t9 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n1 13.2317
R12233 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n3 12.5023
R12234 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t4 11.3259
R12235 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t3 11.146
R12236 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t11 7.3005
R12237 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t7 7.3005
R12238 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n4 5.87653
R12239 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t2 5.47387
R12240 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t0 5.28011
R12241 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t1 4.65398
R12242 7b_counter_0.MDFF_4.QB.n1 7b_counter_0.MDFF_4.QB.t7 53.2571
R12243 7b_counter_0.MDFF_4.QB.n4 7b_counter_0.MDFF_4.QB.t6 38.8649
R12244 7b_counter_0.MDFF_4.QB.n3 7b_counter_0.MDFF_4.QB.t4 28.8568
R12245 7b_counter_0.MDFF_4.tspc2_magic_0.QB 7b_counter_0.MDFF_4.QB.n2 23.3781
R12246 7b_counter_0.MDFF_4.tspc2_magic_0.QB 7b_counter_0.MDFF_4.mux_magic_0.IN1 19.5471
R12247 7b_counter_0.MDFF_4.QB.n2 7b_counter_0.MDFF_4.QB.t8 17.1425
R12248 7b_counter_0.MDFF_4.QB.t6 7b_counter_0.MDFF_4.QB.n3 17.0773
R12249 7b_counter_0.MDFF_4.QB.n2 7b_counter_0.MDFF_4.QB.t5 14.405
R12250 7b_counter_0.MDFF_4.QB.n3 7b_counter_0.MDFF_4.QB.t2 11.6023
R12251 7b_counter_0.MDFF_4.mux_magic_0.IN1 7b_counter_0.MDFF_4.QB.n4 9.4273
R12252 7b_counter_0.MDFF_4.QB.n1 7b_counter_0.MDFF_4.QB.n0 8.57932
R12253 7b_counter_0.MDFF_4.QB.n4 7b_counter_0.MDFF_4.QB.t3 7.3005
R12254 7b_counter_0.MDFF_4.QB.t5 7b_counter_0.MDFF_4.QB.n1 7.3005
R12255 7b_counter_0.MDFF_4.QB.n0 7b_counter_0.MDFF_4.QB.t0 3.62007
R12256 7b_counter_0.MDFF_4.QB.n0 7b_counter_0.MDFF_4.QB.t1 3.15478
R12257 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t20 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t22 47.8944
R12258 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t17 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t15 47.8944
R12259 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n1 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t21 47.3388
R12260 7b_counter_0.DFF_magic_0.tg_magic_2.CLK 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t14 47.2524
R12261 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n10 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t12 38.7949
R12262 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n11 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t19 38.7949
R12263 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n7 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t10 38.7949
R12264 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n6 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t23 38.7949
R12265 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n11 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n10 31.4949
R12266 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n7 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n6 31.4949
R12267 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n9 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t16 26.9781
R12268 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n9 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t13 26.9781
R12269 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n5 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t7 26.9781
R12270 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n5 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t18 26.9781
R12271 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n0 7b_counter_0.DFF_magic_0.tg_magic_2.CLK 20.617
R12272 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n12 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t6 17.9416
R12273 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n8 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t11 17.9416
R12274 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n12 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t20 11.957
R12275 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n8 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t17 11.957
R12276 7b_counter_0.DFF_magic_0.tg_magic_2.CLK 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n12 10.0908
R12277 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n1 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n8 9.77618
R12278 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n10 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t8 7.3005
R12279 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t6 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n11 7.3005
R12280 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t14 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n9 7.3005
R12281 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n6 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t9 7.3005
R12282 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t11 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n7 7.3005
R12283 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t21 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n5 7.3005
R12284 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n0 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n2 3.6455
R12285 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n0 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n3 3.31072
R12286 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n0 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n4 2.90572
R12287 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n0 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n1 1.72041
R12288 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n3 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t0 1.6255
R12289 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n3 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t1 1.6255
R12290 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n4 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t3 1.6255
R12291 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n4 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t2 1.6255
R12292 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n2 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t5 1.463
R12293 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n2 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t4 1.463
R12294 Q4.t22 Q4.t21 48.3065
R12295 Q4.t20 Q4.t16 47.8944
R12296 Q4.t29 Q4.t25 47.8944
R12297 Q4.t12 Q4.t7 47.5387
R12298 Q4.t23 Q4.t18 47.5387
R12299 Q4.n18 Q4.n17 46.7373
R12300 Q4.n16 Q4.t3 38.8649
R12301 Q4.n6 Q4.t19 38.7949
R12302 Q4.n5 Q4.t10 38.7949
R12303 Q4.n10 Q4.t28 38.7949
R12304 Q4.n9 Q4.t24 38.7949
R12305 Q4.t21 Q4.t13 31.5469
R12306 Q4.t14 Q4.t22 31.5469
R12307 Q4.n6 Q4.n5 31.4949
R12308 Q4.n10 Q4.n9 31.4949
R12309 Q4.n15 Q4.t4 28.8568
R12310 Q4.n1 Q4.n0 24.5972
R12311 Q4.n14 Q4.n8 24.309
R12312 Q4.n14 Q4.n13 20.7075
R12313 Q4.n18 Q4.n14 20.3093
R12314 Q4 Q4.n1 19.8717
R12315 Q4.n0 Q4.t14 18.2505
R12316 Q4.n7 Q4.t5 17.9416
R12317 Q4.n11 Q4.t15 17.9416
R12318 Q4.t3 Q4.n15 17.0773
R12319 Q4.n4 Q4.t12 15.7085
R12320 Q4.n12 Q4.t23 15.7085
R12321 Q4.n4 Q4.t6 13.4273
R12322 Q4.n12 Q4.t17 13.4273
R12323 Q4.n7 Q4.t20 11.957
R12324 Q4.n11 Q4.t29 11.957
R12325 Q4.n15 Q4.t27 11.6023
R12326 Q4.n0 Q4.t11 11.4067
R12327 Q4 Q4.n7 9.94647
R12328 Q4 Q4.n11 9.94647
R12329 Q4 Q4.n16 9.27587
R12330 Q4 Q4.n4 8.08021
R12331 Q4 Q4.n12 8.08021
R12332 Q4.n16 Q4.t9 7.3005
R12333 Q4.n5 Q4.t26 7.3005
R12334 Q4.t5 Q4.n6 7.3005
R12335 Q4.n9 Q4.t8 7.3005
R12336 Q4.t15 Q4.n10 7.3005
R12337 Q4.n2 Q4.t2 5.47387
R12338 Q4.n3 Q4.t0 4.65398
R12339 Q4.n2 Q4.t1 4.2255
R12340 Q4.n13 Q4 3.06276
R12341 Q4.n19 Q4.n18 2.54473
R12342 Q4.n8 Q4 2.48223
R12343 Q4.n8 Q4 0.602011
R12344 Q4.n3 Q4.n2 0.427022
R12345 Q4.n19 Q4 0.291564
R12346 Q4 Q4.n3 0.257096
R12347 Q4.n17 Q4 0.167977
R12348 Q4.n1 Q4 0.103357
R12349 Q4.n19 Q4 0.0713511
R12350 Q4.n13 Q4 0.0618636
R12351 Q4.n17 Q4 0.0156948
R12352 Q4 Q4.n19 0.00915385
R12353 OR_magic_2.A.t11 OR_magic_2.A.t16 47.8944
R12354 OR_magic_2.A.t6 OR_magic_2.A.t19 44.6331
R12355 OR_magic_2.A.t18 OR_magic_2.A.t15 44.6331
R12356 OR_magic_2.A.n3 OR_magic_2.A.t14 38.7949
R12357 OR_magic_2.A.n4 OR_magic_2.A.t17 38.7949
R12358 OR_magic_2.A.t10 OR_magic_2.A.t20 31.5469
R12359 OR_magic_2.A.t13 OR_magic_2.A.t21 31.5469
R12360 OR_magic_2.A.n4 OR_magic_2.A.n3 31.4949
R12361 OR_magic_2.A.t20 OR_magic_2.A.t9 28.6791
R12362 OR_magic_2.A.t21 OR_magic_2.A.t12 28.6791
R12363 OR_magic_2.A.n6 OR_magic_2.A.t6 19.4237
R12364 OR_magic_2.A.n2 OR_magic_2.A.t18 19.4237
R12365 OR_magic_2.A.n5 OR_magic_2.A.t7 17.9416
R12366 OR_magic_2.A.n0 OR_magic_2.A 13.8488
R12367 OR_magic_2.A.n6 OR_magic_2.A.t10 12.1237
R12368 OR_magic_2.A.n2 OR_magic_2.A.t13 12.1237
R12369 OR_magic_2.A.n5 OR_magic_2.A.t11 11.957
R12370 OR_magic_2.A OR_magic_2.A.n5 9.95929
R12371 OR_magic_2.A OR_magic_2.A.n6 8.23754
R12372 OR_magic_2.A OR_magic_2.A.n2 8.22853
R12373 OR_magic_2.A.n3 OR_magic_2.A.t8 7.3005
R12374 OR_magic_2.A.t7 OR_magic_2.A.n4 7.3005
R12375 OR_magic_2.A.n1 OR_magic_2.A.n7 3.6455
R12376 OR_magic_2.A.n1 OR_magic_2.A.n8 3.31072
R12377 OR_magic_2.A.n1 OR_magic_2.A.n9 2.90572
R12378 OR_magic_2.A.n8 OR_magic_2.A.t2 1.6255
R12379 OR_magic_2.A.n8 OR_magic_2.A.t1 1.6255
R12380 OR_magic_2.A.n9 OR_magic_2.A.t0 1.6255
R12381 OR_magic_2.A.n9 OR_magic_2.A.t3 1.6255
R12382 OR_magic_2.A.n7 OR_magic_2.A.t5 1.463
R12383 OR_magic_2.A.n7 OR_magic_2.A.t4 1.463
R12384 OR_magic_2.A.n0 OR_magic_2.A 1.25072
R12385 OR_magic_2.A.n1 OR_magic_2.A.n0 1.22536
R12386 p2_gen_magic_0.3_inp_AND_magic_0.C.n1 p2_gen_magic_0.3_inp_AND_magic_0.C.t5 39.1562
R12387 p2_gen_magic_0.3_inp_AND_magic_0.C.t1 p2_gen_magic_0.3_inp_AND_magic_0.C.t2 28.8746
R12388 p2_gen_magic_0.3_inp_AND_magic_0.C.t5 p2_gen_magic_0.3_inp_AND_magic_0.C.t3 23.4648
R12389 p2_gen_magic_0.3_inp_AND_magic_0.C.n0 p2_gen_magic_0.3_inp_AND_magic_0.C.t4 14.1443
R12390 p2_gen_magic_0.3_inp_AND_magic_0.C.n0 p2_gen_magic_0.3_inp_AND_magic_0.C.t1 13.8835
R12391 p2_gen_magic_0.3_inp_AND_magic_0.C.n1 p2_gen_magic_0.3_inp_AND_magic_0.C.n0 12.5017
R12392 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.3_inp_AND_magic_0.C.n1 5.35629
R12393 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.3_inp_AND_magic_0.C.t0 3.46108
R12394 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t3 15.4558
R12395 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n0 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t10 5.68115
R12396 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 5.47974
R12397 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t0 4.928
R12398 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t5 4.66963
R12399 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t6 4.2255
R12400 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n0 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 3.1505
R12401 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t4 p3_gen_magic_0.3_inp_AND_magic_0.VOUT 3.12083
R12402 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n0 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 2.6005
R12403 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n0 2.31651
R12404 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t8 1.6255
R12405 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t9 1.6255
R12406 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t1 1.463
R12407 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t2 1.463
R12408 OR_magic_1.VOUT.t13 OR_magic_1.VOUT.t15 47.8944
R12409 OR_magic_1.VOUT.t24 OR_magic_1.VOUT.t17 47.8944
R12410 OR_magic_1.VOUT.t22 OR_magic_1.VOUT.t14 47.8944
R12411 OR_magic_1.VOUT.n0 OR_magic_1.VOUT.t23 47.3388
R12412 OR_magic_1.VOUT.n9 OR_magic_1.VOUT.t3 38.7949
R12413 OR_magic_1.VOUT.n10 OR_magic_1.VOUT.t19 38.7949
R12414 OR_magic_1.VOUT.n6 OR_magic_1.VOUT.t20 38.7949
R12415 OR_magic_1.VOUT.n5 OR_magic_1.VOUT.t8 38.7949
R12416 OR_magic_1.VOUT.n2 OR_magic_1.VOUT.t10 38.7949
R12417 OR_magic_1.VOUT.n1 OR_magic_1.VOUT.t4 38.7949
R12418 OR_magic_1.VOUT.n10 OR_magic_1.VOUT.n9 31.4949
R12419 OR_magic_1.VOUT.n6 OR_magic_1.VOUT.n5 31.4949
R12420 OR_magic_1.VOUT.n2 OR_magic_1.VOUT.n1 31.4949
R12421 OR_magic_1.VOUT OR_magic_1.VOUT.t11 31.3561
R12422 OR_magic_1.VOUT.n8 OR_magic_1.VOUT.t9 26.9781
R12423 OR_magic_1.VOUT.n8 OR_magic_1.VOUT.t25 26.9781
R12424 OR_magic_1.VOUT.n4 OR_magic_1.VOUT.t5 26.9781
R12425 OR_magic_1.VOUT.n4 OR_magic_1.VOUT.t21 26.9781
R12426 OR_magic_1.VOUT.n11 OR_magic_1.VOUT.t7 17.9416
R12427 OR_magic_1.VOUT.n7 OR_magic_1.VOUT.t18 17.9416
R12428 OR_magic_1.VOUT.n3 OR_magic_1.VOUT.t16 17.9416
R12429 OR_magic_1.VOUT.n0 OR_magic_1.VOUT 12.5623
R12430 OR_magic_1.VOUT.n11 OR_magic_1.VOUT.t13 11.957
R12431 OR_magic_1.VOUT.n7 OR_magic_1.VOUT.t24 11.957
R12432 OR_magic_1.VOUT.n3 OR_magic_1.VOUT.t22 11.957
R12433 OR_magic_1.VOUT OR_magic_1.VOUT.n11 10.0013
R12434 OR_magic_1.VOUT OR_magic_1.VOUT.n3 9.96162
R12435 OR_magic_1.VOUT.n0 OR_magic_1.VOUT.n7 9.77618
R12436 OR_magic_1.VOUT.n12 OR_magic_1.VOUT.n0 8.71923
R12437 OR_magic_1.VOUT.n9 OR_magic_1.VOUT.t2 7.3005
R12438 OR_magic_1.VOUT.t7 OR_magic_1.VOUT.n10 7.3005
R12439 OR_magic_1.VOUT.t11 OR_magic_1.VOUT.n8 7.3005
R12440 OR_magic_1.VOUT.n5 OR_magic_1.VOUT.t12 7.3005
R12441 OR_magic_1.VOUT.t18 OR_magic_1.VOUT.n6 7.3005
R12442 OR_magic_1.VOUT.t23 OR_magic_1.VOUT.n4 7.3005
R12443 OR_magic_1.VOUT.n1 OR_magic_1.VOUT.t6 7.3005
R12444 OR_magic_1.VOUT.t16 OR_magic_1.VOUT.n2 7.3005
R12445 OR_magic_1.VOUT OR_magic_1.VOUT.t1 5.47387
R12446 OR_magic_1.VOUT OR_magic_1.VOUT.t0 4.2255
R12447 OR_magic_1.VOUT.n12 OR_magic_1.VOUT 3.44007
R12448 OR_magic_1.VOUT OR_magic_1.VOUT.n12 2.96809
R12449 divide_by_2_0.tg_magic_3.IN.t20 divide_by_2_0.tg_magic_3.IN.t22 47.8944
R12450 divide_by_2_0.tg_magic_3.IN.n5 divide_by_2_0.tg_magic_3.IN.t18 38.7949
R12451 divide_by_2_0.tg_magic_3.IN.n4 divide_by_2_0.tg_magic_3.IN.t23 38.7949
R12452 divide_by_2_0.tg_magic_3.IN.n5 divide_by_2_0.tg_magic_3.IN.n4 31.4949
R12453 divide_by_2_0.tg_magic_3.IN.n6 divide_by_2_0.tg_magic_3.IN.t21 17.9416
R12454 divide_by_2_0.tg_magic_3.IN.n6 divide_by_2_0.tg_magic_3.IN.t20 11.957
R12455 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.n6 9.96162
R12456 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.n3 9.59884
R12457 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.n11 9.59884
R12458 divide_by_2_0.tg_magic_3.IN.n4 divide_by_2_0.tg_magic_3.IN.t19 7.3005
R12459 divide_by_2_0.tg_magic_3.IN.t21 divide_by_2_0.tg_magic_3.IN.n5 7.3005
R12460 divide_by_2_0.tg_magic_3.IN.n0 divide_by_2_0.tg_magic_3.IN.t16 5.68115
R12461 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.t1 5.34258
R12462 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.t14 4.96909
R12463 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.t8 4.96909
R12464 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.t5 4.928
R12465 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.t10 4.8305
R12466 divide_by_2_0.tg_magic_3.IN.n3 divide_by_2_0.tg_magic_3.IN.n1 3.99516
R12467 divide_by_2_0.tg_magic_3.IN.n11 divide_by_2_0.tg_magic_3.IN.n10 3.99516
R12468 divide_by_2_0.tg_magic_3.IN.n0 divide_by_2_0.tg_magic_3.IN.n8 3.1505
R12469 divide_by_2_0.tg_magic_3.IN.n3 divide_by_2_0.tg_magic_3.IN.n2 2.60841
R12470 divide_by_2_0.tg_magic_3.IN.n11 divide_by_2_0.tg_magic_3.IN.n9 2.60841
R12471 divide_by_2_0.tg_magic_3.IN.n0 divide_by_2_0.tg_magic_3.IN.n7 2.6005
R12472 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_3.IN.n0 2.31898
R12473 divide_by_2_0.tg_magic_3.IN.n7 divide_by_2_0.tg_magic_3.IN.t15 1.6255
R12474 divide_by_2_0.tg_magic_3.IN.n7 divide_by_2_0.tg_magic_3.IN.t17 1.6255
R12475 divide_by_2_0.tg_magic_3.IN.n2 divide_by_2_0.tg_magic_3.IN.t12 1.6255
R12476 divide_by_2_0.tg_magic_3.IN.n2 divide_by_2_0.tg_magic_3.IN.t11 1.6255
R12477 divide_by_2_0.tg_magic_3.IN.n9 divide_by_2_0.tg_magic_3.IN.t0 1.6255
R12478 divide_by_2_0.tg_magic_3.IN.n9 divide_by_2_0.tg_magic_3.IN.t2 1.6255
R12479 divide_by_2_0.tg_magic_3.IN.n8 divide_by_2_0.tg_magic_3.IN.t4 1.463
R12480 divide_by_2_0.tg_magic_3.IN.n8 divide_by_2_0.tg_magic_3.IN.t6 1.463
R12481 divide_by_2_0.tg_magic_3.IN.n1 divide_by_2_0.tg_magic_3.IN.t7 1.463
R12482 divide_by_2_0.tg_magic_3.IN.n1 divide_by_2_0.tg_magic_3.IN.t9 1.463
R12483 divide_by_2_0.tg_magic_3.IN.n10 divide_by_2_0.tg_magic_3.IN.t3 1.463
R12484 divide_by_2_0.tg_magic_3.IN.n10 divide_by_2_0.tg_magic_3.IN.t13 1.463
R12485 a_27567_8496.n1 a_27567_8496.t17 39.6673
R12486 a_27567_8496.t15 a_27567_8496.n1 39.6673
R12487 a_27567_8496.n2 a_27567_8496.t9 39.3349
R12488 a_27567_8496.t13 a_27567_8496.n2 39.3349
R12489 a_27567_8496.t10 a_27567_8496.t15 31.0255
R12490 a_27567_8496.t16 a_27567_8496.t12 31.0255
R12491 a_27567_8496.t9 a_27567_8496.t10 29.1353
R12492 a_27567_8496.t12 a_27567_8496.t11 29.1353
R12493 a_27567_8496.t14 a_27567_8496.t13 29.1353
R12494 a_27567_8496.n3 a_27567_8496.t17 13.6103
R12495 a_27567_8496.n3 a_27567_8496.t14 12.9295
R12496 a_27567_8496.n6 a_27567_8496.n4 9.66932
R12497 a_27567_8496.n11 a_27567_8496.n10 9.63981
R12498 a_27567_8496.n0 a_27567_8496.n3 8.42281
R12499 a_27567_8496.n1 a_27567_8496.t16 7.3005
R12500 a_27567_8496.n2 a_27567_8496.t11 7.3005
R12501 a_27567_8496.n11 a_27567_8496.t8 4.62001
R12502 a_27567_8496.n4 a_27567_8496.t2 4.2255
R12503 a_27567_8496.t5 a_27567_8496.n0 4.2255
R12504 a_27567_8496.n10 a_27567_8496.n9 3.16569
R12505 a_27567_8496.n6 a_27567_8496.n5 2.6005
R12506 a_27567_8496.n8 a_27567_8496.n7 2.6005
R12507 a_27567_8496.n7 a_27567_8496.t4 1.6255
R12508 a_27567_8496.n7 a_27567_8496.t3 1.6255
R12509 a_27567_8496.n5 a_27567_8496.t1 1.6255
R12510 a_27567_8496.n5 a_27567_8496.t0 1.6255
R12511 a_27567_8496.n9 a_27567_8496.t7 1.463
R12512 a_27567_8496.n9 a_27567_8496.t6 1.463
R12513 a_27567_8496.n8 a_27567_8496.n6 0.913343
R12514 a_27567_8496.n0 a_27567_8496.n11 0.832606
R12515 a_27567_8496.n10 a_27567_8496.n8 0.818911
R12516 a_27567_8496.n4 a_27567_8496.n0 0.810801
R12517 a_31440_8496.n1 a_31440_8496.t9 39.6673
R12518 a_31440_8496.t16 a_31440_8496.n1 39.6673
R12519 a_31440_8496.n2 a_31440_8496.t10 39.3349
R12520 a_31440_8496.t14 a_31440_8496.n2 39.3349
R12521 a_31440_8496.t11 a_31440_8496.t16 31.0255
R12522 a_31440_8496.t17 a_31440_8496.t13 31.0255
R12523 a_31440_8496.t10 a_31440_8496.t11 29.1353
R12524 a_31440_8496.t13 a_31440_8496.t12 29.1353
R12525 a_31440_8496.t15 a_31440_8496.t14 29.1353
R12526 a_31440_8496.n3 a_31440_8496.t9 13.6103
R12527 a_31440_8496.n3 a_31440_8496.t15 12.9295
R12528 a_31440_8496.n6 a_31440_8496.n4 9.66932
R12529 a_31440_8496.n11 a_31440_8496.n10 9.63981
R12530 a_31440_8496.n0 a_31440_8496.n3 8.42281
R12531 a_31440_8496.n1 a_31440_8496.t17 7.3005
R12532 a_31440_8496.n2 a_31440_8496.t12 7.3005
R12533 a_31440_8496.n11 a_31440_8496.t8 4.62001
R12534 a_31440_8496.n4 a_31440_8496.t2 4.2255
R12535 a_31440_8496.t5 a_31440_8496.n0 4.2255
R12536 a_31440_8496.n10 a_31440_8496.n9 3.16569
R12537 a_31440_8496.n6 a_31440_8496.n5 2.6005
R12538 a_31440_8496.n8 a_31440_8496.n7 2.6005
R12539 a_31440_8496.n7 a_31440_8496.t4 1.6255
R12540 a_31440_8496.n7 a_31440_8496.t3 1.6255
R12541 a_31440_8496.n5 a_31440_8496.t1 1.6255
R12542 a_31440_8496.n5 a_31440_8496.t0 1.6255
R12543 a_31440_8496.n9 a_31440_8496.t7 1.463
R12544 a_31440_8496.n9 a_31440_8496.t6 1.463
R12545 a_31440_8496.n8 a_31440_8496.n6 0.913343
R12546 a_31440_8496.n0 a_31440_8496.n11 0.832606
R12547 a_31440_8496.n10 a_31440_8496.n8 0.818911
R12548 a_31440_8496.n4 a_31440_8496.n0 0.810801
R12549 p3_gen_magic_0.xnor_magic_5.OUT.t3 p3_gen_magic_0.xnor_magic_5.OUT.t5 144.929
R12550 p3_gen_magic_0.xnor_magic_5.OUT.n0 p3_gen_magic_0.xnor_magic_5.OUT.t4 24.9839
R12551 p3_gen_magic_0.xnor_magic_5.OUT.n2 p3_gen_magic_0.xnor_magic_5.OUT 24.6161
R12552 p3_gen_magic_0.xnor_magic_5.OUT.n1 p3_gen_magic_0.xnor_magic_5.OUT.t3 14.7678
R12553 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_5.OUT.n1 13.7481
R12554 p3_gen_magic_0.xnor_magic_5.OUT.n0 p3_gen_magic_0.xnor_magic_5.OUT.t2 11.3906
R12555 p3_gen_magic_0.xnor_magic_5.OUT.n2 p3_gen_magic_0.xnor_magic_5.OUT.t1 9.23184
R12556 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_5.OUT.n2 5.86488
R12557 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_5.OUT.t0 2.96833
R12558 p3_gen_magic_0.xnor_magic_5.OUT.n1 p3_gen_magic_0.xnor_magic_5.OUT.n0 2.45537
R12559 divide_by_2_1.tg_magic_3.IN.t23 divide_by_2_1.tg_magic_3.IN.t20 47.8944
R12560 divide_by_2_1.tg_magic_3.IN.n5 divide_by_2_1.tg_magic_3.IN.t22 38.7949
R12561 divide_by_2_1.tg_magic_3.IN.n4 divide_by_2_1.tg_magic_3.IN.t18 38.7949
R12562 divide_by_2_1.tg_magic_3.IN.n5 divide_by_2_1.tg_magic_3.IN.n4 31.4949
R12563 divide_by_2_1.tg_magic_3.IN.n6 divide_by_2_1.tg_magic_3.IN.t21 17.9416
R12564 divide_by_2_1.tg_magic_3.IN.n6 divide_by_2_1.tg_magic_3.IN.t23 11.957
R12565 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.n6 9.96162
R12566 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.n11 9.59884
R12567 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.n3 9.59884
R12568 divide_by_2_1.tg_magic_3.IN.n4 divide_by_2_1.tg_magic_3.IN.t19 7.3005
R12569 divide_by_2_1.tg_magic_3.IN.t21 divide_by_2_1.tg_magic_3.IN.n5 7.3005
R12570 divide_by_2_1.tg_magic_3.IN.n0 divide_by_2_1.tg_magic_3.IN.t15 5.68115
R12571 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.t2 5.34258
R12572 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.t4 4.96909
R12573 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.t13 4.96909
R12574 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.t9 4.928
R12575 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.t8 4.8305
R12576 divide_by_2_1.tg_magic_3.IN.n11 divide_by_2_1.tg_magic_3.IN.n10 3.99516
R12577 divide_by_2_1.tg_magic_3.IN.n3 divide_by_2_1.tg_magic_3.IN.n1 3.99516
R12578 divide_by_2_1.tg_magic_3.IN.n0 divide_by_2_1.tg_magic_3.IN.n8 3.1505
R12579 divide_by_2_1.tg_magic_3.IN.n11 divide_by_2_1.tg_magic_3.IN.n9 2.60841
R12580 divide_by_2_1.tg_magic_3.IN.n3 divide_by_2_1.tg_magic_3.IN.n2 2.60841
R12581 divide_by_2_1.tg_magic_3.IN.n0 divide_by_2_1.tg_magic_3.IN.n7 2.6005
R12582 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_3.IN.n0 2.31898
R12583 divide_by_2_1.tg_magic_3.IN.n9 divide_by_2_1.tg_magic_3.IN.t1 1.6255
R12584 divide_by_2_1.tg_magic_3.IN.n9 divide_by_2_1.tg_magic_3.IN.t0 1.6255
R12585 divide_by_2_1.tg_magic_3.IN.n7 divide_by_2_1.tg_magic_3.IN.t17 1.6255
R12586 divide_by_2_1.tg_magic_3.IN.n7 divide_by_2_1.tg_magic_3.IN.t16 1.6255
R12587 divide_by_2_1.tg_magic_3.IN.n2 divide_by_2_1.tg_magic_3.IN.t6 1.6255
R12588 divide_by_2_1.tg_magic_3.IN.n2 divide_by_2_1.tg_magic_3.IN.t7 1.6255
R12589 divide_by_2_1.tg_magic_3.IN.n10 divide_by_2_1.tg_magic_3.IN.t3 1.463
R12590 divide_by_2_1.tg_magic_3.IN.n10 divide_by_2_1.tg_magic_3.IN.t5 1.463
R12591 divide_by_2_1.tg_magic_3.IN.n8 divide_by_2_1.tg_magic_3.IN.t11 1.463
R12592 divide_by_2_1.tg_magic_3.IN.n8 divide_by_2_1.tg_magic_3.IN.t10 1.463
R12593 divide_by_2_1.tg_magic_3.IN.n1 divide_by_2_1.tg_magic_3.IN.t12 1.463
R12594 divide_by_2_1.tg_magic_3.IN.n1 divide_by_2_1.tg_magic_3.IN.t14 1.463
R12595 mux_magic_0.IN1.t8 mux_magic_0.IN1.t11 47.8944
R12596 mux_magic_0.IN1.n1 mux_magic_0.IN1.t12 38.8649
R12597 mux_magic_0.IN1.n2 mux_magic_0.IN1.t14 38.7949
R12598 mux_magic_0.IN1.n3 mux_magic_0.IN1.t13 38.7949
R12599 mux_magic_0.IN1.n3 mux_magic_0.IN1.n2 31.4949
R12600 mux_magic_0.IN1.n0 mux_magic_0.IN1.t6 28.8568
R12601 mux_magic_0.IN1.n4 mux_magic_0.IN1.t10 17.9416
R12602 mux_magic_0.IN1.t12 mux_magic_0.IN1.n0 17.0773
R12603 mux_magic_0.IN1.n4 mux_magic_0.IN1.t8 11.957
R12604 mux_magic_0.IN1.n0 mux_magic_0.IN1.t7 11.6023
R12605 mux_magic_0.IN1 mux_magic_0.IN1.n4 9.95929
R12606 mux_magic_0.IN1 mux_magic_0.IN1.n1 9.40996
R12607 mux_magic_0.IN1.n1 mux_magic_0.IN1.t15 7.3005
R12608 mux_magic_0.IN1.n2 mux_magic_0.IN1.t9 7.3005
R12609 mux_magic_0.IN1.t10 mux_magic_0.IN1.n3 7.3005
R12610 mux_magic_0.IN1 mux_magic_0.IN1.n5 3.6455
R12611 mux_magic_0.IN1 mux_magic_0.IN1.n6 3.31072
R12612 mux_magic_0.IN1 mux_magic_0.IN1.n7 2.90572
R12613 mux_magic_0.IN1.n6 mux_magic_0.IN1.t1 1.6255
R12614 mux_magic_0.IN1.n6 mux_magic_0.IN1.t0 1.6255
R12615 mux_magic_0.IN1.n7 mux_magic_0.IN1.t3 1.6255
R12616 mux_magic_0.IN1.n7 mux_magic_0.IN1.t2 1.6255
R12617 mux_magic_0.IN1.n5 mux_magic_0.IN1.t5 1.463
R12618 mux_magic_0.IN1.n5 mux_magic_0.IN1.t4 1.463
R12619 p3_gen_magic_0.xnor_magic_3.OUT.n0 p3_gen_magic_0.xnor_magic_3.OUT.t5 39.1562
R12620 p3_gen_magic_0.xnor_magic_3.OUT.t3 p3_gen_magic_0.xnor_magic_3.OUT.t2 28.8746
R12621 p3_gen_magic_0.xnor_magic_3.OUT.t5 p3_gen_magic_0.xnor_magic_3.OUT.t6 23.4648
R12622 p3_gen_magic_0.xnor_magic_3.OUT.n2 p3_gen_magic_0.xnor_magic_3.OUT.n0 17.1813
R12623 p3_gen_magic_0.xnor_magic_3.OUT.n1 p3_gen_magic_0.xnor_magic_3.OUT.t4 14.1443
R12624 p3_gen_magic_0.xnor_magic_3.OUT.n1 p3_gen_magic_0.xnor_magic_3.OUT.t3 13.8835
R12625 p3_gen_magic_0.xnor_magic_3.OUT.n0 p3_gen_magic_0.xnor_magic_3.OUT.n1 12.5017
R12626 p3_gen_magic_0.xnor_magic_3.OUT.n2 p3_gen_magic_0.xnor_magic_3.OUT.t1 9.23184
R12627 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.OUT.n2 5.86488
R12628 p3_gen_magic_0.xnor_magic_3.OUT.n0 p3_gen_magic_0.xnor_magic_3.OUT 5.43085
R12629 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.OUT.t0 3.11311
R12630 Q5.n18 Q5.n17 52.1474
R12631 Q5.t4 Q5.t14 48.5227
R12632 Q5.t13 Q5.t9 47.8944
R12633 Q5.t23 Q5.t17 47.8944
R12634 Q5.t16 Q5.t10 47.5387
R12635 Q5.t24 Q5.t19 47.5387
R12636 Q5.n3 Q5.t28 38.8649
R12637 Q5.n14 Q5.t11 38.7949
R12638 Q5.n13 Q5.t12 38.7949
R12639 Q5.n9 Q5.t21 38.7949
R12640 Q5.n8 Q5.t22 38.7949
R12641 Q5.n19 Q5 34.8562
R12642 Q5.n5 Q5.n4 32.6541
R12643 Q5.t14 Q5.t5 31.5469
R12644 Q5.n14 Q5.n13 31.4949
R12645 Q5.n9 Q5.n8 31.4949
R12646 Q5.t5 Q5.t3 29.6567
R12647 Q5.n2 Q5.t7 28.8568
R12648 Q5 Q5.n7 18.475
R12649 Q5.n15 Q5.t25 17.9416
R12650 Q5.n10 Q5.t6 17.9416
R12651 Q5.t28 Q5.n2 17.0773
R12652 Q5.n7 Q5.t4 16.8166
R12653 Q5.n16 Q5.t16 15.7085
R12654 Q5.n11 Q5.t24 15.7085
R12655 Q5.n7 Q5.t27 14.7309
R12656 Q5.n16 Q5.t8 13.4273
R12657 Q5.n11 Q5.t18 13.4273
R12658 Q5.n19 Q5.n18 12.6085
R12659 Q5.n15 Q5.t13 11.957
R12660 Q5.n10 Q5.t23 11.957
R12661 Q5.n2 Q5.t15 11.6023
R12662 Q5.n18 Q5.n12 10.443
R12663 Q5 Q5.n15 9.94647
R12664 Q5 Q5.n10 9.94647
R12665 Q5 Q5.n3 9.27587
R12666 Q5 Q5.n16 8.08021
R12667 Q5 Q5.n11 8.08021
R12668 Q5.n3 Q5.t26 7.3005
R12669 Q5.n13 Q5.t20 7.3005
R12670 Q5.t25 Q5.n14 7.3005
R12671 Q5.n8 Q5.t29 7.3005
R12672 Q5.t6 Q5.n9 7.3005
R12673 Q5.n0 Q5.t2 5.47387
R12674 Q5.n1 Q5.t1 4.65398
R12675 Q5.n0 Q5.t0 4.2255
R12676 Q5.n12 Q5 2.12624
R12677 Q5.n17 Q5 1.96503
R12678 Q5 Q5.n19 1.43232
R12679 Q5.n17 Q5 1.15959
R12680 Q5.n12 Q5 0.939564
R12681 Q5.n1 Q5.n0 0.427022
R12682 Q5 Q5.n1 0.257096
R12683 Q5 Q5.n6 0.113409
R12684 Q5.n5 Q5 0.02675
R12685 Q5.n6 Q5 0.02425
R12686 Q5.n4 Q5 0.0182778
R12687 Q5.n6 Q5.n5 0.00925
R12688 Q5.n4 Q5 0.00161111
R12689 DFF_magic_0.tg_magic_3.CLK.t18 DFF_magic_0.tg_magic_3.CLK.t16 47.8944
R12690 DFF_magic_0.tg_magic_3.CLK.t15 DFF_magic_0.tg_magic_3.CLK.t11 47.8944
R12691 DFF_magic_0.tg_magic_3.CLK.n1 DFF_magic_0.tg_magic_3.CLK.t14 47.3388
R12692 DFF_magic_0.tg_magic_2.CLK DFF_magic_0.tg_magic_3.CLK.t13 47.2524
R12693 DFF_magic_0.tg_magic_3.CLK.n10 DFF_magic_0.tg_magic_3.CLK.t20 38.7949
R12694 DFF_magic_0.tg_magic_3.CLK.n11 DFF_magic_0.tg_magic_3.CLK.t23 38.7949
R12695 DFF_magic_0.tg_magic_3.CLK.n7 DFF_magic_0.tg_magic_3.CLK.t22 38.7949
R12696 DFF_magic_0.tg_magic_3.CLK.n6 DFF_magic_0.tg_magic_3.CLK.t19 38.7949
R12697 DFF_magic_0.tg_magic_3.CLK.n11 DFF_magic_0.tg_magic_3.CLK.n10 31.4949
R12698 DFF_magic_0.tg_magic_3.CLK.n7 DFF_magic_0.tg_magic_3.CLK.n6 31.4949
R12699 DFF_magic_0.tg_magic_3.CLK.n9 DFF_magic_0.tg_magic_3.CLK.t17 26.9781
R12700 DFF_magic_0.tg_magic_3.CLK.n9 DFF_magic_0.tg_magic_3.CLK.t10 26.9781
R12701 DFF_magic_0.tg_magic_3.CLK.n5 DFF_magic_0.tg_magic_3.CLK.t6 26.9781
R12702 DFF_magic_0.tg_magic_3.CLK.n5 DFF_magic_0.tg_magic_3.CLK.t9 26.9781
R12703 DFF_magic_0.tg_magic_3.CLK.n0 DFF_magic_0.tg_magic_2.CLK 20.617
R12704 DFF_magic_0.tg_magic_3.CLK.n12 DFF_magic_0.tg_magic_3.CLK.t12 17.9416
R12705 DFF_magic_0.tg_magic_3.CLK.n8 DFF_magic_0.tg_magic_3.CLK.t7 17.9416
R12706 DFF_magic_0.tg_magic_3.CLK.n12 DFF_magic_0.tg_magic_3.CLK.t18 11.957
R12707 DFF_magic_0.tg_magic_3.CLK.n8 DFF_magic_0.tg_magic_3.CLK.t15 11.957
R12708 DFF_magic_0.tg_magic_2.CLK DFF_magic_0.tg_magic_3.CLK.n12 10.0908
R12709 DFF_magic_0.tg_magic_3.CLK.n1 DFF_magic_0.tg_magic_3.CLK.n8 9.77618
R12710 DFF_magic_0.tg_magic_3.CLK.n10 DFF_magic_0.tg_magic_3.CLK.t8 7.3005
R12711 DFF_magic_0.tg_magic_3.CLK.t12 DFF_magic_0.tg_magic_3.CLK.n11 7.3005
R12712 DFF_magic_0.tg_magic_3.CLK.t13 DFF_magic_0.tg_magic_3.CLK.n9 7.3005
R12713 DFF_magic_0.tg_magic_3.CLK.n6 DFF_magic_0.tg_magic_3.CLK.t21 7.3005
R12714 DFF_magic_0.tg_magic_3.CLK.t7 DFF_magic_0.tg_magic_3.CLK.n7 7.3005
R12715 DFF_magic_0.tg_magic_3.CLK.t14 DFF_magic_0.tg_magic_3.CLK.n5 7.3005
R12716 DFF_magic_0.tg_magic_3.CLK.n0 DFF_magic_0.tg_magic_3.CLK.n3 3.6455
R12717 DFF_magic_0.tg_magic_3.CLK.n0 DFF_magic_0.tg_magic_3.CLK.n4 3.31072
R12718 DFF_magic_0.tg_magic_3.CLK.n0 DFF_magic_0.tg_magic_3.CLK.n2 2.90572
R12719 DFF_magic_0.tg_magic_3.CLK.n0 DFF_magic_0.tg_magic_3.CLK.n1 1.72041
R12720 DFF_magic_0.tg_magic_3.CLK.n2 DFF_magic_0.tg_magic_3.CLK.t2 1.6255
R12721 DFF_magic_0.tg_magic_3.CLK.n2 DFF_magic_0.tg_magic_3.CLK.t1 1.6255
R12722 DFF_magic_0.tg_magic_3.CLK.n4 DFF_magic_0.tg_magic_3.CLK.t3 1.6255
R12723 DFF_magic_0.tg_magic_3.CLK.n4 DFF_magic_0.tg_magic_3.CLK.t0 1.6255
R12724 DFF_magic_0.tg_magic_3.CLK.n3 DFF_magic_0.tg_magic_3.CLK.t5 1.463
R12725 DFF_magic_0.tg_magic_3.CLK.n3 DFF_magic_0.tg_magic_3.CLK.t4 1.463
R12726 7b_counter_0.MDFF_7.QB.n1 7b_counter_0.MDFF_7.QB.t2 53.0329
R12727 7b_counter_0.MDFF_7.QB.n4 7b_counter_0.MDFF_7.QB.t6 38.8649
R12728 7b_counter_0.MDFF_7.QB.n3 7b_counter_0.MDFF_7.QB.t4 28.8568
R12729 7b_counter_0.MDFF_7.tspc2_magic_0.QB 7b_counter_0.MDFF_7.QB.n2 23.3781
R12730 7b_counter_0.MDFF_7.tspc2_magic_0.QB 7b_counter_0.MDFF_7.mux_magic_0.IN1 20.673
R12731 7b_counter_0.MDFF_7.QB.n2 7b_counter_0.MDFF_7.QB.t8 17.2076
R12732 7b_counter_0.MDFF_7.QB.t6 7b_counter_0.MDFF_7.QB.n3 17.0773
R12733 7b_counter_0.MDFF_7.QB.n2 7b_counter_0.MDFF_7.QB.t5 14.3398
R12734 7b_counter_0.MDFF_7.QB.n3 7b_counter_0.MDFF_7.QB.t3 11.6023
R12735 7b_counter_0.MDFF_7.mux_magic_0.IN1 7b_counter_0.MDFF_7.QB.n4 9.4249
R12736 7b_counter_0.MDFF_7.QB.n1 7b_counter_0.MDFF_7.QB.n0 8.57932
R12737 7b_counter_0.MDFF_7.QB.n4 7b_counter_0.MDFF_7.QB.t7 7.3005
R12738 7b_counter_0.MDFF_7.QB.t5 7b_counter_0.MDFF_7.QB.n1 7.3005
R12739 7b_counter_0.MDFF_7.QB.n0 7b_counter_0.MDFF_7.QB.t0 3.62007
R12740 7b_counter_0.MDFF_7.QB.n0 7b_counter_0.MDFF_7.QB.t1 3.15478
R12741 p3_gen_magic_0.xnor_magic_1.OUT.n2 p3_gen_magic_0.xnor_magic_1.OUT 39.3953
R12742 p3_gen_magic_0.xnor_magic_1.OUT.n1 p3_gen_magic_0.xnor_magic_1.OUT.t4 38.8649
R12743 p3_gen_magic_0.xnor_magic_1.OUT.n0 p3_gen_magic_0.xnor_magic_1.OUT.t5 28.8568
R12744 p3_gen_magic_0.xnor_magic_1.OUT.t4 p3_gen_magic_0.xnor_magic_1.OUT.n0 17.0773
R12745 p3_gen_magic_0.xnor_magic_1.OUT.n0 p3_gen_magic_0.xnor_magic_1.OUT.t6 11.6023
R12746 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_1.OUT.n1 9.27587
R12747 p3_gen_magic_0.xnor_magic_1.OUT.n2 p3_gen_magic_0.xnor_magic_1.OUT.t1 9.23184
R12748 p3_gen_magic_0.xnor_magic_1.OUT.n1 p3_gen_magic_0.xnor_magic_1.OUT.t3 7.3005
R12749 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_1.OUT.n2 5.86488
R12750 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_1.OUT.t2 3.10137
R12751 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_1.OUT.t0 2.96833
R12752 7b_counter_0.MDFF_1.QB.n3 7b_counter_0.MDFF_1.QB.t8 53.2954
R12753 7b_counter_0.MDFF_1.QB.n1 7b_counter_0.MDFF_1.QB.t6 38.8649
R12754 7b_counter_0.MDFF_1.QB.n0 7b_counter_0.MDFF_1.QB.t5 28.8568
R12755 7b_counter_0.MDFF_1.tspc2_magic_0.QB 7b_counter_0.MDFF_1.QB.n4 23.3781
R12756 7b_counter_0.MDFF_1.tspc2_magic_0.QB 7b_counter_0.MDFF_1.mux_magic_0.IN1 19.4019
R12757 7b_counter_0.MDFF_1.QB.n4 7b_counter_0.MDFF_1.QB.t2 17.1425
R12758 7b_counter_0.MDFF_1.QB.t6 7b_counter_0.MDFF_1.QB.n0 17.0773
R12759 7b_counter_0.MDFF_1.QB.n4 7b_counter_0.MDFF_1.QB.t4 14.405
R12760 7b_counter_0.MDFF_1.QB.n0 7b_counter_0.MDFF_1.QB.t3 11.6023
R12761 7b_counter_0.MDFF_1.mux_magic_0.IN1 7b_counter_0.MDFF_1.QB.n1 9.42776
R12762 7b_counter_0.MDFF_1.QB.n3 7b_counter_0.MDFF_1.QB.n2 8.51584
R12763 7b_counter_0.MDFF_1.QB.n1 7b_counter_0.MDFF_1.QB.t7 7.3005
R12764 7b_counter_0.MDFF_1.QB.t4 7b_counter_0.MDFF_1.QB.n3 7.3005
R12765 7b_counter_0.MDFF_1.QB.n2 7b_counter_0.MDFF_1.QB.t0 3.62007
R12766 7b_counter_0.MDFF_1.QB.n2 7b_counter_0.MDFF_1.QB.t1 3.15478
R12767 OR_magic_2.VOUT.t9 OR_magic_2.VOUT.t21 47.8944
R12768 OR_magic_2.VOUT.t17 OR_magic_2.VOUT.t3 47.8944
R12769 OR_magic_2.VOUT.t22 OR_magic_2.VOUT.t10 47.8944
R12770 OR_magic_2.VOUT.n0 OR_magic_2.VOUT.t6 47.3388
R12771 OR_magic_2.VOUT.n3 OR_magic_2.VOUT.t25 38.7949
R12772 OR_magic_2.VOUT.n2 OR_magic_2.VOUT.t24 38.7949
R12773 OR_magic_2.VOUT.n10 OR_magic_2.VOUT.t12 38.7949
R12774 OR_magic_2.VOUT.n11 OR_magic_2.VOUT.t5 38.7949
R12775 OR_magic_2.VOUT.n7 OR_magic_2.VOUT.t18 38.7949
R12776 OR_magic_2.VOUT.n6 OR_magic_2.VOUT.t13 38.7949
R12777 OR_magic_2.VOUT.n3 OR_magic_2.VOUT.n2 31.4949
R12778 OR_magic_2.VOUT.n11 OR_magic_2.VOUT.n10 31.4949
R12779 OR_magic_2.VOUT.n7 OR_magic_2.VOUT.n6 31.4949
R12780 divide_by_2_0.tg_magic_0.CLK OR_magic_2.VOUT.t20 31.3561
R12781 OR_magic_2.VOUT.n9 OR_magic_2.VOUT.t8 26.9781
R12782 OR_magic_2.VOUT.n9 OR_magic_2.VOUT.t14 26.9781
R12783 OR_magic_2.VOUT.n5 OR_magic_2.VOUT.t16 26.9781
R12784 OR_magic_2.VOUT.n5 OR_magic_2.VOUT.t26 26.9781
R12785 OR_magic_2.VOUT.n4 OR_magic_2.VOUT.t15 17.9416
R12786 OR_magic_2.VOUT.n12 OR_magic_2.VOUT.t11 17.9416
R12787 OR_magic_2.VOUT.n8 OR_magic_2.VOUT.t7 17.9416
R12788 OR_magic_2.VOUT.n0 divide_by_2_0.tg_magic_0.CLK 12.5623
R12789 OR_magic_2.VOUT.n4 OR_magic_2.VOUT.t9 11.957
R12790 OR_magic_2.VOUT.n12 OR_magic_2.VOUT.t17 11.957
R12791 OR_magic_2.VOUT.n8 OR_magic_2.VOUT.t22 11.957
R12792 OR_magic_2.VOUT.n0 OR_magic_2.VOUT.n8 10.9096
R12793 divide_by_2_0.inverter_magic_5.VIN OR_magic_2.VOUT.n0 10.5271
R12794 divide_by_2_0.tg_magic_0.CLK OR_magic_2.VOUT.n12 10.0013
R12795 divide_by_2_0.inverter_magic_5.VIN OR_magic_2.VOUT.n4 9.96162
R12796 OR_magic_2.VOUT.n2 OR_magic_2.VOUT.t4 7.3005
R12797 OR_magic_2.VOUT.t15 OR_magic_2.VOUT.n3 7.3005
R12798 OR_magic_2.VOUT.n10 OR_magic_2.VOUT.t23 7.3005
R12799 OR_magic_2.VOUT.t11 OR_magic_2.VOUT.n11 7.3005
R12800 OR_magic_2.VOUT.t20 OR_magic_2.VOUT.n9 7.3005
R12801 OR_magic_2.VOUT.n6 OR_magic_2.VOUT.t19 7.3005
R12802 OR_magic_2.VOUT.t7 OR_magic_2.VOUT.n7 7.3005
R12803 OR_magic_2.VOUT.t6 OR_magic_2.VOUT.n5 7.3005
R12804 OR_magic_2.VOUT.n1 OR_magic_2.VOUT.t2 5.47387
R12805 OR_magic_2.VOUT.n1 OR_magic_2.VOUT.t1 4.65398
R12806 OR_magic_2.VOUT.n1 OR_magic_2.VOUT.t0 4.2255
R12807 OR_magic_2.VOUT.n1 divide_by_2_0.inverter_magic_5.VIN 2.72976
R12808 OUT1.n8 OUT1.t2 5.47387
R12809 OUT1.n9 OUT1.t0 4.65398
R12810 OUT1.n7 OUT1.n0 4.5005
R12811 OUT1.n6 OUT1.n5 4.5005
R12812 OUT1.n7 OUT1.n6 4.5005
R12813 OUT1.n8 OUT1.t1 4.2255
R12814 OUT1 OUT1.n7 3.93486
R12815 OUT1.n4 OUT1.n1 2.25472
R12816 OUT1.n5 OUT1.n4 2.24764
R12817 OUT1.n3 OUT1.n2 2.24764
R12818 OUT1.n9 OUT1.n8 0.427022
R12819 OUT1 OUT1.n9 0.257096
R12820 OUT1.n5 OUT1.n3 0.014526
R12821 OUT1.n7 OUT1.n1 0.00800207
R12822 OUT1.n3 OUT1.n1 0.00800207
R12823 OUT1.n6 OUT1.n2 0.00772311
R12824 OUT1.n4 OUT1.n0 0.00772311
R12825 OUT1.n2 OUT1.n0 0.00772311
R12826 7b_counter_0.MDFF_5.QB.n1 7b_counter_0.MDFF_5.QB.t8 53.2571
R12827 7b_counter_0.MDFF_5.QB.n4 7b_counter_0.MDFF_5.QB.t5 38.8649
R12828 7b_counter_0.MDFF_5.QB.n3 7b_counter_0.MDFF_5.QB.t6 28.8568
R12829 7b_counter_0.MDFF_5.tspc2_magic_0.QB 7b_counter_0.MDFF_5.QB.n2 23.3781
R12830 7b_counter_0.MDFF_5.tspc2_magic_0.QB 7b_counter_0.MDFF_5.mux_magic_0.IN1 20.3676
R12831 7b_counter_0.MDFF_5.QB.n2 7b_counter_0.MDFF_5.QB.t7 17.1425
R12832 7b_counter_0.MDFF_5.QB.t5 7b_counter_0.MDFF_5.QB.n3 17.0773
R12833 7b_counter_0.MDFF_5.QB.n2 7b_counter_0.MDFF_5.QB.t4 14.405
R12834 7b_counter_0.MDFF_5.QB.n3 7b_counter_0.MDFF_5.QB.t2 11.6023
R12835 7b_counter_0.MDFF_5.mux_magic_0.IN1 7b_counter_0.MDFF_5.QB.n4 9.4273
R12836 7b_counter_0.MDFF_5.QB.n1 7b_counter_0.MDFF_5.QB.n0 8.57932
R12837 7b_counter_0.MDFF_5.QB.n4 7b_counter_0.MDFF_5.QB.t3 7.3005
R12838 7b_counter_0.MDFF_5.QB.t4 7b_counter_0.MDFF_5.QB.n1 7.3005
R12839 7b_counter_0.MDFF_5.QB.n0 7b_counter_0.MDFF_5.QB.t0 3.62007
R12840 7b_counter_0.MDFF_5.QB.n0 7b_counter_0.MDFF_5.QB.t1 3.15478
R12841 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t10 130.41
R12842 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n5 36.752
R12843 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t7 35.3186
R12844 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t4 33.5023
R12845 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t11 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n2 33.5023
R12846 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t5 32.2349
R12847 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n1 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n0 27.7405
R12848 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t3 26.3866
R12849 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t11 16.3786
R12850 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t3 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n1 13.2317
R12851 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n4 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n3 12.5023
R12852 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n3 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t9 11.3259
R12853 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n0 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t8 11.146
R12854 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n5 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t6 7.3005
R12855 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n2 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t12 7.3005
R12856 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n4 5.87653
R12857 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t2 5.47387
R12858 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t1 5.28011
R12859 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t0 4.65398
C0 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_7 0.028849f
C1 a_2749_10148# D2_7 2.25e-19
C2 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q3 4.44e-19
C3 a_15865_7470# Q1 3.82e-19
C4 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_12387_575# 1.37e-19
C5 a_1975_n1973# a_1541_n3597# 3.04e-19
C6 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A D2_6 0.060358f
C7 a_11279_1124# a_12387_575# 7.54e-20
C8 a_23258_575# a_23802_1059# 0.29829f
C9 a_26038_684# a_27234_575# 0.002003f
C10 a_9059_n1973# VDD 0.001798f
C11 a_8955_3363# Q5 3.88e-19
C12 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A Q6 0.023217f
C13 mux_magic_0.OR_magic_0.B mux_magic_0.IN2 0.002402f
C14 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n6024# 0.063645f
C15 a_15865_4557# a_15865_3363# 0.005574f
C16 a_1209_7469# VDD 0.807784f
C17 7b_counter_0.NAND_magic_0.VOUT CLK 0.678238f
C18 a_2749_3524# Q6 0.010505f
C19 Q1 D2_3 1.18919f
C20 a_4651_3947# a_5515_3947# 0.009722f
C21 a_23207_5885# Q6 2.99e-21
C22 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 0.003149f
C23 a_16065_9774# CLK 0.132735f
C24 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.LD 3.09e-20
C25 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C26 a_8523_n3150# D2_5 6.39e-20
C27 a_8523_n7648# a_8523_n8095# 0.014233f
C28 a_12174_n7648# p3_gen_magic_0.AND2_magic_1.A 0.09365f
C29 a_1409_4557# a_1409_3363# 0.020635f
C30 a_19152_6440# 7b_counter_0.MDFF_1.tspc2_magic_0.Q 0.001156f
C31 mux_magic_0.IN1 a_32816_n1264# 0.128819f
C32 a_8955_8580# VDD 0.085691f
C33 divide_by_2_1.tg_magic_3.IN VDD 2.62211f
C34 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8411_4513# 7.48e-20
C35 a_17405_2092# a_19152_739# 1.39e-20
C36 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 2.64e-19
C37 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_1209_1059# 1.63e-20
C38 7b_counter_0.MDFF_4.tspc2_magic_0.CLK p2_gen_magic_0.xnor_magic_3.OUT 2.45e-19
C39 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_17405_3524# 2.4e-20
C40 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VDD 1.23101f
C41 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B p2_gen_magic_0.xnor_magic_4.OUT 1e-19
C42 a_15865_9774# Q1 3.56e-19
C43 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VDD 1.25834f
C44 7b_counter_0.MDFF_5.tspc2_magic_0.CLK VDD 2.19889f
C45 a_2749_8740# a_4496_10093# 1.39e-20
C46 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.272186f
C47 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 0.00561f
C48 a_1559_n5540# D2_4 0.007723f
C49 a_18891_1669# CLK 0.004836f
C50 7b_counter_0.MDFF_4.LD a_19152_1223# 0.006779f
C51 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 6.94e-21
C52 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN Q4 0.008109f
C53 a_12387_575# VDD 0.91743f
C54 a_4496_4877# VDD 0.768234f
C55 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n1973# 0.009408f
C56 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_5 0.026134f
C57 a_1209_7469# LD 0.224216f
C58 7b_counter_0.MDFF_5.LD 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.015326f
C59 a_17405_2092# p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 6.42e-22
C60 p2_gen_magic_0.xnor_magic_3.OUT a_1559_n1526# 0.371619f
C61 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD 1.06874f
C62 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.001081f
C63 p3_gen_magic_0.xnor_magic_3.OUT a_1559_n6471# 0.09365f
C64 a_12387_5792# D2_6 3.05e-20
C65 p2_gen_magic_0.xnor_magic_1.OUT a_16186_n3644# 0.276806f
C66 a_2749_7308# Q7 0.010424f
C67 a_23985_7877# Q5 5.61e-19
C68 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.VOUT 3.5e-19
C69 p3_gen_magic_0.xnor_magic_4.OUT Q4 0.001267f
C70 7b_counter_0.NAND_magic_0.A 7b_counter_0.NAND_magic_0.VOUT 1.26949f
C71 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_5900# 0.189314f
C72 p2_gen_magic_0.3_inp_AND_magic_0.C D2_6 0.01833f
C73 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_20041_8580# 0.016967f
C74 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN Q4 0.00524f
C75 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_1209_1059# 1.93e-19
C76 a_1409_2253# a_1409_1059# 0.020635f
C77 a_27234_1769# a_27778_2253# 0.299584f
C78 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_1 5.14e-19
C79 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_2.IN 6.95e-19
C80 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A Q1 3.35e-19
C81 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_6 0.055831f
C82 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n5540# 0.090721f
C83 DFF_magic_0.tg_magic_0.IN CLK 0.628351f
C84 a_5470_n1973# Q2 2.48e-20
C85 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A LD 1.1e-20
C86 a_11191_684# D2_2 0.015291f
C87 a_2749_5900# CLK 0.00119f
C88 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.003149f
C89 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B Q1 0.007617f
C90 a_1559_n5540# Q2 0.014303f
C91 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B D2_2 0.003799f
C92 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.001131f
C93 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q6 0.003899f
C94 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.003851f
C95 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 4.02e-20
C96 a_11279_6341# CLK 0.0096f
C97 p2_gen_magic_0.xnor_magic_3.OUT VDD 2.87991f
C98 p2_gen_magic_0.3_inp_AND_magic_0.C a_13553_n2115# 0.001361f
C99 a_5036_n8095# D2_3 3.01e-19
C100 a_32616_n2458# a_32816_n2458# 0.299584f
C101 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.008196f
C102 p3_gen_magic_0.P3 a_23352_n5390# 0.191862f
C103 a_8523_n7648# Q1 0.008025f
C104 7b_counter_0.MDFF_3.QB Q2 2.58597f
C105 p2_gen_magic_0.xnor_magic_3.OUT D2_1 0.028169f
C106 a_23985_7877# D2_4 0.011147f
C107 a_12931_6276# CLK 0.00519f
C108 7b_counter_0.MDFF_4.LD a_15865_6276# 0.001019f
C109 a_34156_n2297# a_32616_n2458# 0.001529f
C110 a_21381_8741# Q2 5.13e-19
C111 a_15865_7470# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.001985f
C112 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_5185_1059# 1.93e-19
C113 7b_counter_0.NAND_magic_0.A 7b_counter_0.3_inp_AND_magic_0.B 0.001911f
C114 a_5385_7469# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 5.46e-20
C115 p2_gen_magic_0.3_inp_AND_magic_0.B a_16186_n3644# 0.04408f
C116 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 2.24e-19
C117 7b_counter_0.MDFF_4.LD a_19841_4557# 3.96e-19
C118 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_4 0.002731f
C119 p2_gen_magic_0.xnor_magic_1.OUT a_1957_n3150# 0.06406f
C120 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_6725_7308# 0.001347f
C121 p2_gen_magic_0.xnor_magic_3.OUT LD 2.3e-19
C122 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B 9.4e-20
C123 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A D2_3 0.014468f
C124 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.AND2_magic_1.A 0.257594f
C125 a_12387_1769# 7b_counter_0.MDFF_4.tspc2_magic_0.D 7.57e-20
C126 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.001415f
C127 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_17405_4932# 0.414018f
C128 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 0.008877f
C129 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_6725_2092# 0.036613f
C130 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_7 0.153151f
C131 p2_gen_magic_0.xnor_magic_0.OUT Q5 1.12e-19
C132 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.tspc2_magic_0.Q 0.121479f
C133 a_12387_5792# D2_2 0.012673f
C134 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 0.178114f
C135 a_23985_7877# Q2 4.81e-19
C136 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q5 2.57e-19
C137 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.B 3.82e-19
C138 a_1559_n1973# a_1541_n3597# 5.1e-19
C139 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q3 2.56e-19
C140 a_24059_4877# CLK 0.001181f
C141 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 8.78e-21
C142 a_8643_n1973# VDD 0.001396f
C143 a_11292_n6613# a_11708_n6613# 0.278913f
C144 a_5054_n1973# Q5 0.045953f
C145 a_16186_n3644# CLK 0.002493f
C146 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A CLK 0.074544f
C147 a_19841_3363# Q5 6.91e-20
C148 a_12387_575# Q3 2.12e-19
C149 a_1559_n6471# a_1541_n7648# 0.012783f
C150 a_24401_7877# VDD 0.021978f
C151 mux_magic_0.IN1 a_32816_n2458# 0.002005f
C152 a_2749_4932# Q6 0.016404f
C153 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 0.005939f
C154 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_17405_684# 3.58e-20
C155 a_22991_5885# Q6 2.81e-19
C156 a_5470_n6471# D2_4 0.005899f
C157 a_5515_9163# CLK 0.003088f
C158 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.xnor_magic_1.OUT 0.022718f
C159 p2_gen_magic_0.xnor_magic_0.OUT D2_4 0.0038f
C160 divide_by_2_0.tg_magic_0.IN VDD 0.995698f
C161 a_5452_n3150# D2_5 0.002782f
C162 p3_gen_magic_0.xnor_magic_6.OUT a_12590_n7648# 0.002939f
C163 a_19841_8580# VDD 0.921956f
C164 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_15865_2253# 5.28e-20
C165 a_18891_6886# 7b_counter_0.MDFF_1.tspc2_magic_0.Q 9.59e-20
C166 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 0.16497f
C167 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A D2_4 0.012116f
C168 a_23258_1769# VDD 0.937997f
C169 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.001313f
C170 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_22062_684# 0.414018f
C171 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_3524# 1e-20
C172 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_20041_9774# 0.128771f
C173 mux_magic_0.IN2 divide_by_2_0.tg_magic_3.IN 0.348508f
C174 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.001081f
C175 a_19841_8580# D2_1 0.243646f
C176 a_8955_4557# VDD 0.098457f
C177 a_17405_10149# VDD 1.55669f
C178 p2_gen_magic_0.xnor_magic_3.OUT Q3 1.2893f
C179 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5385_6275# 0.128771f
C180 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B VDD 1.19253f
C181 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11279_3480# 0.036613f
C182 7b_counter_0.MDFF_4.LD a_18891_1669# 1.61e-20
C183 7b_counter_0.MDFF_1.tspc2_magic_0.D p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.001257f
C184 a_17405_3524# a_15865_3363# 0.001529f
C185 a_1409_4557# VDD 0.05951f
C186 a_27778_2253# VDD 0.012214f
C187 a_23258_1769# a_23802_2253# 0.297401f
C188 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B CLK 0.01272f
C189 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q4 0.001319f
C190 a_8939_n7648# Q5 2.48e-20
C191 a_5470_n6471# Q2 2.48e-20
C192 a_17405_10149# D2_1 0.016115f
C193 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5470_n6471# 0.005701f
C194 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A D2_2 0.004052f
C195 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B D2_1 0.022439f
C196 p3_gen_magic_0.xnor_magic_1.OUT VDD 1.58618f
C197 p3_gen_magic_0.xnor_magic_3.OUT a_5054_n6024# 1.65e-19
C198 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 2.4e-20
C199 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q2 2.21e-19
C200 p2_gen_magic_0.xnor_magic_1.OUT a_14556_n3644# 0.021868f
C201 p2_gen_magic_0.3_inp_AND_magic_0.A D2_3 0.009584f
C202 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.3_inp_AND_magic_0.C 1.28495f
C203 p2_gen_magic_0.3_inp_AND_magic_0.A a_13353_n2115# 0.48198f
C204 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q5 5.26e-19
C205 a_1209_2253# a_1409_1059# 0.003083f
C206 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_0.IN 0.311939f
C207 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n3150# 0.107246f
C208 a_5185_7469# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 0.001985f
C209 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5036_n3150# 5.22e-19
C210 p3_gen_magic_0.xnor_magic_1.OUT D2_1 0.002381f
C211 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7 0.53521f
C212 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_4932# 1.52e-21
C213 a_2749_7308# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 1.01e-20
C214 a_17405_8741# Q1 0.043594f
C215 a_5054_n1973# Q2 0.305824f
C216 a_8955_8580# a_8713_6842# 5.39e-19
C217 7b_counter_0.MDFF_5.tspc2_magic_0.D 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 8.78e-21
C218 a_6725_7308# CLK 9.8e-20
C219 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B LD 6.07e-19
C220 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7215_10149# 0.414018f
C221 a_1409_4557# LD 0.003068f
C222 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A Q1 0.002402f
C223 a_16386_n8142# D2_6 0.010335f
C224 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_8411_9730# 1.93e-19
C225 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B Q6 0.053881f
C226 p3_gen_magic_0.3_inp_AND_magic_0.C D2_6 0.059955f
C227 a_5452_n3150# D2_7 0.007843f
C228 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8713_6842# 0.514308f
C229 DFF_magic_0.D a_30365_3514# 0.003744f
C230 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 3.55e-20
C231 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A D2_4 8.97e-19
C232 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.001139f
C233 a_12387_5792# CLK 0.016029f
C234 a_34156_n889# a_32616_n2458# 7.51e-20
C235 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A Q6 3.87e-19
C236 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 2.07e-19
C237 a_1559_n1526# p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 7.02e-19
C238 p2_gen_magic_0.3_inp_AND_magic_0.C CLK 0.670422f
C239 p2_gen_magic_0.3_inp_AND_magic_0.B a_14556_n3644# 0.146828f
C240 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n4081# 0.064529f
C241 p3_gen_magic_0.xnor_magic_3.OUT VDD 2.86103f
C242 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 0.043481f
C243 a_19152_6440# Q1 0.012641f
C244 7b_counter_0.NAND_magic_0.A 7b_counter_0.3_inp_AND_magic_0.VOUT 0.097055f
C245 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 0.178114f
C246 a_15865_6276# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 1.39e-19
C247 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 0.475387f
C248 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n4081# 0.092231f
C249 a_8713_1625# Q1 0.060197f
C250 a_24401_7877# Q3 7.62e-20
C251 a_9689_6886# a_9412_5956# 0.001643f
C252 a_1541_n3150# a_1957_n3150# 0.002223f
C253 p3_gen_magic_0.xnor_magic_3.OUT D2_1 1.58539f
C254 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.AND2_magic_1.A 3.88e-19
C255 a_5054_n6471# Q5 0.578984f
C256 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VDD 1.17128f
C257 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.18088f
C258 a_23258_1769# Q3 1.56e-19
C259 7b_counter_0.MDFF_4.LD a_8411_4513# 3.96e-19
C260 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD 1.03143f
C261 7b_counter_0.MDFF_5.LD 7b_counter_0.3_inp_AND_magic_0.A 7.88e-20
C262 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A Q5 6.14e-19
C263 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q2 3.98e-20
C264 a_5185_2253# Q5 0.00124f
C265 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 0.00112f
C266 a_9412_739# Q1 0.003124f
C267 a_2749_8740# 7b_counter_0.MDFF_3.tspc2_magic_0.D 0.134004f
C268 a_32816_n1264# VDD 0.056754f
C269 p3_gen_magic_0.xnor_magic_5.OUT D2_6 0.465654f
C270 DFF_magic_0.D a_27234_1769# 6.41e-19
C271 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_1 1.14674f
C272 7b_counter_0.MDFF_7.tspc2_magic_0.D 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B 0.001711f
C273 7b_counter_0.MDFF_1.tspc2_magic_0.D D2_3 0.003663f
C274 a_11292_n6613# a_11492_n6613# 0.522094f
C275 a_22150_1124# CLK 0.095912f
C276 a_8643_n1526# Q5 6.51e-20
C277 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.Q 8.23e-20
C278 a_14556_n3644# CLK 0.003888f
C279 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 8.54e-19
C280 7b_counter_0.MDFF_0.tspc2_magic_0.D VDD 1.451f
C281 a_21504_5904# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 3.96e-19
C282 a_27778_2253# Q3 0.002005f
C283 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 0.002118f
C284 a_24185_7877# VDD 0.020979f
C285 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.00222f
C286 p3_gen_magic_0.xnor_magic_0.OUT Q5 4.41e-20
C287 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B CLK 1.23e-19
C288 a_32816_n1264# D2_1 0.003068f
C289 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1 0.68028f
C290 7b_counter_0.MDFF_6.tspc2_magic_0.Q Q2 7.43e-19
C291 7b_counter_0.MDFF_3.tspc2_magic_0.Q Q7 0.100405f
C292 a_5054_n6471# D2_4 0.008877f
C293 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1541_n3597# 6.14e-19
C294 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19841_8580# 6.68e-20
C295 a_4651_9163# CLK 0.002867f
C296 a_9212_739# Q4 1.76e-20
C297 p3_gen_magic_0.xnor_magic_1.OUT Q3 1.22e-20
C298 a_26038_684# DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.9e-19
C299 a_5452_n7648# a_5036_n8095# 0.013021f
C300 a_7215_4932# a_8411_3319# 7.51e-20
C301 p2_gen_magic_0.AND2_magic_1.A VDD 1.36527f
C302 7b_counter_0.DFF_magic_0.tg_magic_3.OUT LD 0.018595f
C303 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.xnor_magic_6.OUT 0.039667f
C304 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A CLK 0.083594f
C305 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8411_3319# 0.001985f
C306 a_22150_1124# a_22062_684# 0.479729f
C307 a_17405_2092# a_15865_1059# 7.54e-20
C308 a_17405_7309# Q1 1.7e-19
C309 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.025041f
C310 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.099076f
C311 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 0.435114f
C312 p2_gen_magic_0.AND2_magic_1.A D2_1 1.92e-19
C313 a_1409_2253# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 0.001034f
C314 Q7 D2_5 0.831367f
C315 a_4496_4393# VDD 1.07616f
C316 a_27778_4557# D2_4 0.003998f
C317 a_19841_9774# VDD 0.902903f
C318 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 2.63e-19
C319 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5185_6275# 0.243646f
C320 7b_counter_0.MDFF_0.tspc2_magic_0.D LD 0.008524f
C321 a_1409_1059# CLK 0.003964f
C322 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_11191_4932# 0.414018f
C323 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.3_inp_AND_magic_0.C 0.235618f
C324 7b_counter_0.MDFF_5.LD D2_6 0.09231f
C325 a_7215_4932# VDD 1.55679f
C326 a_20171_1669# VDD 0.083906f
C327 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VDD 1.26056f
C328 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n6471# 0.00265f
C329 a_5054_n6471# Q2 0.305824f
C330 a_12387_4513# D2_2 0.012673f
C331 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_26038_684# 0.414018f
C332 a_1541_n7648# VDD 0.013993f
C333 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12931_1059# 0.037614f
C334 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A Q2 0.353472f
C335 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12387_3319# 0.001985f
C336 p3_gen_magic_0.xnor_magic_3.OUT a_1559_n6024# 0.371619f
C337 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8955_3363# 5.46e-20
C338 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_4496_9609# 0.012464f
C339 a_1209_7469# a_2749_5900# 7.51e-20
C340 DFF_magic_0.D P2 0.627139f
C341 a_1209_2253# a_1209_1059# 0.005574f
C342 p3_gen_magic_0.xnor_magic_3.OUT Q3 0.148989f
C343 a_5054_n1973# a_5470_n1973# 5.82e-19
C344 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_2.IN 0.973398f
C345 a_12931_9774# Q1 0.128771f
C346 a_4496_4393# LD 0.00664f
C347 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VDD 1.23245f
C348 a_19841_9774# LD 4.93e-19
C349 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9412_5956# 0.120019f
C350 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1541_n7648# 9.19e-19
C351 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q6 0.212702f
C352 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT 1.75e-19
C353 a_15865_7470# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.001158f
C354 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.09061f
C355 a_14756_n8142# D2_6 0.013925f
C356 p3_gen_magic_0.3_inp_AND_magic_0.A D2_3 0.01949f
C357 DFF_magic_0.D a_30365_4922# 0.016244f
C358 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_11279_6341# 0.009039f
C359 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 2.83e-20
C360 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT D2_1 0.007318f
C361 7b_counter_0.MDFF_4.LD a_12387_5792# 0.001019f
C362 a_12387_9730# Q6 3.01e-19
C363 a_9212_739# p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 4.12e-20
C364 7b_counter_0.MDFF_4.LD p2_gen_magic_0.3_inp_AND_magic_0.C 9.4e-19
C365 a_8523_n3597# D2_6 0.238982f
C366 D2_7 Q7 0.777755f
C367 a_18891_6886# Q1 0.002472f
C368 a_6725_684# VDD 1.55925f
C369 7b_counter_0.MDFF_5.LD a_11279_8697# 0.001152f
C370 7b_counter_0.MDFF_4.tspc2_magic_0.D D2_3 5.71e-19
C371 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.VOUT 3.5e-19
C372 a_24185_7877# Q3 1.32e-19
C373 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8523_n8095# 1.63e-19
C374 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.xnor_magic_5.OUT 5.78e-19
C375 7b_counter_0.MDFF_5.LD D2_2 0.535811f
C376 a_32616_n1264# a_32816_n1264# 0.29829f
C377 DFF_magic_0.D VDD 8.66413f
C378 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.08338f
C379 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n7648# 0.009154f
C380 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_5 0.091602f
C381 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_19841_8580# 0.001158f
C382 a_8643_n6024# Q5 6.51e-20
C383 7b_counter_0.MDFF_5.tspc2_magic_0.Q 7b_counter_0.MDFF_5.LD 0.121479f
C384 a_27778_3363# CLK 0.002092f
C385 p3_gen_magic_0.3_inp_AND_magic_0.C CLK 0.686729f
C386 a_32816_n2458# VDD 0.012214f
C387 a_11279_3480# Q5 0.032844f
C388 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 5.04e-22
C389 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 0.00112f
C390 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT D2_1 0.001243f
C391 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_7309# 0.036613f
C392 a_2749_10148# 7b_counter_0.MDFF_3.tspc2_magic_0.D 1.08e-19
C393 7b_counter_0.MDFF_4.LD a_20041_4557# 1.1e-19
C394 7b_counter_0.DFF_magic_0.tg_magic_0.IN D2_4 0.00268f
C395 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A Q5 0.002209f
C396 a_32816_n2458# D2_1 0.040868f
C397 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8955_4557# 0.128771f
C398 p3_gen_magic_0.xnor_magic_6.OUT D2_5 0.134516f
C399 a_34156_n2297# VDD 0.938506f
C400 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 9.4e-20
C401 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VDD 1.25061f
C402 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A CLK 0.001266f
C403 p2_gen_magic_0.AND2_magic_1.A a_16386_n3644# 3.84e-19
C404 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B CLK 0.012705f
C405 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8411_4513# 2.09e-19
C406 a_1541_n3597# a_1541_n4081# 0.033537f
C407 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_3.OUT 6.9e-21
C408 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 1.64e-19
C409 a_17405_2092# CLK 2.46e-19
C410 a_2749_3524# VDD 0.954212f
C411 mux_magic_0.OR_magic_0.B a_32616_n2458# 0.146237f
C412 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_5385_2253# 0.007492f
C413 a_23207_5885# VDD 0.164609f
C414 a_1559_n6024# a_1541_n7648# 0.001207f
C415 a_4496_9609# D2_7 5.51e-20
C416 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_9212_739# 7.16e-19
C417 a_5054_n1042# Q1 8.14e-20
C418 DFF_magic_0.D LD 0.477933f
C419 p3_gen_magic_0.xnor_magic_1.OUT a_8523_n8579# 0.010037f
C420 a_1541_n7648# Q3 1.88e-19
C421 a_1541_n3597# VDD 0.183944f
C422 a_12387_4513# CLK 0.016029f
C423 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 0.445675f
C424 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 5.37e-19
C425 a_21381_4932# Q4 0.003039f
C426 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.OUT 0.224325f
C427 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A D2_4 0.023258f
C428 a_1209_2253# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 0.001158f
C429 a_1541_n3597# D2_1 0.239111f
C430 a_8523_n3597# D2_2 3.13e-19
C431 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1409_6275# 0.037614f
C432 Q6 Q5 0.353381f
C433 7b_counter_0.3_inp_AND_magic_0.B a_24401_7877# 0.062631f
C434 a_15865_4557# VDD 0.944161f
C435 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.00112f
C436 a_1975_n1973# D2_4 0.005701f
C437 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A LD 1.1e-20
C438 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q1 0.655594f
C439 a_19307_1669# VDD 0.003613f
C440 a_12931_4557# a_12387_3319# 0.003083f
C441 OR_magic_2.A divide_by_2_0.tg_magic_3.IN 0.001359f
C442 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B D2_5 0.007521f
C443 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7 1.18088f
C444 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 0.27167f
C445 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_12387_575# 0.279825f
C446 a_26126_1124# a_26038_684# 0.479729f
C447 a_6725_2092# a_6725_684# 0.479729f
C448 p2_gen_magic_0.xnor_magic_5.OUT p2_gen_magic_0.AND2_magic_1.A 0.424155f
C449 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_1209_8579# 5.28e-20
C450 a_4235_9163# a_4496_9609# 0.301553f
C451 D2_5 D2_3 3.47391f
C452 a_13353_n2115# D2_5 4.86e-20
C453 a_19152_1223# a_20171_1669# 0.043767f
C454 a_11191_684# a_12387_575# 0.002003f
C455 mux_magic_0.IN1 mux_magic_0.OR_magic_0.B 1.06e-19
C456 OR_magic_2.A OR_magic_1.VOUT 0.058198f
C457 p3_gen_magic_0.xnor_magic_6.OUT D2_7 0.001806f
C458 Q6 D2_4 1.66999f
C459 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VDD 1.26783f
C460 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_18891_6886# 3.22e-21
C461 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.008597f
C462 a_1209_3363# Q6 0.00186f
C463 7b_counter_0.MDFF_5.LD CLK 0.959252f
C464 DFF_magic_0.D Q3 0.320053f
C465 a_16186_n8142# D2_6 0.018747f
C466 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK Q4 0.011368f
C467 a_11292_n2115# D2_2 0.036571f
C468 a_15865_7470# 7b_counter_0.MDFF_6.tspc2_magic_0.D 7.57e-20
C469 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C470 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN CLK 0.612651f
C471 a_23793_5904# Q5 0.543517f
C472 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.12089f
C473 Q2 Q6 1.37834f
C474 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q6 0.016176f
C475 p3_gen_magic_0.3_inp_AND_magic_0.B a_16386_n8142# 6.81e-19
C476 7b_counter_0.MDFF_5.LD a_11191_10149# 0.002672f
C477 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.3_inp_AND_magic_0.C 1.28709f
C478 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.854418f
C479 p3_gen_magic_0.3_inp_AND_magic_0.A a_13353_n6613# 0.48198f
C480 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_12387_5792# 1.37e-19
C481 a_23207_5885# Q3 0.205896f
C482 mux_magic_0.AND2_magic_0.A a_32816_n1264# 0.037583f
C483 a_32616_n1264# a_34156_n2297# 7.54e-20
C484 7b_counter_0.MDFF_6.tspc2_magic_0.D D2_3 0.09871f
C485 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1541_n3150# 4.77e-19
C486 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C487 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5452_n3150# 0.005701f
C488 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.0037f
C489 p2_gen_magic_0.xnor_magic_6.OUT Q4 0.385788f
C490 a_1409_8579# VDD 0.012214f
C491 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q4 1.64e-19
C492 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n8095# 0.063777f
C493 a_20041_3363# CLK 3.99e-19
C494 7b_counter_0.MDFF_4.LD a_27778_3363# 0.037786f
C495 p3_gen_magic_0.xnor_magic_0.OUT a_12174_n7648# 0.001986f
C496 a_8411_9730# 7b_counter_0.MDFF_5.LD 3.96e-19
C497 a_15865_4557# a_17405_4932# 0.002003f
C498 a_1541_n3597# Q3 6.69e-21
C499 a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 1.93e-19
C500 D2_7 D2_3 0.012129f
C501 a_27234_4513# 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.279825f
C502 7b_counter_0.NAND_magic_0.A 7b_counter_0.MDFF_5.LD 0.168841f
C503 DFF_magic_0.D 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 2.35e-19
C504 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_19841_9774# 0.279825f
C505 a_2749_10148# a_2749_8740# 0.479729f
C506 a_23793_5904# D2_4 0.006832f
C507 a_8411_4513# a_8955_4557# 0.29829f
C508 a_8523_n7648# D2_5 0.013609f
C509 a_34156_n889# VDD 1.55668f
C510 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 1.1e-20
C511 a_2749_4932# VDD 1.55786f
C512 a_8643_n6471# p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.001598f
C513 7b_counter_0.MDFF_7.tspc2_magic_0.D D2_4 0.087353f
C514 p2_gen_magic_0.AND2_magic_1.A a_14756_n3644# 0.037687f
C515 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 2.36e-19
C516 a_12387_3319# Q5 0.043281f
C517 a_23258_1769# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 0.001985f
C518 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_2749_2092# 0.132169f
C519 a_23560_3728# Q5 7.87e-19
C520 a_1541_n8095# Q6 1.35e-19
C521 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A D2_7 0.013653f
C522 a_22991_5885# VDD 1.07263f
C523 7b_counter_0.MDFF_1.tspc2_magic_0.CLK D2_3 0.069738f
C524 a_8523_n4081# Q5 1.41e-19
C525 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A CLK 0.011567f
C526 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1409_8579# 7.81e-19
C527 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_4.tspc2_magic_0.Q 0.002402f
C528 a_1409_8579# LD 0.037687f
C529 a_1975_n6471# D2_4 0.005701f
C530 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.3_inp_AND_magic_0.C 0.008265f
C531 a_11292_n2115# p2_gen_magic_0.3_inp_AND_magic_0.B 0.002342f
C532 p2_gen_magic_0.xnor_magic_4.OUT D2_3 0.165551f
C533 a_12174_n3150# VDD 0.001396f
C534 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.xnor_magic_5.OUT 0.048563f
C535 7b_counter_0.MDFF_4.LD a_12387_4513# 0.002086f
C536 a_5054_n6471# a_5470_n6471# 5.82e-19
C537 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n7648# 0.107246f
C538 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1209_6275# 0.279825f
C539 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B Q4 0.001088f
C540 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q3 0.003764f
C541 7b_counter_0.3_inp_AND_magic_0.B a_24185_7877# 0.123074f
C542 a_1559_n1973# D2_4 0.101104f
C543 a_11292_n2115# a_11708_n2115# 0.278913f
C544 p3_gen_magic_0.3_inp_AND_magic_0.A a_13769_n6613# 0.02473f
C545 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_2092# 0.431521f
C546 a_5054_n5540# Q1 5.54e-20
C547 a_23560_3728# D2_4 0.019531f
C548 7b_counter_0.3_inp_AND_magic_0.VOUT a_24401_7877# 0.200301f
C549 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n1526# 0.082315f
C550 a_1209_6275# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 1.39e-19
C551 a_17405_684# VDD 1.55668f
C552 OR_magic_2.A a_23352_n6798# 0.036613f
C553 p2_gen_magic_0.xnor_magic_0.OUT a_8643_n1526# 0.417891f
C554 mux_magic_0.OR_magic_0.A a_32616_n2458# 0.001985f
C555 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_6 0.081414f
C556 7b_counter_0.MDFF_7.tspc2_magic_0.CLK CLK 0.042625f
C557 a_1975_n6471# Q2 7.44e-19
C558 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_5.tspc2_magic_0.D 0.001711f
C559 p2_gen_magic_0.xnor_magic_1.OUT a_5036_n3597# 1.79e-22
C560 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n1042# 0.063097f
C561 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B VDD 1.20888f
C562 a_4496_10093# a_4496_9609# 0.014143f
C563 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VDD 1.2392f
C564 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VDD 1.24206f
C565 a_19152_1223# a_19307_1669# 0.240883f
C566 a_18891_1669# a_20171_1669# 0.007202f
C567 7b_counter_0.MDFF_4.tspc2_magic_0.D a_8713_1625# 0.037942f
C568 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.006771f
C569 a_17405_3524# VDD 0.941683f
C570 divide_by_2_0.tg_magic_1.IN VDD 1.85417f
C571 p3_gen_magic_0.P3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 0.314216f
C572 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A D2_1 0.005423f
C573 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B VDD 1.19433f
C574 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.001777f
C575 a_7303_8697# CLK 0.016426f
C576 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_4.LD 0.035182f
C577 a_14556_n8142# D2_6 0.065394f
C578 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VDD 1.25655f
C579 a_8643_n1973# p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.81e-19
C580 a_8825_6886# Q7 0.002019f
C581 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9412_739# 0.120019f
C582 a_13353_n6613# D2_5 0.025567f
C583 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B D2_1 0.002402f
C584 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VDD 1.31149f
C585 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN 0.340787f
C586 a_1975_n6471# a_1541_n8095# 3.04e-19
C587 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 0.001081f
C588 a_8713_1625# a_9689_1669# 0.240883f
C589 mux_magic_0.AND2_magic_0.A a_32816_n2458# 0.001034f
C590 a_5470_n1973# Q6 8.88e-19
C591 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A LD 5.6e-19
C592 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A D2_1 3.54e-19
C593 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.OUT 2.58e-20
C594 p3_gen_magic_0.3_inp_AND_magic_0.B a_14756_n8142# 0.007767f
C595 7b_counter_0.NAND_magic_0.VOUT DFF_magic_0.D 0.00552f
C596 a_15865_6276# a_15865_4557# 0.005698f
C597 a_5185_2253# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 0.001158f
C598 a_22991_5885# Q3 0.032029f
C599 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.08438f
C600 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A D2_3 0.196349f
C601 mux_magic_0.AND2_magic_0.A a_34156_n2297# 2.4e-20
C602 a_32616_n1264# a_34156_n889# 0.002003f
C603 a_17405_7309# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 2.4e-20
C604 mux_magic_0.IN1 mux_magic_0.OR_magic_0.A 0.002509f
C605 OR_magic_1.VOUT mux_magic_0.IN1 0.006372f
C606 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B LD 6.96e-19
C607 a_1209_4557# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 1.37e-19
C608 7b_counter_0.MDFF_3.QB Q6 0.12363f
C609 a_8411_8536# VDD 0.921905f
C610 a_11292_n6613# D2_2 0.002579f
C611 a_9689_1669# a_9412_739# 0.001643f
C612 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A Q5 0.002247f
C613 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD 1.18294f
C614 a_8411_9730# a_7303_8697# 7.54e-20
C615 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.030838f
C616 p3_gen_magic_0.xnor_magic_0.OUT a_8939_n7648# 1.73e-19
C617 7b_counter_0.MDFF_4.LD a_20041_3363# 0.036926f
C618 a_27234_3319# CLK 0.007722f
C619 a_1559_n6471# Q5 0.582233f
C620 a_5515_3947# Q7 0.005231f
C621 a_21381_8741# Q6 0.15441f
C622 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT a_23352_n6798# 1.08e-20
C623 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A LD 6.12e-19
C624 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_1 4.07e-19
C625 a_6725_5900# 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B 4.85e-19
C626 p2_gen_magic_0.xnor_magic_1.OUT a_11292_n6613# 1.35e-19
C627 a_5054_n1526# Q5 0.008164f
C628 a_23258_1769# a_22150_1124# 0.001529f
C629 a_20041_8580# VDD 0.085691f
C630 a_8411_4513# a_7215_4932# 0.002003f
C631 a_5036_n4081# Q5 1.88e-19
C632 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8411_4513# 0.149276f
C633 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A D2_4 0.020305f
C634 a_1559_n6471# D2_4 0.057124f
C635 p3_gen_magic_0.xnor_magic_1.OUT a_1541_n8579# 0.340948f
C636 7b_counter_0.MDFF_7.tspc2_magic_0.Q 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.267492f
C637 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN 0.973393f
C638 a_17405_4932# a_17405_3524# 0.479729f
C639 a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 0.149276f
C640 a_20041_8580# D2_1 0.128625f
C641 a_8939_n3150# VDD 0.001798f
C642 a_15865_8580# VDD 0.821356f
C643 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1957_n3150# 6.1e-19
C644 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_3524# 0.431521f
C645 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B Q4 5.49e-19
C646 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q5 7.7e-19
C647 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A Q3 1.93e-19
C648 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 3.69e-19
C649 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 4e-20
C650 a_15865_8580# D2_1 0.002785f
C651 7b_counter_0.3_inp_AND_magic_0.B a_23207_5885# 0.047377f
C652 a_9059_n6471# a_8523_n8095# 1.25e-19
C653 a_23258_575# Q4 5.48e-20
C654 p3_gen_magic_0.3_inp_AND_magic_0.A a_13553_n6613# 0.075783f
C655 a_11292_n2115# a_11492_n2115# 0.522094f
C656 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26126_3480# 0.431521f
C657 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 1.09743f
C658 7b_counter_0.3_inp_AND_magic_0.VOUT a_24185_7877# 1.9e-20
C659 p3_gen_magic_0.xnor_magic_4.OUT D2_3 0.178008f
C660 a_1209_6275# a_1209_4557# 0.005708f
C661 mux_magic_0.OR_magic_0.B VDD 1.18037f
C662 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_11279_3480# 2.07e-19
C663 a_1209_3363# a_1409_3363# 0.299584f
C664 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 0.084688f
C665 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT 1.98e-19
C666 a_21381_3524# CLK 0.003249f
C667 a_1559_n6471# Q2 5.68e-19
C668 OR_magic_2.A mux_magic_0.IN2 0.010823f
C669 a_12931_7470# Q2 0.072957f
C670 a_8523_n3150# p2_gen_magic_0.xnor_magic_6.OUT 0.09365f
C671 p2_gen_magic_0.xnor_magic_3.OUT a_12174_n3597# 2.99e-20
C672 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4 1.2134f
C673 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8523_n3150# 3.55e-19
C674 a_1209_9773# VDD 0.91502f
C675 a_18891_1669# a_19307_1669# 0.16113f
C676 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8955_9774# 9.27e-19
C677 a_30365_3514# OR_magic_1.VOUT 0.137791f
C678 7b_counter_0.MDFF_6.tspc2_magic_0.D a_19152_6440# 0.036963f
C679 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n1042# 0.093592f
C680 a_5452_n7648# D2_7 0.006494f
C681 a_12931_4557# VDD 0.059235f
C682 a_5054_n1526# Q2 0.08832f
C683 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD 1.50347f
C684 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.02429f
C685 a_1209_9773# D2_1 0.009386f
C686 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT D2_6 0.001989f
C687 a_5036_n4081# p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 1.66e-20
C688 a_5470_n6471# Q6 0.001991f
C689 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 0.00112f
C690 7b_counter_0.MDFF_5.LD a_8955_8580# 0.036926f
C691 a_6725_5900# Q7 0.015269f
C692 p2_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 2.73e-19
C693 a_27234_1769# D2_4 0.01192f
C694 a_12387_9730# VDD 0.915238f
C695 a_1559_n6471# a_1541_n8095# 5.02e-19
C696 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A Q6 8.78e-21
C697 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q2 0.023012f
C698 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1209_9773# 0.279393f
C699 a_8713_1625# a_8825_1669# 0.043767f
C700 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_1209_6275# 1.63e-20
C701 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.AND2_magic_1.A 0.004277f
C702 a_5054_n1973# Q6 0.008976f
C703 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 0.084688f
C704 a_1209_1059# p2_gen_magic_0.xnor_magic_3.OUT 1.9e-19
C705 a_1209_9773# LD 8.88e-19
C706 a_12387_9730# D2_1 2.73e-19
C707 a_9059_n6471# Q1 6.09e-19
C708 p3_gen_magic_0.3_inp_AND_magic_0.B a_16186_n8142# 0.04408f
C709 mux_magic_0.AND2_magic_0.A a_34156_n889# 3.58e-20
C710 a_6725_5900# a_5185_6275# 0.002003f
C711 a_20041_9774# VDD 0.087905f
C712 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 0.252991f
C713 7b_counter_0.MDFF_4.tspc2_magic_0.CLK Q5 0.306933f
C714 a_9059_n1973# a_8523_n3597# 1.25e-19
C715 a_11279_1124# Q5 5.93e-19
C716 a_4651_3947# Q7 0.003587f
C717 a_24536_3947# CLK 1.38e-20
C718 7b_counter_0.MDFF_4.LD a_27234_3319# 0.224216f
C719 a_9212_5956# a_9689_6886# 0.16113f
C720 a_17405_7309# 7b_counter_0.MDFF_6.tspc2_magic_0.D 0.134004f
C721 DFF_magic_0.tg_magic_2.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.270406f
C722 a_12387_9730# LD 4.93e-19
C723 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.007492f
C724 DFF_magic_0.tg_magic_3.OUT CLK 0.458019f
C725 p3_gen_magic_0.AND2_magic_1.A VDD 1.36853f
C726 p2_gen_magic_0.AND2_magic_1.A a_14556_n3644# 0.232114f
C727 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 0.006183f
C728 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_20041_8580# 0.007392f
C729 OR_magic_2.A DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.001277f
C730 a_8411_3319# Q5 7.41e-19
C731 a_16065_8580# VDD 0.017121f
C732 a_2749_684# D2_4 0.008711f
C733 7b_counter_0.3_inp_AND_magic_0.VOUT DFF_magic_0.D 2.51e-20
C734 7b_counter_0.MDFF_4.tspc2_magic_0.CLK D2_4 0.001262f
C735 a_7215_10149# Q7 0.026618f
C736 a_11279_1124# D2_4 0.008528f
C737 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A Q7 0.024842f
C738 a_13553_n6613# D2_5 0.004092f
C739 a_5054_n6024# D2_4 0.10441f
C740 a_21381_10149# a_19841_8580# 7.51e-20
C741 p3_gen_magic_0.xnor_magic_1.OUT a_16386_n8142# 0.140317f
C742 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q6 0.042685f
C743 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.015506f
C744 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_15865_8580# 1.18e-19
C745 a_32616_n1264# mux_magic_0.OR_magic_0.B 1.93e-19
C746 a_12387_8536# VDD 0.808402f
C747 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.167732f
C748 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.xnor_magic_1.OUT 0.018814f
C749 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4496_9609# 0.038362f
C750 a_22150_1124# a_20171_1669# 1.2e-20
C751 VDD Q5 20.6027f
C752 a_8411_8536# a_8713_6842# 3.03e-19
C753 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q3 0.001141f
C754 7b_counter_0.3_inp_AND_magic_0.B a_22991_5885# 0.036617f
C755 p3_gen_magic_0.3_inp_AND_magic_0.A a_11708_n6613# 0.200301f
C756 7b_counter_0.MDFF_3.QB a_5185_7469# 2.1e-19
C757 OR_magic_1.VOUT P2 0.014566f
C758 a_1559_n1526# D2_4 0.238982f
C759 mux_magic_0.IN2 a_32616_n2458# 0.243646f
C760 a_8643_n6471# a_8523_n8095# 3.68e-19
C761 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_24259_4877# 1.29e-19
C762 7b_counter_0.MDFF_6.tspc2_magic_0.Q Q6 0.197372f
C763 a_1209_2253# a_2749_2092# 0.001529f
C764 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5385_2253# 0.016967f
C765 a_5385_1059# D2_5 0.00754f
C766 D2_1 Q5 0.430153f
C767 a_1559_n1042# a_1559_n1526# 0.033537f
C768 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.96823f
C769 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n6024# 0.076813f
C770 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_15865_3363# 0.001158f
C771 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q5 0.002112f
C772 a_5054_n6024# Q2 0.08832f
C773 p3_gen_magic_0.xnor_magic_0.OUT a_8643_n6024# 0.417891f
C774 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_6725_7308# 0.036613f
C775 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.226055f
C776 a_12387_6986# 7b_counter_0.MDFF_5.tspc2_magic_0.D 7.57e-20
C777 a_1957_n3150# a_1541_n3597# 0.013021f
C778 VDD D2_4 7.56276f
C779 a_5054_n1526# a_5470_n1973# 0.011514f
C780 a_19152_6440# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 6.92e-19
C781 a_5054_n1042# D2_5 0.050765f
C782 LD Q5 0.135035f
C783 7b_counter_0.MDFF_6.tspc2_magic_0.D a_18891_6886# 0.282223f
C784 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 1.75e-19
C785 a_11292_n6613# p3_gen_magic_0.3_inp_AND_magic_0.B 0.002342f
C786 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.3_inp_AND_magic_0.C 0.008265f
C787 a_1559_n1042# VDD 0.428164f
C788 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5036_n7648# 5.22e-19
C789 a_1209_3363# VDD 0.807784f
C790 divide_by_2_0.tg_magic_3.IN VDD 2.32307f
C791 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_5.OUT 1.3524f
C792 D2_1 D2_4 0.772998f
C793 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A Q1 0.002736f
C794 a_5054_n6471# Q6 0.034129f
C795 a_1541_n4081# Q2 0.002712f
C796 a_8523_n8095# D2_6 0.247611f
C797 7b_counter_0.MDFF_5.LD a_19841_8580# 0.224142f
C798 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_18891_1669# 3.22e-21
C799 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_4 1.02589f
C800 a_23802_2253# D2_4 0.128625f
C801 divide_by_2_0.tg_magic_3.IN D2_1 1.18541f
C802 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT Q4 0.020027f
C803 a_5185_2253# Q6 0.001407f
C804 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9212_5956# 0.281948f
C805 OR_magic_1.VOUT VDD 7.8931f
C806 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_5 0.105932f
C807 mux_magic_0.OR_magic_0.A VDD 1.23982f
C808 7b_counter_0.3_inp_AND_magic_0.A Q1 9.16e-20
C809 VDD Q2 9.58279f
C810 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VDD 1.36642f
C811 7b_counter_0.MDFF_5.LD a_17405_10149# 0.033168f
C812 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_5 0.004491f
C813 p3_gen_magic_0.AND2_magic_1.A a_12174_n8579# 0.616639f
C814 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 0.03034f
C815 LD D2_4 0.11201f
C816 mux_magic_0.IN1 mux_magic_0.IN2 0.003895f
C817 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 2.8e-19
C818 7b_counter_0.3_inp_AND_magic_0.C Q4 0.070001f
C819 p3_gen_magic_0.3_inp_AND_magic_0.B a_14556_n8142# 0.146828f
C820 a_8643_n6471# Q1 0.306431f
C821 7b_counter_0.MDFF_1.tspc2_magic_0.Q CLK 0.246829f
C822 mux_magic_0.OR_magic_0.A D2_1 1.1e-20
C823 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_20041_8580# 5.46e-20
C824 a_1209_3363# LD 0.224216f
C825 a_17405_5901# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 1.51e-21
C826 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT 9.88e-19
C827 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_1 7.64e-19
C828 Q2 D2_1 1.21457f
C829 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C830 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n5540# 0.063097f
C831 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6 1.17747f
C832 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK 2.41e-19
C833 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A CLK 0.022918f
C834 a_24003_10051# VDD 0.036385f
C835 p2_gen_magic_0.xnor_magic_3.OUT a_11292_n2115# 0.473167f
C836 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 4.28e-19
C837 a_23672_3947# CLK 1.93e-20
C838 a_6725_2092# Q5 0.166603f
C839 a_21381_4932# Q7 0.002782f
C840 a_8643_n1973# a_8523_n3597# 3.68e-19
C841 p3_gen_magic_0.xnor_magic_4.OUT a_5452_n7648# 7.38e-19
C842 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q2 0.058324f
C843 a_1559_n6024# Q5 7.45e-19
C844 p2_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.3_inp_AND_magic_0.C 4.5e-19
C845 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_1.IN 0.340787f
C846 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_6725_5900# 3.58e-20
C847 a_9212_5956# a_8825_6886# 0.007202f
C848 Q7 Q4 0.045256f
C849 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A Q2 0.112612f
C850 Q3 Q5 1.45629f
C851 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_3.OUT 0.001138f
C852 LD Q2 11.240499f
C853 a_1541_n8095# VDD 0.183131f
C854 p2_gen_magic_0.AND2_magic_1.A a_12174_n3597# 0.371679f
C855 a_12931_8580# VDD 0.012214f
C856 Q1 D2_6 0.897757f
C857 a_8523_n8095# D2_2 3.13e-19
C858 a_6725_2092# D2_4 0.00548f
C859 a_11708_n6613# D2_5 0.018884f
C860 a_1559_n6024# D2_4 0.247128f
C861 a_24003_10051# LD 0.023983f
C862 a_16065_9774# a_15865_8580# 0.003083f
C863 p3_gen_magic_0.xnor_magic_1.OUT a_14756_n8142# 1.75e-19
C864 p2_gen_magic_0.3_inp_AND_magic_0.VOUT Q4 0.139242f
C865 p2_gen_magic_0.xnor_magic_4.OUT a_5054_n1042# 0.299642f
C866 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1541_n8095# 5.59e-19
C867 a_15865_2253# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 0.146237f
C868 a_2749_8740# a_4496_9609# 7.92e-19
C869 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.AND2_magic_1.A 0.2354f
C870 7b_counter_0.MDFF_5.tspc2_magic_0.Q 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B 4.47e-20
C871 Q3 D2_4 2.85514f
C872 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_7 1.0525f
C873 a_12387_1769# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 0.146237f
C874 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 0.178114f
C875 a_19841_9774# a_21381_10149# 0.002003f
C876 a_1559_n1042# Q3 0.001176f
C877 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B D2_6 0.009023f
C878 p3_gen_magic_0.3_inp_AND_magic_0.A a_11492_n6613# 1.9e-20
C879 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_24059_4877# 7.16e-19
C880 a_26126_3480# D2_4 0.085237f
C881 a_2749_7308# a_1209_6275# 7.54e-20
C882 a_26038_684# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 3.58e-20
C883 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23802_1059# 0.037614f
C884 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8955_3363# 0.007492f
C885 a_5185_1059# D2_5 0.0193f
C886 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_2749_2092# 0.001371f
C887 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_2 0.011361f
C888 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_20041_4557# 9.27e-19
C889 a_1209_8579# D2_7 0.4436f
C890 a_1559_n6024# Q2 0.004225f
C891 a_19152_1223# Q5 8.58e-19
C892 OR_magic_2.A DFF_magic_0.tg_magic_2.IN 0.329918f
C893 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_23258_1769# 4.65e-19
C894 Q2 Q3 2.42882f
C895 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 0.178114f
C896 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT Q4 0.023826f
C897 7b_counter_0.MDFF_1.tspc2_magic_0.D a_19152_739# 0.120019f
C898 OR_magic_1.VOUT a_32616_n1264# 4.71e-19
C899 a_18891_6886# 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 5.62e-20
C900 a_32616_n1264# mux_magic_0.OR_magic_0.A 0.149276f
C901 a_5054_n1526# a_5054_n1973# 0.013665f
C902 p2_gen_magic_0.xnor_magic_5.OUT Q5 0.032187f
C903 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.001317f
C904 a_8411_3319# a_8955_3363# 0.297401f
C905 a_23352_n6798# VDD 0.990428f
C906 a_7303_3480# a_5515_3947# 2.9e-20
C907 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B p2_gen_magic_0.xnor_magic_3.OUT 1.55e-19
C908 p2_gen_magic_0.3_inp_AND_magic_0.A a_13769_n2115# 0.02473f
C909 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_20041_9774# 0.037614f
C910 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 4.61e-20
C911 DFF_magic_0.D a_27778_3363# 0.002281f
C912 Q1 D2_2 0.723103f
C913 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B D2_4 0.00379f
C914 a_23352_n6798# D2_1 0.024287f
C915 a_19152_1223# D2_4 0.042867f
C916 a_8955_3363# VDD 0.085691f
C917 OR_magic_1.VOUT divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 2.41e-19
C918 a_5470_n1973# VDD 0.003971f
C919 a_5054_n5540# D2_5 0.038932f
C920 p3_gen_magic_0.xnor_magic_6.OUT Q4 0.22793f
C921 a_1559_n5540# VDD 0.427807f
C922 7b_counter_0.MDFF_5.LD a_19841_9774# 0.00185f
C923 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11279_8697# 0.431521f
C924 p2_gen_magic_0.xnor_magic_5.OUT D2_4 0.007615f
C925 a_1541_n8095# Q3 6.69e-21
C926 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B D2_2 0.004429f
C927 a_1409_7469# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 0.001034f
C928 p2_gen_magic_0.xnor_magic_1.OUT Q1 0.010765f
C929 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.tspc2_magic_0.Q 0.114739f
C930 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_21504_5904# 0.022245f
C931 a_27778_1059# CLK 0.006119f
C932 7b_counter_0.MDFF_3.QB VDD 5.26059f
C933 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5036_n3150# 0.002803f
C934 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q7 0.005739f
C935 a_21381_8741# VDD 0.956678f
C936 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 4e-20
C937 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n5540# 0.093592f
C938 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 9.88e-19
C939 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_7215_10149# 3.58e-20
C940 a_16065_3363# CLK 0.180772f
C941 7b_counter_0.MDFF_3.QB D2_1 0.052739f
C942 7b_counter_0.MDFF_4.LD a_23672_3947# 8.49e-19
C943 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 0.001081f
C944 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B CLK 7.16e-20
C945 a_1209_4557# CLK 0.001676f
C946 a_8523_n8579# Q5 1.41e-19
C947 7b_counter_0.MDFF_4.tspc2_magic_0.Q Q5 0.428297f
C948 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 1.99e-20
C949 p2_gen_magic_0.xnor_magic_5.OUT Q2 1.22e-20
C950 a_12174_n7648# VDD 0.001396f
C951 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_8411_8536# 0.146237f
C952 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_3.QB 0.385018f
C953 a_16065_9774# a_16065_8580# 0.020635f
C954 a_20041_3363# a_20171_1669# 0.005699f
C955 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n4081# 0.092057f
C956 a_24259_4877# Q5 8.26e-19
C957 a_23985_7877# VDD 1.1229f
C958 7b_counter_0.MDFF_3.QB LD 0.050802f
C959 OR_magic_2.A p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.002713f
C960 a_12931_3363# D2_2 0.0012f
C961 a_8713_6842# Q2 0.00818f
C962 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT Q4 0.002358f
C963 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_4235_3947# 3.22e-21
C964 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A Q2 0.052982f
C965 p3_gen_magic_0.xnor_magic_1.OUT a_16186_n8142# 0.274615f
C966 a_11492_n6613# D2_5 0.028948f
C967 a_21381_8741# LD 1.6e-20
C968 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.OUT 5.45e-19
C969 Q4 D2_3 0.555579f
C970 a_13353_n2115# Q4 0.019766f
C971 a_12387_5792# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 1.39e-19
C972 a_15865_2253# a_16065_2253# 0.299584f
C973 a_5054_n6024# a_5470_n6471# 0.011514f
C974 7b_counter_0.MDFF_4.tspc2_magic_0.CLK p2_gen_magic_0.xnor_magic_0.OUT 2.76e-20
C975 mux_magic_0.IN2 P2 4.03e-19
C976 a_17405_2092# a_19307_1669# 2.34e-20
C977 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.0887f
C978 7b_counter_0.MDFF_4.tspc2_magic_0.Q D2_4 4.33e-19
C979 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_2749_684# 0.414018f
C980 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 0.254308f
C981 a_5385_2253# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 1.77e-19
C982 a_15865_6276# Q2 1.29e-19
C983 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 0.003149f
C984 a_11191_4932# a_11279_3480# 0.479729f
C985 a_24259_4877# D2_4 0.007614f
C986 7b_counter_0.MDFF_5.LD DFF_magic_0.D 0.467673f
C987 7b_counter_0.MDFF_3.tspc2_magic_0.CLK CLK 0.047656f
C988 p3_gen_magic_0.3_inp_AND_magic_0.VOUT Q4 0.195804f
C989 a_23985_7877# LD 0.008129f
C990 a_18891_1669# Q5 3.37e-20
C991 7b_counter_0.NAND_magic_0.VOUT D2_4 0.061114f
C992 a_1559_n5540# a_1559_n6024# 0.033537f
C993 Q1 CLK 1.16778f
C994 a_11279_3480# a_12387_3319# 0.001529f
C995 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A Q6 0.023134f
C996 7b_counter_0.3_inp_AND_magic_0.B Q5 8.09e-19
C997 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A Q2 8.26e-19
C998 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1541_n3597# 1.73e-19
C999 a_1559_n5540# Q3 1.41e-19
C1000 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B Q4 0.002457f
C1001 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 8.27e-20
C1002 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8411_3319# 0.001158f
C1003 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT LD 0.00146f
C1004 a_1559_n1973# a_1975_n1973# 0.002223f
C1005 mux_magic_0.AND2_magic_0.A mux_magic_0.OR_magic_0.A 0.001081f
C1006 OR_magic_1.VOUT mux_magic_0.AND2_magic_0.A 8.74e-19
C1007 a_5036_n3150# Q5 3.01e-19
C1008 7b_counter_0.MDFF_5.LD a_23207_5885# 1.42e-19
C1009 a_5470_n6471# VDD 0.003218f
C1010 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.170054f
C1011 p3_gen_magic_0.xnor_magic_1.OUT a_1957_n7648# 0.064748f
C1012 p2_gen_magic_0.xnor_magic_0.OUT VDD 0.592075f
C1013 p2_gen_magic_0.3_inp_AND_magic_0.A a_13553_n2115# 0.075783f
C1014 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B CLK 0.015123f
C1015 mux_magic_0.IN2 VDD 2.00141f
C1016 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VDD 1.23996f
C1017 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.017061f
C1018 a_18891_1669# D2_4 0.016347f
C1019 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 7.14e-19
C1020 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 0.001081f
C1021 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VDD 1.33411f
C1022 7b_counter_0.MDFF_0.tspc2_magic_0.CLK D2_5 0.110195f
C1023 7b_counter_0.3_inp_AND_magic_0.B D2_4 0.006272f
C1024 a_5054_n1973# VDD 0.033235f
C1025 mux_magic_0.IN2 D2_1 0.291291f
C1026 a_19841_3363# VDD 0.92192f
C1027 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VDD 1.17678f
C1028 a_8713_1625# a_9212_739# 0.301553f
C1029 a_13353_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.038495f
C1030 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 0.246208f
C1031 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_3 3.04e-19
C1032 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_11191_10149# 0.189314f
C1033 p2_gen_magic_0.xnor_magic_6.OUT D2_3 0.140213f
C1034 7b_counter_0.NAND_magic_0.VOUT a_24003_10051# 0.78696f
C1035 a_1209_7469# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 0.001158f
C1036 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8939_n3150# 0.005701f
C1037 7b_counter_0.MDFF_4.LD a_27778_1059# 0.004065f
C1038 a_23985_7877# Q3 0.00167f
C1039 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C1040 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT P2 0.001425f
C1041 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.08559f
C1042 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A LD 0.00221f
C1043 a_9212_739# a_9412_739# 0.655098f
C1044 a_12931_3363# CLK 0.133959f
C1045 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1541_n7648# 0.002829f
C1046 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.062422f
C1047 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B D2_5 0.016568f
C1048 7b_counter_0.MDFF_4.LD a_16065_3363# 0.037789f
C1049 7b_counter_0.3_inp_AND_magic_0.B Q2 0.176093f
C1050 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_9412_5956# 1.29e-19
C1051 a_5385_7469# CLK 0.001267f
C1052 p2_gen_magic_0.3_inp_AND_magic_0.A D2_2 0.005997f
C1053 a_5036_n8579# Q5 1.88e-19
C1054 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN VDD 2.03971f
C1055 7b_counter_0.MDFF_7.tspc2_magic_0.Q CLK 0.070476f
C1056 a_5036_n3150# Q2 0.001359f
C1057 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A Q7 6.76e-19
C1058 p3_gen_magic_0.xnor_magic_4.OUT a_11708_n6613# 0.058012f
C1059 OR_magic_1.VOUT divide_by_2_1.tg_magic_2.IN 0.001114f
C1060 a_8939_n7648# VDD 0.001798f
C1061 a_12174_n3150# a_12174_n3597# 0.013884f
C1062 a_24003_10051# 7b_counter_0.3_inp_AND_magic_0.B 2.19e-20
C1063 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN D2_1 0.059695f
C1064 a_24059_4877# Q5 0.001975f
C1065 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A Q5 1.03e-21
C1066 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VDD 1.38749f
C1067 a_11279_6341# Q2 0.132132f
C1068 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B D2_3 4.21e-19
C1069 p3_gen_magic_0.xnor_magic_1.OUT a_14556_n8142# 0.019501f
C1070 a_9059_n6471# D2_5 0.002313f
C1071 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_0.IN 0.311939f
C1072 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n7648# 0.107246f
C1073 a_23352_n5390# a_23352_n6798# 0.479729f
C1074 a_5054_n6024# a_5054_n6471# 0.013665f
C1075 a_17405_2092# a_17405_684# 0.479729f
C1076 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.671219f
C1077 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.08682f
C1078 7b_counter_0.MDFF_5.tspc2_magic_0.D a_11191_5901# 1.08e-19
C1079 p3_gen_magic_0.xnor_magic_3.OUT a_11292_n6613# 0.473167f
C1080 a_23793_5904# a_23560_3728# 4.74e-19
C1081 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_20041_3363# 1.77e-19
C1082 a_12931_6276# Q2 0.02984f
C1083 7b_counter_0.MDFF_6.tspc2_magic_0.Q VDD 1.161f
C1084 7b_counter_0.MDFF_7.tspc2_magic_0.D a_23560_3728# 0.037942f
C1085 p2_gen_magic_0.xnor_magic_0.OUT Q3 0.005062f
C1086 a_24059_4877# D2_4 0.05466f
C1087 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A Q5 0.002209f
C1088 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q3 0.0014f
C1089 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 0.178114f
C1090 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 0.178114f
C1091 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A D2_4 0.020759f
C1092 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_17405_2092# 0.036613f
C1093 a_13353_n6613# Q4 0.020727f
C1094 7b_counter_0.MDFF_6.tspc2_magic_0.Q D2_1 0.169003f
C1095 divide_by_2_1.tg_magic_3.IN OUT1 2.8e-19
C1096 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A LD 0.43461f
C1097 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 1.05e-19
C1098 7b_counter_0.MDFF_4.LD Q1 0.194224f
C1099 a_5185_7469# Q6 2.54e-19
C1100 a_11191_4932# a_12387_3319# 7.51e-20
C1101 a_17405_3524# a_17405_2092# 0.00112f
C1102 a_19841_3363# Q3 1.56e-19
C1103 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.B 0.312144f
C1104 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q1 0.018895f
C1105 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8955_3363# 0.016967f
C1106 a_8643_n1042# D2_6 0.018623f
C1107 a_21504_5904# Q6 0.302465f
C1108 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n8579# 0.064529f
C1109 7b_counter_0.MDFF_1.tspc2_magic_0.D a_15865_1059# 1.63e-20
C1110 OR_magic_2.A a_30365_3514# 0.046739f
C1111 7b_counter_0.MDFF_5.LD a_22991_5885# 1.46e-19
C1112 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_1.IN 0.340787f
C1113 a_5054_n6471# VDD 0.027539f
C1114 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_739# 0.365826f
C1115 a_1541_n7648# a_1957_n7648# 0.002223f
C1116 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT a_16386_n8142# 2.88e-19
C1117 p3_gen_magic_0.xnor_magic_4.OUT a_5054_n5540# 0.299642f
C1118 7b_counter_0.MDFF_6.tspc2_magic_0.Q LD 5.47e-19
C1119 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_10149# 0.189314f
C1120 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12931_4557# 0.037614f
C1121 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A D2_4 0.028914f
C1122 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_21381_8741# 2.4e-20
C1123 p2_gen_magic_0.3_inp_AND_magic_0.A a_11708_n2115# 0.200301f
C1124 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VDD 1.38168f
C1125 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.001424f
C1126 a_1559_n6471# Q6 7.08e-19
C1127 DFF_magic_0.D a_27234_3319# 7.25e-19
C1128 a_5185_2253# VDD 0.959921f
C1129 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 0.00112f
C1130 a_20041_8580# a_20171_6886# 0.005699f
C1131 a_11191_684# D2_4 0.014358f
C1132 a_1209_6275# D2_7 0.001168f
C1133 p2_gen_magic_0.AND2_magic_1.A a_11292_n6613# 1.51e-19
C1134 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12387_4513# 0.149276f
C1135 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1975_n1973# 6.1e-19
C1136 a_27778_4557# VDD 0.064271f
C1137 a_8643_n1526# VDD 0.183902f
C1138 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT D2_7 0.004921f
C1139 7b_counter_0.3_inp_AND_magic_0.VOUT D2_4 0.031443f
C1140 a_5054_n1526# Q6 1.77e-20
C1141 a_1409_9773# a_1209_8579# 0.00289f
C1142 a_13353_n6613# p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 1.26e-20
C1143 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 2.07e-19
C1144 p3_gen_magic_0.xnor_magic_0.OUT VDD 0.592422f
C1145 a_6725_2092# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 2.4e-20
C1146 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n3597# 0.083665f
C1147 a_12387_5792# Q5 1.29e-19
C1148 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_684# 0.189314f
C1149 a_5036_n4081# Q6 0.014859f
C1150 p2_gen_magic_0.3_inp_AND_magic_0.C Q5 6.77e-20
C1151 7b_counter_0.MDFF_4.tspc2_magic_0.D D2_6 0.044265f
C1152 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_7308# 0.431521f
C1153 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q3 3.01e-19
C1154 p3_gen_magic_0.xnor_magic_0.OUT D2_1 0.005056f
C1155 a_13769_n6613# Q4 0.009167f
C1156 a_19841_3363# a_19152_1223# 3.03e-19
C1157 a_5385_6275# Q7 0.009309f
C1158 a_8713_1625# Q4 0.001125f
C1159 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5 0.553421f
C1160 a_5185_2253# LD 0.224142f
C1161 7b_counter_0.MDFF_4.LD a_12931_3363# 0.037687f
C1162 a_1409_2253# D2_5 0.078828f
C1163 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B Q2 0.004929f
C1164 a_12387_6986# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 0.001158f
C1165 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.025092f
C1166 a_2749_7308# CLK 0.010623f
C1167 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_3 0.002723f
C1168 a_8643_n1042# D2_2 0.008527f
C1169 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.009823f
C1170 a_1541_n8579# Q5 0.004247f
C1171 7b_counter_0.3_inp_AND_magic_0.VOUT Q2 3.64e-20
C1172 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.tspc2_magic_0.Q 0.111883f
C1173 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_16065_3363# 1.77e-19
C1174 7b_counter_0.NAND_magic_0.VOUT a_23985_7877# 2.05e-19
C1175 p3_gen_magic_0.xnor_magic_4.OUT a_11492_n6613# 0.116764f
C1176 a_8955_9774# Q7 0.026338f
C1177 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B 0.002977f
C1178 a_9689_1669# D2_6 0.011621f
C1179 a_8713_6842# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 6.16e-19
C1180 p2_gen_magic_0.3_inp_AND_magic_0.C D2_4 0.002177f
C1181 p2_gen_magic_0.AND2_magic_1.A a_12590_n3150# 0.06406f
C1182 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B Q7 0.025895f
C1183 a_5185_6275# a_5385_6275# 0.29829f
C1184 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B D2_3 0.00732f
C1185 a_22150_1124# Q5 0.00127f
C1186 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 0.445787f
C1187 7b_counter_0.3_inp_AND_magic_0.VOUT a_24003_10051# 0.187014f
C1188 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1409_4557# 9.27e-19
C1189 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.255796f
C1190 p3_gen_magic_0.3_inp_AND_magic_0.A D2_2 1.71e-20
C1191 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_19152_5956# 1.29e-19
C1192 a_8643_n6471# D2_5 0.063427f
C1193 a_6725_7308# Q2 4.35e-19
C1194 a_27234_575# CLK 0.007499f
C1195 a_15865_2253# D2_3 0.267131f
C1196 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.001131f
C1197 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5452_n3150# 6.1e-19
C1198 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q5 4.71e-19
C1199 DFF_magic_0.tg_magic_2.IN P2 0.008207f
C1200 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q4 1.6e-19
C1201 a_12387_1769# a_12931_2253# 0.299584f
C1202 a_1559_n6471# a_1975_n6471# 0.002223f
C1203 a_9059_n1973# Q1 0.001283f
C1204 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_17405_4932# 3.58e-20
C1205 a_11279_3480# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 0.132169f
C1206 a_11279_3480# a_11279_1124# 0.00112f
C1207 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 0.006421f
C1208 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_1209_7469# 1.18e-19
C1209 a_5185_2253# a_6725_2092# 0.001529f
C1210 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A Q5 0.289682f
C1211 a_4496_4393# a_5385_2253# 5.39e-19
C1212 a_12387_5792# Q2 0.029793f
C1213 7b_counter_0.3_inp_AND_magic_0.B a_23985_7877# 0.326499f
C1214 OR_magic_2.A P2 0.921344f
C1215 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 0.011087f
C1216 7b_counter_0.MDFF_1.tspc2_magic_0.D CLK 0.001202f
C1217 7b_counter_0.MDFF_5.LD a_8411_8536# 0.224142f
C1218 7b_counter_0.MDFF_4.tspc2_magic_0.D D2_2 0.139822f
C1219 a_19841_4557# a_19841_3363# 0.005574f
C1220 a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 1.93e-19
C1221 a_22150_1124# D2_4 0.012823f
C1222 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5054_n5540# 1.66e-20
C1223 a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 0.149276f
C1224 a_8643_n6471# p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 7.47e-19
C1225 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C1226 7b_counter_0.MDFF_4.tspc2_magic_0.Q 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.27167f
C1227 a_1409_2253# D2_7 0.009158f
C1228 mux_magic_0.AND2_magic_0.A mux_magic_0.IN2 0.01312f
C1229 7b_counter_0.DFF_magic_0.tg_magic_0.IN VDD 0.995698f
C1230 7b_counter_0.MDFF_3.tspc2_magic_0.D a_1209_8579# 7.57e-20
C1231 a_19152_5956# Q6 1.13e-20
C1232 7b_counter_0.3_inp_AND_magic_0.C Q7 1.56e-19
C1233 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q1 0.007097f
C1234 D2_5 D2_6 0.029001f
C1235 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A Q1 0.006453f
C1236 p3_gen_magic_0.xnor_magic_3.OUT a_12174_n8095# 2.99e-20
C1237 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8523_n7648# 3.55e-19
C1238 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_23258_575# 1.93e-19
C1239 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.311939f
C1240 a_1559_n1526# a_1975_n1973# 0.013021f
C1241 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.006256f
C1242 7b_counter_0.MDFF_5.LD a_20041_8580# 0.036926f
C1243 OR_magic_2.A a_30365_4922# 0.313772f
C1244 a_8643_n6024# VDD 0.183902f
C1245 a_12387_4513# a_12931_4557# 0.29829f
C1246 DFF_magic_0.tg_magic_2.IN VDD 1.0454f
C1247 p2_gen_magic_0.3_inp_AND_magic_0.A a_11492_n2115# 1.9e-20
C1248 a_5054_n6024# Q6 0.033582f
C1249 a_11279_3480# VDD 0.941683f
C1250 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B VDD 1.21109f
C1251 7b_counter_0.MDFF_5.LD a_15865_8580# 0.22516f
C1252 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q1 0.01485f
C1253 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VDD 1.37702f
C1254 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n1973# 0.107246f
C1255 DFF_magic_0.D DFF_magic_0.tg_magic_3.OUT 0.830938f
C1256 a_1975_n1973# VDD 0.001798f
C1257 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B D2_1 0.00732f
C1258 a_15865_3363# VDD 0.821263f
C1259 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B 0.005939f
C1260 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_6 1.05502f
C1261 OR_magic_2.A VDD 5.46716f
C1262 p3_gen_magic_0.AND2_magic_1.A a_16386_n8142# 3.84e-19
C1263 a_1541_n8095# a_1541_n8579# 0.033537f
C1264 a_12174_n4081# VDD 0.38976f
C1265 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A Q2 0.001167f
C1266 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_21381_3524# 0.036613f
C1267 a_8411_3319# Q6 1.7e-19
C1268 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.OUT 6.31e-19
C1269 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.02485f
C1270 7b_counter_0.MDFF_3.QB a_5515_9163# 0.183194f
C1271 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.AND2_magic_1.A 0.004455f
C1272 p2_gen_magic_0.xnor_magic_3.OUT Q1 0.143901f
C1273 OR_magic_2.A D2_1 0.256323f
C1274 a_13553_n6613# Q4 0.004585f
C1275 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.164969f
C1276 a_5185_6275# Q7 0.037698f
C1277 a_1209_2253# D2_5 0.04928f
C1278 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19841_4557# 7.48e-20
C1279 VDD Q6 9.770889f
C1280 a_5054_n1973# a_5036_n3150# 0.07324f
C1281 a_8643_n1973# p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 7.47e-19
C1282 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_20171_1669# 0.001268f
C1283 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_6.tspc2_magic_0.Q 0.27167f
C1284 D2_2 D2_5 0.296912f
C1285 a_27778_2253# a_27778_1059# 0.020635f
C1286 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B 0.001758f
C1287 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_9412_739# 1.29e-19
C1288 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN 4.63e-20
C1289 a_4496_9609# Q7 5.19e-19
C1290 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A CLK 0.003072f
C1291 D2_1 Q6 2.17141f
C1292 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_0.OUT 6.89e-21
C1293 a_8825_1669# D2_6 7.93e-19
C1294 a_8939_n3150# a_8523_n3597# 0.013021f
C1295 a_16065_2253# D2_3 0.184192f
C1296 a_27234_575# DFF_magic_0.tg_magic_1.IN 5.2e-21
C1297 7b_counter_0.MDFF_5.LD a_12387_9730# 0.002086f
C1298 a_1209_4557# a_1409_4557# 0.29829f
C1299 a_15865_6276# 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 1.27e-19
C1300 7b_counter_0.3_inp_AND_magic_0.VOUT a_21381_8741# 4.62e-22
C1301 a_8643_n5540# D2_2 0.016545f
C1302 a_23802_1059# CLK 0.005196f
C1303 p2_gen_magic_0.xnor_magic_1.OUT D2_5 0.29534f
C1304 p3_gen_magic_0.xnor_magic_1.OUT a_8523_n8095# 0.003763f
C1305 7b_counter_0.MDFF_4.LD a_27234_575# 0.002843f
C1306 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.AND2_magic_1.A 0.424599f
C1307 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5385_6275# 0.037614f
C1308 a_9212_5956# a_9412_5956# 0.655098f
C1309 p2_gen_magic_0.xnor_magic_4.OUT D2_6 0.042411f
C1310 a_32616_n2458# P2 3.9e-19
C1311 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_0.IN 0.010522f
C1312 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_2 0.001008f
C1313 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD 1.03559f
C1314 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_27234_3319# 0.146237f
C1315 a_27778_3363# D2_4 0.176474f
C1316 LD Q6 1.54473f
C1317 a_8643_n1973# Q1 0.323493f
C1318 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_4932# 4.22e-19
C1319 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 0.006183f
C1320 a_12387_4513# Q5 0.243965f
C1321 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 0.0069f
C1322 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_5515_3947# 0.125951f
C1323 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VDD 1.37768f
C1324 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_1 4.17e-19
C1325 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.tspc2_magic_0.D 0.001213f
C1326 7b_counter_0.MDFF_5.LD a_20041_9774# 0.001095f
C1327 a_7303_8697# a_8411_8536# 0.001529f
C1328 7b_counter_0.3_inp_AND_magic_0.VOUT a_23985_7877# 0.125366f
C1329 a_17405_4932# a_15865_3363# 7.51e-20
C1330 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A D2_4 0.017349f
C1331 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_12387_3319# 1.18e-19
C1332 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_15865_3363# 0.146237f
C1333 a_17405_2092# D2_4 0.01081f
C1334 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.716951f
C1335 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VDD 1.25654f
C1336 p3_gen_magic_0.xnor_magic_5.OUT Q5 0.029587f
C1337 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT D2_1 0.079192f
C1338 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A Q3 0.001508f
C1339 a_1209_1059# Q5 2.32e-19
C1340 a_19841_8580# Q1 0.003448f
C1341 a_8411_4513# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.279825f
C1342 a_1209_2253# D2_7 0.012171f
C1343 a_23793_5904# VDD 1.10023f
C1344 a_1975_n1973# Q3 2.06e-19
C1345 7b_counter_0.MDFF_7.tspc2_magic_0.D VDD 1.41986f
C1346 p2_gen_magic_0.3_inp_AND_magic_0.B D2_5 6.85e-21
C1347 a_2749_8740# a_1209_8579# 0.001529f
C1348 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.3_inp_AND_magic_0.B 0.002474f
C1349 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C1350 a_8955_4557# Q1 6.2e-19
C1351 a_1559_n1526# a_1559_n1973# 0.014233f
C1352 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q5 0.002122f
C1353 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B Q1 0.005199f
C1354 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT D2_3 3.26e-20
C1355 7b_counter_0.MDFF_5.LD a_16065_8580# 0.037687f
C1356 a_1975_n6471# VDD 0.001798f
C1357 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_3.IN 0.805432f
C1358 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_15865_1059# 1.37e-19
C1359 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5452_n7648# 0.005701f
C1360 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT a_16186_n8142# 8.71e-20
C1361 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 0.005939f
C1362 a_32616_n2458# VDD 0.807784f
C1363 a_6725_2092# Q6 0.07537f
C1364 a_11191_4932# VDD 1.55695f
C1365 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B Q2 8.2e-19
C1366 a_16065_7470# VDD 0.018978f
C1367 7b_counter_0.MDFF_3.tspc2_magic_0.Q CLK 0.052924f
C1368 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C1369 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_17405_8741# 0.036613f
C1370 7b_counter_0.MDFF_5.LD a_12387_8536# 0.224216f
C1371 mux_magic_0.IN1 P2 0.047467f
C1372 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A LD 0.00221f
C1373 p2_gen_magic_0.xnor_magic_1.OUT D2_7 0.065228f
C1374 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.240827f
C1375 p2_gen_magic_0.xnor_magic_4.OUT D2_2 0.243893f
C1376 a_32616_n2458# D2_1 0.225381f
C1377 Q3 Q6 0.040639f
C1378 a_1559_n1973# VDD 0.01507f
C1379 a_12387_3319# VDD 0.808402f
C1380 a_16065_7470# D2_1 0.176474f
C1381 a_1209_1059# a_1559_n1042# 7.12e-20
C1382 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1975_n6471# 6.1e-19
C1383 a_23560_3728# VDD 0.784341f
C1384 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.04e-19
C1385 a_11191_684# p2_gen_magic_0.xnor_magic_0.OUT 2.31e-20
C1386 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B Q7 0.016336f
C1387 OR_magic_2.A DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 7.82e-19
C1388 a_8523_n4081# VDD 0.42741f
C1389 p3_gen_magic_0.AND2_magic_1.A a_14756_n8142# 0.037687f
C1390 CLK D2_5 2.04471f
C1391 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_4 0.049044f
C1392 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8523_n3150# 0.002613f
C1393 a_1559_n1973# D2_1 3.7e-19
C1394 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8955_9774# 0.037614f
C1395 7b_counter_0.MDFF_3.QB a_4651_9163# 1.9e-20
C1396 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.B 0.312144f
C1397 a_11708_n6613# Q4 2.92e-19
C1398 a_1209_4557# 7b_counter_0.MDFF_0.tspc2_magic_0.D 1.63e-20
C1399 a_1209_7469# a_2749_7308# 0.001529f
C1400 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n1042# 0.066064f
C1401 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_2749_3524# 0.036613f
C1402 a_9689_6886# D2_6 0.00512f
C1403 p3_gen_magic_0.xnor_magic_5.OUT Q2 1.22e-20
C1404 Q7 D2_3 0.059868f
C1405 a_23560_3728# a_23802_2253# 5.39e-19
C1406 a_1209_1059# Q2 2.01e-19
C1407 7b_counter_0.MDFF_6.tspc2_magic_0.CLK Q6 2.96e-19
C1408 a_12387_575# p2_gen_magic_0.3_inp_AND_magic_0.A 1.55e-20
C1409 7b_counter_0.MDFF_0.tspc2_magic_0.Q D2_5 0.213817f
C1410 7b_counter_0.MDFF_5.LD D2_4 0.10331f
C1411 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A Q7 0.085038f
C1412 p2_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 2.24e-19
C1413 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19307_1669# 0.004104f
C1414 p3_gen_magic_0.xnor_magic_3.OUT Q1 0.298279f
C1415 a_5185_1059# Q4 9.11e-19
C1416 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q2 0.014093f
C1417 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23258_1769# 0.029386f
C1418 a_15865_9774# Q7 6e-19
C1419 p3_gen_magic_0.xnor_magic_4.OUT a_8643_n6471# 7.46e-19
C1420 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.001326f
C1421 a_2749_3524# a_2749_2092# 0.00112f
C1422 mux_magic_0.IN1 VDD 6.47339f
C1423 p2_gen_magic_0.3_inp_AND_magic_0.VOUT D2_3 0.126921f
C1424 a_13353_n2115# p2_gen_magic_0.3_inp_AND_magic_0.VOUT 0.123738f
C1425 a_12174_n3150# a_12590_n3150# 0.002223f
C1426 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_7215_4932# 4.85e-19
C1427 a_8523_n3597# Q5 0.08832f
C1428 a_16065_7470# a_16065_6276# 0.020635f
C1429 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_15865_6276# 1.93e-19
C1430 mux_magic_0.IN1 D2_1 0.052209f
C1431 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.3_inp_AND_magic_0.A 0.913677f
C1432 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.3_inp_AND_magic_0.B 0.004678f
C1433 7b_counter_0.MDFF_4.LD a_23802_1059# 1.1e-19
C1434 a_23793_5904# Q3 0.001578f
C1435 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 0.002402f
C1436 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_5185_6275# 0.279825f
C1437 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.0037f
C1438 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B D2_7 0.004014f
C1439 7b_counter_0.MDFF_5.LD Q2 3.80013f
C1440 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q5 2.97e-19
C1441 a_11279_1124# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.036613f
C1442 a_34156_n2297# OUT1 0.138356f
C1443 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.42e-19
C1444 p2_gen_magic_0.xnor_magic_5.OUT Q6 0.301347f
C1445 a_1559_n6024# a_1975_n6471# 0.013021f
C1446 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN D2_6 6.77e-19
C1447 CLK D2_7 0.690409f
C1448 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_4651_3947# 0.069391f
C1449 7b_counter_0.MDFF_7.tspc2_magic_0.D a_26126_3480# 0.134004f
C1450 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A Q7 0.097202f
C1451 a_1975_n6471# Q3 2.48e-20
C1452 a_30365_3514# P2 0.497716f
C1453 p2_gen_magic_0.xnor_magic_4.OUT a_11708_n2115# 0.058012f
C1454 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK 0.005192f
C1455 a_8713_6842# Q6 1.07e-20
C1456 7b_counter_0.MDFF_5.LD a_24003_10051# 0.221427f
C1457 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_11279_3480# 0.001371f
C1458 a_9689_6886# D2_2 8.15e-21
C1459 p3_gen_magic_0.xnor_magic_4.OUT D2_6 3.57e-20
C1460 a_5036_n7648# Q5 0.689995f
C1461 a_5185_7469# VDD 0.959921f
C1462 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_11292_n6613# 2.84e-20
C1463 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT D2_3 4.44e-19
C1464 7b_counter_0.MDFF_1.tspc2_magic_0.CLK CLK 0.118636f
C1465 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 0.0069f
C1466 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN D2_6 0.026749f
C1467 OR_magic_2.A a_23352_n5390# 0.396399f
C1468 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_9689_6886# 1.32e-19
C1469 a_32616_n1264# a_32616_n2458# 0.005574f
C1470 a_21504_5904# VDD 1.13183f
C1471 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5036_n3597# 6.98e-21
C1472 a_1559_n1973# Q3 0.309627f
C1473 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A Q7 0.023977f
C1474 7b_counter_0.MDFF_7.tspc2_magic_0.CLK Q5 0.012426f
C1475 a_2749_10148# a_1209_8579# 7.51e-20
C1476 a_23560_3728# Q3 0.004225f
C1477 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_3 1.35e-19
C1478 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 3.73e-20
C1479 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1559_n1042# 5.58e-20
C1480 a_30365_4922# a_30365_3514# 0.479677f
C1481 a_19841_9774# Q1 1.63e-20
C1482 a_11292_n2115# Q5 6.77e-20
C1483 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VDD 1.24096f
C1484 OR_magic_2.A mux_magic_0.AND2_magic_0.A 0.003211f
C1485 7b_counter_0.MDFF_5.LD a_12931_8580# 0.037789f
C1486 a_26126_3480# a_23560_3728# 6.34e-20
C1487 a_1559_n6471# VDD 0.01507f
C1488 a_20171_1669# Q1 0.002438f
C1489 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A Q1 2.58e-19
C1490 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A CLK 0.015982f
C1491 7b_counter_0.MDFF_5.tspc2_magic_0.D D2_6 0.079906f
C1492 a_4235_9163# CLK 0.008175f
C1493 7b_counter_0.MDFF_0.tspc2_magic_0.Q p2_gen_magic_0.xnor_magic_4.OUT 4.61e-20
C1494 a_12931_7470# VDD 0.002522f
C1495 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A Q4 8.78e-21
C1496 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_19841_3363# 0.146237f
C1497 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A Q6 4.09e-19
C1498 p3_gen_magic_0.3_inp_AND_magic_0.B D2_5 0.031674f
C1499 a_5185_7469# LD 0.224142f
C1500 a_1541_n3150# D2_7 0.001642f
C1501 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q2 0.100114f
C1502 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n1526# 0.063777f
C1503 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 0.002584f
C1504 7b_counter_0.MDFF_4.tspc2_magic_0.Q Q6 2.13e-19
C1505 a_5054_n1526# VDD 0.236943f
C1506 7b_counter_0.MDFF_7.tspc2_magic_0.CLK D2_4 0.248686f
C1507 a_30365_3514# VDD 1.17434f
C1508 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n6471# 0.107246f
C1509 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q5 0.011033f
C1510 a_1409_3363# VDD 0.012214f
C1511 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7303_3480# 0.431521f
C1512 a_11191_5901# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 3.58e-20
C1513 a_5036_n4081# VDD 0.508913f
C1514 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_4235_3947# 6.31e-20
C1515 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12590_n3150# 0.005701f
C1516 a_12387_6986# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 0.146237f
C1517 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 0.178114f
C1518 a_11292_n2115# D2_4 0.006368f
C1519 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_1409_1059# 9.27e-19
C1520 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_5 0.045037f
C1521 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_2749_4932# 0.414018f
C1522 a_1209_4557# a_2749_3524# 7.54e-20
C1523 a_21381_10149# a_21381_8741# 0.479729f
C1524 p3_gen_magic_0.xnor_magic_4.OUT D2_2 0.162528f
C1525 a_8825_6886# D2_6 5.11e-19
C1526 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD 1.03776f
C1527 a_5036_n7648# Q2 1.88e-19
C1528 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5036_n7648# 1.55e-19
C1529 mux_magic_0.IN1 a_32616_n1264# 0.412086f
C1530 a_15865_7470# D2_3 0.002075f
C1531 a_4235_3947# D2_5 0.033779f
C1532 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_4 0.07307f
C1533 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT a_23352_n5390# 1.09e-19
C1534 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_1 5.05e-21
C1535 a_1409_3363# LD 0.037687f
C1536 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_4932# 1.51e-21
C1537 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_9212_5956# 4.79e-21
C1538 a_6725_684# Q1 0.007505f
C1539 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_4.OUT 1.35e-19
C1540 mux_magic_0.IN1 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 0.004003f
C1541 a_27234_1769# VDD 0.807784f
C1542 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 2.42e-19
C1543 a_13353_n2115# D2_3 0.021243f
C1544 7b_counter_0.MDFF_5.tspc2_magic_0.D D2_2 0.012265f
C1545 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_14756_n3644# 0.002513f
C1546 a_23352_n6798# p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 0.003963f
C1547 a_5036_n3597# Q5 2.14e-20
C1548 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A CLK 1.75e-19
C1549 a_9689_6886# CLK 0.00188f
C1550 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_6.tspc2_magic_0.D 0.008512f
C1551 7b_counter_0.3_inp_AND_magic_0.B Q6 0.065627f
C1552 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT LD 1.2e-19
C1553 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.025171f
C1554 a_8523_n7648# p3_gen_magic_0.xnor_magic_6.OUT 0.103719f
C1555 a_21504_5904# Q3 0.190794f
C1556 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_17405_3524# 1.23e-19
C1557 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_11279_1124# 0.018271f
C1558 a_1409_7469# D2_7 0.034642f
C1559 a_7303_8697# Q2 0.172018f
C1560 a_5036_n3150# Q6 0.332475f
C1561 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q2 0.067441f
C1562 a_27234_3319# D2_4 0.26156f
C1563 a_1559_n6024# a_1559_n6471# 0.014233f
C1564 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q5 0.021475f
C1565 p3_gen_magic_0.3_inp_AND_magic_0.VOUT D2_3 0.007114f
C1566 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_1.IN 4.63e-20
C1567 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_6 0.059388f
C1568 7b_counter_0.MDFF_4.tspc2_magic_0.D a_12387_575# 1.63e-20
C1569 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.025047f
C1570 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A Q3 2.33e-19
C1571 a_1559_n6471# Q3 0.306674f
C1572 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24259_4877# 0.120019f
C1573 p2_gen_magic_0.xnor_magic_4.OUT a_11492_n2115# 0.116764f
C1574 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN Q4 0.013263f
C1575 a_30365_4922# P2 0.189462f
C1576 a_23207_5885# Q1 0.005661f
C1577 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_7 0.002161f
C1578 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 8.64e-19
C1579 7b_counter_0.MDFF_4.LD a_8825_1669# 8.49e-19
C1580 a_2749_5900# Q6 0.014805f
C1581 a_1209_6275# 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A 1.28e-19
C1582 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 0.002753f
C1583 a_7303_3480# Q7 0.039081f
C1584 a_8643_n1526# p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.86e-20
C1585 a_8825_6886# D2_2 4.45e-19
C1586 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8411_3319# 4.65e-19
C1587 a_1957_n7648# Q5 0.001196f
C1588 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 0.086059f
C1589 a_16065_4557# CLK 0.00402f
C1590 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A Q7 0.012645f
C1591 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_0.OUT 6.88e-21
C1592 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_21504_5904# 1.75e-21
C1593 mux_magic_0.AND2_magic_0.A a_32616_n2458# 0.001158f
C1594 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8825_6886# 0.001268f
C1595 a_19152_5956# VDD 0.725343f
C1596 a_21381_3524# Q5 0.005555f
C1597 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B D2_4 0.011275f
C1598 VDD P2 4.88028f
C1599 a_15865_4557# Q1 8.5e-19
C1600 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1541_n8095# 1.73e-19
C1601 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.205429f
C1602 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN CLK 0.001114f
C1603 a_2749_684# VDD 1.55812f
C1604 7b_counter_0.MDFF_4.tspc2_magic_0.D p2_gen_magic_0.xnor_magic_3.OUT 2.45e-19
C1605 7b_counter_0.MDFF_4.tspc2_magic_0.CLK VDD 2.19796f
C1606 a_19152_6440# Q7 4.12e-19
C1607 a_11279_1124# VDD 0.94863f
C1608 7b_counter_0.MDFF_5.LD a_23985_7877# 7.97e-20
C1609 a_24259_4877# a_23560_3728# 0.014143f
C1610 a_5054_n6024# VDD 0.225572f
C1611 a_19307_1669# Q1 0.00207f
C1612 D2_1 P2 0.529739f
C1613 a_26126_1124# CLK 0.063008f
C1614 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.003053f
C1615 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q3 0.006143f
C1616 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q4 0.001088f
C1617 a_5036_n3597# Q2 6.69e-21
C1618 a_5036_n8579# Q6 1.79e-19
C1619 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN CLK 0.709192f
C1620 a_8411_4513# Q6 4.96e-20
C1621 a_30365_4922# VDD 1.59406f
C1622 a_1559_n1526# VDD 0.183944f
C1623 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q5 0.542565f
C1624 a_8411_3319# VDD 0.921912f
C1625 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_5900# 0.414018f
C1626 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.003249f
C1627 p3_gen_magic_0.AND2_magic_1.A a_14556_n8142# 0.232114f
C1628 a_1541_n4081# VDD 0.425848f
C1629 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_1209_1059# 0.149276f
C1630 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q1 0.046247f
C1631 a_5385_7469# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 1.77e-19
C1632 a_27234_1769# Q3 2.98e-19
C1633 a_1559_n1526# D2_1 5.31e-19
C1634 a_2749_684# LD 0.002672f
C1635 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q4 8.46e-19
C1636 a_13353_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.038495f
C1637 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_20171_6886# 0.001268f
C1638 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.001478f
C1639 a_1209_4557# a_2749_4932# 0.002003f
C1640 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A D2_5 4.23e-19
C1641 a_1541_n4081# D2_1 0.09803f
C1642 mux_magic_0.IN1 mux_magic_0.AND2_magic_0.A 0.497755f
C1643 7b_counter_0.MDFF_5.tspc2_magic_0.D CLK 0.003746f
C1644 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.014848f
C1645 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.014655f
C1646 a_1541_n4081# p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 1.57e-20
C1647 VDD D2_1 8.86669f
C1648 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_5 0.085517f
C1649 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12931_7470# 1.77e-19
C1650 p2_gen_magic_0.xnor_magic_5.OUT a_5036_n4081# 0.417238f
C1651 a_23802_2253# VDD 0.087968f
C1652 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VDD 1.03134f
C1653 a_9212_739# D2_6 0.064777f
C1654 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT 0.169047f
C1655 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B Q6 6.05e-19
C1656 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 0.434557f
C1657 a_8825_6886# CLK 0.002315f
C1658 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VDD 1.27697f
C1659 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_1 3.98e-19
C1660 a_1957_n7648# a_1541_n8095# 0.013021f
C1661 VDD LD 20.47f
C1662 a_27234_1769# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 0.146237f
C1663 a_1209_7469# D2_7 0.019201f
C1664 p2_gen_magic_0.xnor_magic_3.OUT D2_5 0.041341f
C1665 7b_counter_0.3_inp_AND_magic_0.VOUT Q6 1.06e-20
C1666 a_24536_3947# D2_4 0.009911f
C1667 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n5540# 0.066064f
C1668 Q3 P2 0.016451f
C1669 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A D2_1 0.009291f
C1670 a_13353_n6613# D2_3 0.015364f
C1671 LD D2_1 0.917349f
C1672 a_2749_684# Q3 3.98e-19
C1673 a_23793_5904# a_24059_4877# 2.1e-21
C1674 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.287011f
C1675 7b_counter_0.MDFF_4.tspc2_magic_0.CLK Q3 4.75e-19
C1676 7b_counter_0.MDFF_3.QB a_7303_8697# 0.003632f
C1677 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_15865_4557# 1.39e-19
C1678 a_13769_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.002312f
C1679 a_12931_9774# Q7 0.026338f
C1680 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24059_4877# 0.282223f
C1681 a_13769_n2115# Q4 0.007219f
C1682 7b_counter_0.MDFF_5.LD 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.002173f
C1683 a_22991_5885# Q1 0.216721f
C1684 a_6725_7308# Q6 0.25224f
C1685 mux_magic_0.IN1 divide_by_2_1.tg_magic_2.IN 0.327622f
C1686 7b_counter_0.MDFF_4.LD a_16065_4557# 0.003356f
C1687 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_5956# 0.363339f
C1688 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A LD 0.443289f
C1689 a_19841_3363# a_20041_3363# 0.297401f
C1690 a_27778_4557# a_27778_3363# 0.020635f
C1691 a_13353_n6613# p3_gen_magic_0.3_inp_AND_magic_0.VOUT 0.123693f
C1692 a_16065_6276# VDD 0.065403f
C1693 a_1559_n1526# Q3 0.08832f
C1694 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT Q4 8.43e-19
C1695 p2_gen_magic_0.xnor_magic_0.OUT a_8523_n3597# 0.011792f
C1696 7b_counter_0.MDFF_1.tspc2_magic_0.D a_20171_1669# 2.1e-20
C1697 a_17405_8741# D2_3 0.00152f
C1698 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_7 6.27e-21
C1699 a_16065_6276# D2_1 0.003998f
C1700 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 0.004678f
C1701 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT P2 0.001425f
C1702 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 0.913677f
C1703 a_17405_4932# VDD 1.55668f
C1704 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 6.95e-19
C1705 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 0.001081f
C1706 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK 1.35031f
C1707 a_9212_739# D2_2 0.001077f
C1708 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5515_3947# 0.001268f
C1709 a_6725_2092# VDD 0.955478f
C1710 a_1559_n6024# VDD 0.183944f
C1711 a_24059_4877# a_23560_3728# 0.301553f
C1712 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B VDD 1.21103f
C1713 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27778_4557# 9.27e-19
C1714 a_17405_684# Q1 0.001194f
C1715 7b_counter_0.MDFF_4.LD a_26126_1124# 0.001152f
C1716 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 9.92e-19
C1717 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_11279_3480# 2.4e-20
C1718 7b_counter_0.3_inp_AND_magic_0.B a_21504_5904# 0.900342f
C1719 a_12174_n8579# VDD 0.392783f
C1720 a_1409_9773# CLK 4.61e-19
C1721 a_1409_2253# Q4 0.002005f
C1722 VDD Q3 9.25996f
C1723 a_15865_9774# a_17405_8741# 7.54e-20
C1724 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A a_23258_575# 0.279825f
C1725 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.0037f
C1726 a_1541_n8579# Q6 1.74e-19
C1727 p2_gen_magic_0.xnor_magic_3.OUT D2_7 0.047478f
C1728 a_32616_n1264# VDD 0.914128f
C1729 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A Q1 0.004342f
C1730 D2_1 Q3 0.153356f
C1731 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1559_n6024# 0.063777f
C1732 a_26126_3480# VDD 0.955854f
C1733 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.tspc2_magic_0.Q 0.125613f
C1734 a_13769_n6613# D2_3 0.001839f
C1735 a_19152_6440# D2_3 0.026411f
C1736 a_17405_3524# Q1 0.017029f
C1737 a_8713_1625# D2_3 2.66e-19
C1738 a_16386_n3644# VDD 0.024812f
C1739 p3_gen_magic_0.AND2_magic_1.A a_12174_n8095# 0.371679f
C1740 7b_counter_0.3_inp_AND_magic_0.A Q4 0.045521f
C1741 a_23802_2253# Q3 4.83e-19
C1742 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q3 0.005773f
C1743 a_32616_n1264# D2_1 3.96e-19
C1744 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B Q1 0.007329f
C1745 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19307_6886# 1.2e-19
C1746 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.005763f
C1747 p2_gen_magic_0.xnor_magic_0.OUT a_11292_n2115# 0.394147f
C1748 7b_counter_0.MDFF_6.tspc2_magic_0.CLK VDD 2.20412f
C1749 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A D2_2 0.002102f
C1750 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A Q1 0.00647f
C1751 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_3.OUT 0.871612f
C1752 DFF_magic_0.D a_27234_575# 1.85e-19
C1753 a_16386_n3644# D2_1 0.023133f
C1754 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q6 0.001431f
C1755 7b_counter_0.MDFF_1.tspc2_magic_0.Q Q5 0.476265f
C1756 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_5.tspc2_magic_0.D 0.008512f
C1757 a_13769_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.002312f
C1758 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VDD 1.08651f
C1759 LD Q3 0.010453f
C1760 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A Q1 0.302946f
C1761 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_5.tspc2_magic_0.Q 0.002402f
C1762 p3_gen_magic_0.3_inp_AND_magic_0.VOUT a_13769_n6613# 0.200301f
C1763 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.07839f
C1764 p2_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.3_inp_AND_magic_0.A 3.55e-20
C1765 a_1409_4557# D2_5 0.004183f
C1766 7b_counter_0.MDFF_6.tspc2_magic_0.CLK D2_1 0.124591f
C1767 a_15865_7470# a_17405_7309# 0.001529f
C1768 p3_gen_magic_0.xnor_magic_1.OUT D2_5 3.68e-19
C1769 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B VDD 1.19227f
C1770 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 1.19e-19
C1771 a_19152_1223# VDD 0.764146f
C1772 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VDD 1.03888f
C1773 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_14556_n3644# 0.008182f
C1774 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_3 9.74e-19
C1775 7b_counter_0.MDFF_1.tspc2_magic_0.Q D2_4 0.00648f
C1776 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8939_n3150# 6.1e-19
C1777 p2_gen_magic_0.xnor_magic_5.OUT VDD 1.9483f
C1778 a_17405_7309# D2_3 0.029476f
C1779 Q4 D2_6 3.18631f
C1780 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B a_17405_4932# 0.189314f
C1781 a_23672_3947# D2_4 6.09e-19
C1782 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.010798f
C1783 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_9689_6886# 0.069391f
C1784 p2_gen_magic_0.xnor_magic_5.OUT D2_1 1.51101f
C1785 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n7648# 0.011524f
C1786 a_8713_6842# VDD 0.767425f
C1787 a_13553_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.011362f
C1788 7b_counter_0.MDFF_4.tspc2_magic_0.Q 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 0.005065f
C1789 a_1559_n6024# Q3 0.08832f
C1790 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VDD 1.25149f
C1791 p2_gen_magic_0.xnor_magic_4.OUT a_8643_n1973# 7.46e-19
C1792 a_13553_n2115# Q4 0.00847f
C1793 mux_magic_0.AND2_magic_0.A P2 0.009922f
C1794 a_20041_8580# Q1 0.00357f
C1795 7b_counter_0.MDFF_3.tspc2_magic_0.D CLK 0.00841f
C1796 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1209_3363# 0.001985f
C1797 OR_magic_1.VOUT divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 1.3249f
C1798 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 1.32477f
C1799 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12931_3363# 1.77e-19
C1800 p3_gen_magic_0.xnor_magic_3.OUT D2_5 0.124584f
C1801 a_8939_n3150# Q1 0.006998f
C1802 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n4081# 0.066064f
C1803 a_15865_8580# Q1 0.015458f
C1804 a_15865_6276# VDD 0.944161f
C1805 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A Q2 0.095215f
C1806 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8411_3319# 0.029386f
C1807 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_16065_4557# 9.27e-19
C1808 a_20171_6886# Q6 1.27e-19
C1809 a_2749_2092# D2_4 0.004216f
C1810 7b_counter_0.MDFF_1.tspc2_magic_0.D a_19307_1669# 0.004574f
C1811 p3_gen_magic_0.xnor_magic_1.OUT D2_7 1.68414f
C1812 a_15865_6276# D2_1 2.51e-19
C1813 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_19152_739# 1.29e-19
C1814 a_17405_2092# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 2.4e-20
C1815 a_19841_4557# VDD 0.941676f
C1816 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_4651_3947# 0.004104f
C1817 a_4235_3947# a_5515_3947# 0.007202f
C1818 a_23352_n5390# VDD 1.56587f
C1819 a_5054_n1973# a_5036_n3597# 6.43e-20
C1820 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK D2_6 0.29354f
C1821 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VDD 1.3105f
C1822 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11191_5901# 0.189314f
C1823 a_7215_10149# CLK 0.001996f
C1824 a_8523_n8579# VDD 0.430465f
C1825 a_12387_4513# a_11279_3480# 7.54e-20
C1826 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_11191_4932# 3.58e-20
C1827 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A CLK 0.006122f
C1828 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 0.001081f
C1829 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_9059_n6471# 6.1e-19
C1830 a_15865_1059# Q4 4.47e-19
C1831 a_12174_n3597# a_12174_n4081# 0.033537f
C1832 a_23352_n5390# D2_1 0.011324f
C1833 7b_counter_0.MDFF_0.tspc2_magic_0.D D2_5 0.003828f
C1834 a_1209_9773# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 1.37e-19
C1835 7b_counter_0.MDFF_4.tspc2_magic_0.Q VDD 1.22618f
C1836 D2_2 Q4 0.471976f
C1837 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11191_684# 0.414018f
C1838 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A D2_1 0.012926f
C1839 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.001864f
C1840 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_4496_4393# 0.001157f
C1841 mux_magic_0.AND2_magic_0.A VDD 1.29314f
C1842 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12387_3319# 0.001158f
C1843 a_24259_4877# VDD 0.732917f
C1844 a_13553_n6613# D2_3 8.12e-19
C1845 a_18891_6886# D2_3 0.042648f
C1846 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_27778_2253# 1.77e-19
C1847 a_12931_4557# Q1 6.2e-19
C1848 p2_gen_magic_0.xnor_magic_6.OUT D2_6 0.223057f
C1849 p2_gen_magic_0.AND2_magic_1.A D2_5 0.276014f
C1850 a_14756_n3644# VDD 0.050613f
C1851 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B Q3 0.017749f
C1852 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_6 0.127562f
C1853 a_5185_7469# a_6725_7308# 0.001529f
C1854 a_19152_1223# Q3 8.01e-20
C1855 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n8579# 0.092057f
C1856 7b_counter_0.NAND_magic_0.VOUT VDD 1.39876f
C1857 mux_magic_0.AND2_magic_0.A D2_1 0.43595f
C1858 p3_gen_magic_0.xnor_magic_3.OUT D2_7 0.370036f
C1859 a_16065_9774# VDD 0.061661f
C1860 p2_gen_magic_0.xnor_magic_1.OUT Q4 0.184223f
C1861 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_1.IN 4.63e-20
C1862 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A LD 6.12e-19
C1863 a_4496_4393# D2_5 5.51e-20
C1864 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.OUT 5.45e-19
C1865 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.205497f
C1866 a_13553_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.011362f
C1867 a_12387_9730# Q1 0.243714f
C1868 a_8411_9730# a_7215_10149# 0.002003f
C1869 a_21381_10149# Q6 0.058283f
C1870 p3_gen_magic_0.3_inp_AND_magic_0.VOUT a_13553_n6613# 1.9e-20
C1871 a_13353_n6613# a_13769_n6613# 0.278913f
C1872 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8411_9730# 0.149276f
C1873 a_21381_3524# a_19841_3363# 0.001529f
C1874 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A CLK 0.012578f
C1875 a_15865_6276# a_16065_6276# 0.29829f
C1876 a_8523_n8095# Q5 0.08832f
C1877 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.tspc2_magic_0.D 0.414986f
C1878 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1975_n1973# 0.005701f
C1879 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT Q4 8.15e-19
C1880 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_7 0.037541f
C1881 p2_gen_magic_0.xnor_magic_5.OUT a_16386_n3644# 0.037687f
C1882 a_18891_1669# VDD 0.975666f
C1883 p3_gen_magic_0.xnor_magic_5.OUT Q6 0.16189f
C1884 7b_counter_0.NAND_magic_0.VOUT LD 0.081141f
C1885 7b_counter_0.3_inp_AND_magic_0.B VDD 0.672452f
C1886 a_5054_n1042# D2_3 0.008663f
C1887 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_12387_9730# 1.93e-19
C1888 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n3597# 0.063777f
C1889 a_8955_8580# a_8825_6886# 0.005699f
C1890 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_15865_4557# 1.27e-19
C1891 p2_gen_magic_0.3_inp_AND_magic_0.B Q4 0.050853f
C1892 a_5036_n3150# VDD 0.042066f
C1893 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B D2_6 0.008024f
C1894 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q5 0.005773f
C1895 divide_by_2_1.tg_magic_2.IN VDD 1.04065f
C1896 a_11292_n6613# p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.001281f
C1897 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8825_6886# 0.125951f
C1898 p2_gen_magic_0.xnor_magic_6.OUT D2_2 0.200027f
C1899 DFF_magic_0.tg_magic_0.IN VDD 0.995698f
C1900 a_19841_4557# Q3 4.85e-20
C1901 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2 0.970617f
C1902 OR_magic_2.A p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 1.49e-19
C1903 a_2749_5900# VDD 1.55812f
C1904 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_3 6.21e-19
C1905 a_12931_4557# a_12931_3363# 0.020635f
C1906 a_11708_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.006564f
C1907 a_11279_6341# VDD 0.93439f
C1908 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_26038_4932# 0.189314f
C1909 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_6725_2092# 0.001342f
C1910 a_11708_n2115# Q4 0.008537f
C1911 a_16065_8580# Q1 0.050153f
C1912 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A CLK 0.018587f
C1913 a_2749_8740# CLK 0.016052f
C1914 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_3 1.35e-19
C1915 a_1209_4557# a_1209_3363# 0.005574f
C1916 a_21504_5904# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 5.98e-19
C1917 7b_counter_0.3_inp_AND_magic_0.B LD 0.009811f
C1918 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A P2 5.23e-20
C1919 7b_counter_0.MDFF_5.LD Q6 0.157166f
C1920 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 1.08482f
C1921 a_12387_8536# Q1 0.015128f
C1922 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_15865_6276# 1.37e-19
C1923 a_12931_6276# VDD 0.057637f
C1924 a_27778_4557# a_27234_3319# 0.003083f
C1925 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.079909f
C1926 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 3.27e-20
C1927 CLK Q4 1.39104f
C1928 7b_counter_0.MDFF_3.tspc2_magic_0.Q 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 0.002402f
C1929 Q1 Q5 0.827613f
C1930 a_16065_3363# Q2 0.002005f
C1931 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B Q2 1.74e-19
C1932 a_8411_4513# a_8411_3319# 0.005574f
C1933 7b_counter_0.MDFF_1.tspc2_magic_0.D a_17405_684# 1.08e-19
C1934 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19841_4557# 2.09e-19
C1935 a_1541_n7648# D2_7 4.31e-19
C1936 mux_magic_0.AND2_magic_0.A a_32616_n1264# 0.240798f
C1937 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8939_n7648# 0.005701f
C1938 a_4235_3947# a_4651_3947# 0.16113f
C1939 a_2749_5900# LD 0.002672f
C1940 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_20171_1669# 0.125951f
C1941 a_24259_4877# a_26126_3480# 1.39e-20
C1942 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 0.003149f
C1943 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A D2_2 0.015198f
C1944 a_17405_8741# a_17405_7309# 0.00112f
C1945 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B a_12387_8536# 0.146237f
C1946 a_5185_2253# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B 0.146237f
C1947 a_8713_1625# a_9412_739# 0.014143f
C1948 a_15865_2253# a_16065_1059# 0.003083f
C1949 a_12387_4513# a_11191_4932# 0.002003f
C1950 a_5036_n8579# VDD 0.490263f
C1951 a_11279_1124# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 2.4e-20
C1952 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q4 9.85e-19
C1953 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n6471# 0.107246f
C1954 a_14756_n3644# a_16386_n3644# 0.003333f
C1955 a_8411_4513# VDD 0.937845f
C1956 a_2749_3524# D2_5 0.042236f
C1957 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.272186f
C1958 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B D2_2 0.022957f
C1959 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_11191_684# 0.00215f
C1960 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5054_n5540# 1.54e-20
C1961 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 0.001081f
C1962 Q1 D2_4 0.073837f
C1963 a_11279_1124# a_11191_684# 0.479729f
C1964 a_24059_4877# VDD 0.982676f
C1965 a_12387_4513# a_12387_3319# 0.005574f
C1966 a_11708_n6613# D2_3 0.001839f
C1967 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.xnor_magic_6.OUT 0.197787f
C1968 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 6.36e-20
C1969 a_12174_n7648# a_12174_n8095# 0.013884f
C1970 a_16186_n3644# VDD 0.819774f
C1971 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VDD 1.31563f
C1972 a_8523_n3150# D2_6 0.121793f
C1973 7b_counter_0.3_inp_AND_magic_0.B Q3 0.282789f
C1974 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8523_n7648# 1.55e-19
C1975 a_17405_7309# a_19152_6440# 6.34e-20
C1976 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 0.979103f
C1977 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK CLK 0.876599f
C1978 a_16186_n3644# D2_1 0.01697f
C1979 a_5515_9163# VDD 0.097366f
C1980 a_11708_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.006564f
C1981 7b_counter_0.MDFF_3.tspc2_magic_0.CLK Q2 0.002813f
C1982 a_13353_n6613# a_13553_n6613# 0.522094f
C1983 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_23802_2253# 1.77e-19
C1984 a_5185_1059# D2_3 0.001472f
C1985 Q1 Q2 0.496306f
C1986 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_6 1.86e-19
C1987 a_1559_n1526# a_1957_n3150# 3.01e-19
C1988 a_5036_n8095# Q5 5.75e-19
C1989 a_12931_3363# Q5 0.066427f
C1990 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VDD 1.29631f
C1991 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n1973# 0.011524f
C1992 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12931_9774# 9.27e-19
C1993 DFF_magic_0.D DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.313982f
C1994 a_8713_6842# 7b_counter_0.MDFF_4.tspc2_magic_0.Q 0.001156f
C1995 p2_gen_magic_0.xnor_magic_5.OUT a_14756_n3644# 0.028482f
C1996 p2_gen_magic_0.xnor_magic_6.OUT CLK 8.13e-19
C1997 a_11191_684# VDD 1.55668f
C1998 7b_counter_0.MDFF_5.LD a_16065_7470# 0.037789f
C1999 7b_counter_0.MDFF_0.tspc2_magic_0.CLK Q7 0.045901f
C2000 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B VDD 1.19335f
C2001 a_5036_n7648# Q6 0.319301f
C2002 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q5 0.147667f
C2003 a_9412_5956# D2_6 0.041406f
C2004 a_5385_2253# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 5.46e-20
C2005 7b_counter_0.3_inp_AND_magic_0.VOUT VDD 2.52333f
C2006 a_5515_9163# LD 8.49e-19
C2007 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B Q2 8.23e-19
C2008 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_5901# 0.189314f
C2009 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B D2_1 3.46e-19
C2010 a_1957_n3150# VDD 0.001798f
C2011 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.014172f
C2012 a_11191_5901# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 4.22e-19
C2013 a_18891_1669# a_19152_1223# 0.301553f
C2014 divide_by_2_1.tg_magic_2.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 0.270406f
C2015 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_3.OUT 0.871612f
C2016 p3_gen_magic_0.xnor_magic_0.OUT a_11292_n6613# 0.394147f
C2017 a_5185_6275# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 2.1e-19
C2018 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.42e-19
C2019 a_1541_n3597# D2_7 0.002133f
C2020 a_8523_n3150# D2_2 5.07e-19
C2021 a_1957_n3150# D2_1 0.005701f
C2022 a_19152_5956# a_20041_4557# 3.41e-19
C2023 a_5054_n5540# D2_3 0.010876f
C2024 DFF_magic_0.tg_magic_0.IN DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.272186f
C2025 a_11492_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.00991f
C2026 DFF_magic_0.D 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 2.04e-19
C2027 a_6725_7308# VDD 0.954322f
C2028 7b_counter_0.MDFF_7.tspc2_magic_0.Q D2_4 0.360297f
C2029 a_12931_8580# Q1 0.006533f
C2030 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q7 0.027307f
C2031 a_11492_n2115# Q4 0.009572f
C2032 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.439554f
C2033 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19841_3363# 0.029386f
C2034 a_2749_10148# CLK 0.002001f
C2035 a_27234_4513# CLK 6.38e-19
C2036 p3_gen_magic_0.3_inp_AND_magic_0.B Q4 0.090642f
C2037 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A CLK 0.06685f
C2038 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B LD 6.07e-19
C2039 a_7303_8697# Q6 6.49e-19
C2040 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 0.00112f
C2041 a_13553_n6613# a_13769_n6613# 0.329078f
C2042 7b_counter_0.3_inp_AND_magic_0.VOUT LD 0.163419f
C2043 a_18891_6886# a_19152_6440# 0.301553f
C2044 a_12387_5792# VDD 0.9315f
C2045 a_5036_n3150# p2_gen_magic_0.xnor_magic_5.OUT 0.09365f
C2046 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_2 1.04315f
C2047 7b_counter_0.MDFF_4.LD Q4 3.32919f
C2048 a_5036_n8095# Q2 6.69e-21
C2049 a_24059_4877# Q3 0.002091f
C2050 p2_gen_magic_0.3_inp_AND_magic_0.C VDD 2.56477f
C2051 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5036_n8095# 9.93e-20
C2052 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n8095# 0.083665f
C2053 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A CLK 0.026514f
C2054 a_15865_4557# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 1.63e-20
C2055 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.859117f
C2056 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A Q3 0.001691f
C2057 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q4 1.64e-19
C2058 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD 1.18306f
C2059 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_15865_1059# 1.93e-19
C2060 a_16065_2253# a_16065_1059# 0.020635f
C2061 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 8.78e-21
C2062 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19307_1669# 0.069391f
C2063 a_4496_4877# a_4651_3947# 0.001643f
C2064 a_24059_4877# a_26126_3480# 0.002118f
C2065 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q2 2.32e-20
C2066 p2_gen_magic_0.3_inp_AND_magic_0.C D2_1 0.004759f
C2067 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q7 0.71602f
C2068 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A a_2749_2092# 0.036613f
C2069 a_5185_2253# a_5385_2253# 0.297401f
C2070 a_12387_6986# a_11191_5901# 7.51e-20
C2071 a_15865_2253# a_15865_1059# 0.005574f
C2072 a_1541_n8579# VDD 0.428164f
C2073 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_1 3.49e-19
C2074 a_8523_n3597# a_8523_n4081# 0.033537f
C2075 a_16186_n3644# a_16386_n3644# 0.300637f
C2076 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.3_inp_AND_magic_0.A 1.4e-19
C2077 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 2.34e-19
C2078 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8955_8580# 1.77e-19
C2079 a_23793_5904# 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 0.001078f
C2080 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.P3 3.85e-19
C2081 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.D 0.423451f
C2082 p2_gen_magic_0.3_inp_AND_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.238377f
C2083 OR_magic_1.VOUT divide_by_2_1.tg_magic_0.IN 0.628351f
C2084 a_11279_6341# a_8713_6842# 6.34e-20
C2085 a_11279_6341# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.03261f
C2086 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A Q3 4.82e-20
C2087 a_20041_4557# VDD 0.10656f
C2088 a_11492_n6613# D2_3 8.12e-19
C2089 a_22150_1124# VDD 1.03166f
C2090 a_12174_n3150# D2_5 0.05756f
C2091 a_14556_n3644# VDD 0.896865f
C2092 p3_gen_magic_0.AND2_magic_1.A a_12590_n7648# 0.06406f
C2093 p2_gen_magic_0.3_inp_AND_magic_0.A Q5 6.77e-20
C2094 a_5036_n3597# Q6 0.091427f
C2095 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B VDD 1.21361f
C2096 a_17405_7309# a_18891_6886# 0.002118f
C2097 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12931_6276# 9.27e-19
C2098 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.IN 0.304333f
C2099 a_4651_9163# VDD 0.051184f
C2100 a_14556_n3644# D2_1 5.58e-19
C2101 7b_counter_0.3_inp_AND_magic_0.VOUT Q3 1.6e-21
C2102 a_11492_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.00991f
C2103 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5452_n7648# 6.1e-19
C2104 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VDD 1.32065f
C2105 a_8955_3363# Q1 0.011816f
C2106 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q6 0.087309f
C2107 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_23560_3728# 0.515297f
C2108 a_1409_8579# D2_7 0.201402f
C2109 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.083376f
C2110 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.177041f
C2111 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK 1.33354f
C2112 a_1209_1059# p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 4.97e-19
C2113 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1975_n6471# 0.005701f
C2114 a_8713_6842# a_8411_4513# 1.73e-19
C2115 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT 1.98e-19
C2116 p2_gen_magic_0.xnor_magic_5.OUT a_16186_n3644# 0.229104f
C2117 OR_magic_1.VOUT divide_by_2_1.tg_magic_3.OUT 0.429603f
C2118 a_1409_1059# VDD 0.056754f
C2119 a_8643_n6024# p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 1.86e-20
C2120 p2_gen_magic_0.3_inp_AND_magic_0.A D2_4 0.006951f
C2121 7b_counter_0.MDFF_5.LD a_12931_7470# 0.033946f
C2122 a_21381_8741# Q1 0.137741f
C2123 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 2.07e-19
C2124 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.005939f
C2125 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN 0.010522f
C2126 a_21381_3524# Q6 2e-20
C2127 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.024156f
C2128 a_12387_1769# D2_6 0.261924f
C2129 7b_counter_0.MDFF_7.tspc2_magic_0.D a_27234_3319# 7.57e-20
C2130 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13769_n2115# 0.200301f
C2131 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.007087f
C2132 p2_gen_magic_0.3_inp_AND_magic_0.C Q3 0.196726f
C2133 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B D2_6 0.003901f
C2134 7b_counter_0.MDFF_0.tspc2_magic_0.D a_5515_3947# 2.1e-20
C2135 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.3_inp_AND_magic_0.C 0.226806f
C2136 a_26038_4932# D2_4 0.016305f
C2137 a_1409_2253# Q7 0.008754f
C2138 7b_counter_0.MDFF_4.LD a_27234_4513# 3.96e-19
C2139 a_1409_1059# LD 0.004065f
C2140 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A Q7 7.71e-19
C2141 p2_gen_magic_0.3_inp_AND_magic_0.C a_16386_n3644# 0.002635f
C2142 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.006652f
C2143 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 0.001326f
C2144 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B CLK 3.4e-19
C2145 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B 0.00112f
C2146 7b_counter_0.MDFF_1.tspc2_magic_0.D Q5 0.002903f
C2147 a_8411_4513# 7b_counter_0.MDFF_4.tspc2_magic_0.Q 0.243646f
C2148 a_20171_6886# VDD 0.084465f
C2149 a_15865_2253# CLK 3.82e-19
C2150 a_15865_4557# a_16065_4557# 0.29829f
C2151 a_4496_4393# a_5515_3947# 0.043767f
C2152 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.44608f
C2153 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_5 0.140212f
C2154 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 0.001081f
C2155 a_23258_575# CLK 0.042758f
C2156 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A CLK 0.002402f
C2157 a_22150_1124# Q3 0.021371f
C2158 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.01819f
C2159 a_20171_6886# D2_1 4.45e-19
C2160 OR_magic_2.A DFF_magic_0.tg_magic_3.OUT 0.007984f
C2161 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT D2_6 0.046372f
C2162 a_12387_4513# 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 1.63e-20
C2163 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q4 0.001013f
C2164 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q3 0.007775f
C2165 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_684# 0.00215f
C2166 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A D2_7 0.004847f
C2167 a_24059_4877# a_24259_4877# 0.655098f
C2168 7b_counter_0.MDFF_3.QB a_5385_7469# 2.39e-21
C2169 a_27778_3363# VDD 0.012214f
C2170 a_16386_n8142# VDD 0.024766f
C2171 7b_counter_0.MDFF_1.tspc2_magic_0.D D2_4 0.017889f
C2172 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 4e-20
C2173 a_16186_n3644# a_14756_n3644# 3.21e-19
C2174 a_14556_n3644# a_16386_n3644# 0.00107f
C2175 a_12387_575# Q4 9.11e-19
C2176 a_22062_684# a_23258_575# 0.002003f
C2177 p3_gen_magic_0.3_inp_AND_magic_0.C VDD 2.52836f
C2178 a_12387_1769# D2_2 0.002048f
C2179 a_2749_684# a_1209_1059# 0.002003f
C2180 a_6725_7308# a_8713_6842# 0.001517f
C2181 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 0.0037f
C2182 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_20041_4557# 0.001027f
C2183 a_16386_n8142# D2_1 0.004827f
C2184 a_8955_9774# D2_2 0.00581f
C2185 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.xnor_magic_5.OUT 0.006999f
C2186 a_17405_3524# 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 0.132169f
C2187 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VDD 1.25206f
C2188 p3_gen_magic_0.3_inp_AND_magic_0.C D2_1 0.281031f
C2189 a_17405_2092# VDD 0.94863f
C2190 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B VDD 1.19294f
C2191 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8955_9774# 0.128771f
C2192 a_8939_n3150# D2_5 7.68e-20
C2193 a_12174_n3597# VDD 0.18391f
C2194 a_8939_n7648# a_8523_n8095# 0.013021f
C2195 a_1409_1059# Q3 5.91e-20
C2196 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.015506f
C2197 p2_gen_magic_0.xnor_magic_0.OUT Q1 0.151292f
C2198 p3_gen_magic_0.P3 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.95e-19
C2199 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_11292_n2115# 1.86e-19
C2200 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12387_5792# 0.149276f
C2201 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B D2_1 0.005419f
C2202 a_21381_10149# VDD 1.56461f
C2203 p2_gen_magic_0.xnor_magic_3.OUT Q4 0.025387f
C2204 Q7 D2_6 0.078755f
C2205 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A Q1 0.004119f
C2206 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_9059_n1973# 6.1e-19
C2207 a_12387_4513# VDD 0.9315f
C2208 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_4235_9163# 3.22e-21
C2209 a_19841_3363# Q1 0.03068f
C2210 a_22150_1124# a_19152_1223# 0.001302f
C2211 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B D2_6 0.008142f
C2212 a_21381_3524# a_23560_3728# 0.001302f
C2213 divide_by_2_0.tg_magic_2.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 0.270406f
C2214 a_19307_6886# a_19152_5956# 0.001643f
C2215 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n1526# 0.082667f
C2216 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.003202f
C2217 p3_gen_magic_0.xnor_magic_5.OUT VDD 2.20512f
C2218 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n6471# 0.011524f
C2219 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B LD 6.05e-19
C2220 p2_gen_magic_0.xnor_magic_5.OUT a_14556_n3644# 0.047822f
C2221 a_1209_1059# VDD 0.915754f
C2222 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.NAND_magic_0.VOUT 0.785314f
C2223 p2_gen_magic_0.3_inp_AND_magic_0.VOUT D2_6 0.18848f
C2224 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q5 0.241344f
C2225 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12590_n3150# 6.1e-19
C2226 a_12931_2253# D2_6 0.180849f
C2227 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1409_4557# 0.037614f
C2228 p3_gen_magic_0.xnor_magic_5.OUT D2_1 0.003889f
C2229 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_5 0.055353f
C2230 7b_counter_0.MDFF_4.tspc2_magic_0.D Q5 0.003851f
C2231 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD 1.18054f
C2232 p2_gen_magic_0.3_inp_AND_magic_0.VOUT a_13553_n2115# 1.9e-20
C2233 a_13353_n2115# a_13769_n2115# 0.278913f
C2234 7b_counter_0.MDFF_7.tspc2_magic_0.D a_24536_3947# 0.004574f
C2235 a_13769_n2115# D2_3 0.008431f
C2236 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_27234_1769# 1.18e-19
C2237 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4651_3947# 0.004574f
C2238 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 0.168057f
C2239 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_1 0.007212f
C2240 a_5470_n6471# a_5036_n8095# 1.26e-19
C2241 a_1209_2253# Q7 0.043431f
C2242 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_16065_3363# 0.001034f
C2243 a_1209_1059# LD 0.002086f
C2244 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.B 0.003762f
C2245 p2_gen_magic_0.3_inp_AND_magic_0.C a_14756_n3644# 0.001117f
C2246 a_11279_8697# Q7 0.006685f
C2247 7b_counter_0.MDFF_5.LD VDD 21.117199f
C2248 D2_2 Q7 0.068322f
C2249 a_19841_4557# a_20041_4557# 0.29829f
C2250 a_9689_1669# Q5 0.001642f
C2251 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 9.09e-19
C2252 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT D2_6 0.116345f
C2253 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_20171_6886# 0.125951f
C2254 7b_counter_0.MDFF_4.tspc2_magic_0.D D2_4 0.002044f
C2255 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B D2_2 0.067425f
C2256 7b_counter_0.MDFF_5.LD D2_1 0.621014f
C2257 7b_counter_0.MDFF_5.tspc2_magic_0.Q Q7 0.197262f
C2258 a_19307_6886# VDD 0.003613f
C2259 7b_counter_0.MDFF_4.LD a_15865_2253# 0.224216f
C2260 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VDD 1.06646f
C2261 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT LD 1.17e-19
C2262 a_23560_3728# a_24536_3947# 0.240883f
C2263 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.05295f
C2264 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.001091f
C2265 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_2749_684# 3.58e-20
C2266 a_19841_4557# 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 1.93e-19
C2267 a_26038_684# CLK 0.006461f
C2268 a_23258_1769# Q4 1.41e-19
C2269 a_23802_1059# D2_4 0.030793f
C2270 p3_gen_magic_0.xnor_magic_0.OUT a_8523_n8095# 0.011792f
C2271 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_17405_3524# 2.07e-19
C2272 7b_counter_0.MDFF_4.LD a_23258_575# 0.001153f
C2273 a_4496_4393# a_4651_3947# 0.240883f
C2274 7b_counter_0.MDFF_6.tspc2_magic_0.Q Q1 0.457711f
C2275 a_8955_9774# CLK 4.55e-19
C2276 a_19307_6886# D2_1 9.21e-20
C2277 a_16065_1059# D2_3 0.003998f
C2278 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN D2_1 0.045993f
C2279 p2_gen_magic_0.xnor_magic_1.OUT Q7 0.192484f
C2280 a_1209_9773# D2_7 0.024506f
C2281 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A Q2 0.028159f
C2282 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26126_3480# 0.036613f
C2283 7b_counter_0.MDFF_5.LD LD 0.809257f
C2284 a_20041_3363# VDD 0.085691f
C2285 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_12387_575# 1.93e-19
C2286 p3_gen_magic_0.xnor_magic_6.OUT D2_6 0.38108f
C2287 a_14756_n8142# VDD 0.05463f
C2288 p3_gen_magic_0.AND2_magic_1.A D2_5 0.197392f
C2289 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_7 0.009795f
C2290 a_14556_n3644# a_14756_n3644# 0.300637f
C2291 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A Q6 0.326151f
C2292 a_5036_n3597# a_5036_n4081# 0.033537f
C2293 a_8643_n1526# p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 2.26e-20
C2294 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_15865_9774# 0.279825f
C2295 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.OUT 1.06e-19
C2296 p3_gen_magic_0.xnor_magic_1.OUT Q4 4.22e-19
C2297 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_0.tspc2_magic_0.Q 4.45e-20
C2298 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A Q6 0.020032f
C2299 a_12174_n7648# a_12590_n7648# 0.002223f
C2300 a_5185_1059# a_5385_1059# 0.29829f
C2301 a_8523_n3597# VDD 0.183943f
C2302 a_27234_3319# a_27234_1769# 0.003291f
C2303 a_8411_9730# a_8955_9774# 0.29829f
C2304 a_1209_1059# Q3 8.39e-19
C2305 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A Q1 0.005261f
C2306 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.237944f
C2307 Q5 D2_5 1.14544f
C2308 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_0.tspc2_magic_0.D 8.78e-21
C2309 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK 1.3249f
C2310 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VDD 1.27789f
C2311 a_11279_6341# a_12387_5792# 7.54e-20
C2312 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B p2_gen_magic_0.xnor_magic_3.OUT 1.04e-20
C2313 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n8095# 0.083086f
C2314 7b_counter_0.MDFF_5.LD a_16065_6276# 0.003068f
C2315 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n1973# 0.107246f
C2316 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3 0.626331f
C2317 a_8643_n1526# Q1 0.088603f
C2318 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A D2_1 0.001155f
C2319 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.3_inp_AND_magic_0.C 7e-19
C2320 a_17405_2092# a_19152_1223# 7.92e-19
C2321 7b_counter_0.3_inp_AND_magic_0.C CLK 0.074279f
C2322 a_12387_5792# a_12931_6276# 0.29829f
C2323 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_6725_5900# 0.414018f
C2324 p3_gen_magic_0.xnor_magic_0.OUT Q1 0.146683f
C2325 7b_counter_0.3_inp_AND_magic_0.B 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 2.65e-20
C2326 a_5036_n7648# VDD 0.044055f
C2327 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT D2_6 0.001483f
C2328 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.3_inp_AND_magic_0.VOUT 0.017858f
C2329 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q5 0.005773f
C2330 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B Q7 0.007491f
C2331 p3_gen_magic_0.xnor_magic_3.OUT Q4 0.002063f
C2332 7b_counter_0.MDFF_5.LD Q3 5.6e-19
C2333 D2_6 D2_3 0.65994f
C2334 a_13353_n2115# D2_6 0.004835f
C2335 D2_5 D2_4 0.08017f
C2336 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 0.001081f
C2337 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A LD 0.446138f
C2338 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.xnor_magic_1.OUT 0.002797f
C2339 7b_counter_0.MDFF_7.tspc2_magic_0.CLK VDD 2.28482f
C2340 p3_gen_magic_0.xnor_magic_6.OUT D2_2 5.59e-20
C2341 a_1209_3363# D2_5 0.262187f
C2342 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.3_inp_AND_magic_0.A 0.001214f
C2343 a_11191_684# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 3.58e-20
C2344 CLK Q7 0.863747f
C2345 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.001335f
C2346 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 0.006194f
C2347 7b_counter_0.MDFF_3.tspc2_magic_0.Q Q2 0.405236f
C2348 a_11292_n2115# VDD 1.12502f
C2349 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 4.5e-19
C2350 7b_counter_0.MDFF_7.tspc2_magic_0.D a_23672_3947# 2.1e-20
C2351 a_13353_n2115# a_13553_n2115# 0.522094f
C2352 a_13553_n2115# D2_3 0.002449f
C2353 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B CLK 0.005646f
C2354 a_1541_n4081# p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 1.66e-20
C2355 p3_gen_magic_0.3_inp_AND_magic_0.VOUT D2_6 0.341574f
C2356 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_23802_2253# 0.007492f
C2357 a_2749_3524# a_4651_3947# 2.34e-20
C2358 a_5054_n6471# a_5036_n8095# 2.84e-19
C2359 a_8643_n6471# a_8523_n7648# 0.186236f
C2360 a_1409_9773# a_1409_8579# 0.014163f
C2361 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 0.088975f
C2362 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q7 0.079555f
C2363 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_12387_4513# 1.39e-19
C2364 D2_7 Q5 0.419511f
C2365 Q2 D2_5 0.094726f
C2366 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_5 4.98e-19
C2367 7b_counter_0.NAND_magic_0.A 7b_counter_0.3_inp_AND_magic_0.C 0.002961f
C2368 p2_gen_magic_0.3_inp_AND_magic_0.C a_16186_n3644# 0.146469f
C2369 p2_gen_magic_0.3_inp_AND_magic_0.VOUT CLK 0.041513f
C2370 a_7303_8697# VDD 0.953498f
C2371 a_11191_10149# Q7 0.009747f
C2372 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VDD 1.18604f
C2373 a_8825_1669# Q5 0.001808f
C2374 7b_counter_0.MDFF_4.LD a_16065_2253# 0.037687f
C2375 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19307_6886# 0.069391f
C2376 a_17405_5901# VDD 1.55668f
C2377 a_8411_9730# Q7 0.02258f
C2378 a_15865_3363# a_16065_3363# 0.299584f
C2379 7b_counter_0.MDFF_1.tspc2_magic_0.CLK Q5 0.005188f
C2380 7b_counter_0.MDFF_4.LD a_12387_1769# 0.224216f
C2381 a_23560_3728# a_23672_3947# 0.043767f
C2382 p2_gen_magic_0.AND2_magic_1.A Q4 0.177246f
C2383 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_9412_5956# 0.365826f
C2384 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_1 3.85e-19
C2385 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12590_n7648# 0.005701f
C2386 7b_counter_0.MDFF_4.LD a_26038_684# 0.002672f
C2387 a_4496_9609# CLK 0.047109f
C2388 p2_gen_magic_0.xnor_magic_4.OUT Q5 0.147155f
C2389 a_15865_1059# D2_3 2.51e-19
C2390 a_5185_6275# 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7.51e-20
C2391 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.025092f
C2392 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B D2_6 0.002292f
C2393 a_1541_n3150# Q7 0.348367f
C2394 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.C 3.08e-19
C2395 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q3 0.006038f
C2396 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.160373f
C2397 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_21381_10149# 3.58e-20
C2398 D2_2 D2_3 0.099585f
C2399 D2_7 D2_4 0.936843f
C2400 a_27234_3319# VDD 0.807784f
C2401 a_16186_n8142# VDD 0.834851f
C2402 a_12387_1769# a_12931_1059# 0.003083f
C2403 a_1559_n1042# D2_7 0.017159f
C2404 a_1209_3363# D2_7 0.012171f
C2405 a_8523_n7648# D2_6 0.057124f
C2406 a_14556_n3644# a_16186_n3644# 4.95e-19
C2407 a_22150_1124# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 0.036613f
C2408 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A D2_6 0.062735f
C2409 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT CLK 0.429321f
C2410 a_27778_2253# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.001034f
C2411 7b_counter_0.MDFF_1.tspc2_magic_0.CLK D2_4 0.02577f
C2412 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B Q6 0.052906f
C2413 mux_magic_0.IN1 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 6.54e-20
C2414 a_1209_4557# Q6 0.024869f
C2415 a_16186_n8142# D2_1 0.010408f
C2416 7b_counter_0.MDFF_5.LD a_8713_6842# 0.00664f
C2417 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN D2_6 0.09995f
C2418 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 1.1e-20
C2419 p2_gen_magic_0.xnor_magic_1.OUT D2_3 0.061061f
C2420 p2_gen_magic_0.xnor_magic_4.OUT D2_4 0.002776f
C2421 a_5036_n3597# VDD 0.241656f
C2422 a_8643_n6024# Q1 0.092777f
C2423 a_20041_3363# a_19152_1223# 5.39e-19
C2424 a_32616_n2458# OUT1 7.57e-20
C2425 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_14756_n8142# 7.91e-19
C2426 a_11279_3480# Q1 0.005125f
C2427 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B Q1 1.46e-19
C2428 Q2 D2_7 2.13323f
C2429 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_2749_3524# 2.4e-20
C2430 a_4651_9163# a_5515_9163# 0.009722f
C2431 7b_counter_0.MDFF_7.tspc2_magic_0.CLK Q3 0.066474f
C2432 7b_counter_0.MDFF_5.LD a_15865_6276# 3.96e-19
C2433 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B VDD 1.1992f
C2434 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A Q1 0.002388f
C2435 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A D2_4 0.001764f
C2436 a_8643_n1973# a_8523_n3150# 0.186236f
C2437 a_11292_n2115# Q3 0.00958f
C2438 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1409_9773# 9.27e-19
C2439 a_15865_3363# Q1 0.021197f
C2440 a_12387_6986# D2_6 5.06e-20
C2441 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT 4.16e-20
C2442 a_17405_2092# a_18891_1669# 0.002118f
C2443 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_17405_8741# 2.4e-20
C2444 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_26126_3480# 0.018983f
C2445 p2_gen_magic_0.xnor_magic_4.OUT Q2 0.136949f
C2446 DFF_magic_0.D 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.007873f
C2447 a_1957_n7648# VDD 0.001798f
C2448 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B D2_2 0.064141f
C2449 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1559_n6024# 0.083665f
C2450 p2_gen_magic_0.3_inp_AND_magic_0.B D2_3 0.158244f
C2451 p2_gen_magic_0.3_inp_AND_magic_0.B a_13353_n2115# 0.385755f
C2452 p2_gen_magic_0.xnor_magic_6.OUT p2_gen_magic_0.AND2_magic_1.A 0.256454f
C2453 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 0.454908f
C2454 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT 0.710655f
C2455 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q3 0.54279f
C2456 7b_counter_0.MDFF_3.tspc2_magic_0.CLK Q6 0.003472f
C2457 a_17405_5901# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 4.22e-19
C2458 a_21381_3524# VDD 0.961727f
C2459 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_11279_8697# 2.07e-19
C2460 a_8523_n7648# D2_2 1.85e-19
C2461 a_1541_n8095# D2_7 1.21e-19
C2462 p2_gen_magic_0.xnor_magic_0.OUT a_8643_n1042# 0.298941f
C2463 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A D2_2 0.086634f
C2464 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 0.006911f
C2465 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1209_4557# 1.39e-19
C2466 Q1 Q6 0.432595f
C2467 a_4235_9163# Q2 1.57e-20
C2468 a_9212_5956# D2_6 0.056002f
C2469 7b_counter_0.MDFF_5.tspc2_magic_0.Q 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 0.27167f
C2470 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 0.001207f
C2471 mux_magic_0.IN1 OUT1 0.079149f
C2472 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.MDFF_5.LD 0.053103f
C2473 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.tspc2_magic_0.Q 0.304572f
C2474 a_5470_n1973# D2_5 0.002137f
C2475 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT CLK 0.329619f
C2476 7b_counter_0.MDFF_5.LD a_16065_9774# 0.033901f
C2477 DFF_magic_0.tg_magic_3.OUT P2 3.51e-19
C2478 a_4235_3947# Q7 0.0116f
C2479 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B Q6 3.81e-19
C2480 a_13353_n2115# CLK 0.001356f
C2481 p2_gen_magic_0.3_inp_AND_magic_0.C a_14556_n3644# 5.23e-19
C2482 7b_counter_0.MDFF_4.LD p2_gen_magic_0.3_inp_AND_magic_0.VOUT 5.18e-20
C2483 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 9.4e-20
C2484 CLK D2_3 1.61325f
C2485 a_11292_n6613# VDD 1.12545f
C2486 a_23207_5885# Q4 0.018848f
C2487 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VDD 1.18701f
C2488 7b_counter_0.MDFF_4.LD a_12931_2253# 0.037687f
C2489 a_11492_n6613# a_11708_n6613# 0.329078f
C2490 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_5901# 0.00215f
C2491 a_12387_6986# D2_2 0.268168f
C2492 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A CLK 7.36e-19
C2493 a_11292_n6613# D2_1 0.009796f
C2494 a_26126_3480# a_27234_3319# 0.001529f
C2495 a_12387_5792# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 1.27e-19
C2496 a_22062_684# p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 1.69e-19
C2497 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 3.27e-20
C2498 a_23258_1769# a_23258_575# 0.005574f
C2499 a_15865_9774# CLK 0.243646f
C2500 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A a_1409_3363# 1.77e-19
C2501 p3_gen_magic_0.3_inp_AND_magic_0.VOUT CLK 0.346875f
C2502 7b_counter_0.MDFF_5.LD 7b_counter_0.3_inp_AND_magic_0.B 7.88e-20
C2503 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B a_6725_2092# 0.428787f
C2504 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.856654f
C2505 7b_counter_0.DFF_magic_0.tg_magic_2.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.270406f
C2506 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 3.17e-19
C2507 a_12931_2253# a_12931_1059# 0.020635f
C2508 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n7648# 0.107246f
C2509 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A D2_6 0.002966f
C2510 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_24059_4877# 3.22e-21
C2511 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.178114f
C2512 a_12387_1769# a_12387_575# 0.005574f
C2513 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_17405_10149# 0.414018f
C2514 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q3 2.94e-19
C2515 a_24536_3947# VDD 0.004521f
C2516 a_14556_n8142# VDD 0.877977f
C2517 a_12174_n7648# D2_5 0.081565f
C2518 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 0.178114f
C2519 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B CLK 0.075385f
C2520 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 6.76e-19
C2521 a_5036_n8095# Q6 0.089626f
C2522 a_9689_6886# Q2 0.030174f
C2523 a_1559_n6024# a_1957_n7648# 3.01e-19
C2524 p3_gen_magic_0.xnor_magic_4.OUT Q5 0.477574f
C2525 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n4081# 0.093592f
C2526 DFF_magic_0.tg_magic_3.OUT VDD 1.1675f
C2527 p3_gen_magic_0.xnor_magic_5.OUT a_5036_n8579# 0.426478f
C2528 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_21381_4932# 0.414018f
C2529 a_12590_n3150# VDD 0.001798f
C2530 a_8713_1625# D2_6 0.025758f
C2531 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.xnor_magic_6.OUT 0.199228f
C2532 a_5470_n1973# D2_7 6.9e-19
C2533 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B CLK 0.003598f
C2534 a_11191_4932# Q1 0.002146f
C2535 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.035743f
C2536 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.005351f
C2537 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q4 0.002221f
C2538 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_2749_4932# 3.58e-20
C2539 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22062_684# 0.189314f
C2540 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.001091f
C2541 a_8955_3363# a_8825_1669# 0.005699f
C2542 a_21381_3524# Q3 0.158586f
C2543 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT DFF_magic_0.tg_magic_2.OUT 0.168057f
C2544 7b_counter_0.MDFF_5.LD a_12931_6276# 0.001799f
C2545 a_5385_2253# VDD 0.109264f
C2546 a_26126_1124# D2_4 0.024037f
C2547 7b_counter_0.MDFF_3.QB D2_7 0.298558f
C2548 a_1209_9773# a_1409_9773# 0.29829f
C2549 a_9412_739# D2_6 0.012302f
C2550 a_12387_3319# Q1 0.021245f
C2551 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A CLK 0.00246f
C2552 p2_gen_magic_0.xnor_magic_1.OUT a_13353_n6613# 1.35e-19
C2553 p3_gen_magic_0.xnor_magic_4.OUT D2_4 0.207572f
C2554 a_16065_4557# Q2 0.128771f
C2555 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_9059_n6471# 0.005701f
C2556 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_24259_4877# 0.365826f
C2557 a_17405_5901# a_15865_6276# 0.002003f
C2558 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN D2_4 0.004512f
C2559 a_8523_n4081# Q1 0.007197f
C2560 p2_gen_magic_0.xnor_magic_4.OUT a_5470_n1973# 0.077238f
C2561 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN CLK 0.001049f
C2562 p2_gen_magic_0.xnor_magic_5.OUT a_5036_n3597# 0.3716f
C2563 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11279_8697# 0.036613f
C2564 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A D2_2 0.001793f
C2565 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_6 0.030321f
C2566 a_5185_7469# 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B 0.146237f
C2567 a_5385_2253# LD 0.036926f
C2568 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT P2 4.95e-19
C2569 DFF_magic_0.D 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.011018f
C2570 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A D2_5 0.002851f
C2571 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.202081f
C2572 p3_gen_magic_0.xnor_magic_4.OUT Q2 0.131678f
C2573 a_12387_6986# CLK 0.031838f
C2574 a_8411_9730# 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 0.279825f
C2575 p3_gen_magic_0.3_inp_AND_magic_0.B D2_3 0.007212f
C2576 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q7 0.003321f
C2577 7b_counter_0.MDFF_3.QB a_4235_9163# 0.027775f
C2578 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK 0.012402f
C2579 a_8643_n1042# a_8643_n1526# 0.033537f
C2580 7b_counter_0.MDFF_5.tspc2_magic_0.CLK Q7 0.00429f
C2581 a_5054_n1973# D2_5 0.075944f
C2582 a_7215_10149# a_8411_8536# 7.51e-20
C2583 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT 6.94e-19
C2584 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 0.002343f
C2585 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_5 0.134312f
C2586 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_8411_8536# 0.001985f
C2587 a_24536_3947# Q3 0.001018f
C2588 7b_counter_0.MDFF_4.LD D2_3 0.902721f
C2589 7b_counter_0.MDFF_4.LD a_13353_n2115# 9.33e-19
C2590 a_22991_5885# Q4 0.006975f
C2591 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3 1.02284f
C2592 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_4235_3947# 7.16e-19
C2593 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.3_inp_AND_magic_0.VOUT 0.023253f
C2594 a_9412_739# D2_2 1.68e-20
C2595 7b_counter_0.MDFF_5.tspc2_magic_0.D Q2 0.108645f
C2596 a_12387_3319# a_12931_3363# 0.299584f
C2597 a_12387_5792# a_12387_4513# 0.005698f
C2598 DFF_magic_0.tg_magic_3.OUT Q3 3.73e-19
C2599 a_9212_5956# CLK 0.003549f
C2600 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 0.007053f
C2601 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1957_n3150# 6.85e-21
C2602 a_26126_3480# a_24536_3947# 2.34e-20
C2603 a_12174_n3150# Q4 0.372511f
C2604 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 0.001214f
C2605 7b_counter_0.MDFF_1.tspc2_magic_0.Q VDD 1.15267f
C2606 a_2749_2092# a_2749_684# 0.479729f
C2607 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_5185_7469# 4.65e-19
C2608 a_13353_n6613# CLK 0.001331f
C2609 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VDD 1.08434f
C2610 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23560_3728# 0.012992f
C2611 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 0.005763f
C2612 p2_gen_magic_0.xnor_magic_3.OUT Q7 0.09063f
C2613 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.09196f
C2614 DFF_magic_0.tg_magic_2.OUT CLK 0.303257f
C2615 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_2 0.05482f
C2616 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.MDFF_5.LD 0.102172f
C2617 a_16065_7470# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 1.77e-19
C2618 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VDD 1.31445f
C2619 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_4235_3947# 5.64e-20
C2620 a_12174_n8095# VDD 0.18391f
C2621 a_8939_n7648# D2_5 0.00143f
C2622 a_23672_3947# VDD 0.089802f
C2623 a_1209_9773# 7b_counter_0.MDFF_3.tspc2_magic_0.D 1.63e-20
C2624 7b_counter_0.NAND_magic_0.A 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.95e-19
C2625 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_2749_8740# 0.036613f
C2626 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT D2_1 0.001753f
C2627 7b_counter_0.MDFF_4.tspc2_magic_0.Q 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B 4.45e-20
C2628 a_21504_5904# Q1 0.048507f
C2629 p2_gen_magic_0.xnor_magic_5.OUT a_11292_n6613# 6.92e-21
C2630 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B 9.09e-19
C2631 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VDD 1.25654f
C2632 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A D2_1 5.31e-20
C2633 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A D2_7 0.00417f
C2634 a_2749_7308# Q6 0.009259f
C2635 a_8825_6886# Q2 0.002191f
C2636 a_27234_1769# a_27778_1059# 0.003083f
C2637 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A D2_5 0.092291f
C2638 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.164969f
C2639 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_4 0.004858f
C2640 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.3_inp_AND_magic_0.VOUT 1.64e-19
C2641 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A Q1 0.004356f
C2642 a_19841_4557# a_21381_3524# 7.54e-20
C2643 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 0.003022f
C2644 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A Q4 4.99e-19
C2645 a_5054_n1973# D2_7 0.495733f
C2646 a_23672_3947# a_23802_2253# 0.005699f
C2647 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_14556_n8142# 0.008174f
C2648 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 0.004701f
C2649 7b_counter_0.MDFF_1.tspc2_magic_0.D 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 8.78e-21
C2650 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8939_n7648# 6.1e-19
C2651 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_4.OUT 0.349856f
C2652 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A CLK 0.006122f
C2653 7b_counter_0.3_inp_AND_magic_0.C a_24401_7877# 0.057f
C2654 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A LD 0.445809f
C2655 7b_counter_0.MDFF_5.LD a_12387_5792# 3.96e-19
C2656 a_2749_2092# VDD 0.947759f
C2657 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19841_3363# 4.65e-19
C2658 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT a_27234_4513# 0.005873f
C2659 a_12387_4513# 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 0.279825f
C2660 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n6471# 0.006378f
C2661 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_24059_4877# 0.671058f
C2662 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A LD 0.001147f
C2663 p2_gen_magic_0.xnor_magic_4.OUT a_5054_n1973# 0.300596f
C2664 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_7303_3480# 0.001342f
C2665 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q2 0.001508f
C2666 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.00222f
C2667 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.002118f
C2668 p2_gen_magic_0.xnor_magic_6.OUT a_12174_n3150# 0.143718f
C2669 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_11191_10149# 0.414018f
C2670 a_5036_n3150# a_5036_n3597# 0.014233f
C2671 VDD OUT1 0.34986f
C2672 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n8579# 0.066064f
C2673 a_5185_7469# a_5385_7469# 0.297401f
C2674 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_2749_7308# 0.036613f
C2675 a_5054_n6471# D2_5 0.079228f
C2676 a_19841_8580# Q7 8.99e-19
C2677 a_2749_2092# LD 0.001152f
C2678 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4 0.686515f
C2679 a_1409_9773# Q2 6.99e-19
C2680 a_5185_2253# D2_5 0.253539f
C2681 a_1209_1059# a_1409_1059# 0.29829f
C2682 7b_counter_0.MDFF_3.QB a_4496_10093# 3.52e-19
C2683 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.003129f
C2684 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_6 2.08e-19
C2685 7b_counter_0.MDFF_7.tspc2_magic_0.D a_26038_4932# 1.08e-19
C2686 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B Q7 7.61e-19
C2687 a_7303_8697# a_5515_9163# 3.09e-20
C2688 a_11191_684# a_11292_n2115# 7.67e-20
C2689 a_12174_n8095# a_12174_n8579# 0.033537f
C2690 p3_gen_magic_0.xnor_magic_0.OUT D2_5 0.171896f
C2691 a_23672_3947# Q3 9.38e-19
C2692 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 1.19e-19
C2693 p3_gen_magic_0.3_inp_AND_magic_0.C a_16386_n8142# 0.002635f
C2694 a_9212_739# Q5 0.007724f
C2695 p3_gen_magic_0.xnor_magic_1.OUT Q7 0.1574f
C2696 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n3597# 0.083665f
C2697 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_4496_4877# 1.29e-19
C2698 a_1209_6275# a_1409_6275# 0.29829f
C2699 p3_gen_magic_0.3_inp_AND_magic_0.B a_13353_n6613# 0.385755f
C2700 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A D2_3 0.00207f
C2701 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A D2_3 0.001346f
C2702 a_24259_4877# a_24536_3947# 0.001643f
C2703 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.tspc2_magic_0.Q 4.46e-19
C2704 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27778_3363# 1.77e-19
C2705 p3_gen_magic_0.xnor_magic_0.OUT a_8643_n5540# 0.298941f
C2706 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 1.42966f
C2707 a_12387_575# D2_3 3.32e-19
C2708 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7303_8697# 0.431521f
C2709 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_2.OUT 1.09743f
C2710 a_27778_1059# VDD 0.056754f
C2711 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.018819f
C2712 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_3 1.02771f
C2713 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B a_27234_4513# 1.93e-19
C2714 a_16065_3363# VDD 0.018978f
C2715 a_8523_n8095# VDD 0.183943f
C2716 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_19841_3363# 0.001158f
C2717 a_5054_n6471# D2_7 1.85e-19
C2718 a_1209_9773# a_2749_8740# 7.54e-20
C2719 a_9212_739# D2_4 2.51e-20
C2720 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_2749_10148# 0.414018f
C2721 a_19152_5956# Q1 1.39e-19
C2722 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B VDD 1.21691f
C2723 a_1209_4557# VDD 0.931274f
C2724 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19152_1223# 0.012895f
C2725 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_7215_4932# 0.189314f
C2726 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 0.178114f
C2727 a_11191_5901# D2_6 0.004909f
C2728 a_7303_8697# a_6725_7308# 1.62e-19
C2729 p3_gen_magic_0.xnor_magic_5.OUT a_16386_n8142# 0.037687f
C2730 7b_counter_0.MDFF_4.tspc2_magic_0.CLK Q1 0.045345f
C2731 p3_gen_magic_0.xnor_magic_3.OUT Q7 6.24e-19
C2732 a_11292_n2115# p2_gen_magic_0.3_inp_AND_magic_0.C 2.24e-19
C2733 p2_gen_magic_0.xnor_magic_3.OUT D2_3 0.081186f
C2734 p2_gen_magic_0.xnor_magic_3.OUT a_13353_n2115# 0.001977f
C2735 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.OUT 0.015247f
C2736 a_11279_1124# Q1 0.010291f
C2737 a_12931_9774# CLK 0.00442f
C2738 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_2 0.079116f
C2739 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.xnor_magic_5.OUT 0.006999f
C2740 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 8.78e-21
C2741 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12174_n8095# 0.063777f
C2742 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q4 2.74e-19
C2743 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD 1.03835f
C2744 7b_counter_0.3_inp_AND_magic_0.C a_24185_7877# 0.001361f
C2745 7b_counter_0.MDFF_5.LD a_20171_6886# 8.49e-19
C2746 7b_counter_0.MDFF_3.tspc2_magic_0.D Q2 0.001097f
C2747 a_32616_n1264# OUT1 1.63e-20
C2748 p3_gen_magic_0.3_inp_AND_magic_0.B a_13769_n6613# 0.121479f
C2749 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q7 0.007952f
C2750 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_1 3.57e-19
C2751 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8955_8580# 5.46e-20
C2752 a_8411_3319# Q1 0.020203f
C2753 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 2.29e-19
C2754 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.3_inp_AND_magic_0.A 3.14e-20
C2755 a_1209_4557# LD 0.00142f
C2756 a_19307_6886# a_20171_6886# 0.009722f
C2757 p2_gen_magic_0.xnor_magic_4.OUT a_8643_n1526# 2.24e-19
C2758 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1409_1059# 0.037614f
C2759 p3_gen_magic_0.xnor_magic_4.OUT a_5470_n6471# 0.077238f
C2760 7b_counter_0.MDFF_0.tspc2_magic_0.D Q7 0.01055f
C2761 p2_gen_magic_0.xnor_magic_6.OUT a_8939_n3150# 0.06406f
C2762 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 0.003149f
C2763 7b_counter_0.MDFF_4.LD a_8713_1625# 0.00664f
C2764 7b_counter_0.MDFF_3.tspc2_magic_0.CLK VDD 2.45781f
C2765 DFF_magic_0.tg_magic_3.OUT DFF_magic_0.tg_magic_0.IN 0.859117f
C2766 VDD Q1 6.49757f
C2767 a_8643_n6024# D2_5 0.004188f
C2768 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.054307f
C2769 7b_counter_0.MDFF_3.tspc2_magic_0.CLK D2_1 0.042272f
C2770 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_19841_4557# 0.243646f
C2771 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A Q2 0.002785f
C2772 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_5385_6275# 9.27e-19
C2773 Q1 D2_1 1.88945f
C2774 a_11708_n6613# D2_2 1.63e-20
C2775 a_11191_5901# D2_2 0.044054f
C2776 a_4496_4393# Q7 0.057609f
C2777 7b_counter_0.MDFF_3.QB a_1409_9773# 0.130365f
C2778 a_19841_9774# Q7 0.050778f
C2779 a_27778_1059# Q3 0.155139f
C2780 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B VDD 1.19144f
C2781 a_8643_n5540# a_8643_n6024# 0.033537f
C2782 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1209_3363# 0.001158f
C2783 p3_gen_magic_0.AND2_magic_1.A Q4 0.467693f
C2784 7b_counter_0.MDFF_5.LD a_21381_10149# 0.006057f
C2785 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_12387_6986# 5.28e-20
C2786 a_7215_4932# Q7 0.020007f
C2787 7b_counter_0.MDFF_3.tspc2_magic_0.CLK LD 0.087022f
C2788 a_14756_n8142# a_16386_n8142# 0.003333f
C2789 7b_counter_0.MDFF_5.tspc2_magic_0.D 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 2.05e-19
C2790 a_1209_1059# p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT 4.61e-20
C2791 a_12174_n4081# D2_5 0.027082f
C2792 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A Q7 0.017326f
C2793 a_19841_8580# D2_3 0.003016f
C2794 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.04e-19
C2795 OR_magic_1.VOUT divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT 0.005192f
C2796 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT mux_magic_0.AND2_magic_0.A 4.32e-20
C2797 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5385_1059# 0.128771f
C2798 a_8643_n6024# p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 2.26e-20
C2799 7b_counter_0.MDFF_3.tspc2_magic_0.Q Q6 0.15616f
C2800 LD Q1 0.00361f
C2801 p3_gen_magic_0.3_inp_AND_magic_0.C a_14756_n8142# 0.00228f
C2802 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B D2_1 3.46e-19
C2803 a_1541_n7648# Q7 0.306674f
C2804 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.0041f
C2805 a_24059_4877# a_24536_3947# 0.16113f
C2806 a_5185_6275# a_4496_4393# 2.33e-20
C2807 a_16065_7470# 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.001034f
C2808 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B D2_3 5.05e-19
C2809 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.05295f
C2810 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A Q2 0.098653f
C2811 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5054_n1042# 6.91e-20
C2812 Q6 D2_5 1.17252f
C2813 Q4 Q5 5.11597f
C2814 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_684# 0.189314f
C2815 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_6.tspc2_magic_0.D 0.001711f
C2816 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_9212_5956# 0.671058f
C2817 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B LD 6.07e-19
C2818 a_15865_2253# a_17405_684# 7.51e-20
C2819 a_15865_9774# a_17405_10149# 0.002003f
C2820 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A D2_4 0.012613f
C2821 a_12931_3363# VDD 0.012214f
C2822 a_5036_n8095# VDD 0.240773f
C2823 a_1209_9773# a_2749_10148# 0.002003f
C2824 a_5385_7469# VDD 0.108951f
C2825 a_15865_9774# 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 1.93e-19
C2826 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_18891_1669# 1.94e-20
C2827 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 0.178114f
C2828 a_23258_1769# 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B 0.146237f
C2829 7b_counter_0.MDFF_7.tspc2_magic_0.Q VDD 1.19031f
C2830 a_15865_2253# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 0.001985f
C2831 p3_gen_magic_0.xnor_magic_5.OUT a_14756_n8142# 0.028482f
C2832 a_17405_4932# Q1 0.002146f
C2833 a_6725_2092# Q1 0.017059f
C2834 a_1209_8579# CLK 0.020048f
C2835 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B Q1 0.013345f
C2836 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_19841_8580# 0.001985f
C2837 Q4 D2_4 0.741648f
C2838 a_6725_684# Q7 8.78e-19
C2839 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5 1.05482f
C2840 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_16065_4557# 0.037614f
C2841 a_1559_n1042# Q4 6.99e-20
C2842 Q1 Q3 0.18695f
C2843 divide_by_2_1.tg_magic_3.OUT P2 3.4e-19
C2844 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23802_2253# 0.016967f
C2845 divide_by_2_1.tg_magic_0.IN VDD 1.02232f
C2846 7b_counter_0.3_inp_AND_magic_0.C a_23207_5885# 0.645415f
C2847 mux_magic_0.AND2_magic_0.A OUT1 8.78e-21
C2848 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VDD 1.25834f
C2849 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_15865_3363# 1.18e-19
C2850 p3_gen_magic_0.3_inp_AND_magic_0.B a_13553_n6613# 0.175285f
C2851 a_5385_7469# LD 0.036926f
C2852 p3_gen_magic_0.xnor_magic_3.OUT D2_3 0.134398f
C2853 a_5054_n1973# p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.002715f
C2854 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 0.0037f
C2855 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.tspc2_magic_0.D 0.003457f
C2856 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A D2_1 0.002134f
C2857 a_21381_3524# a_22150_1124# 7.9e-19
C2858 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_2749_5900# 3.58e-20
C2859 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A a_1209_1059# 0.279825f
C2860 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A Q7 0.032975f
C2861 Q2 Q4 0.026955f
C2862 D2_7 Q6 0.999948f
C2863 p3_gen_magic_0.xnor_magic_4.OUT a_5054_n6471# 0.30189f
C2864 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_3524# 0.431521f
C2865 a_27234_1769# a_27234_575# 0.005574f
C2866 a_2749_3524# Q7 0.020941f
C2867 a_8523_n3150# a_8939_n3150# 0.002223f
C2868 a_2749_5900# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 1.52e-21
C2869 a_23207_5885# Q7 2.42e-19
C2870 7b_counter_0.MDFF_6.tspc2_magic_0.CLK Q1 0.086115f
C2871 p2_gen_magic_0.xnor_magic_6.OUT Q5 0.153944f
C2872 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 3.73e-20
C2873 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_0.tspc2_magic_0.D 0.001711f
C2874 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q5 1.35e-19
C2875 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT 1.64e-19
C2876 a_5036_n7648# p3_gen_magic_0.xnor_magic_5.OUT 0.09365f
C2877 p3_gen_magic_0.xnor_magic_1.OUT a_8523_n7648# 4.75e-19
C2878 a_1541_n3597# Q7 0.090996f
C2879 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN D2_6 0.109473f
C2880 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A a_5185_6275# 0.149276f
C2881 p2_gen_magic_0.xnor_magic_4.OUT Q6 0.010076f
C2882 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_4.OUT 0.348279f
C2883 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_9059_n1973# 0.005701f
C2884 a_11492_n6613# D2_2 2.63e-20
C2885 divide_by_2_1.tg_magic_3.OUT VDD 1.16422f
C2886 7b_counter_0.MDFF_3.QB a_7215_10149# 1.88e-20
C2887 a_19152_1223# Q1 0.039491f
C2888 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_0.tspc2_magic_0.D 2.05e-19
C2889 a_27234_3319# a_27778_3363# 0.299584f
C2890 divide_by_2_1.tg_magic_3.OUT D2_1 9.28e-21
C2891 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 4.63e-20
C2892 a_8523_n4081# D2_5 0.007824f
C2893 a_16186_n8142# a_16386_n8142# 0.300637f
C2894 a_8523_n8095# a_8523_n8579# 0.033537f
C2895 p2_gen_magic_0.AND2_magic_1.A D2_3 0.108856f
C2896 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5185_1059# 0.243646f
C2897 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_4 2.86e-19
C2898 p2_gen_magic_0.xnor_magic_5.OUT Q1 0.030344f
C2899 p3_gen_magic_0.3_inp_AND_magic_0.C a_16186_n8142# 0.146469f
C2900 a_1559_n6471# p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.002741f
C2901 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q5 0.00736f
C2902 a_8643_n6471# a_9059_n6471# 5.82e-19
C2903 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_16065_6276# 9.27e-19
C2904 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n1042# 0.093592f
C2905 a_24059_4877# a_23672_3947# 0.007202f
C2906 p2_gen_magic_0.3_inp_AND_magic_0.A VDD 1.2488f
C2907 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q3 0.478529f
C2908 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A D2_7 0.001764f
C2909 a_19841_9774# D2_3 0.002956f
C2910 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27234_3319# 0.001985f
C2911 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_15865_8580# 0.001985f
C2912 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B Q5 0.002371f
C2913 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_4932# 1.51e-21
C2914 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q7 0.002473f
C2915 a_20171_1669# D2_3 4.45e-19
C2916 p2_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.3_inp_AND_magic_0.VOUT 9.58e-20
C2917 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A a_4496_4393# 2.53e-19
C2918 a_12590_n7648# VDD 0.001798f
C2919 a_27234_4513# D2_4 0.004348f
C2920 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_4 2.45e-19
C2921 a_2749_7308# VDD 0.947759f
C2922 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_2.IN 6.95e-19
C2923 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_1209_2253# 1.18e-19
C2924 a_16065_2253# 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 1.77e-19
C2925 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_6 0.044215f
C2926 a_26038_4932# VDD 1.56756f
C2927 a_9059_n6471# D2_6 1.05e-19
C2928 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B D2_4 0.01395f
C2929 a_19841_4557# Q1 0.013976f
C2930 p3_gen_magic_0.xnor_magic_5.OUT a_16186_n8142# 0.229104f
C2931 a_1559_n1973# D2_7 0.004321f
C2932 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.008398f
C2933 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A D2_4 5.7e-19
C2934 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5185_7469# 0.029386f
C2935 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A CLK 0.029356f
C2936 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A Q1 8.6e-19
C2937 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.0037f
C2938 7b_counter_0.MDFF_4.tspc2_magic_0.Q Q1 0.154085f
C2939 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C2940 a_27234_575# VDD 0.91602f
C2941 7b_counter_0.3_inp_AND_magic_0.C a_22991_5885# 0.019083f
C2942 a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 0.149276f
C2943 a_17405_10149# a_17405_8741# 0.479729f
C2944 p3_gen_magic_0.3_inp_AND_magic_0.B a_11708_n6613# 0.002716f
C2945 a_16065_4557# a_15865_3363# 0.003083f
C2946 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_8741# 0.431521f
C2947 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A Q2 0.050944f
C2948 a_2749_7308# LD 0.001152f
C2949 a_1209_2253# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B 0.146237f
C2950 a_22062_684# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 3.58e-20
C2951 a_6725_684# D2_3 2.92e-20
C2952 p3_gen_magic_0.xnor_magic_4.OUT a_8643_n6024# 2.24e-19
C2953 a_1409_6275# CLK 0.003964f
C2954 a_19841_8580# a_19152_6440# 3.03e-19
C2955 7b_counter_0.MDFF_1.tspc2_magic_0.D VDD 1.40894f
C2956 a_2749_4932# Q7 0.002541f
C2957 a_22991_5885# Q7 3.88e-19
C2958 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8643_n1042# 3.85e-20
C2959 a_16065_9774# Q1 5.64e-20
C2960 a_8523_n3150# Q5 0.307379f
C2961 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_3524# 0.431521f
C2962 p3_gen_magic_0.xnor_magic_3.OUT a_13353_n6613# 0.001977f
C2963 a_11292_n6613# p3_gen_magic_0.3_inp_AND_magic_0.C 2.24e-19
C2964 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n8095# 0.063576f
C2965 p2_gen_magic_0.3_inp_AND_magic_0.A Q3 0.003395f
C2966 a_13769_n2115# D2_6 5.08e-20
C2967 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n1973# 0.009408f
C2968 a_9059_n6471# D2_2 0.005701f
C2969 a_5185_1059# p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 4.61e-20
C2970 a_18891_1669# Q1 0.005605f
C2971 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_5385_1059# 8.53e-19
C2972 a_5054_n1526# D2_5 0.050707f
C2973 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 0.001081f
C2974 7b_counter_0.3_inp_AND_magic_0.B Q1 0.058399f
C2975 a_1409_3363# D2_5 0.17951f
C2976 a_12174_n7648# Q4 0.307963f
C2977 a_13553_n2115# a_13769_n2115# 0.329078f
C2978 a_5036_n4081# D2_5 0.050292f
C2979 a_16186_n8142# a_14756_n8142# 3.21e-19
C2980 a_14556_n8142# a_16386_n8142# 0.00107f
C2981 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_20041_4557# 0.128771f
C2982 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q5 0.003756f
C2983 p3_gen_magic_0.3_inp_AND_magic_0.C a_14556_n8142# 5.36e-19
C2984 7b_counter_0.DFF_magic_0.tg_magic_1.IN CLK 0.857164f
C2985 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_22150_1124# 6.72e-19
C2986 a_23985_7877# Q4 7.55e-20
C2987 p3_gen_magic_0.xnor_magic_4.OUT Q6 0.121503f
C2988 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5452_n3150# 7.77e-21
C2989 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_16065_8580# 1.77e-19
C2990 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_15865_6276# 0.149276f
C2991 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B Q5 0.002223f
C2992 a_8643_n1042# VDD 0.38659f
C2993 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.tspc2_magic_0.D 0.40025f
C2994 a_5185_7469# D2_7 0.243646f
C2995 a_11279_1124# 7b_counter_0.MDFF_4.tspc2_magic_0.D 0.134004f
C2996 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN CLK 0.628351f
C2997 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.249077f
C2998 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.015727f
C2999 a_19307_1669# D2_3 0.007464f
C3000 p2_gen_magic_0.AND2_magic_1.A a_13353_n6613# 3.45e-20
C3001 a_26038_4932# a_26126_3480# 0.479729f
C3002 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B Q7 0.079471f
C3003 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_4 1.59e-20
C3004 a_27234_575# Q3 0.270357f
C3005 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C3006 a_1559_n6471# D2_7 4.11e-19
C3007 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.16497f
C3008 p3_gen_magic_0.3_inp_AND_magic_0.A VDD 1.25088f
C3009 a_12590_n3150# a_12174_n3597# 0.013021f
C3010 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.VOUT 9.99e-20
C3011 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A Q7 0.023977f
C3012 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_9689_1669# 0.069391f
C3013 a_11279_1124# a_9689_1669# 2.34e-20
C3014 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B D2_4 0.013873f
C3015 a_1209_8579# a_1209_7469# 0.003291f
C3016 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.tspc2_magic_0.Q 0.018858f
C3017 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD 1.17931f
C3018 p3_gen_magic_0.3_inp_AND_magic_0.A D2_1 0.003522f
C3019 a_8643_n6471# D2_6 1.85e-19
C3020 7b_counter_0.NAND_magic_0.A 7b_counter_0.DFF_magic_0.tg_magic_1.IN 8.34e-19
C3021 p3_gen_magic_0.xnor_magic_5.OUT a_14556_n8142# 0.050614f
C3022 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VDD 1.38534f
C3023 a_15865_2253# D2_4 0.002007f
C3024 7b_counter_0.MDFF_1.tspc2_magic_0.D Q3 2.79e-19
C3025 p2_gen_magic_0.xnor_magic_3.OUT a_5054_n1042# 0.128084f
C3026 a_23258_575# D2_4 0.029476f
C3027 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B CLK 0.002402f
C3028 a_5054_n1526# D2_7 1.66e-20
C3029 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.006184f
C3030 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.435469f
C3031 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT a_12590_n7648# 6.1e-19
C3032 a_19152_739# CLK 4.53e-22
C3033 a_1409_3363# D2_7 0.009158f
C3034 7b_counter_0.MDFF_4.tspc2_magic_0.D VDD 1.40761f
C3035 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_27234_3319# 5.28e-20
C3036 a_5036_n4081# D2_7 0.007723f
C3037 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A D2_1 0.012638f
C3038 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.001228f
C3039 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 0.005351f
C3040 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q2 7.53e-21
C3041 a_8411_8536# Q7 3.67e-19
C3042 p2_gen_magic_0.xnor_magic_0.OUT Q4 0.027739f
C3043 a_8411_4513# Q1 8.5e-19
C3044 a_23802_1059# VDD 0.098144f
C3045 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q4 0.003415f
C3046 a_21381_4932# a_19841_3363# 7.51e-20
C3047 p3_gen_magic_0.3_inp_AND_magic_0.B a_11492_n6613# 7.27e-19
C3048 a_7303_3480# a_4496_4393# 0.001527f
C3049 a_1209_2253# a_1409_2253# 0.299584f
C3050 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_1209_6275# 1.93e-19
C3051 a_1409_7469# a_1409_6275# 0.020635f
C3052 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_7 0.150658f
C3053 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 8.02e-19
C3054 a_15865_1059# a_16065_1059# 0.29829f
C3055 p2_gen_magic_0.xnor_magic_4.OUT a_5054_n1526# 0.418635f
C3056 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK 0.005192f
C3057 a_7215_4932# a_7303_3480# 0.479729f
C3058 a_19841_3363# Q4 2.73e-20
C3059 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7303_3480# 0.036613f
C3060 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_27234_575# 1.93e-19
C3061 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_5515_9163# 0.125951f
C3062 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT Q4 0.68866f
C3063 a_9689_1669# VDD 0.003613f
C3064 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_7308# 0.431521f
C3065 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A Q2 7.6e-19
C3066 a_2749_684# D2_5 0.002918f
C3067 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_2749_4932# 0.189314f
C3068 a_5515_3947# Q6 0.00148f
C3069 a_5054_n6024# D2_5 0.040424f
C3070 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_11191_5901# 8.42e-19
C3071 p2_gen_magic_0.3_inp_AND_magic_0.B a_13769_n2115# 0.121479f
C3072 7b_counter_0.MDFF_1.tspc2_magic_0.D a_19152_1223# 0.038362f
C3073 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A Q1 0.002388f
C3074 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6 0.672068f
C3075 a_8643_n6471# D2_2 0.054067f
C3076 a_11191_684# Q1 0.001194f
C3077 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_16065_6276# 0.037614f
C3078 DFF_magic_0.D DFF_magic_0.tg_magic_2.OUT 0.06125f
C3079 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_5185_1059# 0.149276f
C3080 7b_counter_0.MDFF_3.tspc2_magic_0.Q VDD 1.38715f
C3081 a_12174_n3150# D2_3 6.39e-19
C3082 a_5036_n8095# a_5036_n8579# 0.033537f
C3083 a_14556_n8142# a_14756_n8142# 0.300637f
C3084 7b_counter_0.3_inp_AND_magic_0.VOUT Q1 1.62e-19
C3085 7b_counter_0.MDFF_6.tspc2_magic_0.D a_19152_5956# 0.120019f
C3086 a_1559_n6024# p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 6.69e-21
C3087 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.006453f
C3088 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q4 0.001089f
C3089 7b_counter_0.MDFF_3.tspc2_magic_0.Q D2_1 0.001093f
C3090 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.148797f
C3091 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.166749f
C3092 a_27234_1769# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.001985f
C3093 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q3 0.001438f
C3094 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.025092f
C3095 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n3150# 0.008799f
C3096 VDD D2_5 4.68562f
C3097 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT a_1957_n7648# 1.46e-20
C3098 a_12387_1769# Q5 3.88e-19
C3099 a_15865_1059# D2_6 3.54e-19
C3100 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_24059_4877# 1.94e-20
C3101 a_11279_8697# D2_6 0.012746f
C3102 7b_counter_0.MDFF_4.tspc2_magic_0.D Q3 4.06e-19
C3103 D2_2 D2_6 3.10857f
C3104 D2_1 D2_5 1.73888f
C3105 7b_counter_0.MDFF_7.tspc2_magic_0.Q 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 0.002402f
C3106 7b_counter_0.MDFF_3.tspc2_magic_0.Q LD 0.121479f
C3107 a_5185_1059# p2_gen_magic_0.xnor_magic_3.OUT 1.44e-19
C3108 p3_gen_magic_0.xnor_magic_3.OUT a_13553_n6613# 3.87e-19
C3109 a_5515_9163# a_5385_7469# 0.005699f
C3110 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK 1.36099f
C3111 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B Q5 4.93e-19
C3112 a_8643_n5540# VDD 0.38659f
C3113 a_5054_n6024# D2_7 6.69e-21
C3114 7b_counter_0.MDFF_5.tspc2_magic_0.Q D2_6 0.043343f
C3115 a_12387_9730# Q7 0.021558f
C3116 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A D2_3 0.002134f
C3117 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 0.691605f
C3118 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 3.8e-19
C3119 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8825_1669# 0.125951f
C3120 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VDD 1.04322f
C3121 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_4235_3947# 0.671058f
C3122 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A D2_5 0.004746f
C3123 a_17405_3524# D2_3 0.006461f
C3124 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q1 0.265028f
C3125 LD D2_5 0.879417f
C3126 a_12387_1769# D2_4 0.002007f
C3127 p2_gen_magic_0.xnor_magic_1.OUT D2_6 0.004994f
C3128 a_1409_2253# CLK 0.128771f
C3129 a_1559_n1526# D2_7 0.015874f
C3130 7b_counter_0.MDFF_4.tspc2_magic_0.CLK p2_gen_magic_0.xnor_magic_4.OUT 1.22e-19
C3131 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n5540# 0.093592f
C3132 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A CLK 0.321291f
C3133 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 0.003022f
C3134 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_24536_3947# 0.069391f
C3135 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27778_4557# 0.037614f
C3136 7b_counter_0.MDFF_6.tspc2_magic_0.D VDD 1.42971f
C3137 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B p2_gen_magic_0.xnor_magic_0.OUT 0.001021f
C3138 a_1541_n4081# D2_7 0.002646f
C3139 a_20041_9774# Q7 0.032924f
C3140 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.OUT 0.009313f
C3141 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT D2_6 0.082793f
C3142 a_6725_5900# Q6 0.027999f
C3143 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 1.99e-20
C3144 a_1209_7469# a_1409_6275# 0.003083f
C3145 7b_counter_0.MDFF_6.tspc2_magic_0.D D2_1 0.008271f
C3146 7b_counter_0.3_inp_AND_magic_0.A CLK 2.69e-19
C3147 a_20041_4557# Q1 0.001912f
C3148 VDD D2_7 5.78611f
C3149 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 5.15e-19
C3150 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 0.240827f
C3151 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_4651_9163# 0.069391f
C3152 a_2749_7308# a_2749_5900# 0.479729f
C3153 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.09324f
C3154 a_11279_8697# D2_2 0.0364f
C3155 7b_counter_0.3_inp_AND_magic_0.C Q5 0.263526f
C3156 p3_gen_magic_0.xnor_magic_0.OUT Q4 0.009371f
C3157 a_2749_2092# a_1209_1059# 7.54e-20
C3158 a_8825_1669# VDD 0.083906f
C3159 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q1 0.074976f
C3160 D2_7 D2_1 0.660979f
C3161 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_3 2.59e-19
C3162 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_11279_8697# 0.001371f
C3163 7b_counter_0.MDFF_1.tspc2_magic_0.CLK VDD 2.19751f
C3164 7b_counter_0.MDFF_5.tspc2_magic_0.Q D2_2 0.418637f
C3165 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT D2_7 7.57e-19
C3166 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A Q1 0.004261f
C3167 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK 0.004079f
C3168 a_4651_3947# Q6 6.65e-19
C3169 a_12387_8536# Q7 2.93e-19
C3170 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.008398f
C3171 p2_gen_magic_0.xnor_magic_4.OUT VDD 1.48171f
C3172 p2_gen_magic_0.3_inp_AND_magic_0.B a_13553_n2115# 0.175285f
C3173 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B 0.178114f
C3174 7b_counter_0.MDFF_1.tspc2_magic_0.D a_18891_1669# 0.282223f
C3175 p3_gen_magic_0.3_inp_AND_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.005707f
C3176 a_12174_n8579# D2_5 0.007723f
C3177 a_15865_8580# a_15865_7470# 0.003291f
C3178 Q3 D2_5 0.043979f
C3179 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A D2_7 0.087718f
C3180 Q7 Q5 0.946424f
C3181 7b_counter_0.MDFF_1.tspc2_magic_0.Q a_20041_3363# 0.016967f
C3182 LD D2_7 1.081f
C3183 p2_gen_magic_0.xnor_magic_1.OUT D2_2 0.005371f
C3184 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 0.178114f
C3185 7b_counter_0.3_inp_AND_magic_0.C D2_4 0.028537f
C3186 a_20041_8580# D2_3 8.6e-19
C3187 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_15865_6276# 0.279825f
C3188 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VDD 1.24097f
C3189 7b_counter_0.NAND_magic_0.A 7b_counter_0.3_inp_AND_magic_0.A 0.001889f
C3190 a_4235_9163# VDD 1.06848f
C3191 CLK D2_6 0.660277f
C3192 a_14556_n8142# a_16186_n8142# 4.95e-19
C3193 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A Q6 3.37e-19
C3194 a_4235_9163# D2_1 0.002097f
C3195 p2_gen_magic_0.xnor_magic_0.OUT a_8523_n3150# 0.037448f
C3196 Q7 D2_4 0.037182f
C3197 a_27234_1769# a_26126_1124# 0.001529f
C3198 7b_counter_0.3_inp_AND_magic_0.C Q2 0.085313f
C3199 a_15865_9774# a_15865_8580# 0.005574f
C3200 a_1209_3363# Q7 0.009728f
C3201 a_1559_n1042# Q7 0.049258f
C3202 a_11191_10149# D2_6 0.005215f
C3203 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.A 0.001004f
C3204 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n1526# 0.063777f
C3205 a_4235_9163# LD 2.62e-21
C3206 p3_gen_magic_0.xnor_magic_3.OUT a_11708_n6613# 0.057f
C3207 7b_counter_0.MDFF_4.LD p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 5.14e-19
C3208 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_8411_8536# 0.001158f
C3209 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_7.tspc2_magic_0.Q 1.17e-20
C3210 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A a_12931_3363# 0.001034f
C3211 a_20171_6886# Q1 0.002353f
C3212 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_5 1.01933f
C3213 p2_gen_magic_0.3_inp_AND_magic_0.VOUT D2_4 0.002487f
C3214 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.271976f
C3215 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_20041_8580# 1.77e-19
C3216 a_6725_2092# a_8825_1669# 2.9e-20
C3217 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_4496_4877# 0.365826f
C3218 a_11708_n2115# D2_2 0.006396f
C3219 Q2 Q7 1.94553f
C3220 D2_7 Q3 1.15394f
C3221 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A Q6 0.01512f
C3222 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT Q5 4.95e-19
C3223 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_3 0.053092f
C3224 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.xnor_magic_1.OUT 0.040944f
C3225 p3_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.AND2_magic_1.A 0.253673f
C3226 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B Q2 0.049621f
C3227 p2_gen_magic_0.xnor_magic_5.OUT D2_5 1.10379f
C3228 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q3 0.003474f
C3229 a_1209_2253# CLK 0.243862f
C3230 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_9689_1669# 0.004104f
C3231 7b_counter_0.MDFF_4.LD a_16065_1059# 0.003068f
C3232 a_15865_1059# CLK 2.28e-19
C3233 a_23258_1769# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.001158f
C3234 a_11279_8697# CLK 0.015935f
C3235 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_6.tspc2_magic_0.D 0.413248f
C3236 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.003202f
C3237 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VDD 1.33085f
C3238 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN P2 0.315149f
C3239 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT Q5 0.014758f
C3240 a_2749_2092# 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A 2.4e-20
C3241 7b_counter_0.MDFF_1.tspc2_magic_0.CLK Q3 4.27e-19
C3242 a_27234_4513# a_27778_4557# 0.29829f
C3243 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_23672_3947# 0.125951f
C3244 a_9689_6886# VDD 0.003613f
C3245 CLK D2_2 0.540858f
C3246 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A OR_magic_2.A 1.39e-19
C3247 7b_counter_0.MDFF_5.tspc2_magic_0.Q CLK 0.070136f
C3248 7b_counter_0.DFF_magic_0.tg_magic_2.IN CLK 0.014697f
C3249 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK 1.34511f
C3250 p2_gen_magic_0.xnor_magic_4.OUT Q3 0.002591f
C3251 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.005939f
C3252 a_1209_7469# a_1209_6275# 0.005574f
C3253 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A Q4 5.53e-19
C3254 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.P3 6.97e-20
C3255 p3_gen_magic_0.xnor_magic_6.OUT Q5 0.150271f
C3256 a_5054_n1526# p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 6.69e-21
C3257 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT D2_4 0.014268f
C3258 a_17405_2092# Q1 0.010647f
C3259 a_1541_n8095# Q7 0.08832f
C3260 a_11191_10149# a_11279_8697# 0.479729f
C3261 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.3_inp_AND_magic_0.C 0.042297f
C3262 p3_gen_magic_0.xnor_magic_4.OUT a_5054_n6024# 0.418635f
C3263 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n4081# 0.066064f
C3264 p2_gen_magic_0.xnor_magic_1.OUT CLK 0.150366f
C3265 a_20041_9774# D2_3 0.001383f
C3266 a_12174_n4081# Q4 0.001608f
C3267 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A Q3 0.015519f
C3268 a_4496_9609# Q2 0.001226f
C3269 a_16065_4557# VDD 0.063712f
C3270 a_12387_4513# Q1 8.5e-19
C3271 a_8411_9730# D2_2 0.018168f
C3272 p3_gen_magic_0.xnor_magic_3.OUT a_5054_n5540# 0.128084f
C3273 a_21381_4932# Q6 4.02e-19
C3274 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.003171f
C3275 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT CLK 0.245998f
C3276 p2_gen_magic_0.3_inp_AND_magic_0.B a_11708_n2115# 0.002716f
C3277 a_8411_9730# 7b_counter_0.MDFF_5.tspc2_magic_0.Q 0.243646f
C3278 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B p2_gen_magic_0.xnor_magic_3.OUT 1.55e-19
C3279 Q6 Q4 0.265604f
C3280 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VDD 1.07013f
C3281 p3_gen_magic_0.3_inp_AND_magic_0.B D2_6 0.045711f
C3282 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_19152_1223# 0.515297f
C3283 p2_gen_magic_0.xnor_magic_5.OUT D2_7 0.142398f
C3284 7b_counter_0.NAND_magic_0.A 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.314216f
C3285 a_26126_1124# VDD 0.941683f
C3286 a_5185_7469# a_6725_5900# 7.51e-20
C3287 a_4496_10093# VDD 0.76895f
C3288 p2_gen_magic_0.3_inp_AND_magic_0.B CLK 2.37e-19
C3289 7b_counter_0.MDFF_4.LD D2_6 1.15154f
C3290 p3_gen_magic_0.xnor_magic_4.OUT VDD 1.4576f
C3291 a_14756_n3644# D2_5 0.001368f
C3292 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 0.001081f
C3293 7b_counter_0.MDFF_6.tspc2_magic_0.D a_15865_6276# 1.63e-20
C3294 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VDD 1.85748f
C3295 a_13353_n2115# Q5 6.77e-20
C3296 Q5 D2_3 0.62529f
C3297 a_4496_10093# D2_1 0.003209f
C3298 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 0.164969f
C3299 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n8579# 0.093592f
C3300 a_1541_n3150# p2_gen_magic_0.xnor_magic_1.OUT 0.09365f
C3301 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.178114f
C3302 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_5.OUT 1.36e-19
C3303 p3_gen_magic_0.xnor_magic_4.OUT D2_1 0.002623f
C3304 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_20041_9774# 8.53e-19
C3305 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 3.27e-21
C3306 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 9.4e-20
C3307 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT Q4 0.025734f
C3308 a_12931_1059# D2_6 0.003998f
C3309 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B CLK 0.011738f
C3310 7b_counter_0.MDFF_5.LD Q1 0.205628f
C3311 7b_counter_0.DFF_magic_0.tg_magic_0.IN a_27234_4513# 2.63e-20
C3312 7b_counter_0.MDFF_5.tspc2_magic_0.D VDD 1.43217f
C3313 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A Q3 8.78e-21
C3314 7b_counter_0.MDFF_7.tspc2_magic_0.D 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 8.78e-21
C3315 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B a_1209_3363# 0.146237f
C3316 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT D2_4 6.16e-19
C3317 p3_gen_magic_0.xnor_magic_3.OUT a_11492_n6613# 0.001361f
C3318 a_19307_6886# Q1 0.015173f
C3319 D2_3 D2_4 1.58757f
C3320 a_13353_n2115# D2_4 0.003065f
C3321 a_21381_8741# 7b_counter_0.3_inp_AND_magic_0.C 7.58e-20
C3322 a_5054_n6471# p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.001716f
C3323 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_9212_739# 3.22e-21
C3324 a_23793_5904# Q4 0.371901f
C3325 a_11492_n2115# D2_2 0.008915f
C3326 a_1559_n5540# Q7 1.35e-19
C3327 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n3597# 0.063777f
C3328 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B Q5 3.04e-19
C3329 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_23802_1059# 9.27e-19
C3330 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B 0.004701f
C3331 a_5036_n3150# D2_5 0.078851f
C3332 a_15865_7470# Q2 5.69e-19
C3333 p3_gen_magic_0.xnor_magic_5.OUT a_5036_n8095# 0.3716f
C3334 a_17405_8741# a_15865_8580# 0.001529f
C3335 7b_counter_0.MDFF_3.QB Q7 5.73e-19
C3336 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8825_1669# 0.001268f
C3337 a_22062_684# CLK 0.028207f
C3338 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 0.007591f
C3339 7b_counter_0.MDFF_4.LD a_15865_1059# 0.001153f
C3340 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.166749f
C3341 a_6725_684# a_5185_1059# 0.002003f
C3342 a_11191_10149# CLK 0.001996f
C3343 a_20041_3363# Q1 0.013109f
C3344 a_8825_6886# VDD 0.084074f
C3345 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.240827f
C3346 a_21381_3524# a_23672_3947# 1.2e-20
C3347 7b_counter_0.MDFF_4.LD D2_2 0.032737f
C3348 a_21381_8741# Q7 0.052722f
C3349 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B Q5 0.00368f
C3350 7b_counter_0.3_inp_AND_magic_0.C a_23985_7877# 0.610315f
C3351 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 2.05e-19
C3352 Q2 D2_3 0.051234f
C3353 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.002684f
C3354 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_3 0.047009f
C3355 a_8411_9730# CLK 6.58e-19
C3356 7b_counter_0.MDFF_4.tspc2_magic_0.D 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 8.78e-21
C3357 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.011269f
C3358 a_20041_8580# a_19152_6440# 5.39e-19
C3359 a_8523_n7648# Q5 0.323606f
C3360 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.286389f
C3361 7b_counter_0.MDFF_4.tspc2_magic_0.D a_11191_684# 1.08e-19
C3362 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B D2_4 0.02303f
C3363 a_8523_n3597# Q1 0.022022f
C3364 7b_counter_0.NAND_magic_0.A CLK 1.32543f
C3365 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 0.207107f
C3366 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 0.003202f
C3367 a_23560_3728# Q4 0.003438f
C3368 OR_magic_2.A 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 2.3e-20
C3369 a_26126_1124# Q3 0.011812f
C3370 a_15865_9774# Q2 6.82e-19
C3371 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.OUT 0.037144f
C3372 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q6 0.0205f
C3373 a_5515_3947# VDD 0.097495f
C3374 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.340787f
C3375 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN Q3 0.065225f
C3376 a_26126_3480# a_26126_1124# 0.00112f
C3377 7b_counter_0.MDFF_3.QB a_4496_9609# 0.119508f
C3378 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD 1.49164f
C3379 p2_gen_magic_0.3_inp_AND_magic_0.B a_11492_n2115# 7.27e-19
C3380 a_9059_n1973# D2_6 0.001146f
C3381 a_12387_8536# a_12387_6986# 0.003291f
C3382 a_8713_6842# a_9689_6886# 0.240883f
C3383 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_18891_1669# 0.671058f
C3384 a_5036_n3150# D2_7 0.642098f
C3385 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_1 0.009715f
C3386 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.0953f
C3387 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12931_9774# 0.037614f
C3388 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5515_9163# 0.001268f
C3389 a_1409_9773# VDD 0.052909f
C3390 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A Q2 7.6e-19
C3391 a_11492_n2115# a_11708_n2115# 0.329078f
C3392 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 1.1e-20
C3393 a_23672_3947# a_24536_3947# 0.009722f
C3394 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_1 0.01666f
C3395 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12387_9730# 0.149276f
C3396 a_5515_3947# LD 8.49e-19
C3397 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8939_n3150# 5.84e-19
C3398 7b_counter_0.MDFF_0.tspc2_magic_0.D 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.423451f
C3399 a_1409_9773# D2_1 0.017468f
C3400 p2_gen_magic_0.xnor_magic_4.OUT a_5036_n3150# 0.034857f
C3401 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26126_1124# 0.431521f
C3402 p3_gen_magic_0.P3 CLK 0.233508f
C3403 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n8579# 0.066064f
C3404 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_19841_4557# 0.279825f
C3405 a_1209_8579# a_1409_8579# 0.299584f
C3406 7b_counter_0.MDFF_5.tspc2_magic_0.CLK D2_6 0.502796f
C3407 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A Q2 8.35e-19
C3408 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_3.tspc2_magic_0.Q 4.47e-20
C3409 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1409_3363# 0.001034f
C3410 a_12387_575# D2_6 3.06e-19
C3411 a_1409_7469# CLK 0.13379f
C3412 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1409_9773# 0.036959f
C3413 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_26038_4932# 0.414018f
C3414 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A Q7 0.031311f
C3415 DFF_magic_0.tg_magic_1.IN CLK 0.699469f
C3416 7b_counter_0.MDFF_7.tspc2_magic_0.D a_27234_4513# 1.63e-20
C3417 a_1409_9773# LD 0.003696f
C3418 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n6024# 0.063777f
C3419 p2_gen_magic_0.xnor_magic_6.OUT a_8523_n4081# 0.465726f
C3420 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_4.OUT 6.89e-21
C3421 7b_counter_0.MDFF_4.LD CLK 1.54694f
C3422 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_4496_4393# 0.515297f
C3423 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2e-19
C3424 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_9212_739# 0.671058f
C3425 a_11279_1124# a_9212_739# 0.002118f
C3426 a_5036_n8579# D2_7 0.037922f
C3427 a_9059_n1973# D2_2 0.005701f
C3428 a_21504_5904# Q4 0.002361f
C3429 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_0.IN 0.859117f
C3430 a_12387_6986# Q2 0.100292f
C3431 p3_gen_magic_0.xnor_magic_6.OUT a_12174_n7648# 0.143702f
C3432 a_5036_n7648# a_5036_n8095# 0.014233f
C3433 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 1.09743f
C3434 p2_gen_magic_0.xnor_magic_3.OUT D2_6 0.043388f
C3435 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A Q4 0.001013f
C3436 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.025064f
C3437 a_6725_5900# VDD 1.55921f
C3438 a_8955_8580# D2_2 0.134289f
C3439 7b_counter_0.MDFF_0.tspc2_magic_0.Q p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 2.24e-19
C3440 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12387_8536# 0.001985f
C3441 7b_counter_0.3_inp_AND_magic_0.A a_24401_7877# 0.02473f
C3442 a_7303_3480# Q5 0.007564f
C3443 a_5470_n1973# D2_3 0.005701f
C3444 p2_gen_magic_0.xnor_magic_3.OUT a_13553_n2115# 3.87e-19
C3445 a_17405_2092# 7b_counter_0.MDFF_1.tspc2_magic_0.D 0.134004f
C3446 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8955_8580# 0.016967f
C3447 a_15865_2253# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.001158f
C3448 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_17405_10149# 3.58e-20
C3449 a_11279_8697# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 0.132169f
C3450 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.tspc2_magic_0.Q 0.003482f
C3451 a_5515_9163# D2_7 4.45e-19
C3452 a_4235_3947# 7b_counter_0.MDFF_0.tspc2_magic_0.Q 1.94e-20
C3453 a_15865_3363# a_15865_2253# 0.003291f
C3454 7b_counter_0.MDFF_5.tspc2_magic_0.D a_8713_6842# 0.036809f
C3455 7b_counter_0.MDFF_5.tspc2_magic_0.CLK D2_2 0.055244f
C3456 7b_counter_0.NAND_magic_0.A 7b_counter_0.MDFF_4.LD 1.05485f
C3457 a_9212_5956# Q2 0.098084f
C3458 a_12387_575# D2_2 0.003327f
C3459 7b_counter_0.MDFF_5.tspc2_magic_0.Q 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 0.004808f
C3460 a_9212_739# VDD 0.975666f
C3461 7b_counter_0.MDFF_3.tspc2_magic_0.D VDD 1.42628f
C3462 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT Q6 0.633261f
C3463 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1209_8579# 0.001985f
C3464 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A Q7 3.39e-19
C3465 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_1.IN 0.013133f
C3466 a_4651_3947# VDD 0.05128f
C3467 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q1 0.012436f
C3468 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n8095# 0.083665f
C3469 a_8713_1625# Q5 0.007615f
C3470 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_5 0.056714f
C3471 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.166649f
C3472 7b_counter_0.MDFF_3.tspc2_magic_0.D D2_1 0.005922f
C3473 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q4 1.64e-19
C3474 a_8643_n1973# D2_6 0.012509f
C3475 a_8713_6842# a_8825_6886# 0.043767f
C3476 a_11279_6341# a_9689_6886# 2.34e-20
C3477 7b_counter_0.MDFF_6.tspc2_magic_0.Q Q7 0.185257f
C3478 a_1957_n3150# D2_7 6.21e-19
C3479 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A Q6 3.37e-19
C3480 a_12387_9730# a_12931_9774# 0.29829f
C3481 p2_gen_magic_0.xnor_magic_3.OUT D2_2 0.190073f
C3482 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8643_n5540# 1.05e-19
C3483 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 2.34e-19
C3484 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_3.tspc2_magic_0.D 8.78e-21
C3485 a_5054_n1973# p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 5.81e-19
C3486 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_4651_9163# 0.004104f
C3487 a_4235_9163# a_5515_9163# 0.007202f
C3488 7b_counter_0.MDFF_3.tspc2_magic_0.D LD 8.18e-19
C3489 a_11191_684# p2_gen_magic_0.xnor_magic_4.OUT 1.2e-19
C3490 a_7215_10149# VDD 1.55668f
C3491 a_21381_3524# Q1 0.111781f
C3492 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_2.IN 6.95e-19
C3493 a_8713_1625# D2_4 7.9e-19
C3494 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VDD 1.23949f
C3495 a_14556_n3644# D2_5 7.76e-19
C3496 p3_gen_magic_0.3_inp_AND_magic_0.A p3_gen_magic_0.3_inp_AND_magic_0.C 0.042297f
C3497 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A Q2 7.6e-19
C3498 a_2749_3524# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.018983f
C3499 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.251813f
C3500 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A a_17405_5901# 0.414018f
C3501 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q5 8.31e-19
C3502 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A D2_1 3.01e-19
C3503 a_8955_4557# D2_6 0.00606f
C3504 a_1209_7469# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 0.146237f
C3505 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_21381_8741# 0.036613f
C3506 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_6.OUT 0.017325f
C3507 a_11191_5901# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 1.51e-21
C3508 a_1209_7469# CLK 0.260912f
C3509 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VDD 1.09061f
C3510 a_5185_2253# Q7 0.011994f
C3511 7b_counter_0.MDFF_4.LD DFF_magic_0.tg_magic_1.IN 8.87e-20
C3512 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT Q1 2.49e-19
C3513 p3_gen_magic_0.xnor_magic_1.OUT D2_6 2.33527f
C3514 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_7 0.001733f
C3515 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A LD 5.51e-19
C3516 a_8955_8580# CLK 0.009907f
C3517 a_1409_1059# D2_5 0.001213f
C3518 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VDD 1.29805f
C3519 divide_by_2_1.tg_magic_3.IN divide_by_2_1.tg_magic_1.IN 1.17013f
C3520 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_4 2.79e-19
C3521 a_1559_n6471# p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 7.35e-19
C3522 a_8643_n1973# D2_2 0.054184f
C3523 a_1541_n8579# D2_7 0.062784f
C3524 a_5470_n6471# D2_3 0.005701f
C3525 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A CLK 0.002249f
C3526 p2_gen_magic_0.xnor_magic_0.OUT a_13353_n2115# 1.73e-20
C3527 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.3_inp_AND_magic_0.B 0.010333f
C3528 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n1042# 0.067344f
C3529 a_11292_n2115# p2_gen_magic_0.3_inp_AND_magic_0.A 0.12467f
C3530 p2_gen_magic_0.xnor_magic_0.OUT D2_3 1.56e-19
C3531 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A D2_1 5.31e-20
C3532 p3_gen_magic_0.xnor_magic_6.OUT a_8939_n7648# 0.06406f
C3533 7b_counter_0.MDFF_5.tspc2_magic_0.CLK CLK 0.037826f
C3534 Q4 P2 0.314629f
C3535 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A a_12931_8580# 1.77e-19
C3536 a_12931_9774# a_12387_8536# 0.003083f
C3537 a_12931_7470# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 5.46e-20
C3538 7b_counter_0.MDFF_4.LD a_12931_1059# 0.003068f
C3539 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.178114f
C3540 a_5452_n3150# Q6 7.91e-19
C3541 7b_counter_0.MDFF_4.tspc2_magic_0.CLK Q4 0.001622f
C3542 a_8523_n4081# p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 1.05e-19
C3543 7b_counter_0.3_inp_AND_magic_0.A a_24185_7877# 0.075783f
C3544 a_19841_3363# D2_3 0.243646f
C3545 a_16065_2253# 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.001034f
C3546 a_5054_n1973# D2_3 0.054067f
C3547 p2_gen_magic_0.xnor_magic_3.OUT a_11708_n2115# 0.057f
C3548 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 0.002402f
C3549 a_21381_3524# 7b_counter_0.MDFF_7.tspc2_magic_0.Q 6.46e-19
C3550 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_26038_4932# 0.00215f
C3551 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A LD 0.445505f
C3552 a_4651_9163# D2_7 0.0074f
C3553 p3_gen_magic_0.xnor_magic_3.OUT D2_6 5.14e-19
C3554 a_19307_1669# a_19152_739# 0.001643f
C3555 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C3556 a_11279_6341# 7b_counter_0.MDFF_5.tspc2_magic_0.D 0.134004f
C3557 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 0.16497f
C3558 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VDD 1.30001f
C3559 a_2749_8740# VDD 0.954212f
C3560 a_1209_9773# a_1209_8579# 0.005574f
C3561 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n3597# 0.083665f
C3562 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_27234_575# 1.63e-20
C3563 a_21381_4932# VDD 1.56584f
C3564 a_5385_6275# Q6 1.77e-19
C3565 a_2749_8740# D2_1 0.002184f
C3566 a_1409_1059# D2_7 0.019488f
C3567 VDD Q4 13.062201f
C3568 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.43627f
C3569 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.OUT 0.175616f
C3570 7b_counter_0.MDFF_0.tspc2_magic_0.Q p2_gen_magic_0.xnor_magic_3.OUT 1.47e-19
C3571 p3_gen_magic_0.3_inp_AND_magic_0.C D2_5 0.006821f
C3572 D2_1 Q4 0.135174f
C3573 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_2749_8740# 2.4e-20
C3574 a_4235_9163# a_4651_9163# 0.16113f
C3575 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 9.4e-20
C3576 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B Q6 0.01038f
C3577 a_27234_1769# 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 0.001158f
C3578 a_12174_n3597# D2_5 0.251387f
C3579 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A a_1209_4557# 1.28e-19
C3580 7b_counter_0.MDFF_6.tspc2_magic_0.D a_20171_6886# 2.1e-20
C3581 7b_counter_0.MDFF_4.tspc2_magic_0.CLK p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 8.78e-19
C3582 a_2749_4932# 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 0.00215f
C3583 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n3150# 0.011524f
C3584 a_5054_n1042# Q5 0.008791f
C3585 a_26038_4932# a_27234_3319# 7.51e-20
C3586 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_24536_3947# 0.004104f
C3587 LD Q4 1.92846f
C3588 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 4e-20
C3589 a_1209_7469# a_1409_7469# 0.299584f
C3590 p3_gen_magic_0.xnor_magic_3.OUT D2_2 0.078371f
C3591 7b_counter_0.MDFF_6.tspc2_magic_0.Q D2_3 0.011531f
C3592 a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 0.149276f
C3593 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.148797f
C3594 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A D2_6 0.002219f
C3595 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VDD 3.58078f
C3596 a_8955_3363# a_8713_1625# 5.39e-19
C3597 a_5185_1059# p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 4.61e-20
C3598 p3_gen_magic_0.xnor_magic_5.OUT D2_5 0.001041f
C3599 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_3.OUT 0.020085f
C3600 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q5 7.94e-22
C3601 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_3480# 1e-20
C3602 a_1209_1059# D2_5 0.001663f
C3603 a_23258_1769# CLK 0.056546f
C3604 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_20041_4557# 0.037614f
C3605 a_5054_n1042# D2_4 1.31e-19
C3606 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK D2_1 0.161265f
C3607 a_1975_n1973# Q7 0.005876f
C3608 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT Q5 0.01303f
C3609 a_12931_9774# a_12931_8580# 0.020635f
C3610 a_5054_n6471# D2_3 0.054067f
C3611 7b_counter_0.MDFF_1.tspc2_magic_0.Q Q1 0.086083f
C3612 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 0.00221f
C3613 a_8523_n7648# a_8939_n7648# 0.002223f
C3614 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 8.78e-21
C3615 p2_gen_magic_0.xnor_magic_6.OUT VDD 1.30086f
C3616 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.LD 3.09e-20
C3617 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD 1.02706f
C3618 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B CLK 0.002402f
C3619 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.150184f
C3620 a_27778_2253# CLK 0.205288f
C3621 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 0.005939f
C3622 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_9212_739# 1.94e-20
C3623 a_1409_4557# CLK 7.14e-19
C3624 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.31462f
C3625 7b_counter_0.MDFF_4.LD a_12387_575# 3.96e-19
C3626 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11279_1124# 0.431521f
C3627 a_23258_1769# a_22062_684# 7.51e-20
C3628 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 4.5e-19
C3629 a_21381_4932# Q3 0.0012f
C3630 p2_gen_magic_0.xnor_magic_6.OUT D2_1 6.06e-19
C3631 p2_gen_magic_0.AND2_magic_1.A D2_2 0.00215f
C3632 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B D2_7 0.009349f
C3633 7b_counter_0.3_inp_AND_magic_0.A a_23207_5885# 2.57e-19
C3634 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_26126_3480# 2.4e-20
C3635 7b_counter_0.MDFF_6.tspc2_magic_0.Q 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 0.002402f
C3636 p2_gen_magic_0.xnor_magic_3.OUT a_11492_n2115# 0.001361f
C3637 a_12174_n8579# Q4 0.036643f
C3638 Q3 Q4 0.491372f
C3639 Q7 Q6 6.56387f
C3640 a_5054_n1042# Q2 0.00341f
C3641 p3_gen_magic_0.xnor_magic_0.OUT D2_3 0.006968f
C3642 a_9212_5956# 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 5.62e-20
C3643 a_12387_575# a_12931_1059# 0.29829f
C3644 a_12387_3319# a_12387_1769# 0.003291f
C3645 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_17405_2092# 0.018983f
C3646 a_4496_4877# a_4235_3947# 0.655098f
C3647 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.OUT 7.54e-20
C3648 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.AND2_magic_1.A 0.010924f
C3649 a_27234_4513# VDD 0.930575f
C3650 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VDD 1.03533f
C3651 a_16386_n3644# Q4 0.011403f
C3652 a_2749_10148# VDD 1.55786f
C3653 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VDD 1.3102f
C3654 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.032187f
C3655 a_5185_6275# Q6 5.54e-19
C3656 7b_counter_0.MDFF_5.tspc2_magic_0.D a_12387_5792# 1.63e-20
C3657 p3_gen_magic_0.xnor_magic_5.OUT D2_7 0.314599f
C3658 a_1209_1059# D2_7 0.016083f
C3659 a_16186_n3644# p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 3.96e-20
C3660 a_2749_10148# D2_1 0.003237f
C3661 a_17405_684# p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.78e-19
C3662 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B VDD 1.19332f
C3663 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.00112f
C3664 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VDD 1.28211f
C3665 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_4235_9163# 7.16e-19
C3666 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.033071f
C3667 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 0.008877f
C3668 7b_counter_0.3_inp_AND_magic_0.C a_23793_5904# 0.054305f
C3669 a_14756_n8142# D2_5 0.003236f
C3670 a_6725_7308# a_8825_6886# 3.09e-20
C3671 a_5185_1059# Q5 0.014407f
C3672 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_7 9.27e-19
C3673 a_4496_9609# Q6 3.63e-19
C3674 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.002381f
C3675 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.973393f
C3676 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A a_17405_5901# 3.58e-20
C3677 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_2749_10148# 3.58e-20
C3678 a_4496_10093# a_4651_9163# 0.001643f
C3679 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_7303_3480# 2.4e-20
C3680 a_1209_8579# Q2 0.003166f
C3681 a_19152_1223# Q4 2.83e-19
C3682 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.AND2_magic_1.A 0.007533f
C3683 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A Q7 0.001074f
C3684 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_2.IN 0.973398f
C3685 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT Q4 0.04535f
C3686 a_8523_n3597# D2_5 0.003217f
C3687 7b_counter_0.DFF_magic_0.tg_magic_3.OUT CLK 0.455905f
C3688 7b_counter_0.MDFF_6.tspc2_magic_0.D a_19307_6886# 0.004574f
C3689 a_23793_5904# Q7 2.05e-20
C3690 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A D2_5 0.012503f
C3691 p2_gen_magic_0.xnor_magic_5.OUT Q4 0.07414f
C3692 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23672_3947# 0.001268f
C3693 p3_gen_magic_0.xnor_magic_0.OUT a_8523_n7648# 0.037448f
C3694 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q3 4.44e-19
C3695 a_5185_1059# D2_4 6.03e-19
C3696 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT Q6 0.007688f
C3697 divide_by_2_1.tg_magic_0.IN divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 0.272186f
C3698 a_11191_5901# Q2 0.046952f
C3699 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_2.IN 0.011009f
C3700 DFF_magic_0.D DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.025829f
C3701 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11191_4932# 4.22e-19
C3702 a_5036_n7648# D2_5 0.003766f
C3703 a_15865_7470# 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 0.146237f
C3704 7b_counter_0.MDFF_4.LD a_23258_1769# 0.224142f
C3705 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.16497f
C3706 a_5054_n6024# p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 6.69e-21
C3707 a_1559_n1973# Q7 0.042034f
C3708 a_1559_n6024# p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 7.02e-19
C3709 a_27234_575# DFF_magic_0.tg_magic_3.OUT 0.002608f
C3710 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.08809f
C3711 7b_counter_0.MDFF_4.LD a_8955_4557# 1.1e-19
C3712 7b_counter_0.NAND_magic_0.A 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.004549f
C3713 a_19841_4557# a_21381_4932# 0.002003f
C3714 a_8523_n3150# VDD 0.001396f
C3715 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8955_8580# 0.007492f
C3716 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_7303_8697# 0.001004f
C3717 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.237983f
C3718 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.xnor_magic_1.OUT 0.046715f
C3719 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B D2_3 0.026146f
C3720 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n3150# 0.107246f
C3721 a_20171_1669# CLK 0.002179f
C3722 a_12387_1769# 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 0.001985f
C3723 7b_counter_0.MDFF_4.LD a_27778_2253# 0.037786f
C3724 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT D2_1 0.017156f
C3725 7b_counter_0.MDFF_1.tspc2_magic_0.CLK a_20041_3363# 0.007492f
C3726 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A D2_3 0.102282f
C3727 a_16065_3363# Q1 0.010754f
C3728 a_8523_n8095# Q1 1.86e-20
C3729 p2_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 1.07e-19
C3730 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1957_n7648# 0.005701f
C3731 7b_counter_0.3_inp_AND_magic_0.A a_22991_5885# 8.94e-20
C3732 a_5054_n5540# D2_4 0.021634f
C3733 a_27234_4513# a_26126_3480# 7.54e-20
C3734 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_17405_8741# 0.001371f
C3735 a_15865_3363# D2_3 4e-19
C3736 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT 0.164969f
C3737 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B Q3 2.69e-19
C3738 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_4496_4393# 0.011612f
C3739 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A D2_7 0.104162f
C3740 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A Q3 0.369964f
C3741 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VDD 1.02775f
C3742 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B Q6 0.013699f
C3743 7b_counter_0.DFF_magic_0.tg_magic_2.OUT CLK 0.381933f
C3744 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VDD 1.49154f
C3745 7b_counter_0.MDFF_3.tspc2_magic_0.D a_5515_9163# 2.1e-20
C3746 p2_gen_magic_0.xnor_magic_1.OUT a_1541_n3597# 0.371458f
C3747 p2_gen_magic_0.xnor_magic_5.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.980376f
C3748 a_14756_n3644# Q4 0.003174f
C3749 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT D2_1 7.76e-19
C3750 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q1 0.099518f
C3751 mux_magic_0.IN2 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT 4.95e-19
C3752 a_9412_5956# VDD 0.725398f
C3753 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B VDD 1.19386f
C3754 a_5036_n7648# D2_7 0.057775f
C3755 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A D2_4 0.101065f
C3756 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_16065_1059# 9.27e-19
C3757 Q6 D2_3 0.098813f
C3758 a_11292_n6613# p3_gen_magic_0.3_inp_AND_magic_0.A 0.12467f
C3759 a_5054_n5540# Q2 0.004397f
C3760 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5054_n5540# 0.064941f
C3761 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 0.010333f
C3762 p3_gen_magic_0.xnor_magic_0.OUT a_13353_n6613# 1.73e-20
C3763 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_1.IN 0.340787f
C3764 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19152_6440# 0.012716f
C3765 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 1.55e-19
C3766 a_15865_2253# VDD 0.821356f
C3767 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_4496_10093# 1.29e-19
C3768 a_23258_575# VDD 0.938137f
C3769 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A Q6 0.006686f
C3770 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VDD 1.24107f
C3771 a_12387_575# p2_gen_magic_0.xnor_magic_3.OUT 2.98e-20
C3772 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11279_3480# 0.431521f
C3773 a_6725_7308# a_6725_5900# 0.479729f
C3774 a_15865_9774# Q6 3.01e-19
C3775 divide_by_2_0.tg_magic_0.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 0.272186f
C3776 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A D2_1 0.014463f
C3777 a_8643_n1973# a_9059_n1973# 5.82e-19
C3778 a_18891_1669# Q4 7.16e-21
C3779 DFF_magic_0.D CLK 0.956771f
C3780 a_2749_7308# 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 2.4e-20
C3781 a_5185_7469# Q7 0.03539f
C3782 a_12590_n7648# a_12174_n8095# 0.013021f
C3783 a_5036_n3597# D2_5 0.050398f
C3784 a_27234_1769# a_26038_684# 7.51e-20
C3785 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 1.64e-20
C3786 7b_counter_0.3_inp_AND_magic_0.B Q4 0.001569f
C3787 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_3 0.018494f
C3788 7b_counter_0.MDFF_6.tspc2_magic_0.D a_17405_5901# 1.08e-19
C3789 7b_counter_0.NAND_magic_0.A 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.341127f
C3790 a_21504_5904# Q7 0.48071f
C3791 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_3524# 1.01e-20
C3792 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT D2_7 0.046858f
C3793 p2_gen_magic_0.xnor_magic_4.OUT a_11292_n2115# 0.318049f
C3794 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B D2_5 0.002674f
C3795 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 0.001081f
C3796 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A CLK 6.07e-20
C3797 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.xnor_magic_5.OUT 1.38e-19
C3798 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A LD 5.51e-19
C3799 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B a_7215_10149# 0.189314f
C3800 7b_counter_0.DFF_magic_0.tg_magic_0.IN 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 4.89e-20
C3801 p2_gen_magic_0.AND2_magic_1.A p3_gen_magic_0.3_inp_AND_magic_0.B 2.51e-20
C3802 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B Q1 7.94e-19
C3803 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 0.178114f
C3804 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A Q6 0.027337f
C3805 a_1559_n6471# Q7 9.27e-19
C3806 a_5185_7469# a_5185_6275# 0.005574f
C3807 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_20041_3363# 5.46e-20
C3808 p2_gen_magic_0.xnor_magic_6.OUT a_14756_n3644# 0.128771f
C3809 a_15865_7470# a_16065_7470# 0.299584f
C3810 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A D2_6 5.9e-19
C3811 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4235_3947# 0.282223f
C3812 a_4496_9609# a_5185_7469# 3.03e-19
C3813 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A Q6 3.87e-19
C3814 7b_counter_0.NAND_magic_0.A DFF_magic_0.D 0.874177f
C3815 a_15865_4557# CLK 3.56e-19
C3816 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_12931_2253# 1.77e-19
C3817 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 0.00112f
C3818 a_5452_n3150# VDD 0.005602f
C3819 7b_counter_0.MDFF_4.LD a_20171_1669# 8.49e-19
C3820 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_12387_1769# 5.28e-20
C3821 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_5385_7469# 0.007492f
C3822 a_19307_1669# CLK 0.002015f
C3823 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT OR_magic_2.A 0.006363f
C3824 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A D2_6 1.41e-19
C3825 a_12387_1769# a_11279_1124# 0.001529f
C3826 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B Q3 2.23e-19
C3827 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_15865_8580# 0.001158f
C3828 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 1.1e-20
C3829 a_12931_3363# Q1 0.011133f
C3830 7b_counter_0.MDFF_0.tspc2_magic_0.CLK D2_4 5.78e-19
C3831 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT Q7 0.026414f
C3832 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q5 2.92e-19
C3833 a_5036_n3597# D2_7 0.250622f
C3834 a_12174_n3150# D2_2 3.26e-19
C3835 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n1526# 0.082959f
C3836 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_1209_3363# 5.28e-20
C3837 a_4235_3947# a_4496_4393# 0.301553f
C3838 a_23258_575# Q3 3.14e-19
C3839 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q1 0.003076f
C3840 a_11292_n6613# D2_5 0.047626f
C3841 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_5 0.053654f
C3842 a_17405_684# a_15865_1059# 0.002003f
C3843 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_2.IN 0.973393f
C3844 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A CLK 2.5e-20
C3845 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.001125f
C3846 a_24059_4877# Q4 3.69e-19
C3847 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4651_9163# 0.004574f
C3848 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT D2_6 0.043402f
C3849 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q5 3.73e-19
C3850 a_1541_n3150# a_1541_n3597# 0.014233f
C3851 p2_gen_magic_0.xnor_magic_4.OUT a_5036_n3597# 0.009286f
C3852 a_16186_n3644# Q4 0.05629f
C3853 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A Q4 5.53e-19
C3854 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_6 2.34e-19
C3855 a_5385_6275# VDD 0.119528f
C3856 a_16065_2253# VDD 0.017748f
C3857 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_8411_3319# 0.146237f
C3858 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B D2_4 0.012496f
C3859 a_19152_739# D2_4 0.01311f
C3860 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A Q1 1.35e-19
C3861 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_15865_1059# 0.149276f
C3862 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN 0.010724f
C3863 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5385_1059# 0.037614f
C3864 OR_magic_2.A DFF_magic_0.tg_magic_2.OUT 0.342811f
C3865 a_12387_1769# VDD 0.808402f
C3866 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.025046f
C3867 a_26038_684# VDD 1.55668f
C3868 a_14556_n8142# D2_5 0.001802f
C3869 a_8955_9774# VDD 0.093707f
C3870 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 1.36e-20
C3871 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_11191_4932# 0.189314f
C3872 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK 1.32578f
C3873 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A Q4 0.001089f
C3874 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B VDD 1.20341f
C3875 DFF_magic_0.D DFF_magic_0.tg_magic_1.IN 0.067419f
C3876 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT D2_4 0.003446f
C3877 a_5054_n1526# p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 7.12e-21
C3878 7b_counter_0.MDFF_5.LD a_8825_6886# 8.49e-19
C3879 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A D2_2 0.037193f
C3880 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5054_n1042# 7.23e-20
C3881 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_11279_8697# 2.4e-20
C3882 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_12387_3319# 0.146237f
C3883 a_1409_8579# CLK 0.009697f
C3884 DFF_magic_0.D 7b_counter_0.MDFF_4.LD 1.04659f
C3885 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n4081# 0.093592f
C3886 a_5385_6275# LD 1.1e-19
C3887 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q2 2.56e-19
C3888 a_8939_n3150# D2_6 0.005701f
C3889 a_12590_n3150# D2_5 0.006365f
C3890 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A D2_2 5.7e-19
C3891 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT D2_4 1.42e-19
C3892 mux_magic_0.IN2 divide_by_2_0.tg_magic_2.IN 0.314216f
C3893 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8939_n7648# 1.05e-19
C3894 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B a_2749_4932# 4.23e-19
C3895 a_8713_6842# a_9412_5956# 0.013434f
C3896 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_7 0.003757f
C3897 a_11279_6341# 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 2.4e-20
C3898 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.032187f
C3899 a_5385_2253# D2_5 0.131565f
C3900 p3_gen_magic_0.xnor_magic_4.OUT a_5036_n7648# 0.035422f
C3901 a_2749_684# Q7 0.009821f
C3902 divide_by_2_1.tg_magic_1.IN a_34156_n889# 5.83e-20
C3903 a_27234_575# a_27778_1059# 0.29829f
C3904 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_26126_1124# 0.132169f
C3905 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.08311f
C3906 a_8411_8536# D2_2 0.31821f
C3907 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_2 0.0177f
C3908 a_7303_3480# Q6 0.152096f
C3909 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12931_6276# 0.037614f
C3910 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8411_8536# 0.029386f
C3911 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A Q6 3.37e-19
C3912 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q2 0.009637f
C3913 a_5185_7469# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 0.001158f
C3914 a_5452_n7648# Q6 0.001582f
C3915 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4496_4877# 0.120019f
C3916 a_1559_n1526# Q7 0.052991f
C3917 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT Q5 3.72e-19
C3918 7b_counter_0.3_inp_AND_magic_0.C VDD 1.44601f
C3919 a_2749_3524# a_4235_3947# 0.002118f
C3920 a_8411_3319# Q7 0.004064f
C3921 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A D2_3 3.7e-19
C3922 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_16065_8580# 0.001034f
C3923 a_1541_n4081# Q7 0.002629f
C3924 7b_counter_0.MDFF_4.LD a_15865_4557# 0.002086f
C3925 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.001313f
C3926 p2_gen_magic_0.3_inp_AND_magic_0.C Q4 0.308838f
C3927 a_19152_6440# Q6 4.92e-19
C3928 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_2749_7308# 0.132169f
C3929 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.161613f
C3930 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT DFF_magic_0.tg_magic_3.OUT 0.175652f
C3931 a_16065_1059# Q5 8.32e-19
C3932 VDD Q7 8.66883f
C3933 a_5054_n1526# D2_3 0.236724f
C3934 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_17405_7309# 0.431521f
C3935 a_4496_4877# a_4496_4393# 0.014143f
C3936 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_17405_10149# 0.189314f
C3937 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_3.tspc2_magic_0.D 0.001711f
C3938 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B VDD 1.20935f
C3939 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT D2_4 1.13e-19
C3940 a_26038_684# Q3 0.01134f
C3941 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B CLK 0.003332f
C3942 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A CLK 0.006101f
C3943 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A CLK 3.05e-19
C3944 7b_counter_0.3_inp_AND_magic_0.C LD 0.054829f
C3945 D2_1 Q7 0.342614f
C3946 a_5054_n6471# p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 5.81e-19
C3947 a_17405_3524# CLK 0.043594f
C3948 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A 1.1e-20
C3949 7b_counter_0.3_inp_AND_magic_0.A Q5 0.270371f
C3950 a_2749_8740# a_4651_9163# 2.34e-20
C3951 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B a_21381_4932# 0.189314f
C3952 p2_gen_magic_0.xnor_magic_5.OUT a_5452_n3150# 0.06406f
C3953 a_22150_1124# Q4 0.136867f
C3954 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_21381_3524# 2.4e-20
C3955 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.AND2_magic_1.A 2.36e-19
C3956 a_14556_n3644# Q4 0.018348f
C3957 p2_gen_magic_0.3_inp_AND_magic_0.VOUT VDD 1.79605f
C3958 a_5185_6275# VDD 0.973561f
C3959 a_8643_n6471# Q5 3.78e-19
C3960 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A CLK 0.001885f
C3961 a_12931_2253# VDD 0.012214f
C3962 a_16065_1059# D2_4 0.004104f
C3963 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q4 0.005634f
C3964 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A DFF_magic_0.tg_magic_3.OUT 0.0013f
C3965 divide_by_2_0.tg_magic_3.OUT divide_by_2_0.tg_magic_3.IN 0.787551f
C3966 LD Q7 0.165025f
C3967 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A CLK 0.01832f
C3968 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_5185_1059# 0.279825f
C3969 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.237983f
C3970 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A a_16065_9774# 9.27e-19
C3971 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A D2_5 1.18e-19
C3972 p3_gen_magic_0.AND2_magic_1.A D2_6 0.093454f
C3973 a_12174_n8095# D2_5 0.248327f
C3974 a_4496_9609# VDD 1.07633f
C3975 a_12931_4557# D2_2 0.0012f
C3976 divide_by_2_1.tg_magic_3.OUT divide_by_2_1.tg_magic_0.IN 0.859117f
C3977 7b_counter_0.3_inp_AND_magic_0.A D2_4 0.012978f
C3978 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_18891_1669# 7.16e-19
C3979 7b_counter_0.MDFF_1.tspc2_magic_0.D Q1 0.006076f
C3980 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A D2_5 0.002134f
C3981 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK 1.83e-19
C3982 a_4496_9609# D2_1 0.001309f
C3983 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_11191_10149# 3.58e-20
C3984 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11191_684# 0.189314f
C3985 a_12387_9730# a_11279_8697# 7.54e-20
C3986 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.xnor_magic_6.OUT 0.026656f
C3987 a_1409_1059# Q4 0.129597f
C3988 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B a_26038_684# 0.189314f
C3989 a_8411_8536# CLK 0.019179f
C3990 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A a_6725_684# 0.414018f
C3991 a_5185_6275# LD 3.96e-19
C3992 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VDD 1.18728f
C3993 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A Q2 8.26e-19
C3994 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.OUT 0.241029f
C3995 7b_counter_0.3_inp_AND_magic_0.C Q3 0.285079f
C3996 7b_counter_0.NAND_magic_0.A 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B 2.36e-20
C3997 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_1.IN 4.63e-20
C3998 Q5 D2_6 1.56929f
C3999 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B a_18891_6886# 7.16e-19
C4000 a_24185_7877# a_24401_7877# 0.329078f
C4001 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD 1.07554f
C4002 a_11279_6341# a_9412_5956# 1.39e-20
C4003 a_2749_2092# D2_5 0.056226f
C4004 OR_magic_1.VOUT divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT 1.34511f
C4005 a_4496_9609# LD 0.007507f
C4006 7b_counter_0.3_inp_AND_magic_0.A Q2 0.001013f
C4007 a_6725_2092# Q7 0.004318f
C4008 a_1559_n6024# Q7 5.03e-21
C4009 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT D2_1 4.97e-19
C4010 a_11492_n6613# p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 5.63e-20
C4011 p3_gen_magic_0.xnor_magic_0.OUT a_11708_n6613# 0.02473f
C4012 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12387_5792# 0.279825f
C4013 a_19152_5956# D2_3 0.06582f
C4014 a_8411_9730# a_8411_8536# 0.005574f
C4015 Q3 Q7 0.92204f
C4016 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT P2 0.337059f
C4017 p3_gen_magic_0.xnor_magic_6.OUT VDD 1.34151f
C4018 p2_gen_magic_0.xnor_magic_6.OUT a_14556_n3644# 0.249081f
C4019 a_12387_6986# a_12931_7470# 0.2945f
C4020 a_5185_2253# a_5185_1059# 0.005574f
C4021 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1559_n5540# 1.66e-20
C4022 a_15865_8580# CLK 0.268792f
C4023 a_24003_10051# 7b_counter_0.3_inp_AND_magic_0.A 2.32e-20
C4024 D2_6 D2_4 1.08902f
C4025 a_8643_n1042# Q1 0.001111f
C4026 a_2749_3524# a_4496_4877# 1.39e-20
C4027 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A D2_7 0.110179f
C4028 7b_counter_0.MDFF_4.tspc2_magic_0.CLK D2_3 6.8e-19
C4029 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 0.0035f
C4030 a_5054_n6024# D2_3 0.238989f
C4031 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n8579# 0.066064f
C4032 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27778_3363# 0.001034f
C4033 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n8579# 0.093592f
C4034 a_19841_9774# a_19841_8580# 0.005574f
C4035 a_18891_6886# Q6 3.53e-20
C4036 p2_gen_magic_0.3_inp_AND_magic_0.VOUT Q3 0.019938f
C4037 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_5.LD 1.1e-20
C4038 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.00989f
C4039 p3_gen_magic_0.xnor_magic_4.OUT a_11292_n6613# 0.318049f
C4040 a_11279_8697# a_12387_8536# 0.001529f
C4041 a_15865_4557# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 0.149276f
C4042 divide_by_2_1.tg_magic_1.IN mux_magic_0.OR_magic_0.B 9.17e-20
C4043 a_15865_1059# Q5 0.001903f
C4044 a_12387_8536# D2_2 0.01192f
C4045 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A 0.001081f
C4046 Q2 D2_6 0.250294f
C4047 D2_2 Q5 0.122757f
C4048 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_8740# 0.431521f
C4049 a_15865_7470# VDD 0.821356f
C4050 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8955_4557# 9.27e-19
C4051 p3_gen_magic_0.3_inp_AND_magic_0.C Q4 0.161047f
C4052 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8643_n6024# 0.082959f
C4053 a_1209_9773# CLK 6.34e-19
C4054 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 8.54e-19
C4055 a_5385_1059# Q6 0.036115f
C4056 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B VDD 1.21143f
C4057 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A Q1 9.62e-19
C4058 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B P2 7.78e-21
C4059 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT 2.29e-19
C4060 7b_counter_0.MDFF_4.LD a_17405_3524# 0.001152f
C4061 a_12931_4557# CLK 0.009154f
C4062 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VDD 1.2623f
C4063 a_15865_7470# D2_1 0.258263f
C4064 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n3597# 0.083042f
C4065 7b_counter_0.MDFF_4.tspc2_magic_0.D Q1 0.003739f
C4066 a_5036_n3150# a_5452_n3150# 0.002223f
C4067 a_12174_n3597# Q4 0.092097f
C4068 a_13353_n2115# VDD 1.13805f
C4069 VDD D2_3 5.80874f
C4070 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.240827f
C4071 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A a_23258_575# 0.149276f
C4072 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A 0.007053f
C4073 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A 0.00221f
C4074 p2_gen_magic_0.xnor_magic_1.OUT Q5 0.003619f
C4075 a_15865_1059# D2_4 0.02504f
C4076 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT Q3 0.137714f
C4077 a_5054_n1042# Q6 0.00443f
C4078 divide_by_2_0.tg_magic_3.OUT a_23352_n6798# 1.86e-20
C4079 a_12387_9730# CLK 6.58e-19
C4080 a_1541_n7648# p3_gen_magic_0.xnor_magic_1.OUT 0.093718f
C4081 a_1209_3363# a_1209_2253# 0.003291f
C4082 D2_1 D2_3 2.17246f
C4083 D2_2 D2_4 0.084075f
C4084 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VDD 1.40826f
C4085 a_8523_n8095# D2_5 0.001848f
C4086 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 0.178114f
C4087 a_15865_9774# VDD 0.927898f
C4088 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B LD 0.001212f
C4089 p3_gen_magic_0.3_inp_AND_magic_0.VOUT VDD 2.05341f
C4090 a_9689_1669# Q1 0.00186f
C4091 a_8713_6842# Q7 0.005475f
C4092 a_1209_4557# D2_5 2.51e-19
C4093 p3_gen_magic_0.xnor_magic_5.OUT Q4 0.064085f
C4094 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK a_16386_n8142# 0.015981f
C4095 a_15865_9774# D2_1 0.003239f
C4096 a_12387_9730# a_11191_10149# 0.002003f
C4097 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.178114f
C4098 p3_gen_magic_0.3_inp_AND_magic_0.VOUT D2_1 0.008654f
C4099 p2_gen_magic_0.xnor_magic_1.OUT D2_4 0.248313f
C4100 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK 0.009273f
C4101 LD D2_3 0.016736f
C4102 a_1209_1059# Q4 0.25171f
C4103 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT Q6 0.006508f
C4104 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B VDD 1.23782f
C4105 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n3150# 0.004631f
C4106 p2_gen_magic_0.3_inp_AND_magic_0.B Q5 6.77e-20
C4107 Q2 D2_2 0.253881f
C4108 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n8095# 0.063777f
C4109 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_5 0.010265f
C4110 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A LD 0.43461f
C4111 a_15865_7470# a_16065_6276# 0.003083f
C4112 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_1.tspc2_magic_0.Q 0.268721f
C4113 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q4 6.58e-19
C4114 7b_counter_0.MDFF_0.tspc2_magic_0.CLK 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 0.003149f
C4115 7b_counter_0.MDFF_5.tspc2_magic_0.Q Q2 0.289359f
C4116 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 7b_counter_0.MDFF_3.tspc2_magic_0.Q 0.018858f
C4117 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VDD 1.23136f
C4118 DFF_magic_0.D a_27778_2253# 0.002281f
C4119 a_15865_9774# LD 4.93e-19
C4120 p2_gen_magic_0.xnor_magic_6.OUT p3_gen_magic_0.3_inp_AND_magic_0.C 1.02e-19
C4121 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B VDD 1.20994f
C4122 a_16065_8580# CLK 0.14486f
C4123 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT P2 1.48e-19
C4124 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A Q7 0.024313f
C4125 7b_counter_0.NAND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.C 0.15193f
C4126 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 2.29e-19
C4127 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8643_n5540# 1.08e-19
C4128 p2_gen_magic_0.xnor_magic_1.OUT Q2 0.018066f
C4129 p3_gen_magic_0.xnor_magic_0.OUT a_11492_n6613# 0.075783f
C4130 7b_counter_0.MDFF_0.tspc2_magic_0.D a_4496_4393# 0.038362f
C4131 a_8523_n7648# VDD 0.001396f
C4132 p2_gen_magic_0.3_inp_AND_magic_0.B D2_4 0.002083f
C4133 p2_gen_magic_0.xnor_magic_6.OUT a_12174_n3597# 0.02352f
C4134 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VDD 1.31418f
C4135 a_12387_8536# CLK 0.26404f
C4136 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT p2_gen_magic_0.xnor_magic_5.OUT 5.85e-19
C4137 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C4138 Q1 D2_5 0.214328f
C4139 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23802_1059# 0.128771f
C4140 CLK Q5 0.219314f
C4141 a_17405_4932# D2_3 0.002473f
C4142 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.xnor_magic_5.OUT 0.004328f
C4143 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 9.4e-20
C4144 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B D2_3 0.005637f
C4145 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VDD 1.00398f
C4146 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B D2_7 0.002402f
C4147 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.001081f
C4148 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A D2_1 3.54e-19
C4149 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_5.OUT 0.171314f
C4150 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT Q3 0.091469f
C4151 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A LD 5.51e-19
C4152 a_7215_10149# a_7303_8697# 0.479729f
C4153 a_12931_8580# D2_2 0.040136f
C4154 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT a_30365_4922# 2.63e-19
C4155 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_6.OUT 0.037167f
C4156 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A a_7303_8697# 0.036613f
C4157 Q3 D2_3 1.97584f
C4158 a_13353_n2115# Q3 0.006483f
C4159 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN D2_1 0.007522f
C4160 a_11191_10149# a_12387_8536# 7.51e-20
C4161 a_8643_n5540# Q1 0.013687f
C4162 7b_counter_0.3_inp_AND_magic_0.A a_23985_7877# 0.397303f
C4163 7b_counter_0.3_inp_AND_magic_0.B 7b_counter_0.3_inp_AND_magic_0.C 0.337623f
C4164 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q5 5.67e-19
C4165 a_8955_3363# D2_6 0.134719f
C4166 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A a_27234_4513# 0.149276f
C4167 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_15865_7470# 5.28e-20
C4168 DFF_magic_0.tg_magic_2.OUT P2 0.01392f
C4169 a_14756_n8142# Q4 0.035148f
C4170 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.270406f
C4171 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_2749_10148# 0.189314f
C4172 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A LD 6.12e-19
C4173 a_12387_6986# VDD 0.807353f
C4174 CLK D2_4 0.924842f
C4175 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_27778_1059# 9.27e-19
C4176 7b_counter_0.MDFF_0.tspc2_magic_0.CLK a_5185_2253# 4.65e-19
C4177 a_5185_1059# Q6 0.056229f
C4178 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.12429f
C4179 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_7215_4932# 0.414018f
C4180 a_1209_3363# CLK 0.002302f
C4181 7b_counter_0.MDFF_4.LD a_12931_4557# 0.004065f
C4182 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B a_8411_4513# 1.93e-19
C4183 7b_counter_0.MDFF_6.tspc2_magic_0.CLK D2_3 0.493301f
C4184 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A 0.00112f
C4185 p2_gen_magic_0.xnor_magic_3.OUT a_12174_n3150# 4.14e-19
C4186 a_22150_1124# a_23258_575# 7.54e-20
C4187 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.024392f
C4188 7b_counter_0.3_inp_AND_magic_0.B Q7 0.265346f
C4189 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.019552f
C4190 7b_counter_0.MDFF_6.tspc2_magic_0.D Q1 3.55e-19
C4191 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_5385_7469# 0.016967f
C4192 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.003202f
C4193 a_5515_3947# a_5385_2253# 0.005699f
C4194 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A a_12387_4513# 1.27e-19
C4195 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_17405_3524# 0.036613f
C4196 7b_counter_0.MDFF_0.tspc2_magic_0.Q D2_4 6.84e-19
C4197 a_22062_684# D2_4 0.021305f
C4198 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B Q3 0.004694f
C4199 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q4 0.313059f
C4200 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN 5.37e-19
C4201 a_8523_n4081# p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 1.09e-19
C4202 7b_counter_0.MDFF_3.tspc2_magic_0.CLK D2_7 0.065845f
C4203 OR_magic_1.VOUT CLK 0.015396f
C4204 OR_magic_1.VOUT divide_by_2_1.tg_magic_1.IN 0.69947f
C4205 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 5.37e-19
C4206 a_9212_5956# VDD 0.97511f
C4207 divide_by_2_1.tg_magic_1.IN mux_magic_0.OR_magic_0.A 0.002507f
C4208 CLK Q2 0.389788f
C4209 a_15865_9774# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 1.63e-20
C4210 a_5036_n8095# D2_5 5.71e-19
C4211 a_1409_2253# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 1.77e-19
C4212 a_19152_1223# D2_3 2.21e-19
C4213 a_13353_n6613# VDD 1.14073f
C4214 a_32816_n1264# a_32816_n2458# 0.020635f
C4215 a_12387_1769# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 0.001158f
C4216 a_2749_5900# Q7 0.002935f
C4217 a_8825_1669# Q1 0.007085f
C4218 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 8.78e-21
C4219 a_19152_6440# a_19152_5956# 0.014143f
C4220 DFF_magic_0.tg_magic_2.OUT VDD 1.25471f
C4221 a_12387_1769# a_11191_684# 7.51e-20
C4222 a_5054_n5540# Q6 0.044657f
C4223 7b_counter_0.MDFF_1.tspc2_magic_0.CLK Q1 0.045202f
C4224 7b_counter_0.NAND_magic_0.A D2_4 0.113315f
C4225 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_11279_6341# 0.429153f
C4226 a_1541_n3150# D2_4 0.041124f
C4227 a_13353_n6613# D2_1 0.006442f
C4228 p2_gen_magic_0.xnor_magic_5.OUT D2_3 0.132137f
C4229 a_8411_8536# a_8955_8580# 0.297401f
C4230 p3_gen_magic_0.xnor_magic_6.OUT a_8523_n8579# 0.465726f
C4231 a_7303_3480# a_8411_3319# 0.001529f
C4232 p3_gen_magic_0.3_inp_AND_magic_0.B p3_gen_magic_0.AND2_magic_1.A 0.007712f
C4233 p2_gen_magic_0.xnor_magic_4.OUT Q1 0.366591f
C4234 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_8713_1625# 0.515029f
C4235 DFF_magic_0.tg_magic_2.OUT D2_1 0.002247f
C4236 a_2749_3524# 7b_counter_0.MDFF_0.tspc2_magic_0.D 0.134004f
C4237 7b_counter_0.MDFF_7.tspc2_magic_0.CLK Q4 0.001101f
C4238 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1541_n3597# 0.063777f
C4239 a_11279_1124# a_8713_1625# 6.34e-20
C4240 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT a_16186_n3644# 8.76e-20
C4241 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_8411_8536# 4.65e-19
C4242 a_15865_7470# a_15865_6276# 0.005574f
C4243 a_11292_n2115# Q4 0.020773f
C4244 a_17405_8741# VDD 0.941683f
C4245 a_8411_9730# Q2 7.66e-19
C4246 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_4235_9163# 0.671058f
C4247 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 0.434645f
C4248 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.3_inp_AND_magic_0.VOUT 1.99e-23
C4249 a_7303_3480# VDD 0.942239f
C4250 7b_counter_0.MDFF_4.tspc2_magic_0.CLK a_9412_739# 0.365826f
C4251 a_12931_8580# CLK 0.139116f
C4252 a_11279_1124# a_9412_739# 1.39e-20
C4253 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VDD 1.23928f
C4254 7b_counter_0.NAND_magic_0.A Q2 1.46e-19
C4255 a_17405_8741# D2_1 0.035246f
C4256 a_8411_3319# a_8713_1625# 3.03e-19
C4257 a_15865_6276# D2_3 0.00245f
C4258 p3_gen_magic_0.xnor_magic_0.OUT a_9059_n6471# 0.077312f
C4259 a_5452_n7648# VDD 0.004613f
C4260 a_2749_3524# a_4496_4393# 7.92e-19
C4261 a_8411_4513# Q7 0.005173f
C4262 7b_counter_0.DFF_magic_0.tg_magic_1.IN 7b_counter_0.DFF_magic_0.tg_magic_0.IN 0.311939f
C4263 p2_gen_magic_0.xnor_magic_6.OUT a_8523_n3597# 0.371622f
C4264 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A D2_1 3.01e-19
C4265 a_17405_7309# a_19152_5956# 1.39e-20
C4266 7b_counter_0.NAND_magic_0.A a_24003_10051# 0.098209f
C4267 a_19841_4557# D2_3 5.4e-19
C4268 7b_counter_0.MDFF_4.LD Q5 2.49055f
C4269 a_5036_n8095# D2_7 0.252183f
C4270 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.090266f
C4271 a_5385_7469# D2_7 0.128625f
C4272 a_13769_n6613# VDD 0.019499f
C4273 a_19152_6440# VDD 0.770257f
C4274 p2_gen_magic_0.xnor_magic_0.OUT D2_6 0.200519f
C4275 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n3150# 0.107246f
C4276 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q5 0.134657f
C4277 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_27234_3319# 0.001158f
C4278 a_8713_1625# VDD 0.76217f
C4279 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 2.64e-19
C4280 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A D2_3 0.029243f
C4281 a_1409_6275# Q6 0.138643f
C4282 a_16065_4557# a_16065_3363# 0.020635f
C4283 a_19152_6440# D2_1 4.14e-19
C4284 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A D2_6 0.105789f
C4285 a_5515_9163# Q7 2.52e-19
C4286 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A LD 5.51e-19
C4287 a_12931_1059# Q5 4.49e-19
C4288 a_5054_n1042# a_5054_n1526# 0.033537f
C4289 a_9412_739# VDD 0.725398f
C4290 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.C 0.410203f
C4291 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT D2_6 0.001135f
C4292 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.247535f
C4293 a_14756_n3644# D2_3 0.026553f
C4294 7b_counter_0.MDFF_4.LD D2_4 0.84277f
C4295 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B a_17405_2092# 0.431521f
C4296 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.164969f
C4297 a_19307_1669# a_20171_1669# 0.009722f
C4298 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_4 2.86e-19
C4299 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_0.IN 0.311939f
C4300 a_23352_n6798# CLK 7.74e-20
C4301 a_15865_2253# a_17405_2092# 0.001529f
C4302 p2_gen_magic_0.3_inp_AND_magic_0.A D2_5 0.006558f
C4303 a_11292_n2115# p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.010995f
C4304 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B Q7 0.037595f
C4305 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_19841_8580# 0.146237f
C4306 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A Q1 0.00816f
C4307 a_11292_n2115# p2_gen_magic_0.xnor_magic_6.OUT 0.022681f
C4308 7b_counter_0.MDFF_3.tspc2_magic_0.Q a_2749_7308# 0.001371f
C4309 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD 1.17663f
C4310 a_12931_1059# D2_4 0.003809f
C4311 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 0.001447f
C4312 a_1957_n3150# Q7 0.003349f
C4313 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.252157f
C4314 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN D2_6 0.010053f
C4315 7b_counter_0.MDFF_4.LD OR_magic_1.VOUT 0.002996f
C4316 a_17405_7309# VDD 0.94863f
C4317 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q4 0.001088f
C4318 a_12931_2253# 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A 0.001034f
C4319 a_7303_3480# a_6725_2092# 1.63e-19
C4320 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 0.001081f
C4321 a_4496_9609# a_5515_9163# 0.043767f
C4322 a_15865_9774# a_16065_9774# 0.29829f
C4323 7b_counter_0.MDFF_4.LD Q2 0.203409f
C4324 a_1209_2253# 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A 0.001985f
C4325 a_8939_n7648# D2_6 0.005701f
C4326 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1409_6275# 9.27e-19
C4327 a_12590_n7648# D2_5 0.008738f
C4328 a_18891_1669# D2_3 0.03354f
C4329 7b_counter_0.MDFF_7.tspc2_magic_0.CLK a_27234_4513# 1.37e-19
C4330 p2_gen_magic_0.xnor_magic_0.OUT D2_2 0.224346f
C4331 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q2 0.00597f
C4332 a_17405_7309# D2_1 0.046434f
C4333 a_12387_9730# 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 1.63e-20
C4334 7b_counter_0.MDFF_3.QB CLK 0.006789f
C4335 a_18891_6886# a_19152_5956# 0.655098f
C4336 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.270406f
C4337 a_6725_7308# Q7 0.175844f
C4338 7b_counter_0.MDFF_0.tspc2_magic_0.CLK Q6 0.023077f
C4339 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_4.OUT 8.59e-20
C4340 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK a_16186_n8142# 0.003314f
C4341 a_16065_4557# Q1 6.2e-19
C4342 a_21381_4932# a_21381_3524# 0.479729f
C4343 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C4344 a_12387_6986# 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.001985f
C4345 a_2749_5900# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 4.23e-19
C4346 a_5036_n3150# D2_3 1.85e-19
C4347 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A D2_2 0.002719f
C4348 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VDD 1.08682f
C4349 a_2749_4932# 7b_counter_0.MDFF_0.tspc2_magic_0.D 1.08e-19
C4350 a_21381_3524# Q4 0.004617f
C4351 a_8643_n6024# a_9059_n6471# 0.011514f
C4352 7b_counter_0.MDFF_7.tspc2_magic_0.CLK 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A 8.78e-21
C4353 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.027154f
C4354 a_6725_2092# a_8713_1625# 0.001527f
C4355 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B a_11292_n2115# 1.08e-19
C4356 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B a_12387_5792# 1.93e-19
C4357 a_17405_8741# 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 0.132169f
C4358 a_12931_9774# VDD 0.056754f
C4359 a_6725_7308# a_5185_6275# 7.54e-20
C4360 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_4496_10093# 0.365826f
C4361 a_8713_1625# Q3 8.58e-20
C4362 p2_gen_magic_0.xnor_magic_5.OUT a_13353_n6613# 6.92e-21
C4363 a_8713_6842# a_9212_5956# 0.301553f
C4364 a_19841_8580# a_20041_8580# 0.297401f
C4365 p3_gen_magic_0.xnor_magic_4.OUT Q1 0.340402f
C4366 a_1541_n8579# Q7 1.41e-19
C4367 p3_gen_magic_0.xnor_magic_0.OUT a_8643_n6471# 0.292076f
C4368 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C4369 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.3_inp_AND_magic_0.VOUT 0.795803f
C4370 a_8523_n3150# a_8523_n3597# 0.014233f
C4371 a_12174_n3150# p2_gen_magic_0.AND2_magic_1.A 0.09365f
C4372 a_11292_n6613# Q4 4.41e-19
C4373 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT 3.44e-20
C4374 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 0.022357f
C4375 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT CLK 0.007327f
C4376 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_19152_6440# 0.514788f
C4377 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.3_inp_AND_magic_0.B 9.01e-19
C4378 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.3_inp_AND_magic_0.A 0.003345f
C4379 a_13553_n6613# VDD 0.017725f
C4380 a_18891_6886# VDD 0.977068f
C4381 a_2749_7308# D2_7 0.036293f
C4382 a_27234_4513# a_27234_3319# 0.005574f
C4383 7b_counter_0.MDFF_5.tspc2_magic_0.CLK a_12387_8536# 1.18e-19
C4384 a_17405_10149# a_15865_8580# 7.51e-20
C4385 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B a_15865_8580# 0.146237f
C4386 a_1209_6275# Q6 0.286048f
C4387 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q5 0.023553f
C4388 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B Q7 0.007212f
C4389 p3_gen_magic_0.P3 a_23352_n6798# 0.349803f
C4390 a_17405_7309# 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 1e-20
C4391 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT Q3 9.74e-19
C4392 a_4651_9163# Q7 1.22e-19
C4393 a_18891_6886# D2_1 0.028916f
C4394 p2_gen_magic_0.xnor_magic_0.OUT a_11708_n2115# 0.02473f
C4395 a_12387_575# Q5 0.001903f
C4396 a_8643_n1526# D2_6 0.016846f
C4397 a_14556_n8142# Q4 0.033942f
C4398 a_9212_5956# 7b_counter_0.MDFF_4.tspc2_magic_0.Q 6.28e-20
C4399 a_5385_1059# VDD 0.109184f
C4400 7b_counter_0.NAND_magic_0.A a_23985_7877# 0.001516f
C4401 p2_gen_magic_0.3_inp_AND_magic_0.C p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT 0.009577f
C4402 a_11279_6341# 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B 1e-20
C4403 p3_gen_magic_0.xnor_magic_0.OUT D2_6 0.01556f
C4404 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q5 0.001402f
C4405 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_3.OUT 7.62e-20
C4406 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9689_1669# 0.004574f
C4407 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN 0.345544f
C4408 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A 0.00112f
C4409 a_5054_n6024# p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT 7.12e-21
C4410 a_1409_1059# Q7 0.010048f
C4411 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A D2_4 0.006661f
C4412 a_12590_n3150# Q4 0.003399f
C4413 7b_counter_0.NAND_magic_0.A 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.00184f
C4414 a_5054_n1042# VDD 0.505153f
C4415 p3_gen_magic_0.xnor_magic_4.OUT a_5036_n8095# 0.016433f
C4416 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 0.008125f
C4417 DFF_magic_0.tg_magic_2.OUT mux_magic_0.AND2_magic_0.A 1.68e-20
C4418 p2_gen_magic_0.xnor_magic_3.OUT Q5 0.097028f
C4419 a_12387_575# D2_4 0.025118f
C4420 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_26126_1124# 1.23e-19
C4421 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_17405_7309# 0.018983f
C4422 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n7648# 0.011524f
C4423 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A a_13353_n2115# 1.84e-20
C4424 a_19841_3363# CLK 0.001414f
C4425 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A D2_3 0.002265f
C4426 7b_counter_0.MDFF_4.LD a_8955_3363# 0.036926f
C4427 a_19841_9774# 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B 1.93e-19
C4428 OR_magic_1.VOUT divide_by_2_1.tg_magic_3.IN 0.635475f
C4429 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1957_n7648# 6.1e-19
C4430 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT D2_4 0.007574f
C4431 a_5385_1059# LD 1.1e-19
C4432 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A a_17405_8741# 2.07e-19
C4433 a_8955_8580# Q2 5.02e-19
C4434 a_4496_9609# a_4651_9163# 0.240883f
C4435 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5470_n1973# 6.1e-19
C4436 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A a_1209_6275# 0.149276f
C4437 p3_gen_magic_0.3_inp_AND_magic_0.A D2_5 0.060291f
C4438 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 7b_counter_0.MDFF_1.tspc2_magic_0.D 0.423451f
C4439 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 0.178114f
C4440 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VDD 1.18058f
C4441 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_16065_1059# 0.037614f
C4442 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A a_27234_575# 0.149276f
C4443 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A Q2 0.002402f
C4444 7b_counter_0.MDFF_5.tspc2_magic_0.CLK Q2 0.237309f
C4445 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT CLK 1.36181f
C4446 a_34156_n889# a_34156_n2297# 0.479729f
C4447 a_12387_6986# a_11279_6341# 0.001529f
C4448 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VDD 1.07323f
C4449 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p2_gen_magic_0.AND2_magic_1.A 0.258463f
C4450 p2_gen_magic_0.xnor_magic_3.OUT D2_4 0.199174f
C4451 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT D2_1 7.09e-19
C4452 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A 0.007064f
C4453 a_8643_n1526# D2_2 0.236724f
C4454 a_19152_6440# a_19841_4557# 1.73e-19
C4455 a_2749_4932# a_2749_3524# 0.479729f
C4456 a_8643_n6024# a_8643_n6471# 0.013685f
C4457 p2_gen_magic_0.xnor_magic_3.OUT a_1559_n1042# 0.457196f
C4458 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN CLK 0.016792f
C4459 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 0.024279f
C4460 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q2 0.00597f
C4461 p3_gen_magic_0.xnor_magic_0.OUT D2_2 0.153546f
C4462 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_1.IN 4.63e-20
C4463 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 0.001081f
C4464 a_12387_6986# a_12931_6276# 0.00152f
C4465 a_22991_5885# a_23207_5885# 0.901612f
C4466 a_1209_8579# VDD 0.807784f
C4467 7b_counter_0.MDFF_4.tspc2_magic_0.Q a_8713_1625# 0.012528f
C4468 a_8643_n1973# Q5 6.4e-19
C4469 a_6725_7308# 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A 2.4e-20
C4470 a_11279_6341# a_9212_5956# 8.2e-19
C4471 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A Q6 3.87e-19
C4472 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_6725_5900# 0.189314f
C4473 a_1559_n1973# p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 1.81e-19
C4474 p2_gen_magic_0.xnor_magic_3.OUT Q2 0.863413f
C4475 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_0.OUT 1.35e-19
C4476 a_24401_7877# Q5 4.38e-20
C4477 p2_gen_magic_0.3_inp_AND_magic_0.C a_13353_n2115# 0.536475f
C4478 p2_gen_magic_0.xnor_magic_6.OUT a_12590_n3150# 0.002939f
C4479 p2_gen_magic_0.3_inp_AND_magic_0.C D2_3 0.294866f
C4480 DFF_magic_0.tg_magic_2.OUT DFF_magic_0.tg_magic_0.IN 0.010522f
C4481 7b_counter_0.MDFF_5.LD a_8955_9774# 1.1e-19
C4482 divide_by_2_0.tg_magic_2.IN VDD 1.0449f
C4483 7b_counter_0.NAND_magic_0.A 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.001908f
C4484 7b_counter_0.MDFF_6.tspc2_magic_0.D 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 8.78e-21
C4485 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT D2_3 3.28e-19
C4486 a_17405_7309# a_15865_6276# 7.54e-20
C4487 7b_counter_0.MDFF_6.tspc2_magic_0.CLK a_18891_6886# 0.671058f
C4488 divide_by_2_0.tg_magic_1.IN divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 0.240827f
C4489 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT CLK 2.41e-19
C4490 p2_gen_magic_0.xnor_magic_4.OUT a_8643_n1042# 0.387036f
C4491 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A a_1209_8579# 0.001158f
C4492 7b_counter_0.MDFF_0.tspc2_magic_0.Q 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 0.27167f
C4493 a_8643_n6024# D2_6 7.09e-20
C4494 a_11191_5901# VDD 1.55477f
C4495 a_11708_n6613# VDD 0.012593f
C4496 p3_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.AND2_magic_1.A 0.001148f
C4497 a_1209_8579# LD 0.224216f
C4498 a_11279_3480# D2_6 0.006161f
C4499 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT D2_7 0.023985f
C4500 7b_counter_0.MDFF_4.tspc2_magic_0.Q p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 1.76e-20
C4501 a_21381_10149# Q7 0.017818f
C4502 a_24401_7877# D2_4 0.005636f
C4503 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A D2_6 0.002317f
C4504 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT Q4 0.004092f
C4505 p2_gen_magic_0.xnor_magic_0.OUT a_11492_n2115# 0.075783f
C4506 a_12174_n8095# Q4 0.095437f
C4507 a_5185_1059# VDD 0.93919f
C4508 7b_counter_0.3_inp_AND_magic_0.B a_19152_6440# 8.75e-21
C4509 a_14556_n3644# D2_3 0.026286f
C4510 a_5054_n5540# a_5054_n6024# 0.033537f
C4511 p3_gen_magic_0.xnor_magic_1.OUT Q5 0.076958f
C4512 7b_counter_0.MDFF_4.tspc2_magic_0.D a_8825_1669# 2.1e-20
C4513 a_23258_1769# D2_4 0.244434f
C4514 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B D2_3 0.002402f
C4515 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_0.IN 0.010522f
C4516 a_1209_1059# Q7 0.044482f
C4517 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A CLK 0.020275f
C4518 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.AND2_magic_1.A 2.36e-19
C4519 a_15865_4557# a_17405_3524# 7.54e-20
C4520 a_27778_2253# D2_4 0.040136f
C4521 Q6 D2_6 0.068021f
C4522 7b_counter_0.MDFF_5.LD 7b_counter_0.3_inp_AND_magic_0.C 0.001107f
C4523 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.43461f
C4524 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q7 0.117721f
C4525 7b_counter_0.MDFF_4.LD a_19841_3363# 0.224142f
C4526 a_27778_4557# CLK 3.73e-20
C4527 a_1409_4557# a_1209_3363# 0.003083f
C4528 a_8825_1669# a_9689_1669# 0.009722f
C4529 7b_counter_0.3_inp_AND_magic_0.A a_23793_5904# 0.898684f
C4530 a_5185_1059# LD 3.96e-19
C4531 a_19841_8580# Q2 1.57e-20
C4532 7b_counter_0.MDFF_3.tspc2_magic_0.D 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.423451f
C4533 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n1973# 0.107012f
C4534 7b_counter_0.MDFF_0.tspc2_magic_0.Q a_5185_2253# 0.029386f
C4535 a_8643_n5540# D2_5 0.001584f
C4536 a_8643_n6024# D2_2 0.245196f
C4537 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.MDFF_7.tspc2_magic_0.D 3.94e-20
C4538 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.168057f
C4539 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B a_22150_1124# 0.431521f
C4540 a_9212_739# Q1 0.007967f
C4541 a_11279_3480# D2_2 0.125313f
C4542 a_5054_n5540# VDD 0.50544f
C4543 a_8411_4513# a_7303_3480# 7.54e-20
C4544 a_26126_1124# a_27234_575# 7.54e-20
C4545 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_5 0.007322f
C4546 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A a_15865_1059# 0.279825f
C4547 p3_gen_magic_0.xnor_magic_3.OUT Q5 5.14e-19
C4548 7b_counter_0.MDFF_5.LD Q7 2.36751f
C4549 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B Q2 8.23e-19
C4550 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 6.05e-21
C4551 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.xnor_magic_6.OUT 0.029015f
C4552 7b_counter_0.MDFF_3.tspc2_magic_0.Q D2_7 0.170444f
C4553 a_11292_n6613# p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.010943f
C4554 a_12174_n4081# D2_2 0.001215f
C4555 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A a_1209_4557# 0.279825f
C4556 OR_magic_2.A DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7.58e-20
C4557 a_19841_9774# a_20041_9774# 0.29829f
C4558 7b_counter_0.DFF_magic_0.tg_magic_2.IN OR_magic_2.A 2.96e-20
C4559 a_12387_6986# a_12387_5792# 0.005574f
C4560 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VDD 1.32361f
C4561 p2_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 1.33e-20
C4562 p3_gen_magic_0.xnor_magic_3.OUT D2_4 0.222873f
C4563 a_6725_2092# a_5185_1059# 7.54e-20
C4564 D2_7 D2_5 0.556163f
C4565 a_20171_6886# D2_3 4.43e-19
C4566 a_24185_7877# Q5 2.88e-19
C4567 D2_2 Q6 0.058991f
C4568 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 2.24e-19
C4569 a_5452_n3150# a_5036_n3597# 0.013021f
C4570 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A a_1409_8579# 1.77e-19
C4571 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.003202f
C4572 a_5185_1059# Q3 2.32e-19
C4573 a_23802_2253# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 5.46e-20
C4574 7b_counter_0.MDFF_5.tspc2_magic_0.Q Q6 0.026528f
C4575 7b_counter_0.DFF_magic_0.tg_magic_3.OUT D2_4 0.009728f
C4576 mux_magic_0.OR_magic_0.B a_34156_n2297# 0.431521f
C4577 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT D2_4 0.167041f
C4578 a_1409_6275# VDD 0.058805f
C4579 a_11492_n6613# VDD 0.014256f
C4580 p3_gen_magic_0.xnor_magic_1.OUT a_1541_n8095# 0.37449f
C4581 p3_gen_magic_0.xnor_magic_5.OUT p3_gen_magic_0.xnor_magic_6.OUT 0.980813f
C4582 a_4235_9163# 7b_counter_0.MDFF_3.tspc2_magic_0.Q 1.94e-20
C4583 p2_gen_magic_0.xnor_magic_4.OUT D2_5 0.09813f
C4584 a_11191_4932# D2_6 0.001168f
C4585 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT 0.026342f
C4586 p2_gen_magic_0.xnor_magic_1.OUT Q6 0.035855f
C4587 p3_gen_magic_0.xnor_magic_3.OUT Q2 0.288947f
C4588 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A Q7 0.021228f
C4589 p3_gen_magic_0.3_inp_AND_magic_0.C D2_3 0.024995f
C4590 a_24185_7877# D2_4 0.003198f
C4591 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT mux_magic_0.IN1 6.97e-20
C4592 7b_counter_0.DFF_magic_0.tg_magic_0.IN CLK 0.639804f
C4593 a_20171_1669# Q5 6.75e-20
C4594 p2_gen_magic_0.xnor_magic_0.OUT a_9059_n1973# 0.077312f
C4595 a_12387_3319# D2_6 4e-19
C4596 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A Q5 8.66e-19
C4597 7b_counter_0.MDFF_0.tspc2_magic_0.D a_1209_3363# 7.57e-20
C4598 a_17405_2092# D2_3 0.041889f
C4599 a_8523_n4081# D2_6 0.007723f
C4600 a_1541_n7648# Q5 0.685195f
C4601 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q2 0.00334f
C4602 p3_gen_magic_0.3_inp_AND_magic_0.C p3_gen_magic_0.3_inp_AND_magic_0.VOUT 0.796727f
C4603 mux_magic_0.OR_magic_0.A a_32816_n1264# 9.27e-19
C4604 a_1409_6275# LD 0.003655f
C4605 DFF_magic_0.tg_magic_2.IN CLK 0.001114f
C4606 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 0.445787f
C4607 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_1.OUT 0.001317f
C4608 7b_counter_0.DFF_magic_0.tg_magic_1.IN VDD 1.89471f
C4609 p3_gen_magic_0.xnor_magic_4.OUT p3_gen_magic_0.3_inp_AND_magic_0.A 0.003345f
C4610 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.3_inp_AND_magic_0.B 9.01e-19
C4611 a_20171_1669# D2_4 0.001536f
C4612 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A a_17405_684# 0.414018f
C4613 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A CLK 0.002994f
C4614 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q4 0.005777f
C4615 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B a_2749_684# 0.189314f
C4616 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A a_11191_5901# 0.414018f
C4617 a_15865_3363# CLK 0.264578f
C4618 7b_counter_0.MDFF_4.LD a_27778_4557# 0.003068f
C4619 OR_magic_2.A CLK 0.516087f
C4620 a_2749_8740# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.018983f
C4621 a_1541_n7648# D2_4 2.58e-19
C4622 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VDD 1.00053f
C4623 7b_counter_0.MDFF_0.tspc2_magic_0.CLK VDD 2.47953f
C4624 7b_counter_0.MDFF_5.tspc2_magic_0.CLK 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.006642f
C4625 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5470_n6471# 6.1e-19
C4626 p2_gen_magic_0.xnor_magic_4.OUT D2_7 0.333879f
C4627 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A Q3 0.08528f
C4628 a_11191_4932# D2_2 0.043904f
C4629 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT 0.001724f
C4630 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B Q6 0.012347f
C4631 a_21381_4932# Q1 0.052391f
C4632 a_19841_9774# Q2 6.82e-19
C4633 a_7303_8697# Q7 0.049781f
C4634 a_6725_684# Q5 0.018493f
C4635 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT a_12174_n3150# 0.00871f
C4636 a_21381_8741# a_19841_8580# 0.001529f
C4637 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT Q7 0.036448f
C4638 p3_gen_magic_0.xnor_magic_6.OUT a_14756_n8142# 0.128771f
C4639 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 2.64e-19
C4640 a_12387_3319# D2_2 0.010654f
C4641 7b_counter_0.MDFF_5.LD a_15865_7470# 0.224216f
C4642 Q1 Q4 0.050579f
C4643 CLK Q6 0.130441f
C4644 a_4235_9163# D2_7 0.033531f
C4645 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_3.OUT 0.041842f
C4646 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT divide_by_2_0.tg_magic_3.IN 0.304333f
C4647 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A a_21381_10149# 0.414018f
C4648 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN a_16386_n8142# 2.98e-19
C4649 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 1.55e-19
C4650 a_23985_7877# a_24401_7877# 0.278913f
C4651 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B VDD 1.19364f
C4652 a_19152_739# VDD 0.725398f
C4653 7b_counter_0.MDFF_5.LD D2_3 0.272049f
C4654 7b_counter_0.MDFF_0.tspc2_magic_0.CLK LD 0.08472f
C4655 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B a_12387_4513# 1.93e-19
C4656 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q6 0.287712f
C4657 a_6725_684# D2_4 0.007364f
C4658 a_1559_n1526# p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 6.69e-21
C4659 a_19307_6886# D2_3 0.003363f
C4660 a_23207_5885# Q5 4.56e-20
C4661 DFF_magic_0.D D2_4 0.040521f
C4662 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 9.4e-20
C4663 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1541_n4081# 0.066064f
C4664 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A 0.001081f
C4665 7b_counter_0.MDFF_5.LD a_15865_9774# 0.031272f
C4666 a_7303_8697# a_4496_9609# 0.001517f
C4667 a_8411_9730# Q6 3.01e-19
C4668 mux_magic_0.OR_magic_0.B a_34156_n889# 0.189314f
C4669 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VDD 1.09731f
C4670 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 0.207107f
C4671 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.OUT 0.200659f
C4672 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT 0.003851f
C4673 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT 7.81e-19
C4674 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A D2_6 0.002294f
C4675 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 0.178114f
C4676 a_9059_n6471# VDD 0.001798f
C4677 a_1209_6275# VDD 0.931274f
C4678 a_1541_n7648# a_1541_n8095# 0.004574f
C4679 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT CLK 0.343704f
C4680 7b_counter_0.NAND_magic_0.A Q6 1.47e-19
C4681 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B LD 0.004701f
C4682 p3_gen_magic_0.xnor_magic_3.OUT a_1559_n5540# 0.457196f
C4683 a_20041_3363# D2_3 0.128625f
C4684 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VDD 1.18466f
C4685 7b_counter_0.MDFF_6.tspc2_magic_0.D 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 2.05e-19
C4686 a_1541_n3150# Q6 0.001916f
C4687 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A CLK 0.004331f
C4688 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27778_1059# 0.037614f
C4689 DFF_magic_0.D OR_magic_1.VOUT 0.00188f
C4690 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B Q7 0.006977f
C4691 p2_gen_magic_0.xnor_magic_0.OUT a_8643_n1973# 0.292076f
C4692 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT D2_1 0.08204f
C4693 7b_counter_0.MDFF_4.LD 7b_counter_0.DFF_magic_0.tg_magic_0.IN 5.63e-20
C4694 a_2749_3524# a_1209_3363# 0.001529f
C4695 mux_magic_0.OR_magic_0.A a_32816_n2458# 1.77e-19
C4696 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT divide_by_2_1.tg_magic_3.OUT 0.175616f
C4697 7b_counter_0.MDFF_7.tspc2_magic_0.D CLK 1.54e-19
C4698 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A 0.001571f
C4699 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT P2 6.97e-20
C4700 p3_gen_magic_0.xnor_magic_4.OUT D2_5 0.139977f
C4701 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT a_1559_n5540# 1.54e-20
C4702 a_1541_n3597# D2_4 5.31e-19
C4703 p2_gen_magic_0.xnor_magic_6.OUT Q1 0.123243f
C4704 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 1.89e-19
C4705 DFF_magic_0.tg_magic_1.IN DFF_magic_0.tg_magic_2.IN 6.95e-19
C4706 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q1 0.009922f
C4707 OR_magic_2.A p3_gen_magic_0.P3 0.218409f
C4708 7b_counter_0.MDFF_7.tspc2_magic_0.Q Q4 0.208805f
C4709 mux_magic_0.OR_magic_0.A a_34156_n2297# 0.036613f
C4710 p3_gen_magic_0.3_inp_AND_magic_0.C a_13353_n6613# 0.536475f
C4711 a_8643_n1526# a_9059_n1973# 0.011514f
C4712 a_1957_n7648# Q7 2.48e-20
C4713 a_1209_6275# LD 0.002086f
C4714 a_26038_684# DFF_magic_0.tg_magic_3.OUT 8.55e-20
C4715 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A Q2 6.29e-19
C4716 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_1.tspc2_magic_0.CLK 0.003149f
C4717 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n8579# 0.093592f
C4718 7b_counter_0.MDFF_4.LD a_11279_3480# 0.001152f
C4719 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A Q5 5.18e-19
C4720 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 0.001207f
C4721 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A 7b_counter_0.MDFF_5.LD 0.43461f
C4722 p3_gen_magic_0.xnor_magic_3.OUT a_12174_n7648# 4.14e-19
C4723 a_21381_3524# Q7 0.001053f
C4724 p3_gen_magic_0.xnor_magic_4.OUT a_8643_n5540# 0.387036f
C4725 a_23207_5885# Q2 0.286536f
C4726 OR_magic_2.A DFF_magic_0.tg_magic_1.IN 0.001036f
C4727 a_19307_1669# D2_4 6.76e-19
C4728 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A 0.443527f
C4729 a_12387_3319# CLK 0.279959f
C4730 a_11279_6341# a_11191_5901# 0.477407f
C4731 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A 0.001081f
C4732 a_5185_2253# 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A 0.001985f
C4733 7b_counter_0.MDFF_4.LD a_15865_3363# 0.224216f
C4734 a_23560_3728# CLK 0.001962f
C4735 7b_counter_0.MDFF_4.LD OR_magic_2.A 1.03891f
C4736 a_13769_n2115# VDD 0.017033f
C4737 a_1541_n3597# Q2 0.001394f
C4738 a_2749_10148# 7b_counter_0.MDFF_3.tspc2_magic_0.CLK 0.00215f
C4739 a_5036_n7648# D2_3 1.85e-19
C4740 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A D2_2 0.014827f
C4741 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_8955_4557# 0.037614f
C4742 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B Q3 2.49e-19
C4743 a_1209_9773# 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 0.149276f
C4744 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n6471# 0.107012f
C4745 a_19152_6440# a_20171_6886# 0.043767f
C4746 a_12931_7470# D2_2 0.17383f
C4747 a_15865_4557# Q2 0.250956f
C4748 a_1409_7469# Q6 0.002005f
C4749 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.08926f
C4750 a_11292_n2115# a_13353_n2115# 6.73e-20
C4751 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A a_8955_3363# 1.77e-19
C4752 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n3597# 0.063777f
C4753 7b_counter_0.MDFF_5.LD a_12387_6986# 0.224216f
C4754 a_11292_n2115# D2_3 1.57e-19
C4755 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B Q1 0.00937f
C4756 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 0.169401f
C4757 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT Q3 0.024716f
C4758 a_26126_1124# DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 5.8e-22
C4759 p3_gen_magic_0.xnor_magic_4.OUT D2_7 0.008943f
C4760 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q6 0.004108f
C4761 a_19841_9774# a_21381_8741# 7.54e-20
C4762 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_1.OUT 1.46e-19
C4763 divide_by_2_0.tg_magic_3.OUT VDD 1.16334f
C4764 a_23985_7877# a_24185_7877# 0.522094f
C4765 a_15865_7470# a_17405_5901# 7.51e-20
C4766 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A a_12931_4557# 9.27e-19
C4767 p3_gen_magic_0.3_inp_AND_magic_0.C a_13769_n6613# 0.056504f
C4768 a_1409_2253# VDD 0.012214f
C4769 a_16065_1059# VDD 0.061661f
C4770 divide_by_2_1.tg_magic_1.IN mux_magic_0.IN1 0.004493f
C4771 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT Q3 7.89e-19
C4772 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT D2_4 0.0036f
C4773 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VDD 1.37922f
C4774 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT p3_gen_magic_0.P3 0.337254f
C4775 a_1559_n1973# a_1541_n3150# 0.190683f
C4776 a_4235_3947# Q6 0.012671f
C4777 divide_by_2_0.tg_magic_3.OUT D2_1 0.029655f
C4778 a_18891_6886# a_20041_4557# 7.7e-19
C4779 a_17405_5901# D2_3 0.016406f
C4780 a_22991_5885# Q5 2.42e-20
C4781 p2_gen_magic_0.xnor_magic_1.OUT a_5036_n4081# 2.1e-19
C4782 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A D2_1 3.54e-19
C4783 a_12387_9730# 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A 0.279825f
C4784 7b_counter_0.3_inp_AND_magic_0.A VDD 0.437145f
C4785 a_19152_1223# a_19152_739# 0.014143f
C4786 a_5515_3947# D2_5 4.45e-19
C4787 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VDD 1.0858f
C4788 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT a_8523_n3150# 0.107246f
C4789 7b_counter_0.MDFF_4.tspc2_magic_0.CLK D2_6 0.261939f
C4790 a_11279_1124# D2_6 0.042524f
C4791 a_26126_1124# 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A 0.036613f
C4792 a_8643_n6471# VDD 0.001396f
C4793 p2_gen_magic_0.3_inp_AND_magic_0.A Q4 0.040595f
C4794 a_1409_7469# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 1.77e-19
C4795 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19841_8580# 0.029386f
C4796 p3_gen_magic_0.xnor_magic_1.OUT a_8939_n7648# 6.88e-19
C4797 p3_gen_magic_0.xnor_magic_5.OUT a_5452_n7648# 0.06406f
C4798 a_4496_10093# a_4235_9163# 0.655098f
C4799 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_5 0.048608f
C4800 a_1409_2253# LD 0.037687f
C4801 a_2749_8740# a_2749_7308# 0.00112f
C4802 p3_gen_magic_0.xnor_magic_3.OUT p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 5.72e-19
C4803 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A LD 6.12e-19
C4804 a_5185_7469# CLK 2.95e-19
C4805 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.10998f
C4806 a_5385_2253# Q7 0.004613f
C4807 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A a_26038_4932# 3.58e-20
C4808 a_2749_4932# a_1209_3363# 7.51e-20
C4809 a_8411_3319# D2_6 0.290761f
C4810 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT 0.00167f
C4811 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.001697f
C4812 a_32816_n1264# mux_magic_0.IN2 0.003964f
C4813 a_12590_n7648# Q4 0.001058f
C4814 7b_counter_0.MDFF_5.LD a_17405_8741# 0.013942f
C4815 7b_counter_0.3_inp_AND_magic_0.A LD 0.004366f
C4816 a_5036_n3597# D2_3 4.88e-20
C4817 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT D2_1 0.015199f
C4818 7b_counter_0.MDFF_4.tspc2_magic_0.D a_9212_739# 0.282223f
C4819 a_8523_n3150# Q1 0.062238f
C4820 a_8643_n1526# a_8643_n1973# 0.013685f
C4821 mux_magic_0.OR_magic_0.A a_34156_n889# 0.414018f
C4822 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A Q5 0.00211f
C4823 7b_counter_0.MDFF_5.LD 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A 0.00221f
C4824 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.AND2_magic_1.A 3.88e-19
C4825 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B D2_3 4.21e-19
C4826 a_12931_7470# CLK 0.010628f
C4827 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 4e-20
C4828 7b_counter_0.MDFF_4.LD a_11191_4932# 0.002672f
C4829 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT Q3 0.024911f
C4830 VDD D2_6 6.1513f
C4831 a_11292_n6613# p3_gen_magic_0.xnor_magic_6.OUT 0.022681f
C4832 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A a_7303_8697# 2.4e-20
C4833 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_6.OUT 0.25446f
C4834 a_17405_684# D2_4 0.01674f
C4835 a_22991_5885# Q2 0.191655f
C4836 a_1209_2253# a_2749_684# 7.51e-20
C4837 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12387_8536# 0.001158f
C4838 a_30365_3514# CLK 0.016585f
C4839 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A Q5 0.004609f
C4840 D2_1 D2_6 0.257184f
C4841 7b_counter_0.MDFF_4.LD a_12387_3319# 0.224216f
C4842 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT Q1 0.01733f
C4843 7b_counter_0.MDFF_5.LD a_19152_6440# 0.006914f
C4844 a_1409_3363# CLK 7.14e-19
C4845 a_13553_n2115# VDD 0.016819f
C4846 7b_counter_0.MDFF_4.LD a_23560_3728# 0.006914f
C4847 a_9212_739# a_9689_1669# 0.16113f
C4848 7b_counter_0.MDFF_4.tspc2_magic_0.CLK D2_2 0.222046f
C4849 a_11279_1124# D2_2 0.044038f
C4850 7b_counter_0.DFF_magic_0.tg_magic_2.IN P2 2.11e-19
C4851 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT D2_7 0.059068f
C4852 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B D2_4 0.031239f
C4853 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A D2_4 0.02022f
C4854 DFF_magic_0.D a_23985_7877# 1.56e-20
C4855 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A a_15865_3363# 0.001985f
C4856 a_11191_5901# a_12387_5792# 0.002003f
C4857 a_19152_6440# a_19307_6886# 0.240883f
C4858 a_18891_6886# a_20171_6886# 0.007202f
C4859 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A a_7215_4932# 3.58e-20
C4860 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B Q1 0.009355f
C4861 a_1209_7469# Q6 0.001165f
C4862 7b_counter_0.MDFF_1.tspc2_magic_0.D Q4 7.41e-19
C4863 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A 0.001081f
C4864 p2_gen_magic_0.3_inp_AND_magic_0.A p2_gen_magic_0.xnor_magic_6.OUT 0.039667f
C4865 p3_gen_magic_0.xnor_magic_6.OUT a_14556_n8142# 0.249104f
C4866 LD D2_6 0.016864f
C4867 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT 0.001837f
C4868 a_15865_2253# Q1 0.015574f
C4869 divide_by_2_0.tg_magic_3.IN divide_by_2_0.tg_magic_1.IN 1.17013f
C4870 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 0.001081f
C4871 7b_counter_0.3_inp_AND_magic_0.A Q3 0.011276f
C4872 a_1409_9773# D2_7 0.009997f
C4873 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A Q1 0.002249f
C4874 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT 0.00105f
C4875 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN a_16186_n8142# 1.97e-20
C4876 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A Q6 0.108985f
C4877 p3_gen_magic_0.3_inp_AND_magic_0.C a_13553_n6613# 0.001361f
C4878 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A Q2 7.57e-19
C4879 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A 7b_counter_0.MDFF_6.tspc2_magic_0.CLK 8.78e-21
C4880 a_27234_1769# CLK 0.290487f
C4881 a_1209_2253# VDD 0.807784f
C4882 a_15865_1059# VDD 0.928771f
C4883 7b_counter_0.MDFF_5.tspc2_magic_0.CLK Q6 1.99e-20
C4884 7b_counter_0.MDFF_5.tspc2_magic_0.D a_9689_6886# 0.004574f
C4885 a_11279_8697# VDD 0.941683f
C4886 a_11292_n6613# D2_3 0.015364f
C4887 a_4496_4877# Q6 0.01249f
C4888 a_15865_8580# a_16065_8580# 0.299584f
C4889 p2_gen_magic_0.xnor_magic_3.OUT a_1975_n1973# 0.06406f
C4890 VDD D2_2 4.19298f
C4891 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B Q2 0.001065f
C4892 p2_gen_magic_0.xnor_magic_1.OUT a_1541_n4081# 0.334897f
C4893 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VDD 1.08725f
C4894 7b_counter_0.DFF_magic_0.tg_magic_2.IN VDD 1.0449f
C4895 7b_counter_0.MDFF_5.tspc2_magic_0.Q VDD 1.21217f
C4896 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT Q6 0.021234f
C4897 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A Q7 0.007832f
C4898 D2_2 D2_1 0.117187f
C4899 a_18891_1669# a_19152_739# 0.655098f
C4900 a_4651_3947# D2_5 0.0074f
C4901 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A Q2 8.26e-19
C4902 a_17405_7309# a_19307_6886# 2.34e-20
C4903 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 0.168057f
C4904 a_8939_n3150# Q5 3.02e-20
C4905 7b_counter_0.MDFF_5.tspc2_magic_0.Q D2_1 3.14e-19
C4906 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN 6.95e-19
C4907 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT a_1541_n3150# 9.19e-19
C4908 a_1209_7469# 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A 0.001985f
C4909 p2_gen_magic_0.xnor_magic_1.OUT VDD 6.76041f
C4910 a_5036_n7648# a_5452_n7648# 0.002223f
C4911 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT a_5036_n8095# 0.083665f
C4912 mux_magic_0.IN2 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT 7.64e-20
C4913 a_1209_2253# LD 0.224216f
C4914 a_8825_6886# a_9689_6886# 0.009722f
C4915 p2_gen_magic_0.xnor_magic_3.OUT Q6 0.045457f
C4916 Q3 D2_6 0.279943f
C4917 p3_gen_magic_0.xnor_magic_0.OUT p3_gen_magic_0.xnor_magic_3.OUT 0.041842f
C4918 mux_magic_0.IN2 a_32816_n2458# 0.128771f
C4919 p2_gen_magic_0.xnor_magic_1.OUT D2_1 0.534259f
C4920 LD D2_2 0.015283f
C4921 7b_counter_0.MDFF_6.tspc2_magic_0.Q a_19841_9774# 0.243646f
C4922 a_2749_2092# Q7 0.014002f
C4923 a_27234_4513# a_26038_4932# 0.002003f
C4924 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VDD 1.16929f
C4925 a_8411_8536# Q2 0.002692f
C4926 p2_gen_magic_0.xnor_magic_1.OUT p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 2.56e-19
C4927 7b_counter_0.MDFF_5.tspc2_magic_0.Q LD 5.47e-19
C4928 p3_gen_magic_0.3_inp_AND_magic_0.A Q4 0.01148f
C4929 7b_counter_0.MDFF_5.LD a_12931_9774# 0.004065f
C4930 a_16386_n3644# D2_6 7.6e-19
C4931 CLK P2 0.153023f
C4932 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT D2_1 0.059121f
C4933 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT a_8523_n3597# 1.63e-19
C4934 7b_counter_0.MDFF_3.QB a_1409_8579# 0.0013f
C4935 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B 0.005062f
C4936 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A 1.1e-20
C4937 DFF_magic_0.D 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT 0.025839f
C4938 7b_counter_0.MDFF_7.tspc2_magic_0.Q a_23258_575# 0.243646f
C4939 p2_gen_magic_0.3_inp_AND_magic_0.B VDD 0.747882f
C4940 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A a_12931_8580# 0.001034f
C4941 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q5 0.002165f
C4942 a_12931_4557# Q5 0.12882f
C4943 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN a_16186_n3644# 2.1e-20
C4944 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT 5.04e-22
C4945 7b_counter_0.MDFF_4.tspc2_magic_0.D Q4 0.001445f
C4946 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT a_8523_n7648# 0.011524f
C4947 7b_counter_0.MDFF_3.tspc2_magic_0.D D2_7 0.003663f
C4948 a_2749_5900# a_1209_6275# 0.002003f
C4949 a_12387_9730# a_12387_8536# 0.005574f
C4950 a_30365_4922# CLK 0.012979f
C4951 7b_counter_0.MDFF_4.LD a_30365_3514# 4.86e-20
C4952 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_12931_1059# 9.27e-19
C4953 a_4496_4393# a_5185_2253# 3.03e-19
C4954 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A a_27234_575# 0.279825f
C4955 a_9212_739# a_8825_1669# 0.007202f
C4956 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A a_6725_684# 3.58e-20
C4957 a_11708_n2115# VDD 0.012593f
C4958 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B 0.00112f
C4959 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A 0.00112f
C4960 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT a_5054_n1526# 0.063645f
C4961 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT D2_6 6.49e-19
C4962 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A D2_5 0.013552f
C4963 a_15865_1059# Q3 1.75e-19
C4964 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B VDD 1.21131f
C4965 a_18891_6886# a_19307_6886# 0.16113f
C4966 D2_2 Q3 0.108995f
C4967 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_4 0.00127f
C4968 a_16065_2253# Q1 0.004958f
C4969 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT a_8643_n1042# 0.090721f
C4970 p2_gen_magic_0.xnor_magic_5.OUT D2_6 6.3e-19
C4971 mux_magic_0.OR_magic_0.A mux_magic_0.OR_magic_0.B 0.178114f
C4972 p3_gen_magic_0.xnor_magic_6.OUT a_12174_n8095# 0.02352f
C4973 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B a_1209_8579# 0.146237f
C4974 VDD CLK 39.2676f
C4975 divide_by_2_1.tg_magic_1.IN VDD 1.85679f
C4976 a_12387_1769# Q1 0.015613f
C4977 a_22150_1124# 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A 2.4e-20
C4978 a_19841_8580# Q6 1.22e-19
C4979 CLK D2_1 1.82303f
C4980 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_5.OUT 0.173858f
C4981 a_8713_6842# D2_6 0.051141f
C4982 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4235_9163# 0.282223f
C4983 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B Q1 0.003442f
C4984 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A D2_6 2.27e-19
C4985 p2_gen_magic_0.xnor_magic_1.OUT Q3 0.001466f
C4986 a_1209_9773# Q2 6.79e-19
C4987 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A a_16065_9774# 0.037614f
C4988 a_23802_2253# CLK 0.067361f
C4989 7b_counter_0.MDFF_4.LD a_27234_1769# 0.224216f
C4990 7b_counter_0.MDFF_0.tspc2_magic_0.Q VDD 1.32846f
C4991 a_22062_684# VDD 1.60068f
C4992 divide_by_2_1.tg_magic_3.IN mux_magic_0.IN1 0.345958f
C4993 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A a_19841_3363# 0.001985f
C4994 7b_counter_0.MDFF_5.tspc2_magic_0.D a_8825_6886# 2.1e-20
C4995 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B LD 0.004701f
C4996 a_11191_10149# VDD 1.55695f
C4997 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B Q6 3.81e-19
C4998 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2 0.54616f
C4999 a_1559_n1526# a_1541_n3150# 0.001207f
C5000 a_1409_4557# Q6 0.003986f
C5001 p2_gen_magic_0.xnor_magic_3.OUT a_1559_n1973# 0.09365f
C5002 7b_counter_0.MDFF_3.QB 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A 0.004842f
C5003 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A CLK 0.003148f
C5004 7b_counter_0.DFF_magic_0.tg_magic_3.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.IN 0.859117f
C5005 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B Q7 0.031064f
C5006 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT p3_gen_magic_0.xnor_magic_4.OUT 1.11e-21
C5007 p2_gen_magic_0.xnor_magic_1.OUT a_16386_n3644# 0.140317f
C5008 a_8411_9730# VDD 0.917295f
C5009 LD CLK 0.666866f
C5010 p3_gen_magic_0.xnor_magic_1.OUT Q6 4.67e-19
C5011 a_1209_4557# Q7 9.91e-19
C5012 a_5185_2253# a_6725_684# 7.51e-20
C5013 7b_counter_0.MDFF_1.tspc2_magic_0.Q D2_3 0.28429f
C5014 a_12387_9730# Q2 6.82e-19
C5015 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT 0.16497f
C5016 a_17405_7309# a_17405_5901# 0.479729f
C5017 7b_counter_0.NAND_magic_0.A VDD 6.60135f
C5018 a_11292_n6613# a_13353_n6613# 6.73e-20
C5019 a_8411_9730# D2_1 2.73e-19
C5020 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 0.178114f
C5021 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B a_21381_8741# 0.428973f
C5022 a_1541_n3150# VDD 0.015101f
C5023 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A D2_7 0.091903f
C5024 Q4 D2_5 0.298048f
C5025 p2_gen_magic_0.3_inp_AND_magic_0.B Q3 0.002386f
C5026 7b_counter_0.MDFF_0.tspc2_magic_0.Q LD 0.121479f
C5027 a_8523_n8579# D2_6 0.017097f
C5028 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B a_5185_6275# 1.93e-19
C5029 7b_counter_0.MDFF_4.tspc2_magic_0.Q D2_6 0.410187f
C5030 a_1541_n3150# D2_1 0.057301f
C5031 p2_gen_magic_0.xnor_magic_5.OUT D2_2 0.065257f
C5032 7b_counter_0.3_inp_AND_magic_0.A 7b_counter_0.3_inp_AND_magic_0.B 0.247423f
C5033 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT 0.019115f
C5034 DFF_magic_0.tg_magic_1.IN P2 0.001931f
C5035 7b_counter_0.3_inp_AND_magic_0.C Q1 0.048749f
C5036 a_8411_9730# LD 4.93e-19
C5037 p2_gen_magic_0.3_inp_AND_magic_0.B a_16386_n3644# 6.81e-19
C5038 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A 0.003249f
C5039 a_8713_6842# D2_2 1.65e-19
C5040 7b_counter_0.MDFF_4.LD P2 0.001814f
C5041 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A D2_2 0.040266f
C5042 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT Q4 0.013327f
C5043 p3_gen_magic_0.xnor_magic_3.OUT Q6 0.038867f
C5044 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_4.tspc2_magic_0.CLK 0.084688f
C5045 7b_counter_0.NAND_magic_0.A LD 0.405505f
C5046 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B CLK 0.007602f
C5047 7b_counter_0.MDFF_5.tspc2_magic_0.Q a_8713_6842# 0.012895f
C5048 Q5 D2_4 0.586581f
C5049 7b_counter_0.MDFF_1.tspc2_magic_0.Q 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B 1.17e-20
C5050 p2_gen_magic_0.xnor_magic_1.OUT p2_gen_magic_0.xnor_magic_5.OUT 1.32582f
C5051 p2_gen_magic_0.xnor_magic_0.OUT a_12174_n3150# 0.001986f
C5052 7b_counter_0.MDFF_3.tspc2_magic_0.CLK Q7 0.020773f
C5053 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT a_1957_n3150# 0.005701f
C5054 CLK Q3 0.8319f
C5055 Q1 Q7 0.167752f
C5056 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_4.tspc2_magic_0.D 0.001711f
C5057 a_2749_8740# D2_7 0.04221f
C5058 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT Q6 0.007876f
C5059 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A a_15865_4557# 0.279825f
C5060 p3_gen_magic_0.P3 VDD 2.65516f
C5061 7b_counter_0.MDFF_4.LD a_30365_4922# 0.02544f
C5062 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A a_12387_575# 0.149276f
C5063 7b_counter_0.MDFF_4.LD a_8411_3319# 0.224142f
C5064 a_26126_3480# CLK 9.95e-19
C5065 a_11492_n2115# VDD 0.014256f
C5066 a_23560_3728# a_23258_1769# 3.03e-19
C5067 a_16386_n3644# CLK 2.19e-20
C5068 p2_gen_magic_0.AND2_magic_1.A a_12174_n4081# 0.616639f
C5069 p3_gen_magic_0.3_inp_AND_magic_0.B VDD 0.772318f
C5070 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B 7b_counter_0.MDFF_1.tspc2_magic_0.D 0.001711f
C5071 7b_counter_0.DFF_magic_0.tg_magic_2.OUT 7b_counter_0.DFF_magic_0.tg_magic_0.IN 0.010522f
C5072 a_22062_684# Q3 0.001205f
C5073 7b_counter_0.MDFF_0.tspc2_magic_0.Q Q3 2.63e-19
C5074 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q5 3.37e-19
C5075 p3_gen_magic_0.P3 D2_1 0.139604f
C5076 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p3_gen_magic_0.xnor_magic_3.OUT 3.07e-20
C5077 D2_7 Q4 0.319779f
C5078 a_1409_7469# VDD 0.012214f
C5079 Q2 Q5 0.609214f
C5080 7b_counter_0.MDFF_0.tspc2_magic_0.D Q6 0.017745f
C5081 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B Q7 0.013153f
C5082 DFF_magic_0.tg_magic_1.IN VDD 1.8556f
C5083 a_15865_2253# 7b_counter_0.MDFF_1.tspc2_magic_0.D 7.57e-20
C5084 a_1559_n1042# D2_4 0.008749f
C5085 a_12931_2253# Q1 0.004958f
C5086 p3_gen_magic_0.3_inp_AND_magic_0.B D2_1 0.002417f
C5087 7b_counter_0.MDFF_4.tspc2_magic_0.Q D2_2 5.09e-20
C5088 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B 0.00112f
C5089 p2_gen_magic_0.3_inp_AND_magic_0.B p2_gen_magic_0.xnor_magic_5.OUT 0.048563f
C5090 p3_gen_magic_0.xnor_magic_6.OUT a_8523_n8095# 0.371622f
C5091 p2_gen_magic_0.xnor_magic_6.OUT D2_5 0.06837f
C5092 7b_counter_0.MDFF_4.LD VDD 32.017803f
C5093 divide_by_2_1.tg_magic_1.IN divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT 0.003202f
C5094 7b_counter_0.MDFF_3.tspc2_magic_0.CLK a_4496_9609# 0.515297f
C5095 7b_counter_0.MDFF_1.tspc2_magic_0.CLK Q4 8.64e-19
C5096 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT CLK 1.32506f
C5097 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VDD 1.06707f
C5098 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A p2_gen_magic_0.xnor_magic_3.OUT 0.001039f
C5099 p2_gen_magic_0.xnor_magic_4.OUT Q4 0.010566f
C5100 a_5036_n4081# p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT 1.57e-20
C5101 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT a_5036_n7648# 0.107246f
C5102 7b_counter_0.MDFF_3.tspc2_magic_0.D a_4496_10093# 0.120019f
C5103 a_2749_8740# a_4235_9163# 0.002118f
C5104 a_1541_n3150# Q3 0.002098f
C5105 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B CLK 0.03641f
C5106 a_11279_6341# D2_6 0.022879f
C5107 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT D2_4 0.759724f
C5108 a_4496_4393# Q6 0.037884f
C5109 a_19152_1223# CLK 0.008343f
C5110 Q2 D2_4 0.616499f
C5111 7b_counter_0.MDFF_4.LD a_23802_2253# 0.036926f
C5112 a_12931_1059# VDD 0.056754f
C5113 a_19841_9774# Q6 3.72e-19
C5114 a_4235_3947# VDD 1.06723f
C5115 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT a_5470_n1973# 0.005701f
C5116 a_1409_7469# LD 0.037687f
C5117 a_1541_n8095# Q5 7.64e-19
C5118 a_7215_4932# Q6 0.002831f
C5119 a_12387_8536# a_12931_8580# 0.299584f
C5120 a_1559_n1042# Q2 2.48e-19
C5121 p2_gen_magic_0.xnor_magic_3.OUT a_5054_n1526# 1.65e-19
C5122 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A Q6 0.007545f
C5123 7b_counter_0.MDFF_3.QB a_1209_9773# 0.252332f
C5124 p3_gen_magic_0.xnor_magic_3.OUT a_1975_n6471# 0.06406f
C5125 p2_gen_magic_0.xnor_magic_1.OUT a_14756_n3644# 0.002538f
C5126 p2_gen_magic_0.xnor_magic_5.OUT CLK 0.002963f
C5127 a_5385_7469# Q7 0.014625f
C5128 a_1541_n7648# Q6 0.001276f
C5129 a_24003_10051# D2_4 0.003424f
C5130 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT p2_gen_magic_0.AND2_magic_1.A 0.23537f
C5131 p2_gen_magic_0.xnor_magic_3.OUT p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT 0.18088f
C5132 a_1209_4557# 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B 1.93e-19
C5133 a_8713_6842# CLK 0.039062f
C5134 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT Q2 0.537996f
C5135 p2_gen_magic_0.xnor_magic_0.OUT p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT 5.4e-19
C5136 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A CLK 0.004865f
C5137 p2_gen_magic_0.3_inp_AND_magic_0.C a_13769_n2115# 0.056504f
C5138 a_1541_n8095# D2_4 5.31e-19
C5139 p3_gen_magic_0.xnor_magic_6.OUT Q1 1.36e-19
C5140 a_8411_4513# D2_6 0.018958f
C5141 p2_gen_magic_0.xnor_magic_6.OUT D2_7 0.001727f
C5142 DFF_magic_0.D OR_magic_2.A 0.39399f
C5143 a_24003_10051# Q2 9.92e-20
C5144 a_32816_n1264# a_32616_n2458# 0.003083f
C5145 7b_counter_0.3_inp_AND_magic_0.VOUT 7b_counter_0.3_inp_AND_magic_0.A 0.001186f
C5146 p2_gen_magic_0.3_inp_AND_magic_0.B a_14756_n3644# 0.002269f
C5147 a_1559_n1973# p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT 7.35e-19
C5148 a_11279_8697# a_11279_6341# 0.00112f
C5149 a_16186_n3644# D2_6 8.9e-19
C5150 a_4496_9609# a_5385_7469# 5.39e-19
C5151 a_11279_6341# D2_2 0.132802f
C5152 7b_counter_0.MDFF_4.LD a_17405_4932# 0.002672f
C5153 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VDD 1.07838f
C5154 7b_counter_0.MDFF_4.LD 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B 0.004701f
C5155 a_6725_684# Q6 0.019469f
C5156 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT D2_3 6.1e-19
C5157 DFF_magic_0.tg_magic_1.IN Q3 1.71e-20
C5158 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A a_21381_4932# 3.58e-20
C5159 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_6.OUT 0.030838f
C5160 p2_gen_magic_0.xnor_magic_0.OUT a_8939_n3150# 1.73e-19
C5161 p2_gen_magic_0.xnor_magic_4.OUT p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT 0.099076f
C5162 7b_counter_0.MDFF_4.LD Q3 0.946651f
C5163 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT 5.61e-19
C5164 a_12931_6276# D2_2 0.00289f
C5165 OUT1 VSS 12.9387f
C5166 D2_4 VSS 15.452547f
C5167 D2_3 VSS 13.985817f
C5168 P2 VSS 8.035014f
C5169 D2_6 VSS 15.855757f
C5170 D2_5 VSS 16.776674f
C5171 Q5 VSS 30.518574f
C5172 Q4 VSS 22.805614f
C5173 Q6 VSS 21.969923f
C5174 Q7 VSS 17.87573f
C5175 Q3 VSS 15.270864f
C5176 D2_1 VSS 31.807589f
C5177 D2_2 VSS 13.32588f
C5178 D2_7 VSS 16.47188f
C5179 Q2 VSS 23.635399f
C5180 CLK VSS 62.804924f
C5181 Q1 VSS 20.457476f
C5182 LD VSS 35.866623f
C5183 VDD VSS 0.828663p
C5184 a_12174_n8579# VSS 0.031036f
C5185 a_8523_n8579# VSS 0.025369f
C5186 a_5036_n8579# VSS 0.042952f
C5187 a_1541_n8579# VSS 0.126953f
C5188 a_16386_n8142# VSS 0.27233f
C5189 a_14756_n8142# VSS 0.257354f
C5190 a_16186_n8142# VSS 0.726698f
C5191 a_14556_n8142# VSS 0.755892f
C5192 a_12174_n8095# VSS 0.089261f
C5193 a_8523_n8095# VSS 0.093912f
C5194 a_5036_n8095# VSS 0.088168f
C5195 a_12590_n7648# VSS 0.097856f
C5196 p3_gen_magic_0.AND2_magic_1.A VSS 1.66309f
C5197 a_1541_n8095# VSS 0.176904f
C5198 a_12174_n7648# VSS 2.58145f
C5199 a_8939_n7648# VSS 0.097615f
C5200 p3_gen_magic_0.xnor_magic_6.OUT VSS 3.62995f
C5201 a_8523_n7648# VSS 1.71307f
C5202 a_5452_n7648# VSS 0.096699f
C5203 p3_gen_magic_0.xnor_magic_5.OUT VSS 4.78274f
C5204 a_5036_n7648# VSS 1.66299f
C5205 a_1957_n7648# VSS 0.104141f
C5206 p3_gen_magic_0.xnor_magic_1.OUT VSS 5.620904f
C5207 a_1541_n7648# VSS 1.71115f
C5208 p3_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VSS 0.959872f
C5209 p3_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS 1.12616f
C5210 p3_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VSS 0.880706f
C5211 p3_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS 1.10575f
C5212 p3_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VSS 0.848569f
C5213 p3_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS 1.13643f
C5214 p3_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VSS 1.08838f
C5215 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS 1.19833f
C5216 divide_by_2_0.tg_magic_2.inverter_magic_0.VOUT VSS 0.312686f
C5217 divide_by_2_0.tg_magic_2.IN VSS 1.30934f
C5218 divide_by_2_0.tg_magic_0.inverter_magic_0.VOUT VSS 0.370986f
C5219 divide_by_2_0.tg_magic_0.IN VSS 1.47407f
C5220 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS 0.329237f
C5221 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.IN VSS 1.34024f
C5222 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS 0.320526f
C5223 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_0.IN VSS 1.42667f
C5224 a_13769_n6613# VSS 0.466221f
C5225 a_13553_n6613# VSS 0.095517f
C5226 a_11708_n6613# VSS 0.480536f
C5227 a_11492_n6613# VSS 0.124455f
C5228 a_9059_n6471# VSS 0.096699f
C5229 a_8643_n6471# VSS 1.68741f
C5230 divide_by_2_0.tg_magic_1.inverter_magic_0.VOUT VSS 0.313625f
C5231 divide_by_2_0.tg_magic_1.IN VSS 3.04057f
C5232 divide_by_2_0.tg_magic_3.IN VSS 5.47415f
C5233 a_23352_n6798# VSS 0.946088f
C5234 a_5470_n6471# VSS 0.096699f
C5235 a_5054_n6471# VSS 1.61057f
C5236 a_8643_n6024# VSS 0.072272f
C5237 a_1975_n6471# VSS 0.103867f
C5238 a_1559_n6471# VSS 1.7168f
C5239 a_5054_n6024# VSS 0.071896f
C5240 a_1559_n6024# VSS 0.177872f
C5241 a_23352_n5390# VSS 0.088525f
C5242 divide_by_2_0.tg_magic_3.OUT VSS 2.62756f
C5243 divide_by_2_0.tg_magic_3.inverter_magic_0.VOUT VSS 0.392517f
C5244 p3_gen_magic_0.P3 VSS 3.452314f
C5245 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_2.OUT VSS 2.98116f
C5246 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS 0.330515f
C5247 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN VSS 3.95458f
C5248 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK VSS 7.729736f
C5249 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.OUT VSS 2.4267f
C5250 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS 0.314806f
C5251 p3_gen_magic_0.3_inp_AND_magic_0.VOUT VSS 2.831018f
C5252 a_13353_n6613# VSS 1.59722f
C5253 p3_gen_magic_0.3_inp_AND_magic_0.C VSS 7.378616f
C5254 p3_gen_magic_0.3_inp_AND_magic_0.B VSS 3.24494f
C5255 p3_gen_magic_0.3_inp_AND_magic_0.A VSS 2.19654f
C5256 a_8643_n5540# VSS 0.025865f
C5257 p3_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS 1.14378f
C5258 p3_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VSS 0.79409f
C5259 a_5054_n5540# VSS 0.03217f
C5260 p3_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS 1.09952f
C5261 p3_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VSS 0.759084f
C5262 a_1559_n5540# VSS 0.093106f
C5263 p3_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS 1.17419f
C5264 p3_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VSS 1.10886f
C5265 a_11292_n6613# VSS 1.80611f
C5266 p3_gen_magic_0.xnor_magic_3.OUT VSS 3.242922f
C5267 p3_gen_magic_0.xnor_magic_4.OUT VSS 2.44693f
C5268 p3_gen_magic_0.xnor_magic_0.OUT VSS 2.85739f
C5269 a_12174_n4081# VSS 0.031036f
C5270 a_8523_n4081# VSS 0.025369f
C5271 a_5036_n4081# VSS 0.041332f
C5272 a_1541_n4081# VSS 0.119637f
C5273 a_16386_n3644# VSS 0.249081f
C5274 a_14756_n3644# VSS 0.251103f
C5275 a_16186_n3644# VSS 0.727616f
C5276 a_14556_n3644# VSS 0.749588f
C5277 a_12174_n3597# VSS 0.089261f
C5278 a_8523_n3597# VSS 0.093912f
C5279 a_5036_n3597# VSS 0.085235f
C5280 a_12590_n3150# VSS 0.097856f
C5281 p2_gen_magic_0.AND2_magic_1.A VSS 1.66564f
C5282 a_1541_n3597# VSS 0.180528f
C5283 a_12174_n3150# VSS 2.58371f
C5284 a_8939_n3150# VSS 0.097615f
C5285 p2_gen_magic_0.xnor_magic_6.OUT VSS 3.61325f
C5286 a_8523_n3150# VSS 1.6985f
C5287 a_5452_n3150# VSS 0.096699f
C5288 p2_gen_magic_0.xnor_magic_5.OUT VSS 2.54197f
C5289 a_5036_n3150# VSS 1.63197f
C5290 a_1957_n3150# VSS 0.104141f
C5291 p2_gen_magic_0.xnor_magic_1.OUT VSS 7.10976f
C5292 a_1541_n3150# VSS 1.90683f
C5293 p2_gen_magic_0.xnor_magic_2.inverter_magic_1.VOUT VSS 0.938049f
C5294 p2_gen_magic_0.xnor_magic_2.inverter_magic_0.VOUT VSS 1.12023f
C5295 p2_gen_magic_0.xnor_magic_6.inverter_magic_1.VOUT VSS 0.849532f
C5296 p2_gen_magic_0.xnor_magic_6.inverter_magic_0.VOUT VSS 1.0462f
C5297 p2_gen_magic_0.xnor_magic_5.inverter_magic_1.VOUT VSS 0.828209f
C5298 p2_gen_magic_0.xnor_magic_5.inverter_magic_0.VOUT VSS 1.05364f
C5299 p2_gen_magic_0.xnor_magic_1.inverter_magic_1.VOUT VSS 1.13095f
C5300 p2_gen_magic_0.xnor_magic_1.inverter_magic_0.VOUT VSS 1.10287f
C5301 a_32816_n2458# VSS 0.320067f
C5302 DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS 0.314579f
C5303 DFF_magic_0.tg_magic_2.IN VSS 1.29396f
C5304 a_32616_n2458# VSS 0.938649f
C5305 mux_magic_0.IN2 VSS 4.931779f
C5306 DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS 0.343218f
C5307 DFF_magic_0.tg_magic_0.IN VSS 1.45806f
C5308 p2_gen_magic_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS 0.326676f
C5309 p2_gen_magic_0.DFF_magic_0.tg_magic_2.IN VSS 1.34411f
C5310 p2_gen_magic_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS 0.315638f
C5311 p2_gen_magic_0.DFF_magic_0.tg_magic_0.IN VSS 1.40607f
C5312 a_13769_n2115# VSS 0.466221f
C5313 a_13553_n2115# VSS 0.095517f
C5314 a_11708_n2115# VSS 0.480536f
C5315 a_11492_n2115# VSS 0.129679f
C5316 a_9059_n1973# VSS 0.096699f
C5317 a_8643_n1973# VSS 1.68741f
C5318 a_32816_n1264# VSS 0.281839f
C5319 a_34156_n2297# VSS 0.970791f
C5320 a_34156_n889# VSS 0.096542f
C5321 mux_magic_0.OR_magic_0.B VSS 0.96309f
C5322 mux_magic_0.OR_magic_0.A VSS 0.707909f
C5323 a_5470_n1973# VSS 0.096699f
C5324 a_5054_n1973# VSS 1.62072f
C5325 a_8643_n1526# VSS 0.072272f
C5326 a_1975_n1973# VSS 0.103867f
C5327 a_1559_n1973# VSS 1.89248f
C5328 a_5054_n1526# VSS 0.071877f
C5329 a_1559_n1526# VSS 0.178355f
C5330 a_32616_n1264# VSS 0.749859f
C5331 mux_magic_0.AND2_magic_0.A VSS 1.44736f
C5332 DFF_magic_0.tg_magic_2.OUT VSS 2.57761f
C5333 DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS 0.311593f
C5334 DFF_magic_0.tg_magic_1.IN VSS 3.06532f
C5335 DFF_magic_0.tg_magic_3.OUT VSS 2.57648f
C5336 DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS 0.326997f
C5337 p2_gen_magic_0.DFF_magic_0.tg_magic_2.OUT VSS 2.71557f
C5338 p2_gen_magic_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS 0.327656f
C5339 p2_gen_magic_0.DFF_magic_0.tg_magic_1.IN VSS 3.16037f
C5340 p2_gen_magic_0.DFF_magic_0.tg_magic_3.OUT VSS 2.39596f
C5341 p2_gen_magic_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS 0.30842f
C5342 p2_gen_magic_0.3_inp_AND_magic_0.VOUT VSS 1.49282f
C5343 a_13353_n2115# VSS 1.59691f
C5344 p2_gen_magic_0.3_inp_AND_magic_0.C VSS 6.654581f
C5345 p2_gen_magic_0.3_inp_AND_magic_0.B VSS 3.27039f
C5346 p2_gen_magic_0.3_inp_AND_magic_0.A VSS 2.19848f
C5347 a_8643_n1042# VSS 0.025865f
C5348 p2_gen_magic_0.xnor_magic_0.inverter_magic_0.VOUT VSS 1.15899f
C5349 p2_gen_magic_0.xnor_magic_0.inverter_magic_1.VOUT VSS 0.861374f
C5350 a_5054_n1042# VSS 0.033257f
C5351 p2_gen_magic_0.xnor_magic_4.inverter_magic_0.VOUT VSS 1.1032f
C5352 p2_gen_magic_0.xnor_magic_4.inverter_magic_1.VOUT VSS 0.851994f
C5353 a_1559_n1042# VSS 0.093378f
C5354 p2_gen_magic_0.xnor_magic_3.inverter_magic_0.VOUT VSS 1.09687f
C5355 p2_gen_magic_0.xnor_magic_3.inverter_magic_1.VOUT VSS 1.13515f
C5356 a_11292_n2115# VSS 1.80832f
C5357 p2_gen_magic_0.xnor_magic_3.OUT VSS 3.233982f
C5358 p2_gen_magic_0.xnor_magic_4.OUT VSS 2.56475f
C5359 p2_gen_magic_0.xnor_magic_0.OUT VSS 2.81928f
C5360 divide_by_2_1.tg_magic_2.inverter_magic_0.VOUT VSS 0.315003f
C5361 divide_by_2_1.tg_magic_2.IN VSS 1.3901f
C5362 divide_by_2_1.tg_magic_0.inverter_magic_0.VOUT VSS 0.353019f
C5363 a_27778_1059# VSS 0.218238f
C5364 divide_by_2_1.tg_magic_0.IN VSS 1.47906f
C5365 a_27234_575# VSS 0.700586f
C5366 a_23802_1059# VSS 0.211935f
C5367 7b_counter_0.MDFF_7.mux_magic_3.AND2_magic_0.A VSS 1.44824f
C5368 a_23258_575# VSS 0.688677f
C5369 a_26038_684# VSS 0.146451f
C5370 7b_counter_0.MDFF_7.mux_magic_2.AND2_magic_0.A VSS 1.43048f
C5371 a_19152_739# VSS 0.107771f
C5372 a_16065_1059# VSS 0.212196f
C5373 a_15865_1059# VSS 0.685294f
C5374 a_22062_684# VSS 0.082089f
C5375 a_12931_1059# VSS 0.2134f
C5376 a_12387_575# VSS 0.698036f
C5377 a_27778_2253# VSS 0.244122f
C5378 a_20171_1669# VSS 0.245122f
C5379 a_19307_1669# VSS 0.28235f
C5380 a_17405_684# VSS 0.085437f
C5381 7b_counter_0.MDFF_1.mux_magic_0.AND2_magic_0.A VSS 1.4219f
C5382 7b_counter_0.MDFF_4.mux_magic_0.AND2_magic_0.A VSS 1.42475f
C5383 a_9412_739# VSS 0.068079f
C5384 a_5385_1059# VSS 0.212913f
C5385 a_5185_1059# VSS 0.687997f
C5386 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.A VSS 0.717439f
C5387 a_26126_1124# VSS 1.05041f
C5388 7b_counter_0.MDFF_7.mux_magic_3.OR_magic_0.B VSS 0.977969f
C5389 mux_magic_0.IN1 VSS 8.655424f
C5390 a_27234_1769# VSS 0.87119f
C5391 a_23802_2253# VSS 0.237594f
C5392 a_19152_1223# VSS 1.47203f
C5393 a_18891_1669# VSS 1.0351f
C5394 a_11191_684# VSS 0.121388f
C5395 a_1409_1059# VSS 0.303301f
C5396 a_1209_1059# VSS 0.744596f
C5397 7b_counter_0.MDFF_1.tspc2_magic_0.D VSS 0.999055f
C5398 a_9689_1669# VSS 0.229253f
C5399 a_8825_1669# VSS 0.239729f
C5400 a_6725_684# VSS 0.078522f
C5401 7b_counter_0.MDFF_0.mux_magic_2.AND2_magic_0.A VSS 1.43045f
C5402 a_9212_739# VSS 0.950743f
C5403 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.A VSS 0.67221f
C5404 a_22150_1124# VSS 0.901791f
C5405 a_17405_2092# VSS 0.885368f
C5406 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.A VSS 0.668821f
C5407 7b_counter_0.MDFF_7.mux_magic_2.OR_magic_0.B VSS 0.918414f
C5408 divide_by_2_1.tg_magic_1.inverter_magic_0.VOUT VSS 0.3143f
C5409 divide_by_2_1.tg_magic_1.IN VSS 3.05428f
C5410 divide_by_2_1.tg_magic_3.IN VSS 6.061936f
C5411 a_23258_1769# VSS 0.844476f
C5412 7b_counter_0.MDFF_1.mux_magic_0.OR_magic_0.B VSS 0.911745f
C5413 a_16065_2253# VSS 0.23428f
C5414 a_12931_2253# VSS 0.237417f
C5415 a_8713_1625# VSS 1.26866f
C5416 a_2749_684# VSS 0.089815f
C5417 7b_counter_0.MDFF_0.mux_magic_3.AND2_magic_0.A VSS 1.46929f
C5418 7b_counter_0.MDFF_4.tspc2_magic_0.D VSS 0.957574f
C5419 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.A VSS 0.6907f
C5420 a_11279_1124# VSS 1.00138f
C5421 a_6725_2092# VSS 0.865581f
C5422 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.A VSS 0.658099f
C5423 7b_counter_0.MDFF_4.mux_magic_0.OR_magic_0.B VSS 0.956551f
C5424 a_15865_2253# VSS 0.855646f
C5425 a_12387_1769# VSS 0.865053f
C5426 7b_counter_0.MDFF_0.mux_magic_2.OR_magic_0.B VSS 0.885889f
C5427 a_5385_2253# VSS 0.238539f
C5428 a_2749_2092# VSS 0.909652f
C5429 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.A VSS 0.689727f
C5430 a_5185_2253# VSS 0.844356f
C5431 7b_counter_0.MDFF_0.mux_magic_3.OR_magic_0.B VSS 0.923546f
C5432 a_1409_2253# VSS 0.322786f
C5433 a_1209_2253# VSS 0.910094f
C5434 divide_by_2_1.tg_magic_3.OUT VSS 2.67464f
C5435 divide_by_2_1.tg_magic_3.inverter_magic_0.VOUT VSS 0.346249f
C5436 a_27778_3363# VSS 0.240272f
C5437 a_20041_3363# VSS 0.244534f
C5438 a_27234_3319# VSS 0.868816f
C5439 a_24536_3947# VSS 0.228367f
C5440 a_23672_3947# VSS 0.246406f
C5441 a_16065_3363# VSS 0.239587f
C5442 a_12931_3363# VSS 0.231918f
C5443 OR_magic_1.VOUT VSS 10.425723f
C5444 a_8955_3363# VSS 0.237708f
C5445 a_19841_3363# VSS 0.862214f
C5446 a_27778_4557# VSS 0.213669f
C5447 a_15865_3363# VSS 0.856173f
C5448 a_12387_3319# VSS 0.851933f
C5449 a_30365_3514# VSS 0.872892f
C5450 a_30365_4922# VSS 0.106976f
C5451 OR_magic_2.A VSS 10.970915f
C5452 a_23560_3728# VSS 1.30739f
C5453 a_1409_3363# VSS 0.305818f
C5454 a_8411_3319# VSS 0.826954f
C5455 a_26126_3480# VSS 1.0149f
C5456 a_24259_4877# VSS 0.06541f
C5457 a_24059_4877# VSS 0.949152f
C5458 a_20041_4557# VSS 0.236673f
C5459 7b_counter_0.MDFF_7.tspc2_magic_0.Q VSS 2.30423f
C5460 a_26038_4932# VSS 0.146329f
C5461 7b_counter_0.MDFF_7.mux_magic_0.AND2_magic_0.A VSS 1.40864f
C5462 a_27234_4513# VSS 0.682316f
C5463 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.A VSS 0.716075f
C5464 7b_counter_0.MDFF_7.mux_magic_0.OR_magic_0.B VSS 0.981615f
C5465 7b_counter_0.MDFF_7.tspc2_magic_0.D VSS 0.973011f
C5466 7b_counter_0.MDFF_7.tspc2_magic_0.CLK VSS 4.455723f
C5467 a_21381_3524# VSS 0.912679f
C5468 7b_counter_0.MDFF_1.tspc2_magic_0.CLK VSS 3.70698f
C5469 a_16065_4557# VSS 0.211168f
C5470 a_5515_3947# VSS 0.24134f
C5471 a_4651_3947# VSS 0.228733f
C5472 a_21381_4932# VSS 0.082032f
C5473 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.B VSS 0.898486f
C5474 7b_counter_0.MDFF_1.mux_magic_2.OR_magic_0.A VSS 0.652921f
C5475 a_17405_3524# VSS 0.906287f
C5476 a_12931_4557# VSS 0.212372f
C5477 a_1209_3363# VSS 0.912889f
C5478 7b_counter_0.MDFF_4.tspc2_magic_0.CLK VSS 4.247447f
C5479 a_17405_4932# VSS 0.085596f
C5480 a_19841_4557# VSS 0.68426f
C5481 7b_counter_0.MDFF_1.tspc2_magic_0.Q VSS 2.50377f
C5482 7b_counter_0.MDFF_1.mux_magic_2.AND2_magic_0.A VSS 1.47367f
C5483 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.B VSS 0.891585f
C5484 7b_counter_0.MDFF_1.mux_magic_3.OR_magic_0.A VSS 0.649664f
C5485 a_8955_4557# VSS 0.209955f
C5486 a_4496_4393# VSS 1.24177f
C5487 a_15865_4557# VSS 0.6671f
C5488 7b_counter_0.MDFF_1.mux_magic_3.AND2_magic_0.A VSS 1.40253f
C5489 a_11279_3480# VSS 1.02124f
C5490 a_11191_4932# VSS 0.121155f
C5491 7b_counter_0.MDFF_4.mux_magic_3.AND2_magic_0.A VSS 1.40462f
C5492 a_12387_4513# VSS 0.677684f
C5493 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.A VSS 0.668515f
C5494 7b_counter_0.MDFF_4.mux_magic_3.OR_magic_0.B VSS 0.926418f
C5495 a_7303_3480# VSS 0.914251f
C5496 7b_counter_0.MDFF_0.tspc2_magic_0.Q VSS 2.73801f
C5497 a_4235_3947# VSS 0.945503f
C5498 a_4496_4877# VSS 0.063782f
C5499 a_1409_4557# VSS 0.285451f
C5500 a_7215_4932# VSS 0.082032f
C5501 7b_counter_0.MDFF_4.mux_magic_2.AND2_magic_0.A VSS 1.41018f
C5502 7b_counter_0.MDFF_4.tspc2_magic_0.Q VSS 2.46654f
C5503 a_8411_4513# VSS 0.669359f
C5504 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.A VSS 0.651956f
C5505 7b_counter_0.MDFF_4.mux_magic_2.OR_magic_0.B VSS 0.894665f
C5506 7b_counter_0.MDFF_0.tspc2_magic_0.CLK VSS 4.453256f
C5507 7b_counter_0.MDFF_0.tspc2_magic_0.D VSS 0.924942f
C5508 a_2749_3524# VSS 0.88582f
C5509 a_2749_4932# VSS 0.089655f
C5510 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.B VSS 0.897789f
C5511 7b_counter_0.MDFF_0.mux_magic_0.OR_magic_0.A VSS 0.668484f
C5512 a_1209_4557# VSS 0.724443f
C5513 7b_counter_0.MDFF_0.mux_magic_0.AND2_magic_0.A VSS 1.4422f
C5514 7b_counter_0.DFF_magic_0.tg_magic_2.inverter_magic_0.VOUT VSS 0.269665f
C5515 7b_counter_0.DFF_magic_0.tg_magic_2.IN VSS 1.30364f
C5516 7b_counter_0.DFF_magic_0.tg_magic_0.inverter_magic_0.VOUT VSS 0.288541f
C5517 7b_counter_0.DFF_magic_0.tg_magic_0.IN VSS 1.40659f
C5518 a_23793_5904# VSS 0.255995f
C5519 a_21504_5904# VSS 0.186261f
C5520 a_19152_5956# VSS 0.10352f
C5521 a_16065_6276# VSS 0.211168f
C5522 a_15865_6276# VSS 0.6671f
C5523 a_12931_6276# VSS 0.211158f
C5524 a_12387_5792# VSS 0.674647f
C5525 a_20171_6886# VSS 0.252268f
C5526 a_19307_6886# VSS 0.278098f
C5527 a_17405_5901# VSS 0.085437f
C5528 7b_counter_0.MDFF_6.mux_magic_0.AND2_magic_0.A VSS 1.40016f
C5529 7b_counter_0.MDFF_5.mux_magic_0.AND2_magic_0.A VSS 1.4012f
C5530 a_9412_5956# VSS 0.067196f
C5531 a_5385_6275# VSS 0.209955f
C5532 a_5185_6275# VSS 0.668863f
C5533 a_19152_6440# VSS 1.5264f
C5534 a_18891_6886# VSS 1.04734f
C5535 a_11191_5901# VSS 0.120465f
C5536 a_1409_6275# VSS 0.288456f
C5537 a_1209_6275# VSS 0.724848f
C5538 7b_counter_0.DFF_magic_0.tg_magic_2.OUT VSS 2.58537f
C5539 7b_counter_0.DFF_magic_0.tg_magic_1.inverter_magic_0.VOUT VSS 0.303145f
C5540 7b_counter_0.DFF_magic_0.tg_magic_1.IN VSS 3.01671f
C5541 7b_counter_0.DFF_magic_0.tg_magic_3.OUT VSS 2.41723f
C5542 7b_counter_0.DFF_magic_0.tg_magic_3.inverter_magic_0.VOUT VSS 0.323634f
C5543 7b_counter_0.MDFF_6.tspc2_magic_0.D VSS 0.957178f
C5544 a_9689_6886# VSS 0.21456f
C5545 a_8825_6886# VSS 0.239156f
C5546 a_6725_5900# VSS 0.082032f
C5547 7b_counter_0.MDFF_3.mux_magic_2.AND2_magic_0.A VSS 1.4047f
C5548 a_9212_5956# VSS 0.918368f
C5549 a_17405_7309# VSS 0.885641f
C5550 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.A VSS 0.648641f
C5551 7b_counter_0.MDFF_6.mux_magic_0.OR_magic_0.B VSS 0.888911f
C5552 a_16065_7470# VSS 0.240907f
C5553 a_12931_7470# VSS 0.23499f
C5554 a_8713_6842# VSS 1.25878f
C5555 a_2749_5900# VSS 0.089815f
C5556 7b_counter_0.MDFF_3.mux_magic_3.AND2_magic_0.A VSS 1.4436f
C5557 7b_counter_0.MDFF_5.tspc2_magic_0.D VSS 0.947881f
C5558 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.A VSS 0.663449f
C5559 a_11279_6341# VSS 0.985633f
C5560 a_6725_7308# VSS 0.831638f
C5561 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.A VSS 0.672171f
C5562 7b_counter_0.MDFF_5.mux_magic_0.OR_magic_0.B VSS 0.923408f
C5563 a_15865_7470# VSS 0.855646f
C5564 a_12387_6986# VSS 0.860111f
C5565 7b_counter_0.MDFF_3.mux_magic_2.OR_magic_0.B VSS 0.883952f
C5566 a_5385_7469# VSS 0.238539f
C5567 a_2749_7308# VSS 0.909652f
C5568 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.A VSS 0.669507f
C5569 a_5185_7469# VSS 0.844353f
C5570 7b_counter_0.MDFF_3.mux_magic_3.OR_magic_0.B VSS 0.900468f
C5571 a_1409_7469# VSS 0.327537f
C5572 a_1209_7469# VSS 0.913205f
C5573 a_24401_7877# VSS 0.469686f
C5574 a_24185_7877# VSS 0.09803f
C5575 a_23207_5885# VSS 0.138927f
C5576 a_22991_5885# VSS 0.136139f
C5577 a_20041_8580# VSS 0.242878f
C5578 a_16065_8580# VSS 0.230526f
C5579 a_12931_8580# VSS 0.246855f
C5580 a_23985_7877# VSS 1.63436f
C5581 7b_counter_0.3_inp_AND_magic_0.C VSS 2.6219f
C5582 7b_counter_0.3_inp_AND_magic_0.B VSS 1.80904f
C5583 7b_counter_0.3_inp_AND_magic_0.A VSS 4.59225f
C5584 7b_counter_0.MDFF_4.LD VSS 50.00047f
C5585 a_8955_8580# VSS 0.237472f
C5586 a_19841_8580# VSS 0.864205f
C5587 a_15865_8580# VSS 0.85571f
C5588 a_12387_8536# VSS 0.865603f
C5589 DFF_magic_0.D VSS 10.856565f
C5590 a_1409_8579# VSS 0.308296f
C5591 a_8411_8536# VSS 0.808374f
C5592 a_20041_9774# VSS 0.220277f
C5593 a_24003_10051# VSS 0.354039f
C5594 a_21381_8741# VSS 0.870004f
C5595 7b_counter_0.MDFF_6.tspc2_magic_0.CLK VSS 3.70461f
C5596 a_16065_9774# VSS 0.213112f
C5597 a_5515_9163# VSS 0.248184f
C5598 a_4651_9163# VSS 0.228733f
C5599 a_21381_10149# VSS 0.078522f
C5600 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.B VSS 0.90284f
C5601 7b_counter_0.MDFF_6.mux_magic_2.OR_magic_0.A VSS 0.663468f
C5602 a_17405_8741# VSS 0.905744f
C5603 a_12931_9774# VSS 0.21697f
C5604 a_1209_8579# VSS 0.868128f
C5605 7b_counter_0.MDFF_5.tspc2_magic_0.CLK VSS 4.287547f
C5606 a_17405_10149# VSS 0.085596f
C5607 a_19841_9774# VSS 0.70538f
C5608 7b_counter_0.MDFF_6.tspc2_magic_0.Q VSS 2.61695f
C5609 7b_counter_0.MDFF_6.mux_magic_2.AND2_magic_0.A VSS 1.51881f
C5610 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.B VSS 0.918307f
C5611 7b_counter_0.MDFF_6.mux_magic_3.OR_magic_0.A VSS 0.674063f
C5612 a_8955_9774# VSS 0.216178f
C5613 a_4496_9609# VSS 1.28266f
C5614 a_15865_9774# VSS 0.689983f
C5615 7b_counter_0.MDFF_6.mux_magic_3.AND2_magic_0.A VSS 1.42844f
C5616 a_11279_8697# VSS 1.03297f
C5617 a_11191_10149# VSS 0.12395f
C5618 7b_counter_0.MDFF_5.mux_magic_3.AND2_magic_0.A VSS 1.4321f
C5619 a_12387_9730# VSS 0.700567f
C5620 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.A VSS 0.697957f
C5621 7b_counter_0.MDFF_5.mux_magic_3.OR_magic_0.B VSS 0.966228f
C5622 7b_counter_0.MDFF_5.LD VSS 28.1624f
C5623 a_7303_8697# VSS 0.868545f
C5624 7b_counter_0.MDFF_3.tspc2_magic_0.Q VSS 2.55225f
C5625 a_4235_9163# VSS 0.945711f
C5626 a_4496_10093# VSS 0.063782f
C5627 a_1409_9773# VSS 0.319976f
C5628 a_7215_10149# VSS 0.082032f
C5629 7b_counter_0.MDFF_5.mux_magic_2.AND2_magic_0.A VSS 1.4334f
C5630 7b_counter_0.MDFF_5.tspc2_magic_0.Q VSS 2.44985f
C5631 a_8411_9730# VSS 0.690148f
C5632 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.A VSS 0.67325f
C5633 7b_counter_0.MDFF_5.mux_magic_2.OR_magic_0.B VSS 0.909109f
C5634 7b_counter_0.MDFF_3.tspc2_magic_0.CLK VSS 4.528266f
C5635 7b_counter_0.MDFF_3.tspc2_magic_0.D VSS 0.95917f
C5636 a_2749_8740# VSS 0.886179f
C5637 a_2749_10148# VSS 0.089922f
C5638 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.B VSS 0.925167f
C5639 7b_counter_0.MDFF_3.mux_magic_0.OR_magic_0.A VSS 0.693838f
C5640 a_1209_9773# VSS 0.752332f
C5641 7b_counter_0.MDFF_3.QB VSS 2.13753f
C5642 7b_counter_0.MDFF_3.mux_magic_0.AND2_magic_0.A VSS 1.47031f
C5643 7b_counter_0.NAND_magic_0.VOUT VSS 2.46686f
C5644 7b_counter_0.3_inp_AND_magic_0.VOUT VSS 2.74417f
C5645 7b_counter_0.NAND_magic_0.A VSS 11.185051f
C5646 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t0 VSS 0.034129f
C5647 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t2 VSS 0.039741f
C5648 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t1 VSS 0.031057f
C5649 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t10 VSS 0.110718f
C5650 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t5 VSS 0.056192f
C5651 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t8 VSS 0.037155f
C5652 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n0 VSS 0.09845f
C5653 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n1 VSS 0.140921f
C5654 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t3 VSS 0.070462f
C5655 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t9 VSS 0.0385f
C5656 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t12 VSS 0.030014f
C5657 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t4 VSS 0.060221f
C5658 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n2 VSS 0.06393f
C5659 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t11 VSS 0.076733f
C5660 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n3 VSS 0.093075f
C5661 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n4 VSS 0.252841f
C5662 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t6 VSS 0.030014f
C5663 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.t7 VSS 0.059765f
C5664 7b_counter_0.MDFF_5.tspc2_magic_0.CLK.n5 VSS 0.059173f
C5665 7b_counter_0.MDFF_5.QB.t1 VSS 0.115287f
C5666 7b_counter_0.MDFF_5.QB.t0 VSS 0.111865f
C5667 7b_counter_0.MDFF_5.mux_magic_0.IN1 VSS 1.10688f
C5668 7b_counter_0.MDFF_5.tspc2_magic_0.QB VSS 1.1185f
C5669 7b_counter_0.MDFF_5.QB.n0 VSS 0.195382f
C5670 7b_counter_0.MDFF_5.QB.t8 VSS 0.185836f
C5671 7b_counter_0.MDFF_5.QB.n1 VSS 0.146385f
C5672 7b_counter_0.MDFF_5.QB.t4 VSS 0.084564f
C5673 7b_counter_0.MDFF_5.QB.t7 VSS 0.101324f
C5674 7b_counter_0.MDFF_5.QB.n2 VSS 0.169388f
C5675 7b_counter_0.MDFF_5.QB.t3 VSS 0.062978f
C5676 7b_counter_0.MDFF_5.QB.t6 VSS 0.119652f
C5677 7b_counter_0.MDFF_5.QB.t2 VSS 0.079739f
C5678 7b_counter_0.MDFF_5.QB.n3 VSS 0.148949f
C5679 7b_counter_0.MDFF_5.QB.t5 VSS 0.150866f
C5680 7b_counter_0.MDFF_5.QB.n4 VSS 0.102403f
C5681 OR_magic_2.VOUT.n0 VSS 1.40514f
C5682 divide_by_2_0.inverter_magic_5.VIN VSS 0.694487f
C5683 OR_magic_2.VOUT.n1 VSS 0.347031f
C5684 divide_by_2_0.tg_magic_0.CLK VSS 0.934611f
C5685 OR_magic_2.VOUT.t4 VSS 0.057561f
C5686 OR_magic_2.VOUT.t24 VSS 0.11207f
C5687 OR_magic_2.VOUT.n2 VSS 0.087968f
C5688 OR_magic_2.VOUT.t25 VSS 0.11207f
C5689 OR_magic_2.VOUT.n3 VSS 0.087968f
C5690 OR_magic_2.VOUT.t15 VSS 0.089632f
C5691 OR_magic_2.VOUT.t21 VSS 0.12124f
C5692 OR_magic_2.VOUT.t9 VSS 0.13222f
C5693 OR_magic_2.VOUT.n4 VSS 0.121562f
C5694 OR_magic_2.VOUT.t26 VSS 0.118496f
C5695 OR_magic_2.VOUT.t16 VSS 0.118496f
C5696 OR_magic_2.VOUT.n5 VSS 0.144053f
C5697 OR_magic_2.VOUT.t6 VSS 0.313065f
C5698 OR_magic_2.VOUT.t19 VSS 0.057561f
C5699 OR_magic_2.VOUT.t13 VSS 0.11207f
C5700 OR_magic_2.VOUT.n6 VSS 0.087968f
C5701 OR_magic_2.VOUT.t18 VSS 0.11207f
C5702 OR_magic_2.VOUT.n7 VSS 0.087968f
C5703 OR_magic_2.VOUT.t7 VSS 0.089632f
C5704 OR_magic_2.VOUT.t10 VSS 0.12124f
C5705 OR_magic_2.VOUT.t22 VSS 0.13222f
C5706 OR_magic_2.VOUT.n8 VSS 0.121165f
C5707 OR_magic_2.VOUT.t14 VSS 0.118496f
C5708 OR_magic_2.VOUT.t8 VSS 0.118496f
C5709 OR_magic_2.VOUT.n9 VSS 0.144053f
C5710 OR_magic_2.VOUT.t20 VSS 0.176264f
C5711 OR_magic_2.VOUT.t3 VSS 0.12124f
C5712 OR_magic_2.VOUT.t17 VSS 0.13222f
C5713 OR_magic_2.VOUT.t5 VSS 0.11207f
C5714 OR_magic_2.VOUT.t23 VSS 0.057561f
C5715 OR_magic_2.VOUT.t12 VSS 0.11207f
C5716 OR_magic_2.VOUT.n10 VSS 0.087968f
C5717 OR_magic_2.VOUT.n11 VSS 0.087968f
C5718 OR_magic_2.VOUT.t11 VSS 0.089632f
C5719 OR_magic_2.VOUT.n12 VSS 0.121165f
C5720 OR_magic_2.VOUT.t2 VSS 0.076215f
C5721 OR_magic_2.VOUT.t0 VSS 0.059561f
C5722 OR_magic_2.VOUT.t1 VSS 0.065453f
C5723 7b_counter_0.MDFF_1.QB.t1 VSS 0.082913f
C5724 7b_counter_0.MDFF_1.QB.t0 VSS 0.080452f
C5725 7b_counter_0.MDFF_1.mux_magic_0.IN1 VSS 0.818433f
C5726 7b_counter_0.MDFF_1.tspc2_magic_0.QB VSS 0.805288f
C5727 7b_counter_0.MDFF_1.QB.t7 VSS 0.045293f
C5728 7b_counter_0.MDFF_1.QB.t5 VSS 0.086052f
C5729 7b_counter_0.MDFF_1.QB.t3 VSS 0.057347f
C5730 7b_counter_0.MDFF_1.QB.n0 VSS 0.107122f
C5731 7b_counter_0.MDFF_1.QB.t6 VSS 0.108501f
C5732 7b_counter_0.MDFF_1.QB.n1 VSS 0.073647f
C5733 7b_counter_0.MDFF_1.QB.t8 VSS 0.133702f
C5734 7b_counter_0.MDFF_1.QB.n2 VSS 0.140411f
C5735 7b_counter_0.MDFF_1.QB.n3 VSS 0.105327f
C5736 7b_counter_0.MDFF_1.QB.t4 VSS 0.060817f
C5737 7b_counter_0.MDFF_1.QB.t2 VSS 0.072871f
C5738 7b_counter_0.MDFF_1.QB.n4 VSS 0.121822f
C5739 p3_gen_magic_0.xnor_magic_1.OUT.t2 VSS 0.042717f
C5740 p3_gen_magic_0.xnor_magic_1.OUT.t0 VSS 0.041601f
C5741 p3_gen_magic_0.xnor_magic_1.OUT.t1 VSS 0.048345f
C5742 p3_gen_magic_0.xnor_magic_1.OUT.t3 VSS 0.023669f
C5743 p3_gen_magic_0.xnor_magic_1.OUT.t5 VSS 0.044969f
C5744 p3_gen_magic_0.xnor_magic_1.OUT.t6 VSS 0.029968f
C5745 p3_gen_magic_0.xnor_magic_1.OUT.n0 VSS 0.055979f
C5746 p3_gen_magic_0.xnor_magic_1.OUT.t4 VSS 0.0567f
C5747 p3_gen_magic_0.xnor_magic_1.OUT.n1 VSS 0.038486f
C5748 p3_gen_magic_0.xnor_magic_1.OUT.n2 VSS 1.08121f
C5749 7b_counter_0.MDFF_7.QB.t1 VSS 0.211255f
C5750 7b_counter_0.MDFF_7.QB.t0 VSS 0.204984f
C5751 7b_counter_0.MDFF_7.mux_magic_0.IN1 VSS 1.43318f
C5752 7b_counter_0.MDFF_7.tspc2_magic_0.QB VSS 2.81497f
C5753 7b_counter_0.MDFF_7.QB.t8 VSS 0.186134f
C5754 7b_counter_0.MDFF_7.QB.n0 VSS 0.358022f
C5755 7b_counter_0.MDFF_7.QB.t2 VSS 0.339976f
C5756 7b_counter_0.MDFF_7.QB.n1 VSS 0.268795f
C5757 7b_counter_0.MDFF_7.QB.t5 VSS 0.154491f
C5758 7b_counter_0.MDFF_7.QB.n2 VSS 0.310391f
C5759 7b_counter_0.MDFF_7.QB.t7 VSS 0.115403f
C5760 7b_counter_0.MDFF_7.QB.t4 VSS 0.219254f
C5761 7b_counter_0.MDFF_7.QB.t3 VSS 0.146115f
C5762 7b_counter_0.MDFF_7.QB.n3 VSS 0.272937f
C5763 7b_counter_0.MDFF_7.QB.t6 VSS 0.276451f
C5764 7b_counter_0.MDFF_7.QB.n4 VSS 0.187647f
C5765 DFF_magic_0.tg_magic_3.CLK.n0 VSS 0.818913f
C5766 DFF_magic_0.tg_magic_2.CLK VSS 0.867848f
C5767 DFF_magic_0.tg_magic_3.CLK.n1 VSS 0.266613f
C5768 DFF_magic_0.tg_magic_3.CLK.t2 VSS 0.015303f
C5769 DFF_magic_0.tg_magic_3.CLK.t1 VSS 0.015303f
C5770 DFF_magic_0.tg_magic_3.CLK.n2 VSS 0.032993f
C5771 DFF_magic_0.tg_magic_3.CLK.t5 VSS 0.015303f
C5772 DFF_magic_0.tg_magic_3.CLK.t4 VSS 0.015303f
C5773 DFF_magic_0.tg_magic_3.CLK.n3 VSS 0.034488f
C5774 DFF_magic_0.tg_magic_3.CLK.t3 VSS 0.015303f
C5775 DFF_magic_0.tg_magic_3.CLK.t0 VSS 0.015303f
C5776 DFF_magic_0.tg_magic_3.CLK.n4 VSS 0.038656f
C5777 DFF_magic_0.tg_magic_3.CLK.t9 VSS 0.075122f
C5778 DFF_magic_0.tg_magic_3.CLK.t6 VSS 0.075122f
C5779 DFF_magic_0.tg_magic_3.CLK.n5 VSS 0.091325f
C5780 DFF_magic_0.tg_magic_3.CLK.t14 VSS 0.198472f
C5781 DFF_magic_0.tg_magic_3.CLK.t21 VSS 0.036492f
C5782 DFF_magic_0.tg_magic_3.CLK.t19 VSS 0.071049f
C5783 DFF_magic_0.tg_magic_3.CLK.n6 VSS 0.055769f
C5784 DFF_magic_0.tg_magic_3.CLK.t22 VSS 0.071049f
C5785 DFF_magic_0.tg_magic_3.CLK.n7 VSS 0.055769f
C5786 DFF_magic_0.tg_magic_3.CLK.t7 VSS 0.056823f
C5787 DFF_magic_0.tg_magic_3.CLK.t11 VSS 0.076862f
C5788 DFF_magic_0.tg_magic_3.CLK.t15 VSS 0.083823f
C5789 DFF_magic_0.tg_magic_3.CLK.n8 VSS 0.076815f
C5790 DFF_magic_0.tg_magic_3.CLK.t10 VSS 0.075122f
C5791 DFF_magic_0.tg_magic_3.CLK.t17 VSS 0.075122f
C5792 DFF_magic_0.tg_magic_3.CLK.n9 VSS 0.091325f
C5793 DFF_magic_0.tg_magic_3.CLK.t13 VSS 0.198163f
C5794 DFF_magic_0.tg_magic_3.CLK.t16 VSS 0.076862f
C5795 DFF_magic_0.tg_magic_3.CLK.t18 VSS 0.083823f
C5796 DFF_magic_0.tg_magic_3.CLK.t23 VSS 0.071049f
C5797 DFF_magic_0.tg_magic_3.CLK.t8 VSS 0.036492f
C5798 DFF_magic_0.tg_magic_3.CLK.t20 VSS 0.071049f
C5799 DFF_magic_0.tg_magic_3.CLK.n10 VSS 0.055769f
C5800 DFF_magic_0.tg_magic_3.CLK.n11 VSS 0.055769f
C5801 DFF_magic_0.tg_magic_3.CLK.t12 VSS 0.056823f
C5802 DFF_magic_0.tg_magic_3.CLK.n12 VSS 0.076815f
C5803 Q5.t2 VSS 0.092338f
C5804 Q5.t0 VSS 0.07216f
C5805 Q5.n0 VSS 0.185688f
C5806 Q5.t1 VSS 0.079299f
C5807 Q5.n1 VSS 0.142097f
C5808 Q5.t26 VSS 0.069738f
C5809 Q5.t7 VSS 0.132495f
C5810 Q5.t15 VSS 0.088297f
C5811 Q5.n2 VSS 0.164936f
C5812 Q5.t28 VSS 0.167059f
C5813 Q5.n3 VSS 0.113395f
C5814 Q5.n4 VSS 1.36866f
C5815 Q5.n5 VSS 1.06497f
C5816 Q5.n6 VSS 0.014226f
C5817 Q5.t27 VSS 0.101795f
C5818 Q5.t3 VSS 0.16619f
C5819 Q5.t5 VSS 0.264048f
C5820 Q5.t14 VSS 0.243058f
C5821 Q5.t4 VSS 0.179507f
C5822 Q5.n7 VSS 0.235331f
C5823 Q5.t17 VSS 0.146887f
C5824 Q5.t23 VSS 0.16019f
C5825 Q5.t29 VSS 0.069738f
C5826 Q5.t22 VSS 0.135778f
C5827 Q5.n8 VSS 0.106577f
C5828 Q5.t21 VSS 0.135778f
C5829 Q5.n9 VSS 0.106577f
C5830 Q5.t6 VSS 0.108593f
C5831 Q5.n10 VSS 0.147237f
C5832 Q5.t18 VSS 0.096098f
C5833 Q5.t19 VSS 0.149438f
C5834 Q5.t24 VSS 0.178964f
C5835 Q5.n11 VSS 0.123864f
C5836 Q5.n12 VSS 0.863654f
C5837 Q5.t9 VSS 0.146887f
C5838 Q5.t13 VSS 0.16019f
C5839 Q5.t20 VSS 0.069738f
C5840 Q5.t12 VSS 0.135778f
C5841 Q5.n13 VSS 0.106577f
C5842 Q5.t11 VSS 0.135778f
C5843 Q5.n14 VSS 0.106577f
C5844 Q5.t25 VSS 0.108593f
C5845 Q5.n15 VSS 0.147237f
C5846 Q5.t8 VSS 0.096098f
C5847 Q5.t10 VSS 0.149438f
C5848 Q5.t16 VSS 0.178964f
C5849 Q5.n16 VSS 0.123864f
C5850 Q5.n17 VSS 4.97086f
C5851 Q5.n18 VSS 6.22016f
C5852 Q5.n19 VSS 3.25604f
C5853 p3_gen_magic_0.xnor_magic_3.OUT.t0 VSS 0.058254f
C5854 p3_gen_magic_0.xnor_magic_3.OUT.t1 VSS 0.06593f
C5855 p3_gen_magic_0.xnor_magic_3.OUT.n0 VSS 1.20048f
C5856 p3_gen_magic_0.xnor_magic_3.OUT.t6 VSS 0.064556f
C5857 p3_gen_magic_0.xnor_magic_3.OUT.t5 VSS 0.158504f
C5858 p3_gen_magic_0.xnor_magic_3.OUT.t4 VSS 0.045944f
C5859 p3_gen_magic_0.xnor_magic_3.OUT.t2 VSS 0.075358f
C5860 p3_gen_magic_0.xnor_magic_3.OUT.t3 VSS 0.08538f
C5861 p3_gen_magic_0.xnor_magic_3.OUT.n1 VSS 0.061699f
C5862 p3_gen_magic_0.xnor_magic_3.OUT.n2 VSS 0.904176f
C5863 mux_magic_0.IN1.t15 VSS 0.084422f
C5864 mux_magic_0.IN1.t6 VSS 0.160393f
C5865 mux_magic_0.IN1.t7 VSS 0.106889f
C5866 mux_magic_0.IN1.n0 VSS 0.199665f
C5867 mux_magic_0.IN1.t12 VSS 0.202236f
C5868 mux_magic_0.IN1.n1 VSS 0.137271f
C5869 mux_magic_0.IN1.t11 VSS 0.177816f
C5870 mux_magic_0.IN1.t8 VSS 0.19392f
C5871 mux_magic_0.IN1.t13 VSS 0.164368f
C5872 mux_magic_0.IN1.t9 VSS 0.084422f
C5873 mux_magic_0.IN1.t14 VSS 0.164368f
C5874 mux_magic_0.IN1.n2 VSS 0.129018f
C5875 mux_magic_0.IN1.n3 VSS 0.129018f
C5876 mux_magic_0.IN1.t10 VSS 0.131458f
C5877 mux_magic_0.IN1.n4 VSS 0.178282f
C5878 mux_magic_0.IN1.t5 VSS 0.035403f
C5879 mux_magic_0.IN1.t4 VSS 0.035403f
C5880 mux_magic_0.IN1.n5 VSS 0.079786f
C5881 mux_magic_0.IN1.t1 VSS 0.035403f
C5882 mux_magic_0.IN1.t0 VSS 0.035403f
C5883 mux_magic_0.IN1.n6 VSS 0.089429f
C5884 mux_magic_0.IN1.t3 VSS 0.035403f
C5885 mux_magic_0.IN1.t2 VSS 0.035403f
C5886 mux_magic_0.IN1.n7 VSS 0.076328f
C5887 divide_by_2_1.tg_magic_3.IN.n0 VSS 0.138246f
C5888 divide_by_2_1.tg_magic_3.IN.t13 VSS 0.030044f
C5889 divide_by_2_1.tg_magic_3.IN.t8 VSS 0.026526f
C5890 divide_by_2_1.tg_magic_3.IN.t12 VSS 0.010743f
C5891 divide_by_2_1.tg_magic_3.IN.t14 VSS 0.010743f
C5892 divide_by_2_1.tg_magic_3.IN.n1 VSS 0.027357f
C5893 divide_by_2_1.tg_magic_3.IN.t6 VSS 0.010743f
C5894 divide_by_2_1.tg_magic_3.IN.t7 VSS 0.010743f
C5895 divide_by_2_1.tg_magic_3.IN.n2 VSS 0.021485f
C5896 divide_by_2_1.tg_magic_3.IN.n3 VSS 0.077892f
C5897 divide_by_2_1.tg_magic_3.IN.t19 VSS 0.025619f
C5898 divide_by_2_1.tg_magic_3.IN.t18 VSS 0.049879f
C5899 divide_by_2_1.tg_magic_3.IN.n4 VSS 0.039152f
C5900 divide_by_2_1.tg_magic_3.IN.t22 VSS 0.049879f
C5901 divide_by_2_1.tg_magic_3.IN.n5 VSS 0.039152f
C5902 divide_by_2_1.tg_magic_3.IN.t21 VSS 0.039892f
C5903 divide_by_2_1.tg_magic_3.IN.t20 VSS 0.05396f
C5904 divide_by_2_1.tg_magic_3.IN.t23 VSS 0.058847f
C5905 divide_by_2_1.tg_magic_3.IN.n6 VSS 0.054104f
C5906 divide_by_2_1.tg_magic_3.IN.t9 VSS 0.029792f
C5907 divide_by_2_1.tg_magic_3.IN.t15 VSS 0.040014f
C5908 divide_by_2_1.tg_magic_3.IN.t17 VSS 0.010743f
C5909 divide_by_2_1.tg_magic_3.IN.t16 VSS 0.010743f
C5910 divide_by_2_1.tg_magic_3.IN.n7 VSS 0.021487f
C5911 divide_by_2_1.tg_magic_3.IN.t11 VSS 0.010743f
C5912 divide_by_2_1.tg_magic_3.IN.t10 VSS 0.010743f
C5913 divide_by_2_1.tg_magic_3.IN.n8 VSS 0.021487f
C5914 divide_by_2_1.tg_magic_3.IN.t4 VSS 0.030044f
C5915 divide_by_2_1.tg_magic_3.IN.t2 VSS 0.026526f
C5916 divide_by_2_1.tg_magic_3.IN.t1 VSS 0.010743f
C5917 divide_by_2_1.tg_magic_3.IN.t0 VSS 0.010743f
C5918 divide_by_2_1.tg_magic_3.IN.n9 VSS 0.021485f
C5919 divide_by_2_1.tg_magic_3.IN.t3 VSS 0.010743f
C5920 divide_by_2_1.tg_magic_3.IN.t5 VSS 0.010743f
C5921 divide_by_2_1.tg_magic_3.IN.n10 VSS 0.027357f
C5922 divide_by_2_1.tg_magic_3.IN.n11 VSS 0.077892f
C5923 p3_gen_magic_0.xnor_magic_5.OUT.t0 VSS 0.047523f
C5924 p3_gen_magic_0.xnor_magic_5.OUT.t1 VSS 0.055227f
C5925 p3_gen_magic_0.xnor_magic_5.OUT.t5 VSS 0.098153f
C5926 p3_gen_magic_0.xnor_magic_5.OUT.t3 VSS 0.108047f
C5927 p3_gen_magic_0.xnor_magic_5.OUT.t4 VSS 0.05203f
C5928 p3_gen_magic_0.xnor_magic_5.OUT.t2 VSS 0.033888f
C5929 p3_gen_magic_0.xnor_magic_5.OUT.n0 VSS 0.042059f
C5930 p3_gen_magic_0.xnor_magic_5.OUT.n1 VSS 0.046059f
C5931 p3_gen_magic_0.xnor_magic_5.OUT.n2 VSS 0.984703f
C5932 a_31440_8496.n0 VSS 0.175921f
C5933 a_31440_8496.t9 VSS 0.12297f
C5934 a_31440_8496.t12 VSS 0.119549f
C5935 a_31440_8496.t13 VSS 0.197395f
C5936 a_31440_8496.t17 VSS 0.125751f
C5937 a_31440_8496.n1 VSS 0.089259f
C5938 a_31440_8496.t16 VSS 0.174488f
C5939 a_31440_8496.t11 VSS 0.197395f
C5940 a_31440_8496.t10 VSS 0.169773f
C5941 a_31440_8496.n2 VSS 0.091907f
C5942 a_31440_8496.t14 VSS 0.169773f
C5943 a_31440_8496.t15 VSS 0.141829f
C5944 a_31440_8496.n3 VSS 0.159639f
C5945 a_31440_8496.t8 VSS 0.058483f
C5946 a_31440_8496.t2 VSS 0.054881f
C5947 a_31440_8496.n4 VSS 0.113139f
C5948 a_31440_8496.t1 VSS 0.022242f
C5949 a_31440_8496.t0 VSS 0.022242f
C5950 a_31440_8496.n5 VSS 0.044484f
C5951 a_31440_8496.n6 VSS 0.115439f
C5952 a_31440_8496.t4 VSS 0.022242f
C5953 a_31440_8496.t3 VSS 0.022242f
C5954 a_31440_8496.n7 VSS 0.044484f
C5955 a_31440_8496.n8 VSS 0.077993f
C5956 a_31440_8496.t7 VSS 0.022242f
C5957 a_31440_8496.t6 VSS 0.022242f
C5958 a_31440_8496.n9 VSS 0.044456f
C5959 a_31440_8496.n10 VSS 0.10201f
C5960 a_31440_8496.n11 VSS 0.120648f
C5961 a_31440_8496.t5 VSS 0.054881f
C5962 a_27567_8496.n0 VSS 0.175921f
C5963 a_27567_8496.t17 VSS 0.12297f
C5964 a_27567_8496.t11 VSS 0.119549f
C5965 a_27567_8496.t12 VSS 0.197395f
C5966 a_27567_8496.t16 VSS 0.125751f
C5967 a_27567_8496.n1 VSS 0.089259f
C5968 a_27567_8496.t15 VSS 0.174488f
C5969 a_27567_8496.t10 VSS 0.197395f
C5970 a_27567_8496.t9 VSS 0.169773f
C5971 a_27567_8496.n2 VSS 0.091907f
C5972 a_27567_8496.t13 VSS 0.169773f
C5973 a_27567_8496.t14 VSS 0.141829f
C5974 a_27567_8496.n3 VSS 0.159639f
C5975 a_27567_8496.t8 VSS 0.058483f
C5976 a_27567_8496.t2 VSS 0.054881f
C5977 a_27567_8496.n4 VSS 0.113139f
C5978 a_27567_8496.t1 VSS 0.022242f
C5979 a_27567_8496.t0 VSS 0.022242f
C5980 a_27567_8496.n5 VSS 0.044484f
C5981 a_27567_8496.n6 VSS 0.115439f
C5982 a_27567_8496.t4 VSS 0.022242f
C5983 a_27567_8496.t3 VSS 0.022242f
C5984 a_27567_8496.n7 VSS 0.044484f
C5985 a_27567_8496.n8 VSS 0.077993f
C5986 a_27567_8496.t7 VSS 0.022242f
C5987 a_27567_8496.t6 VSS 0.022242f
C5988 a_27567_8496.n9 VSS 0.044456f
C5989 a_27567_8496.n10 VSS 0.10201f
C5990 a_27567_8496.n11 VSS 0.120648f
C5991 a_27567_8496.t5 VSS 0.054881f
C5992 divide_by_2_0.tg_magic_3.IN.n0 VSS 0.122295f
C5993 divide_by_2_0.tg_magic_3.IN.t8 VSS 0.026577f
C5994 divide_by_2_0.tg_magic_3.IN.t10 VSS 0.023465f
C5995 divide_by_2_0.tg_magic_3.IN.t7 VSS 0.009504f
C5996 divide_by_2_0.tg_magic_3.IN.t9 VSS 0.009504f
C5997 divide_by_2_0.tg_magic_3.IN.n1 VSS 0.0242f
C5998 divide_by_2_0.tg_magic_3.IN.t12 VSS 0.009504f
C5999 divide_by_2_0.tg_magic_3.IN.t11 VSS 0.009504f
C6000 divide_by_2_0.tg_magic_3.IN.n2 VSS 0.019006f
C6001 divide_by_2_0.tg_magic_3.IN.n3 VSS 0.068905f
C6002 divide_by_2_0.tg_magic_3.IN.t19 VSS 0.022663f
C6003 divide_by_2_0.tg_magic_3.IN.t23 VSS 0.044124f
C6004 divide_by_2_0.tg_magic_3.IN.n4 VSS 0.034634f
C6005 divide_by_2_0.tg_magic_3.IN.t18 VSS 0.044124f
C6006 divide_by_2_0.tg_magic_3.IN.n5 VSS 0.034634f
C6007 divide_by_2_0.tg_magic_3.IN.t21 VSS 0.035289f
C6008 divide_by_2_0.tg_magic_3.IN.t22 VSS 0.047734f
C6009 divide_by_2_0.tg_magic_3.IN.t20 VSS 0.052057f
C6010 divide_by_2_0.tg_magic_3.IN.n6 VSS 0.047861f
C6011 divide_by_2_0.tg_magic_3.IN.t5 VSS 0.026354f
C6012 divide_by_2_0.tg_magic_3.IN.t16 VSS 0.035397f
C6013 divide_by_2_0.tg_magic_3.IN.t15 VSS 0.009504f
C6014 divide_by_2_0.tg_magic_3.IN.t17 VSS 0.009504f
C6015 divide_by_2_0.tg_magic_3.IN.n7 VSS 0.019007f
C6016 divide_by_2_0.tg_magic_3.IN.t4 VSS 0.009504f
C6017 divide_by_2_0.tg_magic_3.IN.t6 VSS 0.009504f
C6018 divide_by_2_0.tg_magic_3.IN.n8 VSS 0.019007f
C6019 divide_by_2_0.tg_magic_3.IN.t14 VSS 0.026577f
C6020 divide_by_2_0.tg_magic_3.IN.t1 VSS 0.023465f
C6021 divide_by_2_0.tg_magic_3.IN.t0 VSS 0.009504f
C6022 divide_by_2_0.tg_magic_3.IN.t2 VSS 0.009504f
C6023 divide_by_2_0.tg_magic_3.IN.n9 VSS 0.019006f
C6024 divide_by_2_0.tg_magic_3.IN.t3 VSS 0.009504f
C6025 divide_by_2_0.tg_magic_3.IN.t13 VSS 0.009504f
C6026 divide_by_2_0.tg_magic_3.IN.n10 VSS 0.0242f
C6027 divide_by_2_0.tg_magic_3.IN.n11 VSS 0.068905f
C6028 OR_magic_1.VOUT.n0 VSS 1.29647f
C6029 OR_magic_1.VOUT.t6 VSS 0.059172f
C6030 OR_magic_1.VOUT.t4 VSS 0.115207f
C6031 OR_magic_1.VOUT.n1 VSS 0.09043f
C6032 OR_magic_1.VOUT.t10 VSS 0.115207f
C6033 OR_magic_1.VOUT.n2 VSS 0.09043f
C6034 OR_magic_1.VOUT.t16 VSS 0.09214f
C6035 OR_magic_1.VOUT.t14 VSS 0.124633f
C6036 OR_magic_1.VOUT.t22 VSS 0.135921f
C6037 OR_magic_1.VOUT.n3 VSS 0.124965f
C6038 OR_magic_1.VOUT.t21 VSS 0.121812f
C6039 OR_magic_1.VOUT.t5 VSS 0.121812f
C6040 OR_magic_1.VOUT.n4 VSS 0.148085f
C6041 OR_magic_1.VOUT.t23 VSS 0.321827f
C6042 OR_magic_1.VOUT.t12 VSS 0.059172f
C6043 OR_magic_1.VOUT.t8 VSS 0.115207f
C6044 OR_magic_1.VOUT.n5 VSS 0.09043f
C6045 OR_magic_1.VOUT.t20 VSS 0.115207f
C6046 OR_magic_1.VOUT.n6 VSS 0.09043f
C6047 OR_magic_1.VOUT.t18 VSS 0.09214f
C6048 OR_magic_1.VOUT.t17 VSS 0.124633f
C6049 OR_magic_1.VOUT.t24 VSS 0.135921f
C6050 OR_magic_1.VOUT.n7 VSS 0.124557f
C6051 OR_magic_1.VOUT.t25 VSS 0.121812f
C6052 OR_magic_1.VOUT.t9 VSS 0.121812f
C6053 OR_magic_1.VOUT.n8 VSS 0.148085f
C6054 OR_magic_1.VOUT.t11 VSS 0.181198f
C6055 OR_magic_1.VOUT.t15 VSS 0.124633f
C6056 OR_magic_1.VOUT.t13 VSS 0.135921f
C6057 OR_magic_1.VOUT.t19 VSS 0.115207f
C6058 OR_magic_1.VOUT.t2 VSS 0.059172f
C6059 OR_magic_1.VOUT.t3 VSS 0.115207f
C6060 OR_magic_1.VOUT.n9 VSS 0.09043f
C6061 OR_magic_1.VOUT.n10 VSS 0.09043f
C6062 OR_magic_1.VOUT.t7 VSS 0.09214f
C6063 OR_magic_1.VOUT.n11 VSS 0.124557f
C6064 OR_magic_1.VOUT.n12 VSS 0.668982f
C6065 OR_magic_1.VOUT.t1 VSS 0.078348f
C6066 OR_magic_1.VOUT.t0 VSS 0.061228f
C6067 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n0 VSS 0.239198f
C6068 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t0 VSS 0.051546f
C6069 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t10 VSS 0.069234f
C6070 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t8 VSS 0.018588f
C6071 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t9 VSS 0.018588f
C6072 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n1 VSS 0.037177f
C6073 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t1 VSS 0.018588f
C6074 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t2 VSS 0.018588f
C6075 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.n2 VSS 0.037177f
C6076 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t3 VSS 0.072331f
C6077 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t4 VSS 0.094887f
C6078 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t5 VSS 0.050609f
C6079 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t7 VSS 0.058782f
C6080 p3_gen_magic_0.3_inp_AND_magic_0.VOUT.t6 VSS 0.045866f
C6081 p2_gen_magic_0.3_inp_AND_magic_0.C.t0 VSS 0.075145f
C6082 p2_gen_magic_0.3_inp_AND_magic_0.C.t3 VSS 0.078354f
C6083 p2_gen_magic_0.3_inp_AND_magic_0.C.t5 VSS 0.192384f
C6084 p2_gen_magic_0.3_inp_AND_magic_0.C.t4 VSS 0.055764f
C6085 p2_gen_magic_0.3_inp_AND_magic_0.C.t2 VSS 0.091466f
C6086 p2_gen_magic_0.3_inp_AND_magic_0.C.t1 VSS 0.10363f
C6087 p2_gen_magic_0.3_inp_AND_magic_0.C.n0 VSS 0.074887f
C6088 p2_gen_magic_0.3_inp_AND_magic_0.C.n1 VSS 0.597027f
C6089 OR_magic_2.A.n0 VSS 0.591818f
C6090 OR_magic_2.A.n1 VSS 0.209532f
C6091 OR_magic_2.A.t15 VSS 0.094181f
C6092 OR_magic_2.A.t18 VSS 0.122432f
C6093 OR_magic_2.A.t12 VSS 0.100447f
C6094 OR_magic_2.A.t21 VSS 0.161133f
C6095 OR_magic_2.A.t13 VSS 0.116839f
C6096 OR_magic_2.A.n2 VSS 0.083748f
C6097 OR_magic_2.A.t16 VSS 0.091092f
C6098 OR_magic_2.A.t11 VSS 0.099342f
C6099 OR_magic_2.A.t17 VSS 0.084203f
C6100 OR_magic_2.A.t8 VSS 0.043248f
C6101 OR_magic_2.A.t14 VSS 0.084203f
C6102 OR_magic_2.A.n3 VSS 0.066094f
C6103 OR_magic_2.A.n4 VSS 0.066094f
C6104 OR_magic_2.A.t7 VSS 0.067344f
C6105 OR_magic_2.A.n5 VSS 0.091331f
C6106 OR_magic_2.A.t19 VSS 0.094181f
C6107 OR_magic_2.A.t6 VSS 0.122432f
C6108 OR_magic_2.A.t9 VSS 0.100447f
C6109 OR_magic_2.A.t20 VSS 0.161133f
C6110 OR_magic_2.A.t10 VSS 0.116839f
C6111 OR_magic_2.A.n6 VSS 0.083778f
C6112 OR_magic_2.A.t5 VSS 0.018136f
C6113 OR_magic_2.A.t4 VSS 0.018136f
C6114 OR_magic_2.A.n7 VSS 0.040873f
C6115 OR_magic_2.A.t2 VSS 0.018136f
C6116 OR_magic_2.A.t1 VSS 0.018136f
C6117 OR_magic_2.A.n8 VSS 0.045813f
C6118 OR_magic_2.A.t0 VSS 0.018136f
C6119 OR_magic_2.A.t3 VSS 0.018136f
C6120 OR_magic_2.A.n9 VSS 0.039102f
C6121 Q4.t11 VSS 0.085483f
C6122 Q4.t13 VSS 0.170416f
C6123 Q4.t21 VSS 0.238131f
C6124 Q4.t22 VSS 0.238131f
C6125 Q4.t14 VSS 0.209997f
C6126 Q4.n0 VSS 0.184173f
C6127 Q4.n1 VSS 1.03679f
C6128 Q4.t2 VSS 0.090257f
C6129 Q4.t1 VSS 0.070534f
C6130 Q4.n2 VSS 0.181503f
C6131 Q4.t0 VSS 0.077512f
C6132 Q4.n3 VSS 0.138895f
C6133 Q4.t6 VSS 0.093933f
C6134 Q4.t7 VSS 0.146071f
C6135 Q4.t12 VSS 0.174932f
C6136 Q4.n4 VSS 0.121073f
C6137 Q4.t16 VSS 0.143578f
C6138 Q4.t20 VSS 0.156581f
C6139 Q4.t26 VSS 0.068167f
C6140 Q4.t10 VSS 0.132719f
C6141 Q4.n5 VSS 0.104176f
C6142 Q4.t19 VSS 0.132719f
C6143 Q4.n6 VSS 0.104176f
C6144 Q4.t5 VSS 0.106146f
C6145 Q4.n7 VSS 0.143919f
C6146 Q4.n8 VSS 2.06922f
C6147 Q4.t25 VSS 0.143578f
C6148 Q4.t29 VSS 0.156581f
C6149 Q4.t8 VSS 0.068167f
C6150 Q4.t24 VSS 0.132719f
C6151 Q4.n9 VSS 0.104176f
C6152 Q4.t28 VSS 0.132719f
C6153 Q4.n10 VSS 0.104176f
C6154 Q4.t15 VSS 0.106146f
C6155 Q4.n11 VSS 0.143919f
C6156 Q4.t17 VSS 0.093933f
C6157 Q4.t18 VSS 0.146071f
C6158 Q4.t23 VSS 0.174932f
C6159 Q4.n12 VSS 0.121073f
C6160 Q4.n13 VSS 1.07244f
C6161 Q4.n14 VSS 4.95909f
C6162 Q4.t9 VSS 0.068167f
C6163 Q4.t4 VSS 0.129509f
C6164 Q4.t27 VSS 0.086308f
C6165 Q4.n15 VSS 0.161219f
C6166 Q4.t3 VSS 0.163295f
C6167 Q4.n16 VSS 0.11084f
C6168 Q4.n17 VSS 2.38309f
C6169 Q4.n18 VSS 4.95738f
C6170 Q4.n19 VSS 0.210031f
C6171 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n0 VSS 0.857909f
C6172 7b_counter_0.DFF_magic_0.tg_magic_2.CLK VSS 0.909175f
C6173 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n1 VSS 0.279308f
C6174 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t5 VSS 0.016032f
C6175 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t4 VSS 0.016032f
C6176 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n2 VSS 0.03613f
C6177 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t0 VSS 0.016032f
C6178 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t1 VSS 0.016032f
C6179 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n3 VSS 0.040497f
C6180 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t3 VSS 0.016032f
C6181 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t2 VSS 0.016032f
C6182 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n4 VSS 0.034564f
C6183 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t18 VSS 0.078699f
C6184 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t7 VSS 0.078699f
C6185 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n5 VSS 0.095673f
C6186 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t21 VSS 0.207923f
C6187 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t9 VSS 0.038229f
C6188 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t23 VSS 0.074432f
C6189 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n6 VSS 0.058424f
C6190 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t10 VSS 0.074432f
C6191 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n7 VSS 0.058424f
C6192 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t11 VSS 0.059529f
C6193 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t15 VSS 0.080522f
C6194 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t17 VSS 0.087815f
C6195 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n8 VSS 0.080473f
C6196 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t13 VSS 0.078699f
C6197 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t16 VSS 0.078699f
C6198 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n9 VSS 0.095673f
C6199 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t14 VSS 0.2076f
C6200 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t22 VSS 0.080522f
C6201 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t20 VSS 0.087815f
C6202 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t19 VSS 0.074432f
C6203 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t8 VSS 0.038229f
C6204 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t12 VSS 0.074432f
C6205 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n10 VSS 0.058424f
C6206 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n11 VSS 0.058424f
C6207 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.t6 VSS 0.059529f
C6208 7b_counter_0.DFF_magic_0.tg_magic_3.CLK.n12 VSS 0.080473f
C6209 7b_counter_0.MDFF_4.QB.t1 VSS 0.083008f
C6210 7b_counter_0.MDFF_4.QB.t0 VSS 0.080545f
C6211 7b_counter_0.MDFF_4.mux_magic_0.IN1 VSS 0.842894f
C6212 7b_counter_0.MDFF_4.tspc2_magic_0.QB VSS 0.879351f
C6213 7b_counter_0.MDFF_4.QB.n0 VSS 0.140678f
C6214 7b_counter_0.MDFF_4.QB.t7 VSS 0.133805f
C6215 7b_counter_0.MDFF_4.QB.n1 VSS 0.1054f
C6216 7b_counter_0.MDFF_4.QB.t5 VSS 0.060887f
C6217 7b_counter_0.MDFF_4.QB.t8 VSS 0.072955f
C6218 7b_counter_0.MDFF_4.QB.n2 VSS 0.121962f
C6219 7b_counter_0.MDFF_4.QB.t3 VSS 0.045345f
C6220 7b_counter_0.MDFF_4.QB.t4 VSS 0.086152f
C6221 7b_counter_0.MDFF_4.QB.t2 VSS 0.057413f
C6222 7b_counter_0.MDFF_4.QB.n3 VSS 0.107246f
C6223 7b_counter_0.MDFF_4.QB.t6 VSS 0.108626f
C6224 7b_counter_0.MDFF_4.QB.n4 VSS 0.073732f
C6225 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t2 VSS 0.039741f
C6226 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t0 VSS 0.031057f
C6227 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t1 VSS 0.034129f
C6228 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t5 VSS 0.110718f
C6229 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t10 VSS 0.056192f
C6230 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t3 VSS 0.037155f
C6231 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n0 VSS 0.09845f
C6232 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n1 VSS 0.140921f
C6233 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t9 VSS 0.070462f
C6234 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t4 VSS 0.0385f
C6235 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t7 VSS 0.030014f
C6236 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t6 VSS 0.060221f
C6237 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n2 VSS 0.06393f
C6238 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t8 VSS 0.076733f
C6239 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n3 VSS 0.093075f
C6240 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n4 VSS 0.252841f
C6241 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t11 VSS 0.030014f
C6242 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.t12 VSS 0.059765f
C6243 7b_counter_0.MDFF_4.tspc2_magic_0.CLK.n5 VSS 0.059173f
C6244 Q7.t9 VSS 0.071154f
C6245 Q7.t10 VSS 0.116166f
C6246 Q7.t11 VSS 0.184568f
C6247 Q7.t19 VSS 0.169896f
C6248 Q7.t17 VSS 0.125474f
C6249 Q7.n0 VSS 0.114017f
C6250 Q7.n1 VSS 2.73712f
C6251 Q7.t16 VSS 0.067172f
C6252 Q7.t12 VSS 0.104457f
C6253 Q7.t24 VSS 0.125095f
C6254 Q7.n2 VSS 0.08658f
C6255 Q7.t21 VSS 0.102674f
C6256 Q7.t25 VSS 0.111972f
C6257 Q7.t5 VSS 0.048746f
C6258 Q7.t13 VSS 0.094908f
C6259 Q7.n3 VSS 0.074497f
C6260 Q7.t14 VSS 0.094908f
C6261 Q7.n4 VSS 0.074497f
C6262 Q7.t8 VSS 0.075906f
C6263 Q7.n5 VSS 0.102918f
C6264 Q7.n6 VSS 1.35497f
C6265 Q7.t4 VSS 0.102674f
C6266 Q7.t7 VSS 0.111972f
C6267 Q7.t15 VSS 0.048746f
C6268 Q7.t22 VSS 0.094908f
C6269 Q7.n7 VSS 0.074497f
C6270 Q7.t23 VSS 0.094908f
C6271 Q7.n8 VSS 0.074497f
C6272 Q7.t18 VSS 0.075906f
C6273 Q7.n9 VSS 0.102918f
C6274 Q7.t3 VSS 0.067172f
C6275 Q7.t20 VSS 0.104457f
C6276 Q7.t6 VSS 0.125095f
C6277 Q7.n10 VSS 0.08658f
C6278 Q7.n11 VSS 0.384844f
C6279 Q7.n12 VSS 3.78064f
C6280 Q7.n13 VSS 5.14303f
C6281 Q7.n14 VSS 0.010199f
C6282 Q7.t2 VSS 0.064544f
C6283 Q7.t0 VSS 0.05044f
C6284 Q7.n15 VSS 0.129795f
C6285 Q7.t1 VSS 0.055429f
C6286 Q7.n16 VSS 0.099325f
C6287 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n0 VSS 0.838411f
C6288 p2_gen_magic_0.DFF_magic_0.tg_magic_2.CLK VSS 0.888512f
C6289 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n1 VSS 0.27296f
C6290 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t4 VSS 0.015667f
C6291 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t5 VSS 0.015667f
C6292 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n2 VSS 0.035309f
C6293 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t1 VSS 0.015667f
C6294 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t0 VSS 0.015667f
C6295 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n3 VSS 0.039577f
C6296 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t2 VSS 0.015667f
C6297 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t3 VSS 0.015667f
C6298 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n4 VSS 0.033779f
C6299 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t8 VSS 0.076911f
C6300 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t15 VSS 0.076911f
C6301 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n5 VSS 0.093499f
C6302 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t7 VSS 0.203197f
C6303 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t13 VSS 0.037361f
C6304 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t14 VSS 0.07274f
C6305 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n6 VSS 0.057096f
C6306 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t21 VSS 0.07274f
C6307 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n7 VSS 0.057096f
C6308 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t20 VSS 0.058176f
C6309 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t19 VSS 0.078692f
C6310 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t23 VSS 0.085819f
C6311 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n8 VSS 0.078644f
C6312 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t10 VSS 0.076911f
C6313 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t16 VSS 0.076911f
C6314 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n9 VSS 0.093499f
C6315 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t12 VSS 0.202882f
C6316 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t6 VSS 0.078692f
C6317 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t17 VSS 0.085819f
C6318 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t22 VSS 0.07274f
C6319 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t18 VSS 0.037361f
C6320 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t9 VSS 0.07274f
C6321 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n10 VSS 0.057096f
C6322 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n11 VSS 0.057096f
C6323 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.t11 VSS 0.058176f
C6324 p2_gen_magic_0.DFF_magic_0.tg_magic_3.CLK.n12 VSS 0.078644f
C6325 divide_by_2_0.tg_magic_3.CLK.t1 VSS 1.21872f
C6326 divide_by_2_0.tg_magic_2.CLK VSS 0.867848f
C6327 divide_by_2_0.tg_magic_3.CLK.t0 VSS 0.064766f
C6328 divide_by_2_0.tg_magic_3.CLK.t17 VSS 0.075122f
C6329 divide_by_2_0.tg_magic_3.CLK.t12 VSS 0.075122f
C6330 divide_by_2_0.tg_magic_3.CLK.n0 VSS 0.091325f
C6331 divide_by_2_0.tg_magic_3.CLK.t9 VSS 0.198472f
C6332 divide_by_2_0.tg_magic_3.CLK.t8 VSS 0.036492f
C6333 divide_by_2_0.tg_magic_3.CLK.t15 VSS 0.071049f
C6334 divide_by_2_0.tg_magic_3.CLK.n1 VSS 0.055769f
C6335 divide_by_2_0.tg_magic_3.CLK.t3 VSS 0.071049f
C6336 divide_by_2_0.tg_magic_3.CLK.n2 VSS 0.055769f
C6337 divide_by_2_0.tg_magic_3.CLK.t11 VSS 0.056823f
C6338 divide_by_2_0.tg_magic_3.CLK.t19 VSS 0.076862f
C6339 divide_by_2_0.tg_magic_3.CLK.t6 VSS 0.083823f
C6340 divide_by_2_0.tg_magic_3.CLK.n3 VSS 0.076815f
C6341 divide_by_2_0.tg_magic_3.CLK.t18 VSS 0.075122f
C6342 divide_by_2_0.tg_magic_3.CLK.t7 VSS 0.075122f
C6343 divide_by_2_0.tg_magic_3.CLK.n4 VSS 0.091325f
C6344 divide_by_2_0.tg_magic_3.CLK.t4 VSS 0.198163f
C6345 divide_by_2_0.tg_magic_3.CLK.t16 VSS 0.076862f
C6346 divide_by_2_0.tg_magic_3.CLK.t10 VSS 0.083823f
C6347 divide_by_2_0.tg_magic_3.CLK.t2 VSS 0.071049f
C6348 divide_by_2_0.tg_magic_3.CLK.t13 VSS 0.036492f
C6349 divide_by_2_0.tg_magic_3.CLK.t14 VSS 0.071049f
C6350 divide_by_2_0.tg_magic_3.CLK.n5 VSS 0.055769f
C6351 divide_by_2_0.tg_magic_3.CLK.n6 VSS 0.055769f
C6352 divide_by_2_0.tg_magic_3.CLK.t5 VSS 0.056823f
C6353 divide_by_2_0.tg_magic_3.CLK.n7 VSS 0.076815f
C6354 Q6.t1 VSS 0.057651f
C6355 Q6.t2 VSS 0.06713f
C6356 Q6.t0 VSS 0.052461f
C6357 Q6.n0 VSS 0.134997f
C6358 Q6.n1 VSS 0.103306f
C6359 Q6.t8 VSS 0.063579f
C6360 Q6.t25 VSS 0.12675f
C6361 Q6.t4 VSS 0.177114f
C6362 Q6.t15 VSS 0.177114f
C6363 Q6.t11 VSS 0.156189f
C6364 Q6.n2 VSS 0.137326f
C6365 Q6.t18 VSS 0.0507f
C6366 Q6.t20 VSS 0.096325f
C6367 Q6.t22 VSS 0.064193f
C6368 Q6.n3 VSS 0.11991f
C6369 Q6.t12 VSS 0.121454f
C6370 Q6.n4 VSS 0.082439f
C6371 Q6.n5 VSS 0.799601f
C6372 Q6.n6 VSS 3.99438f
C6373 Q6.t19 VSS 0.106788f
C6374 Q6.t24 VSS 0.11646f
C6375 Q6.t3 VSS 0.0507f
C6376 Q6.t26 VSS 0.098712f
C6377 Q6.n7 VSS 0.077482f
C6378 Q6.t23 VSS 0.098712f
C6379 Q6.n8 VSS 0.077482f
C6380 Q6.t9 VSS 0.078948f
C6381 Q6.n9 VSS 0.107042f
C6382 Q6.t17 VSS 0.069864f
C6383 Q6.t13 VSS 0.108643f
C6384 Q6.t27 VSS 0.130109f
C6385 Q6.n10 VSS 0.09005f
C6386 Q6.n11 VSS 1.11258f
C6387 Q6.t29 VSS 0.106788f
C6388 Q6.t5 VSS 0.11646f
C6389 Q6.t14 VSS 0.0507f
C6390 Q6.t10 VSS 0.098712f
C6391 Q6.n12 VSS 0.077482f
C6392 Q6.t6 VSS 0.098712f
C6393 Q6.n13 VSS 0.077482f
C6394 Q6.t16 VSS 0.078948f
C6395 Q6.n14 VSS 0.107042f
C6396 Q6.t28 VSS 0.069864f
C6397 Q6.t21 VSS 0.108643f
C6398 Q6.t7 VSS 0.130109f
C6399 Q6.n15 VSS 0.09005f
C6400 Q6.n16 VSS 0.468678f
C6401 Q6.n17 VSS 2.46231f
C6402 divide_by_2_1.inverter_magic_5.VOUT VSS 1.28348f
C6403 divide_by_2_1.tg_magic_2.CLK VSS 0.867848f
C6404 divide_by_2_1.tg_magic_3.CLK.t5 VSS 0.075122f
C6405 divide_by_2_1.tg_magic_3.CLK.t7 VSS 0.075122f
C6406 divide_by_2_1.tg_magic_3.CLK.n0 VSS 0.091325f
C6407 divide_by_2_1.tg_magic_3.CLK.t6 VSS 0.198472f
C6408 divide_by_2_1.tg_magic_3.CLK.t12 VSS 0.036492f
C6409 divide_by_2_1.tg_magic_3.CLK.t8 VSS 0.071049f
C6410 divide_by_2_1.tg_magic_3.CLK.n1 VSS 0.055769f
C6411 divide_by_2_1.tg_magic_3.CLK.t13 VSS 0.071049f
C6412 divide_by_2_1.tg_magic_3.CLK.n2 VSS 0.055769f
C6413 divide_by_2_1.tg_magic_3.CLK.t14 VSS 0.056823f
C6414 divide_by_2_1.tg_magic_3.CLK.t0 VSS 0.076862f
C6415 divide_by_2_1.tg_magic_3.CLK.t1 VSS 0.083823f
C6416 divide_by_2_1.tg_magic_3.CLK.n3 VSS 0.076815f
C6417 divide_by_2_1.tg_magic_3.CLK.t16 VSS 0.075122f
C6418 divide_by_2_1.tg_magic_3.CLK.t9 VSS 0.075122f
C6419 divide_by_2_1.tg_magic_3.CLK.n4 VSS 0.091325f
C6420 divide_by_2_1.tg_magic_3.CLK.t4 VSS 0.198163f
C6421 divide_by_2_1.tg_magic_3.CLK.t11 VSS 0.076862f
C6422 divide_by_2_1.tg_magic_3.CLK.t2 VSS 0.083823f
C6423 divide_by_2_1.tg_magic_3.CLK.t15 VSS 0.071049f
C6424 divide_by_2_1.tg_magic_3.CLK.t3 VSS 0.036492f
C6425 divide_by_2_1.tg_magic_3.CLK.t17 VSS 0.071049f
C6426 divide_by_2_1.tg_magic_3.CLK.n5 VSS 0.055769f
C6427 divide_by_2_1.tg_magic_3.CLK.n6 VSS 0.055769f
C6428 divide_by_2_1.tg_magic_3.CLK.t10 VSS 0.056823f
C6429 divide_by_2_1.tg_magic_3.CLK.n7 VSS 0.076815f
C6430 D2_5.t0 VSS 0.077436f
C6431 D2_5.t24 VSS 0.14712f
C6432 D2_5.t3 VSS 0.098044f
C6433 D2_5.n0 VSS 0.183142f
C6434 D2_5.t15 VSS 0.1855f
C6435 D2_5.n1 VSS 0.125912f
C6436 D2_5.t21 VSS 0.077436f
C6437 D2_5.t25 VSS 0.14712f
C6438 D2_5.t4 VSS 0.098044f
C6439 D2_5.n2 VSS 0.183142f
C6440 D2_5.t14 VSS 0.1855f
C6441 D2_5.n3 VSS 0.125912f
C6442 D2_5.t23 VSS 0.163102f
C6443 D2_5.t5 VSS 0.177873f
C6444 D2_5.t8 VSS 0.077436f
C6445 D2_5.t1 VSS 0.150766f
C6446 D2_5.n4 VSS 0.118342f
C6447 D2_5.t22 VSS 0.150766f
C6448 D2_5.n5 VSS 0.118342f
C6449 D2_5.t12 VSS 0.12058f
C6450 D2_5.n6 VSS 0.163512f
C6451 D2_5.t11 VSS 0.102415f
C6452 D2_5.t13 VSS 0.165934f
C6453 D2_5.t16 VSS 0.203091f
C6454 D2_5.n7 VSS 0.143451f
C6455 D2_5.n8 VSS 1.85466f
C6456 D2_5.t6 VSS 0.163102f
C6457 D2_5.t10 VSS 0.177873f
C6458 D2_5.t17 VSS 0.077436f
C6459 D2_5.t9 VSS 0.150766f
C6460 D2_5.n9 VSS 0.118342f
C6461 D2_5.t7 VSS 0.150766f
C6462 D2_5.n10 VSS 0.118342f
C6463 D2_5.t19 VSS 0.12058f
C6464 D2_5.n11 VSS 0.163512f
C6465 D2_5.t18 VSS 0.102415f
C6466 D2_5.t20 VSS 0.165934f
C6467 D2_5.t2 VSS 0.203091f
C6468 D2_5.n12 VSS 0.143451f
C6469 D2_5.n13 VSS 2.13521f
C6470 D2_5.n14 VSS 7.14352f
C6471 D2_5.n15 VSS -3.90333f
C6472 D2_5.n16 VSS -3.35696f
C6473 p3_gen_magic_0.3_inp_AND_magic_0.C.t0 VSS 0.072255f
C6474 p3_gen_magic_0.3_inp_AND_magic_0.C.t3 VSS 0.075341f
C6475 p3_gen_magic_0.3_inp_AND_magic_0.C.t2 VSS 0.184985f
C6476 p3_gen_magic_0.3_inp_AND_magic_0.C.t5 VSS 0.053619f
C6477 p3_gen_magic_0.3_inp_AND_magic_0.C.t1 VSS 0.087948f
C6478 p3_gen_magic_0.3_inp_AND_magic_0.C.t4 VSS 0.099644f
C6479 p3_gen_magic_0.3_inp_AND_magic_0.C.n0 VSS 0.072007f
C6480 p3_gen_magic_0.3_inp_AND_magic_0.C.n1 VSS 0.574065f
C6481 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t10 VSS 0.034107f
C6482 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t5 VSS 0.068433f
C6483 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n0 VSS 0.072648f
C6484 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t12 VSS 0.087197f
C6485 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t7 VSS 0.04375f
C6486 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n1 VSS 0.105769f
C6487 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t3 VSS 0.125816f
C6488 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t4 VSS 0.063854f
C6489 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t6 VSS 0.042221f
C6490 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n2 VSS 0.111875f
C6491 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n3 VSS 0.160137f
C6492 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t11 VSS 0.080066f
C6493 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n4 VSS 0.287322f
C6494 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t9 VSS 0.034107f
C6495 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t8 VSS 0.067915f
C6496 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.n5 VSS 0.067242f
C6497 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t2 VSS 0.04516f
C6498 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t0 VSS 0.035292f
C6499 7b_counter_0.MDFF_3.tspc2_magic_0.CLK.t1 VSS 0.038783f
C6500 7b_counter_0.MDFF_4.LD.n0 VSS 1.70539f
C6501 7b_counter_0.MDFF_4.LD.n1 VSS 0.146301f
C6502 7b_counter_0.MDFF_4.LD.t0 VSS 0.10268f
C6503 7b_counter_0.MDFF_4.LD.t3 VSS 0.08053f
C6504 7b_counter_0.MDFF_4.LD.t4 VSS 0.075104f
C6505 7b_counter_0.MDFF_4.LD.n2 VSS 0.266922f
C6506 7b_counter_0.MDFF_4.LD.t79 VSS 0.080178f
C6507 7b_counter_0.MDFF_4.LD.t57 VSS 0.080178f
C6508 7b_counter_0.MDFF_4.LD.n3 VSS 0.102651f
C6509 7b_counter_0.MDFF_4.LD.t72 VSS 0.080178f
C6510 7b_counter_0.MDFF_4.LD.t45 VSS 0.080178f
C6511 7b_counter_0.MDFF_4.LD.n4 VSS 0.11396f
C6512 7b_counter_0.MDFF_4.LD.t46 VSS 0.080178f
C6513 7b_counter_0.MDFF_4.LD.n5 VSS 0.102651f
C6514 7b_counter_0.MDFF_4.LD.t19 VSS 0.102253f
C6515 7b_counter_0.MDFF_4.LD.t121 VSS 0.062925f
C6516 7b_counter_0.MDFF_4.LD.t30 VSS 0.121066f
C6517 7b_counter_0.MDFF_4.LD.t108 VSS 0.079119f
C6518 7b_counter_0.MDFF_4.LD.n6 VSS 0.098158f
C6519 7b_counter_0.MDFF_4.LD.t111 VSS 0.228428f
C6520 7b_counter_0.MDFF_4.LD.t67 VSS 0.251201f
C6521 7b_counter_0.MDFF_4.LD.n7 VSS 0.106993f
C6522 7b_counter_0.MDFF_4.LD.t8 VSS 0.168722f
C6523 7b_counter_0.MDFF_4.LD.n8 VSS 0.112096f
C6524 7b_counter_0.MDFF_4.LD.t96 VSS 0.079924f
C6525 7b_counter_0.MDFF_4.LD.n9 VSS 0.0707f
C6526 7b_counter_0.MDFF_4.LD.n10 VSS 0.067288f
C6527 7b_counter_0.MDFF_4.LD.t113 VSS 0.062925f
C6528 7b_counter_0.MDFF_4.LD.t53 VSS 0.071805f
C6529 7b_counter_0.MDFF_4.LD.t70 VSS 0.228428f
C6530 7b_counter_0.MDFF_4.LD.t116 VSS 0.239085f
C6531 7b_counter_0.MDFF_4.LD.t85 VSS 0.117907f
C6532 7b_counter_0.MDFF_4.LD.n11 VSS 0.215352f
C6533 7b_counter_0.MDFF_4.LD.t109 VSS 0.168722f
C6534 7b_counter_0.MDFF_4.LD.n12 VSS 0.112096f
C6535 7b_counter_0.MDFF_4.LD.t106 VSS 0.079924f
C6536 7b_counter_0.MDFF_4.LD.n13 VSS 0.0707f
C6537 7b_counter_0.MDFF_4.LD.t49 VSS 0.080178f
C6538 7b_counter_0.MDFF_4.LD.t87 VSS 0.080178f
C6539 7b_counter_0.MDFF_4.LD.n14 VSS 0.102651f
C6540 7b_counter_0.MDFF_4.LD.t54 VSS 0.080178f
C6541 7b_counter_0.MDFF_4.LD.t112 VSS 0.080178f
C6542 7b_counter_0.MDFF_4.LD.n15 VSS 0.11396f
C6543 7b_counter_0.MDFF_4.LD.t15 VSS 0.080178f
C6544 7b_counter_0.MDFF_4.LD.n16 VSS 0.102651f
C6545 7b_counter_0.MDFF_4.LD.t44 VSS 0.102253f
C6546 7b_counter_0.MDFF_4.LD.n17 VSS 0.067288f
C6547 7b_counter_0.MDFF_4.LD.t10 VSS 0.062925f
C6548 7b_counter_0.MDFF_4.LD.t68 VSS 0.228428f
C6549 7b_counter_0.MDFF_4.LD.t31 VSS 0.251454f
C6550 7b_counter_0.MDFF_4.LD.t118 VSS 0.121066f
C6551 7b_counter_0.MDFF_4.LD.t81 VSS 0.078867f
C6552 7b_counter_0.MDFF_4.LD.n18 VSS 0.097903f
C6553 7b_counter_0.MDFF_4.LD.n19 VSS 0.107248f
C6554 7b_counter_0.MDFF_4.LD.t24 VSS 0.168722f
C6555 7b_counter_0.MDFF_4.LD.n20 VSS 0.112096f
C6556 7b_counter_0.MDFF_4.LD.t105 VSS 0.079924f
C6557 7b_counter_0.MDFF_4.LD.n21 VSS 0.0707f
C6558 7b_counter_0.MDFF_4.LD.t77 VSS 0.080178f
C6559 7b_counter_0.MDFF_4.LD.t66 VSS 0.080178f
C6560 7b_counter_0.MDFF_4.LD.n22 VSS 0.102651f
C6561 7b_counter_0.MDFF_4.LD.t71 VSS 0.080178f
C6562 7b_counter_0.MDFF_4.LD.t88 VSS 0.080178f
C6563 7b_counter_0.MDFF_4.LD.n23 VSS 0.11396f
C6564 7b_counter_0.MDFF_4.LD.t117 VSS 0.080178f
C6565 7b_counter_0.MDFF_4.LD.n24 VSS 0.102651f
C6566 7b_counter_0.MDFF_4.LD.t43 VSS 0.102253f
C6567 7b_counter_0.MDFF_4.LD.n25 VSS 0.067288f
C6568 7b_counter_0.MDFF_4.LD.t41 VSS 0.080178f
C6569 7b_counter_0.MDFF_4.LD.t13 VSS 0.080178f
C6570 7b_counter_0.MDFF_4.LD.n26 VSS 0.102651f
C6571 7b_counter_0.MDFF_4.LD.t80 VSS 0.080178f
C6572 7b_counter_0.MDFF_4.LD.t58 VSS 0.080178f
C6573 7b_counter_0.MDFF_4.LD.n27 VSS 0.11396f
C6574 7b_counter_0.MDFF_4.LD.t83 VSS 0.080178f
C6575 7b_counter_0.MDFF_4.LD.n28 VSS 0.102651f
C6576 7b_counter_0.MDFF_4.LD.t61 VSS 0.102253f
C6577 7b_counter_0.MDFF_4.LD.t9 VSS 0.062925f
C6578 7b_counter_0.MDFF_4.LD.t115 VSS 0.121087f
C6579 7b_counter_0.MDFF_4.LD.t94 VSS 0.079119f
C6580 7b_counter_0.MDFF_4.LD.n29 VSS 0.098138f
C6581 7b_counter_0.MDFF_4.LD.t34 VSS 0.228428f
C6582 7b_counter_0.MDFF_4.LD.t59 VSS 0.251201f
C6583 7b_counter_0.MDFF_4.LD.n30 VSS 0.106993f
C6584 7b_counter_0.MDFF_4.LD.t92 VSS 0.168734f
C6585 7b_counter_0.MDFF_4.LD.n31 VSS 0.112096f
C6586 7b_counter_0.MDFF_4.LD.t21 VSS 0.079924f
C6587 7b_counter_0.MDFF_4.LD.n32 VSS 0.0707f
C6588 7b_counter_0.MDFF_4.LD.n33 VSS 0.067288f
C6589 7b_counter_0.MDFF_4.LD.t42 VSS 0.080178f
C6590 7b_counter_0.MDFF_4.LD.t14 VSS 0.080178f
C6591 7b_counter_0.MDFF_4.LD.n34 VSS 0.102651f
C6592 7b_counter_0.MDFF_4.LD.t52 VSS 0.080178f
C6593 7b_counter_0.MDFF_4.LD.t26 VSS 0.080178f
C6594 7b_counter_0.MDFF_4.LD.n35 VSS 0.11396f
C6595 7b_counter_0.MDFF_4.LD.t84 VSS 0.080178f
C6596 7b_counter_0.MDFF_4.LD.n36 VSS 0.102651f
C6597 7b_counter_0.MDFF_4.LD.t62 VSS 0.102253f
C6598 7b_counter_0.MDFF_4.LD.t102 VSS 0.062925f
C6599 7b_counter_0.MDFF_4.LD.t97 VSS 0.120965f
C6600 7b_counter_0.MDFF_4.LD.t95 VSS 0.079119f
C6601 7b_counter_0.MDFF_4.LD.n37 VSS 0.09826f
C6602 7b_counter_0.MDFF_4.LD.t16 VSS 0.228428f
C6603 7b_counter_0.MDFF_4.LD.t60 VSS 0.251201f
C6604 7b_counter_0.MDFF_4.LD.n38 VSS 0.106993f
C6605 7b_counter_0.MDFF_4.LD.t93 VSS 0.168734f
C6606 7b_counter_0.MDFF_4.LD.n39 VSS 0.112096f
C6607 7b_counter_0.MDFF_4.LD.t23 VSS 0.079924f
C6608 7b_counter_0.MDFF_4.LD.n40 VSS 0.0707f
C6609 7b_counter_0.MDFF_4.LD.n41 VSS 0.067288f
C6610 7b_counter_0.MDFF_4.LD.t110 VSS 0.062925f
C6611 7b_counter_0.MDFF_4.LD.t89 VSS 0.228428f
C6612 7b_counter_0.MDFF_4.LD.t17 VSS 0.251454f
C6613 7b_counter_0.MDFF_4.LD.t64 VSS 0.079336f
C6614 7b_counter_0.MDFF_4.LD.t69 VSS 0.114389f
C6615 7b_counter_0.MDFF_4.LD.n42 VSS 0.102073f
C6616 7b_counter_0.MDFF_4.LD.n43 VSS 0.109269f
C6617 7b_counter_0.MDFF_4.LD.t103 VSS 0.168734f
C6618 7b_counter_0.MDFF_4.LD.n44 VSS 0.112096f
C6619 7b_counter_0.MDFF_4.LD.t32 VSS 0.079924f
C6620 7b_counter_0.MDFF_4.LD.n45 VSS 0.0707f
C6621 7b_counter_0.MDFF_4.LD.t37 VSS 0.080178f
C6622 7b_counter_0.MDFF_4.LD.t73 VSS 0.080178f
C6623 7b_counter_0.MDFF_4.LD.n46 VSS 0.102651f
C6624 7b_counter_0.MDFF_4.LD.t50 VSS 0.080178f
C6625 7b_counter_0.MDFF_4.LD.t56 VSS 0.080178f
C6626 7b_counter_0.MDFF_4.LD.n47 VSS 0.11396f
C6627 7b_counter_0.MDFF_4.LD.t29 VSS 0.080178f
C6628 7b_counter_0.MDFF_4.LD.n48 VSS 0.102651f
C6629 7b_counter_0.MDFF_4.LD.t82 VSS 0.102253f
C6630 7b_counter_0.MDFF_4.LD.n49 VSS 0.067288f
C6631 7b_counter_0.MDFF_4.LD.t65 VSS 0.080178f
C6632 7b_counter_0.MDFF_4.LD.t38 VSS 0.080178f
C6633 7b_counter_0.MDFF_4.LD.n50 VSS 0.102651f
C6634 7b_counter_0.MDFF_4.LD.t51 VSS 0.080178f
C6635 7b_counter_0.MDFF_4.LD.t25 VSS 0.080178f
C6636 7b_counter_0.MDFF_4.LD.n51 VSS 0.11396f
C6637 7b_counter_0.MDFF_4.LD.t40 VSS 0.080178f
C6638 7b_counter_0.MDFF_4.LD.n52 VSS 0.102651f
C6639 7b_counter_0.MDFF_4.LD.t12 VSS 0.102253f
C6640 7b_counter_0.MDFF_4.LD.t100 VSS 0.062925f
C6641 7b_counter_0.MDFF_4.LD.t18 VSS 0.121066f
C6642 7b_counter_0.MDFF_4.LD.t122 VSS 0.079119f
C6643 7b_counter_0.MDFF_4.LD.n53 VSS 0.098158f
C6644 7b_counter_0.MDFF_4.LD.t99 VSS 0.228428f
C6645 7b_counter_0.MDFF_4.LD.t86 VSS 0.251201f
C6646 7b_counter_0.MDFF_4.LD.n54 VSS 0.106993f
C6647 7b_counter_0.MDFF_4.LD.t119 VSS 0.168722f
C6648 7b_counter_0.MDFF_4.LD.n55 VSS 0.112096f
C6649 7b_counter_0.MDFF_4.LD.t91 VSS 0.079924f
C6650 7b_counter_0.MDFF_4.LD.n56 VSS 0.0707f
C6651 7b_counter_0.MDFF_4.LD.n57 VSS 0.067288f
C6652 7b_counter_0.MDFF_4.LD.t48 VSS 0.080178f
C6653 7b_counter_0.MDFF_4.LD.t20 VSS 0.080178f
C6654 7b_counter_0.MDFF_4.LD.n58 VSS 0.102651f
C6655 7b_counter_0.MDFF_4.LD.t78 VSS 0.080178f
C6656 7b_counter_0.MDFF_4.LD.t55 VSS 0.080178f
C6657 7b_counter_0.MDFF_4.LD.n59 VSS 0.11396f
C6658 7b_counter_0.MDFF_4.LD.t39 VSS 0.080178f
C6659 7b_counter_0.MDFF_4.LD.n60 VSS 0.102651f
C6660 7b_counter_0.MDFF_4.LD.t11 VSS 0.102253f
C6661 7b_counter_0.MDFF_4.LD.t7 VSS 0.062925f
C6662 7b_counter_0.MDFF_4.LD.t27 VSS 0.121066f
C6663 7b_counter_0.MDFF_4.LD.t104 VSS 0.079119f
C6664 7b_counter_0.MDFF_4.LD.n61 VSS 0.098158f
C6665 7b_counter_0.MDFF_4.LD.t75 VSS 0.228428f
C6666 7b_counter_0.MDFF_4.LD.t63 VSS 0.251201f
C6667 7b_counter_0.MDFF_4.LD.n62 VSS 0.106993f
C6668 7b_counter_0.MDFF_4.LD.t98 VSS 0.168722f
C6669 7b_counter_0.MDFF_4.LD.n63 VSS 0.112096f
C6670 7b_counter_0.MDFF_4.LD.t90 VSS 0.079924f
C6671 7b_counter_0.MDFF_4.LD.n64 VSS 0.0707f
C6672 7b_counter_0.MDFF_4.LD.n65 VSS 0.067288f
C6673 7b_counter_0.MDFF_4.LD.t22 VSS 0.062925f
C6674 7b_counter_0.MDFF_4.LD.t35 VSS 0.228428f
C6675 7b_counter_0.MDFF_4.LD.t28 VSS 0.251454f
C6676 7b_counter_0.MDFF_4.LD.t114 VSS 0.1227f
C6677 7b_counter_0.MDFF_4.LD.t74 VSS 0.078867f
C6678 7b_counter_0.MDFF_4.LD.n66 VSS 0.096256f
C6679 7b_counter_0.MDFF_4.LD.n67 VSS 0.107248f
C6680 7b_counter_0.MDFF_4.LD.t107 VSS 0.168722f
C6681 7b_counter_0.MDFF_4.LD.n68 VSS 0.112096f
C6682 7b_counter_0.MDFF_4.LD.t101 VSS 0.079924f
C6683 7b_counter_0.MDFF_4.LD.n69 VSS 0.0707f
C6684 7b_counter_0.MDFF_4.LD.t47 VSS 0.080178f
C6685 7b_counter_0.MDFF_4.LD.t6 VSS 0.080178f
C6686 7b_counter_0.MDFF_4.LD.n70 VSS 0.102651f
C6687 7b_counter_0.MDFF_4.LD.t76 VSS 0.080178f
C6688 7b_counter_0.MDFF_4.LD.t120 VSS 0.080178f
C6689 7b_counter_0.MDFF_4.LD.n71 VSS 0.11396f
C6690 7b_counter_0.MDFF_4.LD.t33 VSS 0.080178f
C6691 7b_counter_0.MDFF_4.LD.n72 VSS 0.102651f
C6692 7b_counter_0.MDFF_4.LD.t36 VSS 0.102253f
C6693 7b_counter_0.MDFF_4.LD.n73 VSS 0.067288f
C6694 7b_counter_0.MDFF_4.LD.t5 VSS 0.065111f
C6695 7b_counter_0.MDFF_4.LD.t1 VSS 0.069414f
C6696 7b_counter_0.MDFF_4.LD.t2 VSS 0.065111f
C6697 p3_gen_magic_0.P3.n0 VSS 0.22863f
C6698 p3_gen_magic_0.P3.t11 VSS 0.099501f
C6699 p3_gen_magic_0.P3.t15 VSS 0.108513f
C6700 p3_gen_magic_0.P3.t8 VSS 0.091976f
C6701 p3_gen_magic_0.P3.t9 VSS 0.04724f
C6702 p3_gen_magic_0.P3.t10 VSS 0.091976f
C6703 p3_gen_magic_0.P3.n1 VSS 0.072195f
C6704 p3_gen_magic_0.P3.n2 VSS 0.072195f
C6705 p3_gen_magic_0.P3.t14 VSS 0.07356f
C6706 p3_gen_magic_0.P3.n3 VSS 0.099762f
C6707 p3_gen_magic_0.P3.t12 VSS 0.102875f
C6708 p3_gen_magic_0.P3.t16 VSS 0.194954f
C6709 p3_gen_magic_0.P3.t7 VSS 0.205622f
C6710 p3_gen_magic_0.P3.t13 VSS 0.136197f
C6711 p3_gen_magic_0.P3.t6 VSS 0.065717f
C6712 p3_gen_magic_0.P3.n4 VSS 0.080641f
C6713 p3_gen_magic_0.P3.t5 VSS 0.01981f
C6714 p3_gen_magic_0.P3.t4 VSS 0.01981f
C6715 p3_gen_magic_0.P3.n5 VSS 0.044646f
C6716 p3_gen_magic_0.P3.t1 VSS 0.01981f
C6717 p3_gen_magic_0.P3.t0 VSS 0.01981f
C6718 p3_gen_magic_0.P3.n6 VSS 0.050042f
C6719 p3_gen_magic_0.P3.t3 VSS 0.01981f
C6720 p3_gen_magic_0.P3.t2 VSS 0.01981f
C6721 p3_gen_magic_0.P3.n7 VSS 0.042711f
C6722 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t0 VSS 0.03568f
C6723 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t2 VSS 0.041547f
C6724 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t1 VSS 0.032468f
C6725 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t4 VSS 0.031378f
C6726 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t5 VSS 0.062959f
C6727 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n0 VSS 0.066836f
C6728 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t12 VSS 0.080221f
C6729 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t8 VSS 0.04025f
C6730 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n1 VSS 0.097307f
C6731 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t6 VSS 0.11575f
C6732 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t11 VSS 0.058745f
C6733 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t10 VSS 0.038843f
C6734 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n2 VSS 0.102925f
C6735 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n3 VSS 0.147326f
C6736 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t9 VSS 0.073661f
C6737 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n4 VSS 0.264336f
C6738 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t3 VSS 0.031378f
C6739 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.t7 VSS 0.062482f
C6740 7b_counter_0.MDFF_7.tspc2_magic_0.CLK.n5 VSS 0.061863f
C6741 Q1.t1 VSS 0.018759f
C6742 Q1.t2 VSS 0.021844f
C6743 Q1.t0 VSS 0.017071f
C6744 Q1.n0 VSS 0.043928f
C6745 Q1.n1 VSS 0.033615f
C6746 Q1.n2 VSS 0.01076f
C6747 Q1.t21 VSS 0.02281f
C6748 Q1.t9 VSS 0.036588f
C6749 Q1.t7 VSS 0.059737f
C6750 Q1.t27 VSS 0.064394f
C6751 Q1.t11 VSS 0.064394f
C6752 Q1.t4 VSS 0.064394f
C6753 Q1.t18 VSS 0.04783f
C6754 Q1.n3 VSS 0.029276f
C6755 Q1.t13 VSS 0.016498f
C6756 Q1.t26 VSS 0.031344f
C6757 Q1.t8 VSS 0.020888f
C6758 Q1.n4 VSS 0.039018f
C6759 Q1.t16 VSS 0.039521f
C6760 Q1.n5 VSS 0.026825f
C6761 Q1.n6 VSS 0.368111f
C6762 Q1.t19 VSS 0.035352f
C6763 Q1.t25 VSS 0.042337f
C6764 Q1.t31 VSS 0.022731f
C6765 Q1.n7 VSS 0.029305f
C6766 Q1.t3 VSS 0.016498f
C6767 Q1.t20 VSS 0.032121f
C6768 Q1.n8 VSS 0.025213f
C6769 Q1.t17 VSS 0.032121f
C6770 Q1.n9 VSS 0.025213f
C6771 Q1.t12 VSS 0.025689f
C6772 Q1.t15 VSS 0.034749f
C6773 Q1.t24 VSS 0.037896f
C6774 Q1.n10 VSS 0.034831f
C6775 Q1.n11 VSS 0.38736f
C6776 Q1.n12 VSS 0.447139f
C6777 Q1.t14 VSS 0.016498f
C6778 Q1.t30 VSS 0.032121f
C6779 Q1.n13 VSS 0.025213f
C6780 Q1.t29 VSS 0.032121f
C6781 Q1.n14 VSS 0.025213f
C6782 Q1.t22 VSS 0.025689f
C6783 Q1.t23 VSS 0.034749f
C6784 Q1.t5 VSS 0.037896f
C6785 Q1.n15 VSS 0.034831f
C6786 Q1.t28 VSS 0.035352f
C6787 Q1.t6 VSS 0.042337f
C6788 Q1.t10 VSS 0.022731f
C6789 Q1.n16 VSS 0.029305f
C6790 Q1.n17 VSS 0.095281f
C6791 Q1.n18 VSS 0.022344f
C6792 Q1.n19 VSS 1.51738f
C6793 Q1.n20 VSS 1.73202f
C6794 Q1.n21 VSS 0.107991f
C6795 DFF_magic_0.D.t5 VSS 0.039468f
C6796 DFF_magic_0.D.t0 VSS 0.053011f
C6797 DFF_magic_0.D.t1 VSS 0.014233f
C6798 DFF_magic_0.D.t2 VSS 0.014233f
C6799 DFF_magic_0.D.n0 VSS 0.028466f
C6800 DFF_magic_0.D.n1 VSS 0.122135f
C6801 DFF_magic_0.D.t3 VSS 0.014233f
C6802 DFF_magic_0.D.t4 VSS 0.014233f
C6803 DFF_magic_0.D.n2 VSS 0.028466f
C6804 DFF_magic_0.D.n3 VSS 0.061014f
C6805 DFF_magic_0.D.t36 VSS 0.079061f
C6806 DFF_magic_0.D.t20 VSS 0.076502f
C6807 DFF_magic_0.D.t21 VSS 0.126317f
C6808 DFF_magic_0.D.t35 VSS 0.08047f
C6809 DFF_magic_0.D.n4 VSS 0.056677f
C6810 DFF_magic_0.D.t32 VSS 0.111468f
C6811 DFF_magic_0.D.t19 VSS 0.126317f
C6812 DFF_magic_0.D.t18 VSS 0.108641f
C6813 DFF_magic_0.D.n5 VSS 0.058813f
C6814 DFF_magic_0.D.t22 VSS 0.108641f
C6815 DFF_magic_0.D.t23 VSS 0.089867f
C6816 DFF_magic_0.D.n6 VSS 0.127285f
C6817 DFF_magic_0.D.n7 VSS 2.05474f
C6818 DFF_magic_0.D.t28 VSS 0.079061f
C6819 DFF_magic_0.D.t33 VSS 0.076502f
C6820 DFF_magic_0.D.t34 VSS 0.126317f
C6821 DFF_magic_0.D.t17 VSS 0.08047f
C6822 DFF_magic_0.D.n8 VSS 0.056677f
C6823 DFF_magic_0.D.t16 VSS 0.111468f
C6824 DFF_magic_0.D.t31 VSS 0.126317f
C6825 DFF_magic_0.D.t30 VSS 0.108641f
C6826 DFF_magic_0.D.n9 VSS 0.058813f
C6827 DFF_magic_0.D.t12 VSS 0.108641f
C6828 DFF_magic_0.D.t13 VSS 0.089867f
C6829 DFF_magic_0.D.n10 VSS 0.122705f
C6830 DFF_magic_0.D.n11 VSS 0.351771f
C6831 DFF_magic_0.D.t38 VSS 0.079061f
C6832 DFF_magic_0.D.t24 VSS 0.076502f
C6833 DFF_magic_0.D.t25 VSS 0.126317f
C6834 DFF_magic_0.D.t37 VSS 0.08047f
C6835 DFF_magic_0.D.n12 VSS 0.056677f
C6836 DFF_magic_0.D.t29 VSS 0.111468f
C6837 DFF_magic_0.D.t15 VSS 0.126317f
C6838 DFF_magic_0.D.t14 VSS 0.108641f
C6839 DFF_magic_0.D.n13 VSS 0.058813f
C6840 DFF_magic_0.D.t26 VSS 0.108641f
C6841 DFF_magic_0.D.t27 VSS 0.089867f
C6842 DFF_magic_0.D.n14 VSS 0.111313f
C6843 DFF_magic_0.D.n15 VSS 0.346143f
C6844 DFF_magic_0.D.t8 VSS 0.014233f
C6845 DFF_magic_0.D.t7 VSS 0.014233f
C6846 DFF_magic_0.D.n16 VSS 0.030686f
C6847 DFF_magic_0.D.t10 VSS 0.014233f
C6848 DFF_magic_0.D.t11 VSS 0.014233f
C6849 DFF_magic_0.D.n17 VSS 0.032076f
C6850 DFF_magic_0.D.t9 VSS 0.014233f
C6851 DFF_magic_0.D.t6 VSS 0.014233f
C6852 DFF_magic_0.D.n18 VSS 0.035953f
C6853 7b_counter_0.NAND_magic_0.A.n0 VSS 1.09186f
C6854 7b_counter_0.NAND_magic_0.A.n1 VSS 0.292035f
C6855 7b_counter_0.NAND_magic_0.A.t17 VSS 0.060277f
C6856 7b_counter_0.NAND_magic_0.A.t14 VSS 0.117357f
C6857 7b_counter_0.NAND_magic_0.A.n2 VSS 0.092118f
C6858 7b_counter_0.NAND_magic_0.A.t18 VSS 0.117357f
C6859 7b_counter_0.NAND_magic_0.A.n3 VSS 0.092118f
C6860 7b_counter_0.NAND_magic_0.A.t6 VSS 0.09386f
C6861 7b_counter_0.NAND_magic_0.A.t21 VSS 0.12696f
C6862 7b_counter_0.NAND_magic_0.A.t9 VSS 0.138458f
C6863 7b_counter_0.NAND_magic_0.A.n4 VSS 0.127297f
C6864 7b_counter_0.NAND_magic_0.A.t19 VSS 0.110205f
C6865 7b_counter_0.NAND_magic_0.A.t16 VSS 0.0717f
C6866 7b_counter_0.NAND_magic_0.A.n5 VSS 0.090591f
C6867 7b_counter_0.NAND_magic_0.A.t13 VSS 0.113674f
C6868 7b_counter_0.NAND_magic_0.A.t11 VSS 0.073888f
C6869 7b_counter_0.NAND_magic_0.A.n6 VSS 0.088336f
C6870 7b_counter_0.NAND_magic_0.A.n7 VSS 0.033173f
C6871 7b_counter_0.NAND_magic_0.A.n8 VSS 1.4974f
C6872 7b_counter_0.NAND_magic_0.A.t15 VSS 0.12696f
C6873 7b_counter_0.NAND_magic_0.A.t12 VSS 0.138458f
C6874 7b_counter_0.NAND_magic_0.A.t20 VSS 0.117357f
C6875 7b_counter_0.NAND_magic_0.A.t8 VSS 0.060277f
C6876 7b_counter_0.NAND_magic_0.A.t10 VSS 0.117357f
C6877 7b_counter_0.NAND_magic_0.A.n9 VSS 0.092118f
C6878 7b_counter_0.NAND_magic_0.A.n10 VSS 0.092118f
C6879 7b_counter_0.NAND_magic_0.A.t7 VSS 0.09386f
C6880 7b_counter_0.NAND_magic_0.A.n11 VSS 0.127292f
C6881 7b_counter_0.NAND_magic_0.A.t5 VSS 0.025277f
C6882 7b_counter_0.NAND_magic_0.A.t4 VSS 0.025277f
C6883 7b_counter_0.NAND_magic_0.A.n12 VSS 0.056967f
C6884 7b_counter_0.NAND_magic_0.A.t1 VSS 0.025277f
C6885 7b_counter_0.NAND_magic_0.A.t0 VSS 0.025277f
C6886 7b_counter_0.NAND_magic_0.A.n13 VSS 0.063852f
C6887 7b_counter_0.NAND_magic_0.A.t3 VSS 0.025277f
C6888 7b_counter_0.NAND_magic_0.A.t2 VSS 0.025277f
C6889 7b_counter_0.NAND_magic_0.A.n14 VSS 0.054498f
C6890 mux_magic_0.IN2.t2 VSS 0.061795f
C6891 mux_magic_0.IN2.t0 VSS 0.048886f
C6892 mux_magic_0.IN2.t1 VSS 0.65564f
C6893 mux_magic_0.IN2.t12 VSS 0.034643f
C6894 mux_magic_0.IN2.t9 VSS 0.065817f
C6895 mux_magic_0.IN2.t4 VSS 0.043862f
C6896 mux_magic_0.IN2.n0 VSS 0.081932f
C6897 mux_magic_0.IN2.t8 VSS 0.082987f
C6898 mux_magic_0.IN2.n1 VSS 0.056329f
C6899 mux_magic_0.IN2.t6 VSS 0.072967f
C6900 mux_magic_0.IN2.t3 VSS 0.079575f
C6901 mux_magic_0.IN2.t7 VSS 0.067448f
C6902 mux_magic_0.IN2.t11 VSS 0.034643f
C6903 mux_magic_0.IN2.t5 VSS 0.067448f
C6904 mux_magic_0.IN2.n2 VSS 0.052943f
C6905 mux_magic_0.IN2.n3 VSS 0.052943f
C6906 mux_magic_0.IN2.t10 VSS 0.053944f
C6907 mux_magic_0.IN2.n4 VSS 0.073158f
C6908 D2_7.t23 VSS 0.02269f
C6909 D2_7.t22 VSS 0.043108f
C6910 D2_7.t0 VSS 0.028728f
C6911 D2_7.n0 VSS 0.053663f
C6912 D2_7.t15 VSS 0.054354f
C6913 D2_7.n1 VSS 0.036894f
C6914 D2_7.t20 VSS 0.02269f
C6915 D2_7.t24 VSS 0.043108f
C6916 D2_7.t1 VSS 0.028728f
C6917 D2_7.n2 VSS 0.053663f
C6918 D2_7.t13 VSS 0.054354f
C6919 D2_7.n3 VSS 0.036894f
C6920 D2_7.t19 VSS 0.030009f
C6921 D2_7.t16 VSS 0.048621f
C6922 D2_7.t4 VSS 0.059508f
C6923 D2_7.n4 VSS 0.042033f
C6924 D2_7.t2 VSS 0.047791f
C6925 D2_7.t12 VSS 0.052119f
C6926 D2_7.t9 VSS 0.02269f
C6927 D2_7.t6 VSS 0.044176f
C6928 D2_7.n5 VSS 0.034676f
C6929 D2_7.t3 VSS 0.044176f
C6930 D2_7.n6 VSS 0.034676f
C6931 D2_7.t21 VSS 0.035331f
C6932 D2_7.n7 VSS 0.047911f
C6933 D2_7.n8 VSS 0.909985f
C6934 D2_7.t8 VSS 0.047791f
C6935 D2_7.t18 VSS 0.052119f
C6936 D2_7.t17 VSS 0.02269f
C6937 D2_7.t14 VSS 0.044176f
C6938 D2_7.n9 VSS 0.034676f
C6939 D2_7.t11 VSS 0.044176f
C6940 D2_7.n10 VSS 0.034676f
C6941 D2_7.t7 VSS 0.035331f
C6942 D2_7.n11 VSS 0.047911f
C6943 D2_7.t5 VSS 0.030009f
C6944 D2_7.t25 VSS 0.048621f
C6945 D2_7.t10 VSS 0.059508f
C6946 D2_7.n12 VSS 0.042033f
C6947 D2_7.n13 VSS 0.372945f
C6948 D2_7.n14 VSS 2.08667f
C6949 D2_7.n15 VSS 2.31417f
C6950 D2_7.n16 VSS 0.286147f
C6951 LD.t24 VSS 0.083615f
C6952 LD.t84 VSS 0.083615f
C6953 LD.n0 VSS 0.107052f
C6954 LD.t49 VSS 0.083615f
C6955 LD.t30 VSS 0.083615f
C6956 LD.n1 VSS 0.118845f
C6957 LD.t80 VSS 0.083615f
C6958 LD.n2 VSS 0.107052f
C6959 LD.t38 VSS 0.106636f
C6960 LD.t82 VSS 0.065622f
C6961 LD.t33 VSS 0.126277f
C6962 LD.t59 VSS 0.082511f
C6963 LD.n3 VSS 0.102345f
C6964 LD.t55 VSS 0.23822f
C6965 LD.t26 VSS 0.26197f
C6966 LD.n4 VSS 0.11158f
C6967 LD.t60 VSS 0.175967f
C6968 LD.n5 VSS 0.116902f
C6969 LD.t10 VSS 0.083351f
C6970 LD.n6 VSS 0.073731f
C6971 LD.n7 VSS 0.070173f
C6972 LD.t6 VSS 0.067902f
C6973 LD.n8 VSS 0.148309f
C6974 LD.t0 VSS 0.072389f
C6975 LD.t7 VSS 0.027519f
C6976 LD.t8 VSS 0.027519f
C6977 LD.n9 VSS 0.055038f
C6978 LD.n10 VSS 0.149579f
C6979 LD.t3 VSS 0.027519f
C6980 LD.t5 VSS 0.027519f
C6981 LD.n11 VSS 0.055038f
C6982 LD.n12 VSS 0.09634f
C6983 LD.t2 VSS 0.027519f
C6984 LD.t4 VSS 0.027519f
C6985 LD.n13 VSS 0.054966f
C6986 LD.n14 VSS 0.124249f
C6987 LD.n15 VSS 0.144944f
C6988 LD.t1 VSS 0.067902f
C6989 LD.n16 VSS 0.090954f
C6990 LD.n17 VSS 4.35279f
C6991 LD.n18 VSS 5.29068f
C6992 LD.t64 VSS 0.065622f
C6993 LD.t54 VSS 0.23822f
C6994 LD.t23 VSS 0.262233f
C6995 LD.t39 VSS 0.126277f
C6996 LD.t63 VSS 0.082247f
C6997 LD.n19 VSS 0.102079f
C6998 LD.n20 VSS 0.111845f
C6999 LD.t41 VSS 0.175967f
C7000 LD.n21 VSS 0.116902f
C7001 LD.t9 VSS 0.083351f
C7002 LD.n22 VSS 0.073731f
C7003 LD.t74 VSS 0.083615f
C7004 LD.t13 VSS 0.083615f
C7005 LD.n23 VSS 0.107052f
C7006 LD.t19 VSS 0.083615f
C7007 LD.t57 VSS 0.083615f
C7008 LD.n24 VSS 0.118845f
C7009 LD.t44 VSS 0.083615f
C7010 LD.n25 VSS 0.107052f
C7011 LD.t52 VSS 0.106636f
C7012 LD.n26 VSS 0.070173f
C7013 LD.t73 VSS 0.065622f
C7014 LD.t27 VSS 0.23822f
C7015 LD.t86 VSS 0.262233f
C7016 LD.t15 VSS 0.126277f
C7017 LD.t47 VSS 0.082247f
C7018 LD.n27 VSS 0.102079f
C7019 LD.n28 VSS 0.111845f
C7020 LD.t51 VSS 0.175967f
C7021 LD.n29 VSS 0.116902f
C7022 LD.t75 VSS 0.083351f
C7023 LD.n30 VSS 0.073731f
C7024 LD.t53 VSS 0.077265f
C7025 LD.t29 VSS 0.077265f
C7026 LD.t65 VSS 0.077265f
C7027 LD.t83 VSS 0.077265f
C7028 LD.t77 VSS 0.077265f
C7029 LD.n31 VSS 0.119753f
C7030 LD.n32 VSS 0.131546f
C7031 LD.n33 VSS 0.119753f
C7032 LD.t37 VSS 0.100285f
C7033 LD.n34 VSS 0.070173f
C7034 LD.n35 VSS 1.0159f
C7035 LD.t85 VSS 0.083615f
C7036 LD.t68 VSS 0.083615f
C7037 LD.n36 VSS 0.107052f
C7038 LD.t31 VSS 0.083615f
C7039 LD.t11 VSS 0.083615f
C7040 LD.n37 VSS 0.118845f
C7041 LD.t40 VSS 0.083615f
C7042 LD.n38 VSS 0.107052f
C7043 LD.t17 VSS 0.106636f
C7044 LD.t67 VSS 0.065622f
C7045 LD.t36 VSS 0.126277f
C7046 LD.t61 VSS 0.082511f
C7047 LD.n39 VSS 0.102345f
C7048 LD.t58 VSS 0.23822f
C7049 LD.t34 VSS 0.26197f
C7050 LD.n40 VSS 0.11158f
C7051 LD.t46 VSS 0.175967f
C7052 LD.n41 VSS 0.116902f
C7053 LD.t72 VSS 0.083351f
C7054 LD.n42 VSS 0.073731f
C7055 LD.n43 VSS 0.070173f
C7056 LD.n44 VSS 0.370414f
C7057 LD.t56 VSS 0.065622f
C7058 LD.t50 VSS 0.23822f
C7059 LD.t18 VSS 0.262233f
C7060 LD.t35 VSS 0.126277f
C7061 LD.t62 VSS 0.082247f
C7062 LD.n45 VSS 0.102079f
C7063 LD.n46 VSS 0.111845f
C7064 LD.t32 VSS 0.175967f
C7065 LD.n47 VSS 0.116902f
C7066 LD.t81 VSS 0.083351f
C7067 LD.n48 VSS 0.073731f
C7068 LD.t70 VSS 0.083615f
C7069 LD.t69 VSS 0.083615f
C7070 LD.n49 VSS 0.107052f
C7071 LD.t16 VSS 0.083615f
C7072 LD.t12 VSS 0.083615f
C7073 LD.n50 VSS 0.118845f
C7074 LD.t42 VSS 0.083615f
C7075 LD.n51 VSS 0.107052f
C7076 LD.t48 VSS 0.106636f
C7077 LD.n52 VSS 0.070173f
C7078 LD.n53 VSS 0.961681f
C7079 LD.t66 VSS 0.065622f
C7080 LD.t21 VSS 0.23822f
C7081 LD.t79 VSS 0.262233f
C7082 LD.t14 VSS 0.126277f
C7083 LD.t43 VSS 0.082247f
C7084 LD.n54 VSS 0.102079f
C7085 LD.n55 VSS 0.111845f
C7086 LD.t45 VSS 0.175967f
C7087 LD.n56 VSS 0.116902f
C7088 LD.t71 VSS 0.083351f
C7089 LD.n57 VSS 0.073731f
C7090 LD.t25 VSS 0.077265f
C7091 LD.t22 VSS 0.077265f
C7092 LD.t20 VSS 0.077265f
C7093 LD.t78 VSS 0.077265f
C7094 LD.t76 VSS 0.077265f
C7095 LD.n58 VSS 0.119753f
C7096 LD.n59 VSS 0.131546f
C7097 LD.n60 VSS 0.119753f
C7098 LD.t28 VSS 0.100285f
C7099 LD.n61 VSS 0.070173f
C7100 LD.n62 VSS 0.24105f
C7101 D2_2.t11 VSS 0.0311f
C7102 D2_2.t19 VSS 0.059086f
C7103 D2_2.t21 VSS 0.039376f
C7104 D2_2.n0 VSS 0.073553f
C7105 D2_2.t12 VSS 0.0745f
C7106 D2_2.n1 VSS 0.050568f
C7107 D2_2.t13 VSS 0.0311f
C7108 D2_2.t5 VSS 0.06055f
C7109 D2_2.n2 VSS 0.047528f
C7110 D2_2.t7 VSS 0.06055f
C7111 D2_2.n3 VSS 0.047528f
C7112 D2_2.t24 VSS 0.048427f
C7113 D2_2.t23 VSS 0.065504f
C7114 D2_2.t8 VSS 0.071437f
C7115 D2_2.n4 VSS 0.065669f
C7116 D2_2.t20 VSS 0.066642f
C7117 D2_2.t25 VSS 0.081565f
C7118 D2_2.t4 VSS 0.041132f
C7119 D2_2.n5 VSS 0.057612f
C7120 D2_2.n6 VSS 0.442514f
C7121 D2_2.t22 VSS 0.0311f
C7122 D2_2.t15 VSS 0.06055f
C7123 D2_2.n7 VSS 0.047528f
C7124 D2_2.t18 VSS 0.06055f
C7125 D2_2.n8 VSS 0.047528f
C7126 D2_2.t6 VSS 0.048427f
C7127 D2_2.t3 VSS 0.065504f
C7128 D2_2.t16 VSS 0.071437f
C7129 D2_2.n9 VSS 0.065669f
C7130 D2_2.t1 VSS 0.066642f
C7131 D2_2.t9 VSS 0.081565f
C7132 D2_2.t14 VSS 0.041132f
C7133 D2_2.n10 VSS 0.057612f
C7134 D2_2.n11 VSS 0.09276f
C7135 D2_2.n12 VSS 1.64633f
C7136 D2_2.n13 VSS 1.73802f
C7137 D2_2.n14 VSS 0.073141f
C7138 D2_2.t0 VSS 0.0311f
C7139 D2_2.t10 VSS 0.059086f
C7140 D2_2.t17 VSS 0.039376f
C7141 D2_2.n15 VSS 0.073553f
C7142 D2_2.t2 VSS 0.0745f
C7143 D2_2.n16 VSS 0.050568f
C7144 7b_counter_0.MDFF_5.LD.n0 VSS 0.146141f
C7145 7b_counter_0.MDFF_5.LD.n1 VSS 3.28018f
C7146 7b_counter_0.MDFF_5.LD.n2 VSS 3.28401f
C7147 7b_counter_0.MDFF_5.LD.n3 VSS 0.978211f
C7148 7b_counter_0.MDFF_5.LD.t33 VSS 0.064662f
C7149 7b_counter_0.MDFF_5.LD.t72 VSS 0.234736f
C7150 7b_counter_0.MDFF_5.LD.t68 VSS 0.258399f
C7151 7b_counter_0.MDFF_5.LD.t41 VSS 0.12441f
C7152 7b_counter_0.MDFF_5.LD.t19 VSS 0.081045f
C7153 7b_counter_0.MDFF_5.LD.n4 VSS 0.100607f
C7154 7b_counter_0.MDFF_5.LD.n5 VSS 0.11021f
C7155 7b_counter_0.MDFF_5.LD.t13 VSS 0.173381f
C7156 7b_counter_0.MDFF_5.LD.n6 VSS 0.115192f
C7157 7b_counter_0.MDFF_5.LD.t10 VSS 0.082132f
C7158 7b_counter_0.MDFF_5.LD.n7 VSS 0.072652f
C7159 7b_counter_0.MDFF_5.LD.t51 VSS 0.082392f
C7160 7b_counter_0.MDFF_5.LD.t44 VSS 0.082392f
C7161 7b_counter_0.MDFF_5.LD.n8 VSS 0.105486f
C7162 7b_counter_0.MDFF_5.LD.t75 VSS 0.082392f
C7163 7b_counter_0.MDFF_5.LD.t73 VSS 0.082392f
C7164 7b_counter_0.MDFF_5.LD.n9 VSS 0.117108f
C7165 7b_counter_0.MDFF_5.LD.t39 VSS 0.082392f
C7166 7b_counter_0.MDFF_5.LD.n10 VSS 0.105486f
C7167 7b_counter_0.MDFF_5.LD.t45 VSS 0.105076f
C7168 7b_counter_0.MDFF_5.LD.n11 VSS 0.069147f
C7169 7b_counter_0.MDFF_5.LD.t50 VSS 0.082392f
C7170 7b_counter_0.MDFF_5.LD.t62 VSS 0.082392f
C7171 7b_counter_0.MDFF_5.LD.n12 VSS 0.105486f
C7172 7b_counter_0.MDFF_5.LD.t86 VSS 0.082392f
C7173 7b_counter_0.MDFF_5.LD.t78 VSS 0.082392f
C7174 7b_counter_0.MDFF_5.LD.n13 VSS 0.117108f
C7175 7b_counter_0.MDFF_5.LD.t71 VSS 0.082392f
C7176 7b_counter_0.MDFF_5.LD.n14 VSS 0.105486f
C7177 7b_counter_0.MDFF_5.LD.t55 VSS 0.105076f
C7178 7b_counter_0.MDFF_5.LD.t52 VSS 0.064662f
C7179 7b_counter_0.MDFF_5.LD.t69 VSS 0.12441f
C7180 7b_counter_0.MDFF_5.LD.t36 VSS 0.081304f
C7181 7b_counter_0.MDFF_5.LD.n15 VSS 0.100869f
C7182 7b_counter_0.MDFF_5.LD.t17 VSS 0.234736f
C7183 7b_counter_0.MDFF_5.LD.t11 VSS 0.258139f
C7184 7b_counter_0.MDFF_5.LD.n16 VSS 0.109948f
C7185 7b_counter_0.MDFF_5.LD.t26 VSS 0.173381f
C7186 7b_counter_0.MDFF_5.LD.n17 VSS 0.115192f
C7187 7b_counter_0.MDFF_5.LD.t22 VSS 0.082132f
C7188 7b_counter_0.MDFF_5.LD.n18 VSS 0.072652f
C7189 7b_counter_0.MDFF_5.LD.n19 VSS 0.069147f
C7190 7b_counter_0.MDFF_5.LD.t14 VSS 0.064662f
C7191 7b_counter_0.MDFF_5.LD.t21 VSS 0.234736f
C7192 7b_counter_0.MDFF_5.LD.t61 VSS 0.258399f
C7193 7b_counter_0.MDFF_5.LD.t16 VSS 0.124431f
C7194 7b_counter_0.MDFF_5.LD.t15 VSS 0.081045f
C7195 7b_counter_0.MDFF_5.LD.n20 VSS 0.100586f
C7196 7b_counter_0.MDFF_5.LD.n21 VSS 0.11021f
C7197 7b_counter_0.MDFF_5.LD.t12 VSS 0.173394f
C7198 7b_counter_0.MDFF_5.LD.n22 VSS 0.115192f
C7199 7b_counter_0.MDFF_5.LD.t37 VSS 0.082132f
C7200 7b_counter_0.MDFF_5.LD.n23 VSS 0.072652f
C7201 7b_counter_0.MDFF_5.LD.t47 VSS 0.082392f
C7202 7b_counter_0.MDFF_5.LD.t40 VSS 0.082392f
C7203 7b_counter_0.MDFF_5.LD.n24 VSS 0.105486f
C7204 7b_counter_0.MDFF_5.LD.t53 VSS 0.082392f
C7205 7b_counter_0.MDFF_5.LD.t49 VSS 0.082392f
C7206 7b_counter_0.MDFF_5.LD.n25 VSS 0.117108f
C7207 7b_counter_0.MDFF_5.LD.t76 VSS 0.082392f
C7208 7b_counter_0.MDFF_5.LD.n26 VSS 0.105486f
C7209 7b_counter_0.MDFF_5.LD.t77 VSS 0.105076f
C7210 7b_counter_0.MDFF_5.LD.n27 VSS 0.069147f
C7211 7b_counter_0.MDFF_5.LD.t38 VSS 0.082392f
C7212 7b_counter_0.MDFF_5.LD.t58 VSS 0.082392f
C7213 7b_counter_0.MDFF_5.LD.n28 VSS 0.105486f
C7214 7b_counter_0.MDFF_5.LD.t81 VSS 0.082392f
C7215 7b_counter_0.MDFF_5.LD.t66 VSS 0.082392f
C7216 7b_counter_0.MDFF_5.LD.n29 VSS 0.117108f
C7217 7b_counter_0.MDFF_5.LD.t18 VSS 0.082392f
C7218 7b_counter_0.MDFF_5.LD.n30 VSS 0.105486f
C7219 7b_counter_0.MDFF_5.LD.t85 VSS 0.105076f
C7220 7b_counter_0.MDFF_5.LD.t30 VSS 0.064662f
C7221 7b_counter_0.MDFF_5.LD.t34 VSS 0.124305f
C7222 7b_counter_0.MDFF_5.LD.t32 VSS 0.081304f
C7223 7b_counter_0.MDFF_5.LD.n31 VSS 0.100973f
C7224 7b_counter_0.MDFF_5.LD.t60 VSS 0.234736f
C7225 7b_counter_0.MDFF_5.LD.t83 VSS 0.258139f
C7226 7b_counter_0.MDFF_5.LD.n32 VSS 0.109948f
C7227 7b_counter_0.MDFF_5.LD.t25 VSS 0.173394f
C7228 7b_counter_0.MDFF_5.LD.n33 VSS 0.115192f
C7229 7b_counter_0.MDFF_5.LD.t64 VSS 0.082132f
C7230 7b_counter_0.MDFF_5.LD.n34 VSS 0.072652f
C7231 7b_counter_0.MDFF_5.LD.n35 VSS 0.069147f
C7232 7b_counter_0.MDFF_5.LD.t27 VSS 0.082392f
C7233 7b_counter_0.MDFF_5.LD.t57 VSS 0.082392f
C7234 7b_counter_0.MDFF_5.LD.n36 VSS 0.105486f
C7235 7b_counter_0.MDFF_5.LD.t48 VSS 0.082392f
C7236 7b_counter_0.MDFF_5.LD.t80 VSS 0.082392f
C7237 7b_counter_0.MDFF_5.LD.n37 VSS 0.117108f
C7238 7b_counter_0.MDFF_5.LD.t9 VSS 0.082392f
C7239 7b_counter_0.MDFF_5.LD.n38 VSS 0.105486f
C7240 7b_counter_0.MDFF_5.LD.t84 VSS 0.105076f
C7241 7b_counter_0.MDFF_5.LD.t54 VSS 0.064662f
C7242 7b_counter_0.MDFF_5.LD.t43 VSS 0.124431f
C7243 7b_counter_0.MDFF_5.LD.t31 VSS 0.081304f
C7244 7b_counter_0.MDFF_5.LD.n39 VSS 0.100848f
C7245 7b_counter_0.MDFF_5.LD.t70 VSS 0.234736f
C7246 7b_counter_0.MDFF_5.LD.t82 VSS 0.258139f
C7247 7b_counter_0.MDFF_5.LD.n40 VSS 0.109948f
C7248 7b_counter_0.MDFF_5.LD.t24 VSS 0.173394f
C7249 7b_counter_0.MDFF_5.LD.n41 VSS 0.115192f
C7250 7b_counter_0.MDFF_5.LD.t63 VSS 0.082132f
C7251 7b_counter_0.MDFF_5.LD.n42 VSS 0.072652f
C7252 7b_counter_0.MDFF_5.LD.n43 VSS 0.069147f
C7253 7b_counter_0.MDFF_5.LD.t2 VSS 0.066909f
C7254 7b_counter_0.MDFF_5.LD.t6 VSS 0.027117f
C7255 7b_counter_0.MDFF_5.LD.t8 VSS 0.027117f
C7256 7b_counter_0.MDFF_5.LD.n44 VSS 0.054162f
C7257 7b_counter_0.MDFF_5.LD.t7 VSS 0.071331f
C7258 7b_counter_0.MDFF_5.LD.n45 VSS 0.142824f
C7259 7b_counter_0.MDFF_5.LD.n46 VSS 0.122432f
C7260 7b_counter_0.MDFF_5.LD.t1 VSS 0.027117f
C7261 7b_counter_0.MDFF_5.LD.t3 VSS 0.027117f
C7262 7b_counter_0.MDFF_5.LD.n47 VSS 0.054233f
C7263 7b_counter_0.MDFF_5.LD.n48 VSS 0.094931f
C7264 7b_counter_0.MDFF_5.LD.t4 VSS 0.027117f
C7265 7b_counter_0.MDFF_5.LD.t0 VSS 0.027117f
C7266 7b_counter_0.MDFF_5.LD.n49 VSS 0.054233f
C7267 7b_counter_0.MDFF_5.LD.n50 VSS 0.147391f
C7268 7b_counter_0.MDFF_5.LD.t5 VSS 0.066909f
C7269 7b_counter_0.MDFF_5.LD.t46 VSS 0.082392f
C7270 7b_counter_0.MDFF_5.LD.t74 VSS 0.082392f
C7271 7b_counter_0.MDFF_5.LD.n51 VSS 0.105486f
C7272 7b_counter_0.MDFF_5.LD.t35 VSS 0.082392f
C7273 7b_counter_0.MDFF_5.LD.t65 VSS 0.082392f
C7274 7b_counter_0.MDFF_5.LD.n52 VSS 0.117108f
C7275 7b_counter_0.MDFF_5.LD.t79 VSS 0.082392f
C7276 7b_counter_0.MDFF_5.LD.n53 VSS 0.105486f
C7277 7b_counter_0.MDFF_5.LD.t56 VSS 0.105076f
C7278 7b_counter_0.MDFF_5.LD.t29 VSS 0.064662f
C7279 7b_counter_0.MDFF_5.LD.t67 VSS 0.12441f
C7280 7b_counter_0.MDFF_5.LD.t59 VSS 0.081304f
C7281 7b_counter_0.MDFF_5.LD.n54 VSS 0.100869f
C7282 7b_counter_0.MDFF_5.LD.t28 VSS 0.234736f
C7283 7b_counter_0.MDFF_5.LD.t20 VSS 0.258139f
C7284 7b_counter_0.MDFF_5.LD.n55 VSS 0.109948f
C7285 7b_counter_0.MDFF_5.LD.t42 VSS 0.173381f
C7286 7b_counter_0.MDFF_5.LD.n56 VSS 0.115192f
C7287 7b_counter_0.MDFF_5.LD.t23 VSS 0.082132f
C7288 7b_counter_0.MDFF_5.LD.n57 VSS 0.072652f
C7289 7b_counter_0.MDFF_5.LD.n58 VSS 0.069147f
C7290 a_29512_8496.t3 VSS 0.085676f
C7291 a_29512_8496.n0 VSS 0.345476f
C7292 a_29512_8496.n1 VSS 0.409708f
C7293 a_29512_8496.t1 VSS 0.063303f
C7294 a_29512_8496.t0 VSS 0.067861f
C7295 a_29512_8496.t2 VSS 0.054881f
C7296 a_29512_8496.t14 VSS 0.122971f
C7297 a_29512_8496.t12 VSS 0.119549f
C7298 a_29512_8496.t13 VSS 0.197395f
C7299 a_29512_8496.t7 VSS 0.125751f
C7300 a_29512_8496.n2 VSS 0.089259f
C7301 a_29512_8496.t6 VSS 0.174488f
C7302 a_29512_8496.t11 VSS 0.197395f
C7303 a_29512_8496.t10 VSS 0.169773f
C7304 a_29512_8496.n3 VSS 0.091907f
C7305 a_29512_8496.t8 VSS 0.169773f
C7306 a_29512_8496.t9 VSS 0.141829f
C7307 a_29512_8496.n4 VSS 0.159639f
C7308 a_29512_8496.t5 VSS 0.054881f
C7309 a_29512_8496.t4 VSS 0.058483f
C7310 D2_1.t25 VSS 0.024214f
C7311 D2_1.t30 VSS 0.046004f
C7312 D2_1.t3 VSS 0.030658f
C7313 D2_1.n0 VSS 0.057268f
C7314 D2_1.t23 VSS 0.058005f
C7315 D2_1.n1 VSS 0.039372f
C7316 D2_1.n2 VSS 0.002882f
C7317 D2_1.t10 VSS 0.024214f
C7318 D2_1.t9 VSS 0.046004f
C7319 D2_1.t20 VSS 0.030658f
C7320 D2_1.n3 VSS 0.057268f
C7321 D2_1.t4 VSS 0.058005f
C7322 D2_1.n4 VSS 0.039372f
C7323 D2_1.t16 VSS 0.051001f
C7324 D2_1.t29 VSS 0.05562f
C7325 D2_1.t31 VSS 0.024214f
C7326 D2_1.t14 VSS 0.047144f
C7327 D2_1.n5 VSS 0.037005f
C7328 D2_1.t26 VSS 0.047144f
C7329 D2_1.n6 VSS 0.037005f
C7330 D2_1.t12 VSS 0.037705f
C7331 D2_1.n7 VSS 0.05113f
C7332 D2_1.t35 VSS 0.032025f
C7333 D2_1.t0 VSS 0.051887f
C7334 D2_1.t13 VSS 0.063506f
C7335 D2_1.n8 VSS 0.044857f
C7336 D2_1.n9 VSS 0.097543f
C7337 D2_1.t21 VSS 0.051001f
C7338 D2_1.t28 VSS 0.05562f
C7339 D2_1.t32 VSS 0.024214f
C7340 D2_1.t15 VSS 0.047144f
C7341 D2_1.n10 VSS 0.037005f
C7342 D2_1.t27 VSS 0.047144f
C7343 D2_1.n11 VSS 0.037005f
C7344 D2_1.t5 VSS 0.037705f
C7345 D2_1.n12 VSS 0.05113f
C7346 D2_1.t1 VSS 0.030853f
C7347 D2_1.t8 VSS 0.030853f
C7348 D2_1.n13 VSS 0.039501f
C7349 D2_1.t7 VSS 0.030853f
C7350 D2_1.t22 VSS 0.030853f
C7351 D2_1.n14 VSS 0.043853f
C7352 D2_1.t2 VSS 0.030853f
C7353 D2_1.n15 VSS 0.039501f
C7354 D2_1.t33 VSS 0.039348f
C7355 D2_1.t6 VSS 0.024214f
C7356 D2_1.t19 VSS 0.046595f
C7357 D2_1.t34 VSS 0.030446f
C7358 D2_1.n16 VSS 0.037764f
C7359 D2_1.t11 VSS 0.087901f
C7360 D2_1.t18 VSS 0.096665f
C7361 D2_1.n17 VSS 0.041172f
C7362 D2_1.t24 VSS 0.06493f
C7363 D2_1.n18 VSS 0.043136f
C7364 D2_1.t17 VSS 0.030756f
C7365 D2_1.n19 VSS 0.027206f
C7366 D2_1.n20 VSS 0.025893f
C7367 D2_1.n21 VSS 2.75759f
C7368 D2_1.n22 VSS 3.85644f
C7369 D2_1.n23 VSS 2.56612f
C7370 D2_1.n24 VSS 0.078217f
C7371 D2_6.t20 VSS 0.084926f
C7372 D2_6.t4 VSS 0.092618f
C7373 D2_6.t5 VSS 0.04032f
C7374 D2_6.t23 VSS 0.078503f
C7375 D2_6.n0 VSS 0.06162f
C7376 D2_6.t0 VSS 0.078503f
C7377 D2_6.n1 VSS 0.06162f
C7378 D2_6.t14 VSS 0.062785f
C7379 D2_6.n2 VSS 0.08514f
C7380 D2_6.t7 VSS 0.053327f
C7381 D2_6.t9 VSS 0.086401f
C7382 D2_6.t15 VSS 0.105748f
C7383 D2_6.n3 VSS 0.074694f
C7384 D2_6.n4 VSS 3.31367f
C7385 D2_6.t1 VSS 0.084926f
C7386 D2_6.t11 VSS 0.092618f
C7387 D2_6.t13 VSS 0.04032f
C7388 D2_6.t6 VSS 0.078503f
C7389 D2_6.n5 VSS 0.06162f
C7390 D2_6.t8 VSS 0.078503f
C7391 D2_6.n6 VSS 0.06162f
C7392 D2_6.t22 VSS 0.062785f
C7393 D2_6.n7 VSS 0.08514f
C7394 D2_6.t17 VSS 0.053327f
C7395 D2_6.t19 VSS 0.086401f
C7396 D2_6.t25 VSS 0.105748f
C7397 D2_6.n8 VSS 0.074694f
C7398 D2_6.n9 VSS 0.936568f
C7399 D2_6.t18 VSS 0.04032f
C7400 D2_6.t2 VSS 0.076605f
C7401 D2_6.t3 VSS 0.051051f
C7402 D2_6.n10 VSS 0.095361f
C7403 D2_6.t21 VSS 0.096589f
C7404 D2_6.n11 VSS 0.065562f
C7405 D2_6.n12 VSS 3.00958f
C7406 D2_6.n13 VSS 3.63476f
C7407 D2_6.n14 VSS 0.013784f
C7408 D2_6.t10 VSS 0.04032f
C7409 D2_6.t16 VSS 0.076605f
C7410 D2_6.t24 VSS 0.051051f
C7411 D2_6.n15 VSS 0.095361f
C7412 D2_6.t12 VSS 0.096589f
C7413 D2_6.n16 VSS 0.065562f
C7414 Q2.t0 VSS 0.08777f
C7415 Q2.t2 VSS 0.102202f
C7416 Q2.t1 VSS 0.079869f
C7417 Q2.n0 VSS 0.205524f
C7418 Q2.n1 VSS 0.157277f
C7419 Q2.t31 VSS 0.179897f
C7420 Q2.t25 VSS 0.211955f
C7421 Q2.t16 VSS 0.171182f
C7422 Q2.t13 VSS 0.279494f
C7423 Q2.t6 VSS 0.301281f
C7424 Q2.t18 VSS 0.301281f
C7425 Q2.t10 VSS 0.226771f
C7426 Q2.n2 VSS 0.15603f
C7427 Q2.n3 VSS 2.82875f
C7428 Q2.t17 VSS 0.077188f
C7429 Q2.t5 VSS 0.150283f
C7430 Q2.n4 VSS 0.117962f
C7431 Q2.t4 VSS 0.150283f
C7432 Q2.n5 VSS 0.117962f
C7433 Q2.t24 VSS 0.120193f
C7434 Q2.t28 VSS 0.162579f
C7435 Q2.t7 VSS 0.177303f
C7436 Q2.n6 VSS 0.162965f
C7437 Q2.t29 VSS 0.165402f
C7438 Q2.t8 VSS 0.198083f
C7439 Q2.t11 VSS 0.106353f
C7440 Q2.n7 VSS 0.137108f
C7441 Q2.n8 VSS 1.21664f
C7442 Q2.t9 VSS 0.077188f
C7443 Q2.t23 VSS 0.150283f
C7444 Q2.n9 VSS 0.117962f
C7445 Q2.t22 VSS 0.150283f
C7446 Q2.n10 VSS 0.117962f
C7447 Q2.t14 VSS 0.120193f
C7448 Q2.t19 VSS 0.162579f
C7449 Q2.t26 VSS 0.177303f
C7450 Q2.n11 VSS 0.162965f
C7451 Q2.t20 VSS 0.165402f
C7452 Q2.t27 VSS 0.198083f
C7453 Q2.t3 VSS 0.106353f
C7454 Q2.n12 VSS 0.137108f
C7455 Q2.n13 VSS 1.77966f
C7456 Q2.n14 VSS 6.34216f
C7457 Q2.n15 VSS 5.70428f
C7458 Q2.t15 VSS 0.077188f
C7459 Q2.t21 VSS 0.146649f
C7460 Q2.t30 VSS 0.09773f
C7461 Q2.n16 VSS 0.182555f
C7462 Q2.t12 VSS 0.184906f
C7463 Q2.n17 VSS 0.125508f
C7464 Q2.n18 VSS 2.96361f
C7465 p2_gen_magic_0.xnor_magic_1.OUT.t0 VSS 0.127292f
C7466 p2_gen_magic_0.xnor_magic_1.OUT.t1 VSS 0.144065f
C7467 p2_gen_magic_0.xnor_magic_1.OUT.t3 VSS 0.070532f
C7468 p2_gen_magic_0.xnor_magic_1.OUT.t5 VSS 0.134003f
C7469 p2_gen_magic_0.xnor_magic_1.OUT.t2 VSS 0.089302f
C7470 p2_gen_magic_0.xnor_magic_1.OUT.n0 VSS 0.166813f
C7471 p2_gen_magic_0.xnor_magic_1.OUT.t4 VSS 0.168961f
C7472 p2_gen_magic_0.xnor_magic_1.OUT.n1 VSS 0.114685f
C7473 p2_gen_magic_0.xnor_magic_1.OUT.n2 VSS 3.46427f
C7474 7b_counter_0.MDFF_0.QB.t0 VSS 0.103726f
C7475 7b_counter_0.MDFF_0.QB.t1 VSS 0.100648f
C7476 7b_counter_0.MDFF_0.mux_magic_0.IN1 VSS 1.25182f
C7477 7b_counter_0.MDFF_0.tspc2_magic_0.QB VSS 1.25153f
C7478 7b_counter_0.MDFF_0.QB.t2 VSS 0.056663f
C7479 7b_counter_0.MDFF_0.QB.t4 VSS 0.107654f
C7480 7b_counter_0.MDFF_0.QB.t5 VSS 0.071743f
C7481 7b_counter_0.MDFF_0.QB.n0 VSS 0.134013f
C7482 7b_counter_0.MDFF_0.QB.t7 VSS 0.135738f
C7483 7b_counter_0.MDFF_0.QB.n1 VSS 0.092135f
C7484 7b_counter_0.MDFF_0.QB.t6 VSS 0.091392f
C7485 7b_counter_0.MDFF_0.QB.t8 VSS 0.166994f
C7486 7b_counter_0.MDFF_0.QB.n2 VSS 0.175658f
C7487 7b_counter_0.MDFF_0.QB.n3 VSS 0.132038f
C7488 7b_counter_0.MDFF_0.QB.t3 VSS 0.075855f
C7489 7b_counter_0.MDFF_0.QB.n4 VSS 0.152402f
C7490 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t9 VSS 0.034107f
C7491 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t8 VSS 0.068433f
C7492 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n0 VSS 0.072648f
C7493 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t4 VSS 0.087197f
C7494 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t5 VSS 0.04375f
C7495 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n1 VSS 0.105769f
C7496 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t10 VSS 0.125816f
C7497 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t11 VSS 0.063854f
C7498 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t3 VSS 0.042221f
C7499 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n2 VSS 0.111875f
C7500 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n3 VSS 0.160137f
C7501 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t6 VSS 0.080066f
C7502 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n4 VSS 0.287322f
C7503 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t12 VSS 0.034107f
C7504 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t7 VSS 0.067915f
C7505 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.n5 VSS 0.067242f
C7506 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t0 VSS 0.038783f
C7507 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t2 VSS 0.04516f
C7508 7b_counter_0.MDFF_0.tspc2_magic_0.CLK.t1 VSS 0.035292f
C7509 D2_3.t1 VSS 0.043586f
C7510 D2_3.t3 VSS 0.082808f
C7511 D2_3.t10 VSS 0.055185f
C7512 D2_3.n0 VSS 0.103084f
C7513 D2_3.t0 VSS 0.104411f
C7514 D2_3.n1 VSS 0.070871f
C7515 D2_3.n2 VSS 0.005469f
C7516 D2_3.t16 VSS 0.043586f
C7517 D2_3.t14 VSS 0.082808f
C7518 D2_3.t22 VSS 0.055185f
C7519 D2_3.n3 VSS 0.103084f
C7520 D2_3.t13 VSS 0.104411f
C7521 D2_3.n4 VSS 0.070871f
C7522 D2_3.t25 VSS 0.093398f
C7523 D2_3.t11 VSS 0.114312f
C7524 D2_3.t17 VSS 0.057646f
C7525 D2_3.n5 VSS 0.080743f
C7526 D2_3.t20 VSS 0.043586f
C7527 D2_3.t24 VSS 0.08486f
C7528 D2_3.n6 VSS 0.06661f
C7529 D2_3.t19 VSS 0.08486f
C7530 D2_3.n7 VSS 0.06661f
C7531 D2_3.t5 VSS 0.06787f
C7532 D2_3.t2 VSS 0.091804f
C7533 D2_3.t15 VSS 0.100118f
C7534 D2_3.n8 VSS 0.092035f
C7535 D2_3.n9 VSS 0.877896f
C7536 D2_3.t9 VSS 0.043586f
C7537 D2_3.t12 VSS 0.08486f
C7538 D2_3.n10 VSS 0.06661f
C7539 D2_3.t7 VSS 0.08486f
C7540 D2_3.n11 VSS 0.06661f
C7541 D2_3.t23 VSS 0.06787f
C7542 D2_3.t21 VSS 0.091804f
C7543 D2_3.t6 VSS 0.100118f
C7544 D2_3.n12 VSS 0.092035f
C7545 D2_3.t18 VSS 0.093398f
C7546 D2_3.t4 VSS 0.114312f
C7547 D2_3.t8 VSS 0.057646f
C7548 D2_3.n13 VSS 0.080743f
C7549 D2_3.n14 VSS 1.87275f
C7550 D2_3.n15 VSS 3.15516f
C7551 D2_3.n16 VSS 1.27349f
C7552 D2_3.n17 VSS 0.008524f
C7553 p3_gen_magic_0.xnor_magic_1.inverter_magic_0.VIN VSS 1.8586f
C7554 p3_gen_magic_0.xnor_magic_1.B.t1 VSS 0.128777f
C7555 p3_gen_magic_0.xnor_magic_1.B.t3 VSS 0.14044f
C7556 p3_gen_magic_0.xnor_magic_1.B.t4 VSS 0.06114f
C7557 p3_gen_magic_0.xnor_magic_1.B.t0 VSS 0.119038f
C7558 p3_gen_magic_0.xnor_magic_1.B.n0 VSS 0.093437f
C7559 p3_gen_magic_0.xnor_magic_1.B.t2 VSS 0.119038f
C7560 p3_gen_magic_0.xnor_magic_1.B.n1 VSS 0.093437f
C7561 p3_gen_magic_0.xnor_magic_1.B.t7 VSS 0.095204f
C7562 p3_gen_magic_0.xnor_magic_1.B.n2 VSS 0.129101f
C7563 p3_gen_magic_0.xnor_magic_1.B.t5 VSS 0.080862f
C7564 p3_gen_magic_0.xnor_magic_1.B.t6 VSS 0.131014f
C7565 p3_gen_magic_0.xnor_magic_1.B.t8 VSS 0.160351f
C7566 p3_gen_magic_0.xnor_magic_1.B.n3 VSS 0.112838f
C7567 p3_gen_magic_0.inverter_magic_0.VOUT VSS 3.17673f
C7568 P2.t8 VSS 0.068718f
C7569 P2.t13 VSS 0.074941f
C7570 P2.t14 VSS 0.06352f
C7571 P2.t15 VSS 0.032625f
C7572 P2.t7 VSS 0.06352f
C7573 P2.n0 VSS 0.049859f
C7574 P2.n1 VSS 0.049859f
C7575 P2.t9 VSS 0.050802f
C7576 P2.n2 VSS 0.068898f
C7577 P2.t12 VSS 0.071048f
C7578 P2.t11 VSS 0.134639f
C7579 P2.t6 VSS 0.142007f
C7580 P2.t10 VSS 0.09406f
C7581 P2.t16 VSS 0.045386f
C7582 P2.n3 VSS 0.055692f
C7583 P2.n4 VSS 1.60648f
C7584 P2.t2 VSS 0.013682f
C7585 P2.t0 VSS 0.013682f
C7586 P2.n5 VSS 0.029497f
C7587 P2.t5 VSS 0.013682f
C7588 P2.t4 VSS 0.013682f
C7589 P2.n6 VSS 0.030834f
C7590 P2.t1 VSS 0.013682f
C7591 P2.t3 VSS 0.013682f
C7592 P2.n7 VSS 0.03456f
C7593 P2.n8 VSS 0.09643f
C7594 P2.n9 VSS 0.043893f
C7595 P2.n10 VSS 0.024368f
C7596 p2_gen_magic_0.xnor_magic_3.OUT.t0 VSS 0.058254f
C7597 p2_gen_magic_0.xnor_magic_3.OUT.t1 VSS 0.06593f
C7598 p2_gen_magic_0.xnor_magic_3.OUT.n0 VSS 1.20048f
C7599 p2_gen_magic_0.xnor_magic_3.OUT.t2 VSS 0.064556f
C7600 p2_gen_magic_0.xnor_magic_3.OUT.t3 VSS 0.158504f
C7601 p2_gen_magic_0.xnor_magic_3.OUT.t6 VSS 0.045944f
C7602 p2_gen_magic_0.xnor_magic_3.OUT.t4 VSS 0.075358f
C7603 p2_gen_magic_0.xnor_magic_3.OUT.t5 VSS 0.08538f
C7604 p2_gen_magic_0.xnor_magic_3.OUT.n1 VSS 0.061699f
C7605 p2_gen_magic_0.xnor_magic_3.OUT.n2 VSS 0.904176f
C7606 D2_4.n0 VSS 0.002695f
C7607 D2_4.t12 VSS 0.024065f
C7608 D2_4.t9 VSS 0.046853f
C7609 D2_4.n1 VSS 0.036777f
C7610 D2_4.t7 VSS 0.046853f
C7611 D2_4.n2 VSS 0.036777f
C7612 D2_4.t19 VSS 0.037472f
C7613 D2_4.t21 VSS 0.050687f
C7614 D2_4.t4 VSS 0.055277f
C7615 D2_4.n3 VSS 0.050814f
C7616 D2_4.t18 VSS 0.051567f
C7617 D2_4.t5 VSS 0.063114f
C7618 D2_4.t10 VSS 0.031827f
C7619 D2_4.n4 VSS 0.04458f
C7620 D2_4.n5 VSS 0.607015f
C7621 D2_4.t20 VSS 0.024065f
C7622 D2_4.t16 VSS 0.046853f
C7623 D2_4.n6 VSS 0.036777f
C7624 D2_4.t15 VSS 0.046853f
C7625 D2_4.n7 VSS 0.036777f
C7626 D2_4.t1 VSS 0.037472f
C7627 D2_4.t2 VSS 0.050687f
C7628 D2_4.t13 VSS 0.055277f
C7629 D2_4.n8 VSS 0.050814f
C7630 D2_4.t0 VSS 0.051567f
C7631 D2_4.t14 VSS 0.063114f
C7632 D2_4.t17 VSS 0.031827f
C7633 D2_4.n9 VSS 0.04458f
C7634 D2_4.n10 VSS 0.055741f
C7635 D2_4.n11 VSS 2.48612f
C7636 D2_4.t8 VSS 0.024065f
C7637 D2_4.t25 VSS 0.04572f
C7638 D2_4.t11 VSS 0.030469f
C7639 D2_4.n12 VSS 0.056915f
C7640 D2_4.t24 VSS 0.057648f
C7641 D2_4.n13 VSS 0.039129f
C7642 D2_4.n14 VSS 4.84524f
C7643 D2_4.n15 VSS 0.578724f
C7644 D2_4.t23 VSS 0.024065f
C7645 D2_4.t6 VSS 0.04572f
C7646 D2_4.t3 VSS 0.030469f
C7647 D2_4.n16 VSS 0.056915f
C7648 D2_4.t22 VSS 0.057648f
C7649 D2_4.n17 VSS 0.039129f
C7650 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t14 VSS 0.077899f
C7651 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t15 VSS 0.084954f
C7652 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t17 VSS 0.072008f
C7653 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t12 VSS 0.036984f
C7654 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t16 VSS 0.072008f
C7655 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n0 VSS 0.056521f
C7656 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n1 VSS 0.056521f
C7657 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t13 VSS 0.05759f
C7658 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n2 VSS 0.078106f
C7659 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t9 VSS 0.042992f
C7660 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t1 VSS 0.057766f
C7661 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t0 VSS 0.015509f
C7662 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t2 VSS 0.015509f
C7663 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n3 VSS 0.031019f
C7664 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n4 VSS 0.133091f
C7665 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t11 VSS 0.015509f
C7666 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t10 VSS 0.015509f
C7667 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n5 VSS 0.031019f
C7668 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n6 VSS 0.066219f
C7669 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n7 VSS 0.239497f
C7670 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t7 VSS 0.015509f
C7671 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t8 VSS 0.015509f
C7672 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n8 VSS 0.034953f
C7673 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t5 VSS 0.015509f
C7674 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t3 VSS 0.015509f
C7675 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n9 VSS 0.039178f
C7676 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t4 VSS 0.015509f
C7677 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.t6 VSS 0.015509f
C7678 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.IN.n10 VSS 0.033439f
C7679 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t20 VSS 0.063791f
C7680 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t19 VSS 0.063791f
C7681 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n0 VSS 0.07755f
C7682 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t9 VSS 0.094891f
C7683 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t18 VSS 0.065269f
C7684 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t7 VSS 0.07118f
C7685 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t14 VSS 0.060332f
C7686 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t12 VSS 0.030988f
C7687 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t17 VSS 0.060332f
C7688 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n1 VSS 0.047357f
C7689 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n2 VSS 0.047357f
C7690 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t22 VSS 0.048253f
C7691 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n3 VSS 0.065229f
C7692 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t6 VSS 0.063791f
C7693 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t21 VSS 0.063791f
C7694 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n4 VSS 0.07755f
C7695 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t15 VSS 0.094891f
C7696 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t13 VSS 0.030988f
C7697 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t10 VSS 0.060332f
C7698 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n5 VSS 0.047357f
C7699 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t16 VSS 0.060332f
C7700 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n6 VSS 0.047357f
C7701 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t11 VSS 0.048253f
C7702 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t8 VSS 0.065269f
C7703 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t23 VSS 0.07118f
C7704 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n7 VSS 0.065229f
C7705 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n8 VSS 0.717998f
C7706 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t5 VSS 0.012995f
C7707 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t4 VSS 0.012995f
C7708 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n9 VSS 0.029286f
C7709 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t2 VSS 0.012995f
C7710 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t1 VSS 0.012995f
C7711 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n10 VSS 0.032826f
C7712 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t0 VSS 0.012995f
C7713 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.t3 VSS 0.012995f
C7714 p3_gen_magic_0.neg_DFF_magic_0.tg_magic_1.CLK.n11 VSS 0.028017f
C7715 Q3.t24 VSS 0.107376f
C7716 Q3.t18 VSS 0.172024f
C7717 Q3.t3 VSS 0.133012f
C7718 Q3.t12 VSS 0.102174f
C7719 Q3.t6 VSS 0.166822f
C7720 Q3.t26 VSS 0.179826f
C7721 Q3.t14 VSS 0.136532f
C7722 Q3.n0 VSS 0.144911f
C7723 Q3.t0 VSS 0.052387f
C7724 Q3.t2 VSS 0.061001f
C7725 Q3.t1 VSS 0.047672f
C7726 Q3.n1 VSS 0.122672f
C7727 Q3.n2 VSS 0.093874f
C7728 Q3.t10 VSS 0.046071f
C7729 Q3.t22 VSS 0.087531f
C7730 Q3.t28 VSS 0.058332f
C7731 Q3.n3 VSS 0.108962f
C7732 Q3.t8 VSS 0.110365f
C7733 Q3.n4 VSS 0.074912f
C7734 Q3.n5 VSS 0.287237f
C7735 Q3.t19 VSS 0.098724f
C7736 Q3.t31 VSS 0.11823f
C7737 Q3.t9 VSS 0.063479f
C7738 Q3.n6 VSS 0.081836f
C7739 Q3.t11 VSS 0.046071f
C7740 Q3.t25 VSS 0.0897f
C7741 Q3.n7 VSS 0.070408f
C7742 Q3.t29 VSS 0.0897f
C7743 Q3.n8 VSS 0.070408f
C7744 Q3.t23 VSS 0.07174f
C7745 Q3.t21 VSS 0.097039f
C7746 Q3.t5 VSS 0.105827f
C7747 Q3.n9 VSS 0.097269f
C7748 Q3.n10 VSS 0.633063f
C7749 Q3.n11 VSS 0.67942f
C7750 Q3.t20 VSS 0.046071f
C7751 Q3.t7 VSS 0.0897f
C7752 Q3.n12 VSS 0.070408f
C7753 Q3.t13 VSS 0.0897f
C7754 Q3.n13 VSS 0.070408f
C7755 Q3.t4 VSS 0.07174f
C7756 Q3.t30 VSS 0.097039f
C7757 Q3.t16 VSS 0.105827f
C7758 Q3.n14 VSS 0.097269f
C7759 Q3.t27 VSS 0.098724f
C7760 Q3.t15 VSS 0.11823f
C7761 Q3.t17 VSS 0.063479f
C7762 Q3.n15 VSS 0.081836f
C7763 Q3.n16 VSS 0.236857f
C7764 Q3.n17 VSS 0.078405f
C7765 Q3.n18 VSS 2.66368f
C7766 Q3.n19 VSS 3.87282f
C7767 Q3.n20 VSS 0.499939f
C7768 Q3.n21 VSS 0.010393f
C7769 7b_counter_0.MDFF_6.QB.t0 VSS 0.16662f
C7770 7b_counter_0.MDFF_6.QB.t1 VSS 0.161675f
C7771 7b_counter_0.MDFF_6.mux_magic_0.IN1 VSS 1.43325f
C7772 7b_counter_0.MDFF_6.tspc2_magic_0.QB VSS 2.40197f
C7773 7b_counter_0.MDFF_6.QB.t4 VSS 0.09102f
C7774 7b_counter_0.MDFF_6.QB.t5 VSS 0.172929f
C7775 7b_counter_0.MDFF_6.QB.t7 VSS 0.115243f
C7776 7b_counter_0.MDFF_6.QB.n0 VSS 0.21527f
C7777 7b_counter_0.MDFF_6.QB.t3 VSS 0.218042f
C7778 7b_counter_0.MDFF_6.QB.n1 VSS 0.148f
C7779 7b_counter_0.MDFF_6.QB.t6 VSS 0.268685f
C7780 7b_counter_0.MDFF_6.QB.n2 VSS 0.282166f
C7781 7b_counter_0.MDFF_6.QB.n3 VSS 0.211662f
C7782 7b_counter_0.MDFF_6.QB.t8 VSS 0.122217f
C7783 7b_counter_0.MDFF_6.QB.t2 VSS 0.14644f
C7784 7b_counter_0.MDFF_6.QB.n4 VSS 0.24481f
C7785 CLK.t83 VSS 0.086585f
C7786 CLK.t71 VSS 0.086585f
C7787 CLK.n0 VSS 0.10526f
C7788 CLK.t17 VSS 0.228756f
C7789 CLK.t47 VSS 0.04206f
C7790 CLK.t11 VSS 0.08189f
C7791 CLK.n1 VSS 0.064278f
C7792 CLK.t101 VSS 0.08189f
C7793 CLK.n2 VSS 0.064278f
C7794 CLK.t56 VSS 0.065494f
C7795 CLK.t97 VSS 0.08859f
C7796 CLK.t24 VSS 0.096613f
C7797 CLK.n3 VSS 0.088536f
C7798 CLK.n4 VSS 0.276828f
C7799 CLK.t57 VSS 0.04206f
C7800 CLK.t118 VSS 0.07991f
C7801 CLK.t110 VSS 0.053253f
C7802 CLK.n5 VSS 0.099475f
C7803 CLK.t54 VSS 0.100756f
C7804 CLK.n6 VSS 0.06839f
C7805 CLK.n7 VSS 0.013478f
C7806 CLK.t85 VSS 0.04206f
C7807 CLK.t43 VSS 0.08189f
C7808 CLK.n8 VSS 0.064278f
C7809 CLK.t90 VSS 0.08189f
C7810 CLK.n9 VSS 0.064278f
C7811 CLK.t127 VSS 0.065494f
C7812 CLK.t9 VSS 0.08859f
C7813 CLK.t40 VSS 0.096613f
C7814 CLK.n10 VSS 0.088825f
C7815 CLK.t111 VSS 0.086585f
C7816 CLK.t62 VSS 0.086585f
C7817 CLK.n11 VSS 0.10526f
C7818 CLK.t59 VSS 0.228756f
C7819 CLK.t76 VSS 0.04206f
C7820 CLK.t36 VSS 0.08189f
C7821 CLK.n12 VSS 0.064278f
C7822 CLK.t3 VSS 0.08189f
C7823 CLK.n13 VSS 0.064278f
C7824 CLK.t121 VSS 0.065494f
C7825 CLK.t119 VSS 0.08859f
C7826 CLK.t28 VSS 0.096613f
C7827 CLK.n14 VSS 0.088536f
C7828 CLK.n15 VSS 0.276828f
C7829 CLK.n16 VSS 0.432761f
C7830 CLK.t48 VSS 0.086585f
C7831 CLK.t103 VSS 0.086585f
C7832 CLK.n17 VSS 0.10526f
C7833 CLK.t93 VSS 0.128796f
C7834 CLK.t126 VSS 0.08859f
C7835 CLK.t78 VSS 0.096613f
C7836 CLK.t115 VSS 0.08189f
C7837 CLK.t32 VSS 0.04206f
C7838 CLK.t29 VSS 0.08189f
C7839 CLK.n18 VSS 0.064278f
C7840 CLK.n19 VSS 0.064278f
C7841 CLK.t123 VSS 0.065494f
C7842 CLK.n20 VSS 0.088536f
C7843 CLK.n21 VSS 0.376636f
C7844 CLK.n22 VSS 0.129037f
C7845 CLK.n23 VSS 3.14261f
C7846 CLK.n24 VSS 2.36057f
C7847 CLK.t49 VSS 0.04206f
C7848 CLK.t45 VSS 0.07991f
C7849 CLK.t84 VSS 0.053253f
C7850 CLK.n25 VSS 0.099475f
C7851 CLK.t39 VSS 0.100756f
C7852 CLK.n26 VSS 0.06839f
C7853 CLK.n27 VSS 0.004758f
C7854 CLK.t104 VSS 0.046809f
C7855 CLK.t112 VSS 0.07991f
C7856 CLK.t21 VSS 0.053253f
C7857 CLK.n28 VSS 0.099475f
C7858 CLK.t108 VSS 0.102625f
C7859 CLK.n29 VSS 0.037257f
C7860 CLK.t0 VSS 0.04206f
C7861 CLK.t63 VSS 0.07991f
C7862 CLK.t80 VSS 0.053253f
C7863 CLK.n30 VSS 0.099475f
C7864 CLK.t117 VSS 0.100756f
C7865 CLK.n31 VSS 0.06839f
C7866 CLK.t124 VSS 0.04206f
C7867 CLK.t125 VSS 0.07991f
C7868 CLK.t33 VSS 0.053253f
C7869 CLK.n32 VSS 0.099475f
C7870 CLK.t116 VSS 0.100756f
C7871 CLK.n33 VSS 0.06839f
C7872 CLK.n34 VSS 0.350617f
C7873 CLK.t44 VSS 0.046809f
C7874 CLK.t61 VSS 0.07991f
C7875 CLK.t106 VSS 0.053253f
C7876 CLK.n35 VSS 0.099475f
C7877 CLK.t50 VSS 0.102625f
C7878 CLK.n36 VSS 0.037257f
C7879 CLK.n37 VSS 0.176659f
C7880 CLK.t69 VSS 0.04206f
C7881 CLK.t92 VSS 0.07991f
C7882 CLK.t102 VSS 0.053253f
C7883 CLK.n38 VSS 0.099475f
C7884 CLK.t30 VSS 0.100756f
C7885 CLK.n39 VSS 0.06839f
C7886 CLK.n40 VSS 0.025046f
C7887 CLK.t82 VSS 0.04206f
C7888 CLK.t94 VSS 0.07991f
C7889 CLK.t105 VSS 0.053253f
C7890 CLK.n41 VSS 0.099475f
C7891 CLK.t42 VSS 0.100756f
C7892 CLK.n42 VSS 0.06839f
C7893 CLK.n43 VSS 0.445523f
C7894 CLK.n44 VSS 2.56006f
C7895 CLK.n45 VSS 2.0705f
C7896 CLK.n46 VSS 0.469885f
C7897 CLK.n47 VSS 0.743474f
C7898 CLK.n48 VSS 1.08447f
C7899 CLK.t4 VSS 0.086585f
C7900 CLK.t95 VSS 0.086585f
C7901 CLK.n49 VSS 0.10526f
C7902 CLK.t60 VSS 0.228756f
C7903 CLK.t5 VSS 0.04206f
C7904 CLK.t89 VSS 0.08189f
C7905 CLK.n50 VSS 0.064278f
C7906 CLK.t51 VSS 0.08189f
C7907 CLK.n51 VSS 0.064278f
C7908 CLK.t14 VSS 0.065494f
C7909 CLK.t107 VSS 0.08859f
C7910 CLK.t70 VSS 0.096613f
C7911 CLK.n52 VSS 0.088536f
C7912 CLK.n53 VSS 0.276828f
C7913 CLK.t88 VSS 0.086585f
C7914 CLK.t72 VSS 0.086585f
C7915 CLK.n54 VSS 0.10526f
C7916 CLK.t18 VSS 0.128796f
C7917 CLK.t66 VSS 0.08859f
C7918 CLK.t13 VSS 0.096613f
C7919 CLK.t53 VSS 0.08189f
C7920 CLK.t26 VSS 0.04206f
C7921 CLK.t58 VSS 0.08189f
C7922 CLK.n55 VSS 0.064278f
C7923 CLK.n56 VSS 0.064278f
C7924 CLK.t100 VSS 0.065494f
C7925 CLK.n57 VSS 0.088536f
C7926 CLK.n58 VSS 0.376636f
C7927 CLK.n59 VSS 0.287515f
C7928 CLK.n60 VSS 0.351296f
C7929 CLK.t7 VSS 0.04206f
C7930 CLK.t34 VSS 0.08189f
C7931 CLK.n61 VSS 0.064278f
C7932 CLK.t77 VSS 0.08189f
C7933 CLK.n62 VSS 0.064278f
C7934 CLK.t38 VSS 0.065494f
C7935 CLK.t114 VSS 0.08859f
C7936 CLK.t8 VSS 0.096613f
C7937 CLK.n63 VSS 0.088825f
C7938 CLK.n64 VSS 0.57983f
C7939 CLK.n65 VSS 0.876944f
C7940 CLK.t73 VSS 0.04206f
C7941 CLK.t67 VSS 0.08189f
C7942 CLK.n66 VSS 0.064278f
C7943 CLK.t81 VSS 0.08189f
C7944 CLK.n67 VSS 0.064278f
C7945 CLK.t41 VSS 0.065494f
C7946 CLK.t22 VSS 0.08859f
C7947 CLK.t99 VSS 0.096613f
C7948 CLK.n68 VSS 0.088825f
C7949 CLK.t31 VSS 0.086585f
C7950 CLK.t79 VSS 0.086585f
C7951 CLK.n69 VSS 0.10526f
C7952 CLK.t55 VSS 0.228401f
C7953 CLK.t2 VSS 0.08859f
C7954 CLK.t87 VSS 0.096613f
C7955 CLK.t120 VSS 0.08189f
C7956 CLK.t98 VSS 0.04206f
C7957 CLK.t25 VSS 0.08189f
C7958 CLK.n70 VSS 0.064278f
C7959 CLK.n71 VSS 0.064278f
C7960 CLK.t52 VSS 0.065494f
C7961 CLK.n72 VSS 0.088536f
C7962 CLK.n73 VSS 0.277186f
C7963 CLK.t64 VSS 0.04206f
C7964 CLK.t122 VSS 0.08189f
C7965 CLK.n74 VSS 0.064278f
C7966 CLK.t113 VSS 0.08189f
C7967 CLK.n75 VSS 0.064278f
C7968 CLK.t86 VSS 0.064909f
C7969 CLK.t23 VSS 0.08859f
C7970 CLK.t35 VSS 0.09216f
C7971 CLK.n76 VSS 0.095477f
C7972 CLK.t20 VSS 0.086585f
C7973 CLK.t75 VSS 0.086585f
C7974 CLK.n77 VSS 0.10526f
C7975 CLK.t19 VSS 0.128777f
C7976 CLK.t46 VSS 0.04206f
C7977 CLK.t16 VSS 0.08189f
C7978 CLK.n78 VSS 0.064278f
C7979 CLK.t12 VSS 0.08189f
C7980 CLK.n79 VSS 0.064278f
C7981 CLK.t68 VSS 0.065494f
C7982 CLK.t6 VSS 0.08859f
C7983 CLK.t27 VSS 0.096613f
C7984 CLK.n80 VSS 0.088536f
C7985 CLK.n81 VSS 0.376822f
C7986 CLK.n82 VSS 0.514131f
C7987 CLK.n83 VSS 1.56944f
C7988 CLK.n84 VSS 0.59169f
C7989 CLK.n85 VSS 0.152601f
C7990 CLK.t1 VSS 0.086585f
C7991 CLK.t91 VSS 0.086585f
C7992 CLK.n86 VSS 0.10526f
C7993 CLK.t15 VSS 0.128796f
C7994 CLK.t74 VSS 0.08859f
C7995 CLK.t10 VSS 0.096613f
C7996 CLK.t109 VSS 0.08189f
C7997 CLK.t37 VSS 0.04206f
C7998 CLK.t65 VSS 0.08189f
C7999 CLK.n87 VSS 0.064278f
C8000 CLK.n88 VSS 0.064278f
C8001 CLK.t96 VSS 0.065494f
C8002 CLK.n89 VSS 0.088536f
C8003 CLK.n90 VSS 0.376636f
C8004 CLK.n91 VSS 0.287515f
C8005 CLK.n92 VSS 0.606294f
C8006 VDD.t1929 VSS 0.024488f
C8007 VDD.t1924 VSS 0.01669f
C8008 VDD.n0 VSS 0.056767f
C8009 VDD.n1 VSS 0.037445f
C8010 VDD.t1274 VSS 0.006764f
C8011 VDD.t1276 VSS 0.006764f
C8012 VDD.n2 VSS 0.018431f
C8013 VDD.t1286 VSS 0.006764f
C8014 VDD.t1288 VSS 0.006764f
C8015 VDD.n3 VSS 0.013528f
C8016 VDD.n4 VSS 0.032654f
C8017 VDD.n5 VSS 0.033392f
C8018 VDD.t1925 VSS 0.414138f
C8019 VDD.t1927 VSS 0.264656f
C8020 VDD.t1923 VSS 0.36819f
C8021 VDD.t1269 VSS 0.178275f
C8022 VDD.t1414 VSS 0.024488f
C8023 VDD.t1417 VSS 0.01669f
C8024 VDD.n6 VSS 0.056767f
C8025 VDD.t1415 VSS 0.006764f
C8026 VDD.t1416 VSS 0.006764f
C8027 VDD.n7 VSS 0.018431f
C8028 VDD.t1410 VSS 0.006764f
C8029 VDD.t1412 VSS 0.006764f
C8030 VDD.n8 VSS 0.013528f
C8031 VDD.n9 VSS 0.032654f
C8032 VDD.t1278 VSS 0.023942f
C8033 VDD.t1289 VSS 0.01669f
C8034 VDD.n10 VSS 0.056574f
C8035 VDD.n11 VSS 0.051957f
C8036 VDD.n12 VSS 0.051972f
C8037 VDD.n13 VSS 0.037445f
C8038 VDD.t1285 VSS 0.006764f
C8039 VDD.t1287 VSS 0.006764f
C8040 VDD.n14 VSS 0.018431f
C8041 VDD.t1270 VSS 0.006764f
C8042 VDD.t1272 VSS 0.006764f
C8043 VDD.n15 VSS 0.013528f
C8044 VDD.n16 VSS 0.032654f
C8045 VDD.t1266 VSS 0.023942f
C8046 VDD.t1283 VSS 0.01669f
C8047 VDD.n17 VSS 0.056465f
C8048 VDD.t995 VSS 0.006764f
C8049 VDD.t997 VSS 0.006764f
C8050 VDD.n18 VSS 0.018431f
C8051 VDD.t1000 VSS 0.006764f
C8052 VDD.t1001 VSS 0.006764f
C8053 VDD.n19 VSS 0.013528f
C8054 VDD.n20 VSS 0.032654f
C8055 VDD.n21 VSS 0.049867f
C8056 VDD.t1271 VSS 0.264656f
C8057 VDD.t1265 VSS 0.238926f
C8058 VDD.t1281 VSS 0.414138f
C8059 VDD.t1279 VSS 0.264656f
C8060 VDD.t1267 VSS 0.178275f
C8061 VDD.t999 VSS 0.024488f
C8062 VDD.t1002 VSS 0.01669f
C8063 VDD.n22 VSS 0.056767f
C8064 VDD.n23 VSS 0.037445f
C8065 VDD.t1268 VSS 0.006764f
C8066 VDD.t1280 VSS 0.006764f
C8067 VDD.n24 VSS 0.018431f
C8068 VDD.t1284 VSS 0.006764f
C8069 VDD.t1290 VSS 0.006764f
C8070 VDD.n25 VSS 0.013528f
C8071 VDD.n26 VSS 0.032654f
C8072 VDD.t1282 VSS 0.023942f
C8073 VDD.t1291 VSS 0.01669f
C8074 VDD.n27 VSS 0.059526f
C8075 VDD.t500 VSS 0.019461f
C8076 VDD.n28 VSS 0.006972f
C8077 VDD.n29 VSS 0.015826f
C8078 VDD.t499 VSS 0.161428f
C8079 VDD.t1296 VSS 0.233173f
C8080 VDD.t1302 VSS 0.101755f
C8081 VDD.t498 VSS 0.006764f
C8082 VDD.t1303 VSS 0.006764f
C8083 VDD.n30 VSS 0.015423f
C8084 VDD.n31 VSS 0.025914f
C8085 VDD.t1297 VSS 0.019459f
C8086 VDD.t771 VSS 0.021269f
C8087 VDD.t772 VSS 0.01669f
C8088 VDD.n32 VSS 0.068817f
C8089 VDD.t413 VSS 0.021269f
C8090 VDD.t411 VSS 0.01669f
C8091 VDD.n33 VSS 0.070928f
C8092 VDD.t409 VSS 0.006764f
C8093 VDD.t412 VSS 0.006764f
C8094 VDD.n34 VSS 0.013528f
C8095 VDD.n35 VSS 0.036172f
C8096 VDD.n36 VSS 0.032472f
C8097 VDD.t349 VSS 0.619833f
C8098 VDD.t347 VSS 0.375016f
C8099 VDD.t1704 VSS 0.548156f
C8100 VDD.t1750 VSS 0.006764f
C8101 VDD.t1771 VSS 0.006764f
C8102 VDD.n37 VSS 0.01683f
C8103 VDD.t1715 VSS 0.006764f
C8104 VDD.t1740 VSS 0.006764f
C8105 VDD.n38 VSS 0.013528f
C8106 VDD.n39 VSS 0.027737f
C8107 VDD.n40 VSS 0.015175f
C8108 VDD.t1773 VSS 0.01979f
C8109 VDD.t1705 VSS 0.01669f
C8110 VDD.n41 VSS 0.040346f
C8111 VDD.t371 VSS 0.021269f
C8112 VDD.t370 VSS 0.01669f
C8113 VDD.n42 VSS 0.068817f
C8114 VDD.t808 VSS 0.021269f
C8115 VDD.t807 VSS 0.01669f
C8116 VDD.n43 VSS 0.070928f
C8117 VDD.t809 VSS 0.006764f
C8118 VDD.t810 VSS 0.006764f
C8119 VDD.n44 VSS 0.013528f
C8120 VDD.n45 VSS 0.036172f
C8121 VDD.n46 VSS 0.032472f
C8122 VDD.t369 VSS 0.882358f
C8123 VDD.t425 VSS 0.375016f
C8124 VDD.t1768 VSS 0.138882f
C8125 VDD.t1747 VSS 0.01979f
C8126 VDD.t1762 VSS 0.01669f
C8127 VDD.n47 VSS 0.049398f
C8128 VDD.t1769 VSS 0.006764f
C8129 VDD.t1754 VSS 0.006764f
C8130 VDD.n48 VSS 0.01683f
C8131 VDD.t1775 VSS 0.006764f
C8132 VDD.t1743 VSS 0.006764f
C8133 VDD.n49 VSS 0.013528f
C8134 VDD.n50 VSS 0.027737f
C8135 VDD.t120 VSS 0.018157f
C8136 VDD.t118 VSS 0.006764f
C8137 VDD.t1233 VSS 0.006764f
C8138 VDD.n51 VSS 0.022549f
C8139 VDD.t1252 VSS 0.006764f
C8140 VDD.t1219 VSS 0.006764f
C8141 VDD.n52 VSS 0.022549f
C8142 VDD.t1217 VSS 0.018157f
C8143 VDD.t1221 VSS 0.021269f
C8144 VDD.t1223 VSS 0.01669f
C8145 VDD.n53 VSS 0.070928f
C8146 VDD.t1224 VSS 0.006764f
C8147 VDD.t1222 VSS 0.006764f
C8148 VDD.n54 VSS 0.013528f
C8149 VDD.n55 VSS 0.036172f
C8150 VDD.t1724 VSS 0.214331f
C8151 VDD.t1760 VSS 0.136969f
C8152 VDD.t879 VSS 0.136969f
C8153 VDD.t845 VSS 0.136969f
C8154 VDD.t2019 VSS 0.136969f
C8155 VDD.t2021 VSS 0.141408f
C8156 VDD.t1742 VSS 0.363892f
C8157 VDD.t119 VSS 0.214331f
C8158 VDD.t117 VSS 0.136969f
C8159 VDD.t1232 VSS 0.136969f
C8160 VDD.t1251 VSS 0.136969f
C8161 VDD.t1218 VSS 0.136969f
C8162 VDD.t1216 VSS 0.141408f
C8163 VDD.n56 VSS 0.356736f
C8164 VDD.t1220 VSS 0.408943f
C8165 VDD.t44 VSS 0.219141f
C8166 VDD.t1722 VSS 0.138882f
C8167 VDD.t1749 VSS 0.01979f
C8168 VDD.t1770 VSS 0.01669f
C8169 VDD.n57 VSS 0.040346f
C8170 VDD.t47 VSS 0.021269f
C8171 VDD.t46 VSS 0.01669f
C8172 VDD.n58 VSS 0.068817f
C8173 VDD.n59 VSS 0.072393f
C8174 VDD.n60 VSS 0.037945f
C8175 VDD.t1755 VSS 0.006764f
C8176 VDD.t1764 VSS 0.006764f
C8177 VDD.n61 VSS 0.01683f
C8178 VDD.t1723 VSS 0.006764f
C8179 VDD.t1737 VSS 0.006764f
C8180 VDD.n62 VSS 0.013528f
C8181 VDD.n63 VSS 0.027737f
C8182 VDD.t488 VSS 0.018157f
C8183 VDD.t621 VSS 0.047077f
C8184 VDD.t619 VSS 0.006764f
C8185 VDD.t51 VSS 0.006764f
C8186 VDD.n64 VSS 0.013528f
C8187 VDD.n65 VSS 0.057677f
C8188 VDD.t54 VSS 0.01669f
C8189 VDD.n66 VSS 0.026665f
C8190 VDD.n67 VSS 0.082093f
C8191 VDD.t202 VSS 0.538892f
C8192 VDD.t1147 VSS 0.214331f
C8193 VDD.t1038 VSS 0.136969f
C8194 VDD.t1817 VSS 0.136969f
C8195 VDD.t1815 VSS 0.136969f
C8196 VDD.t640 VSS 0.136969f
C8197 VDD.t638 VSS 0.214331f
C8198 VDD.t580 VSS 0.405502f
C8199 VDD.t1 VSS 0.194353f
C8200 VDD.t167 VSS 0.470286f
C8201 VDD.n68 VSS 0.475102f
C8202 VDD.t586 VSS 0.021269f
C8203 VDD.t581 VSS 0.01669f
C8204 VDD.n69 VSS 0.070928f
C8205 VDD.t585 VSS 0.006764f
C8206 VDD.t583 VSS 0.006764f
C8207 VDD.n70 VSS 0.013528f
C8208 VDD.n71 VSS 0.036172f
C8209 VDD.t577 VSS 0.018157f
C8210 VDD.t524 VSS 0.006764f
C8211 VDD.t603 VSS 0.006764f
C8212 VDD.n72 VSS 0.022549f
C8213 VDD.t605 VSS 0.006764f
C8214 VDD.t579 VSS 0.006764f
C8215 VDD.n73 VSS 0.022549f
C8216 VDD.t526 VSS 0.018157f
C8217 VDD.n74 VSS 0.03146f
C8218 VDD.t1148 VSS 0.018316f
C8219 VDD.t1039 VSS 0.006764f
C8220 VDD.t1818 VSS 0.006764f
C8221 VDD.n75 VSS 0.022549f
C8222 VDD.t1816 VSS 0.006764f
C8223 VDD.t641 VSS 0.006764f
C8224 VDD.n76 VSS 0.022549f
C8225 VDD.t639 VSS 0.025643f
C8226 VDD.n77 VSS 0.104443f
C8227 VDD.n78 VSS 0.044574f
C8228 VDD.t658 VSS 0.047077f
C8229 VDD.t656 VSS 0.006764f
C8230 VDD.t992 VSS 0.006764f
C8231 VDD.n79 VSS 0.013528f
C8232 VDD.n80 VSS 0.057677f
C8233 VDD.t993 VSS 0.01669f
C8234 VDD.n81 VSS 0.026665f
C8235 VDD.t2123 VSS 0.017784f
C8236 VDD.t2124 VSS 0.006764f
C8237 VDD.t1625 VSS 0.006764f
C8238 VDD.n82 VSS 0.020425f
C8239 VDD.n83 VSS 0.059702f
C8240 VDD.t1623 VSS 0.01669f
C8241 VDD.n84 VSS 0.017903f
C8242 VDD.t1628 VSS 0.006764f
C8243 VDD.t1626 VSS 0.006764f
C8244 VDD.n85 VSS 0.020425f
C8245 VDD.n86 VSS 0.039154f
C8246 VDD.n87 VSS 0.095546f
C8247 VDD.t2120 VSS 0.286484f
C8248 VDD.t309 VSS 0.195308f
C8249 VDD.t1366 VSS 0.214331f
C8250 VDD.t1344 VSS 0.136969f
C8251 VDD.t1173 VSS 0.136969f
C8252 VDD.t1191 VSS 0.136969f
C8253 VDD.t1552 VSS 0.136969f
C8254 VDD.t1550 VSS 0.214331f
C8255 VDD.t717 VSS 0.168403f
C8256 VDD.t661 VSS 0.080714f
C8257 VDD.t660 VSS 0.159603f
C8258 VDD.t310 VSS 0.021269f
C8259 VDD.t312 VSS 0.01669f
C8260 VDD.n88 VSS 0.084502f
C8261 VDD.t718 VSS 0.021269f
C8262 VDD.t722 VSS 0.01669f
C8263 VDD.n89 VSS 0.070928f
C8264 VDD.t721 VSS 0.006764f
C8265 VDD.t720 VSS 0.006764f
C8266 VDD.n90 VSS 0.013528f
C8267 VDD.n91 VSS 0.036172f
C8268 VDD.t716 VSS 0.018157f
C8269 VDD.t714 VSS 0.006764f
C8270 VDD.t753 VSS 0.006764f
C8271 VDD.n92 VSS 0.014917f
C8272 VDD.t755 VSS 0.006764f
C8273 VDD.t366 VSS 0.006764f
C8274 VDD.n93 VSS 0.014917f
C8275 VDD.t368 VSS 0.018157f
C8276 VDD.t1374 VSS 0.006764f
C8277 VDD.t1320 VSS 0.006764f
C8278 VDD.n94 VSS 0.01683f
C8279 VDD.t1311 VSS 0.006764f
C8280 VDD.t1359 VSS 0.006764f
C8281 VDD.n95 VSS 0.013528f
C8282 VDD.n96 VSS 0.027737f
C8283 VDD.t1357 VSS 0.01979f
C8284 VDD.t1352 VSS 0.01669f
C8285 VDD.n97 VSS 0.040346f
C8286 VDD.n98 VSS 0.037945f
C8287 VDD.t719 VSS 0.45143f
C8288 VDD.t715 VSS 0.214331f
C8289 VDD.t713 VSS 0.136969f
C8290 VDD.t752 VSS 0.136969f
C8291 VDD.t754 VSS 0.136969f
C8292 VDD.t365 VSS 0.136969f
C8293 VDD.t367 VSS 0.214331f
C8294 VDD.t1310 VSS 0.363892f
C8295 VDD.t1319 VSS 0.138882f
C8296 VDD.t223 VSS 0.219141f
C8297 VDD.t206 VSS 0.021269f
C8298 VDD.t205 VSS 0.01669f
C8299 VDD.n99 VSS 0.068817f
C8300 VDD.n100 VSS 0.072393f
C8301 VDD.t225 VSS 0.021269f
C8302 VDD.t226 VSS 0.01669f
C8303 VDD.n101 VSS 0.070928f
C8304 VDD.t224 VSS 0.006764f
C8305 VDD.t222 VSS 0.006764f
C8306 VDD.n102 VSS 0.013528f
C8307 VDD.n103 VSS 0.036172f
C8308 VDD.t247 VSS 0.018157f
C8309 VDD.t245 VSS 0.006764f
C8310 VDD.t1521 VSS 0.006764f
C8311 VDD.n104 VSS 0.014917f
C8312 VDD.t1547 VSS 0.006764f
C8313 VDD.t482 VSS 0.006764f
C8314 VDD.n105 VSS 0.014917f
C8315 VDD.t484 VSS 0.018157f
C8316 VDD.t1382 VSS 0.006764f
C8317 VDD.t1330 VSS 0.006764f
C8318 VDD.n106 VSS 0.01683f
C8319 VDD.t1378 VSS 0.006764f
C8320 VDD.t1368 VSS 0.006764f
C8321 VDD.n107 VSS 0.013528f
C8322 VDD.n108 VSS 0.027737f
C8323 VDD.t1341 VSS 0.01979f
C8324 VDD.t1358 VSS 0.01669f
C8325 VDD.n109 VSS 0.049398f
C8326 VDD.t1353 VSS 0.214331f
C8327 VDD.t1314 VSS 0.136969f
C8328 VDD.t881 VSS 0.136969f
C8329 VDD.t875 VSS 0.136969f
C8330 VDD.t2160 VSS 0.136969f
C8331 VDD.t2158 VSS 0.141408f
C8332 VDD.t221 VSS 0.408943f
C8333 VDD.n110 VSS 0.356736f
C8334 VDD.t246 VSS 0.141408f
C8335 VDD.t244 VSS 0.136969f
C8336 VDD.t1520 VSS 0.136969f
C8337 VDD.t1546 VSS 0.136969f
C8338 VDD.t481 VSS 0.136969f
C8339 VDD.t483 VSS 0.214331f
C8340 VDD.t1377 VSS 0.363892f
C8341 VDD.t1329 VSS 0.138882f
C8342 VDD.t1340 VSS 0.341283f
C8343 VDD.n111 VSS 0.102565f
C8344 VDD.n112 VSS 0.018755f
C8345 VDD.n113 VSS 0.015175f
C8346 VDD.n114 VSS 0.037558f
C8347 VDD.t882 VSS 0.006764f
C8348 VDD.t1315 VSS 0.006764f
C8349 VDD.n115 VSS 0.014917f
C8350 VDD.t2161 VSS 0.006764f
C8351 VDD.t876 VSS 0.006764f
C8352 VDD.n116 VSS 0.014917f
C8353 VDD.t2159 VSS 0.022409f
C8354 VDD.n117 VSS 0.096335f
C8355 VDD.n118 VSS 0.033732f
C8356 VDD.t1354 VSS 0.018316f
C8357 VDD.n119 VSS 0.096908f
C8358 VDD.n120 VSS 0.07211f
C8359 VDD.n121 VSS 0.033732f
C8360 VDD.n122 VSS 0.0563f
C8361 VDD.n123 VSS 0.056289f
C8362 VDD.n124 VSS 0.032472f
C8363 VDD.n125 VSS -0.002571f
C8364 VDD.n126 VSS 0.189733f
C8365 VDD.t775 VSS 0.375016f
C8366 VDD.t204 VSS 0.882358f
C8367 VDD.t1351 VSS 0.548156f
C8368 VDD.n127 VSS 0.102565f
C8369 VDD.n128 VSS 0.006361f
C8370 VDD.n129 VSS 0.015175f
C8371 VDD.n130 VSS 0.037558f
C8372 VDD.t146 VSS 0.047077f
C8373 VDD.t1865 VSS 0.006764f
C8374 VDD.t148 VSS 0.006764f
C8375 VDD.n131 VSS 0.013528f
C8376 VDD.n132 VSS 0.057677f
C8377 VDD.t1868 VSS 0.01669f
C8378 VDD.n133 VSS 0.026665f
C8379 VDD.n134 VSS 0.075391f
C8380 VDD.t2026 VSS 0.031315f
C8381 VDD.t438 VSS 0.233099f
C8382 VDD.t1373 VSS 0.006764f
C8383 VDD.t1316 VSS 0.006764f
C8384 VDD.n135 VSS 0.01683f
C8385 VDD.t1372 VSS 0.006764f
C8386 VDD.t1309 VSS 0.006764f
C8387 VDD.n136 VSS 0.013528f
C8388 VDD.n137 VSS 0.027737f
C8389 VDD.t241 VSS 0.018157f
C8390 VDD.t67 VSS 0.006764f
C8391 VDD.t243 VSS 0.006764f
C8392 VDD.n138 VSS 0.014917f
C8393 VDD.t685 VSS 0.006764f
C8394 VDD.t69 VSS 0.006764f
C8395 VDD.n139 VSS 0.014917f
C8396 VDD.t687 VSS 0.018157f
C8397 VDD.t182 VSS 0.021269f
C8398 VDD.t187 VSS 0.01669f
C8399 VDD.n140 VSS 0.070928f
C8400 VDD.t184 VSS 0.006764f
C8401 VDD.t186 VSS 0.006764f
C8402 VDD.n141 VSS 0.013528f
C8403 VDD.n142 VSS 0.036172f
C8404 VDD.t780 VSS 0.021269f
C8405 VDD.t781 VSS 0.01669f
C8406 VDD.n143 VSS 0.084502f
C8407 VDD.t183 VSS 0.106074f
C8408 VDD.t456 VSS 0.257368f
C8409 VDD.t2 VSS 0.185753f
C8410 VDD.t457 VSS 0.153301f
C8411 VDD.t0 VSS 0.153301f
C8412 VDD.t779 VSS 0.133961f
C8413 VDD.n144 VSS 0.273232f
C8414 VDD.t1364 VSS 0.214331f
C8415 VDD.t1336 VSS 0.136969f
C8416 VDD.t1951 VSS 0.136969f
C8417 VDD.t1971 VSS 0.136969f
C8418 VDD.t723 VSS 0.136969f
C8419 VDD.t725 VSS 0.214331f
C8420 VDD.t181 VSS 0.106193f
C8421 VDD.t240 VSS 0.241577f
C8422 VDD.t2025 VSS 0.241577f
C8423 VDD.t242 VSS 0.031315f
C8424 VDD.t145 VSS 0.241577f
C8425 VDD.t66 VSS 0.241577f
C8426 VDD.t147 VSS 0.241577f
C8427 VDD.t68 VSS 0.241577f
C8428 VDD.t1864 VSS 0.241577f
C8429 VDD.t684 VSS 0.479799f
C8430 VDD.t686 VSS 0.538793f
C8431 VDD.t185 VSS 0.309392f
C8432 VDD.n145 VSS 0.198052f
C8433 VDD.t455 VSS 0.043838f
C8434 VDD.n146 VSS 0.353833f
C8435 VDD.n147 VSS 0.015297f
C8436 VDD.n148 VSS 0.004321f
C8437 VDD.n149 VSS 0.032472f
C8438 VDD.n150 VSS 0.056289f
C8439 VDD.n151 VSS 0.0563f
C8440 VDD.n152 VSS 0.033732f
C8441 VDD.t461 VSS 0.047077f
C8442 VDD.t62 VSS 0.006764f
C8443 VDD.t459 VSS 0.006764f
C8444 VDD.n153 VSS 0.013528f
C8445 VDD.n154 VSS 0.057677f
C8446 VDD.t63 VSS 0.01669f
C8447 VDD.n155 VSS 0.026665f
C8448 VDD.n156 VSS 0.352884f
C8449 VDD.n157 VSS 0.060215f
C8450 VDD.n158 VSS 0.02382f
C8451 VDD.n159 VSS 0.031299f
C8452 VDD.n160 VSS 0.019625f
C8453 VDD.n161 VSS 0.019349f
C8454 VDD.n162 VSS 0.017137f
C8455 VDD.n163 VSS 0.017552f
C8456 VDD.n164 VSS 0.017552f
C8457 VDD.n165 VSS 0.068756f
C8458 VDD.n166 VSS 0.019902f
C8459 VDD.n167 VSS 0.019902f
C8460 VDD.n168 VSS 1.10032f
C8461 VDD.n169 VSS 0.010248f
C8462 VDD.n170 VSS 0.001108f
C8463 VDD.n171 VSS 0.019487f
C8464 VDD.n172 VSS 0.019625f
C8465 VDD.n173 VSS 0.019349f
C8466 VDD.n174 VSS 0.017137f
C8467 VDD.n175 VSS 2.75668f
C8468 VDD.t948 VSS 0.018157f
C8469 VDD.t160 VSS 0.018157f
C8470 VDD.t1861 VSS 0.006764f
C8471 VDD.t162 VSS 0.006764f
C8472 VDD.n176 VSS 0.014917f
C8473 VDD.t166 VSS 0.006764f
C8474 VDD.t1863 VSS 0.006764f
C8475 VDD.n177 VSS 0.014917f
C8476 VDD.t164 VSS 0.022409f
C8477 VDD.n178 VSS 0.096335f
C8478 VDD.n179 VSS 0.034926f
C8479 VDD.n180 VSS 0.056306f
C8480 VDD.n181 VSS 0.054505f
C8481 VDD.t946 VSS 0.006764f
C8482 VDD.t757 VSS 0.006764f
C8483 VDD.n182 VSS 0.014917f
C8484 VDD.t759 VSS 0.006764f
C8485 VDD.t1632 VSS 0.006764f
C8486 VDD.n183 VSS 0.014917f
C8487 VDD.t1630 VSS 0.018157f
C8488 VDD.t1180 VSS 0.018322f
C8489 VDD.t1184 VSS 0.006764f
C8490 VDD.t1186 VSS 0.006764f
C8491 VDD.n184 VSS 0.015166f
C8492 VDD.t163 VSS 0.214331f
C8493 VDD.t165 VSS 0.136969f
C8494 VDD.t1862 VSS 0.136969f
C8495 VDD.t1860 VSS 0.136969f
C8496 VDD.t161 VSS 0.136969f
C8497 VDD.t159 VSS 0.242866f
C8498 VDD.t947 VSS 0.242866f
C8499 VDD.t945 VSS 0.136969f
C8500 VDD.t756 VSS 0.136969f
C8501 VDD.t758 VSS 0.136969f
C8502 VDD.t1631 VSS 0.136969f
C8503 VDD.t1629 VSS 0.262997f
C8504 VDD.t1179 VSS 0.278568f
C8505 VDD.t1183 VSS 0.114849f
C8506 VDD.t1542 VSS 0.146509f
C8507 VDD.t1536 VSS 0.006764f
C8508 VDD.t1541 VSS 0.006764f
C8509 VDD.n185 VSS 0.018548f
C8510 VDD.t141 VSS 0.006764f
C8511 VDD.t139 VSS 0.006764f
C8512 VDD.n186 VSS 0.013528f
C8513 VDD.n187 VSS 0.032109f
C8514 VDD.t1176 VSS 0.018322f
C8515 VDD.n188 VSS 0.103126f
C8516 VDD.n189 VSS 0.07921f
C8517 VDD.t1543 VSS 0.018294f
C8518 VDD.t1526 VSS 0.006764f
C8519 VDD.t1535 VSS 0.006764f
C8520 VDD.n190 VSS 0.015166f
C8521 VDD.t1525 VSS 0.114849f
C8522 VDD.t1831 VSS 0.103398f
C8523 VDD.t1826 VSS 0.006764f
C8524 VDD.t1832 VSS 0.006764f
C8525 VDD.n191 VSS 0.015166f
C8526 VDD.t1822 VSS 0.018322f
C8527 VDD.t1549 VSS 0.018322f
C8528 VDD.n192 VSS 0.07543f
C8529 VDD.n193 VSS 0.077762f
C8530 VDD.n194 VSS 0.046076f
C8531 VDD.t1824 VSS 0.018322f
C8532 VDD.t2002 VSS 0.006764f
C8533 VDD.t2009 VSS 0.006764f
C8534 VDD.n195 VSS 0.018548f
C8535 VDD.t6 VSS 0.006764f
C8536 VDD.t4 VSS 0.006764f
C8537 VDD.n196 VSS 0.013528f
C8538 VDD.n197 VSS 0.032136f
C8539 VDD.t1823 VSS 0.229878f
C8540 VDD.t423 VSS 0.409363f
C8541 VDD.t422 VSS 0.259137f
C8542 VDD.t5 VSS 0.259137f
C8543 VDD.t3 VSS 0.310025f
C8544 VDD.t1992 VSS 0.103398f
C8545 VDD.t2013 VSS 0.006764f
C8546 VDD.t1993 VSS 0.006764f
C8547 VDD.n198 VSS 0.015166f
C8548 VDD.t2008 VSS 0.018294f
C8549 VDD.n199 VSS 0.058631f
C8550 VDD.n200 VSS 0.045731f
C8551 VDD.t2006 VSS 0.018322f
C8552 VDD.t1964 VSS 0.018322f
C8553 VDD.t1966 VSS 0.006764f
C8554 VDD.t1958 VSS 0.006764f
C8555 VDD.n201 VSS 0.015166f
C8556 VDD.t1962 VSS 0.018322f
C8557 VDD.n202 VSS 0.084648f
C8558 VDD.t2005 VSS 0.266747f
C8559 VDD.t1963 VSS 0.266747f
C8560 VDD.t1965 VSS 0.114849f
C8561 VDD.t1436 VSS 0.146509f
C8562 VDD.t1448 VSS 0.006764f
C8563 VDD.t1433 VSS 0.006764f
C8564 VDD.n203 VSS 0.018548f
C8565 VDD.t176 VSS 0.006764f
C8566 VDD.t174 VSS 0.006764f
C8567 VDD.n204 VSS 0.013528f
C8568 VDD.n205 VSS 0.032136f
C8569 VDD.n206 VSS 0.045582f
C8570 VDD.t1437 VSS 0.018294f
C8571 VDD.t1442 VSS 0.006764f
C8572 VDD.t1445 VSS 0.006764f
C8573 VDD.n207 VSS 0.015166f
C8574 VDD.t1441 VSS 0.114849f
C8575 VDD.t1789 VSS 0.103398f
C8576 VDD.t1807 VSS 0.006764f
C8577 VDD.t1790 VSS 0.006764f
C8578 VDD.n208 VSS 0.015166f
C8579 VDD.t1792 VSS 0.018322f
C8580 VDD.t1432 VSS 0.018322f
C8581 VDD.n209 VSS 0.074239f
C8582 VDD.n210 VSS 0.075804f
C8583 VDD.n211 VSS 0.046076f
C8584 VDD.t1801 VSS 0.018322f
C8585 VDD.t2141 VSS 0.006764f
C8586 VDD.t2127 VSS 0.006764f
C8587 VDD.n212 VSS 0.018548f
C8588 VDD.t433 VSS 0.006764f
C8589 VDD.t435 VSS 0.006764f
C8590 VDD.n213 VSS 0.013528f
C8591 VDD.n214 VSS 0.032136f
C8592 VDD.t1800 VSS 0.229878f
C8593 VDD.t405 VSS 0.409363f
C8594 VDD.t406 VSS 0.259137f
C8595 VDD.t432 VSS 0.259137f
C8596 VDD.t434 VSS 0.310025f
C8597 VDD.t2144 VSS 0.227678f
C8598 VDD.t2139 VSS 0.103398f
C8599 VDD.t2138 VSS 0.006764f
C8600 VDD.t2140 VSS 0.006764f
C8601 VDD.n215 VSS 0.015166f
C8602 VDD.t2143 VSS 0.018294f
C8603 VDD.n216 VSS 0.058631f
C8604 VDD.n217 VSS 0.045731f
C8605 VDD.t2145 VSS 0.018322f
C8606 VDD.t1675 VSS 0.035637f
C8607 VDD.t1683 VSS 0.006764f
C8608 VDD.t1672 VSS 0.006764f
C8609 VDD.n218 VSS 0.015166f
C8610 VDD.t1679 VSS 0.03306f
C8611 VDD.n219 VSS 0.026295f
C8612 VDD.n220 VSS 0.019667f
C8613 VDD.t802 VSS 0.310025f
C8614 VDD.t1690 VSS 0.006764f
C8615 VDD.t1680 VSS 0.006764f
C8616 VDD.n221 VSS 0.018548f
C8617 VDD.t805 VSS 0.006764f
C8618 VDD.t803 VSS 0.006764f
C8619 VDD.n222 VSS 0.013528f
C8620 VDD.n223 VSS 0.032136f
C8621 VDD.t1847 VSS 0.114849f
C8622 VDD.t2051 VSS 0.018322f
C8623 VDD.t2053 VSS 0.006764f
C8624 VDD.t2039 VSS 0.006764f
C8625 VDD.n224 VSS 0.015166f
C8626 VDD.t2059 VSS 0.018322f
C8627 VDD.t1256 VSS 0.018322f
C8628 VDD.t1239 VSS 0.006764f
C8629 VDD.t1248 VSS 0.006764f
C8630 VDD.n225 VSS 0.015166f
C8631 VDD.t1258 VSS 0.034094f
C8632 VDD.n226 VSS 0.042374f
C8633 VDD.n227 VSS 0.030866f
C8634 VDD.n228 VSS 0.030866f
C8635 VDD.n229 VSS 0.02436f
C8636 VDD.n230 VSS 0.031399f
C8637 VDD.t1858 VSS 0.006764f
C8638 VDD.t1842 VSS 0.006764f
C8639 VDD.n231 VSS 0.018548f
C8640 VDD.t326 VSS 0.006764f
C8641 VDD.t324 VSS 0.006764f
C8642 VDD.n232 VSS 0.013528f
C8643 VDD.n233 VSS 0.031682f
C8644 VDD.t1840 VSS 0.028156f
C8645 VDD.t1848 VSS 0.006764f
C8646 VDD.t1856 VSS 0.006764f
C8647 VDD.n234 VSS 0.015166f
C8648 VDD.t1838 VSS 0.018322f
C8649 VDD.t2089 VSS 0.018322f
C8650 VDD.t2093 VSS 0.006764f
C8651 VDD.t2073 VSS 0.006764f
C8652 VDD.n235 VSS 0.015166f
C8653 VDD.t2087 VSS 0.027282f
C8654 VDD.n236 VSS 0.042575f
C8655 VDD.n237 VSS 0.029938f
C8656 VDD.n238 VSS 0.029938f
C8657 VDD.n239 VSS 0.025565f
C8658 VDD.n240 VSS 0.022589f
C8659 VDD.n241 VSS 0.01248f
C8660 VDD.n242 VSS 0.105693f
C8661 VDD.t2052 VSS 0.114849f
C8662 VDD.t302 VSS 0.310025f
C8663 VDD.t1254 VSS 0.006764f
C8664 VDD.t1229 VSS 0.006764f
C8665 VDD.n243 VSS 0.018548f
C8666 VDD.t305 VSS 0.006764f
C8667 VDD.t303 VSS 0.006764f
C8668 VDD.n244 VSS 0.013528f
C8669 VDD.n245 VSS 0.032136f
C8670 VDD.t1396 VSS 0.027262f
C8671 VDD.t1406 VSS 0.006764f
C8672 VDD.t1388 VSS 0.006764f
C8673 VDD.n246 VSS 0.015166f
C8674 VDD.t1400 VSS 0.027282f
C8675 VDD.n247 VSS 0.038369f
C8676 VDD.n248 VSS 0.078978f
C8677 VDD.t1395 VSS 0.227678f
C8678 VDD.t1405 VSS 0.114849f
C8679 VDD.t304 VSS 0.259137f
C8680 VDD.t653 VSS 0.259137f
C8681 VDD.t654 VSS 0.409363f
C8682 VDD.t1399 VSS 0.229878f
C8683 VDD.t1387 VSS 0.103398f
C8684 VDD.n249 VSS 0.061018f
C8685 VDD.n250 VSS -0.010365f
C8686 VDD.t70 VSS 0.470588f
C8687 VDD.t745 VSS 0.331315f
C8688 VDD.t1477 VSS 0.185802f
C8689 VDD.t123 VSS 0.006764f
C8690 VDD.t743 VSS 0.006764f
C8691 VDD.n251 VSS 0.029826f
C8692 VDD.t746 VSS 0.006764f
C8693 VDD.t1478 VSS 0.006764f
C8694 VDD.n252 VSS 0.013528f
C8695 VDD.n253 VSS 0.039293f
C8696 VDD.t122 VSS 0.006764f
C8697 VDD.t744 VSS 0.006764f
C8698 VDD.n254 VSS 0.029015f
C8699 VDD.n255 VSS 0.03765f
C8700 VDD.t747 VSS 0.006764f
C8701 VDD.t1479 VSS 0.006764f
C8702 VDD.n256 VSS 0.013528f
C8703 VDD.n257 VSS 0.008042f
C8704 VDD.t220 VSS 0.034731f
C8705 VDD.t832 VSS 0.018322f
C8706 VDD.n258 VSS -0.073356f
C8707 VDD.t1912 VSS 0.006764f
C8708 VDD.t818 VSS 0.006764f
C8709 VDD.n259 VSS 0.015166f
C8710 VDD.n260 VSS 0.035907f
C8711 VDD.t1492 VSS 0.116433f
C8712 VDD.t1493 VSS 0.006764f
C8713 VDD.t1499 VSS 0.006764f
C8714 VDD.n261 VSS 0.015166f
C8715 VDD.t1495 VSS 0.018322f
C8716 VDD.t795 VSS 0.018322f
C8717 VDD.t801 VSS 0.006764f
C8718 VDD.t797 VSS 0.006764f
C8719 VDD.n262 VSS 0.015166f
C8720 VDD.t799 VSS 0.022391f
C8721 VDD.n263 VSS 0.095048f
C8722 VDD.t1909 VSS 0.116433f
C8723 VDD.t1910 VSS 0.006764f
C8724 VDD.t1897 VSS 0.006764f
C8725 VDD.n264 VSS 0.015166f
C8726 VDD.t864 VSS 0.018322f
C8727 VDD.t1016 VSS 0.028459f
C8728 VDD.t1012 VSS 0.006764f
C8729 VDD.t1014 VSS 0.006764f
C8730 VDD.n265 VSS 0.015166f
C8731 VDD.t1018 VSS 0.028486f
C8732 VDD.n266 VSS 0.034939f
C8733 VDD.t2066 VSS 0.018422f
C8734 VDD.t2063 VSS 0.006764f
C8735 VDD.t2068 VSS 0.006764f
C8736 VDD.n267 VSS 0.015166f
C8737 VDD.n268 VSS 0.029124f
C8738 VDD.t2065 VSS 0.227678f
C8739 VDD.t2062 VSS 0.103398f
C8740 VDD.t1496 VSS 0.116433f
C8741 VDD.t1503 VSS 0.018322f
C8742 VDD.t2061 VSS 0.018313f
C8743 VDD.t1481 VSS 0.018322f
C8744 VDD.n269 VSS 0.071098f
C8745 VDD.t2097 VSS 0.018322f
C8746 VDD.t2103 VSS 0.006764f
C8747 VDD.t2099 VSS 0.006764f
C8748 VDD.n270 VSS 0.015166f
C8749 VDD.t2107 VSS 0.021819f
C8750 VDD.t2102 VSS 0.116433f
C8751 VDD.t418 VSS 0.104645f
C8752 VDD.t421 VSS 0.006764f
C8753 VDD.t419 VSS 0.006764f
C8754 VDD.n271 VSS 0.015166f
C8755 VDD.t417 VSS 0.022156f
C8756 VDD.n272 VSS 0.102857f
C8757 VDD.t415 VSS 0.018322f
C8758 VDD.t1901 VSS 0.018322f
C8759 VDD.t826 VSS 0.006764f
C8760 VDD.t848 VSS 0.006764f
C8761 VDD.n273 VSS 0.015166f
C8762 VDD.t414 VSS 0.213738f
C8763 VDD.t1642 VSS 0.214099f
C8764 VDD.t1643 VSS 0.147505f
C8765 VDD.t1644 VSS 0.230818f
C8766 VDD.t1900 VSS 0.230818f
C8767 VDD.t825 VSS 0.116433f
C8768 VDD.t888 VSS 0.227678f
C8769 VDD.t865 VSS 0.103398f
C8770 VDD.t842 VSS 0.006764f
C8771 VDD.t866 VSS 0.006764f
C8772 VDD.n274 VSS 0.015166f
C8773 VDD.t898 VSS 0.018322f
C8774 VDD.t1905 VSS 0.018322f
C8775 VDD.n275 VSS 0.065852f
C8776 VDD.n276 VSS 0.067095f
C8777 VDD.n277 VSS 0.046857f
C8778 VDD.t889 VSS 0.018335f
C8779 VDD.t2109 VSS 0.018322f
C8780 VDD.t2111 VSS 0.006764f
C8781 VDD.t2101 VSS 0.006764f
C8782 VDD.n278 VSS 0.015166f
C8783 VDD.t2114 VSS 0.103398f
C8784 VDD.t2119 VSS 0.018322f
C8785 VDD.t1899 VSS 0.018322f
C8786 VDD.n279 VSS 0.090004f
C8787 VDD.t829 VSS 0.104824f
C8788 VDD.t902 VSS 0.018322f
C8789 VDD.t1978 VSS 0.018313f
C8790 VDD.t1980 VSS 0.006764f
C8791 VDD.t1976 VSS 0.006764f
C8792 VDD.n280 VSS 0.015166f
C8793 VDD.t1974 VSS 0.018884f
C8794 VDD.n281 VSS 0.015731f
C8795 VDD.t1487 VSS 0.018322f
C8796 VDD.t1485 VSS 0.006764f
C8797 VDD.t1483 VSS 0.006764f
C8798 VDD.n282 VSS 0.015166f
C8799 VDD.n283 VSS 0.019803f
C8800 VDD.n284 VSS 0.009459f
C8801 VDD.t1486 VSS 0.227678f
C8802 VDD.t1484 VSS 0.114849f
C8803 VDD.t2096 VSS 0.230818f
C8804 VDD.t171 VSS 0.230818f
C8805 VDD.t172 VSS 0.147505f
C8806 VDD.t170 VSS 0.230818f
C8807 VDD.t1480 VSS 0.227678f
C8808 VDD.t1482 VSS 0.103398f
C8809 VDD.n285 VSS 0.061018f
C8810 VDD.n286 VSS -0.010477f
C8811 VDD.n287 VSS 0.019011f
C8812 VDD.t689 VSS 0.021269f
C8813 VDD.t690 VSS 0.01669f
C8814 VDD.n288 VSS 0.071804f
C8815 VDD.t1655 VSS 0.018322f
C8816 VDD.n289 VSS -0.073356f
C8817 VDD.t1422 VSS 0.006764f
C8818 VDD.t1659 VSS 0.006764f
C8819 VDD.n290 VSS 0.015166f
C8820 VDD.n291 VSS 0.035907f
C8821 VDD.t1510 VSS 0.116433f
C8822 VDD.t1511 VSS 0.006764f
C8823 VDD.t1513 VSS 0.006764f
C8824 VDD.n292 VSS 0.015166f
C8825 VDD.t1519 VSS 0.018322f
C8826 VDD.t340 VSS 0.018322f
C8827 VDD.t336 VSS 0.006764f
C8828 VDD.t342 VSS 0.006764f
C8829 VDD.n293 VSS 0.015166f
C8830 VDD.t338 VSS 0.022391f
C8831 VDD.n294 VSS 0.095048f
C8832 VDD.t1662 VSS 0.116433f
C8833 VDD.t1663 VSS 0.006764f
C8834 VDD.t1426 VSS 0.006764f
C8835 VDD.n295 VSS 0.015166f
C8836 VDD.t1657 VSS 0.018322f
C8837 VDD.t1983 VSS 0.018322f
C8838 VDD.t1985 VSS 0.006764f
C8839 VDD.t1987 VSS 0.006764f
C8840 VDD.n296 VSS 0.015166f
C8841 VDD.t1989 VSS 0.018322f
C8842 VDD.t1942 VSS 0.018422f
C8843 VDD.t1946 VSS 0.006764f
C8844 VDD.t1948 VSS 0.006764f
C8845 VDD.n297 VSS 0.015166f
C8846 VDD.n298 VSS 0.035894f
C8847 VDD.t1941 VSS 0.227678f
C8848 VDD.t1945 VSS 0.103398f
C8849 VDD.t1514 VSS 0.116433f
C8850 VDD.t1505 VSS 0.018322f
C8851 VDD.t1940 VSS 0.018313f
C8852 VDD.n299 VSS 0.051521f
C8853 VDD.n300 VSS 0.059268f
C8854 VDD.t1509 VSS 0.006764f
C8855 VDD.t1515 VSS 0.006764f
C8856 VDD.n301 VSS 0.015166f
C8857 VDD.t1517 VSS 0.018322f
C8858 VDD.t396 VSS 0.018322f
C8859 VDD.n302 VSS 0.046913f
C8860 VDD.t1516 VSS 0.230818f
C8861 VDD.t1590 VSS 0.230818f
C8862 VDD.t1589 VSS 0.147505f
C8863 VDD.t1588 VSS 0.18404f
C8864 VDD.t397 VSS 0.114849f
C8865 VDD.t392 VSS 0.006764f
C8866 VDD.t398 VSS 0.006764f
C8867 VDD.n303 VSS 0.015166f
C8868 VDD.t394 VSS 0.018322f
C8869 VDD.t1424 VSS 0.018322f
C8870 VDD.t1653 VSS 0.006764f
C8871 VDD.t1665 VSS 0.006764f
C8872 VDD.n304 VSS 0.015166f
C8873 VDD.n305 VSS 0.043025f
C8874 VDD.t393 VSS 0.213305f
C8875 VDD.t1423 VSS 0.216226f
C8876 VDD.t1652 VSS 0.104824f
C8877 VDD.t195 VSS 0.230818f
C8878 VDD.t196 VSS 0.147505f
C8879 VDD.t194 VSS 0.230818f
C8880 VDD.t1654 VSS 0.230818f
C8881 VDD.t1664 VSS 0.116433f
C8882 VDD.n306 VSS 0.062021f
C8883 VDD.n307 VSS -0.011488f
C8884 VDD.n308 VSS 0.05616f
C8885 VDD.n309 VSS 0.048865f
C8886 VDD.n310 VSS 0.035907f
C8887 VDD.n311 VSS -0.010928f
C8888 VDD.n312 VSS 0.061018f
C8889 VDD.t391 VSS 0.103398f
C8890 VDD.t395 VSS 0.168918f
C8891 VDD.n313 VSS 0.202202f
C8892 VDD.n314 VSS 0.090004f
C8893 VDD.n315 VSS 0.043025f
C8894 VDD.n316 VSS -0.011488f
C8895 VDD.n317 VSS 0.062021f
C8896 VDD.t1508 VSS 0.104824f
C8897 VDD.t1504 VSS 0.230818f
C8898 VDD.t1939 VSS 0.227678f
C8899 VDD.t1947 VSS 0.114849f
C8900 VDD.n318 VSS 0.061018f
C8901 VDD.n319 VSS -0.010928f
C8902 VDD.n320 VSS 0.134973f
C8903 VDD.n321 VSS 0.141428f
C8904 VDD.n322 VSS 0.041121f
C8905 VDD.t1988 VSS 0.227678f
C8906 VDD.t1984 VSS 0.114849f
C8907 VDD.t1656 VSS 0.230818f
C8908 VDD.t144 VSS 0.230818f
C8909 VDD.t142 VSS 0.147505f
C8910 VDD.t143 VSS 0.230818f
C8911 VDD.t1982 VSS 0.227678f
C8912 VDD.t1986 VSS 0.103398f
C8913 VDD.n323 VSS 0.061018f
C8914 VDD.n324 VSS -0.010718f
C8915 VDD.n325 VSS 0.08647f
C8916 VDD.n326 VSS 0.090838f
C8917 VDD.n327 VSS 0.043025f
C8918 VDD.t1661 VSS 0.022055f
C8919 VDD.n328 VSS -0.011488f
C8920 VDD.n329 VSS 0.062021f
C8921 VDD.t1425 VSS 0.104824f
C8922 VDD.t1660 VSS 0.283776f
C8923 VDD.t337 VSS 0.283492f
C8924 VDD.t335 VSS 0.116235f
C8925 VDD.t1518 VSS 0.230818f
C8926 VDD.t2017 VSS 0.230818f
C8927 VDD.t2018 VSS 0.147505f
C8928 VDD.t2016 VSS 0.214099f
C8929 VDD.t339 VSS 0.213738f
C8930 VDD.t341 VSS 0.104645f
C8931 VDD.n330 VSS 0.061895f
C8932 VDD.n331 VSS -0.010623f
C8933 VDD.n332 VSS 0.086535f
C8934 VDD.n333 VSS 0.089368f
C8935 VDD.n334 VSS 0.043025f
C8936 VDD.t1507 VSS 0.018322f
C8937 VDD.t1667 VSS 0.018322f
C8938 VDD.n335 VSS 0.050861f
C8939 VDD.n336 VSS 0.058884f
C8940 VDD.n337 VSS -0.011488f
C8941 VDD.n338 VSS 0.062021f
C8942 VDD.t1512 VSS 0.104824f
C8943 VDD.t1506 VSS 0.222623f
C8944 VDD.t1666 VSS 0.222623f
C8945 VDD.t1421 VSS 0.116433f
C8946 VDD.t1668 VSS 0.230818f
C8947 VDD.t1658 VSS 0.104824f
C8948 VDD.n339 VSS 0.062021f
C8949 VDD.n340 VSS -0.010928f
C8950 VDD.t1669 VSS 0.018342f
C8951 VDD.n341 VSS 0.0446f
C8952 VDD.n342 VSS -0.174353f
C8953 VDD.n343 VSS 0.071681f
C8954 VDD.t688 VSS 0.619833f
C8955 VDD.t1981 VSS 0.375016f
C8956 VDD.t1464 VSS 0.619833f
C8957 VDD.t1468 VSS 0.219141f
C8958 VDD.n344 VSS 0.189733f
C8959 VDD.n345 VSS -0.002704f
C8960 VDD.t1476 VSS 0.021269f
C8961 VDD.t1465 VSS 0.01669f
C8962 VDD.n346 VSS 0.070928f
C8963 VDD.t1469 VSS 0.006764f
C8964 VDD.t1472 VSS 0.006764f
C8965 VDD.n347 VSS 0.013528f
C8966 VDD.n348 VSS 0.037088f
C8967 VDD.n349 VSS 0.05886f
C8968 VDD.n350 VSS 0.142084f
C8969 VDD.n351 VSS 0.033784f
C8970 VDD.n352 VSS 0.007227f
C8971 VDD.n353 VSS 0.018257f
C8972 VDD.n354 VSS 0.027316f
C8973 VDD.n355 VSS 0.042731f
C8974 VDD.n356 VSS 0.137686f
C8975 VDD.n357 VSS 0.102628f
C8976 VDD.t1973 VSS 0.227678f
C8977 VDD.t1979 VSS 0.103398f
C8978 VDD.t901 VSS 0.230818f
C8979 VDD.t1977 VSS 0.227678f
C8980 VDD.t1975 VSS 0.114849f
C8981 VDD.n358 VSS 0.061018f
C8982 VDD.n359 VSS -0.010928f
C8983 VDD.n360 VSS 0.035894f
C8984 VDD.n361 VSS 0.051521f
C8985 VDD.n362 VSS 0.059268f
C8986 VDD.t830 VSS 0.006764f
C8987 VDD.t872 VSS 0.006764f
C8988 VDD.n363 VSS 0.015166f
C8989 VDD.n364 VSS 0.043025f
C8990 VDD.n365 VSS -0.011488f
C8991 VDD.n366 VSS 0.062021f
C8992 VDD.t871 VSS 0.116433f
C8993 VDD.t1898 VSS 0.230818f
C8994 VDD.t1933 VSS 0.230818f
C8995 VDD.t1932 VSS 0.147505f
C8996 VDD.t1934 VSS 0.18404f
C8997 VDD.t2118 VSS 0.168918f
C8998 VDD.n367 VSS 0.202202f
C8999 VDD.n368 VSS 0.046913f
C9000 VDD.t2115 VSS 0.006764f
C9001 VDD.t2113 VSS 0.006764f
C9002 VDD.n369 VSS 0.015166f
C9003 VDD.t2117 VSS 0.018322f
C9004 VDD.t2105 VSS 0.018322f
C9005 VDD.n370 VSS 0.05616f
C9006 VDD.n371 VSS 0.048865f
C9007 VDD.n372 VSS 0.035907f
C9008 VDD.n373 VSS -0.010928f
C9009 VDD.n374 VSS 0.061018f
C9010 VDD.t2112 VSS 0.114849f
C9011 VDD.t2116 VSS 0.213305f
C9012 VDD.t2104 VSS 0.216226f
C9013 VDD.t2110 VSS 0.104824f
C9014 VDD.t318 VSS 0.230818f
C9015 VDD.t316 VSS 0.147505f
C9016 VDD.t317 VSS 0.230818f
C9017 VDD.t2108 VSS 0.230818f
C9018 VDD.t2100 VSS 0.116433f
C9019 VDD.n375 VSS 0.062021f
C9020 VDD.n376 VSS -0.011488f
C9021 VDD.n377 VSS 0.043025f
C9022 VDD.n378 VSS 0.212659f
C9023 VDD.t468 VSS 0.006764f
C9024 VDD.t652 VSS 0.006764f
C9025 VDD.n379 VSS 0.029826f
C9026 VDD.t480 VSS 0.006764f
C9027 VDD.t1874 VSS 0.006764f
C9028 VDD.n380 VSS 0.013528f
C9029 VDD.n381 VSS 0.039293f
C9030 VDD.t469 VSS 0.006764f
C9031 VDD.t651 VSS 0.006764f
C9032 VDD.n382 VSS 0.029015f
C9033 VDD.n383 VSS 0.03765f
C9034 VDD.t479 VSS 0.006764f
C9035 VDD.t1875 VSS 0.006764f
C9036 VDD.n384 VSS 0.013528f
C9037 VDD.n385 VSS 0.008042f
C9038 VDD.n386 VSS 0.074425f
C9039 VDD.t208 VSS 0.470588f
C9040 VDD.t478 VSS 0.331315f
C9041 VDD.t1873 VSS 0.185802f
C9042 VDD.t699 VSS 0.400006f
C9043 VDD.t1617 VSS 0.197636f
C9044 VDD.t1619 VSS 0.006764f
C9045 VDD.t701 VSS 0.006764f
C9046 VDD.n387 VSS 0.029826f
C9047 VDD.t765 VSS 0.006764f
C9048 VDD.t1419 VSS 0.006764f
C9049 VDD.n388 VSS 0.013528f
C9050 VDD.n389 VSS 0.039293f
C9051 VDD.t1618 VSS 0.006764f
C9052 VDD.t700 VSS 0.006764f
C9053 VDD.n390 VSS 0.029015f
C9054 VDD.n391 VSS 0.03765f
C9055 VDD.t766 VSS 0.006764f
C9056 VDD.t1420 VSS 0.006764f
C9057 VDD.n392 VSS 0.013528f
C9058 VDD.n393 VSS 0.008042f
C9059 VDD.t216 VSS 0.027971f
C9060 VDD.n394 VSS 0.044989f
C9061 VDD.t218 VSS 0.034731f
C9062 VDD.n395 VSS 0.04544f
C9063 VDD.n396 VSS 0.027244f
C9064 VDD.t1244 VSS 0.006764f
C9065 VDD.t1250 VSS 0.006764f
C9066 VDD.n397 VSS 0.018548f
C9067 VDD.t1936 VSS 0.006764f
C9068 VDD.t1935 VSS 0.006764f
C9069 VDD.n398 VSS 0.013528f
C9070 VDD.n399 VSS 0.032136f
C9071 VDD.t1385 VSS 0.227678f
C9072 VDD.t1393 VSS 0.114849f
C9073 VDD.t1386 VSS 0.027262f
C9074 VDD.t1394 VSS 0.006764f
C9075 VDD.t1408 VSS 0.006764f
C9076 VDD.n400 VSS 0.015166f
C9077 VDD.t1390 VSS 0.027282f
C9078 VDD.n401 VSS 0.038369f
C9079 VDD.n402 VSS 0.078978f
C9080 VDD.n403 VSS -0.010365f
C9081 VDD.n404 VSS 0.061018f
C9082 VDD.t1407 VSS 0.103398f
C9083 VDD.t1389 VSS 0.229878f
C9084 VDD.t562 VSS 0.409363f
C9085 VDD.t563 VSS 0.259137f
C9086 VDD.t1243 VSS 0.259137f
C9087 VDD.t1249 VSS 0.310025f
C9088 VDD.t1236 VSS 0.103398f
C9089 VDD.t1240 VSS 0.3011f
C9090 VDD.t2046 VSS 0.3011f
C9091 VDD.t2042 VSS 0.114849f
C9092 VDD.t1853 VSS 0.146509f
C9093 VDD.t2041 VSS 0.018322f
C9094 VDD.t2043 VSS 0.006764f
C9095 VDD.t2057 VSS 0.006764f
C9096 VDD.n405 VSS 0.015166f
C9097 VDD.t2047 VSS 0.018322f
C9098 VDD.t1241 VSS 0.018322f
C9099 VDD.t1226 VSS 0.006764f
C9100 VDD.t1237 VSS 0.006764f
C9101 VDD.n406 VSS 0.015166f
C9102 VDD.t1246 VSS 0.034094f
C9103 VDD.n407 VSS 0.042374f
C9104 VDD.n408 VSS 0.030866f
C9105 VDD.n409 VSS 0.030866f
C9106 VDD.n410 VSS 0.02436f
C9107 VDD.n411 VSS 0.031399f
C9108 VDD.t1849 VSS 0.006764f
C9109 VDD.t1857 VSS 0.006764f
C9110 VDD.n412 VSS 0.018548f
C9111 VDD.t23 VSS 0.006764f
C9112 VDD.t25 VSS 0.006764f
C9113 VDD.n413 VSS 0.013528f
C9114 VDD.n414 VSS 0.031682f
C9115 VDD.t1854 VSS 0.028156f
C9116 VDD.t1844 VSS 0.006764f
C9117 VDD.t1846 VSS 0.006764f
C9118 VDD.n415 VSS 0.015166f
C9119 VDD.t1852 VSS 0.018322f
C9120 VDD.t2081 VSS 0.018322f
C9121 VDD.t2085 VSS 0.006764f
C9122 VDD.t2091 VSS 0.006764f
C9123 VDD.n416 VSS 0.015166f
C9124 VDD.t2079 VSS 0.027282f
C9125 VDD.n417 VSS 0.042575f
C9126 VDD.n418 VSS 0.029938f
C9127 VDD.n419 VSS 0.029938f
C9128 VDD.n420 VSS 0.025565f
C9129 VDD.n421 VSS 0.022589f
C9130 VDD.n422 VSS 0.01248f
C9131 VDD.n423 VSS 0.105693f
C9132 VDD.t1843 VSS 0.114849f
C9133 VDD.t2090 VSS 0.103398f
C9134 VDD.t1681 VSS 0.006764f
C9135 VDD.t1695 VSS 0.006764f
C9136 VDD.n424 VSS 0.018548f
C9137 VDD.t1634 VSS 0.006764f
C9138 VDD.t1636 VSS 0.006764f
C9139 VDD.n425 VSS 0.013528f
C9140 VDD.n426 VSS 0.032136f
C9141 VDD.t2078 VSS 0.229878f
C9142 VDD.t560 VSS 0.409363f
C9143 VDD.t561 VSS 0.259137f
C9144 VDD.t1633 VSS 0.259137f
C9145 VDD.t1635 VSS 0.310025f
C9146 VDD.t1693 VSS 0.227678f
C9147 VDD.t1686 VSS 0.103398f
C9148 VDD.t1689 VSS 0.035637f
C9149 VDD.t1677 VSS 0.006764f
C9150 VDD.t1687 VSS 0.006764f
C9151 VDD.n427 VSS 0.015166f
C9152 VDD.t1694 VSS 0.03306f
C9153 VDD.n428 VSS 0.026295f
C9154 VDD.n429 VSS 0.019667f
C9155 VDD.t2136 VSS 0.018322f
C9156 VDD.t2126 VSS 0.006764f
C9157 VDD.t2129 VSS 0.006764f
C9158 VDD.n430 VSS 0.015166f
C9159 VDD.n431 VSS 0.045731f
C9160 VDD.t769 VSS 0.310025f
C9161 VDD.t2132 VSS 0.006764f
C9162 VDD.t2146 VSS 0.006764f
C9163 VDD.n432 VSS 0.018548f
C9164 VDD.t768 VSS 0.006764f
C9165 VDD.t770 VSS 0.006764f
C9166 VDD.n433 VSS 0.013528f
C9167 VDD.n434 VSS 0.032136f
C9168 VDD.t2031 VSS 0.018322f
C9169 VDD.t2033 VSS 0.006764f
C9170 VDD.t2035 VSS 0.006764f
C9171 VDD.n435 VSS 0.015166f
C9172 VDD.n436 VSS 0.046076f
C9173 VDD.t1427 VSS 0.114849f
C9174 VDD.t1428 VSS 0.006764f
C9175 VDD.t1435 VSS 0.006764f
C9176 VDD.n437 VSS 0.015166f
C9177 VDD.t1455 VSS 0.018294f
C9178 VDD.t1440 VSS 0.006764f
C9179 VDD.t1456 VSS 0.006764f
C9180 VDD.n438 VSS 0.018548f
C9181 VDD.t299 VSS 0.006764f
C9182 VDD.t301 VSS 0.006764f
C9183 VDD.n439 VSS 0.013528f
C9184 VDD.n440 VSS 0.032136f
C9185 VDD.n441 VSS 0.078479f
C9186 VDD.t1959 VSS 0.114849f
C9187 VDD.t1960 VSS 0.006764f
C9188 VDD.t1968 VSS 0.006764f
C9189 VDD.n442 VSS 0.015166f
C9190 VDD.t1956 VSS 0.018322f
C9191 VDD.t1997 VSS 0.018322f
C9192 VDD.t2004 VSS 0.006764f
C9193 VDD.t2011 VSS 0.006764f
C9194 VDD.n443 VSS 0.015166f
C9195 VDD.n444 VSS 0.045731f
C9196 VDD.t598 VSS 0.310025f
C9197 VDD.t1995 VSS 0.006764f
C9198 VDD.t2001 VSS 0.006764f
C9199 VDD.n445 VSS 0.018548f
C9200 VDD.t601 VSS 0.006764f
C9201 VDD.t599 VSS 0.006764f
C9202 VDD.n446 VSS 0.013528f
C9203 VDD.n447 VSS 0.032136f
C9204 VDD.t1814 VSS 0.018322f
C9205 VDD.t1820 VSS 0.006764f
C9206 VDD.t1828 VSS 0.006764f
C9207 VDD.n448 VSS 0.015166f
C9208 VDD.n449 VSS 0.046076f
C9209 VDD.t1544 VSS 0.114849f
C9210 VDD.t1545 VSS 0.006764f
C9211 VDD.t1523 VSS 0.006764f
C9212 VDD.n450 VSS 0.015166f
C9213 VDD.t1528 VSS 0.018294f
C9214 VDD.t1524 VSS 0.006764f
C9215 VDD.t1529 VSS 0.006764f
C9216 VDD.n451 VSS 0.018548f
C9217 VDD.t239 VSS 0.006764f
C9218 VDD.t237 VSS 0.006764f
C9219 VDD.n452 VSS 0.013528f
C9220 VDD.n453 VSS 0.032109f
C9221 VDD.n454 VSS 0.07921f
C9222 VDD.t1177 VSS 0.114849f
C9223 VDD.t1178 VSS 0.006764f
C9224 VDD.t1182 VSS 0.006764f
C9225 VDD.n455 VSS 0.015166f
C9226 VDD.t1170 VSS 0.018322f
C9227 VDD.t551 VSS 0.018157f
C9228 VDD.t104 VSS 0.006764f
C9229 VDD.t553 VSS 0.006764f
C9230 VDD.n456 VSS 0.014917f
C9231 VDD.t464 VSS 0.006764f
C9232 VDD.t106 VSS 0.006764f
C9233 VDD.n457 VSS 0.014917f
C9234 VDD.t466 VSS 0.018157f
C9235 VDD.t1920 VSS 0.018157f
C9236 VDD.t912 VSS 0.006764f
C9237 VDD.t1922 VSS 0.006764f
C9238 VDD.n458 VSS 0.014917f
C9239 VDD.t1609 VSS 0.006764f
C9240 VDD.t910 VSS 0.006764f
C9241 VDD.n459 VSS 0.014917f
C9242 VDD.t1607 VSS 0.018157f
C9243 VDD.t1803 VSS 0.018322f
C9244 VDD.t1809 VSS 0.006764f
C9245 VDD.t1783 VSS 0.006764f
C9246 VDD.n460 VSS 0.015166f
C9247 VDD.t1794 VSS 0.022873f
C9248 VDD.n461 VSS 0.07781f
C9249 VDD.t1793 VSS 0.227678f
C9250 VDD.t1808 VSS 0.114849f
C9251 VDD.t1169 VSS 0.278568f
C9252 VDD.t550 VSS 0.262997f
C9253 VDD.t552 VSS 0.136969f
C9254 VDD.t103 VSS 0.136969f
C9255 VDD.t105 VSS 0.136969f
C9256 VDD.t463 VSS 0.136969f
C9257 VDD.t465 VSS 0.242866f
C9258 VDD.t1919 VSS 0.242866f
C9259 VDD.t1921 VSS 0.136969f
C9260 VDD.t911 VSS 0.136969f
C9261 VDD.t909 VSS 0.136969f
C9262 VDD.t1608 VSS 0.136969f
C9263 VDD.t1606 VSS 0.255519f
C9264 VDD.t1802 VSS 0.270827f
C9265 VDD.t1782 VSS 0.103398f
C9266 VDD.n462 VSS 0.061018f
C9267 VDD.n463 VSS -0.010928f
C9268 VDD.n464 VSS 0.061147f
C9269 VDD.n465 VSS 0.058012f
C9270 VDD.n466 VSS 0.0563f
C9271 VDD.n467 VSS 0.034926f
C9272 VDD.n468 VSS 0.056306f
C9273 VDD.n469 VSS 0.056306f
C9274 VDD.n470 VSS 0.0563f
C9275 VDD.n471 VSS 0.034926f
C9276 VDD.n472 VSS 0.058754f
C9277 VDD.n473 VSS 0.072611f
C9278 VDD.n474 VSS 0.046076f
C9279 VDD.t1188 VSS 0.018322f
C9280 VDD.n475 VSS 0.103126f
C9281 VDD.n476 VSS -0.010519f
C9282 VDD.n477 VSS 0.061018f
C9283 VDD.t1181 VSS 0.103398f
C9284 VDD.t1187 VSS 0.229878f
C9285 VDD.t549 VSS 0.409363f
C9286 VDD.t548 VSS 0.259137f
C9287 VDD.t238 VSS 0.259137f
C9288 VDD.t236 VSS 0.310025f
C9289 VDD.t1527 VSS 0.146509f
C9290 VDD.n478 VSS 0.193277f
C9291 VDD.n479 VSS 0.017772f
C9292 VDD.n480 VSS 0.058631f
C9293 VDD.n481 VSS 0.045731f
C9294 VDD.t1538 VSS 0.018322f
C9295 VDD.t1834 VSS 0.018322f
C9296 VDD.n482 VSS 0.077762f
C9297 VDD.n483 VSS 0.07543f
C9298 VDD.n484 VSS -0.01053f
C9299 VDD.n485 VSS 0.061018f
C9300 VDD.t1522 VSS 0.103398f
C9301 VDD.t1537 VSS 0.321982f
C9302 VDD.t1833 VSS 0.321982f
C9303 VDD.t1819 VSS 0.114849f
C9304 VDD.t600 VSS 0.259137f
C9305 VDD.t1621 VSS 0.259137f
C9306 VDD.t1620 VSS 0.409363f
C9307 VDD.t1813 VSS 0.229878f
C9308 VDD.t1827 VSS 0.103398f
C9309 VDD.n486 VSS 0.061018f
C9310 VDD.n487 VSS -0.010519f
C9311 VDD.n488 VSS 0.102669f
C9312 VDD.n489 VSS 0.078479f
C9313 VDD.t1999 VSS 0.018294f
C9314 VDD.n490 VSS 0.058631f
C9315 VDD.n491 VSS 0.017781f
C9316 VDD.n492 VSS 0.193277f
C9317 VDD.t1998 VSS 0.146509f
C9318 VDD.t2003 VSS 0.114849f
C9319 VDD.t1955 VSS 0.266747f
C9320 VDD.t1996 VSS 0.266747f
C9321 VDD.t2010 VSS 0.103398f
C9322 VDD.n493 VSS 0.061018f
C9323 VDD.n494 VSS -0.01053f
C9324 VDD.n495 VSS 0.073705f
C9325 VDD.n496 VSS 0.075269f
C9326 VDD.n497 VSS 0.046076f
C9327 VDD.t1954 VSS 0.018322f
C9328 VDD.n498 VSS 0.102669f
C9329 VDD.n499 VSS -0.010519f
C9330 VDD.n500 VSS 0.061018f
C9331 VDD.t1967 VSS 0.103398f
C9332 VDD.t1953 VSS 0.229878f
C9333 VDD.t735 VSS 0.409363f
C9334 VDD.t734 VSS 0.259137f
C9335 VDD.t298 VSS 0.259137f
C9336 VDD.t300 VSS 0.310025f
C9337 VDD.t1454 VSS 0.146509f
C9338 VDD.n501 VSS 0.193277f
C9339 VDD.n502 VSS 0.017781f
C9340 VDD.n503 VSS 0.058631f
C9341 VDD.n504 VSS 0.045731f
C9342 VDD.t1452 VSS 0.018322f
C9343 VDD.t2029 VSS 0.018322f
C9344 VDD.n505 VSS 0.075804f
C9345 VDD.n506 VSS 0.074239f
C9346 VDD.n507 VSS -0.01053f
C9347 VDD.n508 VSS 0.061018f
C9348 VDD.t1434 VSS 0.103398f
C9349 VDD.t1451 VSS 0.269441f
C9350 VDD.t2028 VSS 0.269441f
C9351 VDD.t2032 VSS 0.114849f
C9352 VDD.t767 VSS 0.259137f
C9353 VDD.t773 VSS 0.259137f
C9354 VDD.t774 VSS 0.409363f
C9355 VDD.t2030 VSS 0.229878f
C9356 VDD.t2034 VSS 0.103398f
C9357 VDD.n509 VSS 0.061018f
C9358 VDD.n510 VSS -0.010519f
C9359 VDD.n511 VSS 0.102669f
C9360 VDD.n512 VSS 0.078479f
C9361 VDD.t2134 VSS 0.018294f
C9362 VDD.n513 VSS 0.058631f
C9363 VDD.n514 VSS 0.017781f
C9364 VDD.n515 VSS 0.193277f
C9365 VDD.t2133 VSS 0.146509f
C9366 VDD.t2125 VSS 0.114849f
C9367 VDD.t2135 VSS 0.227678f
C9368 VDD.t2128 VSS 0.103398f
C9369 VDD.n516 VSS 0.061018f
C9370 VDD.n517 VSS -0.01053f
C9371 VDD.n518 VSS 0.47366f
C9372 VDD.n519 VSS 0.18346f
C9373 VDD.n520 VSS 0.020137f
C9374 VDD.n521 VSS 0.061018f
C9375 VDD.t1676 VSS 0.114849f
C9376 VDD.t1688 VSS 0.146509f
C9377 VDD.n522 VSS 0.193277f
C9378 VDD.n523 VSS 0.013114f
C9379 VDD.n524 VSS 0.102239f
C9380 VDD.n525 VSS 0.058379f
C9381 VDD.n526 VSS 0.061018f
C9382 VDD.t2084 VSS 0.114849f
C9383 VDD.t2080 VSS 0.269441f
C9384 VDD.t1851 VSS 0.269441f
C9385 VDD.t1845 VSS 0.103398f
C9386 VDD.n527 VSS 0.061018f
C9387 VDD.n528 VSS 0.020137f
C9388 VDD.n529 VSS 0.035024f
C9389 VDD.n530 VSS 0.193277f
C9390 VDD.t24 VSS 0.310025f
C9391 VDD.t22 VSS 0.259137f
C9392 VDD.t110 VSS 0.259137f
C9393 VDD.t109 VSS 0.409363f
C9394 VDD.t2040 VSS 0.229878f
C9395 VDD.t2056 VSS 0.103398f
C9396 VDD.n531 VSS 0.061018f
C9397 VDD.n532 VSS 0.063729f
C9398 VDD.n533 VSS 0.020137f
C9399 VDD.n534 VSS 0.061018f
C9400 VDD.t1225 VSS 0.114849f
C9401 VDD.t1245 VSS 0.146509f
C9402 VDD.n535 VSS 0.193277f
C9403 VDD.n536 VSS 0.013114f
C9404 VDD.n537 VSS 0.099889f
C9405 VDD.n538 VSS 0.075906f
C9406 VDD.n539 VSS 0.021675f
C9407 VDD.n540 VSS 0.099614f
C9408 VDD.t1418 VSS 0.185802f
C9409 VDD.t764 VSS 0.331315f
C9410 VDD.t217 VSS 0.835558f
C9411 VDD.t650 VSS 0.760366f
C9412 VDD.t467 VSS 0.197636f
C9413 VDD.n541 VSS 0.099614f
C9414 VDD.n542 VSS 0.065197f
C9415 VDD.n543 VSS 0.027244f
C9416 VDD.n544 VSS 0.044892f
C9417 VDD.t207 VSS 0.027971f
C9418 VDD.t209 VSS 0.034731f
C9419 VDD.n545 VSS 0.043291f
C9420 VDD.n546 VSS 0.033552f
C9421 VDD.n547 VSS 1.71725f
C9422 VDD.n548 VSS 0.056179f
C9423 VDD.n549 VSS -0.010488f
C9424 VDD.n550 VSS 0.061018f
C9425 VDD.t841 VSS 0.114849f
C9426 VDD.t897 VSS 0.219653f
C9427 VDD.t1904 VSS 0.222676f
C9428 VDD.t847 VSS 0.104824f
C9429 VDD.n551 VSS 0.062021f
C9430 VDD.n552 VSS -0.011456f
C9431 VDD.n553 VSS 0.046651f
C9432 VDD.n554 VSS 0.109145f
C9433 VDD.n555 VSS 0.106936f
C9434 VDD.n556 VSS -0.010468f
C9435 VDD.n557 VSS 0.061895f
C9436 VDD.t420 VSS 0.116235f
C9437 VDD.t416 VSS 0.283492f
C9438 VDD.t2106 VSS 0.283776f
C9439 VDD.t2098 VSS 0.104824f
C9440 VDD.n558 VSS 0.062021f
C9441 VDD.n559 VSS -0.011434f
C9442 VDD.n560 VSS 0.048981f
C9443 VDD.n561 VSS 0.09878f
C9444 VDD.n562 VSS 0.226065f
C9445 VDD.n563 VSS 0.178553f
C9446 VDD.n564 VSS 0.044459f
C9447 VDD.n565 VSS 0.059268f
C9448 VDD.t1491 VSS 0.006764f
C9449 VDD.t1497 VSS 0.006764f
C9450 VDD.n566 VSS 0.015166f
C9451 VDD.t1489 VSS 0.018322f
C9452 VDD.t1008 VSS 0.018322f
C9453 VDD.n567 VSS 0.046913f
C9454 VDD.t1488 VSS 0.230818f
C9455 VDD.t616 VSS 0.230818f
C9456 VDD.t615 VSS 0.147505f
C9457 VDD.t617 VSS 0.18404f
C9458 VDD.t1005 VSS 0.114849f
C9459 VDD.t1004 VSS 0.006764f
C9460 VDD.t1006 VSS 0.006764f
C9461 VDD.n568 VSS 0.015166f
C9462 VDD.t1010 VSS 0.018322f
C9463 VDD.t836 VSS 0.018322f
C9464 VDD.t878 VSS 0.006764f
C9465 VDD.t1903 VSS 0.006764f
C9466 VDD.n569 VSS 0.015166f
C9467 VDD.n570 VSS 0.043025f
C9468 VDD.t1009 VSS 0.213305f
C9469 VDD.t835 VSS 0.216226f
C9470 VDD.t877 VSS 0.104824f
C9471 VDD.t472 VSS 0.230818f
C9472 VDD.t470 VSS 0.147505f
C9473 VDD.t471 VSS 0.230818f
C9474 VDD.t831 VSS 0.230818f
C9475 VDD.t1902 VSS 0.116433f
C9476 VDD.n571 VSS 0.062021f
C9477 VDD.n572 VSS -0.011488f
C9478 VDD.n573 VSS 0.05616f
C9479 VDD.n574 VSS 0.048865f
C9480 VDD.n575 VSS 0.035907f
C9481 VDD.n576 VSS -0.010928f
C9482 VDD.n577 VSS 0.061018f
C9483 VDD.t1003 VSS 0.103398f
C9484 VDD.t1007 VSS 0.168918f
C9485 VDD.n578 VSS 0.202202f
C9486 VDD.n579 VSS 0.090004f
C9487 VDD.n580 VSS 0.043025f
C9488 VDD.n581 VSS -0.011488f
C9489 VDD.n582 VSS 0.062021f
C9490 VDD.t1490 VSS 0.104824f
C9491 VDD.t1502 VSS 0.230818f
C9492 VDD.t2060 VSS 0.227678f
C9493 VDD.t2067 VSS 0.114849f
C9494 VDD.n583 VSS 0.061018f
C9495 VDD.n584 VSS -0.010928f
C9496 VDD.n585 VSS 0.139296f
C9497 VDD.n586 VSS 0.154135f
C9498 VDD.t849 VSS 0.114849f
C9499 VDD.t850 VSS 0.006764f
C9500 VDD.t816 VSS 0.006764f
C9501 VDD.n587 VSS 0.015166f
C9502 VDD.n588 VSS 0.035907f
C9503 VDD.t854 VSS 0.018342f
C9504 VDD.t840 VSS 0.018322f
C9505 VDD.t874 VSS 0.006764f
C9506 VDD.t820 VSS 0.006764f
C9507 VDD.n589 VSS 0.015166f
C9508 VDD.t792 VSS 0.103398f
C9509 VDD.t789 VSS 0.018322f
C9510 VDD.t964 VSS 0.018322f
C9511 VDD.n590 VSS 0.090004f
C9512 VDD.t959 VSS 0.104824f
C9513 VDD.t970 VSS 0.018322f
C9514 VDD.t1467 VSS 0.018313f
C9515 VDD.t1460 VSS 0.006764f
C9516 VDD.t1462 VSS 0.006764f
C9517 VDD.n591 VSS 0.015166f
C9518 VDD.t1471 VSS 0.018422f
C9519 VDD.t1786 VSS 0.006764f
C9520 VDD.t1799 VSS 0.006764f
C9521 VDD.n592 VSS 0.01683f
C9522 VDD.t1777 VSS 0.006764f
C9523 VDD.t1785 VSS 0.006764f
C9524 VDD.n593 VSS 0.013528f
C9525 VDD.n594 VSS 0.027737f
C9526 VDD.n595 VSS 0.015175f
C9527 VDD.t1811 VSS 0.214331f
C9528 VDD.t1795 VSS 0.136969f
C9529 VDD.t1937 VSS 0.136969f
C9530 VDD.t1943 VSS 0.136969f
C9531 VDD.t925 VSS 0.136969f
C9532 VDD.t923 VSS 0.141408f
C9533 VDD.t381 VSS 0.619833f
C9534 VDD.t400 VSS 0.375016f
C9535 VDD.t383 VSS 0.021269f
C9536 VDD.t382 VSS 0.01669f
C9537 VDD.n596 VSS 0.084502f
C9538 VDD.t614 VSS 0.021269f
C9539 VDD.t612 VSS 0.01669f
C9540 VDD.n597 VSS 0.070928f
C9541 VDD.t613 VSS 0.006764f
C9542 VDD.t611 VSS 0.006764f
C9543 VDD.n598 VSS 0.013528f
C9544 VDD.n599 VSS 0.036172f
C9545 VDD.t590 VSS 0.018157f
C9546 VDD.t588 VSS 0.006764f
C9547 VDD.t1150 VSS 0.006764f
C9548 VDD.n600 VSS 0.014917f
C9549 VDD.t1152 VSS 0.006764f
C9550 VDD.t705 VSS 0.006764f
C9551 VDD.n601 VSS 0.014917f
C9552 VDD.t703 VSS 0.018157f
C9553 VDD.t1561 VSS 0.018322f
C9554 VDD.n602 VSS 0.071416f
C9555 VDD.t88 VSS 0.021269f
C9556 VDD.t87 VSS 0.01669f
C9557 VDD.n603 VSS 0.075369f
C9558 VDD.t1475 VSS 0.021269f
C9559 VDD.t1463 VSS 0.01669f
C9560 VDD.n604 VSS 0.070928f
C9561 VDD.t1474 VSS 0.006764f
C9562 VDD.t1458 VSS 0.006764f
C9563 VDD.n605 VSS 0.013528f
C9564 VDD.n606 VSS 0.044529f
C9565 VDD.t2064 VSS 0.571907f
C9566 VDD.t30 VSS 0.112529f
C9567 VDD.t1040 VSS 0.126155f
C9568 VDD.t677 VSS 0.018322f
C9569 VDD.n607 VSS 0.046913f
C9570 VDD.t683 VSS 0.006764f
C9571 VDD.t679 VSS 0.006764f
C9572 VDD.n608 VSS 0.015166f
C9573 VDD.t1041 VSS 0.01979f
C9574 VDD.t1071 VSS 0.01669f
C9575 VDD.n609 VSS 0.046329f
C9576 VDD.n610 VSS 0.033014f
C9577 VDD.t681 VSS 0.018322f
C9578 VDD.t887 VSS 0.018322f
C9579 VDD.t280 VSS 0.469716f
C9580 VDD.t1089 VSS 1.03797f
C9581 VDD.t1135 VSS 0.214331f
C9582 VDD.t1052 VSS 0.136969f
C9583 VDD.t2074 VSS 0.136969f
C9584 VDD.t2076 VSS 0.136969f
C9585 VDD.t556 VSS 0.136969f
C9586 VDD.t554 VSS 0.141408f
C9587 VDD.t128 VSS 0.109612f
C9588 VDD.t130 VSS 0.134227f
C9589 VDD.t675 VSS 0.021269f
C9590 VDD.t672 VSS 0.01669f
C9591 VDD.n611 VSS 0.070928f
C9592 VDD.t674 VSS 0.006764f
C9593 VDD.t673 VSS 0.006764f
C9594 VDD.n612 VSS 0.013528f
C9595 VDD.n613 VSS 0.036172f
C9596 VDD.t281 VSS 0.018157f
C9597 VDD.t941 VSS 0.006764f
C9598 VDD.t282 VSS 0.006764f
C9599 VDD.n614 VSS 0.014917f
C9600 VDD.t1640 VSS 0.006764f
C9601 VDD.t940 VSS 0.006764f
C9602 VDD.n615 VSS 0.014917f
C9603 VDD.t1070 VSS 0.006764f
C9604 VDD.t1090 VSS 0.006764f
C9605 VDD.n616 VSS 0.01683f
C9606 VDD.t1106 VSS 0.006764f
C9607 VDD.t1115 VSS 0.006764f
C9608 VDD.n617 VSS 0.013528f
C9609 VDD.n618 VSS 0.02771f
C9610 VDD.n619 VSS 0.015251f
C9611 VDD.n620 VSS 0.010816f
C9612 VDD.n621 VSS 0.034081f
C9613 VDD.t678 VSS 0.175608f
C9614 VDD.n622 VSS 0.188728f
C9615 VDD.t1069 VSS 0.071656f
C9616 VDD.t680 VSS 0.209922f
C9617 VDD.n623 VSS 0.188728f
C9618 VDD.n624 VSS 0.016505f
C9619 VDD.t1641 VSS 0.018217f
C9620 VDD.n625 VSS 0.038117f
C9621 VDD.t1136 VSS 0.018316f
C9622 VDD.t1053 VSS 0.006764f
C9623 VDD.t2075 VSS 0.006764f
C9624 VDD.n626 VSS 0.014917f
C9625 VDD.t2077 VSS 0.006764f
C9626 VDD.t557 VSS 0.006764f
C9627 VDD.n627 VSS 0.014917f
C9628 VDD.t555 VSS 0.022409f
C9629 VDD.n628 VSS 0.096335f
C9630 VDD.n629 VSS 0.033732f
C9631 VDD.n630 VSS 0.096908f
C9632 VDD.n631 VSS 0.072642f
C9633 VDD.n632 VSS 0.033732f
C9634 VDD.n633 VSS 0.0563f
C9635 VDD.n634 VSS 0.056289f
C9636 VDD.n635 VSS 0.032472f
C9637 VDD.t132 VSS 0.021269f
C9638 VDD.t133 VSS 0.01669f
C9639 VDD.n636 VSS 0.068817f
C9640 VDD.t1200 VSS 0.017784f
C9641 VDD.t1203 VSS 0.006764f
C9642 VDD.t533 VSS 0.006764f
C9643 VDD.n637 VSS 0.020425f
C9644 VDD.n638 VSS 0.059702f
C9645 VDD.t532 VSS 0.01669f
C9646 VDD.n639 VSS 0.017903f
C9647 VDD.t528 VSS 0.006764f
C9648 VDD.t530 VSS 0.006764f
C9649 VDD.n640 VSS 0.020425f
C9650 VDD.n641 VSS 0.039154f
C9651 VDD.t707 VSS 0.047077f
C9652 VDD.t709 VSS 0.006764f
C9653 VDD.t943 VSS 0.006764f
C9654 VDD.n642 VSS 0.013528f
C9655 VDD.n643 VSS 0.057677f
C9656 VDD.t944 VSS 0.01669f
C9657 VDD.n644 VSS 0.026665f
C9658 VDD.t1585 VSS 0.018157f
C9659 VDD.n645 VSS 0.037558f
C9660 VDD.t1587 VSS 0.006764f
C9661 VDD.t627 VSS 0.006764f
C9662 VDD.n646 VSS 0.014917f
C9663 VDD.t625 VSS 0.006764f
C9664 VDD.t565 VSS 0.006764f
C9665 VDD.n647 VSS 0.014917f
C9666 VDD.t567 VSS 0.018157f
C9667 VDD.t427 VSS 0.021269f
C9668 VDD.t431 VSS 0.01669f
C9669 VDD.n648 VSS 0.070928f
C9670 VDD.t428 VSS 0.006764f
C9671 VDD.t430 VSS 0.006764f
C9672 VDD.n649 VSS 0.013528f
C9673 VDD.n650 VSS 0.036172f
C9674 VDD.t477 VSS 0.021269f
C9675 VDD.t476 VSS 0.01669f
C9676 VDD.n651 VSS 0.084502f
C9677 VDD.t1081 VSS 0.214331f
C9678 VDD.t1123 VSS 0.136969f
C9679 VDD.t2082 VSS 0.136969f
C9680 VDD.t2094 VSS 0.136969f
C9681 VDD.t664 VSS 0.136969f
C9682 VDD.t662 VSS 0.141408f
C9683 VDD.t1036 VSS 0.548156f
C9684 VDD.t1068 VSS 0.01979f
C9685 VDD.t1037 VSS 0.01669f
C9686 VDD.n652 VSS 0.040346f
C9687 VDD.t474 VSS 0.021269f
C9688 VDD.t473 VSS 0.01669f
C9689 VDD.n653 VSS 0.068817f
C9690 VDD.t116 VSS 0.021269f
C9691 VDD.t114 VSS 0.01669f
C9692 VDD.n654 VSS 0.070928f
C9693 VDD.t115 VSS 0.006764f
C9694 VDD.t112 VSS 0.006764f
C9695 VDD.n655 VSS 0.013528f
C9696 VDD.n656 VSS 0.036172f
C9697 VDD.n657 VSS 0.032472f
C9698 VDD.t1117 VSS 0.214331f
C9699 VDD.t1143 VSS 0.136969f
C9700 VDD.t892 VSS 0.136969f
C9701 VDD.t903 VSS 0.136969f
C9702 VDD.t296 VSS 0.136969f
C9703 VDD.t294 VSS 0.141408f
C9704 VDD.t1066 VSS 0.341283f
C9705 VDD.t1067 VSS 0.01979f
C9706 VDD.t1142 VSS 0.01669f
C9707 VDD.n658 VSS 0.049398f
C9708 VDD.t1105 VSS 0.006764f
C9709 VDD.t1113 VSS 0.006764f
C9710 VDD.n659 VSS 0.01683f
C9711 VDD.t1126 VSS 0.006764f
C9712 VDD.t1101 VSS 0.006764f
C9713 VDD.n660 VSS 0.013528f
C9714 VDD.n661 VSS 0.027737f
C9715 VDD.t514 VSS 0.018157f
C9716 VDD.t512 VSS 0.006764f
C9717 VDD.t1692 VSS 0.006764f
C9718 VDD.n662 VSS 0.014917f
C9719 VDD.t1685 VSS 0.006764f
C9720 VDD.t761 VSS 0.006764f
C9721 VDD.n663 VSS 0.014917f
C9722 VDD.t763 VSS 0.018157f
C9723 VDD.n664 VSS 0.056289f
C9724 VDD.n665 VSS 0.0563f
C9725 VDD.n666 VSS 0.033732f
C9726 VDD.t1118 VSS 0.018316f
C9727 VDD.t1144 VSS 0.006764f
C9728 VDD.t893 VSS 0.006764f
C9729 VDD.n667 VSS 0.014917f
C9730 VDD.t904 VSS 0.006764f
C9731 VDD.t297 VSS 0.006764f
C9732 VDD.n668 VSS 0.014917f
C9733 VDD.t295 VSS 0.022409f
C9734 VDD.n669 VSS 0.096335f
C9735 VDD.n670 VSS 0.033732f
C9736 VDD.n671 VSS 0.096908f
C9737 VDD.n672 VSS 0.07211f
C9738 VDD.n673 VSS 0.037558f
C9739 VDD.n674 VSS 0.015175f
C9740 VDD.n675 VSS 0.018755f
C9741 VDD.n676 VSS 0.102565f
C9742 VDD.t1104 VSS 0.138882f
C9743 VDD.t1100 VSS 0.363892f
C9744 VDD.t513 VSS 0.214331f
C9745 VDD.t511 VSS 0.136969f
C9746 VDD.t1691 VSS 0.136969f
C9747 VDD.t1684 VSS 0.136969f
C9748 VDD.t760 VSS 0.136969f
C9749 VDD.t762 VSS 0.141408f
C9750 VDD.n677 VSS 0.356736f
C9751 VDD.t113 VSS 0.408943f
C9752 VDD.t111 VSS 0.219141f
C9753 VDD.t189 VSS 0.882358f
C9754 VDD.t188 VSS 0.375016f
C9755 VDD.n678 VSS 0.189733f
C9756 VDD.n679 VSS -0.002571f
C9757 VDD.n680 VSS 0.072393f
C9758 VDD.n681 VSS 0.037945f
C9759 VDD.t1084 VSS 0.006764f
C9760 VDD.t1076 VSS 0.006764f
C9761 VDD.n682 VSS 0.01683f
C9762 VDD.t1137 VSS 0.006764f
C9763 VDD.t1125 VSS 0.006764f
C9764 VDD.n683 VSS 0.013528f
C9765 VDD.n684 VSS 0.027737f
C9766 VDD.n685 VSS 0.015175f
C9767 VDD.n686 VSS 0.006361f
C9768 VDD.n687 VSS 0.102565f
C9769 VDD.t1083 VSS 0.138882f
C9770 VDD.t1075 VSS 0.363892f
C9771 VDD.t1584 VSS 0.214331f
C9772 VDD.t1586 VSS 0.136969f
C9773 VDD.t626 VSS 0.136969f
C9774 VDD.t624 VSS 0.136969f
C9775 VDD.t564 VSS 0.136969f
C9776 VDD.t566 VSS 0.141408f
C9777 VDD.n688 VSS 0.356736f
C9778 VDD.t426 VSS 0.408943f
C9779 VDD.t429 VSS 0.219141f
C9780 VDD.t475 VSS 0.619833f
C9781 VDD.t666 VSS 0.375016f
C9782 VDD.n689 VSS 0.189733f
C9783 VDD.n690 VSS -0.002571f
C9784 VDD.n691 VSS 0.032472f
C9785 VDD.n692 VSS 0.056289f
C9786 VDD.n693 VSS 0.0563f
C9787 VDD.n694 VSS 0.033732f
C9788 VDD.n695 VSS 0.032867f
C9789 VDD.t1082 VSS 0.018316f
C9790 VDD.t1124 VSS 0.006764f
C9791 VDD.t2083 VSS 0.006764f
C9792 VDD.n696 VSS 0.014917f
C9793 VDD.t2095 VSS 0.006764f
C9794 VDD.t665 VSS 0.006764f
C9795 VDD.n697 VSS 0.014917f
C9796 VDD.t663 VSS 0.022409f
C9797 VDD.n698 VSS 0.096335f
C9798 VDD.n699 VSS 0.033732f
C9799 VDD.n700 VSS 0.044404f
C9800 VDD.n701 VSS 0.378059f
C9801 VDD.n702 VSS 0.235278f
C9802 VDD.t131 VSS 0.16641f
C9803 VDD.n703 VSS 0.251862f
C9804 VDD.t129 VSS 0.721486f
C9805 VDD.t531 VSS 0.726829f
C9806 VDD.t527 VSS 0.288488f
C9807 VDD.t529 VSS 0.317265f
C9808 VDD.t1204 VSS 0.334568f
C9809 VDD.t942 VSS 0.992796f
C9810 VDD.t708 VSS 0.224542f
C9811 VDD.t1990 VSS 0.431017f
C9812 VDD.t1991 VSS 0.231449f
C9813 VDD.t1703 VSS 0.018322f
C9814 VDD.t896 VSS 0.006764f
C9815 VDD.t1906 VSS 0.006764f
C9816 VDD.n704 VSS 0.015166f
C9817 VDD.n705 VSS 0.043025f
C9818 VDD.n706 VSS 0.08163f
C9819 VDD.t868 VSS 0.006764f
C9820 VDD.t906 VSS 0.006764f
C9821 VDD.n707 VSS 0.015166f
C9822 VDD.n708 VSS 0.035907f
C9823 VDD.t975 VSS 0.116433f
C9824 VDD.t976 VSS 0.006764f
C9825 VDD.t980 VSS 0.006764f
C9826 VDD.n709 VSS 0.015166f
C9827 VDD.t986 VSS 0.018322f
C9828 VDD.t506 VSS 0.018322f
C9829 VDD.t508 VSS 0.006764f
C9830 VDD.t504 VSS 0.006764f
C9831 VDD.n710 VSS 0.015166f
C9832 VDD.t510 VSS 0.022391f
C9833 VDD.n711 VSS 0.095048f
C9834 VDD.t851 VSS 0.116433f
C9835 VDD.t852 VSS 0.006764f
C9836 VDD.t900 VSS 0.006764f
C9837 VDD.n712 VSS 0.015166f
C9838 VDD.t812 VSS 0.018322f
C9839 VDD.t950 VSS 0.018322f
C9840 VDD.t954 VSS 0.006764f
C9841 VDD.t952 VSS 0.006764f
C9842 VDD.n713 VSS 0.015166f
C9843 VDD.t956 VSS 0.018322f
C9844 VDD.t1305 VSS 0.018422f
C9845 VDD.t1262 VSS 0.006764f
C9846 VDD.t1264 VSS 0.006764f
C9847 VDD.n714 VSS 0.015166f
C9848 VDD.n715 VSS 0.035894f
C9849 VDD.t1304 VSS 0.227678f
C9850 VDD.t1261 VSS 0.103398f
C9851 VDD.t86 VSS 0.314619f
C9852 VDD.t981 VSS 0.314619f
C9853 VDD.t973 VSS 0.356588f
C9854 VDD.t984 VSS 0.018322f
C9855 VDD.t1293 VSS 0.018313f
C9856 VDD.n716 VSS 0.051521f
C9857 VDD.n717 VSS 0.059268f
C9858 VDD.t972 VSS 0.006764f
C9859 VDD.t974 VSS 0.006764f
C9860 VDD.n718 VSS 0.015166f
C9861 VDD.t982 VSS 0.018322f
C9862 VDD.n719 VSS 0.090004f
C9863 VDD.n720 VSS 0.043025f
C9864 VDD.n721 VSS -0.011488f
C9865 VDD.n722 VSS 0.060717f
C9866 VDD.t971 VSS 0.104824f
C9867 VDD.t983 VSS 0.230818f
C9868 VDD.t1292 VSS 0.227678f
C9869 VDD.t1263 VSS 0.114849f
C9870 VDD.n723 VSS 0.061018f
C9871 VDD.n724 VSS -0.010928f
C9872 VDD.n725 VSS 0.134973f
C9873 VDD.n726 VSS 0.141428f
C9874 VDD.n727 VSS 0.041121f
C9875 VDD.t955 VSS 0.227678f
C9876 VDD.t953 VSS 0.114849f
C9877 VDD.t811 VSS 0.230818f
C9878 VDD.t710 VSS 0.230818f
C9879 VDD.t711 VSS 0.147505f
C9880 VDD.t712 VSS 0.230818f
C9881 VDD.t949 VSS 0.227678f
C9882 VDD.t951 VSS 0.103398f
C9883 VDD.n728 VSS 0.061018f
C9884 VDD.n729 VSS -0.010718f
C9885 VDD.n730 VSS 0.08647f
C9886 VDD.n731 VSS 0.090838f
C9887 VDD.n732 VSS 0.043025f
C9888 VDD.t1895 VSS 0.022055f
C9889 VDD.n733 VSS -0.011488f
C9890 VDD.n734 VSS 0.062021f
C9891 VDD.t899 VSS 0.104824f
C9892 VDD.t1894 VSS 0.283776f
C9893 VDD.t509 VSS 0.283492f
C9894 VDD.t507 VSS 0.116235f
C9895 VDD.t985 VSS 0.230818f
C9896 VDD.t731 VSS 0.230818f
C9897 VDD.t732 VSS 0.147505f
C9898 VDD.t733 VSS 0.214099f
C9899 VDD.t505 VSS 0.213738f
C9900 VDD.t503 VSS 0.104645f
C9901 VDD.n735 VSS 0.061895f
C9902 VDD.n736 VSS -0.010623f
C9903 VDD.n737 VSS 0.086535f
C9904 VDD.n738 VSS 0.089368f
C9905 VDD.n739 VSS 0.043025f
C9906 VDD.t978 VSS 0.018322f
C9907 VDD.t814 VSS 0.018322f
C9908 VDD.n740 VSS 0.050861f
C9909 VDD.n741 VSS 0.058884f
C9910 VDD.n742 VSS -0.011488f
C9911 VDD.n743 VSS 0.062021f
C9912 VDD.t979 VSS 0.104824f
C9913 VDD.t977 VSS 0.222676f
C9914 VDD.t813 VSS 0.219653f
C9915 VDD.t867 VSS 0.114849f
C9916 VDD.t861 VSS 0.227678f
C9917 VDD.t905 VSS 0.103398f
C9918 VDD.n744 VSS 0.061018f
C9919 VDD.n745 VSS -0.010928f
C9920 VDD.t862 VSS 0.018342f
C9921 VDD.n746 VSS -0.094981f
C9922 VDD.n747 VSS -0.163936f
C9923 VDD.t1301 VSS 0.018961f
C9924 VDD.n748 VSS 0.050186f
C9925 VDD.t210 VSS 0.027992f
C9926 VDD.n749 VSS 0.046198f
C9927 VDD.t212 VSS 0.034731f
C9928 VDD.t1639 VSS 0.006764f
C9929 VDD.t314 VSS 0.006764f
C9930 VDD.n750 VSS 0.029826f
C9931 VDD.t2148 VSS 0.006764f
C9932 VDD.t1650 VSS 0.006764f
C9933 VDD.n751 VSS 0.013528f
C9934 VDD.n752 VSS 0.039293f
C9935 VDD.t1638 VSS 0.006764f
C9936 VDD.t315 VSS 0.006764f
C9937 VDD.n753 VSS 0.029015f
C9938 VDD.n754 VSS 0.03765f
C9939 VDD.t2149 VSS 0.006764f
C9940 VDD.t1651 VSS 0.006764f
C9941 VDD.n755 VSS 0.013528f
C9942 VDD.n756 VSS 0.008042f
C9943 VDD.t1294 VSS 0.227678f
C9944 VDD.t1298 VSS 0.114849f
C9945 VDD.t1299 VSS 0.006764f
C9946 VDD.t1260 VSS 0.006764f
C9947 VDD.n757 VSS 0.015166f
C9948 VDD.t1295 VSS 0.022873f
C9949 VDD.n758 VSS 0.07781f
C9950 VDD.n759 VSS -0.010928f
C9951 VDD.n760 VSS 0.061018f
C9952 VDD.t1259 VSS 0.103398f
C9953 VDD.t1300 VSS 0.282698f
C9954 VDD.t211 VSS 0.443429f
C9955 VDD.t501 VSS 0.225027f
C9956 VDD.n761 VSS 0.178745f
C9957 VDD.t2147 VSS 0.162133f
C9958 VDD.t1649 VSS 0.185802f
C9959 VDD.t313 VSS 0.400006f
C9960 VDD.t1637 VSS 0.197636f
C9961 VDD.n762 VSS 0.100515f
C9962 VDD.n763 VSS 0.027244f
C9963 VDD.n764 VSS 0.041492f
C9964 VDD.n765 VSS 0.023102f
C9965 VDD.n766 VSS 0.274776f
C9966 VDD.n767 VSS 0.193896f
C9967 VDD.t1533 VSS 0.006764f
C9968 VDD.t1531 VSS 0.006764f
C9969 VDD.n768 VSS 0.018548f
C9970 VDD.t1540 VSS 0.006764f
C9971 VDD.t1539 VSS 0.006764f
C9972 VDD.n769 VSS 0.013528f
C9973 VDD.n770 VSS 0.044415f
C9974 VDD.n771 VSS 0.024748f
C9975 VDD.n772 VSS 0.129987f
C9976 VDD.t1532 VSS 0.126882f
C9977 VDD.n773 VSS 0.09309f
C9978 VDD.n774 VSS 0.009557f
C9979 VDD.t1242 VSS 0.021269f
C9980 VDD.t1228 VSS 0.01669f
C9981 VDD.n775 VSS 0.05249f
C9982 VDD.t1235 VSS 0.01669f
C9983 VDD.n776 VSS 0.032061f
C9984 VDD.t1253 VSS 0.01669f
C9985 VDD.n777 VSS 0.032061f
C9986 VDD.t1231 VSS 0.01669f
C9987 VDD.n778 VSS 0.030191f
C9988 VDD.t1234 VSS 0.01669f
C9989 VDD.n779 VSS 0.025944f
C9990 VDD.n780 VSS 0.021649f
C9991 VDD.t1670 VSS 0.725035f
C9992 VDD.t1227 VSS 0.725035f
C9993 VDD.t1841 VSS 0.531559f
C9994 VDD.t1438 VSS 0.091458f
C9995 VDD.t1439 VSS 0.006764f
C9996 VDD.t1453 VSS 0.006764f
C9997 VDD.n781 VSS 0.018548f
C9998 VDD.t1443 VSS 0.006764f
C9999 VDD.t1430 VSS 0.006764f
C10000 VDD.n782 VSS 0.013528f
C10001 VDD.n783 VSS 0.043881f
C10002 VDD.t2172 VSS 0.021269f
C10003 VDD.t2171 VSS 0.01669f
C10004 VDD.n784 VSS 0.077501f
C10005 VDD.n785 VSS 0.080632f
C10006 VDD.n786 VSS 0.020433f
C10007 VDD.n787 VSS 0.032519f
C10008 VDD.n788 VSS 0.019487f
C10009 VDD.n789 VSS 0.019625f
C10010 VDD.n790 VSS 0.019349f
C10011 VDD.n791 VSS 0.017137f
C10012 VDD.n792 VSS 0.001662f
C10013 VDD.n793 VSS 0.019902f
C10014 VDD.n794 VSS 0.019487f
C10015 VDD.n795 VSS 0.019625f
C10016 VDD.n796 VSS 0.019349f
C10017 VDD.n797 VSS 0.001938f
C10018 VDD.n798 VSS 0.042208f
C10019 VDD.n799 VSS 0.001384f
C10020 VDD.n800 VSS 0.017137f
C10021 VDD.n801 VSS 0.017552f
C10022 VDD.n802 VSS 0.027927f
C10023 VDD.n803 VSS 0.019902f
C10024 VDD.n804 VSS 0.028993f
C10025 VDD.n805 VSS 0.068756f
C10026 VDD.n806 VSS 0.020531f
C10027 VDD.n807 VSS 0.019349f
C10028 VDD.n808 VSS 0.020242f
C10029 VDD.n809 VSS 0.052094f
C10030 VDD.n810 VSS 0.016155f
C10031 VDD.n811 VSS 0.015483f
C10032 VDD.n812 VSS 0.017552f
C10033 VDD.n813 VSS 0.017137f
C10034 VDD.n814 VSS 0.001108f
C10035 VDD.n815 VSS 0.037417f
C10036 VDD.n816 VSS 0.019625f
C10037 VDD.n817 VSS 0.019487f
C10038 VDD.n818 VSS 3.0154f
C10039 VDD.n819 VSS 0.001662f
C10040 VDD.n820 VSS 0.019902f
C10041 VDD.n821 VSS 0.019487f
C10042 VDD.n822 VSS 0.019625f
C10043 VDD.n823 VSS 0.019349f
C10044 VDD.n824 VSS 0.001938f
C10045 VDD.n825 VSS 0.031624f
C10046 VDD.n826 VSS 0.001384f
C10047 VDD.n827 VSS 0.017137f
C10048 VDD.n828 VSS 0.017552f
C10049 VDD.n829 VSS 0.027927f
C10050 VDD.n830 VSS 0.019902f
C10051 VDD.n831 VSS 0.028993f
C10052 VDD.n832 VSS 0.068756f
C10053 VDD.n833 VSS 0.020531f
C10054 VDD.n834 VSS 0.019349f
C10055 VDD.n835 VSS 0.020242f
C10056 VDD.n836 VSS 0.052094f
C10057 VDD.n837 VSS 0.016155f
C10058 VDD.t29 VSS 0.018219f
C10059 VDD.n838 VSS 0.037783f
C10060 VDD.t1738 VSS 0.006764f
C10061 VDD.t1745 VSS 0.006764f
C10062 VDD.n839 VSS 0.01683f
C10063 VDD.t1729 VSS 0.006764f
C10064 VDD.t1741 VSS 0.006764f
C10065 VDD.n840 VSS 0.013528f
C10066 VDD.n841 VSS 0.027336f
C10067 VDD.n842 VSS 0.015759f
C10068 VDD.t1767 VSS 0.01979f
C10069 VDD.t1766 VSS 0.01669f
C10070 VDD.n843 VSS 0.049398f
C10071 VDD.n844 VSS 0.032342f
C10072 VDD.n845 VSS 0.034081f
C10073 VDD.t1034 VSS 0.566627f
C10074 VDD.t1029 VSS 0.01979f
C10075 VDD.t1062 VSS 0.01669f
C10076 VDD.n846 VSS 0.049398f
C10077 VDD.n847 VSS 0.018755f
C10078 VDD.t1085 VSS 0.302686f
C10079 VDD.n848 VSS 0.016505f
C10080 VDD.t1735 VSS 0.01979f
C10081 VDD.t1728 VSS 0.01669f
C10082 VDD.n849 VSS 0.049398f
C10083 VDD.t1765 VSS 0.006764f
C10084 VDD.t1744 VSS 0.006764f
C10085 VDD.n850 VSS 0.01683f
C10086 VDD.t1763 VSS 0.006764f
C10087 VDD.t1734 VSS 0.006764f
C10088 VDD.n851 VSS 0.013528f
C10089 VDD.n852 VSS 0.02771f
C10090 VDD.t2015 VSS 0.006764f
C10091 VDD.t49 VSS 0.006764f
C10092 VDD.n853 VSS 0.014917f
C10093 VDD.t53 VSS 0.006764f
C10094 VDD.t559 VSS 0.006764f
C10095 VDD.n854 VSS 0.014917f
C10096 VDD.t558 VSS 0.018157f
C10097 VDD.t85 VSS 0.021269f
C10098 VDD.t82 VSS 0.01669f
C10099 VDD.n855 VSS 0.070928f
C10100 VDD.t81 VSS 0.006764f
C10101 VDD.t83 VSS 0.006764f
C10102 VDD.n856 VSS 0.013528f
C10103 VDD.n857 VSS 0.036172f
C10104 VDD.t444 VSS 0.021269f
C10105 VDD.t445 VSS 0.01669f
C10106 VDD.n858 VSS 0.068817f
C10107 VDD.t199 VSS 0.017784f
C10108 VDD.t201 VSS 0.006764f
C10109 VDD.t450 VSS 0.006764f
C10110 VDD.n859 VSS 0.020425f
C10111 VDD.n860 VSS 0.059702f
C10112 VDD.t447 VSS 0.01669f
C10113 VDD.n861 VSS 0.017903f
C10114 VDD.t446 VSS 0.006764f
C10115 VDD.t449 VSS 0.006764f
C10116 VDD.n862 VSS 0.020425f
C10117 VDD.n863 VSS 0.039154f
C10118 VDD.n864 VSS 0.070125f
C10119 VDD.n865 VSS 0.07375f
C10120 VDD.t293 VSS 0.021269f
C10121 VDD.t291 VSS 0.01669f
C10122 VDD.n866 VSS 0.070928f
C10123 VDD.t292 VSS 0.006764f
C10124 VDD.t290 VSS 0.006764f
C10125 VDD.n867 VSS 0.013528f
C10126 VDD.n868 VSS 0.036172f
C10127 VDD.t72 VSS 0.018157f
C10128 VDD.t1592 VSS 0.006764f
C10129 VDD.t2000 VSS 0.006764f
C10130 VDD.n869 VSS 0.022549f
C10131 VDD.t1994 VSS 0.006764f
C10132 VDD.t74 VSS 0.006764f
C10133 VDD.n870 VSS 0.022549f
C10134 VDD.t1594 VSS 0.018157f
C10135 VDD.t1086 VSS 0.006764f
C10136 VDD.t1043 VSS 0.006764f
C10137 VDD.n871 VSS 0.01683f
C10138 VDD.t1114 VSS 0.006764f
C10139 VDD.t1074 VSS 0.006764f
C10140 VDD.n872 VSS 0.013528f
C10141 VDD.n873 VSS 0.027737f
C10142 VDD.n874 VSS 0.015175f
C10143 VDD.n875 VSS 0.037558f
C10144 VDD.t1134 VSS 0.018316f
C10145 VDD.t1049 VSS 0.006764f
C10146 VDD.t1916 VSS 0.006764f
C10147 VDD.n876 VSS 0.022549f
C10148 VDD.t891 VSS 0.006764f
C10149 VDD.t193 VSS 0.006764f
C10150 VDD.n877 VSS 0.022549f
C10151 VDD.t191 VSS 0.025643f
C10152 VDD.n878 VSS 0.104443f
C10153 VDD.n879 VSS 0.097077f
C10154 VDD.n880 VSS 0.072279f
C10155 VDD.n881 VSS 0.057655f
C10156 VDD.n882 VSS 0.066276f
C10157 VDD.n883 VSS 0.032472f
C10158 VDD.n884 VSS -0.002571f
C10159 VDD.t1133 VSS 0.214331f
C10160 VDD.t1048 VSS 0.136969f
C10161 VDD.t1915 VSS 0.136969f
C10162 VDD.t890 VSS 0.136969f
C10163 VDD.t192 VSS 0.136969f
C10164 VDD.t190 VSS 0.214331f
C10165 VDD.n885 VSS 0.26152f
C10166 VDD.t1042 VSS 0.566627f
C10167 VDD.t1593 VSS 0.51934f
C10168 VDD.t1591 VSS 0.331886f
C10169 VDD.t48 VSS 0.331886f
C10170 VDD.t52 VSS 0.331886f
C10171 VDD.t73 VSS 0.331886f
C10172 VDD.t71 VSS 0.51934f
C10173 VDD.t80 VSS 1.13446f
C10174 VDD.t76 VSS 0.433271f
C10175 VDD.t448 VSS 0.293512f
C10176 VDD.t1060 VSS 0.289491f
C10177 VDD.t200 VSS 0.289491f
C10178 VDD.t1044 VSS 0.060311f
C10179 VDD.t1031 VSS 0.01979f
C10180 VDD.t1063 VSS 0.01669f
C10181 VDD.n886 VSS 0.040346f
C10182 VDD.t78 VSS 0.021269f
C10183 VDD.t79 VSS 0.01669f
C10184 VDD.n887 VSS 0.068817f
C10185 VDD.n888 VSS 0.072393f
C10186 VDD.n889 VSS 0.037945f
C10187 VDD.t1045 VSS 0.006764f
C10188 VDD.t1061 VSS 0.006764f
C10189 VDD.n890 VSS 0.01683f
C10190 VDD.t1079 VSS 0.006764f
C10191 VDD.t1099 VSS 0.006764f
C10192 VDD.n891 VSS 0.013528f
C10193 VDD.n892 VSS 0.027737f
C10194 VDD.n893 VSS 0.033352f
C10195 VDD.n894 VSS 0.015175f
C10196 VDD.n895 VSS 0.006361f
C10197 VDD.n896 VSS 0.271763f
C10198 VDD.t198 VSS 0.233201f
C10199 VDD.t1030 VSS 1.19143f
C10200 VDD.t77 VSS 1.73753f
C10201 VDD.t1712 VSS 0.214331f
C10202 VDD.t1730 VSS 0.136969f
C10203 VDD.t1397 VSS 0.136969f
C10204 VDD.t1391 VSS 0.136969f
C10205 VDD.t453 VSS 0.136969f
C10206 VDD.t451 VSS 0.214331f
C10207 VDD.t84 VSS 0.151131f
C10208 VDD.t462 VSS 0.072435f
C10209 VDD.t443 VSS 0.175276f
C10210 VDD.n897 VSS 0.169938f
C10211 VDD.t75 VSS 0.419767f
C10212 VDD.n898 VSS 0.213776f
C10213 VDD.n899 VSS 0.275324f
C10214 VDD.n901 VSS 0.123719f
C10215 VDD.n902 VSS -0.002571f
C10216 VDD.n903 VSS 0.032472f
C10217 VDD.n904 VSS 0.056289f
C10218 VDD.n905 VSS 0.0563f
C10219 VDD.n906 VSS 0.033732f
C10220 VDD.t1713 VSS 0.018316f
C10221 VDD.t1731 VSS 0.006764f
C10222 VDD.t1398 VSS 0.006764f
C10223 VDD.n907 VSS 0.014917f
C10224 VDD.t1392 VSS 0.006764f
C10225 VDD.t454 VSS 0.006764f
C10226 VDD.n908 VSS 0.014917f
C10227 VDD.t452 VSS 0.022409f
C10228 VDD.n909 VSS 0.096335f
C10229 VDD.n910 VSS 0.033732f
C10230 VDD.n911 VSS 0.096908f
C10231 VDD.n912 VSS 0.072636f
C10232 VDD.t2014 VSS 0.018218f
C10233 VDD.n913 VSS 0.038386f
C10234 VDD.n914 VSS 0.015251f
C10235 VDD.n915 VSS 0.032455f
C10236 VDD.n916 VSS 0.034081f
C10237 VDD.n917 VSS 0.247812f
C10238 VDD.t1028 VSS 0.930341f
C10239 VDD.t1095 VSS 0.930341f
C10240 VDD.t1035 VSS 0.006764f
C10241 VDD.t1047 VSS 0.006764f
C10242 VDD.n918 VSS 0.01683f
C10243 VDD.t1065 VSS 0.006764f
C10244 VDD.t1080 VSS 0.006764f
C10245 VDD.n919 VSS 0.013528f
C10246 VDD.n920 VSS 0.027737f
C10247 VDD.t1583 VSS 0.018157f
C10248 VDD.t1859 VSS 0.006764f
C10249 VDD.t1582 VSS 0.006764f
C10250 VDD.n921 VSS 0.014917f
C10251 VDD.t36 VSS 0.006764f
C10252 VDD.t1850 VSS 0.006764f
C10253 VDD.n922 VSS 0.014917f
C10254 VDD.t34 VSS 0.018157f
C10255 VDD.t39 VSS 0.021269f
C10256 VDD.t42 VSS 0.01669f
C10257 VDD.n923 VSS 0.070928f
C10258 VDD.t41 VSS 0.006764f
C10259 VDD.t38 VSS 0.006764f
C10260 VDD.n924 VSS 0.013528f
C10261 VDD.n925 VSS 0.036172f
C10262 VDD.t1129 VSS 0.214331f
C10263 VDD.t1131 VSS 0.136969f
C10264 VDD.t859 VSS 0.136969f
C10265 VDD.t827 VSS 0.136969f
C10266 VDD.t363 VSS 0.136969f
C10267 VDD.t361 VSS 0.214331f
C10268 VDD.t28 VSS 0.51934f
C10269 VDD.t26 VSS 0.331886f
C10270 VDD.t1700 VSS 0.331886f
C10271 VDD.t1698 VSS 0.331886f
C10272 VDD.t35 VSS 0.331886f
C10273 VDD.t33 VSS 0.51934f
C10274 VDD.t37 VSS 1.13446f
C10275 VDD.t40 VSS 0.433271f
C10276 VDD.t235 VSS 0.021269f
C10277 VDD.t233 VSS 0.01669f
C10278 VDD.n927 VSS 0.068817f
C10279 VDD.t2165 VSS 0.017784f
C10280 VDD.t158 VSS 0.006764f
C10281 VDD.t2166 VSS 0.006764f
C10282 VDD.n928 VSS 0.020425f
C10283 VDD.n929 VSS 0.059702f
C10284 VDD.t153 VSS 0.01669f
C10285 VDD.n930 VSS 0.017903f
C10286 VDD.t157 VSS 0.006764f
C10287 VDD.t155 VSS 0.006764f
C10288 VDD.n931 VSS 0.020425f
C10289 VDD.n932 VSS 0.039154f
C10290 VDD.t1872 VSS 0.047077f
C10291 VDD.t1702 VSS 0.006764f
C10292 VDD.t1870 VSS 0.006764f
C10293 VDD.n933 VSS 0.013528f
C10294 VDD.n934 VSS 0.057677f
C10295 VDD.t1697 VSS 0.01669f
C10296 VDD.n935 VSS 0.026665f
C10297 VDD.t1798 VSS 0.006764f
C10298 VDD.t1733 VSS 0.006764f
C10299 VDD.n936 VSS 0.014917f
C10300 VDD.t346 VSS 0.006764f
C10301 VDD.t1788 VSS 0.006764f
C10302 VDD.n937 VSS 0.014917f
C10303 VDD.t344 VSS 0.022409f
C10304 VDD.n938 VSS 0.096335f
C10305 VDD.n939 VSS 0.033732f
C10306 VDD.t1717 VSS 0.018316f
C10307 VDD.n940 VSS 0.044405f
C10308 VDD.t178 VSS 0.006764f
C10309 VDD.t1557 VSS 0.006764f
C10310 VDD.n941 VSS 0.014917f
C10311 VDD.t2176 VSS 0.006764f
C10312 VDD.t180 VSS 0.006764f
C10313 VDD.n942 VSS 0.014917f
C10314 VDD.t2174 VSS 0.018157f
C10315 VDD.n943 VSS 0.056289f
C10316 VDD.n944 VSS 0.0563f
C10317 VDD.n945 VSS 0.033732f
C10318 VDD.t1555 VSS 0.018157f
C10319 VDD.n946 VSS 0.037558f
C10320 VDD.n947 VSS 0.032874f
C10321 VDD.n948 VSS 0.378039f
C10322 VDD.n949 VSS 0.235291f
C10323 VDD.t2164 VSS 0.031331f
C10324 VDD.t230 VSS 0.421066f
C10325 VDD.t234 VSS 0.195308f
C10326 VDD.t1706 VSS 0.214331f
C10327 VDD.t1708 VSS 0.136969f
C10328 VDD.t1780 VSS 0.136969f
C10329 VDD.t1804 VSS 0.136969f
C10330 VDD.t352 VSS 0.136969f
C10331 VDD.t350 VSS 0.214331f
C10332 VDD.t95 VSS 0.168403f
C10333 VDD.t232 VSS 0.080714f
C10334 VDD.n950 VSS 0.152698f
C10335 VDD.n951 VSS 0.45946f
C10336 VDD.t231 VSS 1.73753f
C10337 VDD.t1093 VSS 1.19143f
C10338 VDD.t152 VSS 0.233201f
C10339 VDD.t1033 VSS 0.006764f
C10340 VDD.t1092 VSS 0.006764f
C10341 VDD.n953 VSS 0.01683f
C10342 VDD.t1064 VSS 0.006764f
C10343 VDD.t1116 VSS 0.006764f
C10344 VDD.n954 VSS 0.013528f
C10345 VDD.n955 VSS 0.027737f
C10346 VDD.t1646 VSS 0.018157f
C10347 VDD.t275 VSS 0.006764f
C10348 VDD.t1648 VSS 0.006764f
C10349 VDD.n956 VSS 0.014917f
C10350 VDD.t277 VSS 0.006764f
C10351 VDD.t273 VSS 0.006764f
C10352 VDD.n957 VSS 0.014917f
C10353 VDD.t279 VSS 0.018157f
C10354 VDD.t359 VSS 0.021269f
C10355 VDD.t360 VSS 0.01669f
C10356 VDD.n958 VSS 0.070928f
C10357 VDD.t357 VSS 0.006764f
C10358 VDD.t355 VSS 0.006764f
C10359 VDD.n959 VSS 0.013528f
C10360 VDD.n960 VSS 0.036172f
C10361 VDD.t2170 VSS 0.470286f
C10362 VDD.t1127 VSS 0.214331f
C10363 VDD.t1140 VSS 0.136969f
C10364 VDD.t2054 VSS 0.136969f
C10365 VDD.t2048 VSS 0.136969f
C10366 VDD.t374 VSS 0.136969f
C10367 VDD.t376 VSS 0.214331f
C10368 VDD.t358 VSS 0.405502f
C10369 VDD.t2167 VSS 0.194353f
C10370 VDD.n961 VSS 0.368016f
C10371 VDD.t1645 VSS 0.241701f
C10372 VDD.t2162 VSS 0.241701f
C10373 VDD.t1647 VSS 0.031331f
C10374 VDD.t1871 VSS 0.241701f
C10375 VDD.t274 VSS 0.241701f
C10376 VDD.t1869 VSS 0.241701f
C10377 VDD.t272 VSS 0.241701f
C10378 VDD.t1696 VSS 0.241701f
C10379 VDD.t276 VSS 0.480047f
C10380 VDD.t278 VSS 0.749059f
C10381 VDD.t354 VSS 0.63321f
C10382 VDD.t1429 VSS 0.235179f
C10383 VDD.t356 VSS 0.126299f
C10384 VDD.n962 VSS 0.10927f
C10385 VDD.n963 VSS -0.002571f
C10386 VDD.n964 VSS 0.032472f
C10387 VDD.n965 VSS 0.056289f
C10388 VDD.n966 VSS 0.0563f
C10389 VDD.n967 VSS 0.033732f
C10390 VDD.t595 VSS 0.047077f
C10391 VDD.t937 VSS 0.006764f
C10392 VDD.t597 VSS 0.006764f
C10393 VDD.n968 VSS 0.013528f
C10394 VDD.n969 VSS 0.057677f
C10395 VDD.t933 VSS 0.01669f
C10396 VDD.n970 VSS 0.026665f
C10397 VDD.t569 VSS 0.017784f
C10398 VDD.t545 VSS 0.006764f
C10399 VDD.t572 VSS 0.006764f
C10400 VDD.n971 VSS 0.020425f
C10401 VDD.n972 VSS 0.059702f
C10402 VDD.t543 VSS 0.01669f
C10403 VDD.n973 VSS 0.017903f
C10404 VDD.t539 VSS 0.006764f
C10405 VDD.t541 VSS 0.006764f
C10406 VDD.n974 VSS 0.020425f
C10407 VDD.n975 VSS 0.039154f
C10408 VDD.n976 VSS 0.095546f
C10409 VDD.t932 VSS 0.469879f
C10410 VDD.t570 VSS 0.214331f
C10411 VDD.t573 VSS 0.069436f
C10412 VDD.t936 VSS 0.383891f
C10413 VDD.t596 VSS 0.133959f
C10414 VDD.t594 VSS 0.103955f
C10415 VDD.t574 VSS 0.129766f
C10416 VDD.t544 VSS 0.133959f
C10417 VDD.t571 VSS 0.091476f
C10418 VDD.t536 VSS 0.195308f
C10419 VDD.t1097 VSS 0.214331f
C10420 VDD.t1102 VSS 0.136969f
C10421 VDD.t2044 VSS 0.136969f
C10422 VDD.t2036 VSS 0.136969f
C10423 VDD.t634 VSS 0.136969f
C10424 VDD.t636 VSS 0.214331f
C10425 VDD.t695 VSS 0.168403f
C10426 VDD.t100 VSS 0.080714f
C10427 VDD.n977 VSS 0.152698f
C10428 VDD.t693 VSS 0.20962f
C10429 VDD.t102 VSS 0.100469f
C10430 VDD.n978 VSS 0.179038f
C10431 VDD.t534 VSS 0.379239f
C10432 VDD.t568 VSS 0.321253f
C10433 VDD.t691 VSS 0.075777f
C10434 VDD.t537 VSS 0.021269f
C10435 VDD.t535 VSS 0.01669f
C10436 VDD.n979 VSS 0.068817f
C10437 VDD.n980 VSS 0.07375f
C10438 VDD.t696 VSS 0.021269f
C10439 VDD.t694 VSS 0.01669f
C10440 VDD.n981 VSS 0.070928f
C10441 VDD.t692 VSS 0.006764f
C10442 VDD.t698 VSS 0.006764f
C10443 VDD.n982 VSS 0.013528f
C10444 VDD.n983 VSS 0.036172f
C10445 VDD.t522 VSS 0.018157f
C10446 VDD.t520 VSS 0.006764f
C10447 VDD.t939 VSS 0.006764f
C10448 VDD.n984 VSS 0.014917f
C10449 VDD.t935 VSS 0.006764f
C10450 VDD.t516 VSS 0.006764f
C10451 VDD.n985 VSS 0.014917f
C10452 VDD.t1059 VSS 0.006764f
C10453 VDD.t1078 VSS 0.006764f
C10454 VDD.n986 VSS 0.01683f
C10455 VDD.t1108 VSS 0.006764f
C10456 VDD.t1088 VSS 0.006764f
C10457 VDD.n987 VSS 0.013528f
C10458 VDD.n988 VSS 0.02771f
C10459 VDD.n989 VSS 0.015251f
C10460 VDD.t1120 VSS 0.01979f
C10461 VDD.t1051 VSS 0.01669f
C10462 VDD.n990 VSS 0.047504f
C10463 VDD.n991 VSS 0.034042f
C10464 VDD.n992 VSS 0.009282f
C10465 VDD.n993 VSS 0.034081f
C10466 VDD.t697 VSS 0.214331f
C10467 VDD.t521 VSS 0.214331f
C10468 VDD.t519 VSS 0.136969f
C10469 VDD.t938 VSS 0.136969f
C10470 VDD.t934 VSS 0.136969f
C10471 VDD.t515 VSS 0.136969f
C10472 VDD.t517 VSS 0.214331f
C10473 VDD.t1107 VSS 0.148383f
C10474 VDD.t1058 VSS 0.149561f
C10475 VDD.t1077 VSS 0.095577f
C10476 VDD.t1119 VSS 0.125444f
C10477 VDD.t1072 VSS 0.149561f
C10478 VDD.t1111 VSS 0.095577f
C10479 VDD.t1056 VSS 0.125444f
C10480 VDD.t1145 VSS 0.079264f
C10481 VDD.n994 VSS 0.016505f
C10482 VDD.t1057 VSS 0.01979f
C10483 VDD.t1055 VSS 0.01669f
C10484 VDD.n995 VSS 0.049398f
C10485 VDD.t1112 VSS 0.006764f
C10486 VDD.t1073 VSS 0.006764f
C10487 VDD.n996 VSS 0.01683f
C10488 VDD.t1146 VSS 0.006764f
C10489 VDD.t1027 VSS 0.006764f
C10490 VDD.n997 VSS 0.013528f
C10491 VDD.n998 VSS 0.02771f
C10492 VDD.t1025 VSS 0.006764f
C10493 VDD.t988 VSS 0.006764f
C10494 VDD.n999 VSS 0.014917f
C10495 VDD.t990 VSS 0.006764f
C10496 VDD.t269 VSS 0.006764f
C10497 VDD.n1000 VSS 0.014917f
C10498 VDD.t271 VSS 0.018157f
C10499 VDD.t643 VSS 0.021269f
C10500 VDD.t649 VSS 0.01669f
C10501 VDD.n1001 VSS 0.070928f
C10502 VDD.t645 VSS 0.006764f
C10503 VDD.t647 VSS 0.006764f
C10504 VDD.n1002 VSS 0.013528f
C10505 VDD.n1003 VSS 0.036172f
C10506 VDD.t1616 VSS 0.021269f
C10507 VDD.t1614 VSS 0.01669f
C10508 VDD.n1004 VSS 0.068817f
C10509 VDD.n1005 VSS 0.07375f
C10510 VDD.n1006 VSS 0.068485f
C10511 VDD.t1026 VSS 0.148383f
C10512 VDD.t1022 VSS 0.214331f
C10513 VDD.t1024 VSS 0.136969f
C10514 VDD.t987 VSS 0.136969f
C10515 VDD.t989 VSS 0.136969f
C10516 VDD.t268 VSS 0.136969f
C10517 VDD.t270 VSS 0.214331f
C10518 VDD.t644 VSS 0.214331f
C10519 VDD.t646 VSS 0.075777f
C10520 VDD.t1109 VSS 0.214331f
C10521 VDD.t1138 VSS 0.136969f
C10522 VDD.t1835 VSS 0.136969f
C10523 VDD.t1829 VSS 0.136969f
C10524 VDD.t782 VSS 0.136969f
C10525 VDD.t784 VSS 0.214331f
C10526 VDD.t642 VSS 0.168403f
C10527 VDD.t334 VSS 0.080714f
C10528 VDD.t1615 VSS 0.195308f
C10529 VDD.t648 VSS 0.237099f
C10530 VDD.t333 VSS 0.113639f
C10531 VDD.n1007 VSS 0.145849f
C10532 VDD.t1613 VSS 0.371586f
C10533 VDD.t1624 VSS 0.288488f
C10534 VDD.t1627 VSS 0.288488f
C10535 VDD.t1622 VSS 0.298505f
C10536 VDD.n1008 VSS 0.514195f
C10537 VDD.t332 VSS 0.306898f
C10538 VDD.t331 VSS 0.10241f
C10539 VDD.n1009 VSS 0.174831f
C10540 VDD.n1010 VSS 0.026241f
C10541 VDD.n1011 VSS -0.002571f
C10542 VDD.n1012 VSS 0.032472f
C10543 VDD.n1013 VSS 0.056289f
C10544 VDD.n1014 VSS 0.0563f
C10545 VDD.n1015 VSS 0.033732f
C10546 VDD.t1110 VSS 0.018316f
C10547 VDD.t1139 VSS 0.006764f
C10548 VDD.t1836 VSS 0.006764f
C10549 VDD.n1016 VSS 0.014917f
C10550 VDD.t1830 VSS 0.006764f
C10551 VDD.t783 VSS 0.006764f
C10552 VDD.n1017 VSS 0.014917f
C10553 VDD.t785 VSS 0.022409f
C10554 VDD.n1018 VSS 0.096335f
C10555 VDD.n1019 VSS 0.033732f
C10556 VDD.n1020 VSS 0.096908f
C10557 VDD.n1021 VSS 0.072636f
C10558 VDD.t1023 VSS 0.018218f
C10559 VDD.n1022 VSS 0.038386f
C10560 VDD.n1023 VSS 0.015251f
C10561 VDD.n1024 VSS 0.032455f
C10562 VDD.n1025 VSS 0.034081f
C10563 VDD.n1026 VSS 0.068485f
C10564 VDD.t1054 VSS 0.166455f
C10565 VDD.n1027 VSS 0.377886f
C10566 VDD.t1050 VSS 0.166455f
C10567 VDD.n1028 VSS 0.068485f
C10568 VDD.t1087 VSS 0.079264f
C10569 VDD.n1029 VSS 0.068485f
C10570 VDD.n1030 VSS 0.016505f
C10571 VDD.t518 VSS 0.018219f
C10572 VDD.n1031 VSS 0.03844f
C10573 VDD.t2045 VSS 0.006764f
C10574 VDD.t1103 VSS 0.006764f
C10575 VDD.n1032 VSS 0.014917f
C10576 VDD.t635 VSS 0.006764f
C10577 VDD.t2037 VSS 0.006764f
C10578 VDD.n1033 VSS 0.014917f
C10579 VDD.t637 VSS 0.022409f
C10580 VDD.n1034 VSS 0.096335f
C10581 VDD.n1035 VSS 0.033732f
C10582 VDD.t1098 VSS 0.018316f
C10583 VDD.n1036 VSS 0.096908f
C10584 VDD.n1037 VSS 0.072625f
C10585 VDD.n1038 VSS 0.033732f
C10586 VDD.n1039 VSS 0.0563f
C10587 VDD.n1040 VSS 0.056289f
C10588 VDD.n1041 VSS 0.032472f
C10589 VDD.n1042 VSS -0.002571f
C10590 VDD.n1043 VSS 0.060166f
C10591 VDD.t99 VSS 0.129677f
C10592 VDD.t101 VSS 0.353519f
C10593 VDD.t542 VSS 0.328472f
C10594 VDD.n1044 VSS 0.135464f
C10595 VDD.t540 VSS 0.093532f
C10596 VDD.t538 VSS 0.136969f
C10597 VDD.t575 VSS 0.136018f
C10598 VDD.n1045 VSS -0.083222f
C10599 VDD.n1046 VSS -0.085172f
C10600 VDD.n1047 VSS 0.235291f
C10601 VDD.t2055 VSS 0.006764f
C10602 VDD.t1141 VSS 0.006764f
C10603 VDD.n1048 VSS 0.014917f
C10604 VDD.t375 VSS 0.006764f
C10605 VDD.t2049 VSS 0.006764f
C10606 VDD.n1049 VSS 0.014917f
C10607 VDD.t377 VSS 0.022409f
C10608 VDD.n1050 VSS 0.096335f
C10609 VDD.n1051 VSS 0.033732f
C10610 VDD.t1128 VSS 0.018316f
C10611 VDD.n1052 VSS 0.044405f
C10612 VDD.n1053 VSS 0.378039f
C10613 VDD.n1054 VSS 0.032874f
C10614 VDD.n1055 VSS 0.037558f
C10615 VDD.n1056 VSS 0.015175f
C10616 VDD.t1094 VSS 0.01979f
C10617 VDD.t1121 VSS 0.01669f
C10618 VDD.n1057 VSS 0.040346f
C10619 VDD.t623 VSS 0.021269f
C10620 VDD.t622 VSS 0.01669f
C10621 VDD.n1058 VSS 0.068817f
C10622 VDD.n1059 VSS 0.072393f
C10623 VDD.n1060 VSS 0.037945f
C10624 VDD.n1061 VSS 0.006361f
C10625 VDD.n1062 VSS 0.271763f
C10626 VDD.t1091 VSS 0.060311f
C10627 VDD.t154 VSS 0.289491f
C10628 VDD.t1032 VSS 0.289491f
C10629 VDD.t156 VSS 0.293512f
C10630 VDD.t2163 VSS 0.538892f
C10631 VDD.n1063 VSS 0.083806f
C10632 VDD.n1064 VSS -0.085172f
C10633 VDD.n1065 VSS 0.095546f
C10634 VDD.n1066 VSS 0.07375f
C10635 VDD.t96 VSS 0.021269f
C10636 VDD.t98 VSS 0.01669f
C10637 VDD.n1067 VSS 0.070928f
C10638 VDD.t94 VSS 0.006764f
C10639 VDD.t97 VSS 0.006764f
C10640 VDD.n1068 VSS 0.013528f
C10641 VDD.n1069 VSS 0.036172f
C10642 VDD.t92 VSS 0.018157f
C10643 VDD.t93 VSS 0.006764f
C10644 VDD.t1699 VSS 0.006764f
C10645 VDD.n1070 VSS 0.014917f
C10646 VDD.t1701 VSS 0.006764f
C10647 VDD.t27 VSS 0.006764f
C10648 VDD.n1071 VSS 0.014917f
C10649 VDD.t1781 VSS 0.006764f
C10650 VDD.t1709 VSS 0.006764f
C10651 VDD.n1072 VSS 0.014917f
C10652 VDD.t353 VSS 0.006764f
C10653 VDD.t1805 VSS 0.006764f
C10654 VDD.n1073 VSS 0.014917f
C10655 VDD.t351 VSS 0.022409f
C10656 VDD.n1074 VSS 0.096335f
C10657 VDD.n1075 VSS 0.033732f
C10658 VDD.t1707 VSS 0.018316f
C10659 VDD.n1076 VSS 0.096908f
C10660 VDD.n1077 VSS 0.072625f
C10661 VDD.n1078 VSS 0.033732f
C10662 VDD.n1079 VSS 0.0563f
C10663 VDD.n1080 VSS 0.056289f
C10664 VDD.n1081 VSS 0.032472f
C10665 VDD.n1082 VSS -0.002571f
C10666 VDD.n1083 VSS 0.123719f
C10667 VDD.n1084 VSS -0.002571f
C10668 VDD.n1085 VSS 0.032472f
C10669 VDD.n1086 VSS 0.056289f
C10670 VDD.n1087 VSS 0.0563f
C10671 VDD.n1088 VSS 0.033732f
C10672 VDD.t364 VSS 0.006764f
C10673 VDD.t828 VSS 0.006764f
C10674 VDD.n1089 VSS 0.022549f
C10675 VDD.t860 VSS 0.006764f
C10676 VDD.t1132 VSS 0.006764f
C10677 VDD.n1090 VSS 0.022549f
C10678 VDD.t362 VSS 0.025643f
C10679 VDD.n1091 VSS 0.104443f
C10680 VDD.t1130 VSS 0.018316f
C10681 VDD.n1092 VSS 0.097077f
C10682 VDD.n1093 VSS 0.07211f
C10683 VDD.n1094 VSS 0.037558f
C10684 VDD.n1095 VSS 0.015175f
C10685 VDD.t1096 VSS 0.01979f
C10686 VDD.t1122 VSS 0.01669f
C10687 VDD.n1096 VSS 0.049398f
C10688 VDD.n1097 VSS 0.018755f
C10689 VDD.n1098 VSS 0.247812f
C10690 VDD.t1046 VSS 0.302686f
C10691 VDD.n1099 VSS 0.26152f
C10692 VDD.n1100 VSS 0.016505f
C10693 VDD.n1101 VSS 0.030339f
C10694 VDD.n1102 VSS 3.14558f
C10695 VDD.n1103 VSS 1.68964f
C10696 VDD.n1104 VSS 0.015483f
C10697 VDD.n1105 VSS 0.017552f
C10698 VDD.n1106 VSS 0.017137f
C10699 VDD.n1107 VSS 0.001108f
C10700 VDD.n1108 VSS 0.030684f
C10701 VDD.n1109 VSS 0.019625f
C10702 VDD.n1110 VSS 0.019487f
C10703 VDD.n1111 VSS 0.074233f
C10704 VDD.n1112 VSS 5.517951f
C10705 VDD.n1113 VSS 1.7978f
C10706 VDD.n1114 VSS 0.056192f
C10707 VDD.n1115 VSS 0.038642f
C10708 VDD.n1116 VSS 0.017552f
C10709 VDD.n1117 VSS 0.032095f
C10710 VDD.n1118 VSS 0.028482f
C10711 VDD.n1119 VSS 0.028993f
C10712 VDD.n1120 VSS 0.019902f
C10713 VDD.n1121 VSS 0.019487f
C10714 VDD.n1122 VSS 0.068756f
C10715 VDD.n1123 VSS 0.020531f
C10716 VDD.n1124 VSS 0.020242f
C10717 VDD.n1125 VSS 0.017137f
C10718 VDD.n1126 VSS 0.052094f
C10719 VDD.n1127 VSS 0.016155f
C10720 VDD.n1128 VSS 0.015483f
C10721 VDD.n1129 VSS 0.017552f
C10722 VDD.n1130 VSS 0.015586f
C10723 VDD.n1131 VSS 0.015999f
C10724 VDD.n1132 VSS 0.019349f
C10725 VDD.n1133 VSS 0.019625f
C10726 VDD.n1134 VSS 0.004906f
C10727 VDD.n1135 VSS 1.74767f
C10728 VDD.n1136 VSS 0.001662f
C10729 VDD.n1137 VSS 0.019906f
C10730 VDD.n1138 VSS 0.019487f
C10731 VDD.n1139 VSS 0.019625f
C10732 VDD.n1140 VSS 0.019349f
C10733 VDD.n1141 VSS 0.018256f
C10734 VDD.n1142 VSS 0.032026f
C10735 VDD.n1143 VSS 0.017137f
C10736 VDD.n1144 VSS 0.017552f
C10737 VDD.n1145 VSS 0.027927f
C10738 VDD.n1146 VSS 0.019902f
C10739 VDD.n1147 VSS 0.028993f
C10740 VDD.n1148 VSS 0.068756f
C10741 VDD.n1149 VSS 0.020531f
C10742 VDD.n1150 VSS 0.019349f
C10743 VDD.n1151 VSS 0.020242f
C10744 VDD.n1152 VSS 0.052094f
C10745 VDD.n1153 VSS 0.016155f
C10746 VDD.n1154 VSS 0.015609f
C10747 VDD.n1155 VSS 0.017701f
C10748 VDD.n1156 VSS 0.017137f
C10749 VDD.n1157 VSS 0.048746f
C10750 VDD.n1158 VSS 0.013572f
C10751 VDD.n1159 VSS 0.019625f
C10752 VDD.n1160 VSS 0.019487f
C10753 VDD.n1161 VSS 4.31689f
C10754 VDD.n1162 VSS 5.96049f
C10755 VDD.n1163 VSS 0.053047f
C10756 VDD.n1164 VSS 0.093523f
C10757 VDD.t2169 VSS 0.160053f
C10758 VDD.t2131 VSS 0.235179f
C10759 VDD.t2168 VSS 0.235179f
C10760 VDD.t2130 VSS 0.658108f
C10761 VDD.t1230 VSS 0.483498f
C10762 VDD.n1165 VSS 0.137721f
C10763 VDD.n1166 VSS 0.010735f
C10764 VDD.n1167 VSS 0.006958f
C10765 VDD.n1168 VSS 0.00788f
C10766 VDD.n1169 VSS 0.113471f
C10767 VDD.t1673 VSS 0.408064f
C10768 VDD.t1530 VSS 0.418265f
C10769 VDD.n1170 VSS 0.310939f
C10770 VDD.t706 VSS 0.144348f
C10771 VDD.t1202 VSS 0.195672f
C10772 VDD.t1201 VSS 0.175623f
C10773 VDD.n1171 VSS 0.02151f
C10774 VDD.n1172 VSS -0.085172f
C10775 VDD.n1173 VSS 0.095546f
C10776 VDD.n1174 VSS 0.07375f
C10777 VDD.n1175 VSS -0.002571f
C10778 VDD.n1176 VSS 0.135925f
C10779 VDD.t127 VSS 0.159604f
C10780 VDD.t671 VSS 0.518591f
C10781 VDD.t502 VSS 1.42388f
C10782 VDD.n1177 VSS 0.354217f
C10783 VDD.n1178 VSS 0.05616f
C10784 VDD.n1179 VSS 0.041264f
C10785 VDD.n1180 VSS 0.027622f
C10786 VDD.n1181 VSS 0.024192f
C10787 VDD.n1182 VSS -0.010928f
C10788 VDD.n1183 VSS 0.176997f
C10789 VDD.t682 VSS 0.230102f
C10790 VDD.t676 VSS 0.142531f
C10791 VDD.n1184 VSS 0.130881f
C10792 VDD.n1185 VSS 0.314521f
C10793 VDD.t31 VSS 0.32161f
C10794 VDD.t1457 VSS 0.302034f
C10795 VDD.t32 VSS 0.302034f
C10796 VDD.t1473 VSS 0.058729f
C10797 VDD.n1186 VSS 0.293716f
C10798 VDD.n1187 VSS 0.023676f
C10799 VDD.n1188 VSS 0.129048f
C10800 VDD.t1565 VSS 0.006764f
C10801 VDD.t1575 VSS 0.006764f
C10802 VDD.n1189 VSS 0.015166f
C10803 VDD.n1190 VSS 0.035907f
C10804 VDD.t1882 VSS 0.116433f
C10805 VDD.t1883 VSS 0.006764f
C10806 VDD.t1887 VSS 0.006764f
C10807 VDD.n1191 VSS 0.015166f
C10808 VDD.t1879 VSS 0.018322f
C10809 VDD.t255 VSS 0.018322f
C10810 VDD.t249 VSS 0.006764f
C10811 VDD.t253 VSS 0.006764f
C10812 VDD.n1192 VSS 0.015166f
C10813 VDD.t251 VSS 0.022391f
C10814 VDD.n1193 VSS 0.095048f
C10815 VDD.t1572 VSS 0.116433f
C10816 VDD.t1573 VSS 0.006764f
C10817 VDD.t1577 VSS 0.006764f
C10818 VDD.n1194 VSS 0.015166f
C10819 VDD.t1569 VSS 0.018322f
C10820 VDD.t1168 VSS 0.018322f
C10821 VDD.t1164 VSS 0.006764f
C10822 VDD.t1166 VSS 0.006764f
C10823 VDD.n1195 VSS 0.015166f
C10824 VDD.t1162 VSS 0.018322f
C10825 VDD.t1158 VSS 0.018422f
C10826 VDD.t1156 VSS 0.006764f
C10827 VDD.t1154 VSS 0.006764f
C10828 VDD.n1196 VSS 0.015166f
C10829 VDD.n1197 VSS 0.035894f
C10830 VDD.t1157 VSS 0.227678f
C10831 VDD.t1155 VSS 0.103398f
C10832 VDD.t1876 VSS 0.116433f
C10833 VDD.t1889 VSS 0.018322f
C10834 VDD.t1160 VSS 0.018313f
C10835 VDD.n1198 VSS 0.051521f
C10836 VDD.n1199 VSS 0.059268f
C10837 VDD.t1881 VSS 0.006764f
C10838 VDD.t1877 VSS 0.006764f
C10839 VDD.n1200 VSS 0.015166f
C10840 VDD.t1891 VSS 0.018322f
C10841 VDD.t257 VSS 0.018322f
C10842 VDD.n1201 VSS 0.046913f
C10843 VDD.t1890 VSS 0.230818f
C10844 VDD.t776 VSS 0.230818f
C10845 VDD.t777 VSS 0.147505f
C10846 VDD.t778 VSS 0.18404f
C10847 VDD.t262 VSS 0.114849f
C10848 VDD.t259 VSS 0.006764f
C10849 VDD.t263 VSS 0.006764f
C10850 VDD.n1202 VSS 0.015166f
C10851 VDD.t261 VSS 0.018322f
C10852 VDD.t1579 VSS 0.018322f
C10853 VDD.t1567 VSS 0.006764f
C10854 VDD.t1559 VSS 0.006764f
C10855 VDD.n1203 VSS 0.015166f
C10856 VDD.n1204 VSS 0.043025f
C10857 VDD.t260 VSS 0.213305f
C10858 VDD.t1578 VSS 0.216226f
C10859 VDD.t1566 VSS 0.104824f
C10860 VDD.t389 VSS 0.230818f
C10861 VDD.t390 VSS 0.147505f
C10862 VDD.t388 VSS 0.230818f
C10863 VDD.t1560 VSS 0.230818f
C10864 VDD.t1558 VSS 0.116433f
C10865 VDD.n1205 VSS 0.062021f
C10866 VDD.n1206 VSS -0.011488f
C10867 VDD.n1207 VSS 0.05616f
C10868 VDD.n1208 VSS 0.048865f
C10869 VDD.n1209 VSS 0.035907f
C10870 VDD.n1210 VSS -0.010928f
C10871 VDD.n1211 VSS 0.061018f
C10872 VDD.t258 VSS 0.103398f
C10873 VDD.t256 VSS 0.168918f
C10874 VDD.n1212 VSS 0.202202f
C10875 VDD.n1213 VSS 0.090004f
C10876 VDD.n1214 VSS 0.043025f
C10877 VDD.n1215 VSS -0.011488f
C10878 VDD.n1216 VSS 0.062021f
C10879 VDD.t1880 VSS 0.104824f
C10880 VDD.t1888 VSS 0.230818f
C10881 VDD.t1159 VSS 0.227678f
C10882 VDD.t1153 VSS 0.114849f
C10883 VDD.n1217 VSS 0.061018f
C10884 VDD.n1218 VSS -0.010928f
C10885 VDD.n1219 VSS 0.134973f
C10886 VDD.n1220 VSS 0.141428f
C10887 VDD.n1221 VSS 0.041121f
C10888 VDD.t1161 VSS 0.227678f
C10889 VDD.t1163 VSS 0.114849f
C10890 VDD.t1568 VSS 0.230818f
C10891 VDD.t378 VSS 0.230818f
C10892 VDD.t379 VSS 0.147505f
C10893 VDD.t380 VSS 0.230818f
C10894 VDD.t1167 VSS 0.227678f
C10895 VDD.t1165 VSS 0.103398f
C10896 VDD.n1222 VSS 0.061018f
C10897 VDD.n1223 VSS -0.010718f
C10898 VDD.t1926 VSS 0.006764f
C10899 VDD.t1928 VSS 0.006764f
C10900 VDD.n1224 VSS 0.018431f
C10901 VDD.t1930 VSS 0.006764f
C10902 VDD.t1931 VSS 0.006764f
C10903 VDD.n1225 VSS 0.013528f
C10904 VDD.n1226 VSS 0.032654f
C10905 VDD.n1227 VSS 0.058636f
C10906 VDD.n1228 VSS 0.494509f
C10907 VDD.n1229 VSS 0.074078f
C10908 VDD.n1230 VSS 0.090838f
C10909 VDD.n1231 VSS 0.043025f
C10910 VDD.t1581 VSS 0.022055f
C10911 VDD.n1232 VSS -0.011488f
C10912 VDD.n1233 VSS 0.062021f
C10913 VDD.t1576 VSS 0.104824f
C10914 VDD.t1580 VSS 0.283776f
C10915 VDD.t250 VSS 0.283492f
C10916 VDD.t248 VSS 0.116235f
C10917 VDD.t1878 VSS 0.230818f
C10918 VDD.t1610 VSS 0.230818f
C10919 VDD.t1611 VSS 0.147505f
C10920 VDD.t1612 VSS 0.214099f
C10921 VDD.t254 VSS 0.213738f
C10922 VDD.t252 VSS 0.104645f
C10923 VDD.n1234 VSS 0.061895f
C10924 VDD.n1235 VSS -0.010623f
C10925 VDD.n1236 VSS 0.086535f
C10926 VDD.n1237 VSS 0.089368f
C10927 VDD.n1238 VSS 0.043025f
C10928 VDD.t1885 VSS 0.018322f
C10929 VDD.t1563 VSS 0.018322f
C10930 VDD.n1239 VSS 0.050861f
C10931 VDD.n1240 VSS 0.058884f
C10932 VDD.n1241 VSS -0.011488f
C10933 VDD.n1242 VSS 0.062021f
C10934 VDD.t1886 VSS 0.104824f
C10935 VDD.t1884 VSS 0.222623f
C10936 VDD.t1562 VSS 0.222623f
C10937 VDD.t1564 VSS 0.116433f
C10938 VDD.t1570 VSS 0.230818f
C10939 VDD.t1574 VSS 0.104824f
C10940 VDD.n1243 VSS 0.062021f
C10941 VDD.n1244 VSS -0.010928f
C10942 VDD.t1571 VSS 0.018342f
C10943 VDD.n1245 VSS 0.044599f
C10944 VDD.n1246 VSS -0.078363f
C10945 VDD.n1247 VSS -0.108312f
C10946 VDD.n1248 VSS 0.069514f
C10947 VDD.n1249 VSS 0.036111f
C10948 VDD.t1938 VSS 0.006764f
C10949 VDD.t1796 VSS 0.006764f
C10950 VDD.n1250 VSS 0.014917f
C10951 VDD.t926 VSS 0.006764f
C10952 VDD.t1944 VSS 0.006764f
C10953 VDD.n1251 VSS 0.014917f
C10954 VDD.t924 VSS 0.022409f
C10955 VDD.n1252 VSS 0.096335f
C10956 VDD.n1253 VSS 0.033732f
C10957 VDD.t1812 VSS 0.018316f
C10958 VDD.n1254 VSS 0.096908f
C10959 VDD.n1255 VSS 0.07211f
C10960 VDD.n1256 VSS 0.033732f
C10961 VDD.n1257 VSS 0.0563f
C10962 VDD.n1258 VSS 0.056289f
C10963 VDD.n1259 VSS 0.032472f
C10964 VDD.n1260 VSS -0.002571f
C10965 VDD.n1261 VSS 0.189733f
C10966 VDD.t399 VSS 0.219141f
C10967 VDD.t610 VSS 0.408943f
C10968 VDD.n1262 VSS 0.356736f
C10969 VDD.t589 VSS 0.141408f
C10970 VDD.t587 VSS 0.136969f
C10971 VDD.t1149 VSS 0.136969f
C10972 VDD.t1151 VSS 0.136969f
C10973 VDD.t704 VSS 0.136969f
C10974 VDD.t702 VSS 0.214331f
C10975 VDD.t1776 VSS 0.363892f
C10976 VDD.t1784 VSS 0.138882f
C10977 VDD.t1778 VSS 0.341283f
C10978 VDD.n1263 VSS 0.102565f
C10979 VDD.n1264 VSS 0.004714f
C10980 VDD.t1810 VSS 0.01979f
C10981 VDD.t1779 VSS 0.01669f
C10982 VDD.n1265 VSS 0.045279f
C10983 VDD.n1266 VSS 0.109502f
C10984 VDD.t1209 VSS 0.028459f
C10985 VDD.t1215 VSS 0.006764f
C10986 VDD.t1213 VSS 0.006764f
C10987 VDD.n1267 VSS 0.015166f
C10988 VDD.t1211 VSS 0.028486f
C10989 VDD.n1268 VSS 0.034939f
C10990 VDD.t1208 VSS 0.227678f
C10991 VDD.t1214 VSS 0.114849f
C10992 VDD.t2156 VSS 0.104645f
C10993 VDD.t2155 VSS 0.006764f
C10994 VDD.t2157 VSS 0.006764f
C10995 VDD.n1269 VSS 0.015166f
C10996 VDD.t2151 VSS 0.022391f
C10997 VDD.n1270 VSS 0.095048f
C10998 VDD.t2153 VSS 0.018322f
C10999 VDD.t962 VSS 0.018322f
C11000 VDD.t966 VSS 0.006764f
C11001 VDD.t1893 VSS 0.006764f
C11002 VDD.n1271 VSS 0.015166f
C11003 VDD.t968 VSS 0.018322f
C11004 VDD.t838 VSS 0.018322f
C11005 VDD.n1272 VSS 0.050861f
C11006 VDD.n1273 VSS 0.058884f
C11007 VDD.t2152 VSS 0.213738f
C11008 VDD.t228 VSS 0.214099f
C11009 VDD.t229 VSS 0.147505f
C11010 VDD.t227 VSS 0.230818f
C11011 VDD.t961 VSS 0.230818f
C11012 VDD.t965 VSS 0.116433f
C11013 VDD.t837 VSS 0.219653f
C11014 VDD.t967 VSS 0.222676f
C11015 VDD.t1892 VSS 0.104824f
C11016 VDD.n1274 VSS 0.062021f
C11017 VDD.n1275 VSS -0.011488f
C11018 VDD.n1276 VSS 0.043025f
C11019 VDD.n1277 VSS 0.089368f
C11020 VDD.n1278 VSS 0.086535f
C11021 VDD.n1279 VSS -0.010623f
C11022 VDD.n1280 VSS 0.061895f
C11023 VDD.t2154 VSS 0.116235f
C11024 VDD.t2150 VSS 0.283492f
C11025 VDD.t885 VSS 0.283776f
C11026 VDD.t833 VSS 0.104824f
C11027 VDD.t824 VSS 0.006764f
C11028 VDD.t834 VSS 0.006764f
C11029 VDD.n1281 VSS 0.015166f
C11030 VDD.t1918 VSS 0.018322f
C11031 VDD.n1282 VSS 0.103562f
C11032 VDD.n1283 VSS 0.043025f
C11033 VDD.t886 VSS 0.022055f
C11034 VDD.n1284 VSS -0.011488f
C11035 VDD.n1285 VSS 0.062021f
C11036 VDD.t823 VSS 0.116433f
C11037 VDD.t1917 VSS 0.230818f
C11038 VDD.t89 VSS 0.230818f
C11039 VDD.t90 VSS 0.147505f
C11040 VDD.t91 VSS 0.230818f
C11041 VDD.t1210 VSS 0.227678f
C11042 VDD.t1212 VSS 0.103398f
C11043 VDD.n1286 VSS 0.061018f
C11044 VDD.n1287 VSS -0.01056f
C11045 VDD.n1288 VSS 0.034162f
C11046 VDD.n1289 VSS 0.214861f
C11047 VDD.n1290 VSS 0.137299f
C11048 VDD.t1470 VSS 0.227678f
C11049 VDD.t1459 VSS 0.103398f
C11050 VDD.t969 VSS 0.230818f
C11051 VDD.t1466 VSS 0.227678f
C11052 VDD.t1461 VSS 0.114849f
C11053 VDD.n1291 VSS 0.061018f
C11054 VDD.n1292 VSS -0.010928f
C11055 VDD.n1293 VSS 0.035894f
C11056 VDD.n1294 VSS 0.051521f
C11057 VDD.n1295 VSS 0.059268f
C11058 VDD.t960 VSS 0.006764f
C11059 VDD.t958 VSS 0.006764f
C11060 VDD.n1296 VSS 0.015166f
C11061 VDD.n1297 VSS 0.043025f
C11062 VDD.n1298 VSS -0.011488f
C11063 VDD.n1299 VSS 0.062021f
C11064 VDD.t957 VSS 0.116433f
C11065 VDD.t963 VSS 0.230818f
C11066 VDD.t1206 VSS 0.230818f
C11067 VDD.t1205 VSS 0.147505f
C11068 VDD.t1207 VSS 0.18404f
C11069 VDD.t788 VSS 0.168918f
C11070 VDD.n1300 VSS 0.202202f
C11071 VDD.n1301 VSS 0.046913f
C11072 VDD.t793 VSS 0.006764f
C11073 VDD.t791 VSS 0.006764f
C11074 VDD.n1302 VSS 0.015166f
C11075 VDD.t787 VSS 0.018322f
C11076 VDD.t895 VSS 0.018322f
C11077 VDD.n1303 VSS 0.05616f
C11078 VDD.n1304 VSS 0.048865f
C11079 VDD.n1305 VSS 0.035907f
C11080 VDD.n1306 VSS -0.010928f
C11081 VDD.n1307 VSS 0.061018f
C11082 VDD.t790 VSS 0.114849f
C11083 VDD.t786 VSS 0.213305f
C11084 VDD.t894 VSS 0.216226f
C11085 VDD.t873 VSS 0.104824f
C11086 VDD.t738 VSS 0.230818f
C11087 VDD.t736 VSS 0.147505f
C11088 VDD.t737 VSS 0.230818f
C11089 VDD.t839 VSS 0.230818f
C11090 VDD.t819 VSS 0.116433f
C11091 VDD.n1308 VSS 0.062021f
C11092 VDD.n1309 VSS -0.011488f
C11093 VDD.n1310 VSS 0.043025f
C11094 VDD.n1311 VSS -0.141053f
C11095 VDD.n1312 VSS -0.114529f
C11096 VDD.n1313 VSS -0.010928f
C11097 VDD.n1314 VSS 0.061018f
C11098 VDD.t815 VSS 0.103398f
C11099 VDD.t853 VSS 0.545618f
C11100 VDD.t1015 VSS 0.545618f
C11101 VDD.t1011 VSS 0.114849f
C11102 VDD.t863 VSS 0.230818f
C11103 VDD.t1020 VSS 0.230818f
C11104 VDD.t1019 VSS 0.147505f
C11105 VDD.t1021 VSS 0.230818f
C11106 VDD.t1017 VSS 0.227678f
C11107 VDD.t1013 VSS 0.103398f
C11108 VDD.n1315 VSS 0.061018f
C11109 VDD.n1316 VSS -0.01056f
C11110 VDD.n1317 VSS 0.103562f
C11111 VDD.n1318 VSS 0.043025f
C11112 VDD.t822 VSS 0.022055f
C11113 VDD.n1319 VSS -0.011488f
C11114 VDD.n1320 VSS 0.062021f
C11115 VDD.t1896 VSS 0.104824f
C11116 VDD.t821 VSS 0.283776f
C11117 VDD.t798 VSS 0.283492f
C11118 VDD.t800 VSS 0.116235f
C11119 VDD.t1494 VSS 0.230818f
C11120 VDD.t149 VSS 0.230818f
C11121 VDD.t150 VSS 0.147505f
C11122 VDD.t151 VSS 0.214099f
C11123 VDD.t794 VSS 0.213738f
C11124 VDD.t796 VSS 0.104645f
C11125 VDD.n1321 VSS 0.061895f
C11126 VDD.n1322 VSS -0.010623f
C11127 VDD.n1323 VSS 0.086535f
C11128 VDD.n1324 VSS 0.089368f
C11129 VDD.n1325 VSS 0.043025f
C11130 VDD.t1501 VSS 0.018322f
C11131 VDD.t1914 VSS 0.018322f
C11132 VDD.n1326 VSS 0.050861f
C11133 VDD.n1327 VSS 0.058884f
C11134 VDD.n1328 VSS -0.011488f
C11135 VDD.n1329 VSS 0.062021f
C11136 VDD.t1498 VSS 0.104824f
C11137 VDD.t1500 VSS 0.222676f
C11138 VDD.t1913 VSS 0.219653f
C11139 VDD.t1911 VSS 0.114849f
C11140 VDD.t857 VSS 0.227678f
C11141 VDD.t817 VSS 0.103398f
C11142 VDD.n1330 VSS 0.061018f
C11143 VDD.n1331 VSS -0.010928f
C11144 VDD.t858 VSS 0.018342f
C11145 VDD.n1332 VSS 0.0446f
C11146 VDD.n1333 VSS -0.178123f
C11147 VDD.t219 VSS 0.027971f
C11148 VDD.n1334 VSS 0.043291f
C11149 VDD.n1335 VSS 0.031509f
C11150 VDD.n1336 VSS 0.044892f
C11151 VDD.n1337 VSS 0.027244f
C11152 VDD.t125 VSS 0.006764f
C11153 VDD.t308 VSS 0.006764f
C11154 VDD.n1338 VSS 0.029826f
C11155 VDD.t741 VSS 0.006764f
C11156 VDD.t2070 VSS 0.006764f
C11157 VDD.n1339 VSS 0.013528f
C11158 VDD.n1340 VSS 0.039293f
C11159 VDD.t126 VSS 0.006764f
C11160 VDD.t307 VSS 0.006764f
C11161 VDD.n1341 VSS 0.029015f
C11162 VDD.n1342 VSS 0.03765f
C11163 VDD.t740 VSS 0.006764f
C11164 VDD.t2071 VSS 0.006764f
C11165 VDD.n1343 VSS 0.013528f
C11166 VDD.n1344 VSS 0.008042f
C11167 VDD.n1345 VSS 0.027244f
C11168 VDD.n1346 VSS 0.04544f
C11169 VDD.t213 VSS 0.027971f
C11170 VDD.t215 VSS 0.034731f
C11171 VDD.n1347 VSS 0.044989f
C11172 VDD.n1348 VSS 0.074425f
C11173 VDD.n1349 VSS 0.065197f
C11174 VDD.n1350 VSS 0.099614f
C11175 VDD.t121 VSS 0.197636f
C11176 VDD.t742 VSS 0.760366f
C11177 VDD.t214 VSS 0.835558f
C11178 VDD.t739 VSS 0.331315f
C11179 VDD.t2069 VSS 0.185802f
C11180 VDD.t306 VSS 0.400006f
C11181 VDD.t124 VSS 0.197636f
C11182 VDD.n1351 VSS 0.099614f
C11183 VDD.n1352 VSS 0.021675f
C11184 VDD.n1353 VSS 0.075906f
C11185 VDD.n1354 VSS 0.099889f
C11186 VDD.n1355 VSS 0.013114f
C11187 VDD.n1356 VSS 0.193277f
C11188 VDD.t1257 VSS 0.146509f
C11189 VDD.t1238 VSS 0.114849f
C11190 VDD.t2058 VSS 0.3011f
C11191 VDD.t1255 VSS 0.3011f
C11192 VDD.t1247 VSS 0.103398f
C11193 VDD.n1357 VSS 0.061018f
C11194 VDD.n1358 VSS 0.020137f
C11195 VDD.n1359 VSS 0.063729f
C11196 VDD.n1360 VSS 0.061018f
C11197 VDD.t2038 VSS 0.103398f
C11198 VDD.t2050 VSS 0.229878f
C11199 VDD.t372 VSS 0.409363f
C11200 VDD.t373 VSS 0.259137f
C11201 VDD.t325 VSS 0.259137f
C11202 VDD.t323 VSS 0.310025f
C11203 VDD.t1839 VSS 0.146509f
C11204 VDD.n1361 VSS 0.193277f
C11205 VDD.n1362 VSS 0.035024f
C11206 VDD.n1363 VSS 0.020137f
C11207 VDD.n1364 VSS 0.061018f
C11208 VDD.t1855 VSS 0.103398f
C11209 VDD.t1837 VSS 0.269441f
C11210 VDD.t2088 VSS 0.269441f
C11211 VDD.t2092 VSS 0.114849f
C11212 VDD.t804 VSS 0.259137f
C11213 VDD.t547 VSS 0.259137f
C11214 VDD.t546 VSS 0.409363f
C11215 VDD.t2086 VSS 0.229878f
C11216 VDD.t2072 VSS 0.103398f
C11217 VDD.n1365 VSS 0.061018f
C11218 VDD.n1366 VSS 0.058379f
C11219 VDD.n1367 VSS 0.102239f
C11220 VDD.n1368 VSS 0.013114f
C11221 VDD.n1369 VSS 0.193277f
C11222 VDD.t1674 VSS 0.146509f
C11223 VDD.t1682 VSS 0.114849f
C11224 VDD.t1678 VSS 0.227678f
C11225 VDD.t1671 VSS 0.103398f
C11226 VDD.n1370 VSS 0.061018f
C11227 VDD.n1371 VSS 0.020137f
C11228 VDD.n1372 VSS 0.18346f
C11229 VDD.n1373 VSS 0.47366f
C11230 VDD.n1374 VSS -0.01053f
C11231 VDD.n1375 VSS 0.061018f
C11232 VDD.t2137 VSS 0.114849f
C11233 VDD.t2142 VSS 0.146509f
C11234 VDD.n1376 VSS 0.193277f
C11235 VDD.n1377 VSS 0.017781f
C11236 VDD.n1378 VSS 0.078479f
C11237 VDD.n1379 VSS 0.102669f
C11238 VDD.n1380 VSS -0.010519f
C11239 VDD.n1381 VSS 0.061018f
C11240 VDD.t1806 VSS 0.114849f
C11241 VDD.t1791 VSS 0.269441f
C11242 VDD.t1431 VSS 0.269441f
C11243 VDD.t1444 VSS 0.103398f
C11244 VDD.n1382 VSS 0.061018f
C11245 VDD.n1383 VSS -0.01053f
C11246 VDD.n1384 VSS 0.045731f
C11247 VDD.n1385 VSS 0.058631f
C11248 VDD.n1386 VSS 0.017781f
C11249 VDD.n1387 VSS 0.193277f
C11250 VDD.t173 VSS 0.310025f
C11251 VDD.t175 VSS 0.259137f
C11252 VDD.t108 VSS 0.259137f
C11253 VDD.t107 VSS 0.409363f
C11254 VDD.t1961 VSS 0.229878f
C11255 VDD.t1957 VSS 0.103398f
C11256 VDD.n1388 VSS 0.061018f
C11257 VDD.n1389 VSS -0.010519f
C11258 VDD.n1390 VSS 0.046076f
C11259 VDD.n1391 VSS 0.075269f
C11260 VDD.n1392 VSS 0.073705f
C11261 VDD.n1393 VSS -0.01053f
C11262 VDD.n1394 VSS 0.061018f
C11263 VDD.t2012 VSS 0.114849f
C11264 VDD.t2007 VSS 0.146509f
C11265 VDD.n1395 VSS 0.193277f
C11266 VDD.n1396 VSS 0.017781f
C11267 VDD.n1397 VSS 0.078479f
C11268 VDD.n1398 VSS 0.102669f
C11269 VDD.n1399 VSS -0.010519f
C11270 VDD.n1400 VSS 0.061018f
C11271 VDD.t1825 VSS 0.114849f
C11272 VDD.t1821 VSS 0.321982f
C11273 VDD.t1548 VSS 0.321982f
C11274 VDD.t1534 VSS 0.103398f
C11275 VDD.n1401 VSS 0.061018f
C11276 VDD.n1402 VSS -0.01053f
C11277 VDD.n1403 VSS 0.045731f
C11278 VDD.n1404 VSS 0.058631f
C11279 VDD.n1405 VSS 0.017772f
C11280 VDD.n1406 VSS 0.193277f
C11281 VDD.t138 VSS 0.310025f
C11282 VDD.t140 VSS 0.259137f
C11283 VDD.t407 VSS 0.259137f
C11284 VDD.t408 VSS 0.409363f
C11285 VDD.t1175 VSS 0.229878f
C11286 VDD.t1185 VSS 0.103398f
C11287 VDD.n1407 VSS 0.061018f
C11288 VDD.n1408 VSS -0.010519f
C11289 VDD.n1409 VSS 0.046076f
C11290 VDD.n1410 VSS 0.072611f
C11291 VDD.n1411 VSS 0.058754f
C11292 VDD.n1412 VSS 0.034926f
C11293 VDD.n1413 VSS 0.038435f
C11294 VDD.n1414 VSS 0.031626f
C11295 VDD.n1415 VSS 2.89099f
C11296 VDD.n1416 VSS 1.57773f
C11297 VDD.n1417 VSS 0.028993f
C11298 VDD.n1418 VSS 0.019902f
C11299 VDD.n1419 VSS 0.017552f
C11300 VDD.n1420 VSS 0.017552f
C11301 VDD.n1421 VSS 0.019487f
C11302 VDD.n1422 VSS 0.068756f
C11303 VDD.n1423 VSS 0.020531f
C11304 VDD.n1424 VSS 0.020242f
C11305 VDD.n1425 VSS 0.017137f
C11306 VDD.n1426 VSS 0.052094f
C11307 VDD.n1427 VSS 0.016155f
C11308 VDD.n1428 VSS 0.015487f
C11309 VDD.n1429 VSS 0.031018f
C11310 VDD.n1430 VSS 0.019902f
C11311 VDD.n1431 VSS 0.027927f
C11312 VDD.n1432 VSS 0.001662f
C11313 VDD.n1433 VSS 0.001938f
C11314 VDD.n1434 VSS 0.019349f
C11315 VDD.n1435 VSS 0.019625f
C11316 VDD.n1436 VSS 0.021051f
C11317 VDD.n1437 VSS 2.5771f
C11318 VDD.n1438 VSS 0.028993f
C11319 VDD.n1439 VSS 0.027927f
C11320 VDD.n1440 VSS 1.49902f
C11321 VDD.n1441 VSS 0.039887f
C11322 VDD.n1442 VSS 0.039055f
C11323 VDD.n1443 VSS 0.019487f
C11324 VDD.n1444 VSS 0.019487f
C11325 VDD.n1445 VSS 0.019625f
C11326 VDD.n1446 VSS 0.020531f
C11327 VDD.n1447 VSS 0.020242f
C11328 VDD.n1448 VSS 0.052094f
C11329 VDD.n1449 VSS 0.016155f
C11330 VDD.n1450 VSS 0.015495f
C11331 VDD.n1451 VSS 0.088624f
C11332 VDD.n1452 VSS 0.017137f
C11333 VDD.n1453 VSS 0.019349f
C11334 VDD.n1454 VSS 0.00637f
C11335 VDD.n1455 VSS 1.62039f
C11336 VDD.n1456 VSS 4.27303f
C11337 VDD.n1457 VSS 4.10097f
C11338 VDD.n1458 VSS 1.80749f
C11339 VDD.n1459 VSS 0.075391f
C11340 VDD.t1752 VSS 0.214331f
C11341 VDD.t1758 VSS 0.136969f
C11342 VDD.t1403 VSS 0.136969f
C11343 VDD.t1401 VSS 0.136969f
C11344 VDD.t327 VSS 0.136969f
C11345 VDD.t329 VSS 0.214331f
C11346 VDD.t283 VSS 0.16801f
C11347 VDD.t1597 VSS 0.080526f
C11348 VDD.t1599 VSS 0.194852f
C11349 VDD.t1736 VSS 0.363892f
C11350 VDD.t487 VSS 0.214331f
C11351 VDD.t485 VSS 0.136969f
C11352 VDD.t669 VSS 0.136969f
C11353 VDD.t667 VSS 0.136969f
C11354 VDD.t491 VSS 0.136969f
C11355 VDD.t489 VSS 0.214331f
C11356 VDD.t287 VSS 0.451822f
C11357 VDD.t285 VSS 0.159741f
C11358 VDD.t284 VSS 0.021269f
C11359 VDD.t288 VSS 0.01669f
C11360 VDD.n1460 VSS 0.070928f
C11361 VDD.t289 VSS 0.006764f
C11362 VDD.t286 VSS 0.006764f
C11363 VDD.n1461 VSS 0.013528f
C11364 VDD.n1462 VSS 0.036172f
C11365 VDD.t490 VSS 0.018157f
C11366 VDD.t486 VSS 0.006764f
C11367 VDD.t670 VSS 0.006764f
C11368 VDD.n1463 VSS 0.022549f
C11369 VDD.t668 VSS 0.006764f
C11370 VDD.t492 VSS 0.006764f
C11371 VDD.n1464 VSS 0.022549f
C11372 VDD.n1465 VSS 0.057655f
C11373 VDD.n1466 VSS 0.066276f
C11374 VDD.n1467 VSS 0.032472f
C11375 VDD.t1600 VSS 0.021269f
C11376 VDD.t1598 VSS 0.01669f
C11377 VDD.n1468 VSS 0.084502f
C11378 VDD.n1469 VSS -0.002571f
C11379 VDD.n1470 VSS 0.063865f
C11380 VDD.n1471 VSS 0.236364f
C11381 VDD.t1596 VSS 0.216554f
C11382 VDD.t1595 VSS 1.06616f
C11383 VDD.t61 VSS 1.06535f
C11384 VDD.t458 VSS 0.288488f
C11385 VDD.t460 VSS 0.162942f
C11386 VDD.t1193 VSS 0.162942f
C11387 VDD.t1199 VSS 0.146247f
C11388 VDD.t20 VSS 0.195308f
C11389 VDD.t1360 VSS 0.214331f
C11390 VDD.t1334 VSS 0.136969f
C11391 VDD.t1949 VSS 0.136969f
C11392 VDD.t1969 VSS 0.136969f
C11393 VDD.t136 VSS 0.136969f
C11394 VDD.t134 VSS 0.214331f
C11395 VDD.t920 VSS 0.168403f
C11396 VDD.t16 VSS 0.080714f
C11397 VDD.t18 VSS 0.159603f
C11398 VDD.t21 VSS 0.021269f
C11399 VDD.t19 VSS 0.01669f
C11400 VDD.n1472 VSS 0.068817f
C11401 VDD.t1198 VSS 0.017784f
C11402 VDD.t1605 VSS 0.006764f
C11403 VDD.t1196 VSS 0.006764f
C11404 VDD.n1473 VSS 0.020425f
C11405 VDD.n1474 VSS 0.059702f
C11406 VDD.t1601 VSS 0.01669f
C11407 VDD.n1475 VSS 0.017903f
C11408 VDD.t1604 VSS 0.006764f
C11409 VDD.t1602 VSS 0.006764f
C11410 VDD.n1476 VSS 0.020425f
C11411 VDD.n1477 VSS 0.039154f
C11412 VDD.n1478 VSS 0.087529f
C11413 VDD.n1479 VSS 0.07375f
C11414 VDD.t921 VSS 0.021269f
C11415 VDD.t918 VSS 0.01669f
C11416 VDD.n1480 VSS 0.070928f
C11417 VDD.t922 VSS 0.006764f
C11418 VDD.t919 VSS 0.006764f
C11419 VDD.n1481 VSS 0.013528f
C11420 VDD.n1482 VSS 0.036172f
C11421 VDD.t916 VSS 0.018157f
C11422 VDD.t914 VSS 0.006764f
C11423 VDD.t60 VSS 0.006764f
C11424 VDD.n1483 VSS 0.022549f
C11425 VDD.t65 VSS 0.006764f
C11426 VDD.t496 VSS 0.006764f
C11427 VDD.n1484 VSS 0.022549f
C11428 VDD.t1383 VSS 0.006764f
C11429 VDD.t1332 VSS 0.006764f
C11430 VDD.n1485 VSS 0.01683f
C11431 VDD.t1324 VSS 0.006764f
C11432 VDD.t1356 VSS 0.006764f
C11433 VDD.n1486 VSS 0.013528f
C11434 VDD.n1487 VSS 0.030751f
C11435 VDD.n1488 VSS 0.01223f
C11436 VDD.t1343 VSS 0.01979f
C11437 VDD.t1381 VSS 0.01669f
C11438 VDD.n1489 VSS 0.049398f
C11439 VDD.n1490 VSS 0.03223f
C11440 VDD.n1491 VSS 0.014255f
C11441 VDD.t917 VSS 0.45143f
C11442 VDD.t915 VSS 0.214331f
C11443 VDD.t913 VSS 0.136969f
C11444 VDD.t59 VSS 0.136969f
C11445 VDD.t64 VSS 0.136969f
C11446 VDD.t495 VSS 0.136969f
C11447 VDD.t493 VSS 0.214331f
C11448 VDD.t1323 VSS 0.251925f
C11449 VDD.t1342 VSS 0.341283f
C11450 VDD.n1492 VSS 0.116273f
C11451 VDD.t1331 VSS 0.134575f
C11452 VDD.n1493 VSS 0.116273f
C11453 VDD.n1494 VSS 0.016579f
C11454 VDD.t494 VSS 0.018172f
C11455 VDD.n1495 VSS 0.038281f
C11456 VDD.t137 VSS 0.006764f
C11457 VDD.t1970 VSS 0.006764f
C11458 VDD.n1496 VSS 0.022549f
C11459 VDD.t1950 VSS 0.006764f
C11460 VDD.t1335 VSS 0.006764f
C11461 VDD.n1497 VSS 0.022549f
C11462 VDD.t135 VSS 0.025643f
C11463 VDD.n1498 VSS 0.104443f
C11464 VDD.t1361 VSS 0.018316f
C11465 VDD.n1499 VSS 0.097077f
C11466 VDD.n1500 VSS 0.073072f
C11467 VDD.n1501 VSS 0.057655f
C11468 VDD.n1502 VSS 0.066276f
C11469 VDD.n1503 VSS 0.032472f
C11470 VDD.n1504 VSS -0.002571f
C11471 VDD.n1505 VSS 0.063804f
C11472 VDD.n1506 VSS 0.236503f
C11473 VDD.t15 VSS 0.216366f
C11474 VDD.t17 VSS 0.726829f
C11475 VDD.t1197 VSS 0.726829f
C11476 VDD.t1195 VSS 0.288488f
C11477 VDD.t1603 VSS 0.288488f
C11478 VDD.t1194 VSS 0.286484f
C11479 VDD.n1507 VSS -0.007463f
C11480 VDD.n1508 VSS -0.143553f
C11481 VDD.n1509 VSS 0.235278f
C11482 VDD.t1952 VSS 0.006764f
C11483 VDD.t1337 VSS 0.006764f
C11484 VDD.n1510 VSS 0.014917f
C11485 VDD.t724 VSS 0.006764f
C11486 VDD.t1972 VSS 0.006764f
C11487 VDD.n1511 VSS 0.014917f
C11488 VDD.t726 VSS 0.022409f
C11489 VDD.n1512 VSS 0.096335f
C11490 VDD.n1513 VSS 0.033732f
C11491 VDD.t1365 VSS 0.018316f
C11492 VDD.n1514 VSS 0.044404f
C11493 VDD.n1515 VSS 0.378059f
C11494 VDD.n1516 VSS 0.032867f
C11495 VDD.n1517 VSS 0.037558f
C11496 VDD.n1518 VSS 0.015175f
C11497 VDD.t1355 VSS 0.01979f
C11498 VDD.t1348 VSS 0.01669f
C11499 VDD.n1519 VSS 0.040346f
C11500 VDD.t592 VSS 0.021269f
C11501 VDD.t593 VSS 0.01669f
C11502 VDD.n1520 VSS 0.068817f
C11503 VDD.t630 VSS 0.021269f
C11504 VDD.t633 VSS 0.01669f
C11505 VDD.n1521 VSS 0.070928f
C11506 VDD.t628 VSS 0.006764f
C11507 VDD.t632 VSS 0.006764f
C11508 VDD.n1522 VSS 0.013528f
C11509 VDD.n1523 VSS 0.036172f
C11510 VDD.n1524 VSS 0.032472f
C11511 VDD.t591 VSS 0.175276f
C11512 VDD.t1349 VSS 0.214331f
C11513 VDD.t1312 VSS 0.136969f
C11514 VDD.t883 VSS 0.136969f
C11515 VDD.t869 VSS 0.136969f
C11516 VDD.t57 VSS 0.136969f
C11517 VDD.t55 VSS 0.214331f
C11518 VDD.t629 VSS 0.151131f
C11519 VDD.t401 VSS 0.072435f
C11520 VDD.t1347 VSS 1.19091f
C11521 VDD.t404 VSS 1.5616f
C11522 VDD.t403 VSS 0.420878f
C11523 VDD.t749 VSS 0.195308f
C11524 VDD.t1362 VSS 0.214331f
C11525 VDD.t1338 VSS 0.136969f
C11526 VDD.t1171 VSS 0.136969f
C11527 VDD.t1189 VSS 0.136969f
C11528 VDD.t321 VSS 0.136969f
C11529 VDD.t319 VSS 0.214331f
C11530 VDD.t930 VSS 0.168403f
C11531 VDD.t748 VSS 0.080714f
C11532 VDD.n1526 VSS 0.152698f
C11533 VDD.n1527 VSS 0.459347f
C11534 VDD.t750 VSS 0.021269f
C11535 VDD.t751 VSS 0.01669f
C11536 VDD.n1529 VSS 0.068817f
C11537 VDD.t2027 VSS 0.017784f
C11538 VDD.t440 VSS 0.006764f
C11539 VDD.t2024 VSS 0.006764f
C11540 VDD.n1530 VSS 0.020425f
C11541 VDD.n1531 VSS 0.059702f
C11542 VDD.t439 VSS 0.01669f
C11543 VDD.n1532 VSS 0.017903f
C11544 VDD.t437 VSS 0.006764f
C11545 VDD.t442 VSS 0.006764f
C11546 VDD.n1533 VSS 0.020425f
C11547 VDD.n1534 VSS 0.039154f
C11548 VDD.n1535 VSS 0.087187f
C11549 VDD.n1536 VSS 0.07375f
C11550 VDD.t931 VSS 0.021269f
C11551 VDD.t928 VSS 0.01669f
C11552 VDD.n1537 VSS 0.070928f
C11553 VDD.t927 VSS 0.006764f
C11554 VDD.t929 VSS 0.006764f
C11555 VDD.n1538 VSS 0.013528f
C11556 VDD.n1539 VSS 0.036172f
C11557 VDD.t387 VSS 0.018157f
C11558 VDD.t385 VSS 0.006764f
C11559 VDD.t1866 VSS 0.006764f
C11560 VDD.n1540 VSS 0.022549f
C11561 VDD.t1867 VSS 0.006764f
C11562 VDD.t267 VSS 0.006764f
C11563 VDD.n1541 VSS 0.022549f
C11564 VDD.t265 VSS 0.018172f
C11565 VDD.n1542 VSS 0.034494f
C11566 VDD.t402 VSS 0.360697f
C11567 VDD.t631 VSS 0.982939f
C11568 VDD.t386 VSS 0.518948f
C11569 VDD.t384 VSS 0.331635f
C11570 VDD.t1446 VSS 0.331635f
C11571 VDD.t1449 VSS 0.331635f
C11572 VDD.t266 VSS 0.331635f
C11573 VDD.t264 VSS 0.518948f
C11574 VDD.t1375 VSS 0.359272f
C11575 VDD.t1379 VSS 0.149561f
C11576 VDD.t1327 VSS 0.149561f
C11577 VDD.t1369 VSS 0.149561f
C11578 VDD.t1317 VSS 0.149561f
C11579 VDD.t1325 VSS 0.486435f
C11580 VDD.t1380 VSS 0.006764f
C11581 VDD.t1322 VSS 0.006764f
C11582 VDD.n1543 VSS 0.01683f
C11583 VDD.t1376 VSS 0.006764f
C11584 VDD.t1321 VSS 0.006764f
C11585 VDD.n1544 VSS 0.013528f
C11586 VDD.n1545 VSS 0.027737f
C11587 VDD.t727 VSS 0.018157f
C11588 VDD.t1450 VSS 0.006764f
C11589 VDD.t728 VSS 0.006764f
C11590 VDD.n1546 VSS 0.014917f
C11591 VDD.t729 VSS 0.006764f
C11592 VDD.t1447 VSS 0.006764f
C11593 VDD.n1547 VSS 0.014917f
C11594 VDD.t730 VSS 0.018157f
C11595 VDD.n1548 VSS 0.056289f
C11596 VDD.n1549 VSS 0.0563f
C11597 VDD.n1550 VSS 0.033732f
C11598 VDD.t884 VSS 0.006764f
C11599 VDD.t1313 VSS 0.006764f
C11600 VDD.n1551 VSS 0.014917f
C11601 VDD.t58 VSS 0.006764f
C11602 VDD.t870 VSS 0.006764f
C11603 VDD.n1552 VSS 0.014917f
C11604 VDD.t56 VSS 0.022409f
C11605 VDD.n1553 VSS 0.096335f
C11606 VDD.n1554 VSS 0.033732f
C11607 VDD.t1350 VSS 0.018316f
C11608 VDD.n1555 VSS 0.096908f
C11609 VDD.n1556 VSS 0.07211f
C11610 VDD.n1557 VSS 0.037558f
C11611 VDD.n1558 VSS 0.008485f
C11612 VDD.t1370 VSS 0.006764f
C11613 VDD.t1307 VSS 0.006764f
C11614 VDD.n1559 VSS 0.01683f
C11615 VDD.t1384 VSS 0.006764f
C11616 VDD.t1333 VSS 0.006764f
C11617 VDD.n1560 VSS 0.013528f
C11618 VDD.n1561 VSS 0.033163f
C11619 VDD.n1562 VSS 0.003205f
C11620 VDD.t1318 VSS 0.01979f
C11621 VDD.t1346 VSS 0.01669f
C11622 VDD.n1563 VSS 0.049398f
C11623 VDD.n1564 VSS 0.03223f
C11624 VDD.n1565 VSS 0.025683f
C11625 VDD.n1566 VSS 0.023493f
C11626 VDD.t1328 VSS 0.01979f
C11627 VDD.t1326 VSS 0.01669f
C11628 VDD.n1567 VSS 0.049398f
C11629 VDD.n1568 VSS 0.018476f
C11630 VDD.n1569 VSS 0.15211f
C11631 VDD.t1306 VSS 0.383073f
C11632 VDD.n1570 VSS 0.165818f
C11633 VDD.n1571 VSS 0.016853f
C11634 VDD.n1572 VSS 0.038281f
C11635 VDD.t322 VSS 0.006764f
C11636 VDD.t1190 VSS 0.006764f
C11637 VDD.n1573 VSS 0.022549f
C11638 VDD.t1172 VSS 0.006764f
C11639 VDD.t1339 VSS 0.006764f
C11640 VDD.n1574 VSS 0.022549f
C11641 VDD.t320 VSS 0.025643f
C11642 VDD.n1575 VSS 0.104443f
C11643 VDD.t1363 VSS 0.018316f
C11644 VDD.n1576 VSS 0.097077f
C11645 VDD.n1577 VSS 0.073072f
C11646 VDD.n1578 VSS 0.057655f
C11647 VDD.n1579 VSS 0.066276f
C11648 VDD.n1580 VSS 0.032472f
C11649 VDD.n1581 VSS -0.002571f
C11650 VDD.n1582 VSS 0.123655f
C11651 VDD.n1583 VSS -0.002571f
C11652 VDD.n1584 VSS 0.072393f
C11653 VDD.n1585 VSS 0.037945f
C11654 VDD.n1586 VSS 0.006361f
C11655 VDD.n1587 VSS 0.271638f
C11656 VDD.t1308 VSS 0.060284f
C11657 VDD.t441 VSS 0.289364f
C11658 VDD.t1371 VSS 0.289364f
C11659 VDD.t436 VSS 0.293384f
C11660 VDD.t2023 VSS 0.53864f
C11661 VDD.n1588 VSS 0.083684f
C11662 VDD.n1589 VSS -0.14321f
C11663 VDD.n1590 VSS 0.235278f
C11664 VDD.t1174 VSS 0.006764f
C11665 VDD.t1345 VSS 0.006764f
C11666 VDD.n1591 VSS 0.014917f
C11667 VDD.t1553 VSS 0.006764f
C11668 VDD.t1192 VSS 0.006764f
C11669 VDD.n1592 VSS 0.014917f
C11670 VDD.t1551 VSS 0.022409f
C11671 VDD.n1593 VSS 0.096335f
C11672 VDD.n1594 VSS 0.033732f
C11673 VDD.t1367 VSS 0.018316f
C11674 VDD.n1595 VSS 0.044404f
C11675 VDD.n1596 VSS 0.378059f
C11676 VDD.n1597 VSS 0.032867f
C11677 VDD.n1598 VSS 0.033732f
C11678 VDD.n1599 VSS 0.0563f
C11679 VDD.n1600 VSS 0.056289f
C11680 VDD.n1601 VSS 0.032472f
C11681 VDD.n1602 VSS -0.002571f
C11682 VDD.n1603 VSS 0.063804f
C11683 VDD.n1604 VSS 0.236503f
C11684 VDD.t659 VSS 0.216366f
C11685 VDD.t311 VSS 1.06513f
C11686 VDD.t991 VSS 1.06513f
C11687 VDD.t655 VSS 0.288488f
C11688 VDD.t657 VSS 0.162942f
C11689 VDD.t2121 VSS 0.162942f
C11690 VDD.t2122 VSS 0.146247f
C11691 VDD.n1605 VSS -0.007463f
C11692 VDD.n1606 VSS -0.085172f
C11693 VDD.n1607 VSS 0.235291f
C11694 VDD.n1608 VSS 0.378039f
C11695 VDD.n1609 VSS 0.033043f
C11696 VDD.n1610 VSS 0.057655f
C11697 VDD.n1611 VSS 0.066276f
C11698 VDD.n1612 VSS 0.032472f
C11699 VDD.t168 VSS 0.021269f
C11700 VDD.t169 VSS 0.01669f
C11701 VDD.n1613 VSS 0.084502f
C11702 VDD.n1614 VSS -0.002571f
C11703 VDD.n1615 VSS 0.112532f
C11704 VDD.t582 VSS 0.267439f
C11705 VDD.t584 VSS 0.756439f
C11706 VDD.t576 VSS 0.756439f
C11707 VDD.t578 VSS 0.480047f
C11708 VDD.t50 VSS 0.241701f
C11709 VDD.t604 VSS 0.241701f
C11710 VDD.t618 VSS 0.241701f
C11711 VDD.t602 VSS 0.241701f
C11712 VDD.t620 VSS 0.241701f
C11713 VDD.t523 VSS 0.031331f
C11714 VDD.t197 VSS 0.241701f
C11715 VDD.t525 VSS 0.241701f
C11716 VDD.t203 VSS 0.031331f
C11717 VDD.n1616 VSS 0.083806f
C11718 VDD.n1617 VSS -0.126148f
C11719 VDD.n1618 VSS 0.235291f
C11720 VDD.t1753 VSS 0.018316f
C11721 VDD.t1759 VSS 0.006764f
C11722 VDD.t1404 VSS 0.006764f
C11723 VDD.n1619 VSS 0.022549f
C11724 VDD.t1402 VSS 0.006764f
C11725 VDD.t328 VSS 0.006764f
C11726 VDD.n1620 VSS 0.022549f
C11727 VDD.t330 VSS 0.025643f
C11728 VDD.n1621 VSS 0.104443f
C11729 VDD.n1622 VSS 0.044574f
C11730 VDD.n1623 VSS 0.378039f
C11731 VDD.n1624 VSS 0.033043f
C11732 VDD.n1625 VSS 0.037558f
C11733 VDD.n1626 VSS 0.015175f
C11734 VDD.n1627 VSS 0.006361f
C11735 VDD.n1628 VSS 0.102565f
C11736 VDD.t1748 VSS 0.548156f
C11737 VDD.t45 VSS 0.882358f
C11738 VDD.t43 VSS 0.375016f
C11739 VDD.n1629 VSS 0.189733f
C11740 VDD.n1630 VSS -0.002571f
C11741 VDD.n1631 VSS 0.032472f
C11742 VDD.n1632 VSS 0.066276f
C11743 VDD.n1633 VSS 0.057655f
C11744 VDD.t1725 VSS 0.018316f
C11745 VDD.t1761 VSS 0.006764f
C11746 VDD.t880 VSS 0.006764f
C11747 VDD.n1634 VSS 0.022549f
C11748 VDD.t846 VSS 0.006764f
C11749 VDD.t2020 VSS 0.006764f
C11750 VDD.n1635 VSS 0.022549f
C11751 VDD.t2022 VSS 0.025643f
C11752 VDD.n1636 VSS 0.104443f
C11753 VDD.n1637 VSS 0.097077f
C11754 VDD.n1638 VSS 0.072279f
C11755 VDD.n1639 VSS 0.037558f
C11756 VDD.n1640 VSS 0.015175f
C11757 VDD.n1641 VSS 0.018755f
C11758 VDD.n1642 VSS 0.102565f
C11759 VDD.t1746 VSS 0.471552f
C11760 VDD.t1710 VSS 0.471552f
C11761 VDD.t1751 VSS 0.006764f
C11762 VDD.t1757 VSS 0.006764f
C11763 VDD.n1643 VSS 0.01683f
C11764 VDD.t1727 VSS 0.006764f
C11765 VDD.t1772 VSS 0.006764f
C11766 VDD.n1644 VSS 0.013528f
C11767 VDD.n1645 VSS 0.027737f
C11768 VDD.t8 VSS 0.018157f
C11769 VDD.t856 VSS 0.006764f
C11770 VDD.t10 VSS 0.006764f
C11771 VDD.n1646 VSS 0.014917f
C11772 VDD.t14 VSS 0.006764f
C11773 VDD.t844 VSS 0.006764f
C11774 VDD.n1647 VSS 0.014917f
C11775 VDD.t12 VSS 0.018157f
C11776 VDD.n1648 VSS 0.056289f
C11777 VDD.n1649 VSS 0.0563f
C11778 VDD.n1650 VSS 0.033732f
C11779 VDD.t609 VSS 0.006764f
C11780 VDD.t908 VSS 0.006764f
C11781 VDD.n1651 VSS 0.022549f
C11782 VDD.t1908 VSS 0.006764f
C11783 VDD.t1721 VSS 0.006764f
C11784 VDD.n1652 VSS 0.022549f
C11785 VDD.t607 VSS 0.025643f
C11786 VDD.n1653 VSS 0.104443f
C11787 VDD.t1719 VSS 0.018316f
C11788 VDD.n1654 VSS 0.097077f
C11789 VDD.n1655 VSS 0.07211f
C11790 VDD.n1656 VSS 0.037558f
C11791 VDD.n1657 VSS 0.015175f
C11792 VDD.t1774 VSS 0.01979f
C11793 VDD.t1711 VSS 0.01669f
C11794 VDD.n1658 VSS 0.049398f
C11795 VDD.n1659 VSS 0.018755f
C11796 VDD.n1660 VSS 0.102565f
C11797 VDD.t1756 VSS 0.138882f
C11798 VDD.t1726 VSS 0.363892f
C11799 VDD.t7 VSS 0.214331f
C11800 VDD.t9 VSS 0.136969f
C11801 VDD.t855 VSS 0.136969f
C11802 VDD.t843 VSS 0.136969f
C11803 VDD.t13 VSS 0.136969f
C11804 VDD.t11 VSS 0.141408f
C11805 VDD.t1718 VSS 0.214331f
C11806 VDD.t1720 VSS 0.136969f
C11807 VDD.t1907 VSS 0.136969f
C11808 VDD.t907 VSS 0.136969f
C11809 VDD.t608 VSS 0.136969f
C11810 VDD.t606 VSS 0.141408f
C11811 VDD.n1661 VSS 0.356736f
C11812 VDD.t806 VSS 0.408943f
C11813 VDD.t424 VSS 0.219141f
C11814 VDD.n1662 VSS 0.189733f
C11815 VDD.n1663 VSS -0.002571f
C11816 VDD.n1664 VSS 0.072393f
C11817 VDD.n1665 VSS 0.037945f
C11818 VDD.n1666 VSS 0.006361f
C11819 VDD.n1667 VSS 0.102565f
C11820 VDD.t1739 VSS 0.138882f
C11821 VDD.t1714 VSS 0.363892f
C11822 VDD.t1554 VSS 0.214331f
C11823 VDD.t1556 VSS 0.136969f
C11824 VDD.t177 VSS 0.136969f
C11825 VDD.t179 VSS 0.136969f
C11826 VDD.t2175 VSS 0.136969f
C11827 VDD.t2173 VSS 0.141408f
C11828 VDD.t1716 VSS 0.214331f
C11829 VDD.t1732 VSS 0.136969f
C11830 VDD.t1797 VSS 0.136969f
C11831 VDD.t1787 VSS 0.136969f
C11832 VDD.t345 VSS 0.136969f
C11833 VDD.t343 VSS 0.141408f
C11834 VDD.n1668 VSS 0.356736f
C11835 VDD.t410 VSS 0.408943f
C11836 VDD.t348 VSS 0.219141f
C11837 VDD.n1669 VSS 0.189733f
C11838 VDD.n1670 VSS -0.002571f
C11839 VDD.n1671 VSS 0.155963f
C11840 VDD.n1672 VSS 0.129222f
C11841 VDD.n1673 VSS 0.014817f
C11842 VDD.n1674 VSS 0.012937f
C11843 VDD.n1675 VSS 0.074505f
C11844 VDD.t497 VSS 0.066917f
C11845 VDD.n1676 VSS 0.071746f
C11846 VDD.n1677 VSS 0.054844f
C11847 VDD.n1678 VSS 0.01234f
C11848 VDD.n1679 VSS 0.007064f
C11849 VDD.n1680 VSS 0.114922f
C11850 VDD.n1681 VSS 0.194354f
C11851 VDD.n1682 VSS 0.028935f
C11852 VDD.n1683 VSS -0.002692f
C11853 VDD.n1684 VSS 0.270952f
C11854 VDD.t998 VSS 0.36819f
C11855 VDD.t996 VSS 0.264656f
C11856 VDD.t994 VSS 0.406173f
C11857 VDD.n1685 VSS 0.372359f
C11858 VDD.n1686 VSS 0.028538f
C11859 VDD.n1687 VSS 0.033316f
C11860 VDD.n1688 VSS -0.002692f
C11861 VDD.n1689 VSS 0.270952f
C11862 VDD.t1413 VSS 0.36819f
C11863 VDD.t1411 VSS 0.264656f
C11864 VDD.t1409 VSS 0.502356f
C11865 VDD.t1277 VSS 0.502356f
C11866 VDD.t1275 VSS 0.264656f
C11867 VDD.t1273 VSS 0.178275f
C11868 VDD.n1690 VSS 0.270952f
C11869 VDD.n1691 VSS -0.002692f
.ends

