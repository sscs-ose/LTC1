magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -4385 -1349 4385 1349
<< metal3 >>
rect -3385 344 3385 349
rect -3385 316 -3380 344
rect -3352 316 -3314 344
rect -3286 316 -3248 344
rect -3220 316 -3182 344
rect -3154 316 -3116 344
rect -3088 316 -3050 344
rect -3022 316 -2984 344
rect -2956 316 -2918 344
rect -2890 316 -2852 344
rect -2824 316 -2786 344
rect -2758 316 -2720 344
rect -2692 316 -2654 344
rect -2626 316 -2588 344
rect -2560 316 -2522 344
rect -2494 316 -2456 344
rect -2428 316 -2390 344
rect -2362 316 -2324 344
rect -2296 316 -2258 344
rect -2230 316 -2192 344
rect -2164 316 -2126 344
rect -2098 316 -2060 344
rect -2032 316 -1994 344
rect -1966 316 -1928 344
rect -1900 316 -1862 344
rect -1834 316 -1796 344
rect -1768 316 -1730 344
rect -1702 316 -1664 344
rect -1636 316 -1598 344
rect -1570 316 -1532 344
rect -1504 316 -1466 344
rect -1438 316 -1400 344
rect -1372 316 -1334 344
rect -1306 316 -1268 344
rect -1240 316 -1202 344
rect -1174 316 -1136 344
rect -1108 316 -1070 344
rect -1042 316 -1004 344
rect -976 316 -938 344
rect -910 316 -872 344
rect -844 316 -806 344
rect -778 316 -740 344
rect -712 316 -674 344
rect -646 316 -608 344
rect -580 316 -542 344
rect -514 316 -476 344
rect -448 316 -410 344
rect -382 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 382 344
rect 410 316 448 344
rect 476 316 514 344
rect 542 316 580 344
rect 608 316 646 344
rect 674 316 712 344
rect 740 316 778 344
rect 806 316 844 344
rect 872 316 910 344
rect 938 316 976 344
rect 1004 316 1042 344
rect 1070 316 1108 344
rect 1136 316 1174 344
rect 1202 316 1240 344
rect 1268 316 1306 344
rect 1334 316 1372 344
rect 1400 316 1438 344
rect 1466 316 1504 344
rect 1532 316 1570 344
rect 1598 316 1636 344
rect 1664 316 1702 344
rect 1730 316 1768 344
rect 1796 316 1834 344
rect 1862 316 1900 344
rect 1928 316 1966 344
rect 1994 316 2032 344
rect 2060 316 2098 344
rect 2126 316 2164 344
rect 2192 316 2230 344
rect 2258 316 2296 344
rect 2324 316 2362 344
rect 2390 316 2428 344
rect 2456 316 2494 344
rect 2522 316 2560 344
rect 2588 316 2626 344
rect 2654 316 2692 344
rect 2720 316 2758 344
rect 2786 316 2824 344
rect 2852 316 2890 344
rect 2918 316 2956 344
rect 2984 316 3022 344
rect 3050 316 3088 344
rect 3116 316 3154 344
rect 3182 316 3220 344
rect 3248 316 3286 344
rect 3314 316 3352 344
rect 3380 316 3385 344
rect -3385 278 3385 316
rect -3385 250 -3380 278
rect -3352 250 -3314 278
rect -3286 250 -3248 278
rect -3220 250 -3182 278
rect -3154 250 -3116 278
rect -3088 250 -3050 278
rect -3022 250 -2984 278
rect -2956 250 -2918 278
rect -2890 250 -2852 278
rect -2824 250 -2786 278
rect -2758 250 -2720 278
rect -2692 250 -2654 278
rect -2626 250 -2588 278
rect -2560 250 -2522 278
rect -2494 250 -2456 278
rect -2428 250 -2390 278
rect -2362 250 -2324 278
rect -2296 250 -2258 278
rect -2230 250 -2192 278
rect -2164 250 -2126 278
rect -2098 250 -2060 278
rect -2032 250 -1994 278
rect -1966 250 -1928 278
rect -1900 250 -1862 278
rect -1834 250 -1796 278
rect -1768 250 -1730 278
rect -1702 250 -1664 278
rect -1636 250 -1598 278
rect -1570 250 -1532 278
rect -1504 250 -1466 278
rect -1438 250 -1400 278
rect -1372 250 -1334 278
rect -1306 250 -1268 278
rect -1240 250 -1202 278
rect -1174 250 -1136 278
rect -1108 250 -1070 278
rect -1042 250 -1004 278
rect -976 250 -938 278
rect -910 250 -872 278
rect -844 250 -806 278
rect -778 250 -740 278
rect -712 250 -674 278
rect -646 250 -608 278
rect -580 250 -542 278
rect -514 250 -476 278
rect -448 250 -410 278
rect -382 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 382 278
rect 410 250 448 278
rect 476 250 514 278
rect 542 250 580 278
rect 608 250 646 278
rect 674 250 712 278
rect 740 250 778 278
rect 806 250 844 278
rect 872 250 910 278
rect 938 250 976 278
rect 1004 250 1042 278
rect 1070 250 1108 278
rect 1136 250 1174 278
rect 1202 250 1240 278
rect 1268 250 1306 278
rect 1334 250 1372 278
rect 1400 250 1438 278
rect 1466 250 1504 278
rect 1532 250 1570 278
rect 1598 250 1636 278
rect 1664 250 1702 278
rect 1730 250 1768 278
rect 1796 250 1834 278
rect 1862 250 1900 278
rect 1928 250 1966 278
rect 1994 250 2032 278
rect 2060 250 2098 278
rect 2126 250 2164 278
rect 2192 250 2230 278
rect 2258 250 2296 278
rect 2324 250 2362 278
rect 2390 250 2428 278
rect 2456 250 2494 278
rect 2522 250 2560 278
rect 2588 250 2626 278
rect 2654 250 2692 278
rect 2720 250 2758 278
rect 2786 250 2824 278
rect 2852 250 2890 278
rect 2918 250 2956 278
rect 2984 250 3022 278
rect 3050 250 3088 278
rect 3116 250 3154 278
rect 3182 250 3220 278
rect 3248 250 3286 278
rect 3314 250 3352 278
rect 3380 250 3385 278
rect -3385 212 3385 250
rect -3385 184 -3380 212
rect -3352 184 -3314 212
rect -3286 184 -3248 212
rect -3220 184 -3182 212
rect -3154 184 -3116 212
rect -3088 184 -3050 212
rect -3022 184 -2984 212
rect -2956 184 -2918 212
rect -2890 184 -2852 212
rect -2824 184 -2786 212
rect -2758 184 -2720 212
rect -2692 184 -2654 212
rect -2626 184 -2588 212
rect -2560 184 -2522 212
rect -2494 184 -2456 212
rect -2428 184 -2390 212
rect -2362 184 -2324 212
rect -2296 184 -2258 212
rect -2230 184 -2192 212
rect -2164 184 -2126 212
rect -2098 184 -2060 212
rect -2032 184 -1994 212
rect -1966 184 -1928 212
rect -1900 184 -1862 212
rect -1834 184 -1796 212
rect -1768 184 -1730 212
rect -1702 184 -1664 212
rect -1636 184 -1598 212
rect -1570 184 -1532 212
rect -1504 184 -1466 212
rect -1438 184 -1400 212
rect -1372 184 -1334 212
rect -1306 184 -1268 212
rect -1240 184 -1202 212
rect -1174 184 -1136 212
rect -1108 184 -1070 212
rect -1042 184 -1004 212
rect -976 184 -938 212
rect -910 184 -872 212
rect -844 184 -806 212
rect -778 184 -740 212
rect -712 184 -674 212
rect -646 184 -608 212
rect -580 184 -542 212
rect -514 184 -476 212
rect -448 184 -410 212
rect -382 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 382 212
rect 410 184 448 212
rect 476 184 514 212
rect 542 184 580 212
rect 608 184 646 212
rect 674 184 712 212
rect 740 184 778 212
rect 806 184 844 212
rect 872 184 910 212
rect 938 184 976 212
rect 1004 184 1042 212
rect 1070 184 1108 212
rect 1136 184 1174 212
rect 1202 184 1240 212
rect 1268 184 1306 212
rect 1334 184 1372 212
rect 1400 184 1438 212
rect 1466 184 1504 212
rect 1532 184 1570 212
rect 1598 184 1636 212
rect 1664 184 1702 212
rect 1730 184 1768 212
rect 1796 184 1834 212
rect 1862 184 1900 212
rect 1928 184 1966 212
rect 1994 184 2032 212
rect 2060 184 2098 212
rect 2126 184 2164 212
rect 2192 184 2230 212
rect 2258 184 2296 212
rect 2324 184 2362 212
rect 2390 184 2428 212
rect 2456 184 2494 212
rect 2522 184 2560 212
rect 2588 184 2626 212
rect 2654 184 2692 212
rect 2720 184 2758 212
rect 2786 184 2824 212
rect 2852 184 2890 212
rect 2918 184 2956 212
rect 2984 184 3022 212
rect 3050 184 3088 212
rect 3116 184 3154 212
rect 3182 184 3220 212
rect 3248 184 3286 212
rect 3314 184 3352 212
rect 3380 184 3385 212
rect -3385 146 3385 184
rect -3385 118 -3380 146
rect -3352 118 -3314 146
rect -3286 118 -3248 146
rect -3220 118 -3182 146
rect -3154 118 -3116 146
rect -3088 118 -3050 146
rect -3022 118 -2984 146
rect -2956 118 -2918 146
rect -2890 118 -2852 146
rect -2824 118 -2786 146
rect -2758 118 -2720 146
rect -2692 118 -2654 146
rect -2626 118 -2588 146
rect -2560 118 -2522 146
rect -2494 118 -2456 146
rect -2428 118 -2390 146
rect -2362 118 -2324 146
rect -2296 118 -2258 146
rect -2230 118 -2192 146
rect -2164 118 -2126 146
rect -2098 118 -2060 146
rect -2032 118 -1994 146
rect -1966 118 -1928 146
rect -1900 118 -1862 146
rect -1834 118 -1796 146
rect -1768 118 -1730 146
rect -1702 118 -1664 146
rect -1636 118 -1598 146
rect -1570 118 -1532 146
rect -1504 118 -1466 146
rect -1438 118 -1400 146
rect -1372 118 -1334 146
rect -1306 118 -1268 146
rect -1240 118 -1202 146
rect -1174 118 -1136 146
rect -1108 118 -1070 146
rect -1042 118 -1004 146
rect -976 118 -938 146
rect -910 118 -872 146
rect -844 118 -806 146
rect -778 118 -740 146
rect -712 118 -674 146
rect -646 118 -608 146
rect -580 118 -542 146
rect -514 118 -476 146
rect -448 118 -410 146
rect -382 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 382 146
rect 410 118 448 146
rect 476 118 514 146
rect 542 118 580 146
rect 608 118 646 146
rect 674 118 712 146
rect 740 118 778 146
rect 806 118 844 146
rect 872 118 910 146
rect 938 118 976 146
rect 1004 118 1042 146
rect 1070 118 1108 146
rect 1136 118 1174 146
rect 1202 118 1240 146
rect 1268 118 1306 146
rect 1334 118 1372 146
rect 1400 118 1438 146
rect 1466 118 1504 146
rect 1532 118 1570 146
rect 1598 118 1636 146
rect 1664 118 1702 146
rect 1730 118 1768 146
rect 1796 118 1834 146
rect 1862 118 1900 146
rect 1928 118 1966 146
rect 1994 118 2032 146
rect 2060 118 2098 146
rect 2126 118 2164 146
rect 2192 118 2230 146
rect 2258 118 2296 146
rect 2324 118 2362 146
rect 2390 118 2428 146
rect 2456 118 2494 146
rect 2522 118 2560 146
rect 2588 118 2626 146
rect 2654 118 2692 146
rect 2720 118 2758 146
rect 2786 118 2824 146
rect 2852 118 2890 146
rect 2918 118 2956 146
rect 2984 118 3022 146
rect 3050 118 3088 146
rect 3116 118 3154 146
rect 3182 118 3220 146
rect 3248 118 3286 146
rect 3314 118 3352 146
rect 3380 118 3385 146
rect -3385 80 3385 118
rect -3385 52 -3380 80
rect -3352 52 -3314 80
rect -3286 52 -3248 80
rect -3220 52 -3182 80
rect -3154 52 -3116 80
rect -3088 52 -3050 80
rect -3022 52 -2984 80
rect -2956 52 -2918 80
rect -2890 52 -2852 80
rect -2824 52 -2786 80
rect -2758 52 -2720 80
rect -2692 52 -2654 80
rect -2626 52 -2588 80
rect -2560 52 -2522 80
rect -2494 52 -2456 80
rect -2428 52 -2390 80
rect -2362 52 -2324 80
rect -2296 52 -2258 80
rect -2230 52 -2192 80
rect -2164 52 -2126 80
rect -2098 52 -2060 80
rect -2032 52 -1994 80
rect -1966 52 -1928 80
rect -1900 52 -1862 80
rect -1834 52 -1796 80
rect -1768 52 -1730 80
rect -1702 52 -1664 80
rect -1636 52 -1598 80
rect -1570 52 -1532 80
rect -1504 52 -1466 80
rect -1438 52 -1400 80
rect -1372 52 -1334 80
rect -1306 52 -1268 80
rect -1240 52 -1202 80
rect -1174 52 -1136 80
rect -1108 52 -1070 80
rect -1042 52 -1004 80
rect -976 52 -938 80
rect -910 52 -872 80
rect -844 52 -806 80
rect -778 52 -740 80
rect -712 52 -674 80
rect -646 52 -608 80
rect -580 52 -542 80
rect -514 52 -476 80
rect -448 52 -410 80
rect -382 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 382 80
rect 410 52 448 80
rect 476 52 514 80
rect 542 52 580 80
rect 608 52 646 80
rect 674 52 712 80
rect 740 52 778 80
rect 806 52 844 80
rect 872 52 910 80
rect 938 52 976 80
rect 1004 52 1042 80
rect 1070 52 1108 80
rect 1136 52 1174 80
rect 1202 52 1240 80
rect 1268 52 1306 80
rect 1334 52 1372 80
rect 1400 52 1438 80
rect 1466 52 1504 80
rect 1532 52 1570 80
rect 1598 52 1636 80
rect 1664 52 1702 80
rect 1730 52 1768 80
rect 1796 52 1834 80
rect 1862 52 1900 80
rect 1928 52 1966 80
rect 1994 52 2032 80
rect 2060 52 2098 80
rect 2126 52 2164 80
rect 2192 52 2230 80
rect 2258 52 2296 80
rect 2324 52 2362 80
rect 2390 52 2428 80
rect 2456 52 2494 80
rect 2522 52 2560 80
rect 2588 52 2626 80
rect 2654 52 2692 80
rect 2720 52 2758 80
rect 2786 52 2824 80
rect 2852 52 2890 80
rect 2918 52 2956 80
rect 2984 52 3022 80
rect 3050 52 3088 80
rect 3116 52 3154 80
rect 3182 52 3220 80
rect 3248 52 3286 80
rect 3314 52 3352 80
rect 3380 52 3385 80
rect -3385 14 3385 52
rect -3385 -14 -3380 14
rect -3352 -14 -3314 14
rect -3286 -14 -3248 14
rect -3220 -14 -3182 14
rect -3154 -14 -3116 14
rect -3088 -14 -3050 14
rect -3022 -14 -2984 14
rect -2956 -14 -2918 14
rect -2890 -14 -2852 14
rect -2824 -14 -2786 14
rect -2758 -14 -2720 14
rect -2692 -14 -2654 14
rect -2626 -14 -2588 14
rect -2560 -14 -2522 14
rect -2494 -14 -2456 14
rect -2428 -14 -2390 14
rect -2362 -14 -2324 14
rect -2296 -14 -2258 14
rect -2230 -14 -2192 14
rect -2164 -14 -2126 14
rect -2098 -14 -2060 14
rect -2032 -14 -1994 14
rect -1966 -14 -1928 14
rect -1900 -14 -1862 14
rect -1834 -14 -1796 14
rect -1768 -14 -1730 14
rect -1702 -14 -1664 14
rect -1636 -14 -1598 14
rect -1570 -14 -1532 14
rect -1504 -14 -1466 14
rect -1438 -14 -1400 14
rect -1372 -14 -1334 14
rect -1306 -14 -1268 14
rect -1240 -14 -1202 14
rect -1174 -14 -1136 14
rect -1108 -14 -1070 14
rect -1042 -14 -1004 14
rect -976 -14 -938 14
rect -910 -14 -872 14
rect -844 -14 -806 14
rect -778 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 382 14
rect 410 -14 448 14
rect 476 -14 514 14
rect 542 -14 580 14
rect 608 -14 646 14
rect 674 -14 712 14
rect 740 -14 778 14
rect 806 -14 844 14
rect 872 -14 910 14
rect 938 -14 976 14
rect 1004 -14 1042 14
rect 1070 -14 1108 14
rect 1136 -14 1174 14
rect 1202 -14 1240 14
rect 1268 -14 1306 14
rect 1334 -14 1372 14
rect 1400 -14 1438 14
rect 1466 -14 1504 14
rect 1532 -14 1570 14
rect 1598 -14 1636 14
rect 1664 -14 1702 14
rect 1730 -14 1768 14
rect 1796 -14 1834 14
rect 1862 -14 1900 14
rect 1928 -14 1966 14
rect 1994 -14 2032 14
rect 2060 -14 2098 14
rect 2126 -14 2164 14
rect 2192 -14 2230 14
rect 2258 -14 2296 14
rect 2324 -14 2362 14
rect 2390 -14 2428 14
rect 2456 -14 2494 14
rect 2522 -14 2560 14
rect 2588 -14 2626 14
rect 2654 -14 2692 14
rect 2720 -14 2758 14
rect 2786 -14 2824 14
rect 2852 -14 2890 14
rect 2918 -14 2956 14
rect 2984 -14 3022 14
rect 3050 -14 3088 14
rect 3116 -14 3154 14
rect 3182 -14 3220 14
rect 3248 -14 3286 14
rect 3314 -14 3352 14
rect 3380 -14 3385 14
rect -3385 -52 3385 -14
rect -3385 -80 -3380 -52
rect -3352 -80 -3314 -52
rect -3286 -80 -3248 -52
rect -3220 -80 -3182 -52
rect -3154 -80 -3116 -52
rect -3088 -80 -3050 -52
rect -3022 -80 -2984 -52
rect -2956 -80 -2918 -52
rect -2890 -80 -2852 -52
rect -2824 -80 -2786 -52
rect -2758 -80 -2720 -52
rect -2692 -80 -2654 -52
rect -2626 -80 -2588 -52
rect -2560 -80 -2522 -52
rect -2494 -80 -2456 -52
rect -2428 -80 -2390 -52
rect -2362 -80 -2324 -52
rect -2296 -80 -2258 -52
rect -2230 -80 -2192 -52
rect -2164 -80 -2126 -52
rect -2098 -80 -2060 -52
rect -2032 -80 -1994 -52
rect -1966 -80 -1928 -52
rect -1900 -80 -1862 -52
rect -1834 -80 -1796 -52
rect -1768 -80 -1730 -52
rect -1702 -80 -1664 -52
rect -1636 -80 -1598 -52
rect -1570 -80 -1532 -52
rect -1504 -80 -1466 -52
rect -1438 -80 -1400 -52
rect -1372 -80 -1334 -52
rect -1306 -80 -1268 -52
rect -1240 -80 -1202 -52
rect -1174 -80 -1136 -52
rect -1108 -80 -1070 -52
rect -1042 -80 -1004 -52
rect -976 -80 -938 -52
rect -910 -80 -872 -52
rect -844 -80 -806 -52
rect -778 -80 -740 -52
rect -712 -80 -674 -52
rect -646 -80 -608 -52
rect -580 -80 -542 -52
rect -514 -80 -476 -52
rect -448 -80 -410 -52
rect -382 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 382 -52
rect 410 -80 448 -52
rect 476 -80 514 -52
rect 542 -80 580 -52
rect 608 -80 646 -52
rect 674 -80 712 -52
rect 740 -80 778 -52
rect 806 -80 844 -52
rect 872 -80 910 -52
rect 938 -80 976 -52
rect 1004 -80 1042 -52
rect 1070 -80 1108 -52
rect 1136 -80 1174 -52
rect 1202 -80 1240 -52
rect 1268 -80 1306 -52
rect 1334 -80 1372 -52
rect 1400 -80 1438 -52
rect 1466 -80 1504 -52
rect 1532 -80 1570 -52
rect 1598 -80 1636 -52
rect 1664 -80 1702 -52
rect 1730 -80 1768 -52
rect 1796 -80 1834 -52
rect 1862 -80 1900 -52
rect 1928 -80 1966 -52
rect 1994 -80 2032 -52
rect 2060 -80 2098 -52
rect 2126 -80 2164 -52
rect 2192 -80 2230 -52
rect 2258 -80 2296 -52
rect 2324 -80 2362 -52
rect 2390 -80 2428 -52
rect 2456 -80 2494 -52
rect 2522 -80 2560 -52
rect 2588 -80 2626 -52
rect 2654 -80 2692 -52
rect 2720 -80 2758 -52
rect 2786 -80 2824 -52
rect 2852 -80 2890 -52
rect 2918 -80 2956 -52
rect 2984 -80 3022 -52
rect 3050 -80 3088 -52
rect 3116 -80 3154 -52
rect 3182 -80 3220 -52
rect 3248 -80 3286 -52
rect 3314 -80 3352 -52
rect 3380 -80 3385 -52
rect -3385 -118 3385 -80
rect -3385 -146 -3380 -118
rect -3352 -146 -3314 -118
rect -3286 -146 -3248 -118
rect -3220 -146 -3182 -118
rect -3154 -146 -3116 -118
rect -3088 -146 -3050 -118
rect -3022 -146 -2984 -118
rect -2956 -146 -2918 -118
rect -2890 -146 -2852 -118
rect -2824 -146 -2786 -118
rect -2758 -146 -2720 -118
rect -2692 -146 -2654 -118
rect -2626 -146 -2588 -118
rect -2560 -146 -2522 -118
rect -2494 -146 -2456 -118
rect -2428 -146 -2390 -118
rect -2362 -146 -2324 -118
rect -2296 -146 -2258 -118
rect -2230 -146 -2192 -118
rect -2164 -146 -2126 -118
rect -2098 -146 -2060 -118
rect -2032 -146 -1994 -118
rect -1966 -146 -1928 -118
rect -1900 -146 -1862 -118
rect -1834 -146 -1796 -118
rect -1768 -146 -1730 -118
rect -1702 -146 -1664 -118
rect -1636 -146 -1598 -118
rect -1570 -146 -1532 -118
rect -1504 -146 -1466 -118
rect -1438 -146 -1400 -118
rect -1372 -146 -1334 -118
rect -1306 -146 -1268 -118
rect -1240 -146 -1202 -118
rect -1174 -146 -1136 -118
rect -1108 -146 -1070 -118
rect -1042 -146 -1004 -118
rect -976 -146 -938 -118
rect -910 -146 -872 -118
rect -844 -146 -806 -118
rect -778 -146 -740 -118
rect -712 -146 -674 -118
rect -646 -146 -608 -118
rect -580 -146 -542 -118
rect -514 -146 -476 -118
rect -448 -146 -410 -118
rect -382 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 382 -118
rect 410 -146 448 -118
rect 476 -146 514 -118
rect 542 -146 580 -118
rect 608 -146 646 -118
rect 674 -146 712 -118
rect 740 -146 778 -118
rect 806 -146 844 -118
rect 872 -146 910 -118
rect 938 -146 976 -118
rect 1004 -146 1042 -118
rect 1070 -146 1108 -118
rect 1136 -146 1174 -118
rect 1202 -146 1240 -118
rect 1268 -146 1306 -118
rect 1334 -146 1372 -118
rect 1400 -146 1438 -118
rect 1466 -146 1504 -118
rect 1532 -146 1570 -118
rect 1598 -146 1636 -118
rect 1664 -146 1702 -118
rect 1730 -146 1768 -118
rect 1796 -146 1834 -118
rect 1862 -146 1900 -118
rect 1928 -146 1966 -118
rect 1994 -146 2032 -118
rect 2060 -146 2098 -118
rect 2126 -146 2164 -118
rect 2192 -146 2230 -118
rect 2258 -146 2296 -118
rect 2324 -146 2362 -118
rect 2390 -146 2428 -118
rect 2456 -146 2494 -118
rect 2522 -146 2560 -118
rect 2588 -146 2626 -118
rect 2654 -146 2692 -118
rect 2720 -146 2758 -118
rect 2786 -146 2824 -118
rect 2852 -146 2890 -118
rect 2918 -146 2956 -118
rect 2984 -146 3022 -118
rect 3050 -146 3088 -118
rect 3116 -146 3154 -118
rect 3182 -146 3220 -118
rect 3248 -146 3286 -118
rect 3314 -146 3352 -118
rect 3380 -146 3385 -118
rect -3385 -184 3385 -146
rect -3385 -212 -3380 -184
rect -3352 -212 -3314 -184
rect -3286 -212 -3248 -184
rect -3220 -212 -3182 -184
rect -3154 -212 -3116 -184
rect -3088 -212 -3050 -184
rect -3022 -212 -2984 -184
rect -2956 -212 -2918 -184
rect -2890 -212 -2852 -184
rect -2824 -212 -2786 -184
rect -2758 -212 -2720 -184
rect -2692 -212 -2654 -184
rect -2626 -212 -2588 -184
rect -2560 -212 -2522 -184
rect -2494 -212 -2456 -184
rect -2428 -212 -2390 -184
rect -2362 -212 -2324 -184
rect -2296 -212 -2258 -184
rect -2230 -212 -2192 -184
rect -2164 -212 -2126 -184
rect -2098 -212 -2060 -184
rect -2032 -212 -1994 -184
rect -1966 -212 -1928 -184
rect -1900 -212 -1862 -184
rect -1834 -212 -1796 -184
rect -1768 -212 -1730 -184
rect -1702 -212 -1664 -184
rect -1636 -212 -1598 -184
rect -1570 -212 -1532 -184
rect -1504 -212 -1466 -184
rect -1438 -212 -1400 -184
rect -1372 -212 -1334 -184
rect -1306 -212 -1268 -184
rect -1240 -212 -1202 -184
rect -1174 -212 -1136 -184
rect -1108 -212 -1070 -184
rect -1042 -212 -1004 -184
rect -976 -212 -938 -184
rect -910 -212 -872 -184
rect -844 -212 -806 -184
rect -778 -212 -740 -184
rect -712 -212 -674 -184
rect -646 -212 -608 -184
rect -580 -212 -542 -184
rect -514 -212 -476 -184
rect -448 -212 -410 -184
rect -382 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 382 -184
rect 410 -212 448 -184
rect 476 -212 514 -184
rect 542 -212 580 -184
rect 608 -212 646 -184
rect 674 -212 712 -184
rect 740 -212 778 -184
rect 806 -212 844 -184
rect 872 -212 910 -184
rect 938 -212 976 -184
rect 1004 -212 1042 -184
rect 1070 -212 1108 -184
rect 1136 -212 1174 -184
rect 1202 -212 1240 -184
rect 1268 -212 1306 -184
rect 1334 -212 1372 -184
rect 1400 -212 1438 -184
rect 1466 -212 1504 -184
rect 1532 -212 1570 -184
rect 1598 -212 1636 -184
rect 1664 -212 1702 -184
rect 1730 -212 1768 -184
rect 1796 -212 1834 -184
rect 1862 -212 1900 -184
rect 1928 -212 1966 -184
rect 1994 -212 2032 -184
rect 2060 -212 2098 -184
rect 2126 -212 2164 -184
rect 2192 -212 2230 -184
rect 2258 -212 2296 -184
rect 2324 -212 2362 -184
rect 2390 -212 2428 -184
rect 2456 -212 2494 -184
rect 2522 -212 2560 -184
rect 2588 -212 2626 -184
rect 2654 -212 2692 -184
rect 2720 -212 2758 -184
rect 2786 -212 2824 -184
rect 2852 -212 2890 -184
rect 2918 -212 2956 -184
rect 2984 -212 3022 -184
rect 3050 -212 3088 -184
rect 3116 -212 3154 -184
rect 3182 -212 3220 -184
rect 3248 -212 3286 -184
rect 3314 -212 3352 -184
rect 3380 -212 3385 -184
rect -3385 -250 3385 -212
rect -3385 -278 -3380 -250
rect -3352 -278 -3314 -250
rect -3286 -278 -3248 -250
rect -3220 -278 -3182 -250
rect -3154 -278 -3116 -250
rect -3088 -278 -3050 -250
rect -3022 -278 -2984 -250
rect -2956 -278 -2918 -250
rect -2890 -278 -2852 -250
rect -2824 -278 -2786 -250
rect -2758 -278 -2720 -250
rect -2692 -278 -2654 -250
rect -2626 -278 -2588 -250
rect -2560 -278 -2522 -250
rect -2494 -278 -2456 -250
rect -2428 -278 -2390 -250
rect -2362 -278 -2324 -250
rect -2296 -278 -2258 -250
rect -2230 -278 -2192 -250
rect -2164 -278 -2126 -250
rect -2098 -278 -2060 -250
rect -2032 -278 -1994 -250
rect -1966 -278 -1928 -250
rect -1900 -278 -1862 -250
rect -1834 -278 -1796 -250
rect -1768 -278 -1730 -250
rect -1702 -278 -1664 -250
rect -1636 -278 -1598 -250
rect -1570 -278 -1532 -250
rect -1504 -278 -1466 -250
rect -1438 -278 -1400 -250
rect -1372 -278 -1334 -250
rect -1306 -278 -1268 -250
rect -1240 -278 -1202 -250
rect -1174 -278 -1136 -250
rect -1108 -278 -1070 -250
rect -1042 -278 -1004 -250
rect -976 -278 -938 -250
rect -910 -278 -872 -250
rect -844 -278 -806 -250
rect -778 -278 -740 -250
rect -712 -278 -674 -250
rect -646 -278 -608 -250
rect -580 -278 -542 -250
rect -514 -278 -476 -250
rect -448 -278 -410 -250
rect -382 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 382 -250
rect 410 -278 448 -250
rect 476 -278 514 -250
rect 542 -278 580 -250
rect 608 -278 646 -250
rect 674 -278 712 -250
rect 740 -278 778 -250
rect 806 -278 844 -250
rect 872 -278 910 -250
rect 938 -278 976 -250
rect 1004 -278 1042 -250
rect 1070 -278 1108 -250
rect 1136 -278 1174 -250
rect 1202 -278 1240 -250
rect 1268 -278 1306 -250
rect 1334 -278 1372 -250
rect 1400 -278 1438 -250
rect 1466 -278 1504 -250
rect 1532 -278 1570 -250
rect 1598 -278 1636 -250
rect 1664 -278 1702 -250
rect 1730 -278 1768 -250
rect 1796 -278 1834 -250
rect 1862 -278 1900 -250
rect 1928 -278 1966 -250
rect 1994 -278 2032 -250
rect 2060 -278 2098 -250
rect 2126 -278 2164 -250
rect 2192 -278 2230 -250
rect 2258 -278 2296 -250
rect 2324 -278 2362 -250
rect 2390 -278 2428 -250
rect 2456 -278 2494 -250
rect 2522 -278 2560 -250
rect 2588 -278 2626 -250
rect 2654 -278 2692 -250
rect 2720 -278 2758 -250
rect 2786 -278 2824 -250
rect 2852 -278 2890 -250
rect 2918 -278 2956 -250
rect 2984 -278 3022 -250
rect 3050 -278 3088 -250
rect 3116 -278 3154 -250
rect 3182 -278 3220 -250
rect 3248 -278 3286 -250
rect 3314 -278 3352 -250
rect 3380 -278 3385 -250
rect -3385 -316 3385 -278
rect -3385 -344 -3380 -316
rect -3352 -344 -3314 -316
rect -3286 -344 -3248 -316
rect -3220 -344 -3182 -316
rect -3154 -344 -3116 -316
rect -3088 -344 -3050 -316
rect -3022 -344 -2984 -316
rect -2956 -344 -2918 -316
rect -2890 -344 -2852 -316
rect -2824 -344 -2786 -316
rect -2758 -344 -2720 -316
rect -2692 -344 -2654 -316
rect -2626 -344 -2588 -316
rect -2560 -344 -2522 -316
rect -2494 -344 -2456 -316
rect -2428 -344 -2390 -316
rect -2362 -344 -2324 -316
rect -2296 -344 -2258 -316
rect -2230 -344 -2192 -316
rect -2164 -344 -2126 -316
rect -2098 -344 -2060 -316
rect -2032 -344 -1994 -316
rect -1966 -344 -1928 -316
rect -1900 -344 -1862 -316
rect -1834 -344 -1796 -316
rect -1768 -344 -1730 -316
rect -1702 -344 -1664 -316
rect -1636 -344 -1598 -316
rect -1570 -344 -1532 -316
rect -1504 -344 -1466 -316
rect -1438 -344 -1400 -316
rect -1372 -344 -1334 -316
rect -1306 -344 -1268 -316
rect -1240 -344 -1202 -316
rect -1174 -344 -1136 -316
rect -1108 -344 -1070 -316
rect -1042 -344 -1004 -316
rect -976 -344 -938 -316
rect -910 -344 -872 -316
rect -844 -344 -806 -316
rect -778 -344 -740 -316
rect -712 -344 -674 -316
rect -646 -344 -608 -316
rect -580 -344 -542 -316
rect -514 -344 -476 -316
rect -448 -344 -410 -316
rect -382 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 382 -316
rect 410 -344 448 -316
rect 476 -344 514 -316
rect 542 -344 580 -316
rect 608 -344 646 -316
rect 674 -344 712 -316
rect 740 -344 778 -316
rect 806 -344 844 -316
rect 872 -344 910 -316
rect 938 -344 976 -316
rect 1004 -344 1042 -316
rect 1070 -344 1108 -316
rect 1136 -344 1174 -316
rect 1202 -344 1240 -316
rect 1268 -344 1306 -316
rect 1334 -344 1372 -316
rect 1400 -344 1438 -316
rect 1466 -344 1504 -316
rect 1532 -344 1570 -316
rect 1598 -344 1636 -316
rect 1664 -344 1702 -316
rect 1730 -344 1768 -316
rect 1796 -344 1834 -316
rect 1862 -344 1900 -316
rect 1928 -344 1966 -316
rect 1994 -344 2032 -316
rect 2060 -344 2098 -316
rect 2126 -344 2164 -316
rect 2192 -344 2230 -316
rect 2258 -344 2296 -316
rect 2324 -344 2362 -316
rect 2390 -344 2428 -316
rect 2456 -344 2494 -316
rect 2522 -344 2560 -316
rect 2588 -344 2626 -316
rect 2654 -344 2692 -316
rect 2720 -344 2758 -316
rect 2786 -344 2824 -316
rect 2852 -344 2890 -316
rect 2918 -344 2956 -316
rect 2984 -344 3022 -316
rect 3050 -344 3088 -316
rect 3116 -344 3154 -316
rect 3182 -344 3220 -316
rect 3248 -344 3286 -316
rect 3314 -344 3352 -316
rect 3380 -344 3385 -316
rect -3385 -349 3385 -344
<< via3 >>
rect -3380 316 -3352 344
rect -3314 316 -3286 344
rect -3248 316 -3220 344
rect -3182 316 -3154 344
rect -3116 316 -3088 344
rect -3050 316 -3022 344
rect -2984 316 -2956 344
rect -2918 316 -2890 344
rect -2852 316 -2824 344
rect -2786 316 -2758 344
rect -2720 316 -2692 344
rect -2654 316 -2626 344
rect -2588 316 -2560 344
rect -2522 316 -2494 344
rect -2456 316 -2428 344
rect -2390 316 -2362 344
rect -2324 316 -2296 344
rect -2258 316 -2230 344
rect -2192 316 -2164 344
rect -2126 316 -2098 344
rect -2060 316 -2032 344
rect -1994 316 -1966 344
rect -1928 316 -1900 344
rect -1862 316 -1834 344
rect -1796 316 -1768 344
rect -1730 316 -1702 344
rect -1664 316 -1636 344
rect -1598 316 -1570 344
rect -1532 316 -1504 344
rect -1466 316 -1438 344
rect -1400 316 -1372 344
rect -1334 316 -1306 344
rect -1268 316 -1240 344
rect -1202 316 -1174 344
rect -1136 316 -1108 344
rect -1070 316 -1042 344
rect -1004 316 -976 344
rect -938 316 -910 344
rect -872 316 -844 344
rect -806 316 -778 344
rect -740 316 -712 344
rect -674 316 -646 344
rect -608 316 -580 344
rect -542 316 -514 344
rect -476 316 -448 344
rect -410 316 -382 344
rect -344 316 -316 344
rect -278 316 -250 344
rect -212 316 -184 344
rect -146 316 -118 344
rect -80 316 -52 344
rect -14 316 14 344
rect 52 316 80 344
rect 118 316 146 344
rect 184 316 212 344
rect 250 316 278 344
rect 316 316 344 344
rect 382 316 410 344
rect 448 316 476 344
rect 514 316 542 344
rect 580 316 608 344
rect 646 316 674 344
rect 712 316 740 344
rect 778 316 806 344
rect 844 316 872 344
rect 910 316 938 344
rect 976 316 1004 344
rect 1042 316 1070 344
rect 1108 316 1136 344
rect 1174 316 1202 344
rect 1240 316 1268 344
rect 1306 316 1334 344
rect 1372 316 1400 344
rect 1438 316 1466 344
rect 1504 316 1532 344
rect 1570 316 1598 344
rect 1636 316 1664 344
rect 1702 316 1730 344
rect 1768 316 1796 344
rect 1834 316 1862 344
rect 1900 316 1928 344
rect 1966 316 1994 344
rect 2032 316 2060 344
rect 2098 316 2126 344
rect 2164 316 2192 344
rect 2230 316 2258 344
rect 2296 316 2324 344
rect 2362 316 2390 344
rect 2428 316 2456 344
rect 2494 316 2522 344
rect 2560 316 2588 344
rect 2626 316 2654 344
rect 2692 316 2720 344
rect 2758 316 2786 344
rect 2824 316 2852 344
rect 2890 316 2918 344
rect 2956 316 2984 344
rect 3022 316 3050 344
rect 3088 316 3116 344
rect 3154 316 3182 344
rect 3220 316 3248 344
rect 3286 316 3314 344
rect 3352 316 3380 344
rect -3380 250 -3352 278
rect -3314 250 -3286 278
rect -3248 250 -3220 278
rect -3182 250 -3154 278
rect -3116 250 -3088 278
rect -3050 250 -3022 278
rect -2984 250 -2956 278
rect -2918 250 -2890 278
rect -2852 250 -2824 278
rect -2786 250 -2758 278
rect -2720 250 -2692 278
rect -2654 250 -2626 278
rect -2588 250 -2560 278
rect -2522 250 -2494 278
rect -2456 250 -2428 278
rect -2390 250 -2362 278
rect -2324 250 -2296 278
rect -2258 250 -2230 278
rect -2192 250 -2164 278
rect -2126 250 -2098 278
rect -2060 250 -2032 278
rect -1994 250 -1966 278
rect -1928 250 -1900 278
rect -1862 250 -1834 278
rect -1796 250 -1768 278
rect -1730 250 -1702 278
rect -1664 250 -1636 278
rect -1598 250 -1570 278
rect -1532 250 -1504 278
rect -1466 250 -1438 278
rect -1400 250 -1372 278
rect -1334 250 -1306 278
rect -1268 250 -1240 278
rect -1202 250 -1174 278
rect -1136 250 -1108 278
rect -1070 250 -1042 278
rect -1004 250 -976 278
rect -938 250 -910 278
rect -872 250 -844 278
rect -806 250 -778 278
rect -740 250 -712 278
rect -674 250 -646 278
rect -608 250 -580 278
rect -542 250 -514 278
rect -476 250 -448 278
rect -410 250 -382 278
rect -344 250 -316 278
rect -278 250 -250 278
rect -212 250 -184 278
rect -146 250 -118 278
rect -80 250 -52 278
rect -14 250 14 278
rect 52 250 80 278
rect 118 250 146 278
rect 184 250 212 278
rect 250 250 278 278
rect 316 250 344 278
rect 382 250 410 278
rect 448 250 476 278
rect 514 250 542 278
rect 580 250 608 278
rect 646 250 674 278
rect 712 250 740 278
rect 778 250 806 278
rect 844 250 872 278
rect 910 250 938 278
rect 976 250 1004 278
rect 1042 250 1070 278
rect 1108 250 1136 278
rect 1174 250 1202 278
rect 1240 250 1268 278
rect 1306 250 1334 278
rect 1372 250 1400 278
rect 1438 250 1466 278
rect 1504 250 1532 278
rect 1570 250 1598 278
rect 1636 250 1664 278
rect 1702 250 1730 278
rect 1768 250 1796 278
rect 1834 250 1862 278
rect 1900 250 1928 278
rect 1966 250 1994 278
rect 2032 250 2060 278
rect 2098 250 2126 278
rect 2164 250 2192 278
rect 2230 250 2258 278
rect 2296 250 2324 278
rect 2362 250 2390 278
rect 2428 250 2456 278
rect 2494 250 2522 278
rect 2560 250 2588 278
rect 2626 250 2654 278
rect 2692 250 2720 278
rect 2758 250 2786 278
rect 2824 250 2852 278
rect 2890 250 2918 278
rect 2956 250 2984 278
rect 3022 250 3050 278
rect 3088 250 3116 278
rect 3154 250 3182 278
rect 3220 250 3248 278
rect 3286 250 3314 278
rect 3352 250 3380 278
rect -3380 184 -3352 212
rect -3314 184 -3286 212
rect -3248 184 -3220 212
rect -3182 184 -3154 212
rect -3116 184 -3088 212
rect -3050 184 -3022 212
rect -2984 184 -2956 212
rect -2918 184 -2890 212
rect -2852 184 -2824 212
rect -2786 184 -2758 212
rect -2720 184 -2692 212
rect -2654 184 -2626 212
rect -2588 184 -2560 212
rect -2522 184 -2494 212
rect -2456 184 -2428 212
rect -2390 184 -2362 212
rect -2324 184 -2296 212
rect -2258 184 -2230 212
rect -2192 184 -2164 212
rect -2126 184 -2098 212
rect -2060 184 -2032 212
rect -1994 184 -1966 212
rect -1928 184 -1900 212
rect -1862 184 -1834 212
rect -1796 184 -1768 212
rect -1730 184 -1702 212
rect -1664 184 -1636 212
rect -1598 184 -1570 212
rect -1532 184 -1504 212
rect -1466 184 -1438 212
rect -1400 184 -1372 212
rect -1334 184 -1306 212
rect -1268 184 -1240 212
rect -1202 184 -1174 212
rect -1136 184 -1108 212
rect -1070 184 -1042 212
rect -1004 184 -976 212
rect -938 184 -910 212
rect -872 184 -844 212
rect -806 184 -778 212
rect -740 184 -712 212
rect -674 184 -646 212
rect -608 184 -580 212
rect -542 184 -514 212
rect -476 184 -448 212
rect -410 184 -382 212
rect -344 184 -316 212
rect -278 184 -250 212
rect -212 184 -184 212
rect -146 184 -118 212
rect -80 184 -52 212
rect -14 184 14 212
rect 52 184 80 212
rect 118 184 146 212
rect 184 184 212 212
rect 250 184 278 212
rect 316 184 344 212
rect 382 184 410 212
rect 448 184 476 212
rect 514 184 542 212
rect 580 184 608 212
rect 646 184 674 212
rect 712 184 740 212
rect 778 184 806 212
rect 844 184 872 212
rect 910 184 938 212
rect 976 184 1004 212
rect 1042 184 1070 212
rect 1108 184 1136 212
rect 1174 184 1202 212
rect 1240 184 1268 212
rect 1306 184 1334 212
rect 1372 184 1400 212
rect 1438 184 1466 212
rect 1504 184 1532 212
rect 1570 184 1598 212
rect 1636 184 1664 212
rect 1702 184 1730 212
rect 1768 184 1796 212
rect 1834 184 1862 212
rect 1900 184 1928 212
rect 1966 184 1994 212
rect 2032 184 2060 212
rect 2098 184 2126 212
rect 2164 184 2192 212
rect 2230 184 2258 212
rect 2296 184 2324 212
rect 2362 184 2390 212
rect 2428 184 2456 212
rect 2494 184 2522 212
rect 2560 184 2588 212
rect 2626 184 2654 212
rect 2692 184 2720 212
rect 2758 184 2786 212
rect 2824 184 2852 212
rect 2890 184 2918 212
rect 2956 184 2984 212
rect 3022 184 3050 212
rect 3088 184 3116 212
rect 3154 184 3182 212
rect 3220 184 3248 212
rect 3286 184 3314 212
rect 3352 184 3380 212
rect -3380 118 -3352 146
rect -3314 118 -3286 146
rect -3248 118 -3220 146
rect -3182 118 -3154 146
rect -3116 118 -3088 146
rect -3050 118 -3022 146
rect -2984 118 -2956 146
rect -2918 118 -2890 146
rect -2852 118 -2824 146
rect -2786 118 -2758 146
rect -2720 118 -2692 146
rect -2654 118 -2626 146
rect -2588 118 -2560 146
rect -2522 118 -2494 146
rect -2456 118 -2428 146
rect -2390 118 -2362 146
rect -2324 118 -2296 146
rect -2258 118 -2230 146
rect -2192 118 -2164 146
rect -2126 118 -2098 146
rect -2060 118 -2032 146
rect -1994 118 -1966 146
rect -1928 118 -1900 146
rect -1862 118 -1834 146
rect -1796 118 -1768 146
rect -1730 118 -1702 146
rect -1664 118 -1636 146
rect -1598 118 -1570 146
rect -1532 118 -1504 146
rect -1466 118 -1438 146
rect -1400 118 -1372 146
rect -1334 118 -1306 146
rect -1268 118 -1240 146
rect -1202 118 -1174 146
rect -1136 118 -1108 146
rect -1070 118 -1042 146
rect -1004 118 -976 146
rect -938 118 -910 146
rect -872 118 -844 146
rect -806 118 -778 146
rect -740 118 -712 146
rect -674 118 -646 146
rect -608 118 -580 146
rect -542 118 -514 146
rect -476 118 -448 146
rect -410 118 -382 146
rect -344 118 -316 146
rect -278 118 -250 146
rect -212 118 -184 146
rect -146 118 -118 146
rect -80 118 -52 146
rect -14 118 14 146
rect 52 118 80 146
rect 118 118 146 146
rect 184 118 212 146
rect 250 118 278 146
rect 316 118 344 146
rect 382 118 410 146
rect 448 118 476 146
rect 514 118 542 146
rect 580 118 608 146
rect 646 118 674 146
rect 712 118 740 146
rect 778 118 806 146
rect 844 118 872 146
rect 910 118 938 146
rect 976 118 1004 146
rect 1042 118 1070 146
rect 1108 118 1136 146
rect 1174 118 1202 146
rect 1240 118 1268 146
rect 1306 118 1334 146
rect 1372 118 1400 146
rect 1438 118 1466 146
rect 1504 118 1532 146
rect 1570 118 1598 146
rect 1636 118 1664 146
rect 1702 118 1730 146
rect 1768 118 1796 146
rect 1834 118 1862 146
rect 1900 118 1928 146
rect 1966 118 1994 146
rect 2032 118 2060 146
rect 2098 118 2126 146
rect 2164 118 2192 146
rect 2230 118 2258 146
rect 2296 118 2324 146
rect 2362 118 2390 146
rect 2428 118 2456 146
rect 2494 118 2522 146
rect 2560 118 2588 146
rect 2626 118 2654 146
rect 2692 118 2720 146
rect 2758 118 2786 146
rect 2824 118 2852 146
rect 2890 118 2918 146
rect 2956 118 2984 146
rect 3022 118 3050 146
rect 3088 118 3116 146
rect 3154 118 3182 146
rect 3220 118 3248 146
rect 3286 118 3314 146
rect 3352 118 3380 146
rect -3380 52 -3352 80
rect -3314 52 -3286 80
rect -3248 52 -3220 80
rect -3182 52 -3154 80
rect -3116 52 -3088 80
rect -3050 52 -3022 80
rect -2984 52 -2956 80
rect -2918 52 -2890 80
rect -2852 52 -2824 80
rect -2786 52 -2758 80
rect -2720 52 -2692 80
rect -2654 52 -2626 80
rect -2588 52 -2560 80
rect -2522 52 -2494 80
rect -2456 52 -2428 80
rect -2390 52 -2362 80
rect -2324 52 -2296 80
rect -2258 52 -2230 80
rect -2192 52 -2164 80
rect -2126 52 -2098 80
rect -2060 52 -2032 80
rect -1994 52 -1966 80
rect -1928 52 -1900 80
rect -1862 52 -1834 80
rect -1796 52 -1768 80
rect -1730 52 -1702 80
rect -1664 52 -1636 80
rect -1598 52 -1570 80
rect -1532 52 -1504 80
rect -1466 52 -1438 80
rect -1400 52 -1372 80
rect -1334 52 -1306 80
rect -1268 52 -1240 80
rect -1202 52 -1174 80
rect -1136 52 -1108 80
rect -1070 52 -1042 80
rect -1004 52 -976 80
rect -938 52 -910 80
rect -872 52 -844 80
rect -806 52 -778 80
rect -740 52 -712 80
rect -674 52 -646 80
rect -608 52 -580 80
rect -542 52 -514 80
rect -476 52 -448 80
rect -410 52 -382 80
rect -344 52 -316 80
rect -278 52 -250 80
rect -212 52 -184 80
rect -146 52 -118 80
rect -80 52 -52 80
rect -14 52 14 80
rect 52 52 80 80
rect 118 52 146 80
rect 184 52 212 80
rect 250 52 278 80
rect 316 52 344 80
rect 382 52 410 80
rect 448 52 476 80
rect 514 52 542 80
rect 580 52 608 80
rect 646 52 674 80
rect 712 52 740 80
rect 778 52 806 80
rect 844 52 872 80
rect 910 52 938 80
rect 976 52 1004 80
rect 1042 52 1070 80
rect 1108 52 1136 80
rect 1174 52 1202 80
rect 1240 52 1268 80
rect 1306 52 1334 80
rect 1372 52 1400 80
rect 1438 52 1466 80
rect 1504 52 1532 80
rect 1570 52 1598 80
rect 1636 52 1664 80
rect 1702 52 1730 80
rect 1768 52 1796 80
rect 1834 52 1862 80
rect 1900 52 1928 80
rect 1966 52 1994 80
rect 2032 52 2060 80
rect 2098 52 2126 80
rect 2164 52 2192 80
rect 2230 52 2258 80
rect 2296 52 2324 80
rect 2362 52 2390 80
rect 2428 52 2456 80
rect 2494 52 2522 80
rect 2560 52 2588 80
rect 2626 52 2654 80
rect 2692 52 2720 80
rect 2758 52 2786 80
rect 2824 52 2852 80
rect 2890 52 2918 80
rect 2956 52 2984 80
rect 3022 52 3050 80
rect 3088 52 3116 80
rect 3154 52 3182 80
rect 3220 52 3248 80
rect 3286 52 3314 80
rect 3352 52 3380 80
rect -3380 -14 -3352 14
rect -3314 -14 -3286 14
rect -3248 -14 -3220 14
rect -3182 -14 -3154 14
rect -3116 -14 -3088 14
rect -3050 -14 -3022 14
rect -2984 -14 -2956 14
rect -2918 -14 -2890 14
rect -2852 -14 -2824 14
rect -2786 -14 -2758 14
rect -2720 -14 -2692 14
rect -2654 -14 -2626 14
rect -2588 -14 -2560 14
rect -2522 -14 -2494 14
rect -2456 -14 -2428 14
rect -2390 -14 -2362 14
rect -2324 -14 -2296 14
rect -2258 -14 -2230 14
rect -2192 -14 -2164 14
rect -2126 -14 -2098 14
rect -2060 -14 -2032 14
rect -1994 -14 -1966 14
rect -1928 -14 -1900 14
rect -1862 -14 -1834 14
rect -1796 -14 -1768 14
rect -1730 -14 -1702 14
rect -1664 -14 -1636 14
rect -1598 -14 -1570 14
rect -1532 -14 -1504 14
rect -1466 -14 -1438 14
rect -1400 -14 -1372 14
rect -1334 -14 -1306 14
rect -1268 -14 -1240 14
rect -1202 -14 -1174 14
rect -1136 -14 -1108 14
rect -1070 -14 -1042 14
rect -1004 -14 -976 14
rect -938 -14 -910 14
rect -872 -14 -844 14
rect -806 -14 -778 14
rect -740 -14 -712 14
rect -674 -14 -646 14
rect -608 -14 -580 14
rect -542 -14 -514 14
rect -476 -14 -448 14
rect -410 -14 -382 14
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
rect 52 -14 80 14
rect 118 -14 146 14
rect 184 -14 212 14
rect 250 -14 278 14
rect 316 -14 344 14
rect 382 -14 410 14
rect 448 -14 476 14
rect 514 -14 542 14
rect 580 -14 608 14
rect 646 -14 674 14
rect 712 -14 740 14
rect 778 -14 806 14
rect 844 -14 872 14
rect 910 -14 938 14
rect 976 -14 1004 14
rect 1042 -14 1070 14
rect 1108 -14 1136 14
rect 1174 -14 1202 14
rect 1240 -14 1268 14
rect 1306 -14 1334 14
rect 1372 -14 1400 14
rect 1438 -14 1466 14
rect 1504 -14 1532 14
rect 1570 -14 1598 14
rect 1636 -14 1664 14
rect 1702 -14 1730 14
rect 1768 -14 1796 14
rect 1834 -14 1862 14
rect 1900 -14 1928 14
rect 1966 -14 1994 14
rect 2032 -14 2060 14
rect 2098 -14 2126 14
rect 2164 -14 2192 14
rect 2230 -14 2258 14
rect 2296 -14 2324 14
rect 2362 -14 2390 14
rect 2428 -14 2456 14
rect 2494 -14 2522 14
rect 2560 -14 2588 14
rect 2626 -14 2654 14
rect 2692 -14 2720 14
rect 2758 -14 2786 14
rect 2824 -14 2852 14
rect 2890 -14 2918 14
rect 2956 -14 2984 14
rect 3022 -14 3050 14
rect 3088 -14 3116 14
rect 3154 -14 3182 14
rect 3220 -14 3248 14
rect 3286 -14 3314 14
rect 3352 -14 3380 14
rect -3380 -80 -3352 -52
rect -3314 -80 -3286 -52
rect -3248 -80 -3220 -52
rect -3182 -80 -3154 -52
rect -3116 -80 -3088 -52
rect -3050 -80 -3022 -52
rect -2984 -80 -2956 -52
rect -2918 -80 -2890 -52
rect -2852 -80 -2824 -52
rect -2786 -80 -2758 -52
rect -2720 -80 -2692 -52
rect -2654 -80 -2626 -52
rect -2588 -80 -2560 -52
rect -2522 -80 -2494 -52
rect -2456 -80 -2428 -52
rect -2390 -80 -2362 -52
rect -2324 -80 -2296 -52
rect -2258 -80 -2230 -52
rect -2192 -80 -2164 -52
rect -2126 -80 -2098 -52
rect -2060 -80 -2032 -52
rect -1994 -80 -1966 -52
rect -1928 -80 -1900 -52
rect -1862 -80 -1834 -52
rect -1796 -80 -1768 -52
rect -1730 -80 -1702 -52
rect -1664 -80 -1636 -52
rect -1598 -80 -1570 -52
rect -1532 -80 -1504 -52
rect -1466 -80 -1438 -52
rect -1400 -80 -1372 -52
rect -1334 -80 -1306 -52
rect -1268 -80 -1240 -52
rect -1202 -80 -1174 -52
rect -1136 -80 -1108 -52
rect -1070 -80 -1042 -52
rect -1004 -80 -976 -52
rect -938 -80 -910 -52
rect -872 -80 -844 -52
rect -806 -80 -778 -52
rect -740 -80 -712 -52
rect -674 -80 -646 -52
rect -608 -80 -580 -52
rect -542 -80 -514 -52
rect -476 -80 -448 -52
rect -410 -80 -382 -52
rect -344 -80 -316 -52
rect -278 -80 -250 -52
rect -212 -80 -184 -52
rect -146 -80 -118 -52
rect -80 -80 -52 -52
rect -14 -80 14 -52
rect 52 -80 80 -52
rect 118 -80 146 -52
rect 184 -80 212 -52
rect 250 -80 278 -52
rect 316 -80 344 -52
rect 382 -80 410 -52
rect 448 -80 476 -52
rect 514 -80 542 -52
rect 580 -80 608 -52
rect 646 -80 674 -52
rect 712 -80 740 -52
rect 778 -80 806 -52
rect 844 -80 872 -52
rect 910 -80 938 -52
rect 976 -80 1004 -52
rect 1042 -80 1070 -52
rect 1108 -80 1136 -52
rect 1174 -80 1202 -52
rect 1240 -80 1268 -52
rect 1306 -80 1334 -52
rect 1372 -80 1400 -52
rect 1438 -80 1466 -52
rect 1504 -80 1532 -52
rect 1570 -80 1598 -52
rect 1636 -80 1664 -52
rect 1702 -80 1730 -52
rect 1768 -80 1796 -52
rect 1834 -80 1862 -52
rect 1900 -80 1928 -52
rect 1966 -80 1994 -52
rect 2032 -80 2060 -52
rect 2098 -80 2126 -52
rect 2164 -80 2192 -52
rect 2230 -80 2258 -52
rect 2296 -80 2324 -52
rect 2362 -80 2390 -52
rect 2428 -80 2456 -52
rect 2494 -80 2522 -52
rect 2560 -80 2588 -52
rect 2626 -80 2654 -52
rect 2692 -80 2720 -52
rect 2758 -80 2786 -52
rect 2824 -80 2852 -52
rect 2890 -80 2918 -52
rect 2956 -80 2984 -52
rect 3022 -80 3050 -52
rect 3088 -80 3116 -52
rect 3154 -80 3182 -52
rect 3220 -80 3248 -52
rect 3286 -80 3314 -52
rect 3352 -80 3380 -52
rect -3380 -146 -3352 -118
rect -3314 -146 -3286 -118
rect -3248 -146 -3220 -118
rect -3182 -146 -3154 -118
rect -3116 -146 -3088 -118
rect -3050 -146 -3022 -118
rect -2984 -146 -2956 -118
rect -2918 -146 -2890 -118
rect -2852 -146 -2824 -118
rect -2786 -146 -2758 -118
rect -2720 -146 -2692 -118
rect -2654 -146 -2626 -118
rect -2588 -146 -2560 -118
rect -2522 -146 -2494 -118
rect -2456 -146 -2428 -118
rect -2390 -146 -2362 -118
rect -2324 -146 -2296 -118
rect -2258 -146 -2230 -118
rect -2192 -146 -2164 -118
rect -2126 -146 -2098 -118
rect -2060 -146 -2032 -118
rect -1994 -146 -1966 -118
rect -1928 -146 -1900 -118
rect -1862 -146 -1834 -118
rect -1796 -146 -1768 -118
rect -1730 -146 -1702 -118
rect -1664 -146 -1636 -118
rect -1598 -146 -1570 -118
rect -1532 -146 -1504 -118
rect -1466 -146 -1438 -118
rect -1400 -146 -1372 -118
rect -1334 -146 -1306 -118
rect -1268 -146 -1240 -118
rect -1202 -146 -1174 -118
rect -1136 -146 -1108 -118
rect -1070 -146 -1042 -118
rect -1004 -146 -976 -118
rect -938 -146 -910 -118
rect -872 -146 -844 -118
rect -806 -146 -778 -118
rect -740 -146 -712 -118
rect -674 -146 -646 -118
rect -608 -146 -580 -118
rect -542 -146 -514 -118
rect -476 -146 -448 -118
rect -410 -146 -382 -118
rect -344 -146 -316 -118
rect -278 -146 -250 -118
rect -212 -146 -184 -118
rect -146 -146 -118 -118
rect -80 -146 -52 -118
rect -14 -146 14 -118
rect 52 -146 80 -118
rect 118 -146 146 -118
rect 184 -146 212 -118
rect 250 -146 278 -118
rect 316 -146 344 -118
rect 382 -146 410 -118
rect 448 -146 476 -118
rect 514 -146 542 -118
rect 580 -146 608 -118
rect 646 -146 674 -118
rect 712 -146 740 -118
rect 778 -146 806 -118
rect 844 -146 872 -118
rect 910 -146 938 -118
rect 976 -146 1004 -118
rect 1042 -146 1070 -118
rect 1108 -146 1136 -118
rect 1174 -146 1202 -118
rect 1240 -146 1268 -118
rect 1306 -146 1334 -118
rect 1372 -146 1400 -118
rect 1438 -146 1466 -118
rect 1504 -146 1532 -118
rect 1570 -146 1598 -118
rect 1636 -146 1664 -118
rect 1702 -146 1730 -118
rect 1768 -146 1796 -118
rect 1834 -146 1862 -118
rect 1900 -146 1928 -118
rect 1966 -146 1994 -118
rect 2032 -146 2060 -118
rect 2098 -146 2126 -118
rect 2164 -146 2192 -118
rect 2230 -146 2258 -118
rect 2296 -146 2324 -118
rect 2362 -146 2390 -118
rect 2428 -146 2456 -118
rect 2494 -146 2522 -118
rect 2560 -146 2588 -118
rect 2626 -146 2654 -118
rect 2692 -146 2720 -118
rect 2758 -146 2786 -118
rect 2824 -146 2852 -118
rect 2890 -146 2918 -118
rect 2956 -146 2984 -118
rect 3022 -146 3050 -118
rect 3088 -146 3116 -118
rect 3154 -146 3182 -118
rect 3220 -146 3248 -118
rect 3286 -146 3314 -118
rect 3352 -146 3380 -118
rect -3380 -212 -3352 -184
rect -3314 -212 -3286 -184
rect -3248 -212 -3220 -184
rect -3182 -212 -3154 -184
rect -3116 -212 -3088 -184
rect -3050 -212 -3022 -184
rect -2984 -212 -2956 -184
rect -2918 -212 -2890 -184
rect -2852 -212 -2824 -184
rect -2786 -212 -2758 -184
rect -2720 -212 -2692 -184
rect -2654 -212 -2626 -184
rect -2588 -212 -2560 -184
rect -2522 -212 -2494 -184
rect -2456 -212 -2428 -184
rect -2390 -212 -2362 -184
rect -2324 -212 -2296 -184
rect -2258 -212 -2230 -184
rect -2192 -212 -2164 -184
rect -2126 -212 -2098 -184
rect -2060 -212 -2032 -184
rect -1994 -212 -1966 -184
rect -1928 -212 -1900 -184
rect -1862 -212 -1834 -184
rect -1796 -212 -1768 -184
rect -1730 -212 -1702 -184
rect -1664 -212 -1636 -184
rect -1598 -212 -1570 -184
rect -1532 -212 -1504 -184
rect -1466 -212 -1438 -184
rect -1400 -212 -1372 -184
rect -1334 -212 -1306 -184
rect -1268 -212 -1240 -184
rect -1202 -212 -1174 -184
rect -1136 -212 -1108 -184
rect -1070 -212 -1042 -184
rect -1004 -212 -976 -184
rect -938 -212 -910 -184
rect -872 -212 -844 -184
rect -806 -212 -778 -184
rect -740 -212 -712 -184
rect -674 -212 -646 -184
rect -608 -212 -580 -184
rect -542 -212 -514 -184
rect -476 -212 -448 -184
rect -410 -212 -382 -184
rect -344 -212 -316 -184
rect -278 -212 -250 -184
rect -212 -212 -184 -184
rect -146 -212 -118 -184
rect -80 -212 -52 -184
rect -14 -212 14 -184
rect 52 -212 80 -184
rect 118 -212 146 -184
rect 184 -212 212 -184
rect 250 -212 278 -184
rect 316 -212 344 -184
rect 382 -212 410 -184
rect 448 -212 476 -184
rect 514 -212 542 -184
rect 580 -212 608 -184
rect 646 -212 674 -184
rect 712 -212 740 -184
rect 778 -212 806 -184
rect 844 -212 872 -184
rect 910 -212 938 -184
rect 976 -212 1004 -184
rect 1042 -212 1070 -184
rect 1108 -212 1136 -184
rect 1174 -212 1202 -184
rect 1240 -212 1268 -184
rect 1306 -212 1334 -184
rect 1372 -212 1400 -184
rect 1438 -212 1466 -184
rect 1504 -212 1532 -184
rect 1570 -212 1598 -184
rect 1636 -212 1664 -184
rect 1702 -212 1730 -184
rect 1768 -212 1796 -184
rect 1834 -212 1862 -184
rect 1900 -212 1928 -184
rect 1966 -212 1994 -184
rect 2032 -212 2060 -184
rect 2098 -212 2126 -184
rect 2164 -212 2192 -184
rect 2230 -212 2258 -184
rect 2296 -212 2324 -184
rect 2362 -212 2390 -184
rect 2428 -212 2456 -184
rect 2494 -212 2522 -184
rect 2560 -212 2588 -184
rect 2626 -212 2654 -184
rect 2692 -212 2720 -184
rect 2758 -212 2786 -184
rect 2824 -212 2852 -184
rect 2890 -212 2918 -184
rect 2956 -212 2984 -184
rect 3022 -212 3050 -184
rect 3088 -212 3116 -184
rect 3154 -212 3182 -184
rect 3220 -212 3248 -184
rect 3286 -212 3314 -184
rect 3352 -212 3380 -184
rect -3380 -278 -3352 -250
rect -3314 -278 -3286 -250
rect -3248 -278 -3220 -250
rect -3182 -278 -3154 -250
rect -3116 -278 -3088 -250
rect -3050 -278 -3022 -250
rect -2984 -278 -2956 -250
rect -2918 -278 -2890 -250
rect -2852 -278 -2824 -250
rect -2786 -278 -2758 -250
rect -2720 -278 -2692 -250
rect -2654 -278 -2626 -250
rect -2588 -278 -2560 -250
rect -2522 -278 -2494 -250
rect -2456 -278 -2428 -250
rect -2390 -278 -2362 -250
rect -2324 -278 -2296 -250
rect -2258 -278 -2230 -250
rect -2192 -278 -2164 -250
rect -2126 -278 -2098 -250
rect -2060 -278 -2032 -250
rect -1994 -278 -1966 -250
rect -1928 -278 -1900 -250
rect -1862 -278 -1834 -250
rect -1796 -278 -1768 -250
rect -1730 -278 -1702 -250
rect -1664 -278 -1636 -250
rect -1598 -278 -1570 -250
rect -1532 -278 -1504 -250
rect -1466 -278 -1438 -250
rect -1400 -278 -1372 -250
rect -1334 -278 -1306 -250
rect -1268 -278 -1240 -250
rect -1202 -278 -1174 -250
rect -1136 -278 -1108 -250
rect -1070 -278 -1042 -250
rect -1004 -278 -976 -250
rect -938 -278 -910 -250
rect -872 -278 -844 -250
rect -806 -278 -778 -250
rect -740 -278 -712 -250
rect -674 -278 -646 -250
rect -608 -278 -580 -250
rect -542 -278 -514 -250
rect -476 -278 -448 -250
rect -410 -278 -382 -250
rect -344 -278 -316 -250
rect -278 -278 -250 -250
rect -212 -278 -184 -250
rect -146 -278 -118 -250
rect -80 -278 -52 -250
rect -14 -278 14 -250
rect 52 -278 80 -250
rect 118 -278 146 -250
rect 184 -278 212 -250
rect 250 -278 278 -250
rect 316 -278 344 -250
rect 382 -278 410 -250
rect 448 -278 476 -250
rect 514 -278 542 -250
rect 580 -278 608 -250
rect 646 -278 674 -250
rect 712 -278 740 -250
rect 778 -278 806 -250
rect 844 -278 872 -250
rect 910 -278 938 -250
rect 976 -278 1004 -250
rect 1042 -278 1070 -250
rect 1108 -278 1136 -250
rect 1174 -278 1202 -250
rect 1240 -278 1268 -250
rect 1306 -278 1334 -250
rect 1372 -278 1400 -250
rect 1438 -278 1466 -250
rect 1504 -278 1532 -250
rect 1570 -278 1598 -250
rect 1636 -278 1664 -250
rect 1702 -278 1730 -250
rect 1768 -278 1796 -250
rect 1834 -278 1862 -250
rect 1900 -278 1928 -250
rect 1966 -278 1994 -250
rect 2032 -278 2060 -250
rect 2098 -278 2126 -250
rect 2164 -278 2192 -250
rect 2230 -278 2258 -250
rect 2296 -278 2324 -250
rect 2362 -278 2390 -250
rect 2428 -278 2456 -250
rect 2494 -278 2522 -250
rect 2560 -278 2588 -250
rect 2626 -278 2654 -250
rect 2692 -278 2720 -250
rect 2758 -278 2786 -250
rect 2824 -278 2852 -250
rect 2890 -278 2918 -250
rect 2956 -278 2984 -250
rect 3022 -278 3050 -250
rect 3088 -278 3116 -250
rect 3154 -278 3182 -250
rect 3220 -278 3248 -250
rect 3286 -278 3314 -250
rect 3352 -278 3380 -250
rect -3380 -344 -3352 -316
rect -3314 -344 -3286 -316
rect -3248 -344 -3220 -316
rect -3182 -344 -3154 -316
rect -3116 -344 -3088 -316
rect -3050 -344 -3022 -316
rect -2984 -344 -2956 -316
rect -2918 -344 -2890 -316
rect -2852 -344 -2824 -316
rect -2786 -344 -2758 -316
rect -2720 -344 -2692 -316
rect -2654 -344 -2626 -316
rect -2588 -344 -2560 -316
rect -2522 -344 -2494 -316
rect -2456 -344 -2428 -316
rect -2390 -344 -2362 -316
rect -2324 -344 -2296 -316
rect -2258 -344 -2230 -316
rect -2192 -344 -2164 -316
rect -2126 -344 -2098 -316
rect -2060 -344 -2032 -316
rect -1994 -344 -1966 -316
rect -1928 -344 -1900 -316
rect -1862 -344 -1834 -316
rect -1796 -344 -1768 -316
rect -1730 -344 -1702 -316
rect -1664 -344 -1636 -316
rect -1598 -344 -1570 -316
rect -1532 -344 -1504 -316
rect -1466 -344 -1438 -316
rect -1400 -344 -1372 -316
rect -1334 -344 -1306 -316
rect -1268 -344 -1240 -316
rect -1202 -344 -1174 -316
rect -1136 -344 -1108 -316
rect -1070 -344 -1042 -316
rect -1004 -344 -976 -316
rect -938 -344 -910 -316
rect -872 -344 -844 -316
rect -806 -344 -778 -316
rect -740 -344 -712 -316
rect -674 -344 -646 -316
rect -608 -344 -580 -316
rect -542 -344 -514 -316
rect -476 -344 -448 -316
rect -410 -344 -382 -316
rect -344 -344 -316 -316
rect -278 -344 -250 -316
rect -212 -344 -184 -316
rect -146 -344 -118 -316
rect -80 -344 -52 -316
rect -14 -344 14 -316
rect 52 -344 80 -316
rect 118 -344 146 -316
rect 184 -344 212 -316
rect 250 -344 278 -316
rect 316 -344 344 -316
rect 382 -344 410 -316
rect 448 -344 476 -316
rect 514 -344 542 -316
rect 580 -344 608 -316
rect 646 -344 674 -316
rect 712 -344 740 -316
rect 778 -344 806 -316
rect 844 -344 872 -316
rect 910 -344 938 -316
rect 976 -344 1004 -316
rect 1042 -344 1070 -316
rect 1108 -344 1136 -316
rect 1174 -344 1202 -316
rect 1240 -344 1268 -316
rect 1306 -344 1334 -316
rect 1372 -344 1400 -316
rect 1438 -344 1466 -316
rect 1504 -344 1532 -316
rect 1570 -344 1598 -316
rect 1636 -344 1664 -316
rect 1702 -344 1730 -316
rect 1768 -344 1796 -316
rect 1834 -344 1862 -316
rect 1900 -344 1928 -316
rect 1966 -344 1994 -316
rect 2032 -344 2060 -316
rect 2098 -344 2126 -316
rect 2164 -344 2192 -316
rect 2230 -344 2258 -316
rect 2296 -344 2324 -316
rect 2362 -344 2390 -316
rect 2428 -344 2456 -316
rect 2494 -344 2522 -316
rect 2560 -344 2588 -316
rect 2626 -344 2654 -316
rect 2692 -344 2720 -316
rect 2758 -344 2786 -316
rect 2824 -344 2852 -316
rect 2890 -344 2918 -316
rect 2956 -344 2984 -316
rect 3022 -344 3050 -316
rect 3088 -344 3116 -316
rect 3154 -344 3182 -316
rect 3220 -344 3248 -316
rect 3286 -344 3314 -316
rect 3352 -344 3380 -316
<< metal4 >>
rect -3385 344 3385 349
rect -3385 316 -3380 344
rect -3352 316 -3314 344
rect -3286 316 -3248 344
rect -3220 316 -3182 344
rect -3154 316 -3116 344
rect -3088 316 -3050 344
rect -3022 316 -2984 344
rect -2956 316 -2918 344
rect -2890 316 -2852 344
rect -2824 316 -2786 344
rect -2758 316 -2720 344
rect -2692 316 -2654 344
rect -2626 316 -2588 344
rect -2560 316 -2522 344
rect -2494 316 -2456 344
rect -2428 316 -2390 344
rect -2362 316 -2324 344
rect -2296 316 -2258 344
rect -2230 316 -2192 344
rect -2164 316 -2126 344
rect -2098 316 -2060 344
rect -2032 316 -1994 344
rect -1966 316 -1928 344
rect -1900 316 -1862 344
rect -1834 316 -1796 344
rect -1768 316 -1730 344
rect -1702 316 -1664 344
rect -1636 316 -1598 344
rect -1570 316 -1532 344
rect -1504 316 -1466 344
rect -1438 316 -1400 344
rect -1372 316 -1334 344
rect -1306 316 -1268 344
rect -1240 316 -1202 344
rect -1174 316 -1136 344
rect -1108 316 -1070 344
rect -1042 316 -1004 344
rect -976 316 -938 344
rect -910 316 -872 344
rect -844 316 -806 344
rect -778 316 -740 344
rect -712 316 -674 344
rect -646 316 -608 344
rect -580 316 -542 344
rect -514 316 -476 344
rect -448 316 -410 344
rect -382 316 -344 344
rect -316 316 -278 344
rect -250 316 -212 344
rect -184 316 -146 344
rect -118 316 -80 344
rect -52 316 -14 344
rect 14 316 52 344
rect 80 316 118 344
rect 146 316 184 344
rect 212 316 250 344
rect 278 316 316 344
rect 344 316 382 344
rect 410 316 448 344
rect 476 316 514 344
rect 542 316 580 344
rect 608 316 646 344
rect 674 316 712 344
rect 740 316 778 344
rect 806 316 844 344
rect 872 316 910 344
rect 938 316 976 344
rect 1004 316 1042 344
rect 1070 316 1108 344
rect 1136 316 1174 344
rect 1202 316 1240 344
rect 1268 316 1306 344
rect 1334 316 1372 344
rect 1400 316 1438 344
rect 1466 316 1504 344
rect 1532 316 1570 344
rect 1598 316 1636 344
rect 1664 316 1702 344
rect 1730 316 1768 344
rect 1796 316 1834 344
rect 1862 316 1900 344
rect 1928 316 1966 344
rect 1994 316 2032 344
rect 2060 316 2098 344
rect 2126 316 2164 344
rect 2192 316 2230 344
rect 2258 316 2296 344
rect 2324 316 2362 344
rect 2390 316 2428 344
rect 2456 316 2494 344
rect 2522 316 2560 344
rect 2588 316 2626 344
rect 2654 316 2692 344
rect 2720 316 2758 344
rect 2786 316 2824 344
rect 2852 316 2890 344
rect 2918 316 2956 344
rect 2984 316 3022 344
rect 3050 316 3088 344
rect 3116 316 3154 344
rect 3182 316 3220 344
rect 3248 316 3286 344
rect 3314 316 3352 344
rect 3380 316 3385 344
rect -3385 278 3385 316
rect -3385 250 -3380 278
rect -3352 250 -3314 278
rect -3286 250 -3248 278
rect -3220 250 -3182 278
rect -3154 250 -3116 278
rect -3088 250 -3050 278
rect -3022 250 -2984 278
rect -2956 250 -2918 278
rect -2890 250 -2852 278
rect -2824 250 -2786 278
rect -2758 250 -2720 278
rect -2692 250 -2654 278
rect -2626 250 -2588 278
rect -2560 250 -2522 278
rect -2494 250 -2456 278
rect -2428 250 -2390 278
rect -2362 250 -2324 278
rect -2296 250 -2258 278
rect -2230 250 -2192 278
rect -2164 250 -2126 278
rect -2098 250 -2060 278
rect -2032 250 -1994 278
rect -1966 250 -1928 278
rect -1900 250 -1862 278
rect -1834 250 -1796 278
rect -1768 250 -1730 278
rect -1702 250 -1664 278
rect -1636 250 -1598 278
rect -1570 250 -1532 278
rect -1504 250 -1466 278
rect -1438 250 -1400 278
rect -1372 250 -1334 278
rect -1306 250 -1268 278
rect -1240 250 -1202 278
rect -1174 250 -1136 278
rect -1108 250 -1070 278
rect -1042 250 -1004 278
rect -976 250 -938 278
rect -910 250 -872 278
rect -844 250 -806 278
rect -778 250 -740 278
rect -712 250 -674 278
rect -646 250 -608 278
rect -580 250 -542 278
rect -514 250 -476 278
rect -448 250 -410 278
rect -382 250 -344 278
rect -316 250 -278 278
rect -250 250 -212 278
rect -184 250 -146 278
rect -118 250 -80 278
rect -52 250 -14 278
rect 14 250 52 278
rect 80 250 118 278
rect 146 250 184 278
rect 212 250 250 278
rect 278 250 316 278
rect 344 250 382 278
rect 410 250 448 278
rect 476 250 514 278
rect 542 250 580 278
rect 608 250 646 278
rect 674 250 712 278
rect 740 250 778 278
rect 806 250 844 278
rect 872 250 910 278
rect 938 250 976 278
rect 1004 250 1042 278
rect 1070 250 1108 278
rect 1136 250 1174 278
rect 1202 250 1240 278
rect 1268 250 1306 278
rect 1334 250 1372 278
rect 1400 250 1438 278
rect 1466 250 1504 278
rect 1532 250 1570 278
rect 1598 250 1636 278
rect 1664 250 1702 278
rect 1730 250 1768 278
rect 1796 250 1834 278
rect 1862 250 1900 278
rect 1928 250 1966 278
rect 1994 250 2032 278
rect 2060 250 2098 278
rect 2126 250 2164 278
rect 2192 250 2230 278
rect 2258 250 2296 278
rect 2324 250 2362 278
rect 2390 250 2428 278
rect 2456 250 2494 278
rect 2522 250 2560 278
rect 2588 250 2626 278
rect 2654 250 2692 278
rect 2720 250 2758 278
rect 2786 250 2824 278
rect 2852 250 2890 278
rect 2918 250 2956 278
rect 2984 250 3022 278
rect 3050 250 3088 278
rect 3116 250 3154 278
rect 3182 250 3220 278
rect 3248 250 3286 278
rect 3314 250 3352 278
rect 3380 250 3385 278
rect -3385 212 3385 250
rect -3385 184 -3380 212
rect -3352 184 -3314 212
rect -3286 184 -3248 212
rect -3220 184 -3182 212
rect -3154 184 -3116 212
rect -3088 184 -3050 212
rect -3022 184 -2984 212
rect -2956 184 -2918 212
rect -2890 184 -2852 212
rect -2824 184 -2786 212
rect -2758 184 -2720 212
rect -2692 184 -2654 212
rect -2626 184 -2588 212
rect -2560 184 -2522 212
rect -2494 184 -2456 212
rect -2428 184 -2390 212
rect -2362 184 -2324 212
rect -2296 184 -2258 212
rect -2230 184 -2192 212
rect -2164 184 -2126 212
rect -2098 184 -2060 212
rect -2032 184 -1994 212
rect -1966 184 -1928 212
rect -1900 184 -1862 212
rect -1834 184 -1796 212
rect -1768 184 -1730 212
rect -1702 184 -1664 212
rect -1636 184 -1598 212
rect -1570 184 -1532 212
rect -1504 184 -1466 212
rect -1438 184 -1400 212
rect -1372 184 -1334 212
rect -1306 184 -1268 212
rect -1240 184 -1202 212
rect -1174 184 -1136 212
rect -1108 184 -1070 212
rect -1042 184 -1004 212
rect -976 184 -938 212
rect -910 184 -872 212
rect -844 184 -806 212
rect -778 184 -740 212
rect -712 184 -674 212
rect -646 184 -608 212
rect -580 184 -542 212
rect -514 184 -476 212
rect -448 184 -410 212
rect -382 184 -344 212
rect -316 184 -278 212
rect -250 184 -212 212
rect -184 184 -146 212
rect -118 184 -80 212
rect -52 184 -14 212
rect 14 184 52 212
rect 80 184 118 212
rect 146 184 184 212
rect 212 184 250 212
rect 278 184 316 212
rect 344 184 382 212
rect 410 184 448 212
rect 476 184 514 212
rect 542 184 580 212
rect 608 184 646 212
rect 674 184 712 212
rect 740 184 778 212
rect 806 184 844 212
rect 872 184 910 212
rect 938 184 976 212
rect 1004 184 1042 212
rect 1070 184 1108 212
rect 1136 184 1174 212
rect 1202 184 1240 212
rect 1268 184 1306 212
rect 1334 184 1372 212
rect 1400 184 1438 212
rect 1466 184 1504 212
rect 1532 184 1570 212
rect 1598 184 1636 212
rect 1664 184 1702 212
rect 1730 184 1768 212
rect 1796 184 1834 212
rect 1862 184 1900 212
rect 1928 184 1966 212
rect 1994 184 2032 212
rect 2060 184 2098 212
rect 2126 184 2164 212
rect 2192 184 2230 212
rect 2258 184 2296 212
rect 2324 184 2362 212
rect 2390 184 2428 212
rect 2456 184 2494 212
rect 2522 184 2560 212
rect 2588 184 2626 212
rect 2654 184 2692 212
rect 2720 184 2758 212
rect 2786 184 2824 212
rect 2852 184 2890 212
rect 2918 184 2956 212
rect 2984 184 3022 212
rect 3050 184 3088 212
rect 3116 184 3154 212
rect 3182 184 3220 212
rect 3248 184 3286 212
rect 3314 184 3352 212
rect 3380 184 3385 212
rect -3385 146 3385 184
rect -3385 118 -3380 146
rect -3352 118 -3314 146
rect -3286 118 -3248 146
rect -3220 118 -3182 146
rect -3154 118 -3116 146
rect -3088 118 -3050 146
rect -3022 118 -2984 146
rect -2956 118 -2918 146
rect -2890 118 -2852 146
rect -2824 118 -2786 146
rect -2758 118 -2720 146
rect -2692 118 -2654 146
rect -2626 118 -2588 146
rect -2560 118 -2522 146
rect -2494 118 -2456 146
rect -2428 118 -2390 146
rect -2362 118 -2324 146
rect -2296 118 -2258 146
rect -2230 118 -2192 146
rect -2164 118 -2126 146
rect -2098 118 -2060 146
rect -2032 118 -1994 146
rect -1966 118 -1928 146
rect -1900 118 -1862 146
rect -1834 118 -1796 146
rect -1768 118 -1730 146
rect -1702 118 -1664 146
rect -1636 118 -1598 146
rect -1570 118 -1532 146
rect -1504 118 -1466 146
rect -1438 118 -1400 146
rect -1372 118 -1334 146
rect -1306 118 -1268 146
rect -1240 118 -1202 146
rect -1174 118 -1136 146
rect -1108 118 -1070 146
rect -1042 118 -1004 146
rect -976 118 -938 146
rect -910 118 -872 146
rect -844 118 -806 146
rect -778 118 -740 146
rect -712 118 -674 146
rect -646 118 -608 146
rect -580 118 -542 146
rect -514 118 -476 146
rect -448 118 -410 146
rect -382 118 -344 146
rect -316 118 -278 146
rect -250 118 -212 146
rect -184 118 -146 146
rect -118 118 -80 146
rect -52 118 -14 146
rect 14 118 52 146
rect 80 118 118 146
rect 146 118 184 146
rect 212 118 250 146
rect 278 118 316 146
rect 344 118 382 146
rect 410 118 448 146
rect 476 118 514 146
rect 542 118 580 146
rect 608 118 646 146
rect 674 118 712 146
rect 740 118 778 146
rect 806 118 844 146
rect 872 118 910 146
rect 938 118 976 146
rect 1004 118 1042 146
rect 1070 118 1108 146
rect 1136 118 1174 146
rect 1202 118 1240 146
rect 1268 118 1306 146
rect 1334 118 1372 146
rect 1400 118 1438 146
rect 1466 118 1504 146
rect 1532 118 1570 146
rect 1598 118 1636 146
rect 1664 118 1702 146
rect 1730 118 1768 146
rect 1796 118 1834 146
rect 1862 118 1900 146
rect 1928 118 1966 146
rect 1994 118 2032 146
rect 2060 118 2098 146
rect 2126 118 2164 146
rect 2192 118 2230 146
rect 2258 118 2296 146
rect 2324 118 2362 146
rect 2390 118 2428 146
rect 2456 118 2494 146
rect 2522 118 2560 146
rect 2588 118 2626 146
rect 2654 118 2692 146
rect 2720 118 2758 146
rect 2786 118 2824 146
rect 2852 118 2890 146
rect 2918 118 2956 146
rect 2984 118 3022 146
rect 3050 118 3088 146
rect 3116 118 3154 146
rect 3182 118 3220 146
rect 3248 118 3286 146
rect 3314 118 3352 146
rect 3380 118 3385 146
rect -3385 80 3385 118
rect -3385 52 -3380 80
rect -3352 52 -3314 80
rect -3286 52 -3248 80
rect -3220 52 -3182 80
rect -3154 52 -3116 80
rect -3088 52 -3050 80
rect -3022 52 -2984 80
rect -2956 52 -2918 80
rect -2890 52 -2852 80
rect -2824 52 -2786 80
rect -2758 52 -2720 80
rect -2692 52 -2654 80
rect -2626 52 -2588 80
rect -2560 52 -2522 80
rect -2494 52 -2456 80
rect -2428 52 -2390 80
rect -2362 52 -2324 80
rect -2296 52 -2258 80
rect -2230 52 -2192 80
rect -2164 52 -2126 80
rect -2098 52 -2060 80
rect -2032 52 -1994 80
rect -1966 52 -1928 80
rect -1900 52 -1862 80
rect -1834 52 -1796 80
rect -1768 52 -1730 80
rect -1702 52 -1664 80
rect -1636 52 -1598 80
rect -1570 52 -1532 80
rect -1504 52 -1466 80
rect -1438 52 -1400 80
rect -1372 52 -1334 80
rect -1306 52 -1268 80
rect -1240 52 -1202 80
rect -1174 52 -1136 80
rect -1108 52 -1070 80
rect -1042 52 -1004 80
rect -976 52 -938 80
rect -910 52 -872 80
rect -844 52 -806 80
rect -778 52 -740 80
rect -712 52 -674 80
rect -646 52 -608 80
rect -580 52 -542 80
rect -514 52 -476 80
rect -448 52 -410 80
rect -382 52 -344 80
rect -316 52 -278 80
rect -250 52 -212 80
rect -184 52 -146 80
rect -118 52 -80 80
rect -52 52 -14 80
rect 14 52 52 80
rect 80 52 118 80
rect 146 52 184 80
rect 212 52 250 80
rect 278 52 316 80
rect 344 52 382 80
rect 410 52 448 80
rect 476 52 514 80
rect 542 52 580 80
rect 608 52 646 80
rect 674 52 712 80
rect 740 52 778 80
rect 806 52 844 80
rect 872 52 910 80
rect 938 52 976 80
rect 1004 52 1042 80
rect 1070 52 1108 80
rect 1136 52 1174 80
rect 1202 52 1240 80
rect 1268 52 1306 80
rect 1334 52 1372 80
rect 1400 52 1438 80
rect 1466 52 1504 80
rect 1532 52 1570 80
rect 1598 52 1636 80
rect 1664 52 1702 80
rect 1730 52 1768 80
rect 1796 52 1834 80
rect 1862 52 1900 80
rect 1928 52 1966 80
rect 1994 52 2032 80
rect 2060 52 2098 80
rect 2126 52 2164 80
rect 2192 52 2230 80
rect 2258 52 2296 80
rect 2324 52 2362 80
rect 2390 52 2428 80
rect 2456 52 2494 80
rect 2522 52 2560 80
rect 2588 52 2626 80
rect 2654 52 2692 80
rect 2720 52 2758 80
rect 2786 52 2824 80
rect 2852 52 2890 80
rect 2918 52 2956 80
rect 2984 52 3022 80
rect 3050 52 3088 80
rect 3116 52 3154 80
rect 3182 52 3220 80
rect 3248 52 3286 80
rect 3314 52 3352 80
rect 3380 52 3385 80
rect -3385 14 3385 52
rect -3385 -14 -3380 14
rect -3352 -14 -3314 14
rect -3286 -14 -3248 14
rect -3220 -14 -3182 14
rect -3154 -14 -3116 14
rect -3088 -14 -3050 14
rect -3022 -14 -2984 14
rect -2956 -14 -2918 14
rect -2890 -14 -2852 14
rect -2824 -14 -2786 14
rect -2758 -14 -2720 14
rect -2692 -14 -2654 14
rect -2626 -14 -2588 14
rect -2560 -14 -2522 14
rect -2494 -14 -2456 14
rect -2428 -14 -2390 14
rect -2362 -14 -2324 14
rect -2296 -14 -2258 14
rect -2230 -14 -2192 14
rect -2164 -14 -2126 14
rect -2098 -14 -2060 14
rect -2032 -14 -1994 14
rect -1966 -14 -1928 14
rect -1900 -14 -1862 14
rect -1834 -14 -1796 14
rect -1768 -14 -1730 14
rect -1702 -14 -1664 14
rect -1636 -14 -1598 14
rect -1570 -14 -1532 14
rect -1504 -14 -1466 14
rect -1438 -14 -1400 14
rect -1372 -14 -1334 14
rect -1306 -14 -1268 14
rect -1240 -14 -1202 14
rect -1174 -14 -1136 14
rect -1108 -14 -1070 14
rect -1042 -14 -1004 14
rect -976 -14 -938 14
rect -910 -14 -872 14
rect -844 -14 -806 14
rect -778 -14 -740 14
rect -712 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 52 14
rect 80 -14 118 14
rect 146 -14 184 14
rect 212 -14 250 14
rect 278 -14 316 14
rect 344 -14 382 14
rect 410 -14 448 14
rect 476 -14 514 14
rect 542 -14 580 14
rect 608 -14 646 14
rect 674 -14 712 14
rect 740 -14 778 14
rect 806 -14 844 14
rect 872 -14 910 14
rect 938 -14 976 14
rect 1004 -14 1042 14
rect 1070 -14 1108 14
rect 1136 -14 1174 14
rect 1202 -14 1240 14
rect 1268 -14 1306 14
rect 1334 -14 1372 14
rect 1400 -14 1438 14
rect 1466 -14 1504 14
rect 1532 -14 1570 14
rect 1598 -14 1636 14
rect 1664 -14 1702 14
rect 1730 -14 1768 14
rect 1796 -14 1834 14
rect 1862 -14 1900 14
rect 1928 -14 1966 14
rect 1994 -14 2032 14
rect 2060 -14 2098 14
rect 2126 -14 2164 14
rect 2192 -14 2230 14
rect 2258 -14 2296 14
rect 2324 -14 2362 14
rect 2390 -14 2428 14
rect 2456 -14 2494 14
rect 2522 -14 2560 14
rect 2588 -14 2626 14
rect 2654 -14 2692 14
rect 2720 -14 2758 14
rect 2786 -14 2824 14
rect 2852 -14 2890 14
rect 2918 -14 2956 14
rect 2984 -14 3022 14
rect 3050 -14 3088 14
rect 3116 -14 3154 14
rect 3182 -14 3220 14
rect 3248 -14 3286 14
rect 3314 -14 3352 14
rect 3380 -14 3385 14
rect -3385 -52 3385 -14
rect -3385 -80 -3380 -52
rect -3352 -80 -3314 -52
rect -3286 -80 -3248 -52
rect -3220 -80 -3182 -52
rect -3154 -80 -3116 -52
rect -3088 -80 -3050 -52
rect -3022 -80 -2984 -52
rect -2956 -80 -2918 -52
rect -2890 -80 -2852 -52
rect -2824 -80 -2786 -52
rect -2758 -80 -2720 -52
rect -2692 -80 -2654 -52
rect -2626 -80 -2588 -52
rect -2560 -80 -2522 -52
rect -2494 -80 -2456 -52
rect -2428 -80 -2390 -52
rect -2362 -80 -2324 -52
rect -2296 -80 -2258 -52
rect -2230 -80 -2192 -52
rect -2164 -80 -2126 -52
rect -2098 -80 -2060 -52
rect -2032 -80 -1994 -52
rect -1966 -80 -1928 -52
rect -1900 -80 -1862 -52
rect -1834 -80 -1796 -52
rect -1768 -80 -1730 -52
rect -1702 -80 -1664 -52
rect -1636 -80 -1598 -52
rect -1570 -80 -1532 -52
rect -1504 -80 -1466 -52
rect -1438 -80 -1400 -52
rect -1372 -80 -1334 -52
rect -1306 -80 -1268 -52
rect -1240 -80 -1202 -52
rect -1174 -80 -1136 -52
rect -1108 -80 -1070 -52
rect -1042 -80 -1004 -52
rect -976 -80 -938 -52
rect -910 -80 -872 -52
rect -844 -80 -806 -52
rect -778 -80 -740 -52
rect -712 -80 -674 -52
rect -646 -80 -608 -52
rect -580 -80 -542 -52
rect -514 -80 -476 -52
rect -448 -80 -410 -52
rect -382 -80 -344 -52
rect -316 -80 -278 -52
rect -250 -80 -212 -52
rect -184 -80 -146 -52
rect -118 -80 -80 -52
rect -52 -80 -14 -52
rect 14 -80 52 -52
rect 80 -80 118 -52
rect 146 -80 184 -52
rect 212 -80 250 -52
rect 278 -80 316 -52
rect 344 -80 382 -52
rect 410 -80 448 -52
rect 476 -80 514 -52
rect 542 -80 580 -52
rect 608 -80 646 -52
rect 674 -80 712 -52
rect 740 -80 778 -52
rect 806 -80 844 -52
rect 872 -80 910 -52
rect 938 -80 976 -52
rect 1004 -80 1042 -52
rect 1070 -80 1108 -52
rect 1136 -80 1174 -52
rect 1202 -80 1240 -52
rect 1268 -80 1306 -52
rect 1334 -80 1372 -52
rect 1400 -80 1438 -52
rect 1466 -80 1504 -52
rect 1532 -80 1570 -52
rect 1598 -80 1636 -52
rect 1664 -80 1702 -52
rect 1730 -80 1768 -52
rect 1796 -80 1834 -52
rect 1862 -80 1900 -52
rect 1928 -80 1966 -52
rect 1994 -80 2032 -52
rect 2060 -80 2098 -52
rect 2126 -80 2164 -52
rect 2192 -80 2230 -52
rect 2258 -80 2296 -52
rect 2324 -80 2362 -52
rect 2390 -80 2428 -52
rect 2456 -80 2494 -52
rect 2522 -80 2560 -52
rect 2588 -80 2626 -52
rect 2654 -80 2692 -52
rect 2720 -80 2758 -52
rect 2786 -80 2824 -52
rect 2852 -80 2890 -52
rect 2918 -80 2956 -52
rect 2984 -80 3022 -52
rect 3050 -80 3088 -52
rect 3116 -80 3154 -52
rect 3182 -80 3220 -52
rect 3248 -80 3286 -52
rect 3314 -80 3352 -52
rect 3380 -80 3385 -52
rect -3385 -118 3385 -80
rect -3385 -146 -3380 -118
rect -3352 -146 -3314 -118
rect -3286 -146 -3248 -118
rect -3220 -146 -3182 -118
rect -3154 -146 -3116 -118
rect -3088 -146 -3050 -118
rect -3022 -146 -2984 -118
rect -2956 -146 -2918 -118
rect -2890 -146 -2852 -118
rect -2824 -146 -2786 -118
rect -2758 -146 -2720 -118
rect -2692 -146 -2654 -118
rect -2626 -146 -2588 -118
rect -2560 -146 -2522 -118
rect -2494 -146 -2456 -118
rect -2428 -146 -2390 -118
rect -2362 -146 -2324 -118
rect -2296 -146 -2258 -118
rect -2230 -146 -2192 -118
rect -2164 -146 -2126 -118
rect -2098 -146 -2060 -118
rect -2032 -146 -1994 -118
rect -1966 -146 -1928 -118
rect -1900 -146 -1862 -118
rect -1834 -146 -1796 -118
rect -1768 -146 -1730 -118
rect -1702 -146 -1664 -118
rect -1636 -146 -1598 -118
rect -1570 -146 -1532 -118
rect -1504 -146 -1466 -118
rect -1438 -146 -1400 -118
rect -1372 -146 -1334 -118
rect -1306 -146 -1268 -118
rect -1240 -146 -1202 -118
rect -1174 -146 -1136 -118
rect -1108 -146 -1070 -118
rect -1042 -146 -1004 -118
rect -976 -146 -938 -118
rect -910 -146 -872 -118
rect -844 -146 -806 -118
rect -778 -146 -740 -118
rect -712 -146 -674 -118
rect -646 -146 -608 -118
rect -580 -146 -542 -118
rect -514 -146 -476 -118
rect -448 -146 -410 -118
rect -382 -146 -344 -118
rect -316 -146 -278 -118
rect -250 -146 -212 -118
rect -184 -146 -146 -118
rect -118 -146 -80 -118
rect -52 -146 -14 -118
rect 14 -146 52 -118
rect 80 -146 118 -118
rect 146 -146 184 -118
rect 212 -146 250 -118
rect 278 -146 316 -118
rect 344 -146 382 -118
rect 410 -146 448 -118
rect 476 -146 514 -118
rect 542 -146 580 -118
rect 608 -146 646 -118
rect 674 -146 712 -118
rect 740 -146 778 -118
rect 806 -146 844 -118
rect 872 -146 910 -118
rect 938 -146 976 -118
rect 1004 -146 1042 -118
rect 1070 -146 1108 -118
rect 1136 -146 1174 -118
rect 1202 -146 1240 -118
rect 1268 -146 1306 -118
rect 1334 -146 1372 -118
rect 1400 -146 1438 -118
rect 1466 -146 1504 -118
rect 1532 -146 1570 -118
rect 1598 -146 1636 -118
rect 1664 -146 1702 -118
rect 1730 -146 1768 -118
rect 1796 -146 1834 -118
rect 1862 -146 1900 -118
rect 1928 -146 1966 -118
rect 1994 -146 2032 -118
rect 2060 -146 2098 -118
rect 2126 -146 2164 -118
rect 2192 -146 2230 -118
rect 2258 -146 2296 -118
rect 2324 -146 2362 -118
rect 2390 -146 2428 -118
rect 2456 -146 2494 -118
rect 2522 -146 2560 -118
rect 2588 -146 2626 -118
rect 2654 -146 2692 -118
rect 2720 -146 2758 -118
rect 2786 -146 2824 -118
rect 2852 -146 2890 -118
rect 2918 -146 2956 -118
rect 2984 -146 3022 -118
rect 3050 -146 3088 -118
rect 3116 -146 3154 -118
rect 3182 -146 3220 -118
rect 3248 -146 3286 -118
rect 3314 -146 3352 -118
rect 3380 -146 3385 -118
rect -3385 -184 3385 -146
rect -3385 -212 -3380 -184
rect -3352 -212 -3314 -184
rect -3286 -212 -3248 -184
rect -3220 -212 -3182 -184
rect -3154 -212 -3116 -184
rect -3088 -212 -3050 -184
rect -3022 -212 -2984 -184
rect -2956 -212 -2918 -184
rect -2890 -212 -2852 -184
rect -2824 -212 -2786 -184
rect -2758 -212 -2720 -184
rect -2692 -212 -2654 -184
rect -2626 -212 -2588 -184
rect -2560 -212 -2522 -184
rect -2494 -212 -2456 -184
rect -2428 -212 -2390 -184
rect -2362 -212 -2324 -184
rect -2296 -212 -2258 -184
rect -2230 -212 -2192 -184
rect -2164 -212 -2126 -184
rect -2098 -212 -2060 -184
rect -2032 -212 -1994 -184
rect -1966 -212 -1928 -184
rect -1900 -212 -1862 -184
rect -1834 -212 -1796 -184
rect -1768 -212 -1730 -184
rect -1702 -212 -1664 -184
rect -1636 -212 -1598 -184
rect -1570 -212 -1532 -184
rect -1504 -212 -1466 -184
rect -1438 -212 -1400 -184
rect -1372 -212 -1334 -184
rect -1306 -212 -1268 -184
rect -1240 -212 -1202 -184
rect -1174 -212 -1136 -184
rect -1108 -212 -1070 -184
rect -1042 -212 -1004 -184
rect -976 -212 -938 -184
rect -910 -212 -872 -184
rect -844 -212 -806 -184
rect -778 -212 -740 -184
rect -712 -212 -674 -184
rect -646 -212 -608 -184
rect -580 -212 -542 -184
rect -514 -212 -476 -184
rect -448 -212 -410 -184
rect -382 -212 -344 -184
rect -316 -212 -278 -184
rect -250 -212 -212 -184
rect -184 -212 -146 -184
rect -118 -212 -80 -184
rect -52 -212 -14 -184
rect 14 -212 52 -184
rect 80 -212 118 -184
rect 146 -212 184 -184
rect 212 -212 250 -184
rect 278 -212 316 -184
rect 344 -212 382 -184
rect 410 -212 448 -184
rect 476 -212 514 -184
rect 542 -212 580 -184
rect 608 -212 646 -184
rect 674 -212 712 -184
rect 740 -212 778 -184
rect 806 -212 844 -184
rect 872 -212 910 -184
rect 938 -212 976 -184
rect 1004 -212 1042 -184
rect 1070 -212 1108 -184
rect 1136 -212 1174 -184
rect 1202 -212 1240 -184
rect 1268 -212 1306 -184
rect 1334 -212 1372 -184
rect 1400 -212 1438 -184
rect 1466 -212 1504 -184
rect 1532 -212 1570 -184
rect 1598 -212 1636 -184
rect 1664 -212 1702 -184
rect 1730 -212 1768 -184
rect 1796 -212 1834 -184
rect 1862 -212 1900 -184
rect 1928 -212 1966 -184
rect 1994 -212 2032 -184
rect 2060 -212 2098 -184
rect 2126 -212 2164 -184
rect 2192 -212 2230 -184
rect 2258 -212 2296 -184
rect 2324 -212 2362 -184
rect 2390 -212 2428 -184
rect 2456 -212 2494 -184
rect 2522 -212 2560 -184
rect 2588 -212 2626 -184
rect 2654 -212 2692 -184
rect 2720 -212 2758 -184
rect 2786 -212 2824 -184
rect 2852 -212 2890 -184
rect 2918 -212 2956 -184
rect 2984 -212 3022 -184
rect 3050 -212 3088 -184
rect 3116 -212 3154 -184
rect 3182 -212 3220 -184
rect 3248 -212 3286 -184
rect 3314 -212 3352 -184
rect 3380 -212 3385 -184
rect -3385 -250 3385 -212
rect -3385 -278 -3380 -250
rect -3352 -278 -3314 -250
rect -3286 -278 -3248 -250
rect -3220 -278 -3182 -250
rect -3154 -278 -3116 -250
rect -3088 -278 -3050 -250
rect -3022 -278 -2984 -250
rect -2956 -278 -2918 -250
rect -2890 -278 -2852 -250
rect -2824 -278 -2786 -250
rect -2758 -278 -2720 -250
rect -2692 -278 -2654 -250
rect -2626 -278 -2588 -250
rect -2560 -278 -2522 -250
rect -2494 -278 -2456 -250
rect -2428 -278 -2390 -250
rect -2362 -278 -2324 -250
rect -2296 -278 -2258 -250
rect -2230 -278 -2192 -250
rect -2164 -278 -2126 -250
rect -2098 -278 -2060 -250
rect -2032 -278 -1994 -250
rect -1966 -278 -1928 -250
rect -1900 -278 -1862 -250
rect -1834 -278 -1796 -250
rect -1768 -278 -1730 -250
rect -1702 -278 -1664 -250
rect -1636 -278 -1598 -250
rect -1570 -278 -1532 -250
rect -1504 -278 -1466 -250
rect -1438 -278 -1400 -250
rect -1372 -278 -1334 -250
rect -1306 -278 -1268 -250
rect -1240 -278 -1202 -250
rect -1174 -278 -1136 -250
rect -1108 -278 -1070 -250
rect -1042 -278 -1004 -250
rect -976 -278 -938 -250
rect -910 -278 -872 -250
rect -844 -278 -806 -250
rect -778 -278 -740 -250
rect -712 -278 -674 -250
rect -646 -278 -608 -250
rect -580 -278 -542 -250
rect -514 -278 -476 -250
rect -448 -278 -410 -250
rect -382 -278 -344 -250
rect -316 -278 -278 -250
rect -250 -278 -212 -250
rect -184 -278 -146 -250
rect -118 -278 -80 -250
rect -52 -278 -14 -250
rect 14 -278 52 -250
rect 80 -278 118 -250
rect 146 -278 184 -250
rect 212 -278 250 -250
rect 278 -278 316 -250
rect 344 -278 382 -250
rect 410 -278 448 -250
rect 476 -278 514 -250
rect 542 -278 580 -250
rect 608 -278 646 -250
rect 674 -278 712 -250
rect 740 -278 778 -250
rect 806 -278 844 -250
rect 872 -278 910 -250
rect 938 -278 976 -250
rect 1004 -278 1042 -250
rect 1070 -278 1108 -250
rect 1136 -278 1174 -250
rect 1202 -278 1240 -250
rect 1268 -278 1306 -250
rect 1334 -278 1372 -250
rect 1400 -278 1438 -250
rect 1466 -278 1504 -250
rect 1532 -278 1570 -250
rect 1598 -278 1636 -250
rect 1664 -278 1702 -250
rect 1730 -278 1768 -250
rect 1796 -278 1834 -250
rect 1862 -278 1900 -250
rect 1928 -278 1966 -250
rect 1994 -278 2032 -250
rect 2060 -278 2098 -250
rect 2126 -278 2164 -250
rect 2192 -278 2230 -250
rect 2258 -278 2296 -250
rect 2324 -278 2362 -250
rect 2390 -278 2428 -250
rect 2456 -278 2494 -250
rect 2522 -278 2560 -250
rect 2588 -278 2626 -250
rect 2654 -278 2692 -250
rect 2720 -278 2758 -250
rect 2786 -278 2824 -250
rect 2852 -278 2890 -250
rect 2918 -278 2956 -250
rect 2984 -278 3022 -250
rect 3050 -278 3088 -250
rect 3116 -278 3154 -250
rect 3182 -278 3220 -250
rect 3248 -278 3286 -250
rect 3314 -278 3352 -250
rect 3380 -278 3385 -250
rect -3385 -316 3385 -278
rect -3385 -344 -3380 -316
rect -3352 -344 -3314 -316
rect -3286 -344 -3248 -316
rect -3220 -344 -3182 -316
rect -3154 -344 -3116 -316
rect -3088 -344 -3050 -316
rect -3022 -344 -2984 -316
rect -2956 -344 -2918 -316
rect -2890 -344 -2852 -316
rect -2824 -344 -2786 -316
rect -2758 -344 -2720 -316
rect -2692 -344 -2654 -316
rect -2626 -344 -2588 -316
rect -2560 -344 -2522 -316
rect -2494 -344 -2456 -316
rect -2428 -344 -2390 -316
rect -2362 -344 -2324 -316
rect -2296 -344 -2258 -316
rect -2230 -344 -2192 -316
rect -2164 -344 -2126 -316
rect -2098 -344 -2060 -316
rect -2032 -344 -1994 -316
rect -1966 -344 -1928 -316
rect -1900 -344 -1862 -316
rect -1834 -344 -1796 -316
rect -1768 -344 -1730 -316
rect -1702 -344 -1664 -316
rect -1636 -344 -1598 -316
rect -1570 -344 -1532 -316
rect -1504 -344 -1466 -316
rect -1438 -344 -1400 -316
rect -1372 -344 -1334 -316
rect -1306 -344 -1268 -316
rect -1240 -344 -1202 -316
rect -1174 -344 -1136 -316
rect -1108 -344 -1070 -316
rect -1042 -344 -1004 -316
rect -976 -344 -938 -316
rect -910 -344 -872 -316
rect -844 -344 -806 -316
rect -778 -344 -740 -316
rect -712 -344 -674 -316
rect -646 -344 -608 -316
rect -580 -344 -542 -316
rect -514 -344 -476 -316
rect -448 -344 -410 -316
rect -382 -344 -344 -316
rect -316 -344 -278 -316
rect -250 -344 -212 -316
rect -184 -344 -146 -316
rect -118 -344 -80 -316
rect -52 -344 -14 -316
rect 14 -344 52 -316
rect 80 -344 118 -316
rect 146 -344 184 -316
rect 212 -344 250 -316
rect 278 -344 316 -316
rect 344 -344 382 -316
rect 410 -344 448 -316
rect 476 -344 514 -316
rect 542 -344 580 -316
rect 608 -344 646 -316
rect 674 -344 712 -316
rect 740 -344 778 -316
rect 806 -344 844 -316
rect 872 -344 910 -316
rect 938 -344 976 -316
rect 1004 -344 1042 -316
rect 1070 -344 1108 -316
rect 1136 -344 1174 -316
rect 1202 -344 1240 -316
rect 1268 -344 1306 -316
rect 1334 -344 1372 -316
rect 1400 -344 1438 -316
rect 1466 -344 1504 -316
rect 1532 -344 1570 -316
rect 1598 -344 1636 -316
rect 1664 -344 1702 -316
rect 1730 -344 1768 -316
rect 1796 -344 1834 -316
rect 1862 -344 1900 -316
rect 1928 -344 1966 -316
rect 1994 -344 2032 -316
rect 2060 -344 2098 -316
rect 2126 -344 2164 -316
rect 2192 -344 2230 -316
rect 2258 -344 2296 -316
rect 2324 -344 2362 -316
rect 2390 -344 2428 -316
rect 2456 -344 2494 -316
rect 2522 -344 2560 -316
rect 2588 -344 2626 -316
rect 2654 -344 2692 -316
rect 2720 -344 2758 -316
rect 2786 -344 2824 -316
rect 2852 -344 2890 -316
rect 2918 -344 2956 -316
rect 2984 -344 3022 -316
rect 3050 -344 3088 -316
rect 3116 -344 3154 -316
rect 3182 -344 3220 -316
rect 3248 -344 3286 -316
rect 3314 -344 3352 -316
rect 3380 -344 3385 -316
rect -3385 -349 3385 -344
<< end >>
