magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -1952 -1556 4468 10220
<< mvnmos >>
rect 206 532 436 8132
rect 2080 532 2310 8132
<< mvndiff >>
rect 48 8117 150 8132
rect 48 551 61 8117
rect 107 551 150 8117
rect 48 532 150 551
rect 1192 8117 1324 8132
rect 1192 551 1235 8117
rect 1281 551 1324 8117
rect 1192 532 1324 551
rect 2366 8117 2468 8132
rect 2366 551 2409 8117
rect 2455 551 2468 8117
rect 2366 532 2468 551
<< mvndiffc >>
rect 61 551 107 8117
rect 1235 551 1281 8117
rect 2409 551 2455 8117
<< polysilicon >>
rect 206 8132 436 8220
rect 2080 8132 2310 8220
rect 206 444 436 532
rect 2080 444 2310 532
<< mvndiffres >>
rect 150 532 206 8132
rect 436 532 1192 8132
rect 1324 532 2080 8132
rect 2310 532 2366 8132
<< metal1 >>
rect 61 8117 107 8132
rect 61 532 107 551
rect 1235 8117 1281 8132
rect 1235 532 1281 551
rect 2409 8117 2455 8132
rect 2409 532 2455 551
<< end >>
