magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2002 -2052 4031 3117
<< nwell >>
rect 0 1109 2000 1117
rect 1108 1013 2000 1109
<< pwell >>
rect -2 134 282 494
rect 830 134 1170 492
<< psubdiff >>
rect 1428 21 1661 41
rect 1428 -25 1473 21
rect 1519 -25 1661 21
rect 1428 -40 1661 -25
<< psubdiffcont >>
rect 1473 -25 1519 21
<< polysilicon >>
rect 1282 908 1826 979
rect 1282 616 1394 650
rect 1282 570 1314 616
rect 1360 570 1394 616
rect 1282 550 1394 570
rect 1498 508 1610 529
rect 1498 462 1533 508
rect 1579 462 1610 508
rect 1498 443 1610 462
rect 1282 109 1826 180
<< polycontact >>
rect 1314 570 1360 616
rect 1533 462 1579 508
<< metal1 >>
rect 78 1065 1921 1093
rect 82 1039 1921 1065
rect 82 1020 1192 1039
rect 1207 927 1685 973
rect 1207 663 1253 927
rect 1423 803 1469 881
rect 1396 789 1487 803
rect 1396 737 1416 789
rect 1468 737 1487 789
rect 1396 724 1487 737
rect 1297 616 1373 632
rect 1297 615 1314 616
rect 793 613 1314 615
rect 868 570 1314 613
rect 1360 570 1373 616
rect 868 569 1373 570
rect 1282 560 1373 569
rect 1297 552 1373 560
rect 199 474 265 520
rect 354 519 465 521
rect 354 470 466 519
rect 414 158 466 470
rect 640 475 885 521
rect 640 158 687 475
rect 839 439 885 475
rect 1007 444 1103 457
rect 1007 439 1031 444
rect 839 393 1031 439
rect 1007 392 1031 393
rect 1083 392 1103 444
rect 1007 376 1103 392
rect 414 111 687 158
rect 1207 151 1253 414
rect 1423 202 1469 724
rect 1516 519 1592 527
rect 1516 511 1593 519
rect 1516 459 1532 511
rect 1584 459 1593 511
rect 1516 447 1593 459
rect 1516 442 1592 447
rect 1639 151 1685 927
rect 1855 803 1901 881
rect 1829 789 1919 803
rect 1829 737 1848 789
rect 1900 737 1919 789
rect 1829 723 1919 737
rect 1855 540 1901 723
rect 1855 494 2031 540
rect 1855 202 1901 494
rect 1074 105 1685 151
rect 1065 21 1951 41
rect 1065 -25 1473 21
rect 1519 -25 1951 21
rect 1065 -40 1951 -25
<< via1 >>
rect 1416 737 1468 789
rect 1031 392 1083 444
rect 1532 508 1584 511
rect 1532 462 1533 508
rect 1533 462 1579 508
rect 1579 462 1584 508
rect 1532 459 1584 462
rect 1848 737 1900 789
<< metal2 >>
rect 1396 792 1487 803
rect 1829 792 1919 803
rect 1396 789 1919 792
rect 1396 737 1416 789
rect 1468 737 1848 789
rect 1900 737 1919 789
rect 1396 730 1919 737
rect 1396 724 1487 730
rect 1829 723 1919 730
rect 1512 511 1605 528
rect 1512 459 1532 511
rect 1584 459 1605 511
rect 1007 454 1103 457
rect 1512 454 1605 459
rect 1007 444 1605 454
rect 1007 392 1031 444
rect 1083 440 1605 444
rect 1083 392 1602 440
rect 1007 383 1602 392
rect 1007 376 1103 383
use inverter_magic  inverter_magic_0
timestamp 1713185578
transform 1 0 0 0 1 529
box 0 -569 1108 580
use nmos_3p3_G2UGVV  nmos_3p3_G2UGVV_0
timestamp 1713185578
transform 1 0 1554 0 1 312
box -384 -180 384 180
use pmos_3p3_VRY6F7  pmos_3p3_VRY6F7_0
timestamp 1713185578
transform 1 0 1554 0 1 771
box -446 -242 446 242
<< labels >>
flabel psubdiffcont 1493 -3 1493 -3 0 FreeSans 750 0 0 0 VSS
flabel metal1 s 540 1042 540 1042 0 FreeSans 750 0 0 0 VDD
port 1 nsew
flabel metal1 s 2002 516 2002 516 0 FreeSans 750 0 0 0 OUT
port 2 nsew
flabel metal1 s 1097 125 1097 125 0 FreeSans 750 0 0 0 IN
port 3 nsew
flabel metal1 s 207 496 207 496 0 FreeSans 750 0 0 0 CLK
port 4 nsew
<< end >>
