** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/decoder_2x4_ibr.sch
**.subckt decoder_2x4_ibr IN2 IN1 VSS VDD D0 D1 D2 D3
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin D0
*.opin D1
*.opin D2
*.opin D3
x1 VSS IN1 IN1B VDD inv_my_ibr
x2 VSS IN2 IN2B VDD inv_my_ibr
x3 IN1B VSS VDD D0 IN2B and_2_ibr.
x4 IN1 VSS VDD D1 IN2B and_2_ibr.
x5 IN1B VSS VDD D2 IN2 and_2_ibr.
x6 IN1 VSS VDD D3 IN2 and_2_ibr.
**.ends

* expanding   symbol:  inv_my_ibr.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/inv_my_ibr.sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/inv_my_ibr.sch
.subckt inv_my_ibr VSS IN OUT VDD
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  and_2_ibr..sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/and_2_ibr..sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/and_2_ibr..sch
.subckt and_2_ibr. IN1 VSS VDD OUT IN2
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin OUT
x2 VSS net1 OUT VDD inv_my_ibr
x1 IN1 VSS VDD net1 IN2 NAND_dec_ibr
.ends


* expanding   symbol:  NAND_dec_ibr.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/NAND_dec_ibr.sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/NAND_dec_ibr.sch
.subckt NAND_dec_ibr IN1 VSS VDD OUT IN2
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin OUT
XM3 net1 IN2 VSS VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 OUT IN1 net1 VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 OUT IN1 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN2 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.end
