magic
tech gf180mcuC
magscale 1 10
timestamp 1694922630
<< nwell >>
rect -282 -1534 282 1534
<< pmos >>
rect -108 804 -52 1404
rect 52 804 108 1404
rect -108 68 -52 668
rect 52 68 108 668
rect -108 -668 -52 -68
rect 52 -668 108 -68
rect -108 -1404 -52 -804
rect 52 -1404 108 -804
<< pdiff >>
rect -196 1391 -108 1404
rect -196 817 -183 1391
rect -137 817 -108 1391
rect -196 804 -108 817
rect -52 1391 52 1404
rect -52 817 -23 1391
rect 23 817 52 1391
rect -52 804 52 817
rect 108 1391 196 1404
rect 108 817 137 1391
rect 183 817 196 1391
rect 108 804 196 817
rect -196 655 -108 668
rect -196 81 -183 655
rect -137 81 -108 655
rect -196 68 -108 81
rect -52 655 52 668
rect -52 81 -23 655
rect 23 81 52 655
rect -52 68 52 81
rect 108 655 196 668
rect 108 81 137 655
rect 183 81 196 655
rect 108 68 196 81
rect -196 -81 -108 -68
rect -196 -655 -183 -81
rect -137 -655 -108 -81
rect -196 -668 -108 -655
rect -52 -81 52 -68
rect -52 -655 -23 -81
rect 23 -655 52 -81
rect -52 -668 52 -655
rect 108 -81 196 -68
rect 108 -655 137 -81
rect 183 -655 196 -81
rect 108 -668 196 -655
rect -196 -817 -108 -804
rect -196 -1391 -183 -817
rect -137 -1391 -108 -817
rect -196 -1404 -108 -1391
rect -52 -817 52 -804
rect -52 -1391 -23 -817
rect 23 -1391 52 -817
rect -52 -1404 52 -1391
rect 108 -817 196 -804
rect 108 -1391 137 -817
rect 183 -1391 196 -817
rect 108 -1404 196 -1391
<< pdiffc >>
rect -183 817 -137 1391
rect -23 817 23 1391
rect 137 817 183 1391
rect -183 81 -137 655
rect -23 81 23 655
rect 137 81 183 655
rect -183 -655 -137 -81
rect -23 -655 23 -81
rect 137 -655 183 -81
rect -183 -1391 -137 -817
rect -23 -1391 23 -817
rect 137 -1391 183 -817
<< polysilicon >>
rect -108 1404 -52 1448
rect 52 1404 108 1448
rect -108 760 -52 804
rect 52 760 108 804
rect -108 668 -52 712
rect 52 668 108 712
rect -108 24 -52 68
rect 52 24 108 68
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect -108 -712 -52 -668
rect 52 -712 108 -668
rect -108 -804 -52 -760
rect 52 -804 108 -760
rect -108 -1448 -52 -1404
rect 52 -1448 108 -1404
<< metal1 >>
rect -183 1391 -137 1402
rect -183 806 -137 817
rect -23 1391 23 1402
rect -23 806 23 817
rect 137 1391 183 1402
rect 137 806 183 817
rect -183 655 -137 666
rect -183 70 -137 81
rect -23 655 23 666
rect -23 70 23 81
rect 137 655 183 666
rect 137 70 183 81
rect -183 -81 -137 -70
rect -183 -666 -137 -655
rect -23 -81 23 -70
rect -23 -666 23 -655
rect 137 -81 183 -70
rect 137 -666 183 -655
rect -183 -817 -137 -806
rect -183 -1402 -137 -1391
rect -23 -817 23 -806
rect -23 -1402 23 -1391
rect 137 -817 183 -806
rect 137 -1402 183 -1391
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 4 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
