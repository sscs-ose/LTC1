** sch_path: /home/shahid/GF180Projects/ahmar/5b_divider.sch
**.subckt 5b_divider VDD VSS CLK D2_1 D2_2 D2_3 D2_4 D2_5 LD Q5 Q4 Q2 Q3 Q1 OUT1 P2
*.iopin VDD
*.iopin VSS
*.ipin CLK
*.ipin D2_1
*.ipin D2_2
*.ipin D2_3
*.ipin D2_4
*.ipin D2_5
*.opin LD
*.opin Q5
*.opin Q4
*.opin Q2
*.opin Q3
*.opin Q1
*.opin OUT1
*.opin P2
x1 LD VDD Q4 Q2 Q3 Q1 Q5 D2_3 D2_5 D2_4 D2_2 D2_1 CLK VSS 5b_DC
x4 VDD Q2 b D2_3 VSS XNOR
x5 VDD Q1 a D2_2 VSS XNOR
x6 VDD Q3 c D2_4 VSS XNOR
x7 VDD net1 a b c VSS 3_inp_AND
x2 VDD Q4 d D2_5 VSS XNOR
x3 VDD Q5 e D2_1 VSS XNOR
x9 VDD net2 d e VSS NAND
x10 VDD net2 net3 VSS inverter
x11 VDD net4 net1 net3 VSS NAND
x12 VDD net4 net5 VSS inverter
x13 VDD P0 P2 net6 VSS OR
x14 net6 VDD OUT1 VSS div_by_2
x17 CLK VDD net5 P2 VSS DFF
x8 CLK VDD LD P0 VSS ned_DFF
x15 VDD Q2 c2 D2_3 VSS XNOR
x16 VDD Q1 c1 D2_2 VSS XNOR
x18 VDD Q3 c3 D2_4 VSS XNOR
x19 VDD Q4 c4 D2_5 VSS XNOR
x20 VDD Q5 c5 D2_1B VSS XNOR
x21 VDD D2_1 D2_1B VSS inverter
x22 VDD net7 c1 c2 c3 VSS 3_inp_AND
x23 VDD net8 c4 c5 VSS NAND
x24 VDD net8 net9 VSS inverter
x25 VDD net10 net7 net9 VSS NAND
x26 VDD net10 net11 VSS inverter
x27 CLK VDD net11 P3 VSS DFF
x28 CLK VDD P0 P1 VSS DFF
x29 VDD P1 P3 net12 VSS OR
x30 net12 VDD OUT2 VSS div_by_2
**.ends

* expanding   symbol:  5b_DC.sym # of pins=14
** sym_path: /home/shahid/GF180Projects/ahmar/5b_DC.sym
** sch_path: /home/shahid/GF180Projects/ahmar/5b_DC.sch
.subckt 5b_DC LD VDD Q4 Q2 Q3 Q1 Q5 D2_3 D2_5 D2_4 D2_2 D2_1 CLK VSS
*.iopin VDD
*.iopin VSS
*.opin Q3
*.opin Q1
*.ipin D2_1
*.ipin D2_2
*.ipin D2_3
*.ipin CLK
*.opin Q2
*.opin LD
*.ipin D2_4
*.opin Q4
*.ipin D2_5
*.opin Q5
x1 VDD LD D2_1 VSS CLK Q1 1 1 mod_DFF
x3 VDD LD D2_2 VSS Q1 Q2 2 2 mod_DFF
x4 VDD LD D2_3 VSS Q2 Q3 3 3 mod_DFF
x6 VDD net3 net2 net1 VSS NAND
x2 VDD LD D2_4 VSS Q3 Q4 4 4 mod_DFF
x5 VDD net6 net4 net5 VSS NAND
x11 VDD net6 net1 VSS inverter
x10 VDD LD D2_5 VSS Q4 Q5 5 5 mod_DFF
x12 VDD 1 2 net5 VSS NOR
x9 VDD 3 4 5 net4 VSS 3_inp_NOR
x7 CLK VDD net3 net2 VSS DFF
x8 VDD net2 LD VSS inverter
.ends


* expanding   symbol:  XNOR.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/ahmar/XNOR.sym
** sch_path: /home/shahid/GF180Projects/ahmar/XNOR.sch
.subckt XNOR VDD A OUT B VSS
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin OUT
XM1 OUT A net3 VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 A VDD VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net2 A_bar VDD VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 OUT B net1 VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 OUT B_bar net2 VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 OUT A_bar net4 VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 net3 B_bar VSS VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 net4 B VSS VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VDD A A_bar VSS inverter
x2 VDD B B_bar VSS inverter
.ends


* expanding   symbol:  3_inp_AND.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/ahmar/3_inp_AND.sym
** sch_path: /home/shahid/GF180Projects/ahmar/3_inp_AND.sch
.subckt 3_inp_AND VDD VOUT A B C VSS
*.iopin VSS
*.iopin VDD
*.ipin A
*.ipin B
*.ipin C
*.opin VOUT
XM1 net3 A net1 VSS nfet_03v3 L=0.28u W=1.32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net3 C VDD VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B net2 VSS nfet_03v3 L=0.28u W=1.32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net2 C VSS VSS nfet_03v3 L=0.28u W=1.32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net3 B VDD VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net3 A VDD VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VDD VOUT net3 VSS strong_inv
.ends


* expanding   symbol:  NAND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/ahmar/NAND.sym
** sch_path: /home/shahid/GF180Projects/ahmar/NAND.sch
.subckt NAND VDD VOUT A B VSS
*.iopin VDD
*.iopin VSS
*.ipin A
*.ipin B
*.opin VOUT
XM1 VOUT A net1 VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 VOUT A VDD VDD pfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 VOUT B VDD VDD pfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 B VSS VSS nfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/ahmar/inverter.sym
** sch_path: /home/shahid/GF180Projects/ahmar/inverter.sch
.subckt inverter VDD VIN VOUT VSS
*.iopin VDD
*.ipin VIN
*.opin VOUT
*.iopin VSS
XM4 VOUT VIN VDD VDD pfet_03v3 L=0.28u W=0.44u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VOUT VIN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  OR.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/ahmar/OR.sym
** sch_path: /home/shahid/GF180Projects/ahmar/OR.sch
.subckt OR VDD A B VOUT VSS
*.iopin VSS
*.iopin VDD
*.ipin A
*.ipin B
*.opin VOUT
XM1 net1 A VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 B net2 VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net2 A VDD VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
x1 VDD net1 VOUT VSS inverter
.ends


* expanding   symbol:  div_by_2.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/ahmar/div_by_2.sym
** sch_path: /home/shahid/GF180Projects/ahmar/div_by_2.sch
.subckt div_by_2 CLK VDD Q VSS
*.iopin VDD
*.iopin VSS
*.opin Q
*.ipin CLK
x1 VDD CLKB VSS net2 net1 tg
x3 VDD CLK VSS net2 net5 tg
x4 VDD CLK VSS net4 net3 tg
x5 VDD CLKB VSS net4 net1 tg
x2 VDD net2 net3 VSS inverter
x6 VDD net4 Q VSS inverter
x7 VDD Q net1 VSS inverter
x8 VDD net3 net5 VSS inverter
x9 VDD CLK CLKB VSS inverter
.ends


* expanding   symbol:  DFF.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/ahmar/DFF.sym
** sch_path: /home/shahid/GF180Projects/ahmar/DFF.sch
.subckt DFF CLK VDD D Q VSS
*.ipin D
*.iopin VDD
*.iopin VSS
*.opin Q
*.ipin CLK
x1 VDD CLKB VSS net1 D tg
x3 VDD CLK VSS net1 net5 tg
x4 VDD CLK VSS net3 net2 tg
x5 VDD CLKB VSS net3 net4 tg
x2 VDD net1 net2 VSS inverter
x6 VDD net3 Q VSS inverter
x7 VDD Q net4 VSS inverter
x8 VDD net2 net5 VSS inverter
x9 VDD CLK CLKB VSS inverter
.ends


* expanding   symbol:  ned_DFF.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/ahmar/ned_DFF.sym
** sch_path: /home/shahid/GF180Projects/ahmar/ned_DFF.sch
.subckt ned_DFF CLK VDD D Q VSS
*.ipin D
*.iopin VDD
*.iopin VSS
*.opin Q
*.ipin CLK
x1 VDD CLK VSS net1 D tg
x3 VDD CLKB VSS net1 net5 tg
x4 VDD CLKB VSS net3 net2 tg
x5 VDD CLK VSS net3 net4 tg
x2 VDD net1 net2 VSS inverter
x6 VDD net3 Q VSS inverter
x7 VDD Q net4 VSS inverter
x8 VDD net2 net5 VSS inverter
x9 VDD CLK CLKB VSS inverter
.ends


* expanding   symbol:  mod_DFF.sym # of pins=8
** sym_path: /home/shahid/GF180Projects/ahmar/mod_DFF.sym
** sch_path: /home/shahid/GF180Projects/ahmar/mod_DFF.sch
.subckt mod_DFF VDD LD D2 VSS CLK Q D1 Q-
*.ipin LD
*.ipin D2
*.iopin VDD
*.iopin VSS
*.ipin D1
*.opin Q
*.opin Q-
*.ipin CLK
x1 VDD net6 LD D2 VSS NAND
x2 VDD net5 LD net1 VSS NAND
x4 VDD CLKB VSS net2 D1 tg
x5 VDD net3 net2 net5 VSS NAND
x6 VDD CLK VSS net4 net3 tg
x7 VDD Q net4 net6 VSS NAND
x9 VDD Q Q- VSS inverter
x10 VDD net7 net5 Q VSS NAND
x11 VDD CLKB VSS net4 net7 tg
x12 VDD net8 net6 net3 VSS NAND
x13 VDD CLK VSS net2 net8 tg
x14 VDD D2 net1 VSS inverter
x15 VDD CLK CLKB VSS inverter
.ends


* expanding   symbol:  NOR.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/ahmar/NOR.sym
** sch_path: /home/shahid/GF180Projects/ahmar/NOR.sch
.subckt NOR VDD A B VOUT VSS
*.iopin VSS
*.iopin VDD
*.ipin A
*.ipin B
*.opin VOUT
XM1 VOUT A VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 VOUT B net1 VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 VOUT B VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net1 A VDD VDD pfet_03v3 L=0.28u W=0.88u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  3_inp_NOR.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/ahmar/3_inp_NOR.sym
** sch_path: /home/shahid/GF180Projects/ahmar/3_inp_NOR.sch
.subckt 3_inp_NOR VDD A B C VOUT VSS
*.iopin VSS
*.iopin VDD
*.ipin A
*.ipin B
*.ipin C
*.opin VOUT
XM1 VOUT A VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 B net2 VDD pfet_03v3 L=0.28u W=1.32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 VOUT B VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 VOUT C VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VOUT C net1 VDD pfet_03v3 L=0.28u W=1.32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net2 A VDD VDD pfet_03v3 L=0.28u W=1.32u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  strong_inv.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/ahmar/strong_inv.sym
** sch_path: /home/shahid/GF180Projects/ahmar/strong_inv.sch
.subckt strong_inv VDD VOUT VIN VSS
*.iopin VDD
*.ipin VIN
*.opin VOUT
*.iopin VSS
XM4 VOUT VIN VDD VDD pfet_03v3 L=2u W=4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 VOUT VIN VSS VSS nfet_03v3 L=2u W=2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  tg.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/ahmar/tg.sym
** sch_path: /home/shahid/GF180Projects/ahmar/tg.sch
.subckt tg VDD CLK VSS OUT IN
*.iopin VDD
*.iopin VSS
*.ipin CLK
*.ipin IN
*.opin OUT
x1 VDD CLK net1 VSS inverter
XM1 OUT net1 IN VDD pfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT CLK IN VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.end
