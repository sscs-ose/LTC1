magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2092 -4342 2092 4342
<< polysilicon >>
rect -92 2279 92 2342
rect -92 -2279 -70 2279
rect 70 -2279 92 2279
rect -92 -2342 92 -2279
<< polycontact >>
rect -70 -2279 70 2279
<< metal1 >>
rect -84 2279 84 2334
rect -84 -2279 -70 2279
rect 70 -2279 84 2279
rect -84 -2334 84 -2279
<< end >>
