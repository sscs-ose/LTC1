magic
tech gf180mcuC
magscale 1 10
timestamp 1691411081
<< pwell >>
rect -336 -558 336 558
<< psubdiff >>
rect -312 462 312 534
rect -312 -462 -240 462
rect 240 -462 312 462
rect -312 -534 312 -462
<< polysilicon >>
rect -100 309 100 322
rect -100 263 -87 309
rect 87 263 100 309
rect -100 200 100 263
rect -100 -263 100 -200
rect -100 -309 -87 -263
rect 87 -309 100 -263
rect -100 -322 100 -309
<< polycontact >>
rect -87 263 87 309
rect -87 -309 87 -263
<< nhighres >>
rect -100 -200 100 200
<< metal1 >>
rect -98 263 -87 309
rect 87 263 98 309
rect -98 -309 -87 -263
rect 87 -309 98 -263
<< properties >>
string FIXED_BBOX -276 -498 276 498
string gencell ppolyf_u_1k
string library gf180mcu
string parameters w 1.0 l 2.0 m 1 nx 1 wmin 1.000 lmin 1.000 rho 1000 val 2.0k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0 compatible {ppolyf_u_1k ppolyf_u_1k_6p0}
<< end >>
