magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2083 -2083 4889 4911
<< isosubstrate >>
rect 1197 -83 2889 2911
<< nwell >>
rect -83 1213 857 2911
rect 1197 1213 2889 2911
<< polysilicon >>
rect 317 698 457 1578
rect 1605 1202 1745 1914
rect 1849 1202 1989 1914
rect 1605 991 1989 1202
rect 1605 698 1745 991
rect 1849 698 1989 991
rect 2093 1202 2233 1914
rect 2337 1202 2477 1914
rect 2093 991 2477 1202
rect 2093 698 2233 991
rect 2337 698 2477 991
<< metal1 >>
rect 79 2749 165 2817
rect 227 1622 303 2800
rect 609 2749 695 2817
rect 1359 2749 1445 2817
rect 471 1186 547 2222
rect 1515 1622 1591 2812
rect 1759 1186 1835 2222
rect 2003 1622 2079 2812
rect 471 1008 1699 1186
rect 1759 1008 2187 1186
rect 79 11 165 79
rect 227 42 303 654
rect 471 354 547 1008
rect 609 11 695 79
rect 1359 11 1445 79
rect 1515 39 1591 654
rect 1759 354 1835 1008
rect 2003 39 2079 654
rect 2247 354 2323 2222
rect 2491 1622 2567 2812
rect 2641 2749 2727 2817
rect 2491 39 2567 654
rect 2641 11 2727 79
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_0
timestamp 1713338890
transform 1 0 45 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_1
timestamp 1713338890
transform 1 0 729 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_2
timestamp 1713338890
transform 1 0 1325 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_3
timestamp 1713338890
transform 1 0 2761 0 1 2078
box -128 -833 128 833
use M1_NWELL_CDNS_40661953145273  M1_NWELL_CDNS_40661953145273_0
timestamp 1713338890
transform 1 0 387 0 1 2783
box -316 -128 316 128
use M1_NWELL_CDNS_40661953145274  M1_NWELL_CDNS_40661953145274_0
timestamp 1713338890
transform 1 0 2043 0 1 2783
box -692 -128 692 128
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_0
timestamp 1713338890
transform 1 0 377 0 1 1097
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_1
timestamp 1713338890
transform 1 0 1665 0 1 1097
box -42 -89 42 89
use M1_POLY2_CDNS_69033583165610  M1_POLY2_CDNS_69033583165610_2
timestamp 1713338890
transform 1 0 2153 0 1 1097
box -42 -89 42 89
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_0
timestamp 1713338890
transform 1 0 45 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165609  M1_PSUB_CDNS_69033583165609_1
timestamp 1713338890
transform 1 0 2761 0 -1 515
box -45 -515 45 515
use M1_PSUB_CDNS_69033583165611  M1_PSUB_CDNS_69033583165611_0
timestamp 1713338890
transform 1 0 729 0 -1 468
box -45 -468 45 468
use M1_PSUB_CDNS_69033583165611  M1_PSUB_CDNS_69033583165611_1
timestamp 1713338890
transform 1 0 1325 0 -1 468
box -45 -468 45 468
use M1_PSUB_CDNS_69033583165621  M1_PSUB_CDNS_69033583165621_0
timestamp 1713338890
transform 1 0 387 0 -1 45
box -233 -45 233 45
use M1_PSUB_CDNS_69033583165695  M1_PSUB_CDNS_69033583165695_0
timestamp 1713338890
transform 1 0 2043 0 -1 45
box -609 -45 609 45
use nmos_6p0_CDNS_4066195314530  nmos_6p0_CDNS_4066195314530_0
timestamp 1713338890
transform 1 0 317 0 1 354
box -88 -44 228 344
use nmos_6p0_CDNS_4066195314531  nmos_6p0_CDNS_4066195314531_0
timestamp 1713338890
transform 1 0 1605 0 1 354
box -88 -44 472 344
use nmos_6p0_CDNS_4066195314531  nmos_6p0_CDNS_4066195314531_1
timestamp 1713338890
transform 1 0 2093 0 1 354
box -88 -44 472 344
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1713338890
transform 1 0 317 0 1 1622
box -208 -120 348 720
use pmos_6p0_CDNS_4066195314529  pmos_6p0_CDNS_4066195314529_0
timestamp 1713338890
transform 1 0 1605 0 1 1622
box -208 -120 592 720
use pmos_6p0_CDNS_4066195314529  pmos_6p0_CDNS_4066195314529_1
timestamp 1713338890
transform 1 0 2093 0 1 1622
box -208 -120 592 720
<< labels >>
rlabel metal1 s 2286 1098 2286 1098 4 ZB
port 1 nsew
rlabel metal1 s 350 2788 350 2788 4 VDD
port 2 nsew
rlabel metal1 s 377 1098 377 1098 4 A
port 3 nsew
rlabel metal1 s 2442 2788 2442 2788 4 DVDD
port 4 nsew
rlabel metal1 s 2433 45 2433 45 4 DVSS
port 5 nsew
rlabel metal1 s 263 45 263 45 4 VSS
port 6 nsew
rlabel metal1 s 2031 1098 2031 1098 4 Z
port 7 nsew
<< end >>
