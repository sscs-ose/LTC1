magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1331 1019 1331
<< metal1 >>
rect -19 325 19 331
rect -19 -325 -13 325
rect 13 -325 19 325
rect -19 -331 19 -325
<< via1 >>
rect -13 -325 13 325
<< metal2 >>
rect -19 325 19 331
rect -19 -325 -13 325
rect 13 -325 19 325
rect -19 -331 19 -325
<< end >>
