magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1856 1019 1856
<< metal2 >>
rect -19 851 19 856
rect -19 823 -14 851
rect 14 823 19 851
rect -19 789 19 823
rect -19 761 -14 789
rect 14 761 19 789
rect -19 727 19 761
rect -19 699 -14 727
rect 14 699 19 727
rect -19 665 19 699
rect -19 637 -14 665
rect 14 637 19 665
rect -19 603 19 637
rect -19 575 -14 603
rect 14 575 19 603
rect -19 541 19 575
rect -19 513 -14 541
rect 14 513 19 541
rect -19 479 19 513
rect -19 451 -14 479
rect 14 451 19 479
rect -19 417 19 451
rect -19 389 -14 417
rect 14 389 19 417
rect -19 355 19 389
rect -19 327 -14 355
rect 14 327 19 355
rect -19 293 19 327
rect -19 265 -14 293
rect 14 265 19 293
rect -19 231 19 265
rect -19 203 -14 231
rect 14 203 19 231
rect -19 169 19 203
rect -19 141 -14 169
rect 14 141 19 169
rect -19 107 19 141
rect -19 79 -14 107
rect 14 79 19 107
rect -19 45 19 79
rect -19 17 -14 45
rect 14 17 19 45
rect -19 -17 19 17
rect -19 -45 -14 -17
rect 14 -45 19 -17
rect -19 -79 19 -45
rect -19 -107 -14 -79
rect 14 -107 19 -79
rect -19 -141 19 -107
rect -19 -169 -14 -141
rect 14 -169 19 -141
rect -19 -203 19 -169
rect -19 -231 -14 -203
rect 14 -231 19 -203
rect -19 -265 19 -231
rect -19 -293 -14 -265
rect 14 -293 19 -265
rect -19 -327 19 -293
rect -19 -355 -14 -327
rect 14 -355 19 -327
rect -19 -389 19 -355
rect -19 -417 -14 -389
rect 14 -417 19 -389
rect -19 -451 19 -417
rect -19 -479 -14 -451
rect 14 -479 19 -451
rect -19 -513 19 -479
rect -19 -541 -14 -513
rect 14 -541 19 -513
rect -19 -575 19 -541
rect -19 -603 -14 -575
rect 14 -603 19 -575
rect -19 -637 19 -603
rect -19 -665 -14 -637
rect 14 -665 19 -637
rect -19 -699 19 -665
rect -19 -727 -14 -699
rect 14 -727 19 -699
rect -19 -761 19 -727
rect -19 -789 -14 -761
rect 14 -789 19 -761
rect -19 -823 19 -789
rect -19 -851 -14 -823
rect 14 -851 19 -823
rect -19 -856 19 -851
<< via2 >>
rect -14 823 14 851
rect -14 761 14 789
rect -14 699 14 727
rect -14 637 14 665
rect -14 575 14 603
rect -14 513 14 541
rect -14 451 14 479
rect -14 389 14 417
rect -14 327 14 355
rect -14 265 14 293
rect -14 203 14 231
rect -14 141 14 169
rect -14 79 14 107
rect -14 17 14 45
rect -14 -45 14 -17
rect -14 -107 14 -79
rect -14 -169 14 -141
rect -14 -231 14 -203
rect -14 -293 14 -265
rect -14 -355 14 -327
rect -14 -417 14 -389
rect -14 -479 14 -451
rect -14 -541 14 -513
rect -14 -603 14 -575
rect -14 -665 14 -637
rect -14 -727 14 -699
rect -14 -789 14 -761
rect -14 -851 14 -823
<< metal3 >>
rect -19 851 19 856
rect -19 823 -14 851
rect 14 823 19 851
rect -19 789 19 823
rect -19 761 -14 789
rect 14 761 19 789
rect -19 727 19 761
rect -19 699 -14 727
rect 14 699 19 727
rect -19 665 19 699
rect -19 637 -14 665
rect 14 637 19 665
rect -19 603 19 637
rect -19 575 -14 603
rect 14 575 19 603
rect -19 541 19 575
rect -19 513 -14 541
rect 14 513 19 541
rect -19 479 19 513
rect -19 451 -14 479
rect 14 451 19 479
rect -19 417 19 451
rect -19 389 -14 417
rect 14 389 19 417
rect -19 355 19 389
rect -19 327 -14 355
rect 14 327 19 355
rect -19 293 19 327
rect -19 265 -14 293
rect 14 265 19 293
rect -19 231 19 265
rect -19 203 -14 231
rect 14 203 19 231
rect -19 169 19 203
rect -19 141 -14 169
rect 14 141 19 169
rect -19 107 19 141
rect -19 79 -14 107
rect 14 79 19 107
rect -19 45 19 79
rect -19 17 -14 45
rect 14 17 19 45
rect -19 -17 19 17
rect -19 -45 -14 -17
rect 14 -45 19 -17
rect -19 -79 19 -45
rect -19 -107 -14 -79
rect 14 -107 19 -79
rect -19 -141 19 -107
rect -19 -169 -14 -141
rect 14 -169 19 -141
rect -19 -203 19 -169
rect -19 -231 -14 -203
rect 14 -231 19 -203
rect -19 -265 19 -231
rect -19 -293 -14 -265
rect 14 -293 19 -265
rect -19 -327 19 -293
rect -19 -355 -14 -327
rect 14 -355 19 -327
rect -19 -389 19 -355
rect -19 -417 -14 -389
rect 14 -417 19 -389
rect -19 -451 19 -417
rect -19 -479 -14 -451
rect 14 -479 19 -451
rect -19 -513 19 -479
rect -19 -541 -14 -513
rect 14 -541 19 -513
rect -19 -575 19 -541
rect -19 -603 -14 -575
rect 14 -603 19 -575
rect -19 -637 19 -603
rect -19 -665 -14 -637
rect 14 -665 19 -637
rect -19 -699 19 -665
rect -19 -727 -14 -699
rect 14 -727 19 -699
rect -19 -761 19 -727
rect -19 -789 -14 -761
rect 14 -789 19 -761
rect -19 -823 19 -789
rect -19 -851 -14 -823
rect 14 -851 19 -823
rect -19 -856 19 -851
<< end >>
