magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2109 -3458 2109 3458
<< metal2 >>
rect -109 1448 109 1458
rect -109 1392 -99 1448
rect -43 1392 43 1448
rect 99 1392 109 1448
rect -109 1306 109 1392
rect -109 1250 -99 1306
rect -43 1250 43 1306
rect 99 1250 109 1306
rect -109 1164 109 1250
rect -109 1108 -99 1164
rect -43 1108 43 1164
rect 99 1108 109 1164
rect -109 1022 109 1108
rect -109 966 -99 1022
rect -43 966 43 1022
rect 99 966 109 1022
rect -109 880 109 966
rect -109 824 -99 880
rect -43 824 43 880
rect 99 824 109 880
rect -109 738 109 824
rect -109 682 -99 738
rect -43 682 43 738
rect 99 682 109 738
rect -109 596 109 682
rect -109 540 -99 596
rect -43 540 43 596
rect 99 540 109 596
rect -109 454 109 540
rect -109 398 -99 454
rect -43 398 43 454
rect 99 398 109 454
rect -109 312 109 398
rect -109 256 -99 312
rect -43 256 43 312
rect 99 256 109 312
rect -109 170 109 256
rect -109 114 -99 170
rect -43 114 43 170
rect 99 114 109 170
rect -109 28 109 114
rect -109 -28 -99 28
rect -43 -28 43 28
rect 99 -28 109 28
rect -109 -114 109 -28
rect -109 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 109 -114
rect -109 -256 109 -170
rect -109 -312 -99 -256
rect -43 -312 43 -256
rect 99 -312 109 -256
rect -109 -398 109 -312
rect -109 -454 -99 -398
rect -43 -454 43 -398
rect 99 -454 109 -398
rect -109 -540 109 -454
rect -109 -596 -99 -540
rect -43 -596 43 -540
rect 99 -596 109 -540
rect -109 -682 109 -596
rect -109 -738 -99 -682
rect -43 -738 43 -682
rect 99 -738 109 -682
rect -109 -824 109 -738
rect -109 -880 -99 -824
rect -43 -880 43 -824
rect 99 -880 109 -824
rect -109 -966 109 -880
rect -109 -1022 -99 -966
rect -43 -1022 43 -966
rect 99 -1022 109 -966
rect -109 -1108 109 -1022
rect -109 -1164 -99 -1108
rect -43 -1164 43 -1108
rect 99 -1164 109 -1108
rect -109 -1250 109 -1164
rect -109 -1306 -99 -1250
rect -43 -1306 43 -1250
rect 99 -1306 109 -1250
rect -109 -1392 109 -1306
rect -109 -1448 -99 -1392
rect -43 -1448 43 -1392
rect 99 -1448 109 -1392
rect -109 -1458 109 -1448
<< via2 >>
rect -99 1392 -43 1448
rect 43 1392 99 1448
rect -99 1250 -43 1306
rect 43 1250 99 1306
rect -99 1108 -43 1164
rect 43 1108 99 1164
rect -99 966 -43 1022
rect 43 966 99 1022
rect -99 824 -43 880
rect 43 824 99 880
rect -99 682 -43 738
rect 43 682 99 738
rect -99 540 -43 596
rect 43 540 99 596
rect -99 398 -43 454
rect 43 398 99 454
rect -99 256 -43 312
rect 43 256 99 312
rect -99 114 -43 170
rect 43 114 99 170
rect -99 -28 -43 28
rect 43 -28 99 28
rect -99 -170 -43 -114
rect 43 -170 99 -114
rect -99 -312 -43 -256
rect 43 -312 99 -256
rect -99 -454 -43 -398
rect 43 -454 99 -398
rect -99 -596 -43 -540
rect 43 -596 99 -540
rect -99 -738 -43 -682
rect 43 -738 99 -682
rect -99 -880 -43 -824
rect 43 -880 99 -824
rect -99 -1022 -43 -966
rect 43 -1022 99 -966
rect -99 -1164 -43 -1108
rect 43 -1164 99 -1108
rect -99 -1306 -43 -1250
rect 43 -1306 99 -1250
rect -99 -1448 -43 -1392
rect 43 -1448 99 -1392
<< metal3 >>
rect -109 1448 109 1458
rect -109 1392 -99 1448
rect -43 1392 43 1448
rect 99 1392 109 1448
rect -109 1306 109 1392
rect -109 1250 -99 1306
rect -43 1250 43 1306
rect 99 1250 109 1306
rect -109 1164 109 1250
rect -109 1108 -99 1164
rect -43 1108 43 1164
rect 99 1108 109 1164
rect -109 1022 109 1108
rect -109 966 -99 1022
rect -43 966 43 1022
rect 99 966 109 1022
rect -109 880 109 966
rect -109 824 -99 880
rect -43 824 43 880
rect 99 824 109 880
rect -109 738 109 824
rect -109 682 -99 738
rect -43 682 43 738
rect 99 682 109 738
rect -109 596 109 682
rect -109 540 -99 596
rect -43 540 43 596
rect 99 540 109 596
rect -109 454 109 540
rect -109 398 -99 454
rect -43 398 43 454
rect 99 398 109 454
rect -109 312 109 398
rect -109 256 -99 312
rect -43 256 43 312
rect 99 256 109 312
rect -109 170 109 256
rect -109 114 -99 170
rect -43 114 43 170
rect 99 114 109 170
rect -109 28 109 114
rect -109 -28 -99 28
rect -43 -28 43 28
rect 99 -28 109 28
rect -109 -114 109 -28
rect -109 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 109 -114
rect -109 -256 109 -170
rect -109 -312 -99 -256
rect -43 -312 43 -256
rect 99 -312 109 -256
rect -109 -398 109 -312
rect -109 -454 -99 -398
rect -43 -454 43 -398
rect 99 -454 109 -398
rect -109 -540 109 -454
rect -109 -596 -99 -540
rect -43 -596 43 -540
rect 99 -596 109 -540
rect -109 -682 109 -596
rect -109 -738 -99 -682
rect -43 -738 43 -682
rect 99 -738 109 -682
rect -109 -824 109 -738
rect -109 -880 -99 -824
rect -43 -880 43 -824
rect 99 -880 109 -824
rect -109 -966 109 -880
rect -109 -1022 -99 -966
rect -43 -1022 43 -966
rect 99 -1022 109 -966
rect -109 -1108 109 -1022
rect -109 -1164 -99 -1108
rect -43 -1164 43 -1108
rect 99 -1164 109 -1108
rect -109 -1250 109 -1164
rect -109 -1306 -99 -1250
rect -43 -1306 43 -1250
rect 99 -1306 109 -1250
rect -109 -1392 109 -1306
rect -109 -1448 -99 -1392
rect -43 -1448 43 -1392
rect 99 -1448 109 -1392
rect -109 -1458 109 -1448
<< end >>
