magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2051 -2051 15013 27617
<< polysilicon >>
rect 1237 23733 1437 23873
rect 11525 23733 11725 23873
rect 1421 23489 1437 23629
rect 11525 23489 11541 23629
rect 1421 23245 1437 23385
rect 11525 23245 11541 23385
rect 1421 23001 1437 23141
rect 11525 23001 11541 23141
rect 1421 22757 1437 22897
rect 11525 22757 11541 22897
rect 1421 22513 1437 22653
rect 11525 22513 11541 22653
rect 1421 22269 1437 22409
rect 11525 22269 11541 22409
rect 1421 22025 1437 22165
rect 11525 22025 11541 22165
rect 1421 21781 1437 21921
rect 11525 21781 11541 21921
rect 1421 21537 1437 21677
rect 11525 21537 11541 21677
rect 1421 21293 1437 21433
rect 11525 21293 11541 21433
rect 1421 21049 1437 21189
rect 11525 21049 11541 21189
rect 1421 20805 1437 20945
rect 11525 20805 11541 20945
rect 1421 20561 1437 20701
rect 11525 20561 11541 20701
rect 1421 20317 1437 20457
rect 11525 20317 11541 20457
rect 1421 20073 1437 20213
rect 11525 20073 11541 20213
rect 1421 19829 1437 19969
rect 11525 19829 11541 19969
rect 1421 19585 1437 19725
rect 11525 19585 11541 19725
rect 1421 19341 1437 19481
rect 11525 19341 11541 19481
rect 1237 19097 1437 19237
rect 11525 19097 11725 19237
rect 1237 17861 1437 18001
rect 11525 17861 11725 18001
rect 1421 17617 1437 17757
rect 11525 17617 11541 17757
rect 1421 17373 1437 17513
rect 11525 17373 11541 17513
rect 1421 17129 1437 17269
rect 11525 17129 11541 17269
rect 1421 16885 1437 17025
rect 11525 16885 11541 17025
rect 1421 16641 1437 16781
rect 11525 16641 11541 16781
rect 1421 16397 1437 16537
rect 11525 16397 11541 16537
rect 1421 16153 1437 16293
rect 11525 16153 11541 16293
rect 1421 15909 1437 16049
rect 11525 15909 11541 16049
rect 1421 15665 1437 15805
rect 11525 15665 11541 15805
rect 1421 15421 1437 15561
rect 11525 15421 11541 15561
rect 1421 15177 1437 15317
rect 11525 15177 11541 15317
rect 1421 14933 1437 15073
rect 11525 14933 11541 15073
rect 1421 14689 1437 14829
rect 11525 14689 11541 14829
rect 1421 14445 1437 14585
rect 11525 14445 11541 14585
rect 1421 14201 1437 14341
rect 11525 14201 11541 14341
rect 1421 13957 1437 14097
rect 11525 13957 11541 14097
rect 1421 13713 1437 13853
rect 11525 13713 11541 13853
rect 1421 13469 1437 13609
rect 11525 13469 11541 13609
rect 1237 13225 1437 13365
rect 11525 13225 11725 13365
rect 1237 11989 1437 12129
rect 11525 11989 11725 12129
rect 1421 11745 1437 11885
rect 11525 11745 11541 11885
rect 1421 11501 1437 11641
rect 11525 11501 11541 11641
rect 1421 11257 1437 11397
rect 11525 11257 11541 11397
rect 1421 11013 1437 11153
rect 11525 11013 11541 11153
rect 1421 10769 1437 10909
rect 11525 10769 11541 10909
rect 1421 10525 1437 10665
rect 11525 10525 11541 10665
rect 1421 10281 1437 10421
rect 11525 10281 11541 10421
rect 1421 10037 1437 10177
rect 11525 10037 11541 10177
rect 1421 9793 1437 9933
rect 11525 9793 11541 9933
rect 1421 9549 1437 9689
rect 11525 9549 11541 9689
rect 1421 9305 1437 9445
rect 11525 9305 11541 9445
rect 1421 9061 1437 9201
rect 11525 9061 11541 9201
rect 1421 8817 1437 8957
rect 11525 8817 11541 8957
rect 1421 8573 1437 8713
rect 11525 8573 11541 8713
rect 1421 8329 1437 8469
rect 11525 8329 11541 8469
rect 1421 8085 1437 8225
rect 11525 8085 11541 8225
rect 1421 7841 1437 7981
rect 11525 7841 11541 7981
rect 1421 7597 1437 7737
rect 11525 7597 11541 7737
rect 1237 7353 1437 7493
rect 11525 7353 11725 7493
rect 1237 6117 1437 6257
rect 11525 6117 11725 6257
rect 1421 5873 1437 6013
rect 11525 5873 11541 6013
rect 1421 5629 1437 5769
rect 11525 5629 11541 5769
rect 1421 5385 1437 5525
rect 11525 5385 11541 5525
rect 1421 5141 1437 5281
rect 11525 5141 11541 5281
rect 1421 4897 1437 5037
rect 11525 4897 11541 5037
rect 1421 4653 1437 4793
rect 11525 4653 11541 4793
rect 1421 4409 1437 4549
rect 11525 4409 11541 4549
rect 1421 4165 1437 4305
rect 11525 4165 11541 4305
rect 1421 3921 1437 4061
rect 11525 3921 11541 4061
rect 1421 3677 1437 3817
rect 11525 3677 11541 3817
rect 1421 3433 1437 3573
rect 11525 3433 11541 3573
rect 1421 3189 1437 3329
rect 11525 3189 11541 3329
rect 1421 2945 1437 3085
rect 11525 2945 11541 3085
rect 1421 2701 1437 2841
rect 11525 2701 11541 2841
rect 1421 2457 1437 2597
rect 11525 2457 11541 2597
rect 1421 2213 1437 2353
rect 11525 2213 11541 2353
rect 1421 1969 1437 2109
rect 11525 1969 11541 2109
rect 1421 1725 1437 1865
rect 11525 1725 11541 1865
rect 1237 1481 1437 1621
rect 11525 1481 11725 1621
<< metal1 >>
rect 411 24943 497 25311
rect 12465 24943 12551 25311
rect 961 24343 1047 24711
rect 11915 24343 12001 24711
rect 1213 24053 11749 24253
rect 1213 18920 1413 24053
rect 1481 23887 11481 23963
rect 1481 23643 11481 23719
rect 1481 23399 11481 23475
rect 1481 23155 11481 23231
rect 1481 22911 11481 22987
rect 1481 22667 11481 22743
rect 1481 22423 11481 22499
rect 1481 22179 11481 22255
rect 1481 21935 11481 22011
rect 1481 21691 11481 21767
rect 1481 21447 11481 21523
rect 1481 21203 11481 21279
rect 1481 20959 11481 21035
rect 1481 20715 11481 20791
rect 1481 20471 11481 20547
rect 1481 20227 11481 20303
rect 1481 19983 11481 20059
rect 1481 19739 11481 19815
rect 1481 19495 11481 19571
rect 1481 19251 11481 19327
rect 1481 19007 11481 19083
rect 11549 18920 11749 24053
rect 1213 18720 11749 18920
rect 961 18457 12001 18641
rect 1213 18178 11749 18378
rect 1213 13048 1413 18178
rect 1481 18015 11481 18091
rect 1481 17771 11481 17847
rect 1481 17527 11481 17603
rect 1481 17283 11481 17359
rect 1481 17039 11481 17115
rect 1481 16795 11481 16871
rect 1481 16551 11481 16627
rect 1481 16307 11481 16383
rect 1481 16063 11481 16139
rect 1481 15819 11481 15895
rect 1481 15575 11481 15651
rect 1481 15331 11481 15407
rect 1481 15087 11481 15163
rect 1481 14843 11481 14919
rect 1481 14599 11481 14675
rect 1481 14355 11481 14431
rect 1481 14111 11481 14187
rect 1481 13867 11481 13943
rect 1481 13623 11481 13699
rect 1481 13379 11481 13455
rect 1481 13135 11481 13211
rect 11549 13048 11749 18178
rect 1213 12848 11749 13048
rect 961 12585 12001 12769
rect 1213 12306 11749 12506
rect 1213 7176 1413 12306
rect 1481 12143 11481 12219
rect 1481 11899 11481 11975
rect 1481 11655 11481 11731
rect 1481 11411 11481 11487
rect 1481 11167 11481 11243
rect 1481 10923 11481 10999
rect 1481 10679 11481 10755
rect 1481 10435 11481 10511
rect 1481 10191 11481 10267
rect 1481 9947 11481 10023
rect 1481 9703 11481 9779
rect 1481 9459 11481 9535
rect 1481 9215 11481 9291
rect 1481 8971 11481 9047
rect 1481 8727 11481 8803
rect 1481 8483 11481 8559
rect 1481 8239 11481 8315
rect 1481 7995 11481 8071
rect 1481 7751 11481 7827
rect 1481 7507 11481 7583
rect 1481 7263 11481 7339
rect 11549 7176 11749 12306
rect 1213 6976 11749 7176
rect 961 6713 12001 6897
rect 1213 6434 11749 6634
rect 1213 1298 1413 6434
rect 1481 6271 11481 6347
rect 1481 6027 11481 6103
rect 1481 5783 11481 5859
rect 1481 5539 11481 5615
rect 1481 5295 11481 5371
rect 1481 5051 11481 5127
rect 1481 4807 11481 4883
rect 1481 4563 11481 4639
rect 1481 4319 11481 4395
rect 1481 4075 11481 4151
rect 1481 3831 11481 3907
rect 1481 3587 11481 3663
rect 1481 3343 11481 3419
rect 1481 3099 11481 3175
rect 1481 2855 11481 2931
rect 1481 2611 11481 2687
rect 1481 2367 11481 2443
rect 1481 2123 11481 2199
rect 1481 1879 11481 1955
rect 1481 1635 11481 1711
rect 1481 1391 11481 1467
rect 11549 1298 11749 6434
rect 1213 1098 11749 1298
rect 961 643 1047 1011
rect 11915 643 12001 1011
rect 411 43 497 411
rect 12465 43 12551 411
<< metal2 >>
rect 43 43 1145 25617
rect 1213 1455 1413 25617
rect 1481 43 3309 25617
rect 3409 43 5237 25617
rect 5337 43 6431 25617
rect 6531 43 7625 25617
rect 7725 43 9553 25617
rect 9653 43 11481 25617
rect 11549 1455 11749 25617
rect 11817 43 12919 25617
use M1_NWELL_CDNS_40661953145131  M1_NWELL_CDNS_40661953145131_0
timestamp 1713338890
transform 1 0 12735 0 1 12677
box -278 -12728 278 12728
use M1_NWELL_CDNS_40661953145131  M1_NWELL_CDNS_40661953145131_1
timestamp 1713338890
transform 1 0 227 0 1 12677
box -278 -12728 278 12728
use M1_NWELL_CDNS_40661953145135  M1_NWELL_CDNS_40661953145135_0
timestamp 1713338890
transform 1 0 6481 0 1 227
box -6078 -278 6078 278
use M1_NWELL_CDNS_40661953145135  M1_NWELL_CDNS_40661953145135_1
timestamp 1713338890
transform 1 0 6481 0 1 25127
box -6078 -278 6078 278
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_0
timestamp 1713338890
transform 1 0 1329 0 1 3869
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_1
timestamp 1713338890
transform -1 0 11633 0 1 3869
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_2
timestamp 1713338890
transform 1 0 1329 0 1 9741
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_3
timestamp 1713338890
transform -1 0 11633 0 1 9741
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_4
timestamp 1713338890
transform 1 0 1329 0 1 15613
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_5
timestamp 1713338890
transform -1 0 11633 0 1 15613
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_6
timestamp 1713338890
transform 1 0 1329 0 1 21485
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_7
timestamp 1713338890
transform -1 0 11633 0 1 21485
box -92 -2342 92 2342
use M1_PSUB_CDNS_69033583165354  M1_PSUB_CDNS_69033583165354_0
timestamp 1713338890
transform 1 0 6481 0 1 827
box -5445 -195 5445 195
use M1_PSUB_CDNS_69033583165354  M1_PSUB_CDNS_69033583165354_1
timestamp 1713338890
transform 1 0 6481 0 1 24527
box -5445 -195 5445 195
use M1_PSUB_CDNS_69033583165355  M1_PSUB_CDNS_69033583165355_0
timestamp 1713338890
transform 1 0 777 0 1 12677
box -195 -12045 195 12045
use M1_PSUB_CDNS_69033583165355  M1_PSUB_CDNS_69033583165355_1
timestamp 1713338890
transform 1 0 12185 0 1 12677
box -195 -12045 195 12045
use M1_PSUB_CDNS_69033583165356  M1_PSUB_CDNS_69033583165356_0
timestamp 1713338890
transform 1 0 6481 0 1 6805
box -5445 -95 5445 95
use M1_PSUB_CDNS_69033583165356  M1_PSUB_CDNS_69033583165356_1
timestamp 1713338890
transform 1 0 6481 0 1 12677
box -5445 -95 5445 95
use M1_PSUB_CDNS_69033583165356  M1_PSUB_CDNS_69033583165356_2
timestamp 1713338890
transform 1 0 6481 0 1 18549
box -5445 -95 5445 95
use M2_M1_CDNS_69033583165352  M2_M1_CDNS_69033583165352_0
timestamp 1713338890
transform 1 0 5884 0 1 6805
box -524 -92 524 92
use M2_M1_CDNS_69033583165352  M2_M1_CDNS_69033583165352_1
timestamp 1713338890
transform 1 0 5884 0 1 12677
box -524 -92 524 92
use M2_M1_CDNS_69033583165352  M2_M1_CDNS_69033583165352_2
timestamp 1713338890
transform 1 0 5884 0 1 18549
box -524 -92 524 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_0
timestamp 1713338890
transform 1 0 2395 0 1 6805
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_1
timestamp 1713338890
transform 1 0 8639 0 1 6805
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_2
timestamp 1713338890
transform 1 0 8639 0 1 12677
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_3
timestamp 1713338890
transform 1 0 2395 0 1 12677
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_4
timestamp 1713338890
transform 1 0 2395 0 1 18549
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_5
timestamp 1713338890
transform 1 0 8639 0 1 18549
box -902 -92 902 92
use M2_M1_CDNS_69033583165357  M2_M1_CDNS_69033583165357_0
timestamp 1713338890
transform 1 0 227 0 1 12677
box -146 -12188 146 12188
use M2_M1_CDNS_69033583165358  M2_M1_CDNS_69033583165358_0
timestamp 1713338890
transform 1 0 12185 0 1 12677
box -146 -11972 146 11972
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_0
timestamp 1713338890
transform 1 0 2395 0 1 1673
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_1
timestamp 1713338890
transform 1 0 2395 0 1 2161
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_2
timestamp 1713338890
transform 1 0 2395 0 1 2649
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_3
timestamp 1713338890
transform 1 0 2395 0 1 3137
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_4
timestamp 1713338890
transform 1 0 2395 0 1 3625
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_5
timestamp 1713338890
transform 1 0 2395 0 1 4113
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_6
timestamp 1713338890
transform 1 0 2395 0 1 4601
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_7
timestamp 1713338890
transform 1 0 4323 0 1 1917
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_8
timestamp 1713338890
transform 1 0 4323 0 1 1429
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_9
timestamp 1713338890
transform 1 0 4323 0 1 2405
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_10
timestamp 1713338890
transform 1 0 4323 0 1 2893
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_11
timestamp 1713338890
transform 1 0 4323 0 1 3381
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_12
timestamp 1713338890
transform 1 0 4323 0 1 3869
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_13
timestamp 1713338890
transform 1 0 4323 0 1 4357
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_14
timestamp 1713338890
transform 1 0 4323 0 1 4845
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_15
timestamp 1713338890
transform 1 0 8639 0 1 1673
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_16
timestamp 1713338890
transform 1 0 8639 0 1 2161
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_17
timestamp 1713338890
transform 1 0 8639 0 1 2649
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_18
timestamp 1713338890
transform 1 0 8639 0 1 3137
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_19
timestamp 1713338890
transform 1 0 8639 0 1 3625
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_20
timestamp 1713338890
transform 1 0 8639 0 1 4113
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_21
timestamp 1713338890
transform 1 0 8639 0 1 4601
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_22
timestamp 1713338890
transform 1 0 10567 0 1 1429
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_23
timestamp 1713338890
transform 1 0 10567 0 1 1917
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_24
timestamp 1713338890
transform 1 0 10567 0 1 2405
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_25
timestamp 1713338890
transform 1 0 10567 0 1 2893
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_26
timestamp 1713338890
transform 1 0 10567 0 1 3381
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_27
timestamp 1713338890
transform 1 0 10567 0 1 3869
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_28
timestamp 1713338890
transform 1 0 10567 0 1 4357
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_29
timestamp 1713338890
transform 1 0 10567 0 1 4845
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_30
timestamp 1713338890
transform 1 0 2395 0 1 6065
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_31
timestamp 1713338890
transform 1 0 2395 0 1 5089
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_32
timestamp 1713338890
transform 1 0 2395 0 1 5577
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_33
timestamp 1713338890
transform 1 0 2395 0 1 9009
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_34
timestamp 1713338890
transform 1 0 2395 0 1 9497
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_35
timestamp 1713338890
transform 1 0 2395 0 1 7545
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_36
timestamp 1713338890
transform 1 0 2395 0 1 8033
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_37
timestamp 1713338890
transform 1 0 2395 0 1 8521
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_38
timestamp 1713338890
transform 1 0 4323 0 1 9253
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_39
timestamp 1713338890
transform 1 0 4323 0 1 9741
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_40
timestamp 1713338890
transform 1 0 4323 0 1 6309
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_41
timestamp 1713338890
transform 1 0 4323 0 1 5333
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_42
timestamp 1713338890
transform 1 0 4323 0 1 5821
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_43
timestamp 1713338890
transform 1 0 4323 0 1 7301
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_44
timestamp 1713338890
transform 1 0 4323 0 1 7789
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_45
timestamp 1713338890
transform 1 0 4323 0 1 8277
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_46
timestamp 1713338890
transform 1 0 4323 0 1 8765
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_47
timestamp 1713338890
transform 1 0 8639 0 1 5089
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_48
timestamp 1713338890
transform 1 0 8639 0 1 5577
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_49
timestamp 1713338890
transform 1 0 8639 0 1 6065
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_50
timestamp 1713338890
transform 1 0 8639 0 1 7545
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_51
timestamp 1713338890
transform 1 0 8639 0 1 8033
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_52
timestamp 1713338890
transform 1 0 8639 0 1 8521
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_53
timestamp 1713338890
transform 1 0 8639 0 1 9009
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_54
timestamp 1713338890
transform 1 0 8639 0 1 9497
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_55
timestamp 1713338890
transform 1 0 10567 0 1 5333
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_56
timestamp 1713338890
transform 1 0 10567 0 1 5821
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_57
timestamp 1713338890
transform 1 0 10567 0 1 7301
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_58
timestamp 1713338890
transform 1 0 10567 0 1 7789
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_59
timestamp 1713338890
transform 1 0 10567 0 1 9741
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_60
timestamp 1713338890
transform 1 0 10567 0 1 9253
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_61
timestamp 1713338890
transform 1 0 10567 0 1 8765
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_62
timestamp 1713338890
transform 1 0 10567 0 1 8277
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_63
timestamp 1713338890
transform 1 0 10567 0 1 6309
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_64
timestamp 1713338890
transform 1 0 2395 0 1 9985
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_65
timestamp 1713338890
transform 1 0 8639 0 1 9985
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_66
timestamp 1713338890
transform 1 0 4323 0 1 10229
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_67
timestamp 1713338890
transform 1 0 10567 0 1 10229
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_68
timestamp 1713338890
transform 1 0 2395 0 1 10473
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_69
timestamp 1713338890
transform 1 0 8639 0 1 10473
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_70
timestamp 1713338890
transform 1 0 4323 0 1 10717
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_71
timestamp 1713338890
transform 1 0 10567 0 1 10717
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_72
timestamp 1713338890
transform 1 0 2395 0 1 10961
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_73
timestamp 1713338890
transform 1 0 8639 0 1 10961
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_74
timestamp 1713338890
transform 1 0 4323 0 1 11205
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_75
timestamp 1713338890
transform 1 0 10567 0 1 11205
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_76
timestamp 1713338890
transform 1 0 2395 0 1 11449
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_77
timestamp 1713338890
transform 1 0 8639 0 1 11449
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_78
timestamp 1713338890
transform 1 0 4323 0 1 11693
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_79
timestamp 1713338890
transform 1 0 10567 0 1 11693
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_80
timestamp 1713338890
transform 1 0 2395 0 1 11937
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_81
timestamp 1713338890
transform 1 0 8639 0 1 11937
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_82
timestamp 1713338890
transform 1 0 4323 0 1 12181
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_83
timestamp 1713338890
transform 1 0 10567 0 1 12181
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_84
timestamp 1713338890
transform 1 0 2395 0 1 14393
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_85
timestamp 1713338890
transform 1 0 2395 0 1 14881
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_86
timestamp 1713338890
transform 1 0 2395 0 1 13417
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_87
timestamp 1713338890
transform 1 0 2395 0 1 13905
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_88
timestamp 1713338890
transform 1 0 2395 0 1 15369
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_89
timestamp 1713338890
transform 1 0 2395 0 1 16345
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_90
timestamp 1713338890
transform 1 0 2395 0 1 16833
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_91
timestamp 1713338890
transform 1 0 2395 0 1 17321
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_92
timestamp 1713338890
transform 1 0 2395 0 1 15857
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_93
timestamp 1713338890
transform 1 0 4323 0 1 13173
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_94
timestamp 1713338890
transform 1 0 4323 0 1 13661
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_95
timestamp 1713338890
transform 1 0 4323 0 1 14149
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_96
timestamp 1713338890
transform 1 0 4323 0 1 14637
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_97
timestamp 1713338890
transform 1 0 4323 0 1 15125
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_98
timestamp 1713338890
transform 1 0 4323 0 1 15613
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_99
timestamp 1713338890
transform 1 0 4323 0 1 16101
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_100
timestamp 1713338890
transform 1 0 4323 0 1 16589
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_101
timestamp 1713338890
transform 1 0 4323 0 1 17077
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_102
timestamp 1713338890
transform 1 0 4323 0 1 17565
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_103
timestamp 1713338890
transform 1 0 8639 0 1 13417
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_104
timestamp 1713338890
transform 1 0 8639 0 1 13905
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_105
timestamp 1713338890
transform 1 0 8639 0 1 14393
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_106
timestamp 1713338890
transform 1 0 8639 0 1 14881
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_107
timestamp 1713338890
transform 1 0 8639 0 1 15369
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_108
timestamp 1713338890
transform 1 0 8639 0 1 15857
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_109
timestamp 1713338890
transform 1 0 8639 0 1 16345
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_110
timestamp 1713338890
transform 1 0 8639 0 1 16833
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_111
timestamp 1713338890
transform 1 0 8639 0 1 17321
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_112
timestamp 1713338890
transform 1 0 10567 0 1 13173
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_113
timestamp 1713338890
transform 1 0 10567 0 1 13661
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_114
timestamp 1713338890
transform 1 0 10567 0 1 14149
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_115
timestamp 1713338890
transform 1 0 10567 0 1 14637
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_116
timestamp 1713338890
transform 1 0 10567 0 1 15125
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_117
timestamp 1713338890
transform 1 0 10567 0 1 15613
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_118
timestamp 1713338890
transform 1 0 10567 0 1 16101
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_119
timestamp 1713338890
transform 1 0 10567 0 1 16589
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_120
timestamp 1713338890
transform 1 0 10567 0 1 17077
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_121
timestamp 1713338890
transform 1 0 10567 0 1 17565
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_122
timestamp 1713338890
transform 1 0 2395 0 1 17809
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_123
timestamp 1713338890
transform 1 0 2395 0 1 19289
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_124
timestamp 1713338890
transform 1 0 2395 0 1 19777
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_125
timestamp 1713338890
transform 1 0 2395 0 1 21729
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_126
timestamp 1713338890
transform 1 0 2395 0 1 20265
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_127
timestamp 1713338890
transform 1 0 2395 0 1 20753
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_128
timestamp 1713338890
transform 1 0 2395 0 1 21241
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_129
timestamp 1713338890
transform 1 0 2395 0 1 22217
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_130
timestamp 1713338890
transform 1 0 4323 0 1 19045
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_131
timestamp 1713338890
transform 1 0 4323 0 1 18053
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_132
timestamp 1713338890
transform 1 0 4323 0 1 19533
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_133
timestamp 1713338890
transform 1 0 4323 0 1 20021
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_134
timestamp 1713338890
transform 1 0 4323 0 1 20509
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_135
timestamp 1713338890
transform 1 0 4323 0 1 20997
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_136
timestamp 1713338890
transform 1 0 4323 0 1 21485
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_137
timestamp 1713338890
transform 1 0 4323 0 1 21973
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_138
timestamp 1713338890
transform 1 0 4323 0 1 22461
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_139
timestamp 1713338890
transform 1 0 8639 0 1 17809
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_140
timestamp 1713338890
transform 1 0 8639 0 1 19289
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_141
timestamp 1713338890
transform 1 0 8639 0 1 19777
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_142
timestamp 1713338890
transform 1 0 8639 0 1 20265
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_143
timestamp 1713338890
transform 1 0 8639 0 1 20753
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_144
timestamp 1713338890
transform 1 0 8639 0 1 21241
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_145
timestamp 1713338890
transform 1 0 8639 0 1 21729
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_146
timestamp 1713338890
transform 1 0 8639 0 1 22217
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_147
timestamp 1713338890
transform 1 0 10567 0 1 22461
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_148
timestamp 1713338890
transform 1 0 10567 0 1 21973
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_149
timestamp 1713338890
transform 1 0 10567 0 1 21485
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_150
timestamp 1713338890
transform 1 0 10567 0 1 20997
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_151
timestamp 1713338890
transform 1 0 10567 0 1 20509
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_152
timestamp 1713338890
transform 1 0 10567 0 1 20021
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_153
timestamp 1713338890
transform 1 0 10567 0 1 19045
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_154
timestamp 1713338890
transform 1 0 10567 0 1 19533
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_155
timestamp 1713338890
transform 1 0 10567 0 1 18053
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_156
timestamp 1713338890
transform 1 0 10567 0 1 22949
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_157
timestamp 1713338890
transform 1 0 8639 0 1 22705
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_158
timestamp 1713338890
transform 1 0 2395 0 1 22705
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_159
timestamp 1713338890
transform 1 0 4323 0 1 22949
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_160
timestamp 1713338890
transform 1 0 10567 0 1 23437
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_161
timestamp 1713338890
transform 1 0 8639 0 1 23193
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_162
timestamp 1713338890
transform 1 0 8639 0 1 23681
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_163
timestamp 1713338890
transform 1 0 2395 0 1 23193
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_164
timestamp 1713338890
transform 1 0 4323 0 1 23437
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_165
timestamp 1713338890
transform 1 0 2395 0 1 23681
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_166
timestamp 1713338890
transform 1 0 10567 0 1 23925
box -902 -38 902 38
use M2_M1_CDNS_69033583165359  M2_M1_CDNS_69033583165359_167
timestamp 1713338890
transform 1 0 4323 0 1 23925
box -902 -38 902 38
use M2_M1_CDNS_69033583165360  M2_M1_CDNS_69033583165360_0
timestamp 1713338890
transform 1 0 594 0 1 227
box -524 -146 524 146
use M2_M1_CDNS_69033583165360  M2_M1_CDNS_69033583165360_1
timestamp 1713338890
transform 1 0 5884 0 1 827
box -524 -146 524 146
use M2_M1_CDNS_69033583165360  M2_M1_CDNS_69033583165360_2
timestamp 1713338890
transform 1 0 7078 0 1 227
box -524 -146 524 146
use M2_M1_CDNS_69033583165360  M2_M1_CDNS_69033583165360_3
timestamp 1713338890
transform 1 0 5884 0 1 24527
box -524 -146 524 146
use M2_M1_CDNS_69033583165360  M2_M1_CDNS_69033583165360_4
timestamp 1713338890
transform 1 0 7078 0 1 25127
box -524 -146 524 146
use M2_M1_CDNS_69033583165360  M2_M1_CDNS_69033583165360_5
timestamp 1713338890
transform 1 0 594 0 1 25127
box -524 -146 524 146
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_0
timestamp 1713338890
transform 1 0 1313 0 1 3869
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_1
timestamp 1713338890
transform 1 0 11649 0 1 3869
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_2
timestamp 1713338890
transform 1 0 1313 0 1 9741
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_3
timestamp 1713338890
transform 1 0 11649 0 1 9741
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_4
timestamp 1713338890
transform 1 0 1313 0 1 15613
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_5
timestamp 1713338890
transform 1 0 11649 0 1 15613
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_6
timestamp 1713338890
transform 1 0 1313 0 1 21485
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_7
timestamp 1713338890
transform 1 0 11649 0 1 21485
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165363  M2_M1_CDNS_69033583165363_0
timestamp 1713338890
transform 1 0 2395 0 1 827
box -902 -146 902 146
use M2_M1_CDNS_69033583165363  M2_M1_CDNS_69033583165363_1
timestamp 1713338890
transform 1 0 4323 0 1 227
box -902 -146 902 146
use M2_M1_CDNS_69033583165363  M2_M1_CDNS_69033583165363_2
timestamp 1713338890
transform 1 0 8639 0 1 827
box -902 -146 902 146
use M2_M1_CDNS_69033583165363  M2_M1_CDNS_69033583165363_3
timestamp 1713338890
transform 1 0 10567 0 1 227
box -902 -146 902 146
use M2_M1_CDNS_69033583165363  M2_M1_CDNS_69033583165363_4
timestamp 1713338890
transform 1 0 8639 0 1 24527
box -902 -146 902 146
use M2_M1_CDNS_69033583165363  M2_M1_CDNS_69033583165363_5
timestamp 1713338890
transform 1 0 2395 0 1 24527
box -902 -146 902 146
use M2_M1_CDNS_69033583165363  M2_M1_CDNS_69033583165363_6
timestamp 1713338890
transform 1 0 10567 0 1 25127
box -902 -146 902 146
use M2_M1_CDNS_69033583165363  M2_M1_CDNS_69033583165363_7
timestamp 1713338890
transform 1 0 4323 0 1 25127
box -902 -146 902 146
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_0
timestamp 1713338890
transform 1 0 5884 0 1 4601
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_1
timestamp 1713338890
transform 1 0 5884 0 1 4113
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_2
timestamp 1713338890
transform 1 0 5884 0 1 3625
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_3
timestamp 1713338890
transform 1 0 5884 0 1 3137
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_4
timestamp 1713338890
transform 1 0 5884 0 1 2649
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_5
timestamp 1713338890
transform 1 0 5884 0 1 2161
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_6
timestamp 1713338890
transform 1 0 5884 0 1 1673
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_7
timestamp 1713338890
transform 1 0 7078 0 1 1429
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_8
timestamp 1713338890
transform 1 0 7078 0 1 1917
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_9
timestamp 1713338890
transform 1 0 7078 0 1 2405
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_10
timestamp 1713338890
transform 1 0 7078 0 1 2893
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_11
timestamp 1713338890
transform 1 0 7078 0 1 3381
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_12
timestamp 1713338890
transform 1 0 7078 0 1 3869
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_13
timestamp 1713338890
transform 1 0 7078 0 1 4357
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_14
timestamp 1713338890
transform 1 0 7078 0 1 4845
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_15
timestamp 1713338890
transform 1 0 5884 0 1 6065
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_16
timestamp 1713338890
transform 1 0 5884 0 1 5577
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_17
timestamp 1713338890
transform 1 0 5884 0 1 5089
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_18
timestamp 1713338890
transform 1 0 5884 0 1 9497
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_19
timestamp 1713338890
transform 1 0 5884 0 1 9009
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_20
timestamp 1713338890
transform 1 0 5884 0 1 8521
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_21
timestamp 1713338890
transform 1 0 5884 0 1 8033
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_22
timestamp 1713338890
transform 1 0 5884 0 1 7545
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_23
timestamp 1713338890
transform 1 0 7078 0 1 5333
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_24
timestamp 1713338890
transform 1 0 7078 0 1 5821
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_25
timestamp 1713338890
transform 1 0 7078 0 1 6309
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_26
timestamp 1713338890
transform 1 0 7078 0 1 7301
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_27
timestamp 1713338890
transform 1 0 7078 0 1 7789
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_28
timestamp 1713338890
transform 1 0 7078 0 1 8277
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_29
timestamp 1713338890
transform 1 0 7078 0 1 8765
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_30
timestamp 1713338890
transform 1 0 7078 0 1 9253
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_31
timestamp 1713338890
transform 1 0 7078 0 1 9741
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_32
timestamp 1713338890
transform 1 0 5884 0 1 9985
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_33
timestamp 1713338890
transform 1 0 7078 0 1 10229
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_34
timestamp 1713338890
transform 1 0 5884 0 1 10473
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_35
timestamp 1713338890
transform 1 0 7078 0 1 10717
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_36
timestamp 1713338890
transform 1 0 5884 0 1 10961
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_37
timestamp 1713338890
transform 1 0 7078 0 1 11205
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_38
timestamp 1713338890
transform 1 0 5884 0 1 11449
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_39
timestamp 1713338890
transform 1 0 7078 0 1 11693
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_40
timestamp 1713338890
transform 1 0 5884 0 1 11937
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_41
timestamp 1713338890
transform 1 0 7078 0 1 12181
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_42
timestamp 1713338890
transform 1 0 5884 0 1 17321
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_43
timestamp 1713338890
transform 1 0 5884 0 1 16833
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_44
timestamp 1713338890
transform 1 0 5884 0 1 16345
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_45
timestamp 1713338890
transform 1 0 5884 0 1 15857
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_46
timestamp 1713338890
transform 1 0 5884 0 1 15369
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_47
timestamp 1713338890
transform 1 0 5884 0 1 14881
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_48
timestamp 1713338890
transform 1 0 5884 0 1 14393
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_49
timestamp 1713338890
transform 1 0 5884 0 1 13905
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_50
timestamp 1713338890
transform 1 0 5884 0 1 13417
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_51
timestamp 1713338890
transform 1 0 7078 0 1 13173
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_52
timestamp 1713338890
transform 1 0 7078 0 1 13661
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_53
timestamp 1713338890
transform 1 0 7078 0 1 14149
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_54
timestamp 1713338890
transform 1 0 7078 0 1 14637
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_55
timestamp 1713338890
transform 1 0 7078 0 1 15125
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_56
timestamp 1713338890
transform 1 0 7078 0 1 15613
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_57
timestamp 1713338890
transform 1 0 7078 0 1 16101
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_58
timestamp 1713338890
transform 1 0 7078 0 1 16589
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_59
timestamp 1713338890
transform 1 0 7078 0 1 17077
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_60
timestamp 1713338890
transform 1 0 7078 0 1 17565
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_61
timestamp 1713338890
transform 1 0 5884 0 1 17809
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_62
timestamp 1713338890
transform 1 0 5884 0 1 21241
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_63
timestamp 1713338890
transform 1 0 5884 0 1 22217
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_64
timestamp 1713338890
transform 1 0 5884 0 1 21729
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_65
timestamp 1713338890
transform 1 0 5884 0 1 20753
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_66
timestamp 1713338890
transform 1 0 5884 0 1 20265
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_67
timestamp 1713338890
transform 1 0 5884 0 1 19777
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_68
timestamp 1713338890
transform 1 0 5884 0 1 19289
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_69
timestamp 1713338890
transform 1 0 7078 0 1 18053
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_70
timestamp 1713338890
transform 1 0 7078 0 1 19045
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_71
timestamp 1713338890
transform 1 0 7078 0 1 19533
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_72
timestamp 1713338890
transform 1 0 7078 0 1 20021
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_73
timestamp 1713338890
transform 1 0 7078 0 1 20509
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_74
timestamp 1713338890
transform 1 0 7078 0 1 20997
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_75
timestamp 1713338890
transform 1 0 7078 0 1 21485
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_76
timestamp 1713338890
transform 1 0 7078 0 1 21973
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_77
timestamp 1713338890
transform 1 0 7078 0 1 22461
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_78
timestamp 1713338890
transform 1 0 7078 0 1 22949
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_79
timestamp 1713338890
transform 1 0 5884 0 1 22705
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_80
timestamp 1713338890
transform 1 0 7078 0 1 23437
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_81
timestamp 1713338890
transform 1 0 5884 0 1 23681
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_82
timestamp 1713338890
transform 1 0 5884 0 1 23193
box -524 -38 524 38
use M2_M1_CDNS_69033583165364  M2_M1_CDNS_69033583165364_83
timestamp 1713338890
transform 1 0 7078 0 1 23925
box -524 -38 524 38
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_0
timestamp 1713338890
transform 0 -1 11481 1 0 1481
box -88 -44 4864 10044
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_1
timestamp 1713338890
transform 0 -1 11481 1 0 7353
box -88 -44 4864 10044
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_2
timestamp 1713338890
transform 0 -1 11481 1 0 13225
box -88 -44 4864 10044
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_3
timestamp 1713338890
transform 0 -1 11481 1 0 19097
box -88 -44 4864 10044
<< end >>
