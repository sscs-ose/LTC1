** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/LF.sch
**.subckt LF VSS VCNTL VDD
*.iopin VSS
*.iopin VCNTL
*.iopin VDD
x1 VCNTL net1 VDD res_sch
x2 VSS net1 cap80p
x3 VSS VCNTL cap3p
**.ends

* expanding   symbol:  res_sch.sym # of pins=3
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/res_sch.sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/res_sch.sch
.subckt res_sch A B VDD
*.iopin VDD
*.iopin A
*.iopin B
XR1 B A VDD ppolyf_u r_width=0.8e-6 r_length=100e-6 m=1
.ends


* expanding   symbol:  cap80p.sym # of pins=2
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/cap80p.sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/cap80p.sch
.subckt cap80p N P
*.iopin P
*.iopin N
XC1 P N cap_mim_2f0_m4m5_noshield c_width=25e-6 c_length=25e-6 m=64
.ends


* expanding   symbol:  cap3p.sym # of pins=2
** sym_path: /home/shahid/GF180Projects/Top_test/top/xschem/cap3p.sym
** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/cap3p.sch
.subckt cap3p Nn Pp
*.iopin Pp
*.iopin Nn
XC1 Pp Nn cap_mim_2f0_m4m5_noshield c_width=42.5e-6 c_length=42.5e-6 m=1
.ends

.end
