** sch_path: /home/shahid/GF180Projects/Tapeout/Xschem/Logic_Gates/Inverter.sch
.subckt Inverter IN OUT VDD VSS
*.PININFO IN:I OUT:O VDD:B VSS:B
M1 OUT IN VDD VDD pfet_03v3 L=0.28u W=1u nf=1 m=1
M2 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.5u nf=1 m=1
.ends
.end
