* NGSPICE file created from CLK_div_31_mag_flat.ext - technology: gf180mcuC

.subckt pex_CLK_div_31_mag VSS VDD Q0 Q1 Q2 Q3 Q4 Vdiv31 RST CLK
X0 a_2069_4071# Q0.t3 a_1909_4071# VSS.t142 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X1 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand2_mag_3.IN1 VDD.t213 VDD.t212 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 VDD VDD.t40 JK_FF_mag_3.nand3_mag_2.OUT VDD.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VSS.t172 VSS.t171 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X4 a_1185_4071# JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_1.OUT VSS.t49 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X5 VDD JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.QB VDD.t283 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X6 JK_FF_mag_3.nand3_mag_1.OUT RST.t2 VDD.t153 VDD.t152 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X7 VSS JK_FF_mag_3.nand3_mag_2.OUT a_4405_4070# VSS.t27 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X8 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_3.IN1 VDD.t5 VDD.t4 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X9 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN Q2.t3 a_7993_3052# VSS.t99 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X10 Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VDD.t92 VDD.t91 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X11 VSS JK_FF_mag_2.nand3_mag_1.OUT a_621_4071# VSS.t64 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X12 VDD Q3.t3 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t165 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t189 VSS.t188 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X14 VDD Q3.t4 JK_FF_mag_4.nand3_mag_0.OUT VDD.t168 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X15 JK_FF_mag_4.QB Q4.t3 a_8642_248# VSS.t209 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t309 VDD.t308 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X17 or_2_mag_0.GF_INV_MAG_1.IN or_2_mag_0.IN1 a_11530_2405# VDD.t204 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X18 VDD JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_1.IN1 VDD.t137 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X19 JK_FF_mag_4.nand2_mag_1.IN2 JK_FF_mag_4.nand3_mag_1.IN1 VDD.t128 VDD.t127 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.QB a_3724_1302# VSS.t81 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X21 a_516_196# VDD.t362 VSS.t146 VSS.t145 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X22 VDD RST.t3 JK_FF_mag_4.nand3_mag_1.OUT VDD.t154 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X23 VDD Q3.t5 JK_FF_mag_1.QB VDD.t171 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X24 JK_FF_mag_4.nand2_mag_3.IN1 Q3.t6 VDD.t175 VDD.t174 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X25 a_5416_1346# JK_FF_mag_1.nand2_mag_1.IN2 VSS.t220 VSS.t219 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X26 JK_FF_mag_2.QB Q1.t3 VDD.t265 VDD.t264 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X27 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VDD.t56 VDD.t55 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X28 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_1810_1337# VSS.t71 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X29 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand3_mag_0.OUT VDD.t1 VDD.t0 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X30 or_2_mag_0.IN1 Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VSS.t197 VSS.t196 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X31 JK_FF_mag_4.nand2_mag_4.IN2 JK_FF_mag_4.nand2_mag_3.IN1 a_8078_248# VSS.t216 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X32 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 a_1400_196# VSS.t111 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X33 VDD Q2.t4 JK_FF_mag_0.QB.t0 VDD.t339 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X34 VDD JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand2_mag_1.IN2 VDD.t325 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 a_5570_249# JK_FF_mag_1.nand2_mag_4.IN2 VSS.t214 VSS.t213 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X36 a_6796_1301# Q3.t7 a_6636_1301# VSS.t87 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X37 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_2.OUT VDD.t71 VDD.t70 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X38 VDD Q3.t8 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t176 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X39 VDD JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t78 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X40 Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS.t23 VSS.t22 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X41 a_7514_204# RST.t4 a_7354_204# VSS.t82 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X42 VDD Q1.t4 JK_FF_mag_0.nand3_mag_2.OUT VDD.t266 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X43 a_8944_3063# nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS.t17 VSS.t16 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X44 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 VDD.t203 VDD.t202 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X45 a_4399_2973# JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 VSS.t21 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X46 VDD JK_FF_mag_0.QB.t3 Q2.t1 VDD.t245 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X47 a_5123_2973# CLK.t0 a_4963_2973# VSS.t54 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X48 JK_FF_mag_0.nand2_mag_3.IN1 Q1.t5 VDD.t270 VDD.t269 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X49 a_2528_240# JK_FF_mag_0.nand2_mag_4.IN2 VSS.t97 VSS.t96 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X50 VDD Q3.t9 JK_FF_mag_4.nand3_mag_2.OUT VDD.t179 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X51 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT VDD.t144 VDD.t143 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X52 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 VDD.t132 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X53 VSS CLK.t1 JK_FF_mag_3.nand2_mag_3.IN1 VSS.t58 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X54 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN Q3.t10 a_8944_3063# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X55 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB.t4 VDD.t249 VDD.t248 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X56 VDD Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VDD.t300 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X57 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN Q3.t11 a_7994_3809# VSS.t88 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X58 Q2 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t119 VDD.t118 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X59 Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VSS.t174 VSS.t173 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X60 VDD Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VDD.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X61 a_4282_205# JK_FF_mag_1.nand3_mag_2.OUT VSS.t31 VSS.t30 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X62 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t88 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X63 VDD Q1.t6 JK_FF_mag_0.nand3_mag_0.OUT VDD.t271 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X64 VDD Q2.t5 JK_FF_mag_1.nand3_mag_0.OUT VDD.t342 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X65 VSS Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS.t202 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X66 a_1240_196# JK_FF_mag_0.nand3_mag_2.OUT VSS.t79 VSS.t78 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X67 VSS JK_FF_mag_3.nand3_mag_1.OUT a_3681_4070# VSS.t18 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X68 VDD Q1.t7 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t274 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X69 nand_5_mag_0.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t336 VDD.t335 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X70 VSS Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VSS.t24 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X71 JK_FF_mag_1.nand3_mag_2.OUT VDD.t37 VDD.t39 VDD.t38 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X72 JK_FF_mag_3.QB Q0.t4 VDD.t244 VDD.t243 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X73 VDD JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand3_mag_1.IN1 VDD.t52 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X74 JK_FF_mag_1.nand2_mag_3.IN1 Q2.t6 VDD.t346 VDD.t345 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X75 JK_FF_mag_1.QB Q3.t12 a_5570_249# VSS.t89 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X76 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t77 VDD.t76 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X77 a_7924_1345# JK_FF_mag_4.nand3_mag_1.IN1 VSS.t69 VSS.t68 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X78 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand3_mag_1.OUT a_7360_1345# VSS.t74 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X79 a_4969_4070# Q0.t5 JK_FF_mag_3.nand3_mag_2.OUT VSS.t141 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X80 JK_FF_mag_3.nand3_mag_2.OUT CLK.t2 VDD.t109 VDD.t108 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 VDD JK_FF_mag_2.QB JK_FF_mag_2.nand3_mag_0.OUT VDD.t207 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X82 JK_FF_mag_1.nand3_mag_0.OUT VDD.t34 VDD.t36 VDD.t35 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X83 a_6790_204# Q3.t13 a_6630_204# VSS.t90 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X84 Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VDD.t223 VDD.t222 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X85 VSS JK_FF_mag_3.nand2_mag_4.IN2 a_3117_4070# VSS.t121 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X86 a_3681_4070# JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_4.IN2 VSS.t117 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X87 VSS VDD.t363 a_5129_4070# VSS.t147 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X88 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS.t208 VSS.t207 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X89 VDD VDD.t30 JK_FF_mag_2.nand3_mag_0.OUT VDD.t31 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X90 RST nand_5_mag_0.GF_INV_MAG_0.IN VDD.t358 VDD.t357 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X91 VDD RST.t5 JK_FF_mag_1.nand3_mag_1.OUT VDD.t157 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X92 VDD JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_1.OUT VDD.t102 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X93 VDD JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand2_mag_1.IN2 VDD.t99 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X94 a_4405_4070# RST.t6 a_4245_4070# VSS.t83 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X95 JK_FF_mag_0.nand3_mag_2.OUT Q2.t7 VDD.t348 VDD.t347 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X96 VSS JK_FF_mag_2.nand2_mag_4.IN2 a_57_4071# VSS.t185 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X97 a_621_4071# JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_4.IN2 VSS.t3 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X98 a_7360_1345# JK_FF_mag_4.nand3_mag_0.OUT VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X99 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN Q1.t8 a_9908_3052# VSS.t39 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X100 JK_FF_mag_4.nand3_mag_0.OUT VDD.t27 VDD.t29 VDD.t28 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X101 VDD CLK.t3 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t110 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X102 VDD JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand2_mag_1.IN2 VDD.t96 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X103 JK_FF_mag_2.nand3_mag_0.OUT Q0.t6 VDD.t242 VDD.t241 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X104 nand_5_mag_0.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t222 VSS.t221 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X105 a_11530_2405# Q4.t4 VDD.t311 VDD.t310 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X106 VDD JK_FF_mag_4.QB Q4.t1 VDD.t259 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X107 VDD RST.t7 JK_FF_mag_0.nand3_mag_1.OUT VDD.t160 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X108 JK_FF_mag_4.nand2_mag_1.IN2 JK_FF_mag_4.nand2_mag_3.IN1 a_7924_1345# VSS.t215 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X109 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_2.IN2 VDD.t263 VDD.t262 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X110 and_5_mag_0.VOUT and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD.t185 VDD.t184 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X111 a_3724_1302# Q2.t8 a_3564_1302# VSS.t225 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X112 Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VSS.t46 VSS.t45 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X113 RST nand_5_mag_0.GF_INV_MAG_0.IN VSS.t234 VSS.t233 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X114 JK_FF_mag_4.nand3_mag_2.OUT Q4.t5 VDD.t313 VDD.t312 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X115 VDD JK_FF_mag_2.nand2_mag_1.IN2 Q1.t0 VDD.t44 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X116 JK_FF_mag_4.nand2_mag_3.IN1 Q3.t14 VSS.t92 VSS.t91 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X117 a_3558_205# VDD.t365 VSS.t151 VSS.t150 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X118 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_3.IN1 VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X119 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT a_1246_1337# VSS.t38 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X120 Q4 JK_FF_mag_4.nand2_mag_1.IN2 VDD.t196 VDD.t195 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X121 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X122 a_57_4071# Q1.t9 JK_FF_mag_2.QB VSS.t179 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X123 VDD JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand3_mag_1.OUT VDD.t250 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X124 a_1810_1337# JK_FF_mag_0.nand3_mag_1.IN1 VSS.t110 VSS.t109 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X125 a_3564_1302# VDD.t366 VSS.t153 VSS.t152 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X126 JK_FF_mag_4.QB JK_FF_mag_4.nand2_mag_4.IN2 VDD.t75 VDD.t74 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X127 VDD Q2.t9 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t349 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X128 Vdiv31 or_2_mag_0.GF_INV_MAG_1.IN VDD.t356 VDD.t355 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X129 a_4442_205# RST.t8 a_4282_205# VSS.t84 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X130 Q2 JK_FF_mag_0.QB.t5 a_2374_1337# VSS.t143 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X131 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t228 VDD.t227 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X132 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VDD.t82 VDD.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X133 a_6636_1301# VDD.t367 VSS.t155 VSS.t154 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X134 Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VDD.t221 VDD.t220 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X135 a_5006_249# JK_FF_mag_1.nand3_mag_1.OUT VSS.t77 VSS.t76 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X136 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT VDD.t299 VDD.t298 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X137 a_2374_1337# JK_FF_mag_0.nand2_mag_1.IN2 VSS.t63 VSS.t62 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X138 VDD Q2.t10 JK_FF_mag_1.nand3_mag_2.OUT VDD.t352 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X139 JK_FF_mag_4.nand3_mag_2.OUT Q4.t6 a_6790_204# VSS.t210 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X140 a_9908_3052# nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS.t40 VSS.t39 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X141 VSS or_2_mag_0.IN1 or_2_mag_0.GF_INV_MAG_1.IN VSS.t112 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X142 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_4852_1346# VSS.t44 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X143 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t132 VSS.t131 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X144 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.IN2 VDD.t48 VDD.t47 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X145 a_676_196# Q1.t10 a_516_196# VSS.t180 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X146 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_1.IN1 VDD.t126 VDD.t125 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X147 JK_FF_mag_0.nand2_mag_3.IN1 Q1.t11 VSS.t182 VSS.t181 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X148 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN Q0.t7 VDD.t240 VDD.t239 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X149 a_8945_3798# and_5_mag_0.and2_mag_2.IN2 VSS.t178 VSS.t177 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X150 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK.t4 a_9909_3809# VSS.t9 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X151 VDD JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t140 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X152 VSS JK_FF_mag_2.nand3_mag_0.OUT a_1339_2974# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X153 JK_FF_mag_0.nand3_mag_0.OUT VDD.t24 VDD.t26 VDD.t25 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X154 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand3_mag_1.IN1 VDD.t9 VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X155 a_3718_205# Q2.t11 a_3558_205# VSS.t226 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X156 a_1903_2974# JK_FF_mag_2.QB JK_FF_mag_2.nand3_mag_0.OUT VSS.t115 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X157 or_2_mag_0.GF_INV_MAG_1.IN Q4.t7 VSS.t212 VSS.t211 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X158 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB.t6 a_682_1293# VSS.t144 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X159 Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VDD.t329 VDD.t328 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X160 VSS VDD.t368 a_2063_2974# VSS.t115 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X161 VDD Q4.t8 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t314 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X162 a_7047_3047# Q0.t8 VSS.t140 VSS.t139 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X163 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t84 VDD.t83 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X164 VDD JK_FF_mag_1.QB Q3.t0 VDD.t149 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X165 Q4 JK_FF_mag_4.QB a_8488_1345# VSS.t176 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X166 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN Q0.t9 VDD.t238 VDD.t237 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X167 VSS JK_FF_mag_3.nand3_mag_1.IN1 a_3835_2973# VSS.t51 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X168 VDD Q0.t10 JK_FF_mag_2.nand2_mag_3.IN1 VDD.t234 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X169 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT VDD.t338 VDD.t337 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X170 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN Q2.t12 a_8945_3798# VSS.t177 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X171 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_1.OUT VDD.t124 VDD.t123 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X172 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_1.IN1 a_7514_204# VSS.t67 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X173 a_682_1293# Q1.t12 a_522_1293# VSS.t183 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X174 a_3117_4070# Q0.t11 JK_FF_mag_3.QB VSS.t138 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X175 a_5129_4070# CLK.t5 a_4969_4070# VSS.t61 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X176 VSS JK_FF_mag_2.nand3_mag_1.IN1 a_775_2974# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X177 a_2063_2974# Q0.t12 a_1903_2974# VSS.t115 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X178 JK_FF_mag_1.nand2_mag_3.IN1 Q2.t13 VSS.t228 VSS.t227 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X179 and_5_mag_0.VOUT and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS.t95 VSS.t94 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X180 VDD JK_FF_mag_3.nand2_mag_1.IN2 Q0.t0 VDD.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X181 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_5006_249# VSS.t43 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X182 a_8488_1345# JK_FF_mag_4.nand2_mag_1.IN2 VSS.t105 VSS.t104 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X183 a_4245_4070# JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_1.OUT VSS.t50 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X184 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand2_mag_3.IN1 VDD.t211 VDD.t210 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X185 VDD Q1.t13 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t277 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X186 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN Q4.t9 a_7047_3047# VSS.t139 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X187 Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VSS.t127 VSS.t126 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X188 a_8642_248# JK_FF_mag_4.nand2_mag_4.IN2 VSS.t35 VSS.t34 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X189 and_5_mag_0.and2_mag_1.IN2 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t297 VDD.t296 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X190 VSS JK_FF_mag_2.nand2_mag_1.IN2 a_211_2974# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X191 JK_FF_mag_0.QB Q2.t14 a_2528_240# VSS.t229 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X192 a_775_2974# JK_FF_mag_2.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_1.IN2 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X193 VDD JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.nand3_mag_1.IN1 VDD.t224 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X194 VDD JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_0.OUT VDD.t305 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X195 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_2.OUT VDD.t360 VDD.t359 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X196 Q0 JK_FF_mag_3.QB VDD.t304 VDD.t303 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X197 VDD VDD.t20 JK_FF_mag_3.nand3_mag_0.OUT VDD.t21 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X198 VDD Q1.t14 JK_FF_mag_2.nand3_mag_2.OUT VDD.t280 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X199 a_9909_3809# and_5_mag_0.and2_mag_3.IN2 VSS.t10 VSS.t9 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X200 JK_FF_mag_0.nand3_mag_2.OUT Q2.t15 a_676_196# VSS.t230 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X201 VDD VDD.t16 JK_FF_mag_2.nand3_mag_2.OUT VDD.t17 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X202 and_5_mag_0.and2_mag_3.IN2 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD.t73 VDD.t72 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X203 Q1 JK_FF_mag_2.QB VDD.t206 VDD.t205 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X204 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VDD.t191 VDD.t190 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X205 a_1246_1337# JK_FF_mag_0.nand3_mag_0.OUT VSS.t201 VSS.t200 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X206 JK_FF_mag_2.nand3_mag_1.OUT RST.t9 VDD.t164 VDD.t163 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X207 and_5_mag_0.and2_mag_3.IN2 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS.t33 VSS.t32 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X208 Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VDD.t254 VDD.t253 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X209 a_1400_196# RST.t10 a_1240_196# VSS.t85 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X210 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_4.IN2 VDD.t187 VDD.t186 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X211 VSS JK_FF_mag_2.nand3_mag_2.OUT a_1345_4071# VSS.t168 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X212 JK_FF_mag_2.nand3_mag_2.OUT Q0.t13 VDD.t233 VDD.t232 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X213 Vdiv31 or_2_mag_0.GF_INV_MAG_1.IN VSS.t232 VSS.t231 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X214 JK_FF_mag_4.nand2_mag_4.IN2 JK_FF_mag_4.nand3_mag_1.OUT VDD.t136 VDD.t135 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X215 VDD JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_1.OUT VDD.t93 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X216 a_7993_3052# nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS.t100 VSS.t99 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X217 a_7354_204# JK_FF_mag_4.nand3_mag_2.OUT VSS.t236 VSS.t235 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X218 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_1964_240# VSS.t70 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X219 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t7 VDD.t6 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X220 JK_FF_mag_0.nand3_mag_2.OUT VDD.t13 VDD.t15 VDD.t14 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X221 VDD Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VDD.t214 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X222 VDD JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand3_mag_1.OUT VDD.t67 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X223 VDD JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_4.IN2 VDD.t120 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X224 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_1.IN2 VDD.t189 VDD.t188 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X225 a_7048_3814# Q0.t14 VSS.t137 VSS.t136 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X226 Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VSS.t125 VSS.t124 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X227 JK_FF_mag_4.nand3_mag_0.OUT JK_FF_mag_4.QB VDD.t258 VDD.t257 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X228 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT a_4288_1346# VSS.t75 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X229 a_4852_1346# JK_FF_mag_1.nand3_mag_1.IN1 VSS.t6 VSS.t5 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X230 VSS Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VSS.t118 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X231 or_2_mag_0.IN1 Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VDD.t295 VDD.t294 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X232 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t201 VDD.t200 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X233 VDD Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VDD.t49 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X234 Q3 JK_FF_mag_1.QB a_5416_1346# VSS.t80 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X235 JK_FF_mag_4.nand3_mag_2.OUT VDD.t10 VDD.t12 VDD.t11 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X236 VDD Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VDD.t288 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X237 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN Q1.t15 a_7048_3814# VSS.t136 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X238 a_4288_1346# JK_FF_mag_1.nand3_mag_0.OUT VSS.t224 VSS.t223 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X239 a_1964_240# JK_FF_mag_0.nand3_mag_1.OUT VSS.t37 VSS.t36 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X240 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 a_4442_205# VSS.t4 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X241 VDD Q4.t10 JK_FF_mag_4.QB VDD.t317 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X242 VSS Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VSS.t11 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X243 a_1339_2974# JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X244 Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VDD.t63 VDD.t62 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X245 VDD Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VDD.t192 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X246 VSS Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VSS.t190 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X247 VSS JK_FF_mag_3.nand2_mag_1.IN2 a_3271_2973# VSS.t55 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X248 Q3 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t331 VDD.t330 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X249 JK_FF_mag_4.nand3_mag_0.OUT JK_FF_mag_4.QB a_6796_1301# VSS.t175 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X250 a_3835_2973# JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_1.IN2 VSS.t116 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X251 VDD Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VDD.t291 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X252 and_5_mag_0.and2_mag_1.IN2 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t199 VSS.t198 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X253 VSS Q0.t15 JK_FF_mag_2.nand2_mag_3.IN1 VSS.t133 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X254 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t129 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X255 a_522_1293# VDD.t371 VSS.t159 VSS.t158 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X256 Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VSS.t218 VSS.t217 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X257 a_6630_204# VDD.t372 VSS.t161 VSS.t160 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X258 VDD JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand2_mag_4.IN2 VDD.t322 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X259 JK_FF_mag_1.nand3_mag_2.OUT Q3.t15 VDD.t183 VDD.t182 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X260 VSS JK_FF_mag_3.nand3_mag_0.OUT a_4399_2973# VSS.t128 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X261 a_4963_2973# JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_0.OUT VSS.t206 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X262 VSS Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VSS.t101 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X263 a_3271_2973# JK_FF_mag_3.QB Q0.t2 VSS.t205 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X264 VSS VDD.t373 a_5123_2973# VSS.t162 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X265 Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VDD.t256 VDD.t255 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X266 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_4.IN2 VDD.t321 VDD.t320 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X267 VSS Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VSS.t193 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X268 VDD CLK.t6 JK_FF_mag_3.nand2_mag_3.IN1 VDD.t113 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X269 a_7994_3809# and_5_mag_0.and2_mag_1.IN2 VSS.t98 VSS.t88 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X270 a_211_2974# JK_FF_mag_2.QB Q1.t2 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X271 VDD and_5_mag_0.VOUT Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VDD.t197 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=1u
X272 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t42 VSS.t41 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X273 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_1.OUT VDD.t61 VDD.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X274 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT VDD.t146 VDD.t145 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X275 JK_FF_mag_3.nand3_mag_0.OUT CLK.t7 VDD.t117 VDD.t116 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X276 a_8078_248# JK_FF_mag_4.nand3_mag_1.OUT VSS.t73 VSS.t72 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X277 a_1909_4071# Q1.t16 JK_FF_mag_2.nand3_mag_2.OUT VSS.t184 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X278 VSS and_5_mag_0.VOUT Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VSS.t106 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=1u
X279 VSS VDD.t374 a_2069_4071# VSS.t165 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X280 VDD JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_4.IN2 VDD.t57 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X281 VDD Q2.t16 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t332 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X282 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.QB VDD.t148 VDD.t147 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X283 JK_FF_mag_1.nand3_mag_2.OUT Q3.t16 a_3718_205# VSS.t93 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X284 a_1345_4071# RST.t11 a_1185_4071# VSS.t86 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X285 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD.t287 VDD.t286 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X286 VDD Q0.t16 JK_FF_mag_3.nand3_mag_2.OUT VDD.t229 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X287 VDD JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.QB VDD.t217 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 Q0.n13 Q0.t12 36.935
R1 Q0.n8 Q0.t3 36.935
R2 Q0.n2 Q0.t5 36.935
R3 Q0.n27 Q0.t11 31.4332
R4 Q0.n1 Q0.t7 30.9379
R5 Q0.n0 Q0.t9 30.9379
R6 Q0.n5 Q0.t10 25.4744
R7 Q0.n1 Q0.t8 21.6422
R8 Q0.n0 Q0.t14 21.6422
R9 Q0.n13 Q0.t6 18.1962
R10 Q0.n8 Q0.t13 18.1962
R11 Q0.n2 Q0.t16 18.1962
R12 Q0.n27 Q0.t4 15.3826
R13 Q0.n5 Q0.t15 14.1417
R14 Q0.n25 Q0.t2 7.09905
R15 Q0.n28 Q0.n27 6.86029
R16 Q0.n31 Q0 6.54296
R17 Q0.n31 Q0.n30 4.54543
R18 Q0.n19 Q0.n18 4.50225
R19 Q0.n10 Q0.n7 4.5005
R20 Q0.n12 Q0.n11 4.5005
R21 Q0.n16 Q0.n14 4.5005
R22 Q0.n16 Q0.n15 4.5005
R23 Q0.n22 Q0.n21 4.5005
R24 Q0 Q0.n1 4.11094
R25 Q0 Q0.n0 4.11094
R26 Q0.n30 Q0.n29 3.5302
R27 Q0.n25 Q0.n24 3.25053
R28 Q0.n24 Q0.t0 2.2755
R29 Q0.n24 Q0.n23 2.2755
R30 Q0 Q0.n26 2.25518
R31 Q0.n17 Q0.n6 2.25107
R32 Q0.n20 Q0.n4 2.2505
R33 Q0.n3 Q0.n2 2.13459
R34 Q0.n9 Q0.n8 2.12444
R35 Q0.n14 Q0.n13 2.12188
R36 Q0.n16 Q0.n12 1.71671
R37 Q0.n29 Q0 1.52306
R38 Q0.n9 Q0.n7 1.50503
R39 Q0.n19 Q0.n5 1.42118
R40 Q0.n30 Q0.n3 1.37844
R41 Q0.n29 Q0.n28 1.12067
R42 Q0.n18 Q0.n17 0.932217
R43 Q0 Q0.n22 0.634607
R44 Q0 Q0.n31 0.485557
R45 Q0.n21 Q0 0.1605
R46 Q0.n26 Q0.n25 0.0905
R47 Q0.n28 Q0 0.0857632
R48 Q0.n3 Q0 0.0800273
R49 Q0.n26 Q0 0.073625
R50 Q0.n15 Q0 0.0457995
R51 Q0.n10 Q0 0.0457995
R52 Q0.n12 Q0.n7 0.0386356
R53 Q0.n15 Q0.n6 0.0377414
R54 Q0.n11 Q0.n10 0.0377414
R55 Q0.n21 Q0.n20 0.03175
R56 Q0.n22 Q0.n4 0.03175
R57 Q0.n17 Q0.n16 0.0122182
R58 Q0.n14 Q0.n6 0.00360345
R59 Q0.n11 Q0.n9 0.00203726
R60 Q0.n20 Q0.n19 0.00175
R61 Q0.n18 Q0.n4 0.00100174
R62 VSS.n191 VSS.n170 3.10619e+06
R63 VSS.n193 VSS.n192 160965
R64 VSS.n50 VSS.n49 19500
R65 VSS.t106 VSS.n86 18457.5
R66 VSS.n55 VSS.n50 16250
R67 VSS.n169 VSS.n168 9901.08
R68 VSS.n48 VSS.n47 9750
R69 VSS.n142 VSS.n141 7008.64
R70 VSS.n250 VSS.n249 6332.13
R71 VSS.n264 VSS.t181 6054.76
R72 VSS.n24 VSS.t145 5986.26
R73 VSS.n293 VSS.n292 5115.09
R74 VSS.t133 VSS.n264 4342.23
R75 VSS.n105 VSS.t211 3750
R76 VSS.n170 VSS.n169 3205.8
R77 VSS.n132 VSS.n58 3178.41
R78 VSS.n193 VSS.n57 3124.39
R79 VSS.t196 VSS.n85 2912.27
R80 VSS.t173 VSS.n84 2912.27
R81 VSS.t126 VSS.n82 2912.27
R82 VSS.n125 VSS.t217 2912.27
R83 VSS.n126 VSS.t171 2912.27
R84 VSS.t45 VSS.n83 2906.73
R85 VSS.n247 VSS.n246 2360.75
R86 VSS.t38 VSS.t109 2307.56
R87 VSS.t200 VSS.t144 2307.56
R88 VSS.t219 VSS.t44 2307.56
R89 VSS.t5 VSS.t75 2307.56
R90 VSS.t223 VSS.t81 2307.56
R91 VSS.t206 VSS.t128 2307.56
R92 VSS.t21 VSS.t51 2307.56
R93 VSS.t116 VSS.t55 2307.56
R94 VSS.t74 VSS.t68 2307.56
R95 VSS.t0 VSS.t175 2307.56
R96 VSS.t91 VSS.t154 2307.56
R97 VSS.n141 VSS.t22 2292
R98 VSS.n292 VSS.t229 2117.06
R99 VSS.n292 VSS.t150 2103.79
R100 VSS.t96 VSS.t70 1980.39
R101 VSS.t34 VSS.t216 1956.78
R102 VSS.t235 VSS.t210 1956.78
R103 VSS.t43 VSS.t213 1953.87
R104 VSS.t93 VSS.t30 1953.87
R105 VSS.n141 VSS.t209 1748.51
R106 VSS.n246 VSS.t165 1720.99
R107 VSS.t168 VSS.t184 1694.19
R108 VSS.t185 VSS.t3 1694.19
R109 VSS.t27 VSS.t141 1692.01
R110 VSS.t117 VSS.t121 1692.01
R111 VSS.n196 VSS.n193 1607.58
R112 VSS.n192 VSS.n191 1600.5
R113 VSS.n196 VSS.n195 1597.63
R114 VSS.n168 VSS.t80 1577.93
R115 VSS.n117 VSS.n115 1573.59
R116 VSS.n114 VSS.n113 1405.57
R117 VSS.n249 VSS.n248 1385.25
R118 VSS.n132 VSS.t89 1348.12
R119 VSS.n191 VSS.n190 1282.2
R120 VSS.n24 VSS.t158 1199.47
R121 VSS.t152 VSS.n294 1199.47
R122 VSS.n190 VSS.t162 1199.47
R123 VSS.n246 VSS.t138 1170.91
R124 VSS.n293 VSS.t143 1153.78
R125 VSS.t176 VSS.n142 1153.78
R126 VSS.n158 VSS.n157 1119.51
R127 VSS.t160 VSS.n132 1083.78
R128 VSS.n107 VSS.t101 927.717
R129 VSS.n113 VSS.t190 919.253
R130 VSS.n100 VSS.t118 919.253
R131 VSS.t144 VSS.t183 913.885
R132 VSS.t81 VSS.t225 913.885
R133 VSS.t54 VSS.t206 913.885
R134 VSS.t175 VSS.t87 913.885
R135 VSS.n107 VSS.n106 879.836
R136 VSS.n192 VSS.t147 854.362
R137 VSS.n87 VSS.n57 842.777
R138 VSS.n119 VSS.n118 839.716
R139 VSS.n7 VSS.t227 815.13
R140 VSS.t85 VSS.t111 784.314
R141 VSS.t180 VSS.t230 784.314
R142 VSS.t82 VSS.t67 774.963
R143 VSS.t210 VSS.t90 774.963
R144 VSS.t84 VSS.t4 773.811
R145 VSS.t226 VSS.t93 773.811
R146 VSS.n195 VSS.t233 771.441
R147 VSS.n96 VSS.t112 753.193
R148 VSS.t193 VSS.n114 709.049
R149 VSS.t181 VSS.n25 677.995
R150 VSS.n105 VSS.n65 676.096
R151 VSS.n106 VSS.n61 673.139
R152 VSS.t184 VSS.t142 670.968
R153 VSS.t86 VSS.t49 670.968
R154 VSS.t141 VSS.t61 670.104
R155 VSS.t83 VSS.t50 670.104
R156 VSS.n45 VSS.n44 629.365
R157 VSS.n228 VSS.n227 629.365
R158 VSS.n42 VSS.n41 626.053
R159 VSS.n220 VSS.n219 626.053
R160 VSS.n198 VSS.n197 616.962
R161 VSS.n204 VSS.n203 616.962
R162 VSS.n52 VSS.n51 615.048
R163 VSS.n212 VSS.n211 615.048
R164 VSS.n13 VSS.t143 548.331
R165 VSS.n18 VSS.t71 548.331
R166 VSS.n19 VSS.t38 548.331
R167 VSS.n23 VSS.t183 548.331
R168 VSS.t80 VSS.n167 548.331
R169 VSS.t44 VSS.n166 548.331
R170 VSS.t75 VSS.n165 548.331
R171 VSS.n189 VSS.t54 548.331
R172 VSS.n188 VSS.t21 548.331
R173 VSS.n187 VSS.t116 548.331
R174 VSS.n186 VSS.t205 548.331
R175 VSS.n143 VSS.t176 548.331
R176 VSS.n148 VSS.t215 548.331
R177 VSS.n149 VSS.t74 548.331
R178 VSS.n154 VSS.t87 548.331
R179 VSS.n47 VSS.n45 484.921
R180 VSS.t229 VSS.n291 470.589
R181 VSS.t70 VSS.n290 470.589
R182 VSS.n10 VSS.t85 470.589
R183 VSS.n11 VSS.t180 470.589
R184 VSS.n197 VSS.n196 468.62
R185 VSS.t209 VSS.n140 464.978
R186 VSS.t216 VSS.n139 464.978
R187 VSS.n134 VSS.t82 464.978
R188 VSS.t90 VSS.n133 464.978
R189 VSS.t89 VSS.n2 464.286
R190 VSS.n3 VSS.t43 464.286
R191 VSS.n4 VSS.t84 464.286
R192 VSS.n5 VSS.t226 464.286
R193 VSS.t11 VSS.n57 457.224
R194 VSS.n49 VSS.n42 455
R195 VSS.n204 VSS.n55 448.392
R196 VSS.n251 VSS.n250 434.096
R197 VSS.n51 VSS.n50 430.197
R198 VSS.n212 VSS.n50 426.837
R199 VSS.n155 VSS.n58 420.916
R200 VSS.t142 VSS.n273 402.582
R201 VSS.n274 VSS.t86 402.582
R202 VSS.t3 VSS.n278 402.582
R203 VSS.n279 VSS.t179 402.582
R204 VSS.t61 VSS.n237 402.062
R205 VSS.n238 VSS.t83 402.062
R206 VSS.n241 VSS.t117 402.062
R207 VSS.t138 VSS.n245 402.062
R208 VSS.n173 VSS.t58 372.873
R209 VSS.n13 VSS.t62 365.555
R210 VSS.t109 VSS.n18 365.555
R211 VSS.n19 VSS.t200 365.555
R212 VSS.t158 VSS.n23 365.555
R213 VSS.n167 VSS.t219 365.555
R214 VSS.n166 VSS.t5 365.555
R215 VSS.n165 VSS.t223 365.555
R216 VSS.n295 VSS.t152 365.555
R217 VSS.t162 VSS.n189 365.555
R218 VSS.t128 VSS.n188 365.555
R219 VSS.t51 VSS.n187 365.555
R220 VSS.t55 VSS.n186 365.555
R221 VSS.n143 VSS.t104 365.555
R222 VSS.t68 VSS.n148 365.555
R223 VSS.n149 VSS.t0 365.555
R224 VSS.t154 VSS.n154 365.555
R225 VSS.n108 VSS.n107 347.168
R226 VSS.t136 VSS.t198 337.038
R227 VSS.t139 VSS.t41 337.038
R228 VSS.t88 VSS.t207 335.264
R229 VSS.t99 VSS.t188 335.264
R230 VSS.t9 VSS.t94 330.394
R231 VSS.t39 VSS.t221 330.394
R232 VSS.t177 VSS.t32 329.37
R233 VSS.t16 VSS.t131 329.37
R234 VSS.n291 VSS.t96 313.726
R235 VSS.n290 VSS.t36 313.726
R236 VSS.n10 VSS.t78 313.726
R237 VSS.t145 VSS.n11 313.726
R238 VSS.n140 VSS.t34 309.986
R239 VSS.n139 VSS.t72 309.986
R240 VSS.n134 VSS.t235 309.986
R241 VSS.n133 VSS.t160 309.986
R242 VSS.t213 VSS.n2 309.524
R243 VSS.n3 VSS.t76 309.524
R244 VSS.t30 VSS.n4 309.524
R245 VSS.t150 VSS.n5 309.524
R246 VSS.n273 VSS.t165 268.387
R247 VSS.n274 VSS.t168 268.387
R248 VSS.n278 VSS.t64 268.387
R249 VSS.n279 VSS.t185 268.387
R250 VSS.n237 VSS.t147 268.041
R251 VSS.n238 VSS.t27 268.041
R252 VSS.n241 VSS.t18 268.041
R253 VSS.n245 VSS.t121 268.041
R254 VSS.n168 VSS.n158 204.131
R255 VSS.n44 VSS.t136 196.032
R256 VSS.n227 VSS.t139 196.032
R257 VSS.n41 VSS.t88 195
R258 VSS.n219 VSS.t99 195
R259 VSS.n198 VSS.t9 192.168
R260 VSS.n203 VSS.t39 192.168
R261 VSS.n52 VSS.t177 191.572
R262 VSS.n211 VSS.t16 191.572
R263 VSS.n96 VSS.n65 171.989
R264 VSS.t112 VSS.t231 166.059
R265 VSS.n105 VSS.n104 156.642
R266 VSS.n114 VSS.n61 154.197
R267 VSS.n86 VSS.t196 121.806
R268 VSS.n85 VSS.t173 121.806
R269 VSS.n84 VSS.t45 121.806
R270 VSS.n83 VSS.t126 121.806
R271 VSS.n82 VSS.t124 121.806
R272 VSS.n77 VSS.t217 121.806
R273 VSS.t171 VSS.n125 121.806
R274 VSS.n126 VSS.t22 121.806
R275 VSS.n118 VSS.n117 100.334
R276 VSS.t2 VSS.t133 97.6999
R277 VSS.n265 VSS.n263 87.9034
R278 VSS.n118 VSS.t202 74.768
R279 VSS.n115 VSS.t193 72.8445
R280 VSS.n117 VSS.n116 59.271
R281 VSS.n87 VSS.t106 54.3731
R282 VSS.n90 VSS.t11 54.3731
R283 VSS.n104 VSS.t24 52.2145
R284 VSS.n263 VSS.n251 49.2247
R285 VSS.n294 VSS.n293 47.3306
R286 VSS.n263 VSS.n262 34.9528
R287 VSS.n265 VSS.t115 34.8931
R288 VSS.n294 VSS.n7 26.295
R289 VSS.n155 VSS.t91 22.8476
R290 VSS.t115 VSS.t2 21.933
R291 VSS.n25 VSS.n24 21.8713
R292 VSS.n49 VSS.n48 20.5268
R293 VSS.n196 VSS.n55 16.8573
R294 VSS.n106 VSS.n105 13.8894
R295 VSS.n157 VSS.n155 11.424
R296 VSS.n47 VSS.n46 10.318
R297 VSS.n97 VSS.t232 10.2719
R298 VSS.n190 VSS.n173 9.623
R299 VSS VSS.t212 9.43705
R300 VSS.n156 VSS.t92 9.3736
R301 VSS.n6 VSS.t228 9.3736
R302 VSS.n172 VSS.n171 9.37275
R303 VSS.n266 VSS.n32 9.37275
R304 VSS.n199 VSS.t95 9.3533
R305 VSS.n40 VSS.t208 9.3533
R306 VSS.n218 VSS.t189 9.3533
R307 VSS.n43 VSS.t199 9.35181
R308 VSS.n226 VSS.t42 9.35181
R309 VSS.n88 VSS.n68 9.33837
R310 VSS.n95 VSS.n93 9.3221
R311 VSS.n202 VSS.t222 9.31766
R312 VSS.n53 VSS.t33 9.31744
R313 VSS.n210 VSS.t132 9.31744
R314 VSS.n56 VSS.t234 9.30652
R315 VSS.n281 VSS.t182 9.30652
R316 VSS.n120 VSS.n59 9.30652
R317 VSS.n111 VSS.n110 9.30652
R318 VSS.n109 VSS.n62 9.30652
R319 VSS.n70 VSS.t197 9.30518
R320 VSS.n72 VSS.t174 9.30518
R321 VSS.n74 VSS.t46 9.30518
R322 VSS.n76 VSS.t127 9.30518
R323 VSS.n80 VSS.t125 9.30518
R324 VSS.n78 VSS.t218 9.30518
R325 VSS.n123 VSS.t172 9.30518
R326 VSS.n128 VSS.t23 9.30518
R327 VSS.n102 VSS.n99 9.28776
R328 VSS.n64 VSS.n63 9.26757
R329 VSS.n92 VSS.n66 9.26488
R330 VSS.n89 VSS.n67 9.26488
R331 VSS.n131 VSS.t35 7.19156
R332 VSS.n137 VSS.t73 7.19156
R333 VSS.n243 VSS.n33 7.19156
R334 VSS.n240 VSS.n34 7.19156
R335 VSS.n184 VSS.n183 7.19156
R336 VSS.n181 VSS.n180 7.19156
R337 VSS.n178 VSS.n177 7.19156
R338 VSS.n260 VSS.n259 7.19156
R339 VSS.n257 VSS.n256 7.19156
R340 VSS.n254 VSS.n253 7.19156
R341 VSS.n27 VSS.n26 7.19156
R342 VSS.n276 VSS.n28 7.19156
R343 VSS.n15 VSS.t63 7.19156
R344 VSS.n16 VSS.t110 7.19156
R345 VSS.n21 VSS.t201 7.19156
R346 VSS.n306 VSS.t214 7.19156
R347 VSS.n304 VSS.t77 7.19156
R348 VSS.n160 VSS.t220 7.19156
R349 VSS.n162 VSS.t6 7.19156
R350 VSS.n163 VSS.t224 7.19156
R351 VSS.n145 VSS.t105 7.19156
R352 VSS.n146 VSS.t69 7.19156
R353 VSS.n151 VSS.t1 7.19156
R354 VSS.n9 VSS.t97 7.17823
R355 VSS.n288 VSS.t37 7.17823
R356 VSS.n230 VSS.t137 7.14823
R357 VSS.n231 VSS.t140 7.14823
R358 VSS.n206 VSS.t10 7.13989
R359 VSS.n222 VSS.t98 7.13989
R360 VSS.n223 VSS.t100 7.13989
R361 VSS.n207 VSS.t40 7.13989
R362 VSS.n214 VSS.t178 7.12156
R363 VSS.n215 VSS.t17 7.12156
R364 VSS.n104 VSS.n103 6.82037
R365 VSS.n122 VSS.n121 6.06679
R366 VSS.n135 VSS.t236 5.91399
R367 VSS.n309 VSS.t161 5.91399
R368 VSS.n235 VSS.n234 5.91399
R369 VSS.n233 VSS.n35 5.91399
R370 VSS.n175 VSS.n174 5.91399
R371 VSS.n31 VSS.n30 5.91399
R372 VSS.n271 VSS.n270 5.91399
R373 VSS.n269 VSS.n29 5.91399
R374 VSS.n12 VSS.t159 5.91399
R375 VSS.n302 VSS.t31 5.91399
R376 VSS.n300 VSS.t151 5.91399
R377 VSS.n297 VSS.t153 5.91399
R378 VSS.n152 VSS.t155 5.91399
R379 VSS.n286 VSS.t79 5.90065
R380 VSS.n284 VSS.t146 5.90065
R381 VSS.n115 VSS.n60 5.82215
R382 VSS.n273 VSS.n272 5.2005
R383 VSS.n275 VSS.n274 5.2005
R384 VSS.n278 VSS.n277 5.2005
R385 VSS.n280 VSS.n279 5.2005
R386 VSS.n262 VSS.n261 5.2005
R387 VSS.n262 VSS.n258 5.2005
R388 VSS.n262 VSS.n255 5.2005
R389 VSS.n262 VSS.n252 5.2005
R390 VSS.n266 VSS.n265 5.2005
R391 VSS.n23 VSS.n22 5.2005
R392 VSS.n20 VSS.n19 5.2005
R393 VSS.n18 VSS.n17 5.2005
R394 VSS.n14 VSS.n13 5.2005
R395 VSS.n282 VSS.n25 5.2005
R396 VSS.n291 VSS.n8 5.2005
R397 VSS.n290 VSS.n289 5.2005
R398 VSS.n287 VSS.n10 5.2005
R399 VSS.n285 VSS.n11 5.2005
R400 VSS.n167 VSS.n159 5.2005
R401 VSS.n166 VSS.n161 5.2005
R402 VSS.n165 VSS.n164 5.2005
R403 VSS.n296 VSS.n295 5.2005
R404 VSS.n113 VSS.n112 5.2005
R405 VSS.n86 VSS.n69 5.2005
R406 VSS.n85 VSS.n71 5.2005
R407 VSS.n84 VSS.n73 5.2005
R408 VSS.n83 VSS.n75 5.2005
R409 VSS.n82 VSS.n81 5.2005
R410 VSS.n79 VSS.n77 5.2005
R411 VSS.n127 VSS.n126 5.2005
R412 VSS.n125 VSS.n124 5.2005
R413 VSS.n88 VSS.n87 5.2005
R414 VSS.n91 VSS.n90 5.2005
R415 VSS.n101 VSS.n100 5.2005
R416 VSS.n94 VSS.n65 5.2005
R417 VSS.n97 VSS.n96 5.2005
R418 VSS.n195 VSS.n194 5.2005
R419 VSS.n199 VSS.n198 5.2005
R420 VSS.n203 VSS.n202 5.2005
R421 VSS.n205 VSS.n204 5.2005
R422 VSS.n53 VSS.n52 5.2005
R423 VSS.n213 VSS.n212 5.2005
R424 VSS.n211 VSS.n210 5.2005
R425 VSS.n42 VSS.n38 5.2005
R426 VSS.n41 VSS.n40 5.2005
R427 VSS.n221 VSS.n220 5.2005
R428 VSS.n219 VSS.n218 5.2005
R429 VSS.n45 VSS.n37 5.2005
R430 VSS.n44 VSS.n43 5.2005
R431 VSS.n229 VSS.n228 5.2005
R432 VSS.n227 VSS.n226 5.2005
R433 VSS.n173 VSS.n172 5.2005
R434 VSS.n237 VSS.n236 5.2005
R435 VSS.n239 VSS.n238 5.2005
R436 VSS.n242 VSS.n241 5.2005
R437 VSS.n245 VSS.n244 5.2005
R438 VSS.n186 VSS.n185 5.2005
R439 VSS.n187 VSS.n182 5.2005
R440 VSS.n188 VSS.n179 5.2005
R441 VSS.n189 VSS.n176 5.2005
R442 VSS.n7 VSS.n6 5.2005
R443 VSS.n301 VSS.n5 5.2005
R444 VSS.n303 VSS.n4 5.2005
R445 VSS.n305 VSS.n3 5.2005
R446 VSS.n307 VSS.n2 5.2005
R447 VSS.n157 VSS.n156 5.2005
R448 VSS.n144 VSS.n143 5.2005
R449 VSS.n148 VSS.n147 5.2005
R450 VSS.n150 VSS.n149 5.2005
R451 VSS.n154 VSS.n153 5.2005
R452 VSS.n133 VSS.n0 5.2005
R453 VSS.n136 VSS.n134 5.2005
R454 VSS.n139 VSS.n138 5.2005
R455 VSS.n140 VSS.n130 5.2005
R456 VSS.n232 VSS.n231 4.93566
R457 VSS.n129 VSS 2.96937
R458 VSS.n281 VSS 2.19213
R459 VSS.n251 VSS.n247 0.912828
R460 VSS.n268 VSS.n267 0.889398
R461 VSS.n284 VSS.n283 0.889168
R462 VSS.n299 VSS.n298 0.845914
R463 VSS.n308 VSS.n1 0.845914
R464 VSS.n233 VSS.n232 0.817931
R465 VSS.n268 VSS 0.51022
R466 VSS.n236 VSS.n235 0.480225
R467 VSS.n240 VSS.n239 0.480225
R468 VSS.n272 VSS.n271 0.480225
R469 VSS.n276 VSS.n275 0.480225
R470 VSS.n181 VSS 0.343161
R471 VSS.n184 VSS 0.343161
R472 VSS.n243 VSS 0.343161
R473 VSS.n257 VSS 0.343161
R474 VSS.n260 VSS 0.343161
R475 VSS VSS.n27 0.343161
R476 VSS VSS.n15 0.343161
R477 VSS.n16 VSS 0.343161
R478 VSS VSS.n160 0.343161
R479 VSS VSS.n162 0.343161
R480 VSS VSS.n145 0.343161
R481 VSS.n146 VSS 0.343161
R482 VSS VSS.n176 0.289491
R483 VSS VSS.n252 0.289491
R484 VSS.n22 VSS 0.289491
R485 VSS.n296 VSS 0.289491
R486 VSS.n153 VSS 0.289491
R487 VSS.n308 VSS 0.239649
R488 VSS.n299 VSS 0.229454
R489 VSS.n288 VSS.n287 0.203963
R490 VSS.n286 VSS.n285 0.203963
R491 VSS.n137 VSS.n136 0.203963
R492 VSS.n135 VSS.n0 0.203963
R493 VSS.n304 VSS.n303 0.203174
R494 VSS.n302 VSS.n301 0.203174
R495 VSS.n178 VSS 0.191234
R496 VSS.n254 VSS 0.191234
R497 VSS VSS.n21 0.191234
R498 VSS.n163 VSS 0.191234
R499 VSS VSS.n151 0.191234
R500 VSS VSS.n129 0.153185
R501 VSS.n89 VSS 0.152427
R502 VSS.n92 VSS 0.152427
R503 VSS.n109 VSS 0.151087
R504 VSS VSS.n64 0.150362
R505 VSS VSS.n9 0.145831
R506 VSS VSS.n131 0.145831
R507 VSS.n306 VSS 0.145267
R508 VSS.n269 VSS.n268 0.14417
R509 VSS VSS.n111 0.141998
R510 VSS VSS.n1 0.137685
R511 VSS.n298 VSS 0.137685
R512 VSS VSS.n36 0.137136
R513 VSS.n267 VSS 0.137136
R514 VSS.n95 VSS.n94 0.136634
R515 VSS.n283 VSS.n12 0.135964
R516 VSS.n179 VSS.n178 0.118573
R517 VSS.n182 VSS.n181 0.118573
R518 VSS.n185 VSS.n184 0.118573
R519 VSS.n242 VSS.n240 0.118573
R520 VSS.n244 VSS.n243 0.118573
R521 VSS.n255 VSS.n254 0.118573
R522 VSS.n258 VSS.n257 0.118573
R523 VSS.n261 VSS.n260 0.118573
R524 VSS.n277 VSS.n276 0.118573
R525 VSS.n280 VSS.n27 0.118573
R526 VSS.n15 VSS.n14 0.118573
R527 VSS.n17 VSS.n16 0.118573
R528 VSS.n21 VSS.n20 0.118573
R529 VSS.n160 VSS.n159 0.118573
R530 VSS.n162 VSS.n161 0.118573
R531 VSS.n164 VSS.n163 0.118573
R532 VSS.n145 VSS.n144 0.118573
R533 VSS.n147 VSS.n146 0.118573
R534 VSS.n151 VSS.n150 0.118573
R535 VSS VSS.n175 0.115271
R536 VSS VSS.n233 0.115271
R537 VSS.n235 VSS 0.115271
R538 VSS VSS.n31 0.115271
R539 VSS VSS.n269 0.115271
R540 VSS.n271 VSS 0.115271
R541 VSS VSS.n12 0.115271
R542 VSS.n297 VSS 0.115271
R543 VSS VSS.n152 0.115271
R544 VSS.n121 VSS 0.111993
R545 VSS.n209 VSS.n39 0.103269
R546 VSS.n217 VSS.n38 0.103269
R547 VSS.n225 VSS.n37 0.103269
R548 VSS.n175 VSS.n36 0.10206
R549 VSS.n267 VSS.n31 0.10206
R550 VSS.n298 VSS.n297 0.10206
R551 VSS.n152 VSS.n1 0.10206
R552 VSS VSS.n70 0.09225
R553 VSS VSS.n72 0.09225
R554 VSS.n80 VSS 0.09225
R555 VSS.n78 VSS 0.09225
R556 VSS VSS.n74 0.092
R557 VSS.n98 VSS.n95 0.0844496
R558 VSS.n309 VSS.n308 0.0799942
R559 VSS.n300 VSS.n299 0.079686
R560 VSS.n91 VSS.n89 0.0739862
R561 VSS.n103 VSS.n92 0.0739862
R562 VSS.n108 VSS.n64 0.0739862
R563 VSS.n112 VSS.n109 0.066973
R564 VSS.n120 VSS.n119 0.0666983
R565 VSS.n208 VSS.n207 0.0664039
R566 VSS.n216 VSS.n215 0.0637265
R567 VSS.n111 VSS.n60 0.0618793
R568 VSS.n200 VSS.n54 0.061873
R569 VSS.n122 VSS 0.061
R570 VSS.n232 VSS.n36 0.059582
R571 VSS.n102 VSS.n98 0.0540556
R572 VSS VSS.n223 0.053635
R573 VSS.n129 VSS 0.0523288
R574 VSS.n9 VSS.n8 0.0505778
R575 VSS.n289 VSS.n288 0.0505778
R576 VSS.n131 VSS.n130 0.0505778
R577 VSS.n138 VSS.n137 0.0505778
R578 VSS.n307 VSS.n306 0.0503837
R579 VSS.n305 VSS.n304 0.0503837
R580 VSS.n200 VSS 0.0502725
R581 VSS VSS.n286 0.049177
R582 VSS VSS.n284 0.049177
R583 VSS VSS.n135 0.049177
R584 VSS VSS.n309 0.049177
R585 VSS VSS.n302 0.0489884
R586 VSS VSS.n300 0.0489884
R587 VSS VSS.n76 0.04625
R588 VSS VSS.n128 0.0454173
R589 VSS.n70 VSS.n69 0.04525
R590 VSS.n72 VSS.n71 0.04525
R591 VSS.n74 VSS.n73 0.04525
R592 VSS.n76 VSS.n75 0.04525
R593 VSS.n81 VSS.n80 0.04525
R594 VSS.n79 VSS.n78 0.04525
R595 VSS.n124 VSS.n123 0.04525
R596 VSS.n128 VSS.n127 0.04525
R597 VSS.n201 VSS.n200 0.0423182
R598 VSS.n102 VSS.n101 0.032289
R599 VSS.n123 VSS.n122 0.03175
R600 VSS VSS.n201 0.0311818
R601 VSS.n283 VSS 0.030089
R602 VSS.n201 VSS.n56 0.0295323
R603 VSS.n206 VSS 0.0289211
R604 VSS.n214 VSS 0.0289211
R605 VSS.n222 VSS 0.0289211
R606 VSS.n230 VSS 0.0289211
R607 VSS VSS.n102 0.026922
R608 VSS.n121 VSS.n120 0.0255299
R609 VSS.n282 VSS.n281 0.0248493
R610 VSS.n208 VSS 0.0205495
R611 VSS VSS.n209 0.0205495
R612 VSS VSS.n56 0.0135645
R613 VSS.n224 VSS 0.00935583
R614 VSS.n194 VSS 0.00654839
R615 VSS VSS.n179 0.00545413
R616 VSS VSS.n182 0.00545413
R617 VSS.n185 VSS 0.00545413
R618 VSS VSS.n242 0.00545413
R619 VSS.n244 VSS 0.00545413
R620 VSS VSS.n255 0.00545413
R621 VSS VSS.n258 0.00545413
R622 VSS.n261 VSS 0.00545413
R623 VSS.n277 VSS 0.00545413
R624 VSS VSS.n280 0.00545413
R625 VSS.n14 VSS 0.00545413
R626 VSS.n17 VSS 0.00545413
R627 VSS.n20 VSS 0.00545413
R628 VSS.n159 VSS 0.00545413
R629 VSS.n161 VSS 0.00545413
R630 VSS.n164 VSS 0.00545413
R631 VSS.n144 VSS 0.00545413
R632 VSS.n147 VSS 0.00545413
R633 VSS.n150 VSS 0.00545413
R634 VSS.n98 VSS 0.00427778
R635 VSS.n176 VSS 0.00380275
R636 VSS.n236 VSS 0.00380275
R637 VSS.n239 VSS 0.00380275
R638 VSS.n252 VSS 0.00380275
R639 VSS.n272 VSS 0.00380275
R640 VSS.n275 VSS 0.00380275
R641 VSS.n22 VSS 0.00380275
R642 VSS VSS.n296 0.00380275
R643 VSS.n153 VSS 0.00380275
R644 VSS.n94 VSS 0.00352521
R645 VSS.n216 VSS 0.00286842
R646 VSS VSS.n217 0.00286842
R647 VSS.n224 VSS 0.00279299
R648 VSS VSS.n225 0.00279299
R649 VSS.n8 VSS 0.00260117
R650 VSS.n289 VSS 0.00260117
R651 VSS.n130 VSS 0.00260117
R652 VSS.n138 VSS 0.00260117
R653 VSS VSS.n307 0.00259302
R654 VSS VSS.n305 0.00259302
R655 VSS.n156 VSS 0.00219811
R656 VSS.n6 VSS 0.00219811
R657 VSS.n172 VSS 0.00219811
R658 VSS VSS.n266 0.00219811
R659 VSS.n287 VSS 0.00190078
R660 VSS.n285 VSS 0.00190078
R661 VSS.n136 VSS 0.00190078
R662 VSS VSS.n0 0.00190078
R663 VSS.n303 VSS 0.00189535
R664 VSS.n301 VSS 0.00189535
R665 VSS VSS.n199 0.00168421
R666 VSS.n40 VSS 0.00168421
R667 VSS.n218 VSS 0.00168421
R668 VSS.n43 VSS 0.0016465
R669 VSS.n226 VSS 0.0016465
R670 VSS VSS.n88 0.00132569
R671 VSS VSS.n91 0.00132569
R672 VSS.n103 VSS 0.00132569
R673 VSS.n101 VSS 0.00132569
R674 VSS VSS.n108 0.00132569
R675 VSS.n112 VSS 0.00124689
R676 VSS.n119 VSS 0.0012438
R677 VSS.n60 VSS 0.00118965
R678 VSS VSS.n205 0.00111785
R679 VSS VSS.n213 0.00111785
R680 VSS VSS.n221 0.00111785
R681 VSS VSS.n229 0.00111785
R682 VSS VSS.n282 0.00111644
R683 VSS.n69 VSS 0.001
R684 VSS.n71 VSS 0.001
R685 VSS.n73 VSS 0.001
R686 VSS.n75 VSS 0.001
R687 VSS.n81 VSS 0.001
R688 VSS VSS.n79 0.001
R689 VSS.n124 VSS 0.001
R690 VSS.n127 VSS 0.001
R691 VSS.n194 VSS 0.000983871
R692 VSS.n202 VSS 0.000954545
R693 VSS VSS.n53 0.000945545
R694 VSS.n210 VSS 0.000945545
R695 VSS VSS.n97 0.000944444
R696 VSS.n205 VSS.n54 0.00070595
R697 VSS.n207 VSS.n206 0.00070595
R698 VSS.n209 VSS.n208 0.00070595
R699 VSS.n213 VSS.n39 0.00070595
R700 VSS.n215 VSS.n214 0.00070595
R701 VSS.n217 VSS.n216 0.00070595
R702 VSS.n221 VSS.n38 0.00070595
R703 VSS.n223 VSS.n222 0.00070595
R704 VSS.n225 VSS.n224 0.00070595
R705 VSS.n229 VSS.n37 0.00070595
R706 VSS.n231 VSS.n230 0.00070595
R707 VDD.n143 VDD.t190 13882.6
R708 VDD.n95 VDD.t188 13882.6
R709 VDD.n125 VDD.t55 12382.6
R710 VDD.n92 VDD.t262 12382.6
R711 VDD.n249 VDD.n248 11185.2
R712 VDD.n89 VDD.t47 7208.33
R713 VDD.n120 VDD.t81 7041.67
R714 VDD.t129 VDD.t118 961.905
R715 VDD.t248 VDD.t298 961.905
R716 VDD.t335 VDD.n114 848.615
R717 VDD.n115 VDD.t274 809.492
R718 VDD.t88 VDD.t330 765.152
R719 VDD.t140 VDD.t8 765.152
R720 VDD.t147 VDD.t337 765.152
R721 VDD.t224 VDD.t305 765.152
R722 VDD.t99 VDD.t60 765.152
R723 VDD.t105 VDD.t210 765.152
R724 VDD.t67 VDD.t229 765.152
R725 VDD.t102 VDD.t57 765.152
R726 VDD.t217 VDD.t212 765.152
R727 VDD.t52 VDD.t207 765.152
R728 VDD.t96 VDD.t123 765.152
R729 VDD.t44 VDD.t2 765.152
R730 VDD.t250 VDD.t280 765.152
R731 VDD.t93 VDD.t120 765.152
R732 VDD.t283 VDD.t4 765.152
R733 VDD.t132 VDD.t186 765.152
R734 VDD.t200 VDD.t76 765.152
R735 VDD.t347 VDD.t145 765.152
R736 VDD.t85 VDD.t320 765.152
R737 VDD.t6 VDD.t143 765.152
R738 VDD.t182 VDD.t70 765.152
R739 VDD.t325 VDD.t195 765.152
R740 VDD.t127 VDD.t137 765.152
R741 VDD.t257 VDD.t0 765.152
R742 VDD.t322 VDD.t74 765.152
R743 VDD.t125 VDD.t135 765.152
R744 VDD.t312 VDD.t359 765.152
R745 VDD.n248 VDD.t202 676.191
R746 VDD.t300 VDD.t253 536.798
R747 VDD.t49 VDD.t294 501.002
R748 VDD.t255 VDD.t64 501.002
R749 VDD.t214 VDD.t91 501.002
R750 VDD.n249 VDD.t25 485.714
R751 VDD VDD.n95 451.327
R752 VDD.n143 VDD 448.709
R753 VDD VDD.n92 445.577
R754 VDD VDD.n125 442.993
R755 VDD VDD.n89 431.3
R756 VDD VDD.n199 429.187
R757 VDD VDD.n364 429.187
R758 VDD VDD.n120 428.8
R759 VDD.n82 VDD 427.092
R760 VDD VDD.n178 426.699
R761 VDD VDD.n227 426.699
R762 VDD.t269 VDD.n249 426.44
R763 VDD VDD.n86 425.019
R764 VDD.n199 VDD.t35 386.365
R765 VDD.t21 VDD.n178 386.365
R766 VDD.t31 VDD.n227 386.365
R767 VDD.n364 VDD.t28 386.365
R768 VDD.t271 VDD.t248 380.952
R769 VDD.t314 VDD.n143 378.788
R770 VDD.n125 VDD.t332 378.788
R771 VDD.n120 VDD.t176 378.788
R772 VDD.t110 VDD.n86 378.788
R773 VDD.t349 VDD.n89 378.788
R774 VDD.t165 VDD.n92 378.788
R775 VDD.t277 VDD.n95 378.788
R776 VDD.n36 VDD.t192 362.8
R777 VDD.n38 VDD.t220 362.8
R778 VDD.n40 VDD.t288 359.49
R779 VDD.n12 VDD.t328 359.49
R780 VDD.t204 VDD.n82 309.341
R781 VDD.t342 VDD.t147 303.031
R782 VDD.t305 VDD.t116 303.031
R783 VDD.t229 VDD.t108 303.031
R784 VDD.t152 VDD.t102 303.031
R785 VDD.t207 VDD.t241 303.031
R786 VDD.t280 VDD.t232 303.031
R787 VDD.t163 VDD.t93 303.031
R788 VDD.t160 VDD.t200 303.031
R789 VDD.t266 VDD.t347 303.031
R790 VDD.t157 VDD.t6 303.031
R791 VDD.t352 VDD.t182 303.031
R792 VDD.t168 VDD.t257 303.031
R793 VDD.t154 VDD.t125 303.031
R794 VDD.t179 VDD.t312 303.031
R795 VDD.n13 VDD.t291 296.538
R796 VDD.n248 VDD.t78 285.714
R797 VDD.n230 VDD.t245 242.857
R798 VDD.n236 VDD.t129 242.857
R799 VDD.t78 VDD.n240 242.857
R800 VDD.n245 VDD.t271 242.857
R801 VDD.t222 VDD.n14 227.456
R802 VDD.n181 VDD.t149 193.183
R803 VDD.n187 VDD.t88 193.183
R804 VDD.n191 VDD.t140 193.183
R805 VDD.n196 VDD.t342 193.183
R806 VDD.n201 VDD.t339 193.183
R807 VDD.n203 VDD.t132 193.183
R808 VDD.n206 VDD.t160 193.183
R809 VDD.n209 VDD.t266 193.183
R810 VDD.n152 VDD.t171 193.183
R811 VDD.n154 VDD.t85 193.183
R812 VDD.n157 VDD.t157 193.183
R813 VDD.n160 VDD.t352 193.183
R814 VDD.n135 VDD.t259 193.183
R815 VDD.n136 VDD.t325 193.183
R816 VDD.n149 VDD.t137 193.183
R817 VDD.n150 VDD.t168 193.183
R818 VDD.n49 VDD.t317 193.183
R819 VDD.n51 VDD.t322 193.183
R820 VDD.n54 VDD.t154 193.183
R821 VDD.n57 VDD.t179 193.183
R822 VDD.n144 VDD.t314 193.183
R823 VDD.n142 VDD.t332 193.183
R824 VDD.n124 VDD.t176 193.183
R825 VDD.n119 VDD.t274 193.183
R826 VDD.n88 VDD.t110 193.183
R827 VDD.n91 VDD.t349 193.183
R828 VDD.n94 VDD.t165 193.183
R829 VDD.n97 VDD.t277 193.183
R830 VDD.t116 VDD.n183 191.288
R831 VDD.t60 VDD.n190 191.288
R832 VDD.t210 VDD.n193 191.288
R833 VDD.n198 VDD.t303 191.288
R834 VDD.t108 VDD.n322 191.288
R835 VDD.n323 VDD.t152 191.288
R836 VDD.t212 VDD.n331 191.288
R837 VDD.n332 VDD.t243 191.288
R838 VDD.t241 VDD.n232 191.288
R839 VDD.t123 VDD.n239 191.288
R840 VDD.t2 VDD.n242 191.288
R841 VDD.n247 VDD.t205 191.288
R842 VDD.t232 VDD.n266 191.288
R843 VDD.n267 VDD.t163 191.288
R844 VDD.t4 VDD.n275 191.288
R845 VDD.n276 VDD.t264 191.288
R846 VDD.n36 VDD.n14 167.588
R847 VDD.t118 VDD.n230 138.095
R848 VDD.t202 VDD.n236 138.095
R849 VDD.t298 VDD.n240 138.095
R850 VDD.t25 VDD.n245 138.095
R851 VDD.n83 VDD.t204 137.826
R852 VDD.n39 VDD.n38 119.706
R853 VDD.n40 VDD.n39 118.614
R854 VDD.n183 VDD.t21 111.743
R855 VDD.n190 VDD.t224 111.743
R856 VDD.n193 VDD.t99 111.743
R857 VDD.n198 VDD.t105 111.743
R858 VDD.n322 VDD.t41 111.743
R859 VDD.n323 VDD.t67 111.743
R860 VDD.n331 VDD.t57 111.743
R861 VDD.n332 VDD.t217 111.743
R862 VDD.n232 VDD.t31 111.743
R863 VDD.n239 VDD.t52 111.743
R864 VDD.n242 VDD.t96 111.743
R865 VDD.n247 VDD.t44 111.743
R866 VDD.n266 VDD.t17 111.743
R867 VDD.n267 VDD.t250 111.743
R868 VDD.n275 VDD.t120 111.743
R869 VDD.n276 VDD.t283 111.743
R870 VDD.t330 VDD.n181 109.849
R871 VDD.t8 VDD.n187 109.849
R872 VDD.t337 VDD.n191 109.849
R873 VDD.t35 VDD.n196 109.849
R874 VDD.t186 VDD.n201 109.849
R875 VDD.t76 VDD.n203 109.849
R876 VDD.t145 VDD.n206 109.849
R877 VDD.n209 VDD.t14 109.849
R878 VDD.t320 VDD.n152 109.849
R879 VDD.t143 VDD.n154 109.849
R880 VDD.t70 VDD.n157 109.849
R881 VDD.n160 VDD.t38 109.849
R882 VDD.t195 VDD.n135 109.849
R883 VDD.n136 VDD.t127 109.849
R884 VDD.t0 VDD.n149 109.849
R885 VDD.t28 VDD.n150 109.849
R886 VDD.t74 VDD.n49 109.849
R887 VDD.t135 VDD.n51 109.849
R888 VDD.t359 VDD.n54 109.849
R889 VDD.n57 VDD.t11 109.849
R890 VDD.n144 VDD.t239 109.849
R891 VDD.t190 VDD.n142 109.849
R892 VDD.t55 VDD.n124 109.849
R893 VDD.t81 VDD.n119 109.849
R894 VDD.t47 VDD.n88 109.849
R895 VDD.t262 VDD.n91 109.849
R896 VDD.t188 VDD.n94 109.849
R897 VDD.n97 VDD.t237 109.849
R898 VDD.n83 VDD.t310 107.198
R899 VDD.n13 VDD.n12 100.365
R900 VDD.n143 VDD.t83 65.4455
R901 VDD.n125 VDD.t286 64.6
R902 VDD.n95 VDD.t296 62.8277
R903 VDD.n120 VDD.t227 62.5005
R904 VDD.n178 VDD.t113 62.1896
R905 VDD.n227 VDD.t234 62.1896
R906 VDD.n92 VDD.t308 62.016
R907 VDD.n89 VDD.t72 60.0005
R908 VDD.n199 VDD.t345 59.702
R909 VDD.n364 VDD.t174 59.702
R910 VDD.n82 VDD.t355 59.4064
R911 VDD.n86 VDD.t184 59.1138
R912 VDD.n39 VDD.n14 47.8826
R913 VDD.n312 VDD.t40 30.9379
R914 VDD.n314 VDD.t20 30.9379
R915 VDD.n256 VDD.t16 30.9379
R916 VDD.n257 VDD.t30 30.9379
R917 VDD.n210 VDD.t24 30.9379
R918 VDD.n212 VDD.t13 30.9379
R919 VDD.n161 VDD.t34 30.9379
R920 VDD.n163 VDD.t37 30.9379
R921 VDD.n60 VDD.t10 30.9379
R922 VDD.n58 VDD.t27 30.9379
R923 VDD.n45 VDD.t291 28.139
R924 VDD.t253 VDD.n45 28.139
R925 VDD.n46 VDD.t300 28.139
R926 VDD.n46 VDD.t62 28.139
R927 VDD.n312 VDD.t363 24.5101
R928 VDD.n314 VDD.t373 24.5101
R929 VDD.n256 VDD.t374 24.5101
R930 VDD.n257 VDD.t368 24.5101
R931 VDD.n210 VDD.t371 24.5101
R932 VDD.n212 VDD.t362 24.5101
R933 VDD.n161 VDD.t366 24.5101
R934 VDD.n163 VDD.t365 24.5101
R935 VDD.n60 VDD.t372 24.5101
R936 VDD.n58 VDD.t367 24.5101
R937 VDD.n18 VDD.t197 22.0446
R938 VDD.t294 VDD.n23 22.0446
R939 VDD.n24 VDD.t49 22.0446
R940 VDD.n25 VDD.t255 22.0446
R941 VDD.t64 VDD.n16 22.0446
R942 VDD.t91 VDD.n31 22.0446
R943 VDD.n32 VDD.t214 21.0426
R944 VDD.n33 VDD.t222 21.0426
R945 VDD.n39 VDD.n13 18.2487
R946 VDD VDD.t269 10.5649
R947 VDD.n137 VDD.t84 6.62407
R948 VDD.n266 VDD.n265 6.3005
R949 VDD.n268 VDD.n267 6.3005
R950 VDD.n275 VDD.n274 6.3005
R951 VDD.n277 VDD.n276 6.3005
R952 VDD.n216 VDD.n209 6.3005
R953 VDD.n219 VDD.n206 6.3005
R954 VDD.n222 VDD.n203 6.3005
R955 VDD.n225 VDD.n201 6.3005
R956 VDD.n299 VDD.n232 6.3005
R957 VDD.n292 VDD.n239 6.3005
R958 VDD.n287 VDD.n242 6.3005
R959 VDD.n281 VDD.n247 6.3005
R960 VDD.n284 VDD.n245 6.3005
R961 VDD.n291 VDD.n240 6.3005
R962 VDD.n296 VDD.n236 6.3005
R963 VDD.n302 VDD.n230 6.3005
R964 VDD.n322 VDD.n321 6.3005
R965 VDD.n324 VDD.n323 6.3005
R966 VDD.n331 VDD.n330 6.3005
R967 VDD.n333 VDD.n332 6.3005
R968 VDD.n167 VDD.n160 6.3005
R969 VDD.n170 VDD.n157 6.3005
R970 VDD.n173 VDD.n154 6.3005
R971 VDD.n176 VDD.n152 6.3005
R972 VDD.n356 VDD.n183 6.3005
R973 VDD.n349 VDD.n190 6.3005
R974 VDD.n344 VDD.n193 6.3005
R975 VDD.n338 VDD.n198 6.3005
R976 VDD.n341 VDD.n196 6.3005
R977 VDD.n348 VDD.n191 6.3005
R978 VDD.n353 VDD.n187 6.3005
R979 VDD.n359 VDD.n181 6.3005
R980 VDD.n366 VDD.n150 6.3005
R981 VDD VDD.n18 6.3005
R982 VDD.n23 VDD 6.3005
R983 VDD.n24 VDD 6.3005
R984 VDD VDD.n25 6.3005
R985 VDD VDD.n16 6.3005
R986 VDD.n31 VDD 6.3005
R987 VDD.n32 VDD 6.3005
R988 VDD VDD.n33 6.3005
R989 VDD.n38 VDD 6.3005
R990 VDD VDD.n36 6.3005
R991 VDD.n73 VDD.n49 6.3005
R992 VDD.n70 VDD.n51 6.3005
R993 VDD.n67 VDD.n54 6.3005
R994 VDD.n64 VDD.n57 6.3005
R995 VDD.n98 VDD.n97 6.3005
R996 VDD.n102 VDD.n94 6.3005
R997 VDD.n106 VDD.n91 6.3005
R998 VDD.n110 VDD.n88 6.3005
R999 VDD.n84 VDD.n83 6.3005
R1000 VDD.n114 VDD 6.3005
R1001 VDD VDD.n115 6.3005
R1002 VDD.n119 VDD.n118 6.3005
R1003 VDD.n124 VDD.n123 6.3005
R1004 VDD.n135 VDD.n134 6.3005
R1005 VDD.n142 VDD.n141 6.3005
R1006 VDD.n149 VDD.n148 6.3005
R1007 VDD.n140 VDD.n136 6.3005
R1008 VDD.n145 VDD.n144 6.3005
R1009 VDD.n113 VDD 6.18684
R1010 VDD.n279 VDD.t270 5.85907
R1011 VDD.n336 VDD.t346 5.85907
R1012 VDD.n361 VDD.n179 5.85007
R1013 VDD.n304 VDD.n228 5.85007
R1014 VDD VDD.t238 5.1878
R1015 VDD VDD.n19 5.1552
R1016 VDD VDD.t56 5.1508
R1017 VDD.n358 VDD.n182 5.13287
R1018 VDD.n351 VDD.n188 5.13287
R1019 VDD.n347 VDD.t61 5.13287
R1020 VDD.n345 VDD.n192 5.13287
R1021 VDD.n342 VDD.t211 5.13287
R1022 VDD.n340 VDD.n197 5.13287
R1023 VDD.n337 VDD.t304 5.13287
R1024 VDD.n301 VDD.n231 5.13287
R1025 VDD.n294 VDD.n237 5.13287
R1026 VDD.n290 VDD.t124 5.13287
R1027 VDD.n288 VDD.n241 5.13287
R1028 VDD.n285 VDD.t3 5.13287
R1029 VDD.n283 VDD.n246 5.13287
R1030 VDD.n280 VDD.t206 5.13287
R1031 VDD.n261 VDD.n255 5.13287
R1032 VDD.n254 VDD.n253 5.13287
R1033 VDD.n270 VDD.n250 5.13287
R1034 VDD.n273 VDD.t5 5.13287
R1035 VDD.n272 VDD.n271 5.13287
R1036 VDD.n278 VDD.t265 5.13287
R1037 VDD.n282 VDD.t26 5.13287
R1038 VDD.n289 VDD.t299 5.13287
R1039 VDD.n293 VDD.n238 5.13287
R1040 VDD.n295 VDD.t203 5.13287
R1041 VDD.n298 VDD.n233 5.13287
R1042 VDD.n300 VDD.t119 5.13287
R1043 VDD.n303 VDD.n229 5.13287
R1044 VDD.n215 VDD.t15 5.13287
R1045 VDD.n218 VDD.t146 5.13287
R1046 VDD.n221 VDD.t77 5.13287
R1047 VDD.n223 VDD.n202 5.13287
R1048 VDD.n224 VDD.t187 5.13287
R1049 VDD.n226 VDD.n200 5.13287
R1050 VDD.n317 VDD.n311 5.13287
R1051 VDD.n310 VDD.n309 5.13287
R1052 VDD.n326 VDD.n306 5.13287
R1053 VDD.n329 VDD.t213 5.13287
R1054 VDD.n328 VDD.n327 5.13287
R1055 VDD.n334 VDD.t244 5.13287
R1056 VDD.n339 VDD.t36 5.13287
R1057 VDD.n346 VDD.t338 5.13287
R1058 VDD.n350 VDD.n189 5.13287
R1059 VDD.n352 VDD.t9 5.13287
R1060 VDD.n355 VDD.n184 5.13287
R1061 VDD.n357 VDD.t331 5.13287
R1062 VDD.n360 VDD.n180 5.13287
R1063 VDD.n166 VDD.t39 5.13287
R1064 VDD.n169 VDD.t71 5.13287
R1065 VDD.n172 VDD.t144 5.13287
R1066 VDD.n174 VDD.n153 5.13287
R1067 VDD.n175 VDD.t321 5.13287
R1068 VDD.n177 VDD.n151 5.13287
R1069 VDD.n365 VDD.t29 5.13287
R1070 VDD.n63 VDD.t12 5.13287
R1071 VDD.n66 VDD.t360 5.13287
R1072 VDD.n69 VDD.t136 5.13287
R1073 VDD.n71 VDD.n50 5.13287
R1074 VDD.n72 VDD.t75 5.13287
R1075 VDD.n74 VDD.n48 5.13287
R1076 VDD.n99 VDD.n96 5.13287
R1077 VDD.n101 VDD.t189 5.13287
R1078 VDD.n103 VDD.n93 5.13287
R1079 VDD.n105 VDD.t263 5.13287
R1080 VDD.n107 VDD.n90 5.13287
R1081 VDD.n109 VDD.t48 5.13287
R1082 VDD.n111 VDD.n87 5.13287
R1083 VDD.n117 VDD.n79 5.13287
R1084 VDD.n78 VDD.t82 5.13287
R1085 VDD.n122 VDD.n77 5.13287
R1086 VDD.n133 VDD.t196 5.13287
R1087 VDD.n127 VDD.n126 5.13287
R1088 VDD.n139 VDD.t191 5.13287
R1089 VDD.n3 VDD.n2 5.13287
R1090 VDD.n138 VDD.t128 5.13287
R1091 VDD.n6 VDD.n5 5.13287
R1092 VDD.n147 VDD.n4 5.13287
R1093 VDD.n368 VDD.t240 5.13287
R1094 VDD.n146 VDD.t1 5.13287
R1095 VDD VDD.t287 5.10366
R1096 VDD.n22 VDD.t295 5.09836
R1097 VDD.n21 VDD.n20 5.09836
R1098 VDD.n26 VDD.t256 5.09836
R1099 VDD.n27 VDD.n17 5.09836
R1100 VDD.n30 VDD.t92 5.09836
R1101 VDD.n29 VDD.n28 5.09836
R1102 VDD.n34 VDD.t223 5.09836
R1103 VDD.n35 VDD.n15 5.09836
R1104 VDD.n37 VDD.t221 5.09836
R1105 VDD.n11 VDD.n10 5.09836
R1106 VDD.n42 VDD.t329 5.09836
R1107 VDD.n43 VDD.n9 5.09836
R1108 VDD.n44 VDD.t254 5.09836
R1109 VDD.n8 VDD.n7 5.09836
R1110 VDD.n47 VDD.t63 5.09836
R1111 VDD.n363 VDD.t175 5.09407
R1112 VDD.n100 VDD.t297 5.09407
R1113 VDD.n104 VDD.t309 5.09407
R1114 VDD.n108 VDD.t73 5.09407
R1115 VDD.n112 VDD.t185 5.09407
R1116 VDD.n81 VDD.t356 5.09407
R1117 VDD.n80 VDD.t358 5.09407
R1118 VDD.n116 VDD.t336 5.09407
R1119 VDD.n121 VDD.t228 5.09407
R1120 VDD.n33 VDD.n32 5.01052
R1121 VDD.n132 VDD.n131 4.97242
R1122 VDD.n75 VDD.n47 4.93241
R1123 VDD.n114 VDD.t357 4.26489
R1124 VDD.n115 VDD.t335 4.26489
R1125 VDD.n85 VDD.t311 4.12326
R1126 VDD.n164 VDD.n163 4.08741
R1127 VDD VDD.n256 4.08362
R1128 VDD.n211 VDD.n210 4.07437
R1129 VDD.n61 VDD.n60 4.07346
R1130 VDD.n213 VDD.n212 4.06995
R1131 VDD.n162 VDD.n161 4.06354
R1132 VDD VDD.n312 4.0592
R1133 VDD.n59 VDD.n58 4.05141
R1134 VDD.n315 VDD.n314 4.04913
R1135 VDD.n23 VDD.n18 4.00852
R1136 VDD.n25 VDD.n24 4.00852
R1137 VDD.n31 VDD.n16 4.00852
R1138 VDD.n258 VDD.n257 4.0005
R1139 VDD.n41 VDD.n40 3.1505
R1140 VDD.n41 VDD.n12 3.1505
R1141 VDD.n45 VDD 3.1505
R1142 VDD VDD.n46 3.1505
R1143 VDD.n214 VDD.n211 3.06712
R1144 VDD.n165 VDD.n162 3.0645
R1145 VDD.n316 VDD.n315 3.00562
R1146 VDD.n62 VDD.n59 2.95066
R1147 VDD.n165 VDD.n164 2.92128
R1148 VDD.n260 VDD.n259 2.91332
R1149 VDD.n354 VDD.n186 2.85787
R1150 VDD.n297 VDD.n235 2.85787
R1151 VDD.n264 VDD.n263 2.85787
R1152 VDD.n269 VDD.n252 2.85787
R1153 VDD.n286 VDD.n244 2.85787
R1154 VDD.n217 VDD.n208 2.85787
R1155 VDD.n220 VDD.n205 2.85787
R1156 VDD.n320 VDD.n319 2.85787
R1157 VDD.n325 VDD.n308 2.85787
R1158 VDD.n343 VDD.n195 2.85787
R1159 VDD.n168 VDD.n159 2.85787
R1160 VDD.n171 VDD.n156 2.85787
R1161 VDD.n65 VDD.n56 2.85787
R1162 VDD.n68 VDD.n53 2.85787
R1163 VDD.n367 VDD.n1 2.85787
R1164 VDD.n214 VDD.n213 2.85553
R1165 VDD.n260 VDD 2.82101
R1166 VDD.n316 VDD.n313 2.8124
R1167 VDD.n62 VDD.n61 2.79396
R1168 VDD.n186 VDD.t117 2.2755
R1169 VDD.n186 VDD.n185 2.2755
R1170 VDD.n235 VDD.t242 2.2755
R1171 VDD.n235 VDD.n234 2.2755
R1172 VDD.n263 VDD.t233 2.2755
R1173 VDD.n263 VDD.n262 2.2755
R1174 VDD.n252 VDD.t164 2.2755
R1175 VDD.n252 VDD.n251 2.2755
R1176 VDD.n244 VDD.t249 2.2755
R1177 VDD.n244 VDD.n243 2.2755
R1178 VDD.n208 VDD.t348 2.2755
R1179 VDD.n208 VDD.n207 2.2755
R1180 VDD.n205 VDD.t201 2.2755
R1181 VDD.n205 VDD.n204 2.2755
R1182 VDD.n319 VDD.t109 2.2755
R1183 VDD.n319 VDD.n318 2.2755
R1184 VDD.n308 VDD.t153 2.2755
R1185 VDD.n308 VDD.n307 2.2755
R1186 VDD.n195 VDD.t148 2.2755
R1187 VDD.n195 VDD.n194 2.2755
R1188 VDD.n159 VDD.t183 2.2755
R1189 VDD.n159 VDD.n158 2.2755
R1190 VDD.n156 VDD.t7 2.2755
R1191 VDD.n156 VDD.n155 2.2755
R1192 VDD.n56 VDD.t313 2.2755
R1193 VDD.n56 VDD.n55 2.2755
R1194 VDD.n53 VDD.t126 2.2755
R1195 VDD.n53 VDD.n52 2.2755
R1196 VDD.n1 VDD.t258 2.2755
R1197 VDD.n1 VDD.n0 2.2755
R1198 VDD.n317 VDD.n316 2.27547
R1199 VDD.n261 VDD.n260 2.27315
R1200 VDD.n166 VDD.n165 2.26966
R1201 VDD.n215 VDD.n214 2.26502
R1202 VDD.n63 VDD.n62 2.26153
R1203 VDD VDD.n41 1.5755
R1204 VDD VDD.n113 1.37899
R1205 VDD VDD.n278 1.21661
R1206 VDD.n305 VDD.n226 1.18347
R1207 VDD.n22 VDD.n21 1.13088
R1208 VDD.n27 VDD.n26 1.13088
R1209 VDD.n30 VDD.n29 1.13083
R1210 VDD.n362 VDD.n177 1.12775
R1211 VDD.n335 VDD.n334 1.12407
R1212 VDD.n130 VDD.n75 0.986314
R1213 VDD VDD.n34 0.886596
R1214 VDD.n132 VDD.n130 0.559447
R1215 VDD.n84 VDD.n81 0.388218
R1216 VDD.n133 VDD.n132 0.279974
R1217 VDD.n264 VDD.n254 0.233919
R1218 VDD.n270 VDD.n269 0.233919
R1219 VDD.n221 VDD.n220 0.233919
R1220 VDD.n218 VDD.n217 0.233919
R1221 VDD.n320 VDD.n310 0.233919
R1222 VDD.n326 VDD.n325 0.233919
R1223 VDD.n172 VDD.n171 0.233919
R1224 VDD.n169 VDD.n168 0.233919
R1225 VDD.n69 VDD.n68 0.233919
R1226 VDD.n66 VDD.n65 0.233919
R1227 VDD.n335 VDD.n305 0.178068
R1228 VDD.n363 VDD.n362 0.162742
R1229 VDD.n273 VDD.n272 0.141016
R1230 VDD.n224 VDD.n223 0.141016
R1231 VDD.n329 VDD.n328 0.141016
R1232 VDD.n175 VDD.n174 0.141016
R1233 VDD.n72 VDD.n71 0.141016
R1234 VDD.n109 VDD 0.126036
R1235 VDD VDD.n78 0.126036
R1236 VDD VDD.n80 0.125632
R1237 VDD.n105 VDD 0.12226
R1238 VDD VDD.n258 0.121547
R1239 VDD.n113 VDD.n85 0.119239
R1240 VDD.n101 VDD 0.11887
R1241 VDD.n85 VDD 0.110164
R1242 VDD.n274 VDD.n273 0.107339
R1243 VDD.n278 VDD.n277 0.107339
R1244 VDD.n226 VDD.n225 0.107339
R1245 VDD.n223 VDD.n222 0.107339
R1246 VDD.n330 VDD.n329 0.107339
R1247 VDD.n334 VDD.n333 0.107339
R1248 VDD.n177 VDD.n176 0.107339
R1249 VDD.n174 VDD.n173 0.107339
R1250 VDD.n74 VDD.n73 0.107339
R1251 VDD.n71 VDD.n70 0.107339
R1252 VDD VDD.n264 0.106758
R1253 VDD.n269 VDD 0.106758
R1254 VDD VDD.n320 0.106758
R1255 VDD.n325 VDD 0.106758
R1256 VDD.n220 VDD 0.106177
R1257 VDD.n217 VDD 0.106177
R1258 VDD.n171 VDD 0.106177
R1259 VDD.n168 VDD 0.106177
R1260 VDD.n68 VDD 0.106177
R1261 VDD.n65 VDD 0.106177
R1262 VDD.n44 VDD.n8 0.102798
R1263 VDD.n43 VDD.n42 0.102778
R1264 VDD.n37 VDD.n11 0.0987707
R1265 VDD.n100 VDD.n99 0.0984239
R1266 VDD.n104 VDD.n103 0.0962255
R1267 VDD.n112 VDD.n111 0.0962255
R1268 VDD.n117 VDD.n116 0.0962255
R1269 VDD.n108 VDD.n107 0.0917202
R1270 VDD.n122 VDD.n121 0.0917202
R1271 VDD.n130 VDD.n129 0.0908448
R1272 VDD VDD.n44 0.0815938
R1273 VDD VDD.n43 0.081125
R1274 VDD.n365 VDD 0.0808411
R1275 VDD.n265 VDD.n261 0.080629
R1276 VDD.n268 VDD.n254 0.080629
R1277 VDD.n219 VDD.n218 0.080629
R1278 VDD.n216 VDD.n215 0.080629
R1279 VDD.n321 VDD.n317 0.080629
R1280 VDD.n324 VDD.n310 0.080629
R1281 VDD.n170 VDD.n169 0.080629
R1282 VDD.n167 VDD.n166 0.080629
R1283 VDD.n67 VDD.n66 0.080629
R1284 VDD.n64 VDD.n63 0.080629
R1285 VDD VDD.n224 0.0794677
R1286 VDD VDD.n221 0.0794677
R1287 VDD VDD.n175 0.0794677
R1288 VDD VDD.n172 0.0794677
R1289 VDD VDD.n72 0.0794677
R1290 VDD VDD.n69 0.0794677
R1291 VDD VDD.n270 0.0788871
R1292 VDD.n272 VDD 0.0788871
R1293 VDD VDD.n326 0.0788871
R1294 VDD.n328 VDD 0.0788871
R1295 VDD.n99 VDD.n98 0.0782465
R1296 VDD.n103 VDD.n102 0.0764633
R1297 VDD.n111 VDD.n110 0.0764633
R1298 VDD.n118 VDD.n117 0.0764633
R1299 VDD.n47 VDD 0.0742915
R1300 VDD.n42 VDD 0.0739434
R1301 VDD VDD.n8 0.0738649
R1302 VDD VDD.n11 0.0735189
R1303 VDD.n107 VDD.n106 0.0728144
R1304 VDD.n123 VDD.n122 0.0728144
R1305 VDD VDD.n81 0.0709717
R1306 VDD VDD.n37 0.0594773
R1307 VDD VDD.n35 0.0591364
R1308 VDD VDD.n22 0.0576804
R1309 VDD.n26 VDD 0.0576804
R1310 VDD VDD.n30 0.0576804
R1311 VDD.n21 VDD 0.0573421
R1312 VDD VDD.n27 0.0573421
R1313 VDD.n34 VDD 0.0571292
R1314 VDD.n29 VDD 0.0567921
R1315 VDD VDD.n101 0.0541697
R1316 VDD VDD.n109 0.0541697
R1317 VDD VDD.n78 0.0541697
R1318 VDD.n129 VDD 0.0523961
R1319 VDD.n129 VDD.n76 0.0518793
R1320 VDD VDD.n105 0.0515917
R1321 VDD.n128 VDD 0.0493571
R1322 VDD.n367 VDD 0.0435288
R1323 VDD.n75 VDD.n74 0.0434677
R1324 VDD.n305 VDD 0.0403112
R1325 VDD VDD.n335 0.0394651
R1326 VDD.n362 VDD 0.0394564
R1327 VDD.n138 VDD 0.0392961
R1328 VDD.n360 VDD.n359 0.038569
R1329 VDD.n338 VDD.n337 0.038569
R1330 VDD.n303 VDD.n302 0.0377135
R1331 VDD.n281 VDD.n280 0.0377135
R1332 VDD.n35 VDD 0.0352326
R1333 VDD.n366 VDD.n365 0.0350961
R1334 VDD VDD.n100 0.0339978
R1335 VDD VDD.n104 0.0332632
R1336 VDD VDD.n112 0.0332632
R1337 VDD.n116 VDD 0.0332632
R1338 VDD.n148 VDD.n3 0.0326553
R1339 VDD.n349 VDD.n348 0.0323621
R1340 VDD VDD.n108 0.0317552
R1341 VDD.n121 VDD 0.0317552
R1342 VDD.n146 VDD.n145 0.0313824
R1343 VDD.n295 VDD.n294 0.0312416
R1344 VDD.n289 VDD.n288 0.0312416
R1345 VDD.n352 VDD.n351 0.0282241
R1346 VDD.n346 VDD.n345 0.0282241
R1347 VDD.n292 VDD.n291 0.0280056
R1348 VDD.n354 VDD.n353 0.0273966
R1349 VDD.n344 VDD.n343 0.0273966
R1350 VDD VDD.n355 0.0271897
R1351 VDD.n342 VDD 0.0269828
R1352 VDD.n300 VDD.n299 0.0267921
R1353 VDD.n284 VDD.n283 0.0267921
R1354 VDD VDD.n301 0.0263876
R1355 VDD.n282 VDD 0.0261854
R1356 VDD.n357 VDD.n356 0.0236724
R1357 VDD.n341 VDD.n340 0.0236724
R1358 VDD VDD.n358 0.0232586
R1359 VDD.n297 VDD.n296 0.0231517
R1360 VDD.n287 VDD.n286 0.0231517
R1361 VDD.n339 VDD 0.0230517
R1362 VDD VDD.n298 0.0229494
R1363 VDD.n351 VDD.n350 0.0228448
R1364 VDD.n347 VDD.n346 0.0228448
R1365 VDD.n285 VDD 0.0227472
R1366 VDD.n76 VDD 0.0222241
R1367 VDD.n128 VDD.n127 0.0214709
R1368 VDD VDD.n363 0.0207439
R1369 VDD.n141 VDD.n6 0.0205971
R1370 VDD.n294 VDD.n293 0.0187022
R1371 VDD.n290 VDD.n289 0.0187022
R1372 VDD VDD.n368 0.0186765
R1373 VDD.n315 VDD 0.0181958
R1374 VDD VDD.n352 0.016431
R1375 VDD.n345 VDD 0.0162241
R1376 VDD.n368 VDD.n367 0.0162059
R1377 VDD.n211 VDD 0.0157113
R1378 VDD.n259 VDD 0.0152541
R1379 VDD.n298 VDD.n297 0.0150618
R1380 VDD.n286 VDD.n285 0.0150618
R1381 VDD VDD.n147 0.0137353
R1382 VDD.n61 VDD 0.0133571
R1383 VDD.n59 VDD 0.0132059
R1384 VDD.n127 VDD.n6 0.0125583
R1385 VDD.n139 VDD.n138 0.0125583
R1386 VDD VDD.n295 0.0124326
R1387 VDD.n288 VDD 0.0122303
R1388 VDD VDD.n139 0.0122087
R1389 VDD.n355 VDD.n354 0.0116724
R1390 VDD.n343 VDD.n342 0.0116724
R1391 VDD VDD.n140 0.0111602
R1392 VDD.n162 VDD 0.0110882
R1393 VDD.n134 VDD.n133 0.0105519
R1394 VDD.n213 VDD 0.00981034
R1395 VDD VDD.n290 0.00980337
R1396 VDD.n293 VDD 0.00960112
R1397 VDD VDD.n80 0.00839474
R1398 VDD.n361 VDD.n360 0.0065
R1399 VDD VDD.n347 0.0062931
R1400 VDD.n337 VDD.n336 0.0062931
R1401 VDD.n350 VDD 0.00608621
R1402 VDD.n358 VDD.n357 0.00587931
R1403 VDD.n340 VDD.n339 0.00587931
R1404 VDD.n313 VDD 0.00579412
R1405 VDD VDD.n84 0.00579412
R1406 VDD.n259 VDD.n258 0.00419863
R1407 VDD.n98 VDD 0.00388028
R1408 VDD.n102 VDD 0.00380275
R1409 VDD.n110 VDD 0.00380275
R1410 VDD.n118 VDD 0.00380275
R1411 VDD.n106 VDD 0.0036441
R1412 VDD.n164 VDD 0.00307143
R1413 VDD.n304 VDD.n303 0.00272472
R1414 VDD.n280 VDD.n279 0.00252247
R1415 VDD VDD.n137 0.00242233
R1416 VDD.n274 VDD 0.00224194
R1417 VDD.n277 VDD 0.00224194
R1418 VDD.n330 VDD 0.00224194
R1419 VDD.n333 VDD 0.00224194
R1420 VDD.n301 VDD.n300 0.00211798
R1421 VDD.n283 VDD.n282 0.00211798
R1422 VDD.n147 VDD.n146 0.00208824
R1423 VDD.n145 VDD 0.00191176
R1424 VDD.n141 VDD 0.00189806
R1425 VDD VDD.n3 0.0017233
R1426 VDD.n129 VDD.n128 0.00166883
R1427 VDD.n134 VDD 0.00166883
R1428 VDD.n225 VDD 0.00166129
R1429 VDD.n222 VDD 0.00166129
R1430 VDD VDD.n219 0.00166129
R1431 VDD VDD.n216 0.00166129
R1432 VDD.n176 VDD 0.00166129
R1433 VDD.n173 VDD 0.00166129
R1434 VDD VDD.n170 0.00166129
R1435 VDD VDD.n167 0.00166129
R1436 VDD.n73 VDD 0.00166129
R1437 VDD.n70 VDD 0.00166129
R1438 VDD VDD.n67 0.00166129
R1439 VDD VDD.n64 0.00166129
R1440 VDD.n313 VDD 0.00155882
R1441 VDD VDD.n349 0.00112069
R1442 VDD VDD.n344 0.00112069
R1443 VDD VDD.n338 0.00112069
R1444 VDD VDD.n292 0.00110674
R1445 VDD VDD.n287 0.00110674
R1446 VDD VDD.n281 0.00110674
R1447 VDD.n265 VDD 0.00108064
R1448 VDD VDD.n268 0.00108064
R1449 VDD.n321 VDD 0.00108064
R1450 VDD VDD.n324 0.00108064
R1451 VDD VDD.n366 0.00100139
R1452 VDD VDD.n361 0.000913793
R1453 VDD.n359 VDD 0.000913793
R1454 VDD.n353 VDD 0.000913793
R1455 VDD.n348 VDD 0.000913793
R1456 VDD VDD.n341 0.000913793
R1457 VDD.n336 VDD 0.000913793
R1458 VDD VDD.n304 0.000904494
R1459 VDD.n302 VDD 0.000904494
R1460 VDD.n296 VDD 0.000904494
R1461 VDD.n291 VDD 0.000904494
R1462 VDD VDD.n284 0.000904494
R1463 VDD.n279 VDD 0.000904494
R1464 VDD.n123 VDD.n76 0.000893013
R1465 VDD.n140 VDD 0.000849515
R1466 VDD.n137 VDD 0.000849515
R1467 VDD.n148 VDD 0.000849515
R1468 VDD.n356 VDD 0.000706897
R1469 VDD.n299 VDD 0.000702247
R1470 RST.n31 RST.t10 36.935
R1471 RST.n22 RST.t8 36.935
R1472 RST.n27 RST.t4 36.935
R1473 RST.n1 RST.t6 36.935
R1474 RST.n13 RST.t11 36.935
R1475 RST.n31 RST.t7 18.1962
R1476 RST.n22 RST.t5 18.1962
R1477 RST.n27 RST.t3 18.1962
R1478 RST.n1 RST.t2 18.1962
R1479 RST.n13 RST.t9 18.1962
R1480 RST.n39 RST.n37 9.33985
R1481 RST.n35 RST.n34 6.70742
R1482 RST.n29 RST.n28 5.42044
R1483 RST.n39 RST.n38 5.17836
R1484 RST RST.n0 4.57629
R1485 RST.n15 RST.n11 4.5005
R1486 RST.n15 RST.n14 4.5005
R1487 RST.n17 RST.n16 4.5005
R1488 RST.n33 RST.n32 3.49993
R1489 RST.n40 RST 2.27453
R1490 RST.n6 RST.n4 2.2505
R1491 RST.n18 RST.n17 2.2505
R1492 RST.n28 RST.n27 2.15059
R1493 RST.n32 RST.n31 2.14848
R1494 RST.n2 RST.n1 2.1224
R1495 RST.n14 RST.n13 2.12207
R1496 RST.n23 RST.n22 2.1217
R1497 RST.n34 RST.n21 2.06221
R1498 RST.n34 RST.n33 1.79221
R1499 RST.n21 RST.n8 1.78161
R1500 RST.n33 RST.n30 1.72354
R1501 RST.n21 RST.n20 1.53272
R1502 RST.n41 RST.n40 1.50509
R1503 RST.n30 RST.n26 1.1266
R1504 RST.n8 RST.n7 0.940487
R1505 RST.n43 RST.n0 0.90348
R1506 RST.n25 RST.n24 0.898026
R1507 RST.n43 RST.n42 0.722474
R1508 RST RST.n39 0.109973
R1509 RST.n32 RST 0.0563307
R1510 RST.n28 RST 0.0558741
R1511 RST.n24 RST 0.0553557
R1512 RST.n3 RST 0.0377414
R1513 RST.n4 RST.n3 0.0361897
R1514 RST.n11 RST 0.0348285
R1515 RST.n24 RST.n23 0.0275188
R1516 RST.n41 RST.n35 0.0274231
R1517 RST.n6 RST.n5 0.0267025
R1518 RST.n15 RST.n12 0.0255
R1519 RST.n10 RST.n9 0.0235
R1520 RST.n30 RST.n29 0.0175868
R1521 RST.n42 RST.n41 0.0140977
R1522 RST RST.n43 0.00984233
R1523 RST.n4 RST.n2 0.00515517
R1524 RST.n26 RST.n25 0.00494444
R1525 RST.n7 RST.n6 0.00372575
R1526 RST.n40 RST.n36 0.00217441
R1527 RST.n17 RST.n10 0.0015
R1528 RST.n17 RST.n15 0.0015
R1529 RST.n20 RST.n19 0.0015
R1530 RST.n19 RST.n18 0.0015
R1531 Q2.n18 Q2.t8 36.935
R1532 Q2.n12 Q2.t11 36.935
R1533 Q2.n28 Q2.t15 36.935
R1534 Q2.n4 Q2.t3 31.528
R1535 Q2.n0 Q2.t12 31.528
R1536 Q2.n30 Q2.t14 31.528
R1537 Q2.n23 Q2.t6 25.5364
R1538 Q2.n18 Q2.t5 18.1962
R1539 Q2.n12 Q2.t10 18.1962
R1540 Q2.n28 Q2.t7 18.1962
R1541 Q2.n4 Q2.t16 15.3826
R1542 Q2.n0 Q2.t9 15.3826
R1543 Q2.n30 Q2.t4 15.3826
R1544 Q2.n34 Q2.n9 14.2212
R1545 Q2.n23 Q2.t13 14.0749
R1546 Q2.n1 Q2.n0 7.63656
R1547 Q2.n38 Q2.n35 7.09905
R1548 Q2.n31 Q2.n30 6.86134
R1549 Q2.n5 Q2.n4 5.75592
R1550 Q2.n32 Q2.n29 5.01116
R1551 Q2.n9 Q2.n1 4.925
R1552 Q2.n14 Q2.n11 4.5005
R1553 Q2.n14 Q2.n13 4.5005
R1554 Q2.n17 Q2.n16 4.5005
R1555 Q2.n19 Q2.n16 4.5005
R1556 Q2.n27 Q2.n24 4.5005
R1557 Q2.n27 Q2.n26 4.5005
R1558 Q2.n5 Q2.n2 4.5005
R1559 Q2.n38 Q2.n37 3.25085
R1560 Q2.n8 Q2.n7 2.52083
R1561 Q2.n37 Q2.t1 2.2755
R1562 Q2.n37 Q2.n36 2.2755
R1563 Q2.n8 Q2 2.26388
R1564 Q2.n21 Q2.n20 2.25107
R1565 Q2.n39 Q2.n34 2.2505
R1566 Q2.n3 Q2.n2 2.2473
R1567 Q2.n7 Q2.n6 2.24676
R1568 Q2.n25 Q2.n22 2.2425
R1569 Q2.n29 Q2.n28 2.13398
R1570 Q2.n13 Q2.n12 2.12175
R1571 Q2.n19 Q2.n18 2.12075
R1572 Q2.n16 Q2.n15 1.74297
R1573 Q2.n15 Q2.n10 1.49778
R1574 Q2.n24 Q2.n23 1.42706
R1575 Q2.n33 Q2.n32 1.37495
R1576 Q2.n32 Q2.n31 1.12056
R1577 Q2.n22 Q2.n21 0.966797
R1578 Q2.n33 Q2.n27 0.836389
R1579 Q2.n26 Q2 0.1605
R1580 Q2.n34 Q2.n33 0.110256
R1581 Q2 Q2.n38 0.0862812
R1582 Q2.n31 Q2 0.0857632
R1583 Q2.n29 Q2 0.0810725
R1584 Q2.n1 Q2 0.0809204
R1585 Q2 Q2.n39 0.073625
R1586 Q2.n3 Q2 0.0565129
R1587 Q2.n17 Q2 0.0473512
R1588 Q2.n11 Q2 0.0473512
R1589 Q2.n20 Q2.n17 0.0361897
R1590 Q2.n11 Q2.n10 0.0361897
R1591 Q2.n26 Q2.n25 0.03175
R1592 Q2.n27 Q2.n22 0.0242114
R1593 Q2 Q2.n8 0.0199595
R1594 Q2.n6 Q2.n5 0.0191207
R1595 Q2.n6 Q2.n3 0.0172663
R1596 Q2.n9 Q2 0.0153101
R1597 Q2.n15 Q2.n14 0.0131772
R1598 Q2.n21 Q2.n16 0.0122182
R1599 Q2.n7 Q2.n2 0.0101966
R1600 Q2.n39 Q2 0.006125
R1601 Q2.n20 Q2.n19 0.00515517
R1602 Q2.n13 Q2.n10 0.00515517
R1603 Q2.n25 Q2.n24 0.00175
R1604 Q3.n0 Q3.t16 36.935
R1605 Q3.n30 Q3.t7 36.935
R1606 Q3.n24 Q3.t13 36.935
R1607 Q3.n2 Q3.t12 31.528
R1608 Q3.n7 Q3.t11 31.528
R1609 Q3.n12 Q3.t10 31.528
R1610 Q3.n17 Q3.t6 25.5364
R1611 Q3.n0 Q3.t15 18.1962
R1612 Q3.n30 Q3.t4 18.1962
R1613 Q3.n24 Q3.t9 18.1962
R1614 Q3.n2 Q3.t5 15.3826
R1615 Q3.n7 Q3.t3 15.3826
R1616 Q3.n12 Q3.t8 15.3826
R1617 Q3.n17 Q3.t14 14.0749
R1618 Q3.n13 Q3.n12 7.63631
R1619 Q3.n40 Q3.n37 7.09905
R1620 Q3.n3 Q3.n2 6.86134
R1621 Q3.n15 Q3.n11 6.23913
R1622 Q3.n8 Q3.n7 5.75592
R1623 Q3.n4 Q3.n1 5.01116
R1624 Q3.n14 Q3.n13 4.92545
R1625 Q3.n8 Q3.n5 4.5005
R1626 Q3.n26 Q3.n23 4.5005
R1627 Q3.n26 Q3.n25 4.5005
R1628 Q3.n29 Q3.n28 4.5005
R1629 Q3.n31 Q3.n28 4.5005
R1630 Q3.n18 Q3.n16 4.5005
R1631 Q3.n19 Q3.n16 4.5005
R1632 Q3.n40 Q3.n39 3.25085
R1633 Q3.n15 Q3 2.91397
R1634 Q3.n11 Q3.n10 2.52047
R1635 Q3.n41 Q3.n36 2.36285
R1636 Q3.n39 Q3.t0 2.2755
R1637 Q3.n39 Q3.n38 2.2755
R1638 Q3 Q3.n14 2.26759
R1639 Q3.n33 Q3.n32 2.25107
R1640 Q3.n6 Q3.n5 2.24713
R1641 Q3.n10 Q3.n9 2.24658
R1642 Q3.n21 Q3.n20 2.24235
R1643 Q3.n1 Q3.n0 2.13398
R1644 Q3.n25 Q3.n24 2.12175
R1645 Q3.n31 Q3.n30 2.12075
R1646 Q3.n35 Q3.n15 1.97218
R1647 Q3.n28 Q3.n27 1.74297
R1648 Q3.n27 Q3.n22 1.49778
R1649 Q3.n18 Q3.n17 1.42706
R1650 Q3.n36 Q3.n4 1.32654
R1651 Q3.n4 Q3.n3 1.12056
R1652 Q3.n34 Q3.n33 0.928385
R1653 Q3.n36 Q3.n35 0.57425
R1654 Q3.n35 Q3.n34 0.474184
R1655 Q3.n19 Q3 0.1605
R1656 Q3 Q3.n40 0.0862812
R1657 Q3.n3 Q3 0.0857632
R1658 Q3.n13 Q3 0.0811682
R1659 Q3.n1 Q3 0.0810725
R1660 Q3 Q3.n41 0.073625
R1661 Q3.n6 Q3 0.0565142
R1662 Q3.n29 Q3 0.0473512
R1663 Q3.n23 Q3 0.0473512
R1664 Q3.n34 Q3.n21 0.0435648
R1665 Q3.n32 Q3.n29 0.0361897
R1666 Q3.n23 Q3.n22 0.0361897
R1667 Q3.n20 Q3.n19 0.03175
R1668 Q3.n21 Q3.n16 0.0246174
R1669 Q3.n11 Q3 0.0199595
R1670 Q3.n9 Q3.n8 0.0191207
R1671 Q3.n9 Q3.n6 0.0172651
R1672 Q3.n14 Q3 0.0153101
R1673 Q3.n27 Q3.n26 0.0131772
R1674 Q3.n33 Q3.n28 0.0122182
R1675 Q3.n10 Q3.n5 0.0105495
R1676 Q3.n41 Q3 0.006125
R1677 Q3.n32 Q3.n31 0.00515517
R1678 Q3.n25 Q3.n22 0.00515517
R1679 Q3.n20 Q3.n18 0.00175
R1680 Q4.n4 Q4.t4 40.2519
R1681 Q4.n10 Q4.t6 36.935
R1682 Q4.n6 Q4.t9 31.528
R1683 Q4.n12 Q4.t3 31.528
R1684 Q4.n10 Q4.t5 18.1962
R1685 Q4.n4 Q4.t7 15.3826
R1686 Q4.n6 Q4.t8 15.3826
R1687 Q4.n12 Q4.t10 15.3826
R1688 Q4.n7 Q4.n6 7.63442
R1689 Q4.n3 Q4.n0 7.09905
R1690 Q4.n13 Q4.n12 6.86134
R1691 Q4.n14 Q4.n11 5.01116
R1692 Q4.n9 Q4 4.89286
R1693 Q4.n9 Q4.n5 4.81742
R1694 Q4.n3 Q4.n2 3.25085
R1695 Q4.n2 Q4.t1 2.2755
R1696 Q4.n2 Q4.n1 2.2755
R1697 Q4.n8 Q4 2.26567
R1698 Q4 Q4.n15 2.25751
R1699 Q4.n5 Q4.n4 2.15197
R1700 Q4.n11 Q4.n10 2.13398
R1701 Q4.n15 Q4.n14 1.52188
R1702 Q4.n8 Q4.n7 1.48351
R1703 Q4.n15 Q4.n9 1.36175
R1704 Q4.n14 Q4.n13 1.12056
R1705 Q4 Q4.n3 0.0919062
R1706 Q4.n13 Q4 0.0857632
R1707 Q4.n7 Q4 0.0831009
R1708 Q4.n11 Q4 0.0810725
R1709 Q4.n5 Q4 0.0389209
R1710 Q4 Q4.n8 0.00322727
R1711 Q1.n24 Q1.t12 36.935
R1712 Q1.n18 Q1.t10 36.935
R1713 Q1.n0 Q1.t16 36.935
R1714 Q1.n1 Q1.t15 31.528
R1715 Q1.n4 Q1.t8 31.528
R1716 Q1.n8 Q1.t9 31.4332
R1717 Q1.n11 Q1.t5 25.5364
R1718 Q1.n24 Q1.t6 18.1962
R1719 Q1.n18 Q1.t4 18.1962
R1720 Q1.n0 Q1.t14 18.1962
R1721 Q1.n8 Q1.t3 15.3826
R1722 Q1.n1 Q1.t13 15.3826
R1723 Q1.n4 Q1.t7 15.3826
R1724 Q1.n11 Q1.t11 14.0749
R1725 Q1.n2 Q1.n1 7.63417
R1726 Q1.n5 Q1.n4 7.62076
R1727 Q1.n31 Q1.t2 7.09905
R1728 Q1.n9 Q1.n8 6.86029
R1729 Q1.n35 Q1.n7 6.65668
R1730 Q1.n7 Q1.n3 5.46205
R1731 Q1.n6 Q1.n5 5.05792
R1732 Q1.n7 Q1 4.73586
R1733 Q1.n20 Q1.n17 4.5005
R1734 Q1.n20 Q1.n19 4.5005
R1735 Q1.n23 Q1.n22 4.5005
R1736 Q1.n25 Q1.n22 4.5005
R1737 Q1.n12 Q1.n10 4.5005
R1738 Q1.n13 Q1.n10 4.5005
R1739 Q1.n35 Q1.n34 3.41968
R1740 Q1.n31 Q1.n30 3.25053
R1741 Q1.n30 Q1.t0 2.2755
R1742 Q1.n30 Q1.n29 2.2755
R1743 Q1 Q1.n6 2.25519
R1744 Q1.n33 Q1.n32 2.25167
R1745 Q1.n27 Q1.n26 2.25107
R1746 Q1.n15 Q1.n14 2.24235
R1747 Q1.n36 Q1.n0 2.13459
R1748 Q1.n19 Q1.n18 2.12175
R1749 Q1.n25 Q1.n24 2.12075
R1750 Q1.n33 Q1.n28 2.05551
R1751 Q1.n22 Q1.n21 1.74297
R1752 Q1.n36 Q1.n35 1.5916
R1753 Q1.n34 Q1 1.52423
R1754 Q1.n21 Q1.n16 1.49778
R1755 Q1.n3 Q1.n2 1.48396
R1756 Q1.n12 Q1.n11 1.42706
R1757 Q1.n34 Q1.n9 1.12067
R1758 Q1.n28 Q1.n27 0.928385
R1759 Q1.n13 Q1 0.1605
R1760 Q1.n32 Q1.n31 0.0905
R1761 Q1.n9 Q1 0.0857632
R1762 Q1.n2 Q1 0.0833467
R1763 Q1 Q1.n36 0.0800273
R1764 Q1.n32 Q1 0.073625
R1765 Q1.n23 Q1 0.0473512
R1766 Q1.n17 Q1 0.0473512
R1767 Q1.n28 Q1.n15 0.0435648
R1768 Q1.n26 Q1.n23 0.0361897
R1769 Q1.n17 Q1.n16 0.0361897
R1770 Q1.n14 Q1.n13 0.03175
R1771 Q1.n5 Q1 0.0305
R1772 Q1.n15 Q1.n10 0.0246174
R1773 Q1.n21 Q1.n20 0.0131772
R1774 Q1.n27 Q1.n22 0.0122182
R1775 Q1.n6 Q1 0.0095
R1776 Q1.n26 Q1.n25 0.00515517
R1777 Q1.n19 Q1.n16 0.00515517
R1778 Q1.n3 Q1 0.00322727
R1779 Q1 Q1.n33 0.00283766
R1780 Q1.n14 Q1.n12 0.00175
R1781 JK_FF_mag_0.QB.n2 JK_FF_mag_0.QB.t6 37.1981
R1782 JK_FF_mag_0.QB.n1 JK_FF_mag_0.QB.t5 31.528
R1783 JK_FF_mag_0.QB.n2 JK_FF_mag_0.QB.t4 17.6611
R1784 JK_FF_mag_0.QB.n1 JK_FF_mag_0.QB.t3 15.3826
R1785 JK_FF_mag_0.QB JK_FF_mag_0.QB.n1 7.62751
R1786 JK_FF_mag_0.QB.n3 JK_FF_mag_0.QB 6.09789
R1787 JK_FF_mag_0.QB.n0 JK_FF_mag_0.QB.n5 2.99416
R1788 JK_FF_mag_0.QB.n3 JK_FF_mag_0.QB 2.67866
R1789 JK_FF_mag_0.QB.n5 JK_FF_mag_0.QB.t0 2.2755
R1790 JK_FF_mag_0.QB.n5 JK_FF_mag_0.QB.n4 2.2755
R1791 JK_FF_mag_0.QB.n0 JK_FF_mag_0.QB.n3 2.2505
R1792 JK_FF_mag_0.QB JK_FF_mag_0.QB.n2 1.43706
R1793 JK_FF_mag_0.QB JK_FF_mag_0.QB.n0 0.281955
R1794 CLK.n4 CLK.t0 36.935
R1795 CLK.n8 CLK.t5 36.935
R1796 CLK.n28 CLK.t4 31.528
R1797 CLK.n16 CLK.t6 25.4744
R1798 CLK.n4 CLK.t7 18.1962
R1799 CLK.n8 CLK.t2 18.1962
R1800 CLK.n28 CLK.t3 15.3826
R1801 CLK.n16 CLK.t1 14.1417
R1802 CLK.n29 CLK.n28 7.62171
R1803 CLK.n31 CLK.n30 5.58475
R1804 CLK.n30 CLK.n29 5.0581
R1805 CLK CLK.n32 4.55616
R1806 CLK.n24 CLK.n3 2.26042
R1807 CLK.n15 CLK.n7 2.25107
R1808 CLK.n3 CLK.n2 2.2505
R1809 CLK.n19 CLK.n18 2.24319
R1810 CLK.n23 CLK.n22 2.24244
R1811 CLK.n11 CLK.n8 2.12464
R1812 CLK.n5 CLK.n4 2.12188
R1813 CLK.n14 CLK.n13 1.71671
R1814 CLK.n27 CLK.n26 1.56853
R1815 CLK.n12 CLK.n11 1.50503
R1816 CLK.n17 CLK.n16 1.42118
R1817 CLK.n19 CLK.n15 0.964895
R1818 CLK.n31 CLK.n27 0.903813
R1819 CLK.n2 CLK.n1 0.09875
R1820 CLK.n2 CLK 0.04775
R1821 CLK.n6 CLK 0.0457995
R1822 CLK.n9 CLK 0.0457995
R1823 CLK.n22 CLK.n21 0.0403734
R1824 CLK.n13 CLK.n12 0.0386356
R1825 CLK.n7 CLK.n6 0.0377414
R1826 CLK.n10 CLK.n9 0.0377414
R1827 CLK.n21 CLK.n20 0.03466
R1828 CLK.n26 CLK.n25 0.0328596
R1829 CLK.n29 CLK 0.0316785
R1830 CLK.n20 CLK.n19 0.0207183
R1831 CLK.n24 CLK.n23 0.0181256
R1832 CLK.n15 CLK.n14 0.0122182
R1833 CLK.n30 CLK 0.0095
R1834 CLK CLK.n27 0.00561799
R1835 CLK.n32 CLK.n31 0.00464474
R1836 CLK.n7 CLK.n5 0.00360345
R1837 CLK.n25 CLK.n0 0.00286842
R1838 CLK.n11 CLK.n10 0.00203726
R1839 CLK.n18 CLK.n17 0.00175
R1840 CLK.n25 CLK.n24 0.00151124
R1841 Vdiv31.n2 Vdiv31.n1 9.33985
R1842 Vdiv31.n2 Vdiv31.n0 5.17836
R1843 Vdiv31 Vdiv31.n2 0.0749828
C0 Q4 a_8488_1345# 0.0694f
C1 a_7048_3814# Q0 0.00389f
C2 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.0877f
C3 a_211_2974# JK_FF_mag_2.nand2_mag_4.IN2 4.52e-20
C4 a_1810_1337# JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C5 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C6 JK_FF_mag_4.nand3_mag_0.OUT a_6796_1301# 0.0732f
C7 JK_FF_mag_1.nand2_mag_1.IN2 a_4852_1346# 0.069f
C8 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.00122f
C9 CLK and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0477f
C10 JK_FF_mag_3.nand3_mag_2.OUT CLK 0.242f
C11 a_5129_4070# Q0 0.0117f
C12 a_4442_205# RST 0.00187f
C13 JK_FF_mag_4.nand3_mag_0.OUT JK_FF_mag_4.nand3_mag_1.OUT 0.0622f
C14 JK_FF_mag_0.QB Q0 0.00258f
C15 Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VDD 0.519f
C16 a_8945_3798# and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.05e-20
C17 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C18 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_9909_3809# 8.67e-20
C19 JK_FF_mag_1.nand3_mag_1.OUT RST 0.289f
C20 Q2 JK_FF_mag_0.nand3_mag_1.IN1 0.00392f
C21 a_7354_204# VDD 2.21e-19
C22 JK_FF_mag_4.nand3_mag_0.OUT a_6636_1301# 0.0203f
C23 a_4442_205# Q3 0.0101f
C24 JK_FF_mag_2.QB JK_FF_mag_0.nand2_mag_1.IN2 3.48e-19
C25 JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.402f
C26 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN CLK 0.046f
C27 JK_FF_mag_3.nand2_mag_4.IN2 Q0 0.0635f
C28 a_1964_240# JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C29 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_0.QB 3.01e-20
C30 JK_FF_mag_1.nand3_mag_1.OUT Q3 0.0345f
C31 a_4969_4070# Q0 0.016f
C32 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_1.OUT 3.09e-19
C33 a_1246_1337# Q1 6.43e-21
C34 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 Q1 0.101f
C35 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_2.OUT 0.121f
C36 and_5_mag_0.and2_mag_1.IN2 VDD 0.387f
C37 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_8945_3798# 0.069f
C38 JK_FF_mag_2.QB Q1 1.98f
C39 Q4 nand_5_mag_0.GF_INV_MAG_0.IN 0.00849f
C40 JK_FF_mag_1.nand3_mag_2.OUT a_3558_205# 0.0202f
C41 or_2_mag_0.GF_INV_MAG_1.IN Vdiv31 0.128f
C42 Q0 JK_FF_mag_2.nand3_mag_2.OUT 0.235f
C43 and_5_mag_0.VOUT VDD 0.68f
C44 VDD and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.428f
C45 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.4e-21
C46 a_4405_4070# Q0 0.0102f
C47 JK_FF_mag_1.nand3_mag_1.OUT Q2 0.00182f
C48 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.00517f
C49 JK_FF_mag_4.nand2_mag_1.IN2 RST 0.00889f
C50 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C51 Q4 a_6796_1301# 2.79e-20
C52 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN Q4 5.09e-24
C53 Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 0.112f
C54 and_5_mag_0.and2_mag_2.IN2 VDD 0.388f
C55 a_775_2974# JK_FF_mag_2.nand2_mag_3.IN1 0.011f
C56 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 2.06e-19
C57 JK_FF_mag_4.QB JK_FF_mag_4.nand2_mag_1.IN2 0.0592f
C58 JK_FF_mag_0.nand2_mag_3.IN1 RST 0.071f
C59 JK_FF_mag_2.nand2_mag_1.IN2 a_775_2974# 0.069f
C60 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 4.31e-19
C61 JK_FF_mag_1.QB a_5570_249# 0.0811f
C62 JK_FF_mag_4.nand2_mag_1.IN2 Q3 1.48e-20
C63 a_7048_3814# VDD 3.14e-19
C64 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.129f
C65 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN or_2_mag_0.IN1 2.97e-19
C66 JK_FF_mag_4.nand3_mag_1.OUT Q4 0.0355f
C67 JK_FF_mag_3.nand3_mag_0.OUT Q0 9.41e-19
C68 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_2.OUT 0.121f
C69 JK_FF_mag_2.nand3_mag_1.OUT a_621_4071# 0.00378f
C70 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C71 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 8.46e-19
C72 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 RST 0.00589f
C73 a_4245_4070# Q0 0.0101f
C74 a_1810_1337# JK_FF_mag_2.QB 5e-20
C75 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 3.09e-19
C76 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_1.IN1 0.0385f
C77 a_5129_4070# VDD 0.00108f
C78 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_9908_3052# 8.67e-20
C79 a_5570_249# RST 9.82e-19
C80 JK_FF_mag_2.nand3_mag_0.OUT a_2063_2974# 0.0203f
C81 JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand2_mag_4.IN2 0.321f
C82 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 Q3 0.00525f
C83 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN RST 0.00994f
C84 JK_FF_mag_0.QB VDD 0.915f
C85 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.64e-19
C86 and_5_mag_0.and2_mag_1.IN2 Q1 0.00846f
C87 a_11530_2405# or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C88 JK_FF_mag_4.nand2_mag_1.IN2 Q2 4.94e-20
C89 a_8642_248# VDD 3.14e-19
C90 JK_FF_mag_4.nand3_mag_0.OUT JK_FF_mag_4.nand3_mag_1.IN1 0.122f
C91 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN RST 0.00661f
C92 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.16f
C93 JK_FF_mag_4.QB Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.00185f
C94 a_5570_249# Q3 0.0157f
C95 Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN Vdiv31 2.76e-19
C96 a_3681_4070# Q0 0.00859f
C97 Q1 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.298f
C98 Q2 JK_FF_mag_0.nand2_mag_3.IN1 0.0262f
C99 JK_FF_mag_1.nand3_mag_1.IN1 RST 0.2f
C100 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand3_mag_1.OUT 0.00975f
C101 JK_FF_mag_1.nand3_mag_1.OUT a_4399_2973# 4.61e-20
C102 or_2_mag_0.IN1 Vdiv31 0.00337f
C103 JK_FF_mag_4.nand2_mag_3.IN1 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 1.02e-20
C104 JK_FF_mag_4.nand2_mag_4.IN2 VDD 0.391f
C105 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_3.IN1 3.61e-20
C106 JK_FF_mag_3.nand2_mag_4.IN2 VDD 0.391f
C107 Q0 JK_FF_mag_2.nand2_mag_3.IN1 0.41f
C108 Q3 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0264f
C109 a_3724_1302# JK_FF_mag_0.QB 1.07e-20
C110 JK_FF_mag_2.nand2_mag_1.IN2 Q0 1.48e-20
C111 JK_FF_mag_2.nand3_mag_0.OUT a_1903_2974# 0.0732f
C112 a_7047_3047# nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.91e-21
C113 and_5_mag_0.and2_mag_2.IN2 Q1 1.01e-20
C114 Q2 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.102f
C115 JK_FF_mag_1.nand3_mag_1.IN1 Q3 0.00381f
C116 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_3.QB 9.89e-20
C117 JK_FF_mag_4.nand3_mag_0.OUT Q0 2.86e-19
C118 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_1.OUT 3.61e-20
C119 a_676_196# Q1 0.00164f
C120 a_7048_3814# Q1 0.00353f
C121 JK_FF_mag_1.nand3_mag_2.OUT a_4282_205# 9.1e-19
C122 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VDD 0.769f
C123 a_3117_4070# Q0 0.0157f
C124 VDD JK_FF_mag_2.nand3_mag_2.OUT 0.749f
C125 Vdiv31 RST 0.00235f
C126 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C127 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.429f
C128 and_5_mag_0.and2_mag_3.IN2 VDD 0.385f
C129 or_2_mag_0.IN1 or_2_mag_0.GF_INV_MAG_1.IN 0.208f
C130 a_4405_4070# VDD 2.21e-19
C131 a_3564_1302# JK_FF_mag_0.QB 1.4e-20
C132 Q2 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.318f
C133 JK_FF_mag_2.nand3_mag_0.OUT a_1339_2974# 0.00378f
C134 JK_FF_mag_0.nand3_mag_2.OUT VDD 0.752f
C135 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C136 a_5129_4070# Q1 0.00613f
C137 JK_FF_mag_1.nand3_mag_1.IN1 Q2 0.00273f
C138 JK_FF_mag_0.QB Q1 0.308f
C139 a_3558_205# a_3718_205# 0.0504f
C140 CLK Q0 0.306f
C141 JK_FF_mag_2.nand3_mag_1.IN1 RST 0.154f
C142 JK_FF_mag_3.nand3_mag_0.OUT VDD 0.744f
C143 or_2_mag_0.GF_INV_MAG_1.IN RST 0.0165f
C144 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 6.28e-19
C145 JK_FF_mag_4.nand2_mag_1.IN2 a_8488_1345# 0.00372f
C146 a_8944_3063# VDD 3.14e-19
C147 or_2_mag_0.IN1 a_11530_2405# 0.0144f
C148 CLK nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 8.46e-19
C149 JK_FF_mag_4.nand3_mag_1.IN1 Q4 0.00602f
C150 a_2374_1337# JK_FF_mag_0.QB 0.0114f
C151 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand3_mag_2.OUT 0.00168f
C152 JK_FF_mag_3.nand2_mag_4.IN2 Q1 0.00288f
C153 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C154 a_682_1293# Q2 2.79e-20
C155 a_4969_4070# Q1 0.006f
C156 JK_FF_mag_3.nand3_mag_1.OUT RST 0.273f
C157 a_621_4071# VDD 3.14e-19
C158 a_6790_204# RST 0.00189f
C159 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 8.03e-20
C160 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.11f
C161 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C162 a_7354_204# a_7514_204# 0.0504f
C163 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.OUT 3.58e-19
C164 a_11530_2405# RST 0.00703f
C165 JK_FF_mag_4.nand2_mag_1.IN2 a_7924_1345# 0.069f
C166 Q1 JK_FF_mag_2.nand3_mag_2.OUT 0.349f
C167 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.QB 0.25f
C168 a_6790_204# Q3 0.00214f
C169 a_3681_4070# VDD 3.14e-19
C170 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 7.4e-22
C171 Q4 Q0 0.192f
C172 JK_FF_mag_4.nand3_mag_0.OUT JK_FF_mag_4.nand2_mag_3.IN1 0.0886f
C173 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.00102f
C174 CLK a_9908_3052# 2.43e-19
C175 a_1810_1337# JK_FF_mag_0.QB 2.96e-19
C176 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN Q1 0.046f
C177 and_5_mag_0.and2_mag_3.IN2 Q1 0.0014f
C178 a_4405_4070# Q1 9.09e-19
C179 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN 0.0079f
C180 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C181 Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 7e-19
C182 Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN or_2_mag_0.IN1 0.0181f
C183 VDD JK_FF_mag_2.nand2_mag_3.IN1 1.32f
C184 JK_FF_mag_1.nand2_mag_3.IN1 RST 0.127f
C185 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN a_8488_1345# 6.6e-20
C186 JK_FF_mag_2.nand2_mag_1.IN2 VDD 0.401f
C187 JK_FF_mag_0.nand3_mag_2.OUT Q1 0.235f
C188 Q4 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00556f
C189 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_3.nand2_mag_3.IN1 8.93e-21
C190 a_8488_1345# nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 3.59e-20
C191 JK_FF_mag_4.nand3_mag_0.OUT VDD 0.745f
C192 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 a_7924_1345# 3.59e-20
C193 JK_FF_mag_1.nand3_mag_2.OUT VDD 0.749f
C194 a_1964_240# JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C195 JK_FF_mag_3.nand3_mag_1.OUT Q2 0.00136f
C196 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C197 JK_FF_mag_1.nand2_mag_3.IN1 Q3 0.0245f
C198 a_3117_4070# VDD 3.15e-19
C199 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_3.QB 6.46e-19
C200 JK_FF_mag_3.nand3_mag_0.OUT Q1 2.33e-20
C201 a_2063_2974# Q0 0.0101f
C202 a_1246_1337# JK_FF_mag_0.QB 3.33e-19
C203 a_8944_3063# Q1 7.37e-19
C204 Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN Vdiv31 1.34e-20
C205 a_4245_4070# Q1 9.09e-19
C206 JK_FF_mag_1.QB RST 0.221f
C207 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN a_7924_1345# 2.72e-20
C208 a_9909_3809# VDD 5.2e-19
C209 or_2_mag_0.IN1 RST 0.0122f
C210 a_621_4071# Q1 0.00859f
C211 a_2528_240# VDD 3.14e-19
C212 JK_FF_mag_1.QB JK_FF_mag_4.QB 2.42e-21
C213 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.IN1 0.768f
C214 and_5_mag_0.and2_mag_1.IN2 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.129f
C215 JK_FF_mag_1.nand2_mag_3.IN1 Q2 0.656f
C216 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN RST 0.00657f
C217 JK_FF_mag_1.QB Q3 1.97f
C218 CLK VDD 2.15f
C219 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_3.IN1 0.00279f
C220 a_1903_2974# Q0 0.00939f
C221 JK_FF_mag_1.nand3_mag_1.OUT a_3558_205# 1.17e-20
C222 a_3681_4070# Q1 0.00108f
C223 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_1.IN2 0.00975f
C224 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand2_mag_1.IN2 0.00975f
C225 a_8945_3798# VDD 3.14e-19
C226 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_1.IN2 5.06e-21
C227 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.00122f
C228 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN Q3 0.0129f
C229 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VDD 0.519f
C230 Q1 JK_FF_mag_2.nand2_mag_3.IN1 0.0291f
C231 a_1339_2974# JK_FF_mag_2.nand3_mag_1.OUT 0.0202f
C232 a_7047_3047# nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C233 JK_FF_mag_4.QB RST 0.11f
C234 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00113f
C235 JK_FF_mag_4.nand2_mag_3.IN1 Q4 0.193f
C236 JK_FF_mag_2.nand2_mag_1.IN2 Q1 0.11f
C237 Q3 RST 0.325f
C238 Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VDD 0.511f
C239 JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand3_mag_2.OUT 0.00118f
C240 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C241 JK_FF_mag_2.QB JK_FF_mag_2.nand3_mag_2.OUT 0.103f
C242 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.34e-21
C243 JK_FF_mag_3.QB RST 0.187f
C244 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_1.IN1 8.93e-21
C245 JK_FF_mag_3.nand3_mag_1.OUT a_4399_2973# 0.0202f
C246 a_7047_3047# RST 3.99e-19
C247 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.127f
C248 JK_FF_mag_1.QB Q2 0.321f
C249 JK_FF_mag_4.QB a_8078_248# 0.00964f
C250 Q2 a_516_196# 0.00335f
C251 JK_FF_mag_4.nand3_mag_0.OUT Q1 8.48e-20
C252 and_5_mag_0.and2_mag_3.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0016f
C253 a_1339_2974# Q0 6.43e-21
C254 JK_FF_mag_1.nand2_mag_3.IN1 a_4963_2973# 3.42e-20
C255 a_7994_3809# Q3 0.00943f
C256 a_211_2974# VDD 3.56e-19
C257 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_3.IN1 0.16f
C258 a_7048_3814# and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C259 JK_FF_mag_4.QB Q3 0.308f
C260 a_2374_1337# JK_FF_mag_2.nand2_mag_3.IN1 2.21e-19
C261 a_3117_4070# Q1 0.00108f
C262 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 3.48e-19
C263 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_1.IN2 6.04e-20
C264 Q4 VDD 3.05f
C265 JK_FF_mag_0.nand3_mag_1.OUT VDD 0.998f
C266 JK_FF_mag_4.nand3_mag_2.OUT VDD 0.75f
C267 a_7047_3047# Q3 0.0108f
C268 Q2 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0728f
C269 JK_FF_mag_4.nand2_mag_3.IN1 a_7993_3052# 3.66e-20
C270 a_9909_3809# Q1 2.43e-19
C271 Q2 RST 0.719f
C272 JK_FF_mag_1.nand2_mag_4.IN2 a_5570_249# 0.00372f
C273 a_5123_2973# RST 8.67e-19
C274 JK_FF_mag_1.QB JK_FF_mag_3.nand3_mag_1.IN1 9.89e-20
C275 JK_FF_mag_3.nand3_mag_1.OUT a_3835_2973# 4.52e-20
C276 a_8944_3063# nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 8.97e-21
C277 Q2 a_7994_3809# 0.0114f
C278 CLK Q1 0.666f
C279 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_3.nand2_mag_3.IN1 8.64e-20
C280 nand_5_mag_0.GF_INV_MAG_0.IN Vdiv31 1e-20
C281 JK_FF_mag_4.QB Q2 2.42e-20
C282 a_7993_3052# VDD 3.14e-19
C283 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 0.111f
C284 JK_FF_mag_1.QB JK_FF_mag_3.nand2_mag_1.IN2 3.09e-19
C285 a_2063_2974# VDD 0.00523f
C286 Q2 Q3 2.38f
C287 JK_FF_mag_3.QB Q2 0.0134f
C288 JK_FF_mag_2.QB a_621_4071# 0.00964f
C289 Q2 a_7047_3047# 0.00692f
C290 Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 0.00527f
C291 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN or_2_mag_0.IN1 0.00382f
C292 a_1240_196# RST 8.64e-19
C293 JK_FF_mag_3.nand3_mag_1.IN1 RST 0.205f
C294 Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.112f
C295 a_4963_2973# RST 7.2e-19
C296 Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN or_2_mag_0.IN1 0.118f
C297 a_4282_205# a_4442_205# 0.0504f
C298 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C299 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.00687f
C300 a_1185_4071# JK_FF_mag_2.nand3_mag_1.IN1 8.64e-19
C301 nand_5_mag_0.GF_INV_MAG_0.IN or_2_mag_0.GF_INV_MAG_1.IN 2.08e-19
C302 JK_FF_mag_1.QB JK_FF_mag_3.nand2_mag_3.IN1 6.46e-19
C303 Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN or_2_mag_0.IN1 0.00162f
C304 JK_FF_mag_3.nand2_mag_1.IN2 RST 0.02f
C305 a_211_2974# Q1 0.069f
C306 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN RST 0.0103f
C307 a_682_1293# JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C308 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_1.IN1 0.0386f
C309 JK_FF_mag_1.nand3_mag_1.OUT a_4282_205# 0.0203f
C310 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_2.OUT 0.121f
C311 JK_FF_mag_2.QB JK_FF_mag_2.nand2_mag_3.IN1 0.28f
C312 JK_FF_mag_3.QB a_4963_2973# 0.00392f
C313 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.QB 0.0592f
C314 Q4 Q1 0.775f
C315 JK_FF_mag_0.nand3_mag_1.OUT Q1 9.27e-19
C316 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_3.nand2_mag_3.IN1 0.00103f
C317 a_2069_4071# RST 0.00113f
C318 JK_FF_mag_4.QB Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 1.59e-19
C319 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VDD 0.39f
C320 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_1.IN2 0.0592f
C321 a_4399_2973# RST 3.98e-19
C322 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand3_mag_1.IN1 0.122f
C323 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand2_mag_1.IN2 0.109f
C324 JK_FF_mag_1.QB a_3835_2973# 4.61e-20
C325 Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN RST 0.00191f
C326 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C327 JK_FF_mag_3.nand2_mag_3.IN1 RST 0.0989f
C328 nand_5_mag_0.GF_INV_MAG_0.IN a_11530_2405# 4.15e-20
C329 Q2 a_1240_196# 0.0102f
C330 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_2.nand3_mag_1.IN1 6.28e-19
C331 a_1339_2974# VDD 3.14e-19
C332 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_3.IN2 4.92e-21
C333 Q2 JK_FF_mag_3.nand3_mag_1.IN1 0.00274f
C334 a_8488_1345# RST 6.56e-19
C335 a_4969_4070# a_5129_4070# 0.0504f
C336 JK_FF_mag_3.QB a_4399_2973# 3.29e-19
C337 a_4963_2973# a_5123_2973# 0.0504f
C338 Q3 JK_FF_mag_3.nand2_mag_3.IN1 4.92e-19
C339 a_2063_2974# Q1 4.47e-19
C340 Q4 a_6630_204# 0.00335f
C341 JK_FF_mag_4.nand2_mag_4.IN2 a_8642_248# 0.00372f
C342 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_3.IN1 0.28f
C343 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN RST 5.63e-20
C344 JK_FF_mag_4.nand3_mag_2.OUT a_6630_204# 0.0202f
C345 RST JK_FF_mag_2.nand2_mag_4.IN2 3.44e-19
C346 JK_FF_mag_4.QB a_8488_1345# 0.0114f
C347 a_1909_4071# RST 0.00113f
C348 Q2 JK_FF_mag_3.nand2_mag_1.IN2 0.00641f
C349 JK_FF_mag_0.nand3_mag_2.OUT a_676_196# 0.0731f
C350 JK_FF_mag_4.nand3_mag_1.IN1 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 4.73e-19
C351 a_3835_2973# RST 0.00173f
C352 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_3.IN1 5.53e-19
C353 CLK nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0014f
C354 JK_FF_mag_4.nand3_mag_1.OUT a_6790_204# 1.5e-20
C355 JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.655f
C356 Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VDD 0.519f
C357 JK_FF_mag_0.nand2_mag_4.IN2 RST 0.02f
C358 JK_FF_mag_0.nand2_mag_3.IN1 Q0 0.00133f
C359 a_1810_1337# JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C360 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN a_8642_248# 5.06e-20
C361 a_7924_1345# RST 6.56e-19
C362 JK_FF_mag_1.nand3_mag_1.OUT a_4852_1346# 4.52e-20
C363 JK_FF_mag_3.QB a_3835_2973# 2.96e-19
C364 a_1903_2974# Q1 3.43e-19
C365 Q2 JK_FF_mag_3.nand2_mag_3.IN1 0.243f
C366 a_1345_4071# RST 0.00171f
C367 JK_FF_mag_4.QB a_7924_1345# 2.96e-19
C368 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand3_mag_1.IN1 0.109f
C369 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.QB 0.103f
C370 a_3271_2973# RST 0.00252f
C371 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 Q0 4.09e-19
C372 a_1964_240# RST 9.46e-19
C373 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN JK_FF_mag_4.nand2_mag_4.IN2 3e-20
C374 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 0.321f
C375 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 Q1 0.0512f
C376 a_1400_196# JK_FF_mag_0.QB 0.00696f
C377 a_211_2974# JK_FF_mag_2.QB 0.0114f
C378 a_1246_1337# JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C379 Q2 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00164f
C380 Q4 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.00179f
C381 a_7360_1345# RST 5.43e-19
C382 JK_FF_mag_3.nand3_mag_2.OUT RST 0.0508f
C383 a_4399_2973# JK_FF_mag_3.nand3_mag_1.IN1 0.0697f
C384 JK_FF_mag_1.QB a_6796_1301# 1.33e-20
C385 JK_FF_mag_1.nand3_mag_1.OUT a_4288_1346# 0.0202f
C386 JK_FF_mag_3.QB a_3271_2973# 0.0114f
C387 a_7994_3809# and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C388 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand2_mag_3.IN1 0.233f
C389 JK_FF_mag_1.nand3_mag_1.OUT VDD 0.998f
C390 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 7.87e-19
C391 nand_5_mag_0.GF_INV_MAG_0.IN RST 0.147f
C392 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C393 a_4963_2973# JK_FF_mag_3.nand2_mag_3.IN1 0.00119f
C394 JK_FF_mag_1.nand3_mag_1.OUT a_5006_249# 0.00378f
C395 a_1185_4071# RST 0.00133f
C396 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN Q0 5.52e-20
C397 JK_FF_mag_1.nand2_mag_1.IN2 CLK 1.44e-19
C398 JK_FF_mag_4.QB a_7360_1345# 3.33e-19
C399 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 7.44e-19
C400 a_775_2974# JK_FF_mag_2.nand3_mag_1.IN1 0.0059f
C401 Q2 JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C402 a_7360_1345# Q3 6.43e-21
C403 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1.75e-19
C404 Q3 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.318f
C405 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_2.OUT 0.103f
C406 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand2_mag_3.IN1 0.36f
C407 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_4.IN2 0.199f
C408 Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN or_2_mag_0.IN1 0.0042f
C409 Q3 nand_5_mag_0.GF_INV_MAG_0.IN 3.08e-19
C410 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.00668f
C411 CLK and_5_mag_0.and2_mag_1.IN2 0.0502f
C412 JK_FF_mag_0.nand3_mag_1.IN1 Q1 3.67e-19
C413 a_6796_1301# RST 0.00154f
C414 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN RST 3.56e-20
C415 a_3835_2973# JK_FF_mag_3.nand3_mag_1.IN1 0.0059f
C416 Q2 a_3271_2973# 4.52e-19
C417 JK_FF_mag_1.QB a_6636_1301# 1.72e-20
C418 JK_FF_mag_2.nand3_mag_0.OUT RST 0.00961f
C419 Q2 a_1964_240# 0.00859f
C420 JK_FF_mag_4.nand3_mag_1.OUT nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 8.36e-19
C421 JK_FF_mag_4.nand2_mag_3.IN1 JK_FF_mag_4.nand2_mag_1.IN2 0.36f
C422 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN a_7994_3809# 4.56e-21
C423 and_5_mag_0.VOUT CLK 0.0094f
C424 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C425 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 8.18e-19
C426 CLK and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0454f
C427 a_4399_2973# JK_FF_mag_3.nand2_mag_3.IN1 1.43e-19
C428 JK_FF_mag_4.QB a_6796_1301# 0.00392f
C429 JK_FF_mag_4.nand3_mag_1.OUT RST 0.259f
C430 Q4 a_7514_204# 0.0101f
C431 JK_FF_mag_3.nand2_mag_1.IN2 a_3835_2973# 0.069f
C432 JK_FF_mag_0.QB JK_FF_mag_2.nand2_mag_3.IN1 0.00541f
C433 JK_FF_mag_1.nand2_mag_4.IN2 RST 0.0196f
C434 a_6796_1301# Q3 0.00939f
C435 JK_FF_mag_4.nand3_mag_2.OUT a_7514_204# 2.88e-20
C436 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN Q3 8.75e-19
C437 Q2 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.0264f
C438 Q4 a_7354_204# 0.0102f
C439 Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN RST 0.00191f
C440 JK_FF_mag_4.nand3_mag_2.OUT a_7354_204# 9.1e-19
C441 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_0.QB 3.48e-19
C442 a_57_4071# JK_FF_mag_2.nand2_mag_4.IN2 0.00372f
C443 JK_FF_mag_0.nand3_mag_2.OUT a_1400_196# 2.88e-20
C444 JK_FF_mag_4.nand3_mag_1.OUT a_8078_248# 0.00378f
C445 JK_FF_mag_3.QB JK_FF_mag_2.nand3_mag_0.OUT 2.79e-20
C446 and_5_mag_0.VOUT Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 1.56e-19
C447 a_8944_3063# nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.069f
C448 JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_1.OUT 0.25f
C449 JK_FF_mag_4.nand2_mag_1.IN2 VDD 0.4f
C450 and_5_mag_0.and2_mag_2.IN2 CLK 0.0512f
C451 a_3681_4070# JK_FF_mag_3.nand2_mag_4.IN2 0.069f
C452 a_1909_4071# a_2069_4071# 0.0504f
C453 a_6636_1301# RST 0.00185f
C454 a_4245_4070# a_4405_4070# 0.0504f
C455 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 0.768f
C456 JK_FF_mag_4.nand3_mag_1.OUT Q3 8.12e-19
C457 a_1903_2974# JK_FF_mag_2.QB 0.00392f
C458 JK_FF_mag_1.nand2_mag_4.IN2 Q3 0.0635f
C459 JK_FF_mag_4.nand2_mag_3.IN1 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 1.29e-20
C460 and_5_mag_0.VOUT Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN 0.00527f
C461 a_7048_3814# CLK 2.25e-19
C462 JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.28f
C463 a_3835_2973# JK_FF_mag_3.nand2_mag_3.IN1 0.011f
C464 Q0 JK_FF_mag_2.nand3_mag_1.IN1 9.71e-20
C465 JK_FF_mag_3.nand2_mag_1.IN2 a_3271_2973# 0.00372f
C466 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 4.92e-21
C467 and_5_mag_0.and2_mag_2.IN2 a_8945_3798# 0.00347f
C468 a_6636_1301# Q3 0.0101f
C469 a_1810_1337# JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C470 JK_FF_mag_3.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_2.OUT 0.00166f
C471 Q2 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.314f
C472 JK_FF_mag_4.nand2_mag_3.IN1 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 5.47e-20
C473 and_5_mag_0.VOUT Q4 2.07e-20
C474 JK_FF_mag_1.nand3_mag_1.IN1 a_4852_1346# 0.0059f
C475 Q4 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 9.67e-20
C476 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VDD 0.39f
C477 a_3558_205# RST 0.00189f
C478 a_5129_4070# CLK 0.00201f
C479 a_3117_4070# JK_FF_mag_3.nand2_mag_4.IN2 0.00372f
C480 JK_FF_mag_2.nand3_mag_2.OUT JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C481 a_2528_240# JK_FF_mag_0.QB 0.0811f
C482 JK_FF_mag_4.nand2_mag_3.IN1 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.62e-19
C483 JK_FF_mag_4.nand3_mag_1.OUT Q2 5.76e-22
C484 a_1339_2974# JK_FF_mag_2.QB 3.33e-19
C485 JK_FF_mag_3.nand3_mag_1.OUT Q0 0.0343f
C486 Q2 JK_FF_mag_1.nand2_mag_4.IN2 2.4e-19
C487 Q2 JK_FF_mag_0.nand3_mag_0.OUT 8.97e-19
C488 a_5570_249# VDD 3.15e-19
C489 a_3271_2973# JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C490 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VDD 0.515f
C491 a_3558_205# Q3 0.00335f
C492 a_1246_1337# JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C493 a_676_196# JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C494 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.432f
C495 JK_FF_mag_1.nand3_mag_1.IN1 a_4288_1346# 0.0697f
C496 JK_FF_mag_2.QB JK_FF_mag_0.nand3_mag_1.IN1 1.14e-19
C497 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_3.nand3_mag_1.OUT 1.77e-19
C498 JK_FF_mag_3.nand3_mag_2.OUT JK_FF_mag_3.nand2_mag_3.IN1 0.00118f
C499 JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.655f
C500 a_4969_4070# CLK 0.00194f
C501 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C502 JK_FF_mag_4.nand2_mag_1.IN2 Q1 3.86e-20
C503 and_5_mag_0.and2_mag_3.IN2 a_9909_3809# 0.00347f
C504 Q2 a_3558_205# 0.00185f
C505 JK_FF_mag_0.nand2_mag_3.IN1 Q1 0.427f
C506 a_621_4071# JK_FF_mag_2.nand2_mag_3.IN1 0.0036f
C507 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C508 JK_FF_mag_0.nand2_mag_4.IN2 a_1964_240# 0.069f
C509 Q4 a_8642_248# 0.0157f
C510 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.00102f
C511 JK_FF_mag_4.nand3_mag_1.IN1 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 4.3e-20
C512 CLK nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.09e-19
C513 and_5_mag_0.and2_mag_3.IN2 CLK 0.101f
C514 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand2_mag_3.IN1 0.0886f
C515 a_4405_4070# CLK 1.97e-19
C516 Vdiv31 VDD 0.152f
C517 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_3.nand2_mag_3.IN1 1.73e-20
C518 Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 0.112f
C519 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 Q1 0.0502f
C520 JK_FF_mag_4.nand3_mag_1.IN1 RST 0.162f
C521 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 3.59e-20
C522 a_2374_1337# JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C523 JK_FF_mag_1.QB a_4282_205# 0.00695f
C524 Q4 JK_FF_mag_4.nand2_mag_4.IN2 0.0637f
C525 and_5_mag_0.and2_mag_3.IN2 a_8945_3798# 8.97e-21
C526 JK_FF_mag_1.nand2_mag_3.IN1 a_5416_1346# 0.00118f
C527 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN or_2_mag_0.IN1 0.0104f
C528 Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.112f
C529 JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_1.IN1 0.0388f
C530 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 2.8e-19
C531 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN Q1 2.02e-19
C532 JK_FF_mag_4.nand3_mag_1.IN1 Q3 3.22e-19
C533 JK_FF_mag_3.nand3_mag_0.OUT CLK 0.271f
C534 JK_FF_mag_2.nand3_mag_1.OUT RST 0.256f
C535 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_3.IN1 0.36f
C536 VDD JK_FF_mag_2.nand3_mag_1.IN1 0.655f
C537 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN Q0 0.0943f
C538 Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.112f
C539 and_5_mag_0.and2_mag_2.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.00165f
C540 JK_FF_mag_4.nand2_mag_3.IN1 a_6790_204# 1.46e-19
C541 a_4245_4070# CLK 1.65e-19
C542 a_1185_4071# a_1345_4071# 0.0504f
C543 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C544 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN Q1 0.0477f
C545 or_2_mag_0.GF_INV_MAG_1.IN VDD 0.414f
C546 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 0.0263f
C547 Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN or_2_mag_0.IN1 0.012f
C548 Q0 RST 0.263f
C549 a_4282_205# RST 0.00171f
C550 a_1810_1337# JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C551 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN RST 0.0107f
C552 JK_FF_mag_3.nand3_mag_1.OUT a_4288_1346# 4.61e-20
C553 Q4 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00174f
C554 a_7994_3809# Q0 6.36e-20
C555 and_5_mag_0.and2_mag_3.IN2 Q4 3.13e-22
C556 JK_FF_mag_1.nand2_mag_3.IN1 a_4852_1346# 0.011f
C557 JK_FF_mag_1.QB a_5416_1346# 0.0114f
C558 a_522_1293# a_682_1293# 0.0504f
C559 JK_FF_mag_3.nand3_mag_1.OUT VDD 0.998f
C560 JK_FF_mag_4.QB Q0 6.38e-19
C561 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN RST 0.0152f
C562 Q3 Q0 0.983f
C563 JK_FF_mag_4.nand3_mag_1.OUT a_7924_1345# 4.52e-20
C564 JK_FF_mag_4.nand3_mag_1.IN1 Q2 2.93e-20
C565 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C566 JK_FF_mag_3.QB Q0 1.96f
C567 a_4282_205# Q3 0.0102f
C568 a_7047_3047# Q0 0.00347f
C569 JK_FF_mag_1.nand3_mag_0.OUT RST 0.0231f
C570 a_1400_196# JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C571 a_11530_2405# VDD 0.165f
C572 a_682_1293# Q1 0.00939f
C573 Q3 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00164f
C574 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 2.17e-19
C575 a_1246_1337# JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C576 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C577 a_7993_3052# nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 4.18e-21
C578 a_5416_1346# RST 0.00126f
C579 JK_FF_mag_1.nand2_mag_3.IN1 a_4288_1346# 1.43e-19
C580 JK_FF_mag_1.nand3_mag_0.OUT Q3 8.31e-19
C581 JK_FF_mag_1.QB a_4852_1346# 2.96e-19
C582 JK_FF_mag_2.QB JK_FF_mag_0.nand2_mag_3.IN1 0.00541f
C583 JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.24f
C584 a_9908_3052# RST 9.29e-19
C585 JK_FF_mag_1.nand2_mag_3.IN1 a_5006_249# 0.0036f
C586 JK_FF_mag_4.nand3_mag_1.OUT a_7360_1345# 0.0202f
C587 Q2 Q0 0.664f
C588 a_5123_2973# Q0 5.54e-19
C589 a_5416_1346# Q3 0.069f
C590 JK_FF_mag_1.QB JK_FF_mag_4.nand2_mag_3.IN1 6.23e-20
C591 Q1 JK_FF_mag_2.nand3_mag_1.IN1 0.00393f
C592 Q3 a_9908_3052# 4.35e-19
C593 or_2_mag_0.GF_INV_MAG_1.IN Q1 6.26e-20
C594 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_1.IN1 0.038f
C595 a_4852_1346# RST 0.00126f
C596 Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VDD 0.517f
C597 JK_FF_mag_1.nand3_mag_0.OUT Q2 0.273f
C598 a_211_2974# JK_FF_mag_2.nand2_mag_3.IN1 0.00118f
C599 a_9909_3809# CLK 0.00479f
C600 JK_FF_mag_1.QB a_4288_1346# 3.25e-19
C601 JK_FF_mag_4.nand2_mag_3.IN1 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.36e-20
C602 JK_FF_mag_1.nand2_mag_3.IN1 a_3724_1302# 0.00119f
C603 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 2.91e-19
C604 JK_FF_mag_2.nand2_mag_1.IN2 a_211_2974# 0.00372f
C605 JK_FF_mag_1.QB VDD 0.915f
C606 JK_FF_mag_1.QB a_5006_249# 0.00964f
C607 a_516_196# VDD 0.00108f
C608 or_2_mag_0.IN1 VDD 0.728f
C609 JK_FF_mag_3.nand3_mag_1.IN1 Q0 0.00335f
C610 JK_FF_mag_4.nand2_mag_3.IN1 RST 0.0618f
C611 JK_FF_mag_3.nand3_mag_1.OUT Q1 0.0048f
C612 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 1.97e-19
C613 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.119f
C614 a_4963_2973# Q0 4.21e-19
C615 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_3.IN1 5.53e-19
C616 a_4852_1346# Q3 6.03e-21
C617 Q2 a_5416_1346# 4.6e-19
C618 JK_FF_mag_3.QB a_4852_1346# 4.61e-20
C619 JK_FF_mag_4.nand2_mag_3.IN1 a_8078_248# 0.0036f
C620 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.431f
C621 JK_FF_mag_3.nand2_mag_1.IN2 Q0 0.107f
C622 a_6636_1301# a_6796_1301# 0.0504f
C623 JK_FF_mag_4.nand3_mag_0.OUT Q4 0.00517f
C624 JK_FF_mag_4.QB JK_FF_mag_4.nand2_mag_3.IN1 0.28f
C625 a_11530_2405# Q1 1.78e-19
C626 a_4288_1346# RST 6.86e-19
C627 JK_FF_mag_4.nand3_mag_0.OUT JK_FF_mag_4.nand3_mag_2.OUT 0.00183f
C628 JK_FF_mag_2.nand3_mag_1.OUT a_2069_4071# 1.17e-20
C629 JK_FF_mag_4.nand2_mag_3.IN1 Q3 0.434f
C630 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_3.nand3_mag_1.IN1 6.95e-19
C631 a_8945_3798# CLK 7.37e-19
C632 VDD RST 3.98f
C633 a_5006_249# RST 9.62e-19
C634 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.111f
C635 JK_FF_mag_1.QB a_3724_1302# 0.00392f
C636 a_7994_3809# VDD 3.14e-19
C637 a_2069_4071# Q0 0.00144f
C638 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 a_8944_3063# 0.00347f
C639 a_8078_248# VDD 3.14e-19
C640 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 1.15e-19
C641 a_6630_204# a_6790_204# 0.0504f
C642 JK_FF_mag_4.QB VDD 0.914f
C643 JK_FF_mag_3.nand2_mag_3.IN1 Q0 0.0218f
C644 Q3 VDD 3.01f
C645 a_5006_249# Q3 0.00859f
C646 JK_FF_mag_3.QB VDD 0.917f
C647 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 4.29e-20
C648 a_7047_3047# VDD 3.14e-19
C649 JK_FF_mag_2.nand3_mag_1.OUT a_1909_4071# 1.5e-20
C650 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 and_5_mag_0.and2_mag_1.IN2 0.0016f
C651 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.nand2_mag_4.IN2 0.122f
C652 JK_FF_mag_4.nand3_mag_1.IN1 a_7924_1345# 0.0059f
C653 Q4 CLK 0.00597f
C654 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.0016f
C655 JK_FF_mag_4.nand2_mag_3.IN1 Q2 0.00113f
C656 Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 7e-19
C657 a_3724_1302# RST 0.00229f
C658 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN or_2_mag_0.IN1 0.0829f
C659 a_1400_196# JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C660 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_3.nand2_mag_3.IN1 1.01e-19
C661 a_1909_4071# Q0 0.00169f
C662 Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN or_2_mag_0.IN1 0.108f
C663 a_1903_2974# JK_FF_mag_2.nand2_mag_3.IN1 0.00119f
C664 a_3835_2973# Q0 6.14e-21
C665 Q2 a_4288_1346# 6.43e-21
C666 or_2_mag_0.IN1 Q1 1.64e-19
C667 a_516_196# Q1 0.00117f
C668 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C669 a_3724_1302# Q3 2.79e-20
C670 a_676_196# JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C671 JK_FF_mag_1.nand3_mag_2.OUT a_3718_205# 0.0731f
C672 JK_FF_mag_2.QB JK_FF_mag_2.nand3_mag_1.IN1 0.0381f
C673 Q2 VDD 4.34f
C674 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.00113f
C675 JK_FF_mag_0.nand2_mag_1.IN2 RST 0.01f
C676 a_5123_2973# VDD 0.00503f
C677 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN RST 0.00111f
C678 JK_FF_mag_4.nand3_mag_1.IN1 a_7360_1345# 0.0697f
C679 JK_FF_mag_2.nand3_mag_1.OUT a_1345_4071# 0.0203f
C680 a_3564_1302# RST 0.003f
C681 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN Q1 0.0443f
C682 a_1339_2974# JK_FF_mag_2.nand2_mag_3.IN1 1.43e-19
C683 Q1 RST 0.137f
C684 a_3271_2973# Q0 0.069f
C685 a_1240_196# VDD 2.21e-19
C686 Q4 JK_FF_mag_4.nand3_mag_2.OUT 0.338f
C687 a_7994_3809# Q1 3.11e-21
C688 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_3.IN1 0.28f
C689 a_3724_1302# Q2 0.00939f
C690 JK_FF_mag_3.nand3_mag_1.IN1 VDD 0.655f
C691 JK_FF_mag_4.QB Q1 9.12e-20
C692 JK_FF_mag_2.nand3_mag_1.OUT a_1185_4071# 0.0733f
C693 Q3 Q1 0.813f
C694 JK_FF_mag_4.nand2_mag_1.IN2 JK_FF_mag_4.nand2_mag_4.IN2 8.16e-20
C695 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN Q0 6.3e-20
C696 JK_FF_mag_3.nand3_mag_2.OUT Q0 0.365f
C697 a_2374_1337# RST 0.00157f
C698 JK_FF_mag_3.QB Q1 0.00585f
C699 a_7047_3047# Q1 2.95e-21
C700 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.00103f
C701 JK_FF_mag_3.nand2_mag_1.IN2 VDD 0.402f
C702 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_0.OUT 1.77e-19
C703 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VDD 0.517f
C704 and_5_mag_0.VOUT Vdiv31 4.61e-19
C705 Q2 JK_FF_mag_0.nand2_mag_1.IN2 0.11f
C706 a_57_4071# VDD 3.14e-19
C707 Q4 a_7993_3052# 3.11e-21
C708 a_6630_204# RST 0.00189f
C709 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN nand_5_mag_0.GF_INV_MAG_0.IN 4.48e-19
C710 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand3_mag_1.IN1 0.768f
C711 Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VDD 0.519f
C712 JK_FF_mag_4.nand2_mag_3.IN1 a_8488_1345# 0.00118f
C713 a_3564_1302# Q2 0.0101f
C714 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN nand_5_mag_0.GF_INV_MAG_0.IN 0.128f
C715 a_2069_4071# VDD 0.00108f
C716 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand3_mag_1.OUT 0.0622f
C717 a_4399_2973# VDD 3.14e-19
C718 Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VDD 0.514f
C719 JK_FF_mag_3.nand2_mag_3.IN1 VDD 1.22f
C720 Q2 Q1 0.893f
C721 a_6630_204# Q3 0.00182f
C722 a_1810_1337# RST 0.001f
C723 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_0.OUT 4.31e-19
C724 JK_FF_mag_2.nand3_mag_0.OUT Q0 0.267f
C725 a_8488_1345# VDD 3.56e-19
C726 and_5_mag_0.VOUT or_2_mag_0.GF_INV_MAG_1.IN 1.65e-20
C727 JK_FF_mag_4.nand2_mag_3.IN1 a_7924_1345# 0.011f
C728 a_2374_1337# Q2 0.069f
C729 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C730 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD 0.426f
C731 VDD JK_FF_mag_2.nand2_mag_4.IN2 0.391f
C732 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN 0.00617f
C733 a_3835_2973# VDD 3.14e-19
C734 a_3724_1302# JK_FF_mag_3.nand2_mag_3.IN1 3.42e-20
C735 JK_FF_mag_3.nand3_mag_1.IN1 Q1 7.98e-19
C736 JK_FF_mag_1.nand3_mag_2.OUT a_4442_205# 2.88e-20
C737 Q4 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.00171f
C738 a_1246_1337# RST 4.22e-20
C739 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 4.17e-19
C740 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.11f
C741 a_682_1293# JK_FF_mag_0.QB 0.00392f
C742 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C743 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 RST 0.00941f
C744 JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C745 JK_FF_mag_2.QB RST 0.105f
C746 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C747 a_7924_1345# VDD 3.14e-19
C748 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 0.00529f
C749 JK_FF_mag_3.nand2_mag_1.IN2 Q1 3.27e-20
C750 a_1903_2974# a_2063_2974# 0.0504f
C751 a_1339_2974# JK_FF_mag_0.nand3_mag_1.OUT 5e-20
C752 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN Q1 6.2e-19
C753 JK_FF_mag_4.nand2_mag_3.IN1 a_7360_1345# 1.43e-19
C754 a_57_4071# Q1 0.0157f
C755 a_1810_1337# Q2 1.46e-21
C756 a_1345_4071# VDD 2.21e-19
C757 Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN or_2_mag_0.IN1 0.0123f
C758 Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.112f
C759 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 2.23e-19
C760 a_5416_1346# JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C761 a_3271_2973# VDD 3.56e-19
C762 Q3 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 0.0124f
C763 a_1964_240# VDD 3.14e-19
C764 JK_FF_mag_3.QB JK_FF_mag_2.QB 2.46e-21
C765 a_2069_4071# Q1 0.0122f
C766 JK_FF_mag_0.QB JK_FF_mag_2.nand3_mag_1.IN1 1.14e-19
C767 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C768 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN 1.33e-19
C769 JK_FF_mag_3.nand2_mag_3.IN1 Q1 0.00119f
C770 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C771 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VDD 0.43f
C772 a_7360_1345# VDD 3.14e-19
C773 JK_FF_mag_3.nand3_mag_2.OUT VDD 0.755f
C774 Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN RST 7.05e-19
C775 JK_FF_mag_4.nand2_mag_3.IN1 a_6796_1301# 0.00119f
C776 nand_5_mag_0.GF_INV_MAG_0.IN VDD 0.418f
C777 JK_FF_mag_3.nand3_mag_1.OUT a_5129_4070# 1.17e-20
C778 a_7514_204# RST 0.00147f
C779 a_775_2974# JK_FF_mag_2.nand3_mag_1.OUT 4.52e-20
C780 a_7354_204# RST 0.0017f
C781 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.0822f
C782 and_5_mag_0.VOUT Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.00174f
C783 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN a_8944_3063# 1.05e-20
C784 Q2 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 1.05e-20
C785 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_3.nand3_mag_0.OUT 6.95e-19
C786 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.00279f
C787 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN Q1 8.4e-19
C788 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C789 a_1909_4071# Q1 0.0151f
C790 Q1 JK_FF_mag_2.nand2_mag_4.IN2 0.0635f
C791 JK_FF_mag_4.QB a_7514_204# 0.00696f
C792 and_5_mag_0.VOUT or_2_mag_0.IN1 0.0102f
C793 JK_FF_mag_1.nand2_mag_1.IN2 RST 0.0132f
C794 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand2_mag_3.IN1 0.16f
C795 JK_FF_mag_4.QB a_7354_204# 0.00695f
C796 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VDD 0.429f
C797 JK_FF_mag_2.nand3_mag_0.OUT VDD 0.746f
C798 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand2_mag_4.IN2 0.122f
C799 and_5_mag_0.and2_mag_1.IN2 RST 2.65e-20
C800 JK_FF_mag_3.nand3_mag_1.OUT a_4969_4070# 1.5e-20
C801 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand3_mag_2.OUT 0.00161f
C802 JK_FF_mag_1.nand2_mag_1.IN2 Q3 0.109f
C803 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.00112f
C804 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_3.QB 3.09e-19
C805 JK_FF_mag_4.nand3_mag_1.OUT VDD 0.998f
C806 a_7994_3809# and_5_mag_0.and2_mag_1.IN2 0.00347f
C807 and_5_mag_0.VOUT RST 0.0197f
C808 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_0.QB 7.57e-20
C809 JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.391f
C810 JK_FF_mag_0.nand3_mag_0.OUT VDD 0.744f
C811 a_1345_4071# Q1 0.0102f
C812 Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VDD 0.517f
C813 a_516_196# a_676_196# 0.0504f
C814 JK_FF_mag_1.nand2_mag_4.IN2 a_5006_249# 0.069f
C815 and_5_mag_0.and2_mag_1.IN2 Q3 0.102f
C816 a_2374_1337# JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C817 a_7994_3809# and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 3.85e-20
C818 a_6636_1301# VDD 0.00554f
C819 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN Q1 1.88e-19
C820 Q3 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0725f
C821 and_5_mag_0.and2_mag_2.IN2 RST 4.4e-20
C822 JK_FF_mag_3.nand3_mag_2.OUT Q1 0.00542f
C823 JK_FF_mag_2.QB a_57_4071# 0.0811f
C824 JK_FF_mag_3.nand3_mag_1.OUT a_4405_4070# 0.0203f
C825 JK_FF_mag_2.nand3_mag_1.OUT Q0 6.64e-19
C826 JK_FF_mag_1.nand2_mag_1.IN2 Q2 0.0064f
C827 nand_5_mag_0.GF_INV_MAG_0.IN Q1 0.0103f
C828 JK_FF_mag_1.QB JK_FF_mag_0.QB 2e-21
C829 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00164f
C830 a_1185_4071# Q1 0.0101f
C831 and_5_mag_0.and2_mag_2.IN2 Q3 0.0124f
C832 Q2 and_5_mag_0.and2_mag_1.IN2 0.00542f
C833 a_3558_205# VDD 0.00108f
C834 a_682_1293# JK_FF_mag_2.nand2_mag_3.IN1 3.87e-20
C835 JK_FF_mag_3.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_0.OUT 0.0622f
C836 JK_FF_mag_4.nand2_mag_1.IN2 Q4 0.115f
C837 a_7048_3814# Q3 0.00665f
C838 Q2 and_5_mag_0.VOUT 3.05e-19
C839 a_522_1293# JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C840 a_211_2974# JK_FF_mag_0.nand2_mag_3.IN1 2.21e-19
C841 JK_FF_mag_1.nand3_mag_1.OUT a_3718_205# 1.5e-20
C842 Q2 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0126f
C843 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN Q1 8.11e-19
C844 JK_FF_mag_3.nand3_mag_1.OUT a_4245_4070# 0.0733f
C845 JK_FF_mag_0.QB RST 0.157f
C846 JK_FF_mag_2.nand3_mag_0.OUT Q1 0.00106f
C847 JK_FF_mag_2.QB JK_FF_mag_2.nand2_mag_4.IN2 0.198f
C848 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C849 JK_FF_mag_4.nand3_mag_1.OUT Q1 2.59e-20
C850 JK_FF_mag_0.nand3_mag_0.OUT Q1 0.269f
C851 and_5_mag_0.and2_mag_2.IN2 Q2 0.0782f
C852 JK_FF_mag_2.nand3_mag_1.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.233f
C853 Q3 JK_FF_mag_0.QB 2.1e-19
C854 Q4 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 0.0107f
C855 JK_FF_mag_4.QB a_8642_248# 0.0811f
C856 Q2 a_676_196# 0.00789f
C857 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_3.nand3_mag_0.OUT 1.01e-19
C858 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand3_mag_1.IN1 0.109f
C859 a_775_2974# VDD 3.14e-19
C860 Q2 a_7048_3814# 0.0108f
C861 JK_FF_mag_3.nand2_mag_4.IN2 RST 0.0214f
C862 JK_FF_mag_4.nand2_mag_4.IN2 RST 8.23e-19
C863 JK_FF_mag_3.nand3_mag_1.OUT a_3681_4070# 0.00378f
C864 JK_FF_mag_4.nand3_mag_1.IN1 JK_FF_mag_4.nand2_mag_3.IN1 0.233f
C865 JK_FF_mag_4.nand2_mag_4.IN2 a_8078_248# 0.069f
C866 JK_FF_mag_2.QB a_1345_4071# 0.00695f
C867 JK_FF_mag_4.QB JK_FF_mag_4.nand2_mag_4.IN2 0.199f
C868 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_3.nand2_mag_3.IN1 6.04e-20
C869 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 0.0147f
C870 JK_FF_mag_0.nand3_mag_2.OUT a_516_196# 0.0202f
C871 a_9908_3052# nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.069f
C872 JK_FF_mag_4.nand3_mag_1.OUT a_6630_204# 1.17e-20
C873 JK_FF_mag_3.QB JK_FF_mag_3.nand2_mag_4.IN2 0.199f
C874 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN RST 0.00619f
C875 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 1.9e-21
C876 Q4 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.00237f
C877 RST JK_FF_mag_2.nand3_mag_2.OUT 0.0857f
C878 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 a_7993_3052# 0.00347f
C879 Q2 JK_FF_mag_0.QB 2f
C880 JK_FF_mag_4.nand3_mag_1.IN1 VDD 0.655f
C881 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN RST 0.00751f
C882 and_5_mag_0.and2_mag_3.IN2 RST 1.08e-19
C883 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN a_8078_248# 1.76e-20
C884 a_4405_4070# RST 8.64e-19
C885 JK_FF_mag_4.QB Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN 8.53e-19
C886 JK_FF_mag_4.nand2_mag_3.IN1 Q0 0.00381f
C887 JK_FF_mag_0.nand3_mag_2.OUT RST 0.0494f
C888 a_1903_2974# JK_FF_mag_0.nand2_mag_3.IN1 3.87e-20
C889 JK_FF_mag_2.QB a_1185_4071# 0.00696f
C890 JK_FF_mag_2.nand3_mag_1.OUT VDD 0.998f
C891 Q3 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.314f
C892 a_1400_196# RST 0.00186f
C893 and_5_mag_0.and2_mag_3.IN2 Q3 1.05e-20
C894 Q2 JK_FF_mag_3.nand2_mag_4.IN2 2.33e-19
C895 a_7993_3052# nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.069f
C896 JK_FF_mag_3.QB a_4405_4070# 0.00695f
C897 a_1240_196# JK_FF_mag_0.QB 0.00695f
C898 JK_FF_mag_3.nand3_mag_0.OUT RST 0.012f
C899 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN and_5_mag_0.VOUT 0.119f
C900 VDD Q0 2.56f
C901 a_8944_3063# RST 2.96e-19
C902 a_4282_205# VDD 2.21e-19
C903 JK_FF_mag_3.nand3_mag_1.OUT CLK 0.00317f
C904 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C905 a_4245_4070# RST 0.00187f
C906 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VDD 0.512f
C907 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.QB 0.343f
C908 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN or_2_mag_0.GF_INV_MAG_1.IN 8.18e-19
C909 a_1246_1337# JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C910 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 5.06e-21
C911 JK_FF_mag_1.nand3_mag_1.OUT a_4442_205# 0.0733f
C912 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VDD 0.431f
C913 JK_FF_mag_1.nand3_mag_0.OUT a_4288_1346# 0.00378f
C914 JK_FF_mag_3.QB JK_FF_mag_3.nand3_mag_0.OUT 0.343f
C915 Q2 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 8.87e-19
C916 Q3 a_8944_3063# 0.0193f
C917 JK_FF_mag_1.nand3_mag_0.OUT VDD 0.745f
C918 Q2 and_5_mag_0.and2_mag_3.IN2 0.0127f
C919 Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VDD 0.516f
C920 JK_FF_mag_3.QB a_4245_4070# 0.00696f
C921 Q2 JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C922 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_2.nand3_mag_1.IN1 3.48e-19
C923 JK_FF_mag_1.QB JK_FF_mag_4.nand3_mag_0.OUT 2.74e-20
C924 Q4 or_2_mag_0.GF_INV_MAG_1.IN 0.0403f
C925 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C926 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_3.nand2_mag_4.IN2 8.16e-20
C927 a_3681_4070# RST 9.7e-19
C928 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C929 JK_FF_mag_1.nand2_mag_3.IN1 CLK 6.68e-19
C930 a_5416_1346# VDD 3.56e-19
C931 Q2 a_1400_196# 0.0101f
C932 JK_FF_mag_4.nand3_mag_1.IN1 Q1 4.21e-20
C933 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.128f
C934 and_5_mag_0.and2_mag_1.IN2 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.12f
C935 RST JK_FF_mag_2.nand2_mag_3.IN1 0.0119f
C936 a_9908_3052# VDD 5.19e-19
C937 Q2 JK_FF_mag_3.nand3_mag_0.OUT 0.00627f
C938 JK_FF_mag_3.nand3_mag_0.OUT a_5123_2973# 0.0203f
C939 JK_FF_mag_4.nand3_mag_0.OUT nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 6.2e-20
C940 JK_FF_mag_1.nand3_mag_0.OUT a_3724_1302# 0.0732f
C941 JK_FF_mag_0.nand2_mag_1.IN2 Q0 1.28e-19
C942 Q2 a_8944_3063# 9.22e-21
C943 Q4 a_6790_204# 0.00789f
C944 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 2.23e-19
C945 JK_FF_mag_4.nand3_mag_2.OUT a_6790_204# 0.0731f
C946 JK_FF_mag_3.QB a_3681_4070# 0.00964f
C947 JK_FF_mag_2.nand3_mag_1.OUT Q1 0.0346f
C948 JK_FF_mag_0.nand3_mag_2.OUT a_1240_196# 9.1e-19
C949 JK_FF_mag_4.nand3_mag_0.OUT RST 0.0173f
C950 JK_FF_mag_4.nand3_mag_1.OUT a_7514_204# 0.0733f
C951 Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 0.112f
C952 and_5_mag_0.VOUT nand_5_mag_0.GF_INV_MAG_0.IN 5.16e-20
C953 JK_FF_mag_3.nand2_mag_4.IN2 JK_FF_mag_3.nand2_mag_3.IN1 0.321f
C954 JK_FF_mag_4.nand3_mag_1.OUT a_7354_204# 0.0203f
C955 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 1.03e-19
C956 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN 0.108f
C957 JK_FF_mag_1.nand3_mag_2.OUT RST 0.0859f
C958 Q4 a_11530_2405# 8.64e-19
C959 a_1240_196# a_1400_196# 0.0504f
C960 a_3117_4070# RST 9.87e-19
C961 JK_FF_mag_3.QB JK_FF_mag_2.nand2_mag_3.IN1 3.21e-19
C962 a_4852_1346# VDD 3.14e-19
C963 JK_FF_mag_1.QB CLK 2.15e-19
C964 Q0 Q1 2.08f
C965 a_8488_1345# JK_FF_mag_4.nand2_mag_4.IN2 4.52e-20
C966 JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_0.OUT 0.343f
C967 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.128f
C968 a_2069_4071# JK_FF_mag_2.nand3_mag_2.OUT 0.0202f
C969 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_4.IN2 8.16e-20
C970 JK_FF_mag_4.nand3_mag_0.OUT Q3 0.269f
C971 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.nand3_mag_1.IN1 0.122f
C972 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.QB 0.199f
C973 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN 0.112f
C974 JK_FF_mag_1.nand3_mag_2.OUT Q3 0.338f
C975 a_9909_3809# RST 6.53e-20
C976 JK_FF_mag_3.nand3_mag_0.OUT a_4963_2973# 0.0732f
C977 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.107f
C978 JK_FF_mag_1.nand3_mag_0.OUT a_3564_1302# 0.0203f
C979 a_7048_3814# and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 4.6e-21
C980 JK_FF_mag_4.nand2_mag_3.IN1 VDD 1.25f
C981 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN and_5_mag_0.VOUT 5.82e-21
C982 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN Q1 0.3f
C983 a_4245_4070# JK_FF_mag_3.nand3_mag_1.IN1 8.64e-19
C984 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK 0.00127f
C985 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 1.9e-21
C986 JK_FF_mag_3.QB a_3117_4070# 0.0811f
C987 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN or_2_mag_0.IN1 0.0405f
C988 Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN 0.00527f
C989 a_2528_240# RST 9.7e-19
C990 CLK RST 0.0304f
C991 Q2 JK_FF_mag_2.nand2_mag_3.IN1 0.00127f
C992 a_1964_240# JK_FF_mag_0.QB 0.00964f
C993 Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN or_2_mag_0.IN1 0.207f
C994 a_4288_1346# VDD 3.14e-19
C995 a_775_2974# JK_FF_mag_2.QB 2.96e-19
C996 a_5006_249# VDD 3.14e-19
C997 a_5129_4070# JK_FF_mag_3.nand3_mag_2.OUT 0.0202f
C998 and_5_mag_0.and2_mag_2.IN2 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.119f
C999 a_1909_4071# JK_FF_mag_2.nand3_mag_2.OUT 0.0731f
C1000 JK_FF_mag_4.nand3_mag_0.OUT Q2 3.91e-20
C1001 JK_FF_mag_3.nand3_mag_0.OUT a_4399_2973# 0.00378f
C1002 Q2 JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C1003 CLK Q3 0.198f
C1004 and_5_mag_0.and2_mag_3.IN2 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.118f
C1005 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN RST 0.00145f
C1006 JK_FF_mag_1.QB Q4 1.34e-19
C1007 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.nand2_mag_3.IN1 0.089f
C1008 a_9908_3052# Q1 0.00479f
C1009 Q4 or_2_mag_0.IN1 0.0716f
C1010 a_3271_2973# JK_FF_mag_3.nand2_mag_4.IN2 4.52e-20
C1011 JK_FF_mag_3.QB CLK 0.311f
C1012 a_7047_3047# CLK 2.26e-19
C1013 a_516_196# JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C1014 a_1339_2974# JK_FF_mag_2.nand3_mag_1.IN1 0.0697f
C1015 JK_FF_mag_1.nand3_mag_1.IN1 a_4442_205# 8.64e-19
C1016 Q2 a_9909_3809# 4.35e-19
C1017 a_8945_3798# Q3 9.22e-21
C1018 Q4 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.3f
C1019 JK_FF_mag_1.nand2_mag_3.IN1 a_3718_205# 1.46e-19
C1020 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C1021 a_4969_4070# JK_FF_mag_3.nand3_mag_2.OUT 0.0731f
C1022 a_1345_4071# JK_FF_mag_2.nand3_mag_2.OUT 9.1e-19
C1023 JK_FF_mag_3.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_3.IN1 1.93e-19
C1024 a_1246_1337# JK_FF_mag_2.nand3_mag_1.OUT 5e-20
C1025 Q2 a_2528_240# 0.0157f
C1026 Q4 RST 0.744f
C1027 JK_FF_mag_0.nand3_mag_1.OUT RST 0.262f
C1028 JK_FF_mag_4.nand3_mag_2.OUT RST 0.0826f
C1029 Q2 CLK 0.324f
C1030 a_5123_2973# CLK 0.0113f
C1031 JK_FF_mag_2.nand3_mag_1.OUT JK_FF_mag_2.QB 0.25f
C1032 Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN or_2_mag_0.GF_INV_MAG_1.IN 2.44e-21
C1033 Q4 a_8078_248# 0.00859f
C1034 JK_FF_mag_4.nand2_mag_1.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 2.66e-19
C1035 JK_FF_mag_4.nand2_mag_3.IN1 Q1 7.52e-19
C1036 JK_FF_mag_4.QB Q4 1.97f
C1037 a_522_1293# VDD 0.00533f
C1038 JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.401f
C1039 a_3681_4070# JK_FF_mag_3.nand2_mag_3.IN1 0.0036f
C1040 a_621_4071# JK_FF_mag_2.nand2_mag_4.IN2 0.069f
C1041 JK_FF_mag_4.QB JK_FF_mag_4.nand3_mag_2.OUT 0.103f
C1042 Q4 Q3 0.259f
C1043 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C1044 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VDD 0.517f
C1045 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_7993_3052# 3.85e-20
C1046 JK_FF_mag_2.QB Q0 0.307f
C1047 Q2 a_8945_3798# 0.0193f
C1048 JK_FF_mag_4.nand3_mag_2.OUT Q3 0.235f
C1049 Q4 a_7047_3047# 0.00353f
C1050 a_3564_1302# VDD 0.00519f
C1051 and_5_mag_0.and2_mag_3.IN2 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 1.97e-19
C1052 JK_FF_mag_3.nand2_mag_3.IN1 JK_FF_mag_2.nand2_mag_3.IN1 0.00229f
C1053 a_4405_4070# JK_FF_mag_3.nand3_mag_2.OUT 9.1e-19
C1054 a_1185_4071# JK_FF_mag_2.nand3_mag_2.OUT 2.88e-20
C1055 JK_FF_mag_4.nand2_mag_1.IN2 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN 2.63e-20
C1056 Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VDD 0.519f
C1057 a_7993_3052# RST 3.66e-19
C1058 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN nand_5_mag_0.GF_INV_MAG_0.IN 5.82e-21
C1059 JK_FF_mag_4.nand3_mag_1.IN1 a_7514_204# 8.64e-19
C1060 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN 0.118f
C1061 a_2063_2974# RST 0.00177f
C1062 VDD Q1 3.73f
C1063 JK_FF_mag_3.nand3_mag_1.IN1 CLK 0.00182f
C1064 a_4963_2973# CLK 0.0102f
C1065 JK_FF_mag_4.nand3_mag_1.OUT JK_FF_mag_4.nand2_mag_4.IN2 0.122f
C1066 JK_FF_mag_4.nand2_mag_1.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 3.68e-19
C1067 a_1909_4071# JK_FF_mag_2.nand2_mag_3.IN1 8.66e-20
C1068 JK_FF_mag_2.nand2_mag_4.IN2 JK_FF_mag_2.nand2_mag_3.IN1 0.321f
C1069 a_7993_3052# Q3 0.0114f
C1070 JK_FF_mag_3.nand3_mag_0.OUT JK_FF_mag_3.nand3_mag_2.OUT 0.00183f
C1071 JK_FF_mag_3.nand2_mag_1.IN2 CLK 1.48e-20
C1072 a_3564_1302# a_3724_1302# 0.0504f
C1073 Q2 Q4 0.195f
C1074 JK_FF_mag_3.QB a_2063_2974# 1.76e-20
C1075 JK_FF_mag_2.nand3_mag_0.OUT JK_FF_mag_2.nand3_mag_2.OUT 0.00183f
C1076 Q2 JK_FF_mag_0.nand3_mag_1.OUT 0.0345f
C1077 JK_FF_mag_2.nand2_mag_1.IN2 JK_FF_mag_2.nand2_mag_4.IN2 8.16e-20
C1078 a_3718_205# RST 0.00189f
C1079 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN 0.00116f
C1080 a_2374_1337# VDD 3.56e-19
C1081 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN and_5_mag_0.and2_mag_3.IN2 0.127f
C1082 a_4245_4070# JK_FF_mag_3.nand3_mag_2.OUT 2.88e-20
C1083 a_1903_2974# RST 0.00132f
C1084 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 a_9908_3052# 0.00347f
C1085 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN 8.99e-19
C1086 a_6630_204# VDD 0.00108f
C1087 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 3.34e-21
C1088 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN 0.12f
C1089 a_4399_2973# CLK 1.4e-19
C1090 a_3718_205# Q3 0.00789f
C1091 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN 1.56e-21
C1092 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_3.nand3_mag_1.OUT 4.98e-19
C1093 CLK JK_FF_mag_3.nand2_mag_3.IN1 0.414f
C1094 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 RST 0.00628f
C1095 Q2 a_7993_3052# 0.00952f
C1096 a_1240_196# JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C1097 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C1098 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN a_9909_3809# 0.069f
C1099 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN 6.85e-19
C1100 JK_FF_mag_3.QB a_1903_2974# 1.35e-20
C1101 a_522_1293# Q1 0.0101f
C1102 JK_FF_mag_0.nand2_mag_1.IN2 Q1 1.48e-20
C1103 a_1810_1337# VDD 3.14e-19
C1104 a_682_1293# JK_FF_mag_0.nand2_mag_3.IN1 0.00119f
C1105 JK_FF_mag_4.QB nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 3.95e-19
C1106 and_5_mag_0.and2_mag_1.IN2 Q0 5.32e-19
C1107 Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN or_2_mag_0.IN1 0.0836f
C1108 a_1339_2974# RST 3.66e-19
C1109 Q3 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0781f
C1110 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN CLK 0.3f
C1111 a_775_2974# JK_FF_mag_0.QB 5e-20
C1112 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN 0.0075f
C1113 Q2 a_3718_205# 0.00216f
C1114 Q0 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.0957f
C1115 a_2374_1337# JK_FF_mag_0.nand2_mag_1.IN2 0.00372f
C1116 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C1117 JK_FF_mag_4.nand3_mag_0.OUT a_7360_1345# 0.00378f
C1118 JK_FF_mag_0.nand2_mag_4.IN2 a_2528_240# 0.00372f
C1119 JK_FF_mag_1.nand2_mag_1.IN2 a_5416_1346# 0.00372f
C1120 a_1246_1337# VDD 3.14e-19
C1121 JK_FF_mag_0.nand3_mag_1.IN1 RST 0.196f
C1122 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_2.nand3_mag_1.IN1 0.00103f
C1123 Q4 Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN 0.00223f
C1124 Q4 JK_FF_mag_3.nand2_mag_3.IN1 6.74e-19
C1125 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VDD 0.385f
C1126 JK_FF_mag_2.QB VDD 0.912f
C1127 and_5_mag_0.VOUT Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN 0.106f
C1128 Q2 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 0.0127f
C1129 JK_FF_mag_1.QB a_4442_205# 0.00696f
C1130 a_8642_248# VSS 0.0675f
C1131 a_8078_248# VSS 0.0676f
C1132 a_7514_204# VSS 0.0343f
C1133 a_7354_204# VSS 0.0881f
C1134 a_6790_204# VSS 0.0343f
C1135 a_6630_204# VSS 0.0881f
C1136 a_5570_249# VSS 0.0675f
C1137 a_5006_249# VSS 0.0676f
C1138 a_4442_205# VSS 0.0343f
C1139 a_4282_205# VSS 0.0881f
C1140 a_3718_205# VSS 0.0343f
C1141 a_3558_205# VSS 0.0881f
C1142 a_2528_240# VSS 0.0686f
C1143 a_1964_240# VSS 0.0687f
C1144 a_1400_196# VSS 0.036f
C1145 a_1240_196# VSS 0.0898f
C1146 a_676_196# VSS 0.036f
C1147 a_516_196# VSS 0.0899f
C1148 Buffer_Delayed1_mag_0.Inverter_delayed_mag_7.IN VSS 0.678f
C1149 Buffer_Delayed1_mag_0.Inverter_delayed_mag_6.IN VSS 0.66f
C1150 Buffer_Delayed1_mag_0.Inverter_delayed_mag_5.IN VSS 0.66f
C1151 Buffer_Delayed1_mag_0.Inverter_delayed_mag_4.IN VSS 0.66f
C1152 Buffer_Delayed1_mag_0.Inverter_delayed_mag_3.IN VSS 0.665f
C1153 Buffer_Delayed1_mag_0.Inverter_delayed_mag_0.IN VSS 0.675f
C1154 Buffer_Delayed1_mag_0.Inverter_delayed_mag_2.IN VSS 0.76f
C1155 JK_FF_mag_4.nand2_mag_4.IN2 VSS 0.416f
C1156 JK_FF_mag_4.nand3_mag_2.OUT VSS 0.54f
C1157 JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.416f
C1158 JK_FF_mag_1.nand3_mag_2.OUT VSS 0.54f
C1159 JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.418f
C1160 JK_FF_mag_0.nand3_mag_2.OUT VSS 0.545f
C1161 Buffer_Delayed1_mag_0.Inverter_delayed_mag_14.IN VSS 0.71f
C1162 Buffer_Delayed1_mag_0.Inverter_delayed_mag_13.IN VSS 0.698f
C1163 Buffer_Delayed1_mag_0.Inverter_delayed_mag_12.IN VSS 0.698f
C1164 Buffer_Delayed1_mag_0.Inverter_delayed_mag_11.IN VSS 0.708f
C1165 Buffer_Delayed1_mag_0.Inverter_delayed_mag_9.IN VSS 0.681f
C1166 a_8488_1345# VSS 0.0676f
C1167 a_7924_1345# VSS 0.0676f
C1168 a_7360_1345# VSS 0.0676f
C1169 a_6796_1301# VSS 0.0343f
C1170 a_6636_1301# VSS 0.0881f
C1171 Buffer_Delayed1_mag_0.Inverter_delayed_mag_8.IN VSS 0.761f
C1172 Buffer_Delayed1_mag_0.Inverter_delayed_mag_1.IN VSS 1.68f
C1173 Buffer_Delayed1_mag_0.Inverter_delayed_mag_10.IN VSS 0.703f
C1174 a_5416_1346# VSS 0.0676f
C1175 a_4852_1346# VSS 0.0676f
C1176 a_4288_1346# VSS 0.0676f
C1177 a_3724_1302# VSS 0.0343f
C1178 a_3564_1302# VSS 0.0881f
C1179 a_2374_1337# VSS 0.0676f
C1180 a_1810_1337# VSS 0.0676f
C1181 a_1246_1337# VSS 0.0676f
C1182 a_682_1293# VSS 0.0343f
C1183 a_522_1293# VSS 0.0881f
C1184 JK_FF_mag_4.nand2_mag_1.IN2 VSS 0.413f
C1185 JK_FF_mag_4.nand2_mag_3.IN1 VSS 0.716f
C1186 JK_FF_mag_4.nand3_mag_1.IN1 VSS 0.723f
C1187 JK_FF_mag_4.nand3_mag_1.OUT VSS 0.808f
C1188 JK_FF_mag_4.nand3_mag_0.OUT VSS 0.507f
C1189 JK_FF_mag_4.QB VSS 0.929f
C1190 JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.412f
C1191 JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.69f
C1192 JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C1193 JK_FF_mag_1.nand3_mag_1.OUT VSS 0.808f
C1194 JK_FF_mag_1.nand3_mag_0.OUT VSS 0.507f
C1195 JK_FF_mag_1.QB VSS 0.886f
C1196 JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.413f
C1197 JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.739f
C1198 JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C1199 JK_FF_mag_0.nand3_mag_1.OUT VSS 0.813f
C1200 JK_FF_mag_0.nand3_mag_0.OUT VSS 0.507f
C1201 JK_FF_mag_0.QB VSS 1.61f
C1202 Vdiv31 VSS 0.315f
C1203 or_2_mag_0.GF_INV_MAG_1.IN VSS 0.602f
C1204 a_11530_2405# VSS 0.0247f
C1205 or_2_mag_0.IN1 VSS 1.37f
C1206 nand_5_mag_0.GF_INV_MAG_0.IN VSS 0.413f
C1207 nand_5_mag_0.and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.446f
C1208 a_9908_3052# VSS 0.073f
C1209 nand_5_mag_0.and_5_mag_0.and2_mag_3.IN2 VSS 0.4f
C1210 nand_5_mag_0.and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.451f
C1211 a_8944_3063# VSS 0.0757f
C1212 nand_5_mag_0.and_5_mag_0.and2_mag_2.IN2 VSS 0.397f
C1213 nand_5_mag_0.and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.443f
C1214 a_7993_3052# VSS 0.073f
C1215 nand_5_mag_0.and_5_mag_0.and2_mag_1.IN2 VSS 0.393f
C1216 nand_5_mag_0.and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.445f
C1217 a_7047_3047# VSS 0.072f
C1218 a_5123_2973# VSS 0.0881f
C1219 a_4963_2973# VSS 0.0343f
C1220 a_4399_2973# VSS 0.0676f
C1221 a_3835_2973# VSS 0.0676f
C1222 a_3271_2973# VSS 0.0676f
C1223 JK_FF_mag_3.nand3_mag_0.OUT VSS 0.507f
C1224 JK_FF_mag_3.nand2_mag_1.IN2 VSS 0.412f
C1225 Q4 VSS 3.04f
C1226 a_2063_2974# VSS 0.0881f
C1227 a_1903_2974# VSS 0.0343f
C1228 a_1339_2974# VSS 0.0676f
C1229 a_775_2974# VSS 0.0676f
C1230 a_211_2974# VSS 0.0676f
C1231 JK_FF_mag_2.nand3_mag_0.OUT VSS 0.506f
C1232 JK_FF_mag_2.nand2_mag_1.IN2 VSS 0.413f
C1233 a_9909_3809# VSS 0.073f
C1234 a_8945_3798# VSS 0.0757f
C1235 a_7994_3809# VSS 0.073f
C1236 and_5_mag_0.VOUT VSS 3.27f
C1237 a_7048_3814# VSS 0.0717f
C1238 and_5_mag_0.and2_mag_3.GF_INV_MAG_0.IN VSS 0.465f
C1239 and_5_mag_0.and2_mag_3.IN2 VSS 0.4f
C1240 and_5_mag_0.and2_mag_2.GF_INV_MAG_0.IN VSS 0.451f
C1241 Q2 VSS 5.04f
C1242 and_5_mag_0.and2_mag_2.IN2 VSS 0.398f
C1243 a_5129_4070# VSS 0.0881f
C1244 a_4969_4070# VSS 0.0343f
C1245 a_4405_4070# VSS 0.0881f
C1246 a_4245_4070# VSS 0.0343f
C1247 a_3681_4070# VSS 0.0676f
C1248 a_3117_4070# VSS 0.0675f
C1249 JK_FF_mag_3.QB VSS 0.887f
C1250 JK_FF_mag_3.nand3_mag_1.OUT VSS 0.807f
C1251 JK_FF_mag_3.nand2_mag_3.IN1 VSS 0.698f
C1252 JK_FF_mag_3.nand2_mag_4.IN2 VSS 0.415f
C1253 and_5_mag_0.and2_mag_1.GF_INV_MAG_0.IN VSS 0.445f
C1254 Q3 VSS 4.36f
C1255 and_5_mag_0.and2_mag_1.IN2 VSS 0.395f
C1256 CLK VSS 2.61f
C1257 JK_FF_mag_3.nand3_mag_2.OUT VSS 0.536f
C1258 JK_FF_mag_3.nand3_mag_1.IN1 VSS 0.722f
C1259 a_2069_4071# VSS 0.0881f
C1260 a_1909_4071# VSS 0.0343f
C1261 a_1345_4071# VSS 0.0881f
C1262 a_1185_4071# VSS 0.0343f
C1263 a_621_4071# VSS 0.0676f
C1264 a_57_4071# VSS 0.0675f
C1265 JK_FF_mag_2.QB VSS 0.923f
C1266 JK_FF_mag_2.nand3_mag_1.OUT VSS 0.807f
C1267 JK_FF_mag_2.nand2_mag_3.IN1 VSS 0.716f
C1268 JK_FF_mag_2.nand2_mag_4.IN2 VSS 0.415f
C1269 JK_FF_mag_2.nand3_mag_2.OUT VSS 0.539f
C1270 RST VSS 5.59f
C1271 JK_FF_mag_2.nand3_mag_1.IN1 VSS 0.722f
C1272 and_5_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.448f
C1273 Q1 VSS 5.56f
C1274 Q0 VSS 3.67f
C1275 VDD VSS 96.6f
C1276 CLK.n0 VSS 0.0044f
C1277 CLK.n1 VSS 0.0114f
C1278 CLK.n2 VSS 0.0139f
C1279 CLK.n3 VSS 0.0116f
C1280 CLK.t0 VSS 0.025f
C1281 CLK.t7 VSS 0.0165f
C1282 CLK.n4 VSS 0.0442f
C1283 CLK.n5 VSS 0.00577f
C1284 CLK.n6 VSS 0.00415f
C1285 CLK.n7 VSS 0.00205f
C1286 CLK.t5 VSS 0.025f
C1287 CLK.t2 VSS 0.0165f
C1288 CLK.n8 VSS 0.0442f
C1289 CLK.n9 VSS 0.00415f
C1290 CLK.n10 VSS 0.00207f
C1291 CLK.n11 VSS 0.00577f
C1292 CLK.n12 VSS 0.00816f
C1293 CLK.n13 VSS 0.0829f
C1294 CLK.n14 VSS 0.0817f
C1295 CLK.n15 VSS 0.0521f
C1296 CLK.t6 VSS 0.0206f
C1297 CLK.t1 VSS 0.00534f
C1298 CLK.n16 VSS 0.0342f
C1299 CLK.n17 VSS 0.00726f
C1300 CLK.n18 VSS 0.00253f
C1301 CLK.n19 VSS 0.0526f
C1302 CLK.n20 VSS 0.0105f
C1303 CLK.n21 VSS 0.00828f
C1304 CLK.n22 VSS 0.00533f
C1305 CLK.n23 VSS 0.00558f
C1306 CLK.n24 VSS 0.00426f
C1307 CLK.n25 VSS 0.00791f
C1308 CLK.n26 VSS 0.19f
C1309 CLK.n27 VSS 0.216f
C1310 CLK.t3 VSS 0.0144f
C1311 CLK.t4 VSS 0.018f
C1312 CLK.n28 VSS 0.0425f
C1313 CLK.n29 VSS 0.309f
C1314 CLK.n30 VSS 0.55f
C1315 CLK.n31 VSS 0.166f
C1316 CLK.n32 VSS 0.0244f
C1317 JK_FF_mag_0.QB.n0 VSS 0.123f
C1318 JK_FF_mag_0.QB.t3 VSS 0.0265f
C1319 JK_FF_mag_0.QB.t5 VSS 0.0332f
C1320 JK_FF_mag_0.QB.n1 VSS 0.0786f
C1321 JK_FF_mag_0.QB.t4 VSS 0.0297f
C1322 JK_FF_mag_0.QB.t6 VSS 0.0466f
C1323 JK_FF_mag_0.QB.n2 VSS 0.0825f
C1324 JK_FF_mag_0.QB.n3 VSS 0.763f
C1325 JK_FF_mag_0.QB.t0 VSS 0.0207f
C1326 JK_FF_mag_0.QB.n4 VSS 0.0207f
C1327 JK_FF_mag_0.QB.n5 VSS 0.0489f
C1328 Q1.t16 VSS 0.035f
C1329 Q1.t14 VSS 0.0231f
C1330 Q1.n0 VSS 0.0621f
C1331 Q1.t13 VSS 0.0201f
C1332 Q1.t15 VSS 0.0252f
C1333 Q1.n1 VSS 0.0596f
C1334 Q1.n2 VSS 0.0614f
C1335 Q1.n3 VSS 0.191f
C1336 Q1.t7 VSS 0.0201f
C1337 Q1.t8 VSS 0.0252f
C1338 Q1.n4 VSS 0.0595f
C1339 Q1.n5 VSS 0.433f
C1340 Q1.n6 VSS 0.584f
C1341 Q1.n7 VSS 1.05f
C1342 Q1.t9 VSS 0.0251f
C1343 Q1.t3 VSS 0.0201f
C1344 Q1.n8 VSS 0.0583f
C1345 Q1.n9 VSS 0.0362f
C1346 Q1.n10 VSS 0.01f
C1347 Q1.t5 VSS 0.0289f
C1348 Q1.t11 VSS 0.00739f
C1349 Q1.n11 VSS 0.0479f
C1350 Q1.n12 VSS 0.0102f
C1351 Q1.n13 VSS 0.0208f
C1352 Q1.n14 VSS 0.00353f
C1353 Q1.n15 VSS 0.00313f
C1354 Q1.n16 VSS 0.0029f
C1355 Q1.n17 VSS 0.00581f
C1356 Q1.t4 VSS 0.0231f
C1357 Q1.t10 VSS 0.035f
C1358 Q1.n18 VSS 0.0618f
C1359 Q1.n19 VSS 0.00797f
C1360 Q1.n20 VSS 0.0113f
C1361 Q1.n21 VSS 0.114f
C1362 Q1.n22 VSS 0.116f
C1363 Q1.n23 VSS 0.00581f
C1364 Q1.t6 VSS 0.0231f
C1365 Q1.t12 VSS 0.035f
C1366 Q1.n24 VSS 0.0618f
C1367 Q1.n25 VSS 0.00797f
C1368 Q1.n26 VSS 0.00287f
C1369 Q1.n27 VSS 0.0701f
C1370 Q1.n28 VSS 0.209f
C1371 Q1.t2 VSS 0.0191f
C1372 Q1.t0 VSS 0.0157f
C1373 Q1.n29 VSS 0.0157f
C1374 Q1.n30 VSS 0.0377f
C1375 Q1.n31 VSS 0.118f
C1376 Q1.n32 VSS 0.014f
C1377 Q1.n33 VSS 0.153f
C1378 Q1.n34 VSS 0.364f
C1379 Q1.n35 VSS 0.789f
C1380 Q1.n36 VSS 0.029f
C1381 Q4.n0 VSS 0.0185f
C1382 Q4.t1 VSS 0.0152f
C1383 Q4.n1 VSS 0.0152f
C1384 Q4.n2 VSS 0.0419f
C1385 Q4.n3 VSS 0.135f
C1386 Q4.t4 VSS 0.0557f
C1387 Q4.t7 VSS 0.00804f
C1388 Q4.n4 VSS 0.0464f
C1389 Q4.n5 VSS 0.234f
C1390 Q4.t8 VSS 0.0195f
C1391 Q4.t9 VSS 0.0244f
C1392 Q4.n6 VSS 0.0578f
C1393 Q4.n7 VSS 0.0596f
C1394 Q4.n8 VSS 0.0926f
C1395 Q4.n9 VSS 0.703f
C1396 Q4.t5 VSS 0.0224f
C1397 Q4.t6 VSS 0.034f
C1398 Q4.n10 VSS 0.0603f
C1399 Q4.n11 VSS 0.237f
C1400 Q4.t10 VSS 0.0195f
C1401 Q4.t3 VSS 0.0244f
C1402 Q4.n12 VSS 0.0565f
C1403 Q4.n13 VSS 0.0351f
C1404 Q4.n14 VSS 0.45f
C1405 Q4.n15 VSS 0.205f
C1406 Q3.t15 VSS 0.0264f
C1407 Q3.t16 VSS 0.0401f
C1408 Q3.n0 VSS 0.0711f
C1409 Q3.n1 VSS 0.279f
C1410 Q3.t5 VSS 0.023f
C1411 Q3.t12 VSS 0.0288f
C1412 Q3.n2 VSS 0.0666f
C1413 Q3.n3 VSS 0.0414f
C1414 Q3.n4 VSS 0.515f
C1415 Q3.n5 VSS 0.0222f
C1416 Q3.n6 VSS 0.00403f
C1417 Q3.t3 VSS 0.023f
C1418 Q3.t11 VSS 0.0288f
C1419 Q3.n7 VSS 0.066f
C1420 Q3.n8 VSS 0.0272f
C1421 Q3.n9 VSS 0.00417f
C1422 Q3.n10 VSS 0.205f
C1423 Q3.n11 VSS 0.31f
C1424 Q3.t8 VSS 0.023f
C1425 Q3.t10 VSS 0.0288f
C1426 Q3.n12 VSS 0.0682f
C1427 Q3.n13 VSS 0.33f
C1428 Q3.n14 VSS 0.382f
C1429 Q3.n15 VSS 0.724f
C1430 Q3.n16 VSS 0.0115f
C1431 Q3.t6 VSS 0.0331f
C1432 Q3.t14 VSS 0.00846f
C1433 Q3.n17 VSS 0.0548f
C1434 Q3.n18 VSS 0.0116f
C1435 Q3.n19 VSS 0.0238f
C1436 Q3.n20 VSS 0.00404f
C1437 Q3.n21 VSS 0.00358f
C1438 Q3.n22 VSS 0.00332f
C1439 Q3.n23 VSS 0.00665f
C1440 Q3.t9 VSS 0.0264f
C1441 Q3.t13 VSS 0.0401f
C1442 Q3.n24 VSS 0.0707f
C1443 Q3.n25 VSS 0.00912f
C1444 Q3.n26 VSS 0.0129f
C1445 Q3.n27 VSS 0.131f
C1446 Q3.n28 VSS 0.133f
C1447 Q3.n29 VSS 0.00665f
C1448 Q3.t4 VSS 0.0264f
C1449 Q3.t7 VSS 0.0401f
C1450 Q3.n30 VSS 0.0707f
C1451 Q3.n31 VSS 0.00912f
C1452 Q3.n32 VSS 0.00328f
C1453 Q3.n33 VSS 0.0802f
C1454 Q3.n34 VSS 0.113f
C1455 Q3.n35 VSS 0.368f
C1456 Q3.n36 VSS 0.187f
C1457 Q3.n37 VSS 0.0218f
C1458 Q3.t0 VSS 0.018f
C1459 Q3.n38 VSS 0.018f
C1460 Q3.n39 VSS 0.0494f
C1461 Q3.n40 VSS 0.159f
C1462 Q3.n41 VSS 0.00887f
C1463 Q2.t9 VSS 0.0332f
C1464 Q2.t12 VSS 0.0416f
C1465 Q2.n0 VSS 0.0985f
C1466 Q2.n1 VSS 0.477f
C1467 Q2.n2 VSS 0.0317f
C1468 Q2.n3 VSS 0.00582f
C1469 Q2.t16 VSS 0.0332f
C1470 Q2.t3 VSS 0.0416f
C1471 Q2.n4 VSS 0.0953f
C1472 Q2.n5 VSS 0.0392f
C1473 Q2.n6 VSS 0.00602f
C1474 Q2.n7 VSS 0.296f
C1475 Q2.n8 VSS 0.291f
C1476 Q2.n9 VSS 1.47f
C1477 Q2.n10 VSS 0.0048f
C1478 Q2.n11 VSS 0.0096f
C1479 Q2.t10 VSS 0.0381f
C1480 Q2.t11 VSS 0.0579f
C1481 Q2.n12 VSS 0.102f
C1482 Q2.n13 VSS 0.0132f
C1483 Q2.n14 VSS 0.0187f
C1484 Q2.n15 VSS 0.189f
C1485 Q2.n16 VSS 0.192f
C1486 Q2.n17 VSS 0.0096f
C1487 Q2.t5 VSS 0.0381f
C1488 Q2.t8 VSS 0.0579f
C1489 Q2.n18 VSS 0.102f
C1490 Q2.n19 VSS 0.0132f
C1491 Q2.n20 VSS 0.00474f
C1492 Q2.n21 VSS 0.121f
C1493 Q2.n22 VSS 0.12f
C1494 Q2.t6 VSS 0.0478f
C1495 Q2.t13 VSS 0.0122f
C1496 Q2.n23 VSS 0.0791f
C1497 Q2.n24 VSS 0.0168f
C1498 Q2.n25 VSS 0.00584f
C1499 Q2.n26 VSS 0.0344f
C1500 Q2.n27 VSS 0.106f
C1501 Q2.t7 VSS 0.0381f
C1502 Q2.t15 VSS 0.0579f
C1503 Q2.n28 VSS 0.103f
C1504 Q2.n29 VSS 0.403f
C1505 Q2.t4 VSS 0.0332f
C1506 Q2.t14 VSS 0.0416f
C1507 Q2.n30 VSS 0.0963f
C1508 Q2.n31 VSS 0.0598f
C1509 Q2.n32 VSS 0.75f
C1510 Q2.n33 VSS 0.28f
C1511 Q2.n34 VSS 1.47f
C1512 Q2.n35 VSS 0.0315f
C1513 Q2.t1 VSS 0.026f
C1514 Q2.n36 VSS 0.026f
C1515 Q2.n37 VSS 0.0713f
C1516 Q2.n38 VSS 0.229f
C1517 Q2.n39 VSS 0.0112f
C1518 RST.n0 VSS 0.131f
C1519 RST.t6 VSS 0.0145f
C1520 RST.t2 VSS 0.00954f
C1521 RST.n1 VSS 0.0256f
C1522 RST.n2 VSS 0.00348f
C1523 RST.n3 VSS 0.00213f
C1524 RST.n4 VSS 0.00118f
C1525 RST.n5 VSS 0.00261f
C1526 RST.n6 VSS 0.0016f
C1527 RST.n7 VSS 0.00653f
C1528 RST.n8 VSS 0.111f
C1529 RST.n9 VSS 0.00473f
C1530 RST.n10 VSS 0.00169f
C1531 RST.n11 VSS 0.00204f
C1532 RST.n12 VSS 0.00445f
C1533 RST.t11 VSS 0.0145f
C1534 RST.t9 VSS 0.00954f
C1535 RST.n13 VSS 0.0256f
C1536 RST.n14 VSS 0.00352f
C1537 RST.n15 VSS 0.00183f
C1538 RST.n16 VSS 0.00131f
C1539 RST.n17 VSS 1.41e-19
C1540 RST.n18 VSS 0.00637f
C1541 RST.n19 VSS 1.41e-19
C1542 RST.n20 VSS 0.0935f
C1543 RST.n21 VSS 0.297f
C1544 RST.t5 VSS 0.00954f
C1545 RST.t8 VSS 0.0145f
C1546 RST.n22 VSS 0.0256f
C1547 RST.n23 VSS 0.00449f
C1548 RST.n24 VSS 0.00171f
C1549 RST.n25 VSS 0.00526f
C1550 RST.n26 VSS 0.00628f
C1551 RST.t3 VSS 0.00954f
C1552 RST.t4 VSS 0.0145f
C1553 RST.n27 VSS 0.0256f
C1554 RST.n28 VSS 0.141f
C1555 RST.n29 VSS 0.248f
C1556 RST.n30 VSS 0.0872f
C1557 RST.t7 VSS 0.00954f
C1558 RST.t10 VSS 0.0145f
C1559 RST.n31 VSS 0.0256f
C1560 RST.n32 VSS 0.0683f
C1561 RST.n33 VSS 0.319f
C1562 RST.n34 VSS 1f
C1563 RST.n35 VSS 0.81f
C1564 RST.n36 VSS 0.00983f
C1565 RST.n37 VSS 0.00488f
C1566 RST.n38 VSS 0.0162f
C1567 RST.n39 VSS 0.0561f
C1568 RST.n40 VSS 0.0104f
C1569 RST.n41 VSS 0.00487f
C1570 RST.n42 VSS 0.0951f
C1571 RST.n43 VSS 0.112f
C1572 VDD.t240 VSS 0.00585f
C1573 VDD.t258 VSS 0.0024f
C1574 VDD.n0 VSS 0.0024f
C1575 VDD.n1 VSS 0.00525f
C1576 VDD.t137 VSS 0.0772f
C1577 VDD.n2 VSS 0.00584f
C1578 VDD.n3 VSS 0.0383f
C1579 VDD.n4 VSS 0.00584f
C1580 VDD.t1 VSS 0.00585f
C1581 VDD.t83 VSS 0.0491f
C1582 VDD.t332 VSS 0.0461f
C1583 VDD.n5 VSS 0.00584f
C1584 VDD.n6 VSS 0.0373f
C1585 VDD.t259 VSS 0.0761f
C1586 VDD.t196 VSS 0.00585f
C1587 VDD.t63 VSS 0.00582f
C1588 VDD.n7 VSS 0.00582f
C1589 VDD.n8 VSS 0.0321f
C1590 VDD.t291 VSS 0.0801f
C1591 VDD.n9 VSS 0.00582f
C1592 VDD.t329 VSS 0.00582f
C1593 VDD.n10 VSS 0.00582f
C1594 VDD.n11 VSS 0.0319f
C1595 VDD.t328 VSS 0.0977f
C1596 VDD.n12 VSS 0.0399f
C1597 VDD.t288 VSS 0.0977f
C1598 VDD.n13 VSS 0.0834f
C1599 VDD.n14 VSS 0.0838f
C1600 VDD.n15 VSS 0.00582f
C1601 VDD.t223 VSS 0.00582f
C1602 VDD.n16 VSS 0.0152f
C1603 VDD.n17 VSS 0.00582f
C1604 VDD.t256 VSS 0.00582f
C1605 VDD.t197 VSS 0.122f
C1606 VDD.n18 VSS 0.0152f
C1607 VDD.n19 VSS 0.00614f
C1608 VDD.t295 VSS 0.00582f
C1609 VDD.n20 VSS 0.00582f
C1610 VDD.n21 VSS 0.042f
C1611 VDD.n22 VSS 0.0295f
C1612 VDD.n23 VSS 0.0152f
C1613 VDD.t294 VSS 0.151f
C1614 VDD.t49 VSS 0.151f
C1615 VDD.n24 VSS 0.0152f
C1616 VDD.t64 VSS 0.151f
C1617 VDD.t255 VSS 0.151f
C1618 VDD.n25 VSS 0.0152f
C1619 VDD.n26 VSS 0.0295f
C1620 VDD.n27 VSS 0.042f
C1621 VDD.t92 VSS 0.00582f
C1622 VDD.n28 VSS 0.00582f
C1623 VDD.n29 VSS 0.042f
C1624 VDD.n30 VSS 0.0295f
C1625 VDD.n31 VSS 0.0152f
C1626 VDD.t91 VSS 0.151f
C1627 VDD.t214 VSS 0.15f
C1628 VDD.n32 VSS 0.0152f
C1629 VDD.t222 VSS 0.0715f
C1630 VDD.n33 VSS 0.0152f
C1631 VDD.n34 VSS 0.0292f
C1632 VDD.n35 VSS 0.0295f
C1633 VDD.t192 VSS 0.0968f
C1634 VDD.n36 VSS 0.0528f
C1635 VDD.t221 VSS 0.00582f
C1636 VDD.n37 VSS 0.0358f
C1637 VDD.t220 VSS 0.0968f
C1638 VDD.n38 VSS 0.0488f
C1639 VDD.n39 VSS 0.0262f
C1640 VDD.n40 VSS 0.0415f
C1641 VDD.n41 VSS 0.0393f
C1642 VDD.n42 VSS 0.0322f
C1643 VDD.n43 VSS 0.0306f
C1644 VDD.t254 VSS 0.00582f
C1645 VDD.n44 VSS 0.0306f
C1646 VDD.n45 VSS 0.0317f
C1647 VDD.t253 VSS 0.139f
C1648 VDD.t300 VSS 0.133f
C1649 VDD.t62 VSS 0.111f
C1650 VDD.n46 VSS 0.0335f
C1651 VDD.n47 VSS 0.0472f
C1652 VDD.n48 VSS 0.00584f
C1653 VDD.t317 VSS 0.0761f
C1654 VDD.n49 VSS 0.0363f
C1655 VDD.t75 VSS 0.00585f
C1656 VDD.n50 VSS 0.00584f
C1657 VDD.t74 VSS 0.0705f
C1658 VDD.t322 VSS 0.0772f
C1659 VDD.n51 VSS 0.0363f
C1660 VDD.t136 VSS 0.00585f
C1661 VDD.t126 VSS 0.0024f
C1662 VDD.n52 VSS 0.0024f
C1663 VDD.n53 VSS 0.00525f
C1664 VDD.t135 VSS 0.0705f
C1665 VDD.t125 VSS 0.086f
C1666 VDD.t154 VSS 0.04f
C1667 VDD.n54 VSS 0.0363f
C1668 VDD.t360 VSS 0.00585f
C1669 VDD.t313 VSS 0.0024f
C1670 VDD.n55 VSS 0.0024f
C1671 VDD.n56 VSS 0.00525f
C1672 VDD.t359 VSS 0.0705f
C1673 VDD.t312 VSS 0.086f
C1674 VDD.t179 VSS 0.04f
C1675 VDD.t11 VSS 0.0703f
C1676 VDD.n57 VSS 0.0363f
C1677 VDD.t12 VSS 0.00585f
C1678 VDD.t27 VSS 0.00502f
C1679 VDD.t367 VSS 0.0038f
C1680 VDD.n58 VSS 0.00984f
C1681 VDD.n59 VSS 0.00906f
C1682 VDD.t10 VSS 0.00502f
C1683 VDD.t372 VSS 0.0038f
C1684 VDD.n60 VSS 0.00985f
C1685 VDD.n61 VSS 0.00735f
C1686 VDD.n62 VSS 0.0469f
C1687 VDD.n63 VSS 0.0272f
C1688 VDD.n64 VSS 0.0181f
C1689 VDD.n65 VSS 0.0333f
C1690 VDD.n66 VSS 0.0342f
C1691 VDD.n67 VSS 0.0181f
C1692 VDD.n68 VSS 0.0333f
C1693 VDD.n69 VSS 0.0341f
C1694 VDD.n70 VSS 0.0202f
C1695 VDD.n71 VSS 0.029f
C1696 VDD.n72 VSS 0.0269f
C1697 VDD.n73 VSS 0.0202f
C1698 VDD.n74 VSS 0.0214f
C1699 VDD.n75 VSS 0.0478f
C1700 VDD.t56 VSS 0.0059f
C1701 VDD.n76 VSS 0.0161f
C1702 VDD.t287 VSS 0.00585f
C1703 VDD.t286 VSS 0.0498f
C1704 VDD.t176 VSS 0.0461f
C1705 VDD.n77 VSS 0.00584f
C1706 VDD.t228 VSS 0.00582f
C1707 VDD.t82 VSS 0.00585f
C1708 VDD.n78 VSS 0.0388f
C1709 VDD.t227 VSS 0.0514f
C1710 VDD.t274 VSS 0.0769f
C1711 VDD.n79 VSS 0.00584f
C1712 VDD.t336 VSS 0.00582f
C1713 VDD.t358 VSS 0.00582f
C1714 VDD.n80 VSS 0.033f
C1715 VDD.t357 VSS 0.055f
C1716 VDD.t311 VSS 0.014f
C1717 VDD.t356 VSS 0.00582f
C1718 VDD.n81 VSS 0.0313f
C1719 VDD.t355 VSS 0.0518f
C1720 VDD.n82 VSS 0.0614f
C1721 VDD.t204 VSS 0.0551f
C1722 VDD.t310 VSS 0.0894f
C1723 VDD.n83 VSS 0.043f
C1724 VDD.n84 VSS 0.0311f
C1725 VDD.n85 VSS 0.026f
C1726 VDD.t184 VSS 0.0521f
C1727 VDD.n86 VSS 0.0539f
C1728 VDD.t185 VSS 0.00582f
C1729 VDD.n87 VSS 0.00584f
C1730 VDD.t110 VSS 0.0461f
C1731 VDD.n88 VSS 0.0363f
C1732 VDD.t48 VSS 0.00585f
C1733 VDD.t47 VSS 0.0686f
C1734 VDD.t72 VSS 0.0513f
C1735 VDD.n89 VSS 0.0561f
C1736 VDD.t73 VSS 0.00582f
C1737 VDD.n90 VSS 0.00584f
C1738 VDD.t349 VSS 0.0461f
C1739 VDD.n91 VSS 0.0363f
C1740 VDD.t263 VSS 0.00585f
C1741 VDD.t262 VSS 0.0698f
C1742 VDD.t308 VSS 0.0496f
C1743 VDD.n92 VSS 0.054f
C1744 VDD.t309 VSS 0.00582f
C1745 VDD.n93 VSS 0.00584f
C1746 VDD.t165 VSS 0.0461f
C1747 VDD.n94 VSS 0.0363f
C1748 VDD.t189 VSS 0.00585f
C1749 VDD.t188 VSS 0.0699f
C1750 VDD.t296 VSS 0.049f
C1751 VDD.n95 VSS 0.0536f
C1752 VDD.t297 VSS 0.00582f
C1753 VDD.n96 VSS 0.00584f
C1754 VDD.t277 VSS 0.0461f
C1755 VDD.t237 VSS 0.0703f
C1756 VDD.n97 VSS 0.0363f
C1757 VDD.t238 VSS 0.00619f
C1758 VDD.n98 VSS 0.0237f
C1759 VDD.n99 VSS 0.0358f
C1760 VDD.n100 VSS 0.0314f
C1761 VDD.n101 VSS 0.0366f
C1762 VDD.n102 VSS 0.024f
C1763 VDD.n103 VSS 0.0364f
C1764 VDD.n104 VSS 0.0319f
C1765 VDD.n105 VSS 0.039f
C1766 VDD.n106 VSS 0.0246f
C1767 VDD.n107 VSS 0.0377f
C1768 VDD.n108 VSS 0.0329f
C1769 VDD.n109 VSS 0.0388f
C1770 VDD.n110 VSS 0.024f
C1771 VDD.n111 VSS 0.0364f
C1772 VDD.n112 VSS 0.0319f
C1773 VDD.n113 VSS 0.106f
C1774 VDD.n114 VSS 0.0619f
C1775 VDD.t335 VSS 0.0542f
C1776 VDD.n115 VSS 0.0624f
C1777 VDD.n116 VSS 0.0319f
C1778 VDD.n117 VSS 0.0364f
C1779 VDD.n118 VSS 0.024f
C1780 VDD.n119 VSS 0.0363f
C1781 VDD.t81 VSS 0.0686f
C1782 VDD.n120 VSS 0.0561f
C1783 VDD.n121 VSS 0.0329f
C1784 VDD.n122 VSS 0.0377f
C1785 VDD.n123 VSS 0.0241f
C1786 VDD.n124 VSS 0.0363f
C1787 VDD.t55 VSS 0.0698f
C1788 VDD.n125 VSS 0.054f
C1789 VDD.n126 VSS 0.00584f
C1790 VDD.n127 VSS 0.038f
C1791 VDD.n128 VSS 0.0417f
C1792 VDD.n129 VSS 0.0562f
C1793 VDD.n130 VSS 0.0438f
C1794 VDD.n131 VSS 0.00556f
C1795 VDD.n132 VSS 0.00853f
C1796 VDD.n133 VSS 0.0161f
C1797 VDD.n134 VSS 0.0172f
C1798 VDD.n135 VSS 0.0363f
C1799 VDD.t195 VSS 0.0705f
C1800 VDD.t325 VSS 0.0772f
C1801 VDD.t127 VSS 0.0705f
C1802 VDD.n136 VSS 0.0363f
C1803 VDD.t191 VSS 0.00585f
C1804 VDD.t128 VSS 0.00585f
C1805 VDD.t84 VSS 0.00842f
C1806 VDD.n137 VSS 0.0113f
C1807 VDD.n138 VSS 0.0533f
C1808 VDD.n139 VSS 0.0302f
C1809 VDD.n140 VSS 0.0212f
C1810 VDD.n141 VSS 0.0302f
C1811 VDD.n142 VSS 0.0363f
C1812 VDD.t190 VSS 0.0699f
C1813 VDD.n143 VSS 0.0536f
C1814 VDD.t314 VSS 0.0461f
C1815 VDD.t239 VSS 0.0703f
C1816 VDD.n144 VSS 0.0363f
C1817 VDD.n145 VSS 0.0388f
C1818 VDD.n146 VSS 0.0371f
C1819 VDD.n147 VSS 0.0223f
C1820 VDD.n148 VSS 0.0395f
C1821 VDD.n149 VSS 0.0363f
C1822 VDD.t0 VSS 0.0705f
C1823 VDD.t257 VSS 0.086f
C1824 VDD.t168 VSS 0.04f
C1825 VDD.n150 VSS 0.0363f
C1826 VDD.t29 VSS 0.00585f
C1827 VDD.t175 VSS 0.00582f
C1828 VDD.n151 VSS 0.00584f
C1829 VDD.t171 VSS 0.0761f
C1830 VDD.n152 VSS 0.0363f
C1831 VDD.t321 VSS 0.00585f
C1832 VDD.n153 VSS 0.00584f
C1833 VDD.t320 VSS 0.0705f
C1834 VDD.t85 VSS 0.0772f
C1835 VDD.n154 VSS 0.0363f
C1836 VDD.t144 VSS 0.00585f
C1837 VDD.t7 VSS 0.0024f
C1838 VDD.n155 VSS 0.0024f
C1839 VDD.n156 VSS 0.00525f
C1840 VDD.t143 VSS 0.0705f
C1841 VDD.t6 VSS 0.086f
C1842 VDD.t157 VSS 0.04f
C1843 VDD.n157 VSS 0.0363f
C1844 VDD.t71 VSS 0.00585f
C1845 VDD.t183 VSS 0.0024f
C1846 VDD.n158 VSS 0.0024f
C1847 VDD.n159 VSS 0.00525f
C1848 VDD.t70 VSS 0.0705f
C1849 VDD.t182 VSS 0.086f
C1850 VDD.t352 VSS 0.04f
C1851 VDD.t38 VSS 0.0703f
C1852 VDD.n160 VSS 0.0363f
C1853 VDD.t39 VSS 0.00585f
C1854 VDD.t34 VSS 0.00502f
C1855 VDD.t366 VSS 0.0038f
C1856 VDD.n161 VSS 0.00985f
C1857 VDD.n162 VSS 0.00922f
C1858 VDD.t37 VSS 0.00502f
C1859 VDD.t365 VSS 0.0038f
C1860 VDD.n163 VSS 0.00987f
C1861 VDD.n164 VSS 0.0074f
C1862 VDD.n165 VSS 0.0386f
C1863 VDD.n166 VSS 0.0272f
C1864 VDD.n167 VSS 0.0181f
C1865 VDD.n168 VSS 0.0333f
C1866 VDD.n169 VSS 0.0342f
C1867 VDD.n170 VSS 0.0181f
C1868 VDD.n171 VSS 0.0333f
C1869 VDD.n172 VSS 0.0341f
C1870 VDD.n173 VSS 0.0202f
C1871 VDD.n174 VSS 0.029f
C1872 VDD.n175 VSS 0.0269f
C1873 VDD.n176 VSS 0.0202f
C1874 VDD.n177 VSS 0.052f
C1875 VDD.t113 VSS 0.0517f
C1876 VDD.n178 VSS 0.0543f
C1877 VDD.n179 VSS 0.00734f
C1878 VDD.n180 VSS 0.00584f
C1879 VDD.t149 VSS 0.0761f
C1880 VDD.n181 VSS 0.0363f
C1881 VDD.n182 VSS 0.00585f
C1882 VDD.t331 VSS 0.00585f
C1883 VDD.t21 VSS 0.0401f
C1884 VDD.n183 VSS 0.0363f
C1885 VDD.n184 VSS 0.00584f
C1886 VDD.t117 VSS 0.0024f
C1887 VDD.n185 VSS 0.0024f
C1888 VDD.n186 VSS 0.00525f
C1889 VDD.t330 VSS 0.0705f
C1890 VDD.t88 VSS 0.0772f
C1891 VDD.n187 VSS 0.0363f
C1892 VDD.t9 VSS 0.00585f
C1893 VDD.n188 VSS 0.00585f
C1894 VDD.n189 VSS 0.00584f
C1895 VDD.t116 VSS 0.0398f
C1896 VDD.t305 VSS 0.086f
C1897 VDD.t224 VSS 0.0706f
C1898 VDD.n190 VSS 0.0363f
C1899 VDD.t8 VSS 0.0705f
C1900 VDD.t140 VSS 0.0772f
C1901 VDD.n191 VSS 0.0363f
C1902 VDD.t61 VSS 0.00584f
C1903 VDD.t338 VSS 0.00585f
C1904 VDD.n192 VSS 0.00585f
C1905 VDD.t60 VSS 0.077f
C1906 VDD.t99 VSS 0.0706f
C1907 VDD.n193 VSS 0.0363f
C1908 VDD.t148 VSS 0.0024f
C1909 VDD.n194 VSS 0.0024f
C1910 VDD.n195 VSS 0.00525f
C1911 VDD.t211 VSS 0.00584f
C1912 VDD.t337 VSS 0.0705f
C1913 VDD.t147 VSS 0.086f
C1914 VDD.t342 VSS 0.04f
C1915 VDD.n196 VSS 0.0363f
C1916 VDD.n197 VSS 0.00585f
C1917 VDD.t36 VSS 0.00585f
C1918 VDD.t210 VSS 0.077f
C1919 VDD.t105 VSS 0.0706f
C1920 VDD.t303 VSS 0.0759f
C1921 VDD.n198 VSS 0.0363f
C1922 VDD.t304 VSS 0.00584f
C1923 VDD.t346 VSS 0.00735f
C1924 VDD.t345 VSS 0.0516f
C1925 VDD.t35 VSS 0.04f
C1926 VDD.n199 VSS 0.0543f
C1927 VDD.n200 VSS 0.00584f
C1928 VDD.t339 VSS 0.0761f
C1929 VDD.n201 VSS 0.0363f
C1930 VDD.t187 VSS 0.00585f
C1931 VDD.n202 VSS 0.00584f
C1932 VDD.t186 VSS 0.0705f
C1933 VDD.t132 VSS 0.0772f
C1934 VDD.n203 VSS 0.0363f
C1935 VDD.t77 VSS 0.00585f
C1936 VDD.t201 VSS 0.0024f
C1937 VDD.n204 VSS 0.0024f
C1938 VDD.n205 VSS 0.00525f
C1939 VDD.t76 VSS 0.0705f
C1940 VDD.t200 VSS 0.086f
C1941 VDD.t160 VSS 0.04f
C1942 VDD.n206 VSS 0.0363f
C1943 VDD.t146 VSS 0.00585f
C1944 VDD.t348 VSS 0.0024f
C1945 VDD.n207 VSS 0.0024f
C1946 VDD.n208 VSS 0.00525f
C1947 VDD.t145 VSS 0.0705f
C1948 VDD.t347 VSS 0.086f
C1949 VDD.t266 VSS 0.04f
C1950 VDD.t14 VSS 0.0703f
C1951 VDD.n209 VSS 0.0363f
C1952 VDD.t15 VSS 0.00585f
C1953 VDD.t24 VSS 0.00502f
C1954 VDD.t371 VSS 0.0038f
C1955 VDD.n210 VSS 0.00985f
C1956 VDD.n211 VSS 0.00814f
C1957 VDD.t13 VSS 0.00502f
C1958 VDD.t362 VSS 0.0038f
C1959 VDD.n212 VSS 0.00985f
C1960 VDD.n213 VSS 0.00783f
C1961 VDD.n214 VSS 0.0401f
C1962 VDD.n215 VSS 0.0272f
C1963 VDD.n216 VSS 0.0181f
C1964 VDD.n217 VSS 0.0333f
C1965 VDD.n218 VSS 0.0342f
C1966 VDD.n219 VSS 0.0181f
C1967 VDD.n220 VSS 0.0333f
C1968 VDD.n221 VSS 0.0341f
C1969 VDD.n222 VSS 0.0202f
C1970 VDD.n223 VSS 0.029f
C1971 VDD.n224 VSS 0.0269f
C1972 VDD.n225 VSS 0.0202f
C1973 VDD.n226 VSS 0.0528f
C1974 VDD.t234 VSS 0.0517f
C1975 VDD.n227 VSS 0.0543f
C1976 VDD.n228 VSS 0.00734f
C1977 VDD.n229 VSS 0.00584f
C1978 VDD.t245 VSS 0.0614f
C1979 VDD.n230 VSS 0.0313f
C1980 VDD.n231 VSS 0.00585f
C1981 VDD.t119 VSS 0.00585f
C1982 VDD.t31 VSS 0.0401f
C1983 VDD.n232 VSS 0.0363f
C1984 VDD.n233 VSS 0.00584f
C1985 VDD.t242 VSS 0.0024f
C1986 VDD.n234 VSS 0.0024f
C1987 VDD.n235 VSS 0.00525f
C1988 VDD.t118 VSS 0.0561f
C1989 VDD.t129 VSS 0.0614f
C1990 VDD.n236 VSS 0.0313f
C1991 VDD.t203 VSS 0.00585f
C1992 VDD.n237 VSS 0.00585f
C1993 VDD.n238 VSS 0.00584f
C1994 VDD.t241 VSS 0.0398f
C1995 VDD.t207 VSS 0.086f
C1996 VDD.t52 VSS 0.0706f
C1997 VDD.n239 VSS 0.0363f
C1998 VDD.n240 VSS 0.0313f
C1999 VDD.t124 VSS 0.00584f
C2000 VDD.t299 VSS 0.00585f
C2001 VDD.n241 VSS 0.00585f
C2002 VDD.t123 VSS 0.077f
C2003 VDD.t96 VSS 0.0706f
C2004 VDD.n242 VSS 0.0363f
C2005 VDD.t249 VSS 0.0024f
C2006 VDD.n243 VSS 0.0024f
C2007 VDD.n244 VSS 0.00525f
C2008 VDD.t3 VSS 0.00584f
C2009 VDD.t298 VSS 0.0561f
C2010 VDD.t248 VSS 0.0684f
C2011 VDD.t271 VSS 0.0318f
C2012 VDD.n245 VSS 0.0313f
C2013 VDD.n246 VSS 0.00585f
C2014 VDD.t26 VSS 0.00585f
C2015 VDD.t2 VSS 0.077f
C2016 VDD.t44 VSS 0.0706f
C2017 VDD.t205 VSS 0.0759f
C2018 VDD.n247 VSS 0.0363f
C2019 VDD.t206 VSS 0.00584f
C2020 VDD.t270 VSS 0.00735f
C2021 VDD.t25 VSS 0.0318f
C2022 VDD.t202 VSS 0.0415f
C2023 VDD.t78 VSS 0.0269f
C2024 VDD.n248 VSS 0.162f
C2025 VDD.n249 VSS 0.0896f
C2026 VDD.t269 VSS 0.0644f
C2027 VDD.t265 VSS 0.00584f
C2028 VDD.t120 VSS 0.0706f
C2029 VDD.n250 VSS 0.00585f
C2030 VDD.t164 VSS 0.0024f
C2031 VDD.n251 VSS 0.0024f
C2032 VDD.n252 VSS 0.00525f
C2033 VDD.n253 VSS 0.00585f
C2034 VDD.n254 VSS 0.0342f
C2035 VDD.t17 VSS 0.0704f
C2036 VDD.n255 VSS 0.00585f
C2037 VDD.t374 VSS 0.0038f
C2038 VDD.t16 VSS 0.00502f
C2039 VDD.n256 VSS 0.00986f
C2040 VDD.t368 VSS 0.0038f
C2041 VDD.t30 VSS 0.00502f
C2042 VDD.n257 VSS 0.00979f
C2043 VDD.n258 VSS 0.00149f
C2044 VDD.n259 VSS 0.00887f
C2045 VDD.n260 VSS 0.0484f
C2046 VDD.n261 VSS 0.0273f
C2047 VDD.t233 VSS 0.0024f
C2048 VDD.n262 VSS 0.0024f
C2049 VDD.n263 VSS 0.00525f
C2050 VDD.n264 VSS 0.0333f
C2051 VDD.n265 VSS 0.0181f
C2052 VDD.n266 VSS 0.0363f
C2053 VDD.t232 VSS 0.0398f
C2054 VDD.t280 VSS 0.086f
C2055 VDD.t250 VSS 0.0706f
C2056 VDD.t93 VSS 0.086f
C2057 VDD.t163 VSS 0.0398f
C2058 VDD.n267 VSS 0.0363f
C2059 VDD.n268 VSS 0.0181f
C2060 VDD.n269 VSS 0.0333f
C2061 VDD.n270 VSS 0.034f
C2062 VDD.t5 VSS 0.00584f
C2063 VDD.n271 VSS 0.00585f
C2064 VDD.n272 VSS 0.0269f
C2065 VDD.n273 VSS 0.029f
C2066 VDD.n274 VSS 0.0202f
C2067 VDD.n275 VSS 0.0363f
C2068 VDD.t4 VSS 0.077f
C2069 VDD.t283 VSS 0.0706f
C2070 VDD.t264 VSS 0.0759f
C2071 VDD.n276 VSS 0.0363f
C2072 VDD.n277 VSS 0.0202f
C2073 VDD.n278 VSS 0.0546f
C2074 VDD.n279 VSS 0.0131f
C2075 VDD.n280 VSS 0.0348f
C2076 VDD.n281 VSS 0.0359f
C2077 VDD.n282 VSS 0.0273f
C2078 VDD.n283 VSS 0.0277f
C2079 VDD.n284 VSS 0.0288f
C2080 VDD.n285 VSS 0.0333f
C2081 VDD.n286 VSS 0.0308f
C2082 VDD.n287 VSS 0.0267f
C2083 VDD.n288 VSS 0.037f
C2084 VDD.n289 VSS 0.0411f
C2085 VDD.n290 VSS 0.0274f
C2086 VDD.n291 VSS 0.0296f
C2087 VDD.n292 VSS 0.0297f
C2088 VDD.n293 VSS 0.0272f
C2089 VDD.n294 VSS 0.0411f
C2090 VDD.n295 VSS 0.0371f
C2091 VDD.n296 VSS 0.0265f
C2092 VDD.n297 VSS 0.0308f
C2093 VDD.n298 VSS 0.0334f
C2094 VDD.n299 VSS 0.0287f
C2095 VDD.n300 VSS 0.0277f
C2096 VDD.n301 VSS 0.0275f
C2097 VDD.n302 VSS 0.0358f
C2098 VDD.n303 VSS 0.0349f
C2099 VDD.n304 VSS 0.0133f
C2100 VDD.n305 VSS 0.0631f
C2101 VDD.t244 VSS 0.00584f
C2102 VDD.t57 VSS 0.0706f
C2103 VDD.n306 VSS 0.00585f
C2104 VDD.t153 VSS 0.0024f
C2105 VDD.n307 VSS 0.0024f
C2106 VDD.n308 VSS 0.00525f
C2107 VDD.n309 VSS 0.00585f
C2108 VDD.n310 VSS 0.0342f
C2109 VDD.t41 VSS 0.0704f
C2110 VDD.n311 VSS 0.00585f
C2111 VDD.t363 VSS 0.0038f
C2112 VDD.t40 VSS 0.00502f
C2113 VDD.n312 VSS 0.00985f
C2114 VDD.n313 VSS 0.00274f
C2115 VDD.t373 VSS 0.0038f
C2116 VDD.t20 VSS 0.00502f
C2117 VDD.n314 VSS 0.00983f
C2118 VDD.n315 VSS 0.00801f
C2119 VDD.n316 VSS 0.0436f
C2120 VDD.n317 VSS 0.0273f
C2121 VDD.t109 VSS 0.0024f
C2122 VDD.n318 VSS 0.0024f
C2123 VDD.n319 VSS 0.00525f
C2124 VDD.n320 VSS 0.0333f
C2125 VDD.n321 VSS 0.0181f
C2126 VDD.n322 VSS 0.0363f
C2127 VDD.t108 VSS 0.0398f
C2128 VDD.t229 VSS 0.086f
C2129 VDD.t67 VSS 0.0706f
C2130 VDD.t102 VSS 0.086f
C2131 VDD.t152 VSS 0.0398f
C2132 VDD.n323 VSS 0.0363f
C2133 VDD.n324 VSS 0.0181f
C2134 VDD.n325 VSS 0.0333f
C2135 VDD.n326 VSS 0.034f
C2136 VDD.t213 VSS 0.00584f
C2137 VDD.n327 VSS 0.00585f
C2138 VDD.n328 VSS 0.0269f
C2139 VDD.n329 VSS 0.029f
C2140 VDD.n330 VSS 0.0202f
C2141 VDD.n331 VSS 0.0363f
C2142 VDD.t212 VSS 0.077f
C2143 VDD.t217 VSS 0.0706f
C2144 VDD.t243 VSS 0.0759f
C2145 VDD.n332 VSS 0.0363f
C2146 VDD.n333 VSS 0.0202f
C2147 VDD.n334 VSS 0.0519f
C2148 VDD.n335 VSS 0.0602f
C2149 VDD.n336 VSS 0.0154f
C2150 VDD.n337 VSS 0.0365f
C2151 VDD.n338 VSS 0.0354f
C2152 VDD.n339 VSS 0.027f
C2153 VDD.n340 VSS 0.0273f
C2154 VDD.n341 VSS 0.0262f
C2155 VDD.n342 VSS 0.0328f
C2156 VDD.n343 VSS 0.0303f
C2157 VDD.n344 VSS 0.0286f
C2158 VDD.n345 VSS 0.0364f
C2159 VDD.n346 VSS 0.0404f
C2160 VDD.n347 VSS 0.027f
C2161 VDD.n348 VSS 0.0315f
C2162 VDD.n349 VSS 0.0316f
C2163 VDD.n350 VSS 0.0268f
C2164 VDD.n351 VSS 0.0404f
C2165 VDD.n352 VSS 0.0365f
C2166 VDD.n353 VSS 0.0285f
C2167 VDD.n354 VSS 0.0303f
C2168 VDD.n355 VSS 0.0329f
C2169 VDD.n356 VSS 0.0261f
C2170 VDD.n357 VSS 0.0273f
C2171 VDD.n358 VSS 0.0271f
C2172 VDD.n359 VSS 0.0352f
C2173 VDD.n360 VSS 0.0366f
C2174 VDD.n361 VSS 0.0155f
C2175 VDD.n362 VSS 0.0619f
C2176 VDD.n363 VSS 0.0563f
C2177 VDD.t174 VSS 0.0516f
C2178 VDD.t28 VSS 0.04f
C2179 VDD.n364 VSS 0.0543f
C2180 VDD.n365 VSS 0.0583f
C2181 VDD.n366 VSS 0.0264f
C2182 VDD.n367 VSS 0.0429f
C2183 VDD.n368 VSS 0.0383f
C2184 Q0.t9 VSS 0.045f
C2185 Q0.t14 VSS 0.0246f
C2186 Q0.n0 VSS 0.0855f
C2187 Q0.t8 VSS 0.0246f
C2188 Q0.t7 VSS 0.045f
C2189 Q0.n1 VSS 0.0855f
C2190 Q0.t5 VSS 0.0481f
C2191 Q0.t16 VSS 0.0317f
C2192 Q0.n2 VSS 0.0854f
C2193 Q0.n3 VSS 0.0288f
C2194 Q0.n4 VSS 0.00529f
C2195 Q0.t10 VSS 0.0396f
C2196 Q0.t15 VSS 0.0103f
C2197 Q0.n5 VSS 0.0657f
C2198 Q0.n6 VSS 0.00394f
C2199 Q0.n7 VSS 0.0157f
C2200 Q0.t3 VSS 0.0481f
C2201 Q0.t13 VSS 0.0317f
C2202 Q0.n8 VSS 0.0849f
C2203 Q0.n9 VSS 0.0111f
C2204 Q0.n10 VSS 0.00798f
C2205 Q0.n11 VSS 0.00398f
C2206 Q0.n12 VSS 0.159f
C2207 Q0.t12 VSS 0.0481f
C2208 Q0.t6 VSS 0.0317f
C2209 Q0.n13 VSS 0.0849f
C2210 Q0.n14 VSS 0.0111f
C2211 Q0.n15 VSS 0.00798f
C2212 Q0.n16 VSS 0.157f
C2213 Q0.n17 VSS 0.0971f
C2214 Q0.n18 VSS 0.106f
C2215 Q0.n19 VSS 0.014f
C2216 Q0.n20 VSS 0.00486f
C2217 Q0.n21 VSS 0.0286f
C2218 Q0.n22 VSS 0.0882f
C2219 Q0.t2 VSS 0.0262f
C2220 Q0.t0 VSS 0.0216f
C2221 Q0.n23 VSS 0.0216f
C2222 Q0.n24 VSS 0.0518f
C2223 Q0.n25 VSS 0.162f
C2224 Q0.n26 VSS 0.0193f
C2225 Q0.t11 VSS 0.0345f
C2226 Q0.t4 VSS 0.0276f
C2227 Q0.n27 VSS 0.0801f
C2228 Q0.n28 VSS 0.0497f
C2229 Q0.n29 VSS 0.51f
C2230 Q0.n30 VSS 0.74f
C2231 Q0.n31 VSS 0.489f
.ends

