magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2541 -2975 2541 2975
<< psubdiff >>
rect -541 953 541 975
rect -541 907 -519 953
rect -473 907 -395 953
rect -349 907 -271 953
rect -225 907 -147 953
rect -101 907 -23 953
rect 23 907 101 953
rect 147 907 225 953
rect 271 907 349 953
rect 395 907 473 953
rect 519 907 541 953
rect -541 829 541 907
rect -541 783 -519 829
rect -473 783 -395 829
rect -349 783 -271 829
rect -225 783 -147 829
rect -101 783 -23 829
rect 23 783 101 829
rect 147 783 225 829
rect 271 783 349 829
rect 395 783 473 829
rect 519 783 541 829
rect -541 705 541 783
rect -541 659 -519 705
rect -473 659 -395 705
rect -349 659 -271 705
rect -225 659 -147 705
rect -101 659 -23 705
rect 23 659 101 705
rect 147 659 225 705
rect 271 659 349 705
rect 395 659 473 705
rect 519 659 541 705
rect -541 581 541 659
rect -541 535 -519 581
rect -473 535 -395 581
rect -349 535 -271 581
rect -225 535 -147 581
rect -101 535 -23 581
rect 23 535 101 581
rect 147 535 225 581
rect 271 535 349 581
rect 395 535 473 581
rect 519 535 541 581
rect -541 457 541 535
rect -541 411 -519 457
rect -473 411 -395 457
rect -349 411 -271 457
rect -225 411 -147 457
rect -101 411 -23 457
rect 23 411 101 457
rect 147 411 225 457
rect 271 411 349 457
rect 395 411 473 457
rect 519 411 541 457
rect -541 333 541 411
rect -541 287 -519 333
rect -473 287 -395 333
rect -349 287 -271 333
rect -225 287 -147 333
rect -101 287 -23 333
rect 23 287 101 333
rect 147 287 225 333
rect 271 287 349 333
rect 395 287 473 333
rect 519 287 541 333
rect -541 209 541 287
rect -541 163 -519 209
rect -473 163 -395 209
rect -349 163 -271 209
rect -225 163 -147 209
rect -101 163 -23 209
rect 23 163 101 209
rect 147 163 225 209
rect 271 163 349 209
rect 395 163 473 209
rect 519 163 541 209
rect -541 85 541 163
rect -541 39 -519 85
rect -473 39 -395 85
rect -349 39 -271 85
rect -225 39 -147 85
rect -101 39 -23 85
rect 23 39 101 85
rect 147 39 225 85
rect 271 39 349 85
rect 395 39 473 85
rect 519 39 541 85
rect -541 -39 541 39
rect -541 -85 -519 -39
rect -473 -85 -395 -39
rect -349 -85 -271 -39
rect -225 -85 -147 -39
rect -101 -85 -23 -39
rect 23 -85 101 -39
rect 147 -85 225 -39
rect 271 -85 349 -39
rect 395 -85 473 -39
rect 519 -85 541 -39
rect -541 -163 541 -85
rect -541 -209 -519 -163
rect -473 -209 -395 -163
rect -349 -209 -271 -163
rect -225 -209 -147 -163
rect -101 -209 -23 -163
rect 23 -209 101 -163
rect 147 -209 225 -163
rect 271 -209 349 -163
rect 395 -209 473 -163
rect 519 -209 541 -163
rect -541 -287 541 -209
rect -541 -333 -519 -287
rect -473 -333 -395 -287
rect -349 -333 -271 -287
rect -225 -333 -147 -287
rect -101 -333 -23 -287
rect 23 -333 101 -287
rect 147 -333 225 -287
rect 271 -333 349 -287
rect 395 -333 473 -287
rect 519 -333 541 -287
rect -541 -411 541 -333
rect -541 -457 -519 -411
rect -473 -457 -395 -411
rect -349 -457 -271 -411
rect -225 -457 -147 -411
rect -101 -457 -23 -411
rect 23 -457 101 -411
rect 147 -457 225 -411
rect 271 -457 349 -411
rect 395 -457 473 -411
rect 519 -457 541 -411
rect -541 -535 541 -457
rect -541 -581 -519 -535
rect -473 -581 -395 -535
rect -349 -581 -271 -535
rect -225 -581 -147 -535
rect -101 -581 -23 -535
rect 23 -581 101 -535
rect 147 -581 225 -535
rect 271 -581 349 -535
rect 395 -581 473 -535
rect 519 -581 541 -535
rect -541 -659 541 -581
rect -541 -705 -519 -659
rect -473 -705 -395 -659
rect -349 -705 -271 -659
rect -225 -705 -147 -659
rect -101 -705 -23 -659
rect 23 -705 101 -659
rect 147 -705 225 -659
rect 271 -705 349 -659
rect 395 -705 473 -659
rect 519 -705 541 -659
rect -541 -783 541 -705
rect -541 -829 -519 -783
rect -473 -829 -395 -783
rect -349 -829 -271 -783
rect -225 -829 -147 -783
rect -101 -829 -23 -783
rect 23 -829 101 -783
rect 147 -829 225 -783
rect 271 -829 349 -783
rect 395 -829 473 -783
rect 519 -829 541 -783
rect -541 -907 541 -829
rect -541 -953 -519 -907
rect -473 -953 -395 -907
rect -349 -953 -271 -907
rect -225 -953 -147 -907
rect -101 -953 -23 -907
rect 23 -953 101 -907
rect 147 -953 225 -907
rect 271 -953 349 -907
rect 395 -953 473 -907
rect 519 -953 541 -907
rect -541 -975 541 -953
<< psubdiffcont >>
rect -519 907 -473 953
rect -395 907 -349 953
rect -271 907 -225 953
rect -147 907 -101 953
rect -23 907 23 953
rect 101 907 147 953
rect 225 907 271 953
rect 349 907 395 953
rect 473 907 519 953
rect -519 783 -473 829
rect -395 783 -349 829
rect -271 783 -225 829
rect -147 783 -101 829
rect -23 783 23 829
rect 101 783 147 829
rect 225 783 271 829
rect 349 783 395 829
rect 473 783 519 829
rect -519 659 -473 705
rect -395 659 -349 705
rect -271 659 -225 705
rect -147 659 -101 705
rect -23 659 23 705
rect 101 659 147 705
rect 225 659 271 705
rect 349 659 395 705
rect 473 659 519 705
rect -519 535 -473 581
rect -395 535 -349 581
rect -271 535 -225 581
rect -147 535 -101 581
rect -23 535 23 581
rect 101 535 147 581
rect 225 535 271 581
rect 349 535 395 581
rect 473 535 519 581
rect -519 411 -473 457
rect -395 411 -349 457
rect -271 411 -225 457
rect -147 411 -101 457
rect -23 411 23 457
rect 101 411 147 457
rect 225 411 271 457
rect 349 411 395 457
rect 473 411 519 457
rect -519 287 -473 333
rect -395 287 -349 333
rect -271 287 -225 333
rect -147 287 -101 333
rect -23 287 23 333
rect 101 287 147 333
rect 225 287 271 333
rect 349 287 395 333
rect 473 287 519 333
rect -519 163 -473 209
rect -395 163 -349 209
rect -271 163 -225 209
rect -147 163 -101 209
rect -23 163 23 209
rect 101 163 147 209
rect 225 163 271 209
rect 349 163 395 209
rect 473 163 519 209
rect -519 39 -473 85
rect -395 39 -349 85
rect -271 39 -225 85
rect -147 39 -101 85
rect -23 39 23 85
rect 101 39 147 85
rect 225 39 271 85
rect 349 39 395 85
rect 473 39 519 85
rect -519 -85 -473 -39
rect -395 -85 -349 -39
rect -271 -85 -225 -39
rect -147 -85 -101 -39
rect -23 -85 23 -39
rect 101 -85 147 -39
rect 225 -85 271 -39
rect 349 -85 395 -39
rect 473 -85 519 -39
rect -519 -209 -473 -163
rect -395 -209 -349 -163
rect -271 -209 -225 -163
rect -147 -209 -101 -163
rect -23 -209 23 -163
rect 101 -209 147 -163
rect 225 -209 271 -163
rect 349 -209 395 -163
rect 473 -209 519 -163
rect -519 -333 -473 -287
rect -395 -333 -349 -287
rect -271 -333 -225 -287
rect -147 -333 -101 -287
rect -23 -333 23 -287
rect 101 -333 147 -287
rect 225 -333 271 -287
rect 349 -333 395 -287
rect 473 -333 519 -287
rect -519 -457 -473 -411
rect -395 -457 -349 -411
rect -271 -457 -225 -411
rect -147 -457 -101 -411
rect -23 -457 23 -411
rect 101 -457 147 -411
rect 225 -457 271 -411
rect 349 -457 395 -411
rect 473 -457 519 -411
rect -519 -581 -473 -535
rect -395 -581 -349 -535
rect -271 -581 -225 -535
rect -147 -581 -101 -535
rect -23 -581 23 -535
rect 101 -581 147 -535
rect 225 -581 271 -535
rect 349 -581 395 -535
rect 473 -581 519 -535
rect -519 -705 -473 -659
rect -395 -705 -349 -659
rect -271 -705 -225 -659
rect -147 -705 -101 -659
rect -23 -705 23 -659
rect 101 -705 147 -659
rect 225 -705 271 -659
rect 349 -705 395 -659
rect 473 -705 519 -659
rect -519 -829 -473 -783
rect -395 -829 -349 -783
rect -271 -829 -225 -783
rect -147 -829 -101 -783
rect -23 -829 23 -783
rect 101 -829 147 -783
rect 225 -829 271 -783
rect 349 -829 395 -783
rect 473 -829 519 -783
rect -519 -953 -473 -907
rect -395 -953 -349 -907
rect -271 -953 -225 -907
rect -147 -953 -101 -907
rect -23 -953 23 -907
rect 101 -953 147 -907
rect 225 -953 271 -907
rect 349 -953 395 -907
rect 473 -953 519 -907
<< metal1 >>
rect -530 953 530 964
rect -530 907 -519 953
rect -473 907 -395 953
rect -349 907 -271 953
rect -225 907 -147 953
rect -101 907 -23 953
rect 23 907 101 953
rect 147 907 225 953
rect 271 907 349 953
rect 395 907 473 953
rect 519 907 530 953
rect -530 829 530 907
rect -530 783 -519 829
rect -473 783 -395 829
rect -349 783 -271 829
rect -225 783 -147 829
rect -101 783 -23 829
rect 23 783 101 829
rect 147 783 225 829
rect 271 783 349 829
rect 395 783 473 829
rect 519 783 530 829
rect -530 705 530 783
rect -530 659 -519 705
rect -473 659 -395 705
rect -349 659 -271 705
rect -225 659 -147 705
rect -101 659 -23 705
rect 23 659 101 705
rect 147 659 225 705
rect 271 659 349 705
rect 395 659 473 705
rect 519 659 530 705
rect -530 581 530 659
rect -530 535 -519 581
rect -473 535 -395 581
rect -349 535 -271 581
rect -225 535 -147 581
rect -101 535 -23 581
rect 23 535 101 581
rect 147 535 225 581
rect 271 535 349 581
rect 395 535 473 581
rect 519 535 530 581
rect -530 457 530 535
rect -530 411 -519 457
rect -473 411 -395 457
rect -349 411 -271 457
rect -225 411 -147 457
rect -101 411 -23 457
rect 23 411 101 457
rect 147 411 225 457
rect 271 411 349 457
rect 395 411 473 457
rect 519 411 530 457
rect -530 333 530 411
rect -530 287 -519 333
rect -473 287 -395 333
rect -349 287 -271 333
rect -225 287 -147 333
rect -101 287 -23 333
rect 23 287 101 333
rect 147 287 225 333
rect 271 287 349 333
rect 395 287 473 333
rect 519 287 530 333
rect -530 209 530 287
rect -530 163 -519 209
rect -473 163 -395 209
rect -349 163 -271 209
rect -225 163 -147 209
rect -101 163 -23 209
rect 23 163 101 209
rect 147 163 225 209
rect 271 163 349 209
rect 395 163 473 209
rect 519 163 530 209
rect -530 85 530 163
rect -530 39 -519 85
rect -473 39 -395 85
rect -349 39 -271 85
rect -225 39 -147 85
rect -101 39 -23 85
rect 23 39 101 85
rect 147 39 225 85
rect 271 39 349 85
rect 395 39 473 85
rect 519 39 530 85
rect -530 -39 530 39
rect -530 -85 -519 -39
rect -473 -85 -395 -39
rect -349 -85 -271 -39
rect -225 -85 -147 -39
rect -101 -85 -23 -39
rect 23 -85 101 -39
rect 147 -85 225 -39
rect 271 -85 349 -39
rect 395 -85 473 -39
rect 519 -85 530 -39
rect -530 -163 530 -85
rect -530 -209 -519 -163
rect -473 -209 -395 -163
rect -349 -209 -271 -163
rect -225 -209 -147 -163
rect -101 -209 -23 -163
rect 23 -209 101 -163
rect 147 -209 225 -163
rect 271 -209 349 -163
rect 395 -209 473 -163
rect 519 -209 530 -163
rect -530 -287 530 -209
rect -530 -333 -519 -287
rect -473 -333 -395 -287
rect -349 -333 -271 -287
rect -225 -333 -147 -287
rect -101 -333 -23 -287
rect 23 -333 101 -287
rect 147 -333 225 -287
rect 271 -333 349 -287
rect 395 -333 473 -287
rect 519 -333 530 -287
rect -530 -411 530 -333
rect -530 -457 -519 -411
rect -473 -457 -395 -411
rect -349 -457 -271 -411
rect -225 -457 -147 -411
rect -101 -457 -23 -411
rect 23 -457 101 -411
rect 147 -457 225 -411
rect 271 -457 349 -411
rect 395 -457 473 -411
rect 519 -457 530 -411
rect -530 -535 530 -457
rect -530 -581 -519 -535
rect -473 -581 -395 -535
rect -349 -581 -271 -535
rect -225 -581 -147 -535
rect -101 -581 -23 -535
rect 23 -581 101 -535
rect 147 -581 225 -535
rect 271 -581 349 -535
rect 395 -581 473 -535
rect 519 -581 530 -535
rect -530 -659 530 -581
rect -530 -705 -519 -659
rect -473 -705 -395 -659
rect -349 -705 -271 -659
rect -225 -705 -147 -659
rect -101 -705 -23 -659
rect 23 -705 101 -659
rect 147 -705 225 -659
rect 271 -705 349 -659
rect 395 -705 473 -659
rect 519 -705 530 -659
rect -530 -783 530 -705
rect -530 -829 -519 -783
rect -473 -829 -395 -783
rect -349 -829 -271 -783
rect -225 -829 -147 -783
rect -101 -829 -23 -783
rect 23 -829 101 -783
rect 147 -829 225 -783
rect 271 -829 349 -783
rect 395 -829 473 -783
rect 519 -829 530 -783
rect -530 -907 530 -829
rect -530 -953 -519 -907
rect -473 -953 -395 -907
rect -349 -953 -271 -907
rect -225 -953 -147 -907
rect -101 -953 -23 -907
rect 23 -953 101 -907
rect 147 -953 225 -907
rect 271 -953 349 -907
rect 395 -953 473 -907
rect 519 -953 530 -907
rect -530 -964 530 -953
<< end >>
