magic
tech gf180mcuC
magscale 1 10
timestamp 1692680230
<< nwell >>
rect -762 -330 762 330
<< pmos >>
rect -588 -200 -532 200
rect -428 -200 -372 200
rect -268 -200 -212 200
rect -108 -200 -52 200
rect 52 -200 108 200
rect 212 -200 268 200
rect 372 -200 428 200
rect 532 -200 588 200
<< pdiff >>
rect -676 187 -588 200
rect -676 -187 -663 187
rect -617 -187 -588 187
rect -676 -200 -588 -187
rect -532 187 -428 200
rect -532 -187 -503 187
rect -457 -187 -428 187
rect -532 -200 -428 -187
rect -372 187 -268 200
rect -372 -187 -343 187
rect -297 -187 -268 187
rect -372 -200 -268 -187
rect -212 187 -108 200
rect -212 -187 -183 187
rect -137 -187 -108 187
rect -212 -200 -108 -187
rect -52 187 52 200
rect -52 -187 -23 187
rect 23 -187 52 187
rect -52 -200 52 -187
rect 108 187 212 200
rect 108 -187 137 187
rect 183 -187 212 187
rect 108 -200 212 -187
rect 268 187 372 200
rect 268 -187 297 187
rect 343 -187 372 187
rect 268 -200 372 -187
rect 428 187 532 200
rect 428 -187 457 187
rect 503 -187 532 187
rect 428 -200 532 -187
rect 588 187 676 200
rect 588 -187 617 187
rect 663 -187 676 187
rect 588 -200 676 -187
<< pdiffc >>
rect -663 -187 -617 187
rect -503 -187 -457 187
rect -343 -187 -297 187
rect -183 -187 -137 187
rect -23 -187 23 187
rect 137 -187 183 187
rect 297 -187 343 187
rect 457 -187 503 187
rect 617 -187 663 187
<< polysilicon >>
rect -588 200 -532 244
rect -428 200 -372 244
rect -268 200 -212 244
rect -108 200 -52 244
rect 52 200 108 244
rect 212 200 268 244
rect 372 200 428 244
rect 532 200 588 244
rect -588 -244 -532 -200
rect -428 -244 -372 -200
rect -268 -244 -212 -200
rect -108 -244 -52 -200
rect 52 -244 108 -200
rect 212 -244 268 -200
rect 372 -244 428 -200
rect 532 -244 588 -200
<< metal1 >>
rect -663 187 -617 198
rect -663 -198 -617 -187
rect -503 187 -457 198
rect -503 -198 -457 -187
rect -343 187 -297 198
rect -343 -198 -297 -187
rect -183 187 -137 198
rect -183 -198 -137 -187
rect -23 187 23 198
rect -23 -198 23 -187
rect 137 187 183 198
rect 137 -198 183 -187
rect 297 187 343 198
rect 297 -198 343 -187
rect 457 187 503 198
rect 457 -198 503 -187
rect 617 187 663 198
rect 617 -198 663 -187
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2 l 0.280 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
