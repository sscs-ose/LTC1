magic
tech gf180mcuC
magscale 1 10
timestamp 1714558796
<< nwell >>
rect 4392 3239 4912 3247
rect 4392 3191 4924 3239
rect 4404 3183 4924 3191
rect 4821 3164 4846 3183
rect 4763 3092 4869 3164
rect 4821 2824 4838 3092
rect 4821 2719 4870 2824
rect 4829 2558 4870 2719
rect 2818 1620 3058 2089
rect 1555 561 1567 599
<< pwell >>
rect 4356 2497 4479 2608
rect 4677 2502 4707 2507
rect 4746 2502 4790 2691
rect 4670 2498 4895 2502
rect 4670 2355 4907 2498
rect 5341 2336 5454 2502
<< psubdiff >>
rect 5387 2234 5478 2298
<< metal1 >>
rect 3639 3093 3867 3249
rect 4824 3164 4846 3188
rect 5476 3185 5528 3211
rect 2945 1983 3047 2089
rect 3639 2039 3795 3093
rect 4763 3092 4869 3164
rect 4820 2581 4875 2746
rect 5143 2624 5225 2644
rect 4820 2566 4905 2581
rect 5143 2572 5156 2624
rect 5208 2572 5225 2624
rect 5143 2568 5225 2572
rect 4820 2535 4995 2566
rect 4859 2520 4995 2535
rect 5714 2527 5798 2585
rect 4516 2317 4836 2319
rect 4516 2271 4843 2317
rect 4517 2201 4843 2271
rect 5361 2200 6160 2305
rect 85 1603 119 1643
rect 2806 1544 2834 1591
rect 5840 1549 5851 1582
rect 491 505 549 725
rect 1555 561 1567 599
rect 491 468 542 505
rect 2377 438 2433 494
rect 6057 109 6160 2200
rect 2856 0 3295 109
rect 5873 0 6160 109
rect 6050 -1 6160 0
<< via1 >>
rect 4257 2745 4309 2797
rect 3999 2639 4051 2691
rect 5156 2572 5208 2624
rect 546 1544 598 1596
rect 3563 1544 3615 1596
rect 1485 552 1537 604
rect 4502 549 4554 601
rect 542 453 594 505
rect 3563 454 3615 506
<< metal2 >>
rect 4255 2797 4311 2809
rect 4255 2745 4257 2797
rect 4309 2745 4311 2797
rect 3997 2691 4053 2703
rect 3997 2639 3999 2691
rect 4051 2639 4053 2691
rect 3773 2306 3829 2319
rect 3997 2306 4053 2639
rect 3829 2250 4053 2306
rect 3773 2249 4053 2250
rect 3773 2238 3829 2249
rect 4255 2181 4311 2745
rect 5143 2624 5225 2644
rect 5143 2572 5156 2624
rect 5208 2572 5225 2624
rect 5143 2568 5225 2572
rect 3560 2179 4311 2181
rect 3560 2123 3572 2179
rect 3628 2123 4311 2179
rect 3560 2122 4311 2123
rect 5154 2177 5210 2568
rect 5154 2121 5835 2177
rect 21 2009 5684 2065
rect 21 1529 77 2009
rect 133 1890 3207 1947
rect 133 1587 190 1890
rect 544 1596 601 1608
rect 544 1544 546 1596
rect 598 1544 601 1596
rect 3150 1587 3207 1890
rect 3560 1596 3619 1608
rect 544 1529 601 1544
rect 3560 1544 3563 1596
rect 3615 1544 3619 1596
rect 5628 1580 5684 2009
rect 3560 1541 3619 1544
rect 3560 1531 3561 1541
rect 21 1473 601 1529
rect 2744 1485 3561 1531
rect 3617 1485 3619 1541
rect 2744 1475 3619 1485
rect 5779 1480 5835 2121
rect 1474 604 1549 616
rect 1474 552 1485 604
rect 1537 552 1549 604
rect 540 505 596 517
rect 540 453 542 505
rect 594 453 596 505
rect 540 153 596 453
rect 1474 494 1549 552
rect 4499 601 4556 613
rect 4499 549 4502 601
rect 4554 549 4556 601
rect 3561 506 3617 518
rect 1474 438 2427 494
rect 2483 438 2553 494
rect 1474 437 2553 438
rect 3561 454 3563 506
rect 3615 454 3617 506
rect 4499 494 4556 549
rect 3561 153 3617 454
rect 4183 493 4556 494
rect 4183 437 4193 493
rect 4249 437 4556 493
rect 540 97 3617 153
<< via2 >>
rect 3773 2250 3829 2306
rect 3572 2123 3628 2179
rect 3773 1570 3829 1626
rect 3561 1485 3617 1541
rect 2427 438 2483 494
rect 4193 437 4249 493
<< metal3 >>
rect 3773 2306 3829 2319
rect 3560 2179 3638 2181
rect 3560 2123 3572 2179
rect 3628 2123 3638 2179
rect 3560 2122 3638 2123
rect 3560 1541 3619 2122
rect 3773 1626 3829 2250
rect 3773 1560 3829 1570
rect 3560 1485 3561 1541
rect 3617 1485 3619 1541
rect 3560 1475 3619 1485
rect 2405 438 2427 494
rect 2483 493 4259 494
rect 2483 438 4193 493
rect 2405 437 4193 438
rect 4249 437 4259 493
use and2_mag  and2_mag_0
timestamp 1714558667
transform 1 0 3919 0 1 2384
box -70 -188 1009 863
use JK_FF_mag  JK_FF_mag_0
timestamp 1714558667
transform 1 0 3407 0 1 0
box -430 0 2603 2148
use JK_FF_mag  JK_FF_mag_1
timestamp 1714558667
transform 1 0 390 0 1 0
box -430 0 2603 2148
use or_2  or_2_0
timestamp 1714126980
transform 1 0 6460 0 1 1250
box 0 0 1 1
use or_2_mag  or_2_mag_0
timestamp 1714558667
transform 1 0 4500 0 1 1690
box 330 510 1401 1521
<< labels >>
flabel metal1 3687 2882 3687 2882 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal1 3089 47 3089 47 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal1 2819 1564 2819 1564 0 FreeSans 320 0 0 0 Q1
port 4 nsew
flabel metal1 5845 1571 5845 1571 0 FreeSans 320 0 0 0 Q0
port 5 nsew
flabel metal1 5763 2560 5763 2560 0 FreeSans 800 0 0 0 Vdiv3
port 6 nsew
flabel metal1 101 1623 101 1623 0 FreeSans 800 0 0 0 CLK
port 7 nsew
flabel via1 1504 577 1504 577 0 FreeSans 800 0 0 0 RST
port 8 nsew
<< end >>
