magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -3398 -1319 3398 1319
<< metal4 >>
rect -2395 311 2395 316
rect -2395 283 -2390 311
rect -2362 283 -2324 311
rect -2296 283 -2258 311
rect -2230 283 -2192 311
rect -2164 283 -2126 311
rect -2098 283 -2060 311
rect -2032 283 -1994 311
rect -1966 283 -1928 311
rect -1900 283 -1862 311
rect -1834 283 -1796 311
rect -1768 283 -1730 311
rect -1702 283 -1664 311
rect -1636 283 -1598 311
rect -1570 283 -1532 311
rect -1504 283 -1466 311
rect -1438 283 -1400 311
rect -1372 283 -1334 311
rect -1306 283 -1268 311
rect -1240 283 -1202 311
rect -1174 283 -1136 311
rect -1108 283 -1070 311
rect -1042 283 -1004 311
rect -976 283 -938 311
rect -910 283 -872 311
rect -844 283 -806 311
rect -778 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 778 311
rect 806 283 844 311
rect 872 283 910 311
rect 938 283 976 311
rect 1004 283 1042 311
rect 1070 283 1108 311
rect 1136 283 1174 311
rect 1202 283 1240 311
rect 1268 283 1306 311
rect 1334 283 1372 311
rect 1400 283 1438 311
rect 1466 283 1504 311
rect 1532 283 1570 311
rect 1598 283 1636 311
rect 1664 283 1702 311
rect 1730 283 1768 311
rect 1796 283 1834 311
rect 1862 283 1900 311
rect 1928 283 1966 311
rect 1994 283 2032 311
rect 2060 283 2098 311
rect 2126 283 2164 311
rect 2192 283 2230 311
rect 2258 283 2296 311
rect 2324 283 2362 311
rect 2390 283 2395 311
rect -2395 245 2395 283
rect -2395 217 -2390 245
rect -2362 217 -2324 245
rect -2296 217 -2258 245
rect -2230 217 -2192 245
rect -2164 217 -2126 245
rect -2098 217 -2060 245
rect -2032 217 -1994 245
rect -1966 217 -1928 245
rect -1900 217 -1862 245
rect -1834 217 -1796 245
rect -1768 217 -1730 245
rect -1702 217 -1664 245
rect -1636 217 -1598 245
rect -1570 217 -1532 245
rect -1504 217 -1466 245
rect -1438 217 -1400 245
rect -1372 217 -1334 245
rect -1306 217 -1268 245
rect -1240 217 -1202 245
rect -1174 217 -1136 245
rect -1108 217 -1070 245
rect -1042 217 -1004 245
rect -976 217 -938 245
rect -910 217 -872 245
rect -844 217 -806 245
rect -778 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 778 245
rect 806 217 844 245
rect 872 217 910 245
rect 938 217 976 245
rect 1004 217 1042 245
rect 1070 217 1108 245
rect 1136 217 1174 245
rect 1202 217 1240 245
rect 1268 217 1306 245
rect 1334 217 1372 245
rect 1400 217 1438 245
rect 1466 217 1504 245
rect 1532 217 1570 245
rect 1598 217 1636 245
rect 1664 217 1702 245
rect 1730 217 1768 245
rect 1796 217 1834 245
rect 1862 217 1900 245
rect 1928 217 1966 245
rect 1994 217 2032 245
rect 2060 217 2098 245
rect 2126 217 2164 245
rect 2192 217 2230 245
rect 2258 217 2296 245
rect 2324 217 2362 245
rect 2390 217 2395 245
rect -2395 179 2395 217
rect -2395 151 -2390 179
rect -2362 151 -2324 179
rect -2296 151 -2258 179
rect -2230 151 -2192 179
rect -2164 151 -2126 179
rect -2098 151 -2060 179
rect -2032 151 -1994 179
rect -1966 151 -1928 179
rect -1900 151 -1862 179
rect -1834 151 -1796 179
rect -1768 151 -1730 179
rect -1702 151 -1664 179
rect -1636 151 -1598 179
rect -1570 151 -1532 179
rect -1504 151 -1466 179
rect -1438 151 -1400 179
rect -1372 151 -1334 179
rect -1306 151 -1268 179
rect -1240 151 -1202 179
rect -1174 151 -1136 179
rect -1108 151 -1070 179
rect -1042 151 -1004 179
rect -976 151 -938 179
rect -910 151 -872 179
rect -844 151 -806 179
rect -778 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 778 179
rect 806 151 844 179
rect 872 151 910 179
rect 938 151 976 179
rect 1004 151 1042 179
rect 1070 151 1108 179
rect 1136 151 1174 179
rect 1202 151 1240 179
rect 1268 151 1306 179
rect 1334 151 1372 179
rect 1400 151 1438 179
rect 1466 151 1504 179
rect 1532 151 1570 179
rect 1598 151 1636 179
rect 1664 151 1702 179
rect 1730 151 1768 179
rect 1796 151 1834 179
rect 1862 151 1900 179
rect 1928 151 1966 179
rect 1994 151 2032 179
rect 2060 151 2098 179
rect 2126 151 2164 179
rect 2192 151 2230 179
rect 2258 151 2296 179
rect 2324 151 2362 179
rect 2390 151 2395 179
rect -2395 113 2395 151
rect -2395 85 -2390 113
rect -2362 85 -2324 113
rect -2296 85 -2258 113
rect -2230 85 -2192 113
rect -2164 85 -2126 113
rect -2098 85 -2060 113
rect -2032 85 -1994 113
rect -1966 85 -1928 113
rect -1900 85 -1862 113
rect -1834 85 -1796 113
rect -1768 85 -1730 113
rect -1702 85 -1664 113
rect -1636 85 -1598 113
rect -1570 85 -1532 113
rect -1504 85 -1466 113
rect -1438 85 -1400 113
rect -1372 85 -1334 113
rect -1306 85 -1268 113
rect -1240 85 -1202 113
rect -1174 85 -1136 113
rect -1108 85 -1070 113
rect -1042 85 -1004 113
rect -976 85 -938 113
rect -910 85 -872 113
rect -844 85 -806 113
rect -778 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 778 113
rect 806 85 844 113
rect 872 85 910 113
rect 938 85 976 113
rect 1004 85 1042 113
rect 1070 85 1108 113
rect 1136 85 1174 113
rect 1202 85 1240 113
rect 1268 85 1306 113
rect 1334 85 1372 113
rect 1400 85 1438 113
rect 1466 85 1504 113
rect 1532 85 1570 113
rect 1598 85 1636 113
rect 1664 85 1702 113
rect 1730 85 1768 113
rect 1796 85 1834 113
rect 1862 85 1900 113
rect 1928 85 1966 113
rect 1994 85 2032 113
rect 2060 85 2098 113
rect 2126 85 2164 113
rect 2192 85 2230 113
rect 2258 85 2296 113
rect 2324 85 2362 113
rect 2390 85 2395 113
rect -2395 47 2395 85
rect -2395 19 -2390 47
rect -2362 19 -2324 47
rect -2296 19 -2258 47
rect -2230 19 -2192 47
rect -2164 19 -2126 47
rect -2098 19 -2060 47
rect -2032 19 -1994 47
rect -1966 19 -1928 47
rect -1900 19 -1862 47
rect -1834 19 -1796 47
rect -1768 19 -1730 47
rect -1702 19 -1664 47
rect -1636 19 -1598 47
rect -1570 19 -1532 47
rect -1504 19 -1466 47
rect -1438 19 -1400 47
rect -1372 19 -1334 47
rect -1306 19 -1268 47
rect -1240 19 -1202 47
rect -1174 19 -1136 47
rect -1108 19 -1070 47
rect -1042 19 -1004 47
rect -976 19 -938 47
rect -910 19 -872 47
rect -844 19 -806 47
rect -778 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 778 47
rect 806 19 844 47
rect 872 19 910 47
rect 938 19 976 47
rect 1004 19 1042 47
rect 1070 19 1108 47
rect 1136 19 1174 47
rect 1202 19 1240 47
rect 1268 19 1306 47
rect 1334 19 1372 47
rect 1400 19 1438 47
rect 1466 19 1504 47
rect 1532 19 1570 47
rect 1598 19 1636 47
rect 1664 19 1702 47
rect 1730 19 1768 47
rect 1796 19 1834 47
rect 1862 19 1900 47
rect 1928 19 1966 47
rect 1994 19 2032 47
rect 2060 19 2098 47
rect 2126 19 2164 47
rect 2192 19 2230 47
rect 2258 19 2296 47
rect 2324 19 2362 47
rect 2390 19 2395 47
rect -2395 -19 2395 19
rect -2395 -47 -2390 -19
rect -2362 -47 -2324 -19
rect -2296 -47 -2258 -19
rect -2230 -47 -2192 -19
rect -2164 -47 -2126 -19
rect -2098 -47 -2060 -19
rect -2032 -47 -1994 -19
rect -1966 -47 -1928 -19
rect -1900 -47 -1862 -19
rect -1834 -47 -1796 -19
rect -1768 -47 -1730 -19
rect -1702 -47 -1664 -19
rect -1636 -47 -1598 -19
rect -1570 -47 -1532 -19
rect -1504 -47 -1466 -19
rect -1438 -47 -1400 -19
rect -1372 -47 -1334 -19
rect -1306 -47 -1268 -19
rect -1240 -47 -1202 -19
rect -1174 -47 -1136 -19
rect -1108 -47 -1070 -19
rect -1042 -47 -1004 -19
rect -976 -47 -938 -19
rect -910 -47 -872 -19
rect -844 -47 -806 -19
rect -778 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 778 -19
rect 806 -47 844 -19
rect 872 -47 910 -19
rect 938 -47 976 -19
rect 1004 -47 1042 -19
rect 1070 -47 1108 -19
rect 1136 -47 1174 -19
rect 1202 -47 1240 -19
rect 1268 -47 1306 -19
rect 1334 -47 1372 -19
rect 1400 -47 1438 -19
rect 1466 -47 1504 -19
rect 1532 -47 1570 -19
rect 1598 -47 1636 -19
rect 1664 -47 1702 -19
rect 1730 -47 1768 -19
rect 1796 -47 1834 -19
rect 1862 -47 1900 -19
rect 1928 -47 1966 -19
rect 1994 -47 2032 -19
rect 2060 -47 2098 -19
rect 2126 -47 2164 -19
rect 2192 -47 2230 -19
rect 2258 -47 2296 -19
rect 2324 -47 2362 -19
rect 2390 -47 2395 -19
rect -2395 -85 2395 -47
rect -2395 -113 -2390 -85
rect -2362 -113 -2324 -85
rect -2296 -113 -2258 -85
rect -2230 -113 -2192 -85
rect -2164 -113 -2126 -85
rect -2098 -113 -2060 -85
rect -2032 -113 -1994 -85
rect -1966 -113 -1928 -85
rect -1900 -113 -1862 -85
rect -1834 -113 -1796 -85
rect -1768 -113 -1730 -85
rect -1702 -113 -1664 -85
rect -1636 -113 -1598 -85
rect -1570 -113 -1532 -85
rect -1504 -113 -1466 -85
rect -1438 -113 -1400 -85
rect -1372 -113 -1334 -85
rect -1306 -113 -1268 -85
rect -1240 -113 -1202 -85
rect -1174 -113 -1136 -85
rect -1108 -113 -1070 -85
rect -1042 -113 -1004 -85
rect -976 -113 -938 -85
rect -910 -113 -872 -85
rect -844 -113 -806 -85
rect -778 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 778 -85
rect 806 -113 844 -85
rect 872 -113 910 -85
rect 938 -113 976 -85
rect 1004 -113 1042 -85
rect 1070 -113 1108 -85
rect 1136 -113 1174 -85
rect 1202 -113 1240 -85
rect 1268 -113 1306 -85
rect 1334 -113 1372 -85
rect 1400 -113 1438 -85
rect 1466 -113 1504 -85
rect 1532 -113 1570 -85
rect 1598 -113 1636 -85
rect 1664 -113 1702 -85
rect 1730 -113 1768 -85
rect 1796 -113 1834 -85
rect 1862 -113 1900 -85
rect 1928 -113 1966 -85
rect 1994 -113 2032 -85
rect 2060 -113 2098 -85
rect 2126 -113 2164 -85
rect 2192 -113 2230 -85
rect 2258 -113 2296 -85
rect 2324 -113 2362 -85
rect 2390 -113 2395 -85
rect -2395 -151 2395 -113
rect -2395 -179 -2390 -151
rect -2362 -179 -2324 -151
rect -2296 -179 -2258 -151
rect -2230 -179 -2192 -151
rect -2164 -179 -2126 -151
rect -2098 -179 -2060 -151
rect -2032 -179 -1994 -151
rect -1966 -179 -1928 -151
rect -1900 -179 -1862 -151
rect -1834 -179 -1796 -151
rect -1768 -179 -1730 -151
rect -1702 -179 -1664 -151
rect -1636 -179 -1598 -151
rect -1570 -179 -1532 -151
rect -1504 -179 -1466 -151
rect -1438 -179 -1400 -151
rect -1372 -179 -1334 -151
rect -1306 -179 -1268 -151
rect -1240 -179 -1202 -151
rect -1174 -179 -1136 -151
rect -1108 -179 -1070 -151
rect -1042 -179 -1004 -151
rect -976 -179 -938 -151
rect -910 -179 -872 -151
rect -844 -179 -806 -151
rect -778 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 778 -151
rect 806 -179 844 -151
rect 872 -179 910 -151
rect 938 -179 976 -151
rect 1004 -179 1042 -151
rect 1070 -179 1108 -151
rect 1136 -179 1174 -151
rect 1202 -179 1240 -151
rect 1268 -179 1306 -151
rect 1334 -179 1372 -151
rect 1400 -179 1438 -151
rect 1466 -179 1504 -151
rect 1532 -179 1570 -151
rect 1598 -179 1636 -151
rect 1664 -179 1702 -151
rect 1730 -179 1768 -151
rect 1796 -179 1834 -151
rect 1862 -179 1900 -151
rect 1928 -179 1966 -151
rect 1994 -179 2032 -151
rect 2060 -179 2098 -151
rect 2126 -179 2164 -151
rect 2192 -179 2230 -151
rect 2258 -179 2296 -151
rect 2324 -179 2362 -151
rect 2390 -179 2395 -151
rect -2395 -217 2395 -179
rect -2395 -245 -2390 -217
rect -2362 -245 -2324 -217
rect -2296 -245 -2258 -217
rect -2230 -245 -2192 -217
rect -2164 -245 -2126 -217
rect -2098 -245 -2060 -217
rect -2032 -245 -1994 -217
rect -1966 -245 -1928 -217
rect -1900 -245 -1862 -217
rect -1834 -245 -1796 -217
rect -1768 -245 -1730 -217
rect -1702 -245 -1664 -217
rect -1636 -245 -1598 -217
rect -1570 -245 -1532 -217
rect -1504 -245 -1466 -217
rect -1438 -245 -1400 -217
rect -1372 -245 -1334 -217
rect -1306 -245 -1268 -217
rect -1240 -245 -1202 -217
rect -1174 -245 -1136 -217
rect -1108 -245 -1070 -217
rect -1042 -245 -1004 -217
rect -976 -245 -938 -217
rect -910 -245 -872 -217
rect -844 -245 -806 -217
rect -778 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 778 -217
rect 806 -245 844 -217
rect 872 -245 910 -217
rect 938 -245 976 -217
rect 1004 -245 1042 -217
rect 1070 -245 1108 -217
rect 1136 -245 1174 -217
rect 1202 -245 1240 -217
rect 1268 -245 1306 -217
rect 1334 -245 1372 -217
rect 1400 -245 1438 -217
rect 1466 -245 1504 -217
rect 1532 -245 1570 -217
rect 1598 -245 1636 -217
rect 1664 -245 1702 -217
rect 1730 -245 1768 -217
rect 1796 -245 1834 -217
rect 1862 -245 1900 -217
rect 1928 -245 1966 -217
rect 1994 -245 2032 -217
rect 2060 -245 2098 -217
rect 2126 -245 2164 -217
rect 2192 -245 2230 -217
rect 2258 -245 2296 -217
rect 2324 -245 2362 -217
rect 2390 -245 2395 -217
rect -2395 -283 2395 -245
rect -2395 -311 -2390 -283
rect -2362 -311 -2324 -283
rect -2296 -311 -2258 -283
rect -2230 -311 -2192 -283
rect -2164 -311 -2126 -283
rect -2098 -311 -2060 -283
rect -2032 -311 -1994 -283
rect -1966 -311 -1928 -283
rect -1900 -311 -1862 -283
rect -1834 -311 -1796 -283
rect -1768 -311 -1730 -283
rect -1702 -311 -1664 -283
rect -1636 -311 -1598 -283
rect -1570 -311 -1532 -283
rect -1504 -311 -1466 -283
rect -1438 -311 -1400 -283
rect -1372 -311 -1334 -283
rect -1306 -311 -1268 -283
rect -1240 -311 -1202 -283
rect -1174 -311 -1136 -283
rect -1108 -311 -1070 -283
rect -1042 -311 -1004 -283
rect -976 -311 -938 -283
rect -910 -311 -872 -283
rect -844 -311 -806 -283
rect -778 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 778 -283
rect 806 -311 844 -283
rect 872 -311 910 -283
rect 938 -311 976 -283
rect 1004 -311 1042 -283
rect 1070 -311 1108 -283
rect 1136 -311 1174 -283
rect 1202 -311 1240 -283
rect 1268 -311 1306 -283
rect 1334 -311 1372 -283
rect 1400 -311 1438 -283
rect 1466 -311 1504 -283
rect 1532 -311 1570 -283
rect 1598 -311 1636 -283
rect 1664 -311 1702 -283
rect 1730 -311 1768 -283
rect 1796 -311 1834 -283
rect 1862 -311 1900 -283
rect 1928 -311 1966 -283
rect 1994 -311 2032 -283
rect 2060 -311 2098 -283
rect 2126 -311 2164 -283
rect 2192 -311 2230 -283
rect 2258 -311 2296 -283
rect 2324 -311 2362 -283
rect 2390 -311 2395 -283
rect -2395 -316 2395 -311
<< via4 >>
rect -2390 283 -2362 311
rect -2324 283 -2296 311
rect -2258 283 -2230 311
rect -2192 283 -2164 311
rect -2126 283 -2098 311
rect -2060 283 -2032 311
rect -1994 283 -1966 311
rect -1928 283 -1900 311
rect -1862 283 -1834 311
rect -1796 283 -1768 311
rect -1730 283 -1702 311
rect -1664 283 -1636 311
rect -1598 283 -1570 311
rect -1532 283 -1504 311
rect -1466 283 -1438 311
rect -1400 283 -1372 311
rect -1334 283 -1306 311
rect -1268 283 -1240 311
rect -1202 283 -1174 311
rect -1136 283 -1108 311
rect -1070 283 -1042 311
rect -1004 283 -976 311
rect -938 283 -910 311
rect -872 283 -844 311
rect -806 283 -778 311
rect -740 283 -712 311
rect -674 283 -646 311
rect -608 283 -580 311
rect -542 283 -514 311
rect -476 283 -448 311
rect -410 283 -382 311
rect -344 283 -316 311
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect 316 283 344 311
rect 382 283 410 311
rect 448 283 476 311
rect 514 283 542 311
rect 580 283 608 311
rect 646 283 674 311
rect 712 283 740 311
rect 778 283 806 311
rect 844 283 872 311
rect 910 283 938 311
rect 976 283 1004 311
rect 1042 283 1070 311
rect 1108 283 1136 311
rect 1174 283 1202 311
rect 1240 283 1268 311
rect 1306 283 1334 311
rect 1372 283 1400 311
rect 1438 283 1466 311
rect 1504 283 1532 311
rect 1570 283 1598 311
rect 1636 283 1664 311
rect 1702 283 1730 311
rect 1768 283 1796 311
rect 1834 283 1862 311
rect 1900 283 1928 311
rect 1966 283 1994 311
rect 2032 283 2060 311
rect 2098 283 2126 311
rect 2164 283 2192 311
rect 2230 283 2258 311
rect 2296 283 2324 311
rect 2362 283 2390 311
rect -2390 217 -2362 245
rect -2324 217 -2296 245
rect -2258 217 -2230 245
rect -2192 217 -2164 245
rect -2126 217 -2098 245
rect -2060 217 -2032 245
rect -1994 217 -1966 245
rect -1928 217 -1900 245
rect -1862 217 -1834 245
rect -1796 217 -1768 245
rect -1730 217 -1702 245
rect -1664 217 -1636 245
rect -1598 217 -1570 245
rect -1532 217 -1504 245
rect -1466 217 -1438 245
rect -1400 217 -1372 245
rect -1334 217 -1306 245
rect -1268 217 -1240 245
rect -1202 217 -1174 245
rect -1136 217 -1108 245
rect -1070 217 -1042 245
rect -1004 217 -976 245
rect -938 217 -910 245
rect -872 217 -844 245
rect -806 217 -778 245
rect -740 217 -712 245
rect -674 217 -646 245
rect -608 217 -580 245
rect -542 217 -514 245
rect -476 217 -448 245
rect -410 217 -382 245
rect -344 217 -316 245
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect 316 217 344 245
rect 382 217 410 245
rect 448 217 476 245
rect 514 217 542 245
rect 580 217 608 245
rect 646 217 674 245
rect 712 217 740 245
rect 778 217 806 245
rect 844 217 872 245
rect 910 217 938 245
rect 976 217 1004 245
rect 1042 217 1070 245
rect 1108 217 1136 245
rect 1174 217 1202 245
rect 1240 217 1268 245
rect 1306 217 1334 245
rect 1372 217 1400 245
rect 1438 217 1466 245
rect 1504 217 1532 245
rect 1570 217 1598 245
rect 1636 217 1664 245
rect 1702 217 1730 245
rect 1768 217 1796 245
rect 1834 217 1862 245
rect 1900 217 1928 245
rect 1966 217 1994 245
rect 2032 217 2060 245
rect 2098 217 2126 245
rect 2164 217 2192 245
rect 2230 217 2258 245
rect 2296 217 2324 245
rect 2362 217 2390 245
rect -2390 151 -2362 179
rect -2324 151 -2296 179
rect -2258 151 -2230 179
rect -2192 151 -2164 179
rect -2126 151 -2098 179
rect -2060 151 -2032 179
rect -1994 151 -1966 179
rect -1928 151 -1900 179
rect -1862 151 -1834 179
rect -1796 151 -1768 179
rect -1730 151 -1702 179
rect -1664 151 -1636 179
rect -1598 151 -1570 179
rect -1532 151 -1504 179
rect -1466 151 -1438 179
rect -1400 151 -1372 179
rect -1334 151 -1306 179
rect -1268 151 -1240 179
rect -1202 151 -1174 179
rect -1136 151 -1108 179
rect -1070 151 -1042 179
rect -1004 151 -976 179
rect -938 151 -910 179
rect -872 151 -844 179
rect -806 151 -778 179
rect -740 151 -712 179
rect -674 151 -646 179
rect -608 151 -580 179
rect -542 151 -514 179
rect -476 151 -448 179
rect -410 151 -382 179
rect -344 151 -316 179
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect 316 151 344 179
rect 382 151 410 179
rect 448 151 476 179
rect 514 151 542 179
rect 580 151 608 179
rect 646 151 674 179
rect 712 151 740 179
rect 778 151 806 179
rect 844 151 872 179
rect 910 151 938 179
rect 976 151 1004 179
rect 1042 151 1070 179
rect 1108 151 1136 179
rect 1174 151 1202 179
rect 1240 151 1268 179
rect 1306 151 1334 179
rect 1372 151 1400 179
rect 1438 151 1466 179
rect 1504 151 1532 179
rect 1570 151 1598 179
rect 1636 151 1664 179
rect 1702 151 1730 179
rect 1768 151 1796 179
rect 1834 151 1862 179
rect 1900 151 1928 179
rect 1966 151 1994 179
rect 2032 151 2060 179
rect 2098 151 2126 179
rect 2164 151 2192 179
rect 2230 151 2258 179
rect 2296 151 2324 179
rect 2362 151 2390 179
rect -2390 85 -2362 113
rect -2324 85 -2296 113
rect -2258 85 -2230 113
rect -2192 85 -2164 113
rect -2126 85 -2098 113
rect -2060 85 -2032 113
rect -1994 85 -1966 113
rect -1928 85 -1900 113
rect -1862 85 -1834 113
rect -1796 85 -1768 113
rect -1730 85 -1702 113
rect -1664 85 -1636 113
rect -1598 85 -1570 113
rect -1532 85 -1504 113
rect -1466 85 -1438 113
rect -1400 85 -1372 113
rect -1334 85 -1306 113
rect -1268 85 -1240 113
rect -1202 85 -1174 113
rect -1136 85 -1108 113
rect -1070 85 -1042 113
rect -1004 85 -976 113
rect -938 85 -910 113
rect -872 85 -844 113
rect -806 85 -778 113
rect -740 85 -712 113
rect -674 85 -646 113
rect -608 85 -580 113
rect -542 85 -514 113
rect -476 85 -448 113
rect -410 85 -382 113
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect 382 85 410 113
rect 448 85 476 113
rect 514 85 542 113
rect 580 85 608 113
rect 646 85 674 113
rect 712 85 740 113
rect 778 85 806 113
rect 844 85 872 113
rect 910 85 938 113
rect 976 85 1004 113
rect 1042 85 1070 113
rect 1108 85 1136 113
rect 1174 85 1202 113
rect 1240 85 1268 113
rect 1306 85 1334 113
rect 1372 85 1400 113
rect 1438 85 1466 113
rect 1504 85 1532 113
rect 1570 85 1598 113
rect 1636 85 1664 113
rect 1702 85 1730 113
rect 1768 85 1796 113
rect 1834 85 1862 113
rect 1900 85 1928 113
rect 1966 85 1994 113
rect 2032 85 2060 113
rect 2098 85 2126 113
rect 2164 85 2192 113
rect 2230 85 2258 113
rect 2296 85 2324 113
rect 2362 85 2390 113
rect -2390 19 -2362 47
rect -2324 19 -2296 47
rect -2258 19 -2230 47
rect -2192 19 -2164 47
rect -2126 19 -2098 47
rect -2060 19 -2032 47
rect -1994 19 -1966 47
rect -1928 19 -1900 47
rect -1862 19 -1834 47
rect -1796 19 -1768 47
rect -1730 19 -1702 47
rect -1664 19 -1636 47
rect -1598 19 -1570 47
rect -1532 19 -1504 47
rect -1466 19 -1438 47
rect -1400 19 -1372 47
rect -1334 19 -1306 47
rect -1268 19 -1240 47
rect -1202 19 -1174 47
rect -1136 19 -1108 47
rect -1070 19 -1042 47
rect -1004 19 -976 47
rect -938 19 -910 47
rect -872 19 -844 47
rect -806 19 -778 47
rect -740 19 -712 47
rect -674 19 -646 47
rect -608 19 -580 47
rect -542 19 -514 47
rect -476 19 -448 47
rect -410 19 -382 47
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect 382 19 410 47
rect 448 19 476 47
rect 514 19 542 47
rect 580 19 608 47
rect 646 19 674 47
rect 712 19 740 47
rect 778 19 806 47
rect 844 19 872 47
rect 910 19 938 47
rect 976 19 1004 47
rect 1042 19 1070 47
rect 1108 19 1136 47
rect 1174 19 1202 47
rect 1240 19 1268 47
rect 1306 19 1334 47
rect 1372 19 1400 47
rect 1438 19 1466 47
rect 1504 19 1532 47
rect 1570 19 1598 47
rect 1636 19 1664 47
rect 1702 19 1730 47
rect 1768 19 1796 47
rect 1834 19 1862 47
rect 1900 19 1928 47
rect 1966 19 1994 47
rect 2032 19 2060 47
rect 2098 19 2126 47
rect 2164 19 2192 47
rect 2230 19 2258 47
rect 2296 19 2324 47
rect 2362 19 2390 47
rect -2390 -47 -2362 -19
rect -2324 -47 -2296 -19
rect -2258 -47 -2230 -19
rect -2192 -47 -2164 -19
rect -2126 -47 -2098 -19
rect -2060 -47 -2032 -19
rect -1994 -47 -1966 -19
rect -1928 -47 -1900 -19
rect -1862 -47 -1834 -19
rect -1796 -47 -1768 -19
rect -1730 -47 -1702 -19
rect -1664 -47 -1636 -19
rect -1598 -47 -1570 -19
rect -1532 -47 -1504 -19
rect -1466 -47 -1438 -19
rect -1400 -47 -1372 -19
rect -1334 -47 -1306 -19
rect -1268 -47 -1240 -19
rect -1202 -47 -1174 -19
rect -1136 -47 -1108 -19
rect -1070 -47 -1042 -19
rect -1004 -47 -976 -19
rect -938 -47 -910 -19
rect -872 -47 -844 -19
rect -806 -47 -778 -19
rect -740 -47 -712 -19
rect -674 -47 -646 -19
rect -608 -47 -580 -19
rect -542 -47 -514 -19
rect -476 -47 -448 -19
rect -410 -47 -382 -19
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect 382 -47 410 -19
rect 448 -47 476 -19
rect 514 -47 542 -19
rect 580 -47 608 -19
rect 646 -47 674 -19
rect 712 -47 740 -19
rect 778 -47 806 -19
rect 844 -47 872 -19
rect 910 -47 938 -19
rect 976 -47 1004 -19
rect 1042 -47 1070 -19
rect 1108 -47 1136 -19
rect 1174 -47 1202 -19
rect 1240 -47 1268 -19
rect 1306 -47 1334 -19
rect 1372 -47 1400 -19
rect 1438 -47 1466 -19
rect 1504 -47 1532 -19
rect 1570 -47 1598 -19
rect 1636 -47 1664 -19
rect 1702 -47 1730 -19
rect 1768 -47 1796 -19
rect 1834 -47 1862 -19
rect 1900 -47 1928 -19
rect 1966 -47 1994 -19
rect 2032 -47 2060 -19
rect 2098 -47 2126 -19
rect 2164 -47 2192 -19
rect 2230 -47 2258 -19
rect 2296 -47 2324 -19
rect 2362 -47 2390 -19
rect -2390 -113 -2362 -85
rect -2324 -113 -2296 -85
rect -2258 -113 -2230 -85
rect -2192 -113 -2164 -85
rect -2126 -113 -2098 -85
rect -2060 -113 -2032 -85
rect -1994 -113 -1966 -85
rect -1928 -113 -1900 -85
rect -1862 -113 -1834 -85
rect -1796 -113 -1768 -85
rect -1730 -113 -1702 -85
rect -1664 -113 -1636 -85
rect -1598 -113 -1570 -85
rect -1532 -113 -1504 -85
rect -1466 -113 -1438 -85
rect -1400 -113 -1372 -85
rect -1334 -113 -1306 -85
rect -1268 -113 -1240 -85
rect -1202 -113 -1174 -85
rect -1136 -113 -1108 -85
rect -1070 -113 -1042 -85
rect -1004 -113 -976 -85
rect -938 -113 -910 -85
rect -872 -113 -844 -85
rect -806 -113 -778 -85
rect -740 -113 -712 -85
rect -674 -113 -646 -85
rect -608 -113 -580 -85
rect -542 -113 -514 -85
rect -476 -113 -448 -85
rect -410 -113 -382 -85
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect 382 -113 410 -85
rect 448 -113 476 -85
rect 514 -113 542 -85
rect 580 -113 608 -85
rect 646 -113 674 -85
rect 712 -113 740 -85
rect 778 -113 806 -85
rect 844 -113 872 -85
rect 910 -113 938 -85
rect 976 -113 1004 -85
rect 1042 -113 1070 -85
rect 1108 -113 1136 -85
rect 1174 -113 1202 -85
rect 1240 -113 1268 -85
rect 1306 -113 1334 -85
rect 1372 -113 1400 -85
rect 1438 -113 1466 -85
rect 1504 -113 1532 -85
rect 1570 -113 1598 -85
rect 1636 -113 1664 -85
rect 1702 -113 1730 -85
rect 1768 -113 1796 -85
rect 1834 -113 1862 -85
rect 1900 -113 1928 -85
rect 1966 -113 1994 -85
rect 2032 -113 2060 -85
rect 2098 -113 2126 -85
rect 2164 -113 2192 -85
rect 2230 -113 2258 -85
rect 2296 -113 2324 -85
rect 2362 -113 2390 -85
rect -2390 -179 -2362 -151
rect -2324 -179 -2296 -151
rect -2258 -179 -2230 -151
rect -2192 -179 -2164 -151
rect -2126 -179 -2098 -151
rect -2060 -179 -2032 -151
rect -1994 -179 -1966 -151
rect -1928 -179 -1900 -151
rect -1862 -179 -1834 -151
rect -1796 -179 -1768 -151
rect -1730 -179 -1702 -151
rect -1664 -179 -1636 -151
rect -1598 -179 -1570 -151
rect -1532 -179 -1504 -151
rect -1466 -179 -1438 -151
rect -1400 -179 -1372 -151
rect -1334 -179 -1306 -151
rect -1268 -179 -1240 -151
rect -1202 -179 -1174 -151
rect -1136 -179 -1108 -151
rect -1070 -179 -1042 -151
rect -1004 -179 -976 -151
rect -938 -179 -910 -151
rect -872 -179 -844 -151
rect -806 -179 -778 -151
rect -740 -179 -712 -151
rect -674 -179 -646 -151
rect -608 -179 -580 -151
rect -542 -179 -514 -151
rect -476 -179 -448 -151
rect -410 -179 -382 -151
rect -344 -179 -316 -151
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect 316 -179 344 -151
rect 382 -179 410 -151
rect 448 -179 476 -151
rect 514 -179 542 -151
rect 580 -179 608 -151
rect 646 -179 674 -151
rect 712 -179 740 -151
rect 778 -179 806 -151
rect 844 -179 872 -151
rect 910 -179 938 -151
rect 976 -179 1004 -151
rect 1042 -179 1070 -151
rect 1108 -179 1136 -151
rect 1174 -179 1202 -151
rect 1240 -179 1268 -151
rect 1306 -179 1334 -151
rect 1372 -179 1400 -151
rect 1438 -179 1466 -151
rect 1504 -179 1532 -151
rect 1570 -179 1598 -151
rect 1636 -179 1664 -151
rect 1702 -179 1730 -151
rect 1768 -179 1796 -151
rect 1834 -179 1862 -151
rect 1900 -179 1928 -151
rect 1966 -179 1994 -151
rect 2032 -179 2060 -151
rect 2098 -179 2126 -151
rect 2164 -179 2192 -151
rect 2230 -179 2258 -151
rect 2296 -179 2324 -151
rect 2362 -179 2390 -151
rect -2390 -245 -2362 -217
rect -2324 -245 -2296 -217
rect -2258 -245 -2230 -217
rect -2192 -245 -2164 -217
rect -2126 -245 -2098 -217
rect -2060 -245 -2032 -217
rect -1994 -245 -1966 -217
rect -1928 -245 -1900 -217
rect -1862 -245 -1834 -217
rect -1796 -245 -1768 -217
rect -1730 -245 -1702 -217
rect -1664 -245 -1636 -217
rect -1598 -245 -1570 -217
rect -1532 -245 -1504 -217
rect -1466 -245 -1438 -217
rect -1400 -245 -1372 -217
rect -1334 -245 -1306 -217
rect -1268 -245 -1240 -217
rect -1202 -245 -1174 -217
rect -1136 -245 -1108 -217
rect -1070 -245 -1042 -217
rect -1004 -245 -976 -217
rect -938 -245 -910 -217
rect -872 -245 -844 -217
rect -806 -245 -778 -217
rect -740 -245 -712 -217
rect -674 -245 -646 -217
rect -608 -245 -580 -217
rect -542 -245 -514 -217
rect -476 -245 -448 -217
rect -410 -245 -382 -217
rect -344 -245 -316 -217
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect 316 -245 344 -217
rect 382 -245 410 -217
rect 448 -245 476 -217
rect 514 -245 542 -217
rect 580 -245 608 -217
rect 646 -245 674 -217
rect 712 -245 740 -217
rect 778 -245 806 -217
rect 844 -245 872 -217
rect 910 -245 938 -217
rect 976 -245 1004 -217
rect 1042 -245 1070 -217
rect 1108 -245 1136 -217
rect 1174 -245 1202 -217
rect 1240 -245 1268 -217
rect 1306 -245 1334 -217
rect 1372 -245 1400 -217
rect 1438 -245 1466 -217
rect 1504 -245 1532 -217
rect 1570 -245 1598 -217
rect 1636 -245 1664 -217
rect 1702 -245 1730 -217
rect 1768 -245 1796 -217
rect 1834 -245 1862 -217
rect 1900 -245 1928 -217
rect 1966 -245 1994 -217
rect 2032 -245 2060 -217
rect 2098 -245 2126 -217
rect 2164 -245 2192 -217
rect 2230 -245 2258 -217
rect 2296 -245 2324 -217
rect 2362 -245 2390 -217
rect -2390 -311 -2362 -283
rect -2324 -311 -2296 -283
rect -2258 -311 -2230 -283
rect -2192 -311 -2164 -283
rect -2126 -311 -2098 -283
rect -2060 -311 -2032 -283
rect -1994 -311 -1966 -283
rect -1928 -311 -1900 -283
rect -1862 -311 -1834 -283
rect -1796 -311 -1768 -283
rect -1730 -311 -1702 -283
rect -1664 -311 -1636 -283
rect -1598 -311 -1570 -283
rect -1532 -311 -1504 -283
rect -1466 -311 -1438 -283
rect -1400 -311 -1372 -283
rect -1334 -311 -1306 -283
rect -1268 -311 -1240 -283
rect -1202 -311 -1174 -283
rect -1136 -311 -1108 -283
rect -1070 -311 -1042 -283
rect -1004 -311 -976 -283
rect -938 -311 -910 -283
rect -872 -311 -844 -283
rect -806 -311 -778 -283
rect -740 -311 -712 -283
rect -674 -311 -646 -283
rect -608 -311 -580 -283
rect -542 -311 -514 -283
rect -476 -311 -448 -283
rect -410 -311 -382 -283
rect -344 -311 -316 -283
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
rect 316 -311 344 -283
rect 382 -311 410 -283
rect 448 -311 476 -283
rect 514 -311 542 -283
rect 580 -311 608 -283
rect 646 -311 674 -283
rect 712 -311 740 -283
rect 778 -311 806 -283
rect 844 -311 872 -283
rect 910 -311 938 -283
rect 976 -311 1004 -283
rect 1042 -311 1070 -283
rect 1108 -311 1136 -283
rect 1174 -311 1202 -283
rect 1240 -311 1268 -283
rect 1306 -311 1334 -283
rect 1372 -311 1400 -283
rect 1438 -311 1466 -283
rect 1504 -311 1532 -283
rect 1570 -311 1598 -283
rect 1636 -311 1664 -283
rect 1702 -311 1730 -283
rect 1768 -311 1796 -283
rect 1834 -311 1862 -283
rect 1900 -311 1928 -283
rect 1966 -311 1994 -283
rect 2032 -311 2060 -283
rect 2098 -311 2126 -283
rect 2164 -311 2192 -283
rect 2230 -311 2258 -283
rect 2296 -311 2324 -283
rect 2362 -311 2390 -283
<< metal5 >>
rect -2398 311 2398 319
rect -2398 283 -2390 311
rect -2362 283 -2324 311
rect -2296 283 -2258 311
rect -2230 283 -2192 311
rect -2164 283 -2126 311
rect -2098 283 -2060 311
rect -2032 283 -1994 311
rect -1966 283 -1928 311
rect -1900 283 -1862 311
rect -1834 283 -1796 311
rect -1768 283 -1730 311
rect -1702 283 -1664 311
rect -1636 283 -1598 311
rect -1570 283 -1532 311
rect -1504 283 -1466 311
rect -1438 283 -1400 311
rect -1372 283 -1334 311
rect -1306 283 -1268 311
rect -1240 283 -1202 311
rect -1174 283 -1136 311
rect -1108 283 -1070 311
rect -1042 283 -1004 311
rect -976 283 -938 311
rect -910 283 -872 311
rect -844 283 -806 311
rect -778 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 778 311
rect 806 283 844 311
rect 872 283 910 311
rect 938 283 976 311
rect 1004 283 1042 311
rect 1070 283 1108 311
rect 1136 283 1174 311
rect 1202 283 1240 311
rect 1268 283 1306 311
rect 1334 283 1372 311
rect 1400 283 1438 311
rect 1466 283 1504 311
rect 1532 283 1570 311
rect 1598 283 1636 311
rect 1664 283 1702 311
rect 1730 283 1768 311
rect 1796 283 1834 311
rect 1862 283 1900 311
rect 1928 283 1966 311
rect 1994 283 2032 311
rect 2060 283 2098 311
rect 2126 283 2164 311
rect 2192 283 2230 311
rect 2258 283 2296 311
rect 2324 283 2362 311
rect 2390 283 2398 311
rect -2398 245 2398 283
rect -2398 217 -2390 245
rect -2362 217 -2324 245
rect -2296 217 -2258 245
rect -2230 217 -2192 245
rect -2164 217 -2126 245
rect -2098 217 -2060 245
rect -2032 217 -1994 245
rect -1966 217 -1928 245
rect -1900 217 -1862 245
rect -1834 217 -1796 245
rect -1768 217 -1730 245
rect -1702 217 -1664 245
rect -1636 217 -1598 245
rect -1570 217 -1532 245
rect -1504 217 -1466 245
rect -1438 217 -1400 245
rect -1372 217 -1334 245
rect -1306 217 -1268 245
rect -1240 217 -1202 245
rect -1174 217 -1136 245
rect -1108 217 -1070 245
rect -1042 217 -1004 245
rect -976 217 -938 245
rect -910 217 -872 245
rect -844 217 -806 245
rect -778 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 778 245
rect 806 217 844 245
rect 872 217 910 245
rect 938 217 976 245
rect 1004 217 1042 245
rect 1070 217 1108 245
rect 1136 217 1174 245
rect 1202 217 1240 245
rect 1268 217 1306 245
rect 1334 217 1372 245
rect 1400 217 1438 245
rect 1466 217 1504 245
rect 1532 217 1570 245
rect 1598 217 1636 245
rect 1664 217 1702 245
rect 1730 217 1768 245
rect 1796 217 1834 245
rect 1862 217 1900 245
rect 1928 217 1966 245
rect 1994 217 2032 245
rect 2060 217 2098 245
rect 2126 217 2164 245
rect 2192 217 2230 245
rect 2258 217 2296 245
rect 2324 217 2362 245
rect 2390 217 2398 245
rect -2398 179 2398 217
rect -2398 151 -2390 179
rect -2362 151 -2324 179
rect -2296 151 -2258 179
rect -2230 151 -2192 179
rect -2164 151 -2126 179
rect -2098 151 -2060 179
rect -2032 151 -1994 179
rect -1966 151 -1928 179
rect -1900 151 -1862 179
rect -1834 151 -1796 179
rect -1768 151 -1730 179
rect -1702 151 -1664 179
rect -1636 151 -1598 179
rect -1570 151 -1532 179
rect -1504 151 -1466 179
rect -1438 151 -1400 179
rect -1372 151 -1334 179
rect -1306 151 -1268 179
rect -1240 151 -1202 179
rect -1174 151 -1136 179
rect -1108 151 -1070 179
rect -1042 151 -1004 179
rect -976 151 -938 179
rect -910 151 -872 179
rect -844 151 -806 179
rect -778 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 778 179
rect 806 151 844 179
rect 872 151 910 179
rect 938 151 976 179
rect 1004 151 1042 179
rect 1070 151 1108 179
rect 1136 151 1174 179
rect 1202 151 1240 179
rect 1268 151 1306 179
rect 1334 151 1372 179
rect 1400 151 1438 179
rect 1466 151 1504 179
rect 1532 151 1570 179
rect 1598 151 1636 179
rect 1664 151 1702 179
rect 1730 151 1768 179
rect 1796 151 1834 179
rect 1862 151 1900 179
rect 1928 151 1966 179
rect 1994 151 2032 179
rect 2060 151 2098 179
rect 2126 151 2164 179
rect 2192 151 2230 179
rect 2258 151 2296 179
rect 2324 151 2362 179
rect 2390 151 2398 179
rect -2398 113 2398 151
rect -2398 85 -2390 113
rect -2362 85 -2324 113
rect -2296 85 -2258 113
rect -2230 85 -2192 113
rect -2164 85 -2126 113
rect -2098 85 -2060 113
rect -2032 85 -1994 113
rect -1966 85 -1928 113
rect -1900 85 -1862 113
rect -1834 85 -1796 113
rect -1768 85 -1730 113
rect -1702 85 -1664 113
rect -1636 85 -1598 113
rect -1570 85 -1532 113
rect -1504 85 -1466 113
rect -1438 85 -1400 113
rect -1372 85 -1334 113
rect -1306 85 -1268 113
rect -1240 85 -1202 113
rect -1174 85 -1136 113
rect -1108 85 -1070 113
rect -1042 85 -1004 113
rect -976 85 -938 113
rect -910 85 -872 113
rect -844 85 -806 113
rect -778 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 778 113
rect 806 85 844 113
rect 872 85 910 113
rect 938 85 976 113
rect 1004 85 1042 113
rect 1070 85 1108 113
rect 1136 85 1174 113
rect 1202 85 1240 113
rect 1268 85 1306 113
rect 1334 85 1372 113
rect 1400 85 1438 113
rect 1466 85 1504 113
rect 1532 85 1570 113
rect 1598 85 1636 113
rect 1664 85 1702 113
rect 1730 85 1768 113
rect 1796 85 1834 113
rect 1862 85 1900 113
rect 1928 85 1966 113
rect 1994 85 2032 113
rect 2060 85 2098 113
rect 2126 85 2164 113
rect 2192 85 2230 113
rect 2258 85 2296 113
rect 2324 85 2362 113
rect 2390 85 2398 113
rect -2398 47 2398 85
rect -2398 19 -2390 47
rect -2362 19 -2324 47
rect -2296 19 -2258 47
rect -2230 19 -2192 47
rect -2164 19 -2126 47
rect -2098 19 -2060 47
rect -2032 19 -1994 47
rect -1966 19 -1928 47
rect -1900 19 -1862 47
rect -1834 19 -1796 47
rect -1768 19 -1730 47
rect -1702 19 -1664 47
rect -1636 19 -1598 47
rect -1570 19 -1532 47
rect -1504 19 -1466 47
rect -1438 19 -1400 47
rect -1372 19 -1334 47
rect -1306 19 -1268 47
rect -1240 19 -1202 47
rect -1174 19 -1136 47
rect -1108 19 -1070 47
rect -1042 19 -1004 47
rect -976 19 -938 47
rect -910 19 -872 47
rect -844 19 -806 47
rect -778 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 778 47
rect 806 19 844 47
rect 872 19 910 47
rect 938 19 976 47
rect 1004 19 1042 47
rect 1070 19 1108 47
rect 1136 19 1174 47
rect 1202 19 1240 47
rect 1268 19 1306 47
rect 1334 19 1372 47
rect 1400 19 1438 47
rect 1466 19 1504 47
rect 1532 19 1570 47
rect 1598 19 1636 47
rect 1664 19 1702 47
rect 1730 19 1768 47
rect 1796 19 1834 47
rect 1862 19 1900 47
rect 1928 19 1966 47
rect 1994 19 2032 47
rect 2060 19 2098 47
rect 2126 19 2164 47
rect 2192 19 2230 47
rect 2258 19 2296 47
rect 2324 19 2362 47
rect 2390 19 2398 47
rect -2398 -19 2398 19
rect -2398 -47 -2390 -19
rect -2362 -47 -2324 -19
rect -2296 -47 -2258 -19
rect -2230 -47 -2192 -19
rect -2164 -47 -2126 -19
rect -2098 -47 -2060 -19
rect -2032 -47 -1994 -19
rect -1966 -47 -1928 -19
rect -1900 -47 -1862 -19
rect -1834 -47 -1796 -19
rect -1768 -47 -1730 -19
rect -1702 -47 -1664 -19
rect -1636 -47 -1598 -19
rect -1570 -47 -1532 -19
rect -1504 -47 -1466 -19
rect -1438 -47 -1400 -19
rect -1372 -47 -1334 -19
rect -1306 -47 -1268 -19
rect -1240 -47 -1202 -19
rect -1174 -47 -1136 -19
rect -1108 -47 -1070 -19
rect -1042 -47 -1004 -19
rect -976 -47 -938 -19
rect -910 -47 -872 -19
rect -844 -47 -806 -19
rect -778 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 778 -19
rect 806 -47 844 -19
rect 872 -47 910 -19
rect 938 -47 976 -19
rect 1004 -47 1042 -19
rect 1070 -47 1108 -19
rect 1136 -47 1174 -19
rect 1202 -47 1240 -19
rect 1268 -47 1306 -19
rect 1334 -47 1372 -19
rect 1400 -47 1438 -19
rect 1466 -47 1504 -19
rect 1532 -47 1570 -19
rect 1598 -47 1636 -19
rect 1664 -47 1702 -19
rect 1730 -47 1768 -19
rect 1796 -47 1834 -19
rect 1862 -47 1900 -19
rect 1928 -47 1966 -19
rect 1994 -47 2032 -19
rect 2060 -47 2098 -19
rect 2126 -47 2164 -19
rect 2192 -47 2230 -19
rect 2258 -47 2296 -19
rect 2324 -47 2362 -19
rect 2390 -47 2398 -19
rect -2398 -85 2398 -47
rect -2398 -113 -2390 -85
rect -2362 -113 -2324 -85
rect -2296 -113 -2258 -85
rect -2230 -113 -2192 -85
rect -2164 -113 -2126 -85
rect -2098 -113 -2060 -85
rect -2032 -113 -1994 -85
rect -1966 -113 -1928 -85
rect -1900 -113 -1862 -85
rect -1834 -113 -1796 -85
rect -1768 -113 -1730 -85
rect -1702 -113 -1664 -85
rect -1636 -113 -1598 -85
rect -1570 -113 -1532 -85
rect -1504 -113 -1466 -85
rect -1438 -113 -1400 -85
rect -1372 -113 -1334 -85
rect -1306 -113 -1268 -85
rect -1240 -113 -1202 -85
rect -1174 -113 -1136 -85
rect -1108 -113 -1070 -85
rect -1042 -113 -1004 -85
rect -976 -113 -938 -85
rect -910 -113 -872 -85
rect -844 -113 -806 -85
rect -778 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 778 -85
rect 806 -113 844 -85
rect 872 -113 910 -85
rect 938 -113 976 -85
rect 1004 -113 1042 -85
rect 1070 -113 1108 -85
rect 1136 -113 1174 -85
rect 1202 -113 1240 -85
rect 1268 -113 1306 -85
rect 1334 -113 1372 -85
rect 1400 -113 1438 -85
rect 1466 -113 1504 -85
rect 1532 -113 1570 -85
rect 1598 -113 1636 -85
rect 1664 -113 1702 -85
rect 1730 -113 1768 -85
rect 1796 -113 1834 -85
rect 1862 -113 1900 -85
rect 1928 -113 1966 -85
rect 1994 -113 2032 -85
rect 2060 -113 2098 -85
rect 2126 -113 2164 -85
rect 2192 -113 2230 -85
rect 2258 -113 2296 -85
rect 2324 -113 2362 -85
rect 2390 -113 2398 -85
rect -2398 -151 2398 -113
rect -2398 -179 -2390 -151
rect -2362 -179 -2324 -151
rect -2296 -179 -2258 -151
rect -2230 -179 -2192 -151
rect -2164 -179 -2126 -151
rect -2098 -179 -2060 -151
rect -2032 -179 -1994 -151
rect -1966 -179 -1928 -151
rect -1900 -179 -1862 -151
rect -1834 -179 -1796 -151
rect -1768 -179 -1730 -151
rect -1702 -179 -1664 -151
rect -1636 -179 -1598 -151
rect -1570 -179 -1532 -151
rect -1504 -179 -1466 -151
rect -1438 -179 -1400 -151
rect -1372 -179 -1334 -151
rect -1306 -179 -1268 -151
rect -1240 -179 -1202 -151
rect -1174 -179 -1136 -151
rect -1108 -179 -1070 -151
rect -1042 -179 -1004 -151
rect -976 -179 -938 -151
rect -910 -179 -872 -151
rect -844 -179 -806 -151
rect -778 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 778 -151
rect 806 -179 844 -151
rect 872 -179 910 -151
rect 938 -179 976 -151
rect 1004 -179 1042 -151
rect 1070 -179 1108 -151
rect 1136 -179 1174 -151
rect 1202 -179 1240 -151
rect 1268 -179 1306 -151
rect 1334 -179 1372 -151
rect 1400 -179 1438 -151
rect 1466 -179 1504 -151
rect 1532 -179 1570 -151
rect 1598 -179 1636 -151
rect 1664 -179 1702 -151
rect 1730 -179 1768 -151
rect 1796 -179 1834 -151
rect 1862 -179 1900 -151
rect 1928 -179 1966 -151
rect 1994 -179 2032 -151
rect 2060 -179 2098 -151
rect 2126 -179 2164 -151
rect 2192 -179 2230 -151
rect 2258 -179 2296 -151
rect 2324 -179 2362 -151
rect 2390 -179 2398 -151
rect -2398 -217 2398 -179
rect -2398 -245 -2390 -217
rect -2362 -245 -2324 -217
rect -2296 -245 -2258 -217
rect -2230 -245 -2192 -217
rect -2164 -245 -2126 -217
rect -2098 -245 -2060 -217
rect -2032 -245 -1994 -217
rect -1966 -245 -1928 -217
rect -1900 -245 -1862 -217
rect -1834 -245 -1796 -217
rect -1768 -245 -1730 -217
rect -1702 -245 -1664 -217
rect -1636 -245 -1598 -217
rect -1570 -245 -1532 -217
rect -1504 -245 -1466 -217
rect -1438 -245 -1400 -217
rect -1372 -245 -1334 -217
rect -1306 -245 -1268 -217
rect -1240 -245 -1202 -217
rect -1174 -245 -1136 -217
rect -1108 -245 -1070 -217
rect -1042 -245 -1004 -217
rect -976 -245 -938 -217
rect -910 -245 -872 -217
rect -844 -245 -806 -217
rect -778 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 778 -217
rect 806 -245 844 -217
rect 872 -245 910 -217
rect 938 -245 976 -217
rect 1004 -245 1042 -217
rect 1070 -245 1108 -217
rect 1136 -245 1174 -217
rect 1202 -245 1240 -217
rect 1268 -245 1306 -217
rect 1334 -245 1372 -217
rect 1400 -245 1438 -217
rect 1466 -245 1504 -217
rect 1532 -245 1570 -217
rect 1598 -245 1636 -217
rect 1664 -245 1702 -217
rect 1730 -245 1768 -217
rect 1796 -245 1834 -217
rect 1862 -245 1900 -217
rect 1928 -245 1966 -217
rect 1994 -245 2032 -217
rect 2060 -245 2098 -217
rect 2126 -245 2164 -217
rect 2192 -245 2230 -217
rect 2258 -245 2296 -217
rect 2324 -245 2362 -217
rect 2390 -245 2398 -217
rect -2398 -283 2398 -245
rect -2398 -311 -2390 -283
rect -2362 -311 -2324 -283
rect -2296 -311 -2258 -283
rect -2230 -311 -2192 -283
rect -2164 -311 -2126 -283
rect -2098 -311 -2060 -283
rect -2032 -311 -1994 -283
rect -1966 -311 -1928 -283
rect -1900 -311 -1862 -283
rect -1834 -311 -1796 -283
rect -1768 -311 -1730 -283
rect -1702 -311 -1664 -283
rect -1636 -311 -1598 -283
rect -1570 -311 -1532 -283
rect -1504 -311 -1466 -283
rect -1438 -311 -1400 -283
rect -1372 -311 -1334 -283
rect -1306 -311 -1268 -283
rect -1240 -311 -1202 -283
rect -1174 -311 -1136 -283
rect -1108 -311 -1070 -283
rect -1042 -311 -1004 -283
rect -976 -311 -938 -283
rect -910 -311 -872 -283
rect -844 -311 -806 -283
rect -778 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 778 -283
rect 806 -311 844 -283
rect 872 -311 910 -283
rect 938 -311 976 -283
rect 1004 -311 1042 -283
rect 1070 -311 1108 -283
rect 1136 -311 1174 -283
rect 1202 -311 1240 -283
rect 1268 -311 1306 -283
rect 1334 -311 1372 -283
rect 1400 -311 1438 -283
rect 1466 -311 1504 -283
rect 1532 -311 1570 -283
rect 1598 -311 1636 -283
rect 1664 -311 1702 -283
rect 1730 -311 1768 -283
rect 1796 -311 1834 -283
rect 1862 -311 1900 -283
rect 1928 -311 1966 -283
rect 1994 -311 2032 -283
rect 2060 -311 2098 -283
rect 2126 -311 2164 -283
rect 2192 -311 2230 -283
rect 2258 -311 2296 -283
rect 2324 -311 2362 -283
rect 2390 -311 2398 -283
rect -2398 -319 2398 -311
<< end >>
