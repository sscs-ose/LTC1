magic
tech gf180mcuC
magscale 1 10
timestamp 1692335619
<< pwell >>
rect -700 -579 700 579
<< nmos >>
rect -588 261 -532 511
rect -428 261 -372 511
rect -268 261 -212 511
rect -108 261 -52 511
rect 52 261 108 511
rect 212 261 268 511
rect 372 261 428 511
rect 532 261 588 511
rect -588 -125 -532 125
rect -428 -125 -372 125
rect -268 -125 -212 125
rect -108 -125 -52 125
rect 52 -125 108 125
rect 212 -125 268 125
rect 372 -125 428 125
rect 532 -125 588 125
rect -588 -511 -532 -261
rect -428 -511 -372 -261
rect -268 -511 -212 -261
rect -108 -511 -52 -261
rect 52 -511 108 -261
rect 212 -511 268 -261
rect 372 -511 428 -261
rect 532 -511 588 -261
<< ndiff >>
rect -676 498 -588 511
rect -676 274 -663 498
rect -617 274 -588 498
rect -676 261 -588 274
rect -532 498 -428 511
rect -532 274 -503 498
rect -457 274 -428 498
rect -532 261 -428 274
rect -372 498 -268 511
rect -372 274 -343 498
rect -297 274 -268 498
rect -372 261 -268 274
rect -212 498 -108 511
rect -212 274 -183 498
rect -137 274 -108 498
rect -212 261 -108 274
rect -52 498 52 511
rect -52 274 -23 498
rect 23 274 52 498
rect -52 261 52 274
rect 108 498 212 511
rect 108 274 137 498
rect 183 274 212 498
rect 108 261 212 274
rect 268 498 372 511
rect 268 274 297 498
rect 343 274 372 498
rect 268 261 372 274
rect 428 498 532 511
rect 428 274 457 498
rect 503 274 532 498
rect 428 261 532 274
rect 588 498 676 511
rect 588 274 617 498
rect 663 274 676 498
rect 588 261 676 274
rect -676 112 -588 125
rect -676 -112 -663 112
rect -617 -112 -588 112
rect -676 -125 -588 -112
rect -532 112 -428 125
rect -532 -112 -503 112
rect -457 -112 -428 112
rect -532 -125 -428 -112
rect -372 112 -268 125
rect -372 -112 -343 112
rect -297 -112 -268 112
rect -372 -125 -268 -112
rect -212 112 -108 125
rect -212 -112 -183 112
rect -137 -112 -108 112
rect -212 -125 -108 -112
rect -52 112 52 125
rect -52 -112 -23 112
rect 23 -112 52 112
rect -52 -125 52 -112
rect 108 112 212 125
rect 108 -112 137 112
rect 183 -112 212 112
rect 108 -125 212 -112
rect 268 112 372 125
rect 268 -112 297 112
rect 343 -112 372 112
rect 268 -125 372 -112
rect 428 112 532 125
rect 428 -112 457 112
rect 503 -112 532 112
rect 428 -125 532 -112
rect 588 112 676 125
rect 588 -112 617 112
rect 663 -112 676 112
rect 588 -125 676 -112
rect -676 -274 -588 -261
rect -676 -498 -663 -274
rect -617 -498 -588 -274
rect -676 -511 -588 -498
rect -532 -274 -428 -261
rect -532 -498 -503 -274
rect -457 -498 -428 -274
rect -532 -511 -428 -498
rect -372 -274 -268 -261
rect -372 -498 -343 -274
rect -297 -498 -268 -274
rect -372 -511 -268 -498
rect -212 -274 -108 -261
rect -212 -498 -183 -274
rect -137 -498 -108 -274
rect -212 -511 -108 -498
rect -52 -274 52 -261
rect -52 -498 -23 -274
rect 23 -498 52 -274
rect -52 -511 52 -498
rect 108 -274 212 -261
rect 108 -498 137 -274
rect 183 -498 212 -274
rect 108 -511 212 -498
rect 268 -274 372 -261
rect 268 -498 297 -274
rect 343 -498 372 -274
rect 268 -511 372 -498
rect 428 -274 532 -261
rect 428 -498 457 -274
rect 503 -498 532 -274
rect 428 -511 532 -498
rect 588 -274 676 -261
rect 588 -498 617 -274
rect 663 -498 676 -274
rect 588 -511 676 -498
<< ndiffc >>
rect -663 274 -617 498
rect -503 274 -457 498
rect -343 274 -297 498
rect -183 274 -137 498
rect -23 274 23 498
rect 137 274 183 498
rect 297 274 343 498
rect 457 274 503 498
rect 617 274 663 498
rect -663 -112 -617 112
rect -503 -112 -457 112
rect -343 -112 -297 112
rect -183 -112 -137 112
rect -23 -112 23 112
rect 137 -112 183 112
rect 297 -112 343 112
rect 457 -112 503 112
rect 617 -112 663 112
rect -663 -498 -617 -274
rect -503 -498 -457 -274
rect -343 -498 -297 -274
rect -183 -498 -137 -274
rect -23 -498 23 -274
rect 137 -498 183 -274
rect 297 -498 343 -274
rect 457 -498 503 -274
rect 617 -498 663 -274
<< polysilicon >>
rect -588 511 -532 555
rect -428 511 -372 555
rect -268 511 -212 555
rect -108 511 -52 555
rect 52 511 108 555
rect 212 511 268 555
rect 372 511 428 555
rect 532 511 588 555
rect -588 217 -532 261
rect -428 217 -372 261
rect -268 217 -212 261
rect -108 217 -52 261
rect 52 217 108 261
rect 212 217 268 261
rect 372 217 428 261
rect 532 217 588 261
rect -588 125 -532 169
rect -428 125 -372 169
rect -268 125 -212 169
rect -108 125 -52 169
rect 52 125 108 169
rect 212 125 268 169
rect 372 125 428 169
rect 532 125 588 169
rect -588 -169 -532 -125
rect -428 -169 -372 -125
rect -268 -169 -212 -125
rect -108 -169 -52 -125
rect 52 -169 108 -125
rect 212 -169 268 -125
rect 372 -169 428 -125
rect 532 -169 588 -125
rect -588 -261 -532 -217
rect -428 -261 -372 -217
rect -268 -261 -212 -217
rect -108 -261 -52 -217
rect 52 -261 108 -217
rect 212 -261 268 -217
rect 372 -261 428 -217
rect 532 -261 588 -217
rect -588 -555 -532 -511
rect -428 -555 -372 -511
rect -268 -555 -212 -511
rect -108 -555 -52 -511
rect 52 -555 108 -511
rect 212 -555 268 -511
rect 372 -555 428 -511
rect 532 -555 588 -511
<< metal1 >>
rect -663 498 -617 509
rect -663 263 -617 274
rect -503 498 -457 509
rect -503 263 -457 274
rect -343 498 -297 509
rect -343 263 -297 274
rect -183 498 -137 509
rect -183 263 -137 274
rect -23 498 23 509
rect -23 263 23 274
rect 137 498 183 509
rect 137 263 183 274
rect 297 498 343 509
rect 297 263 343 274
rect 457 498 503 509
rect 457 263 503 274
rect 617 498 663 509
rect 617 263 663 274
rect -663 112 -617 123
rect -663 -123 -617 -112
rect -503 112 -457 123
rect -503 -123 -457 -112
rect -343 112 -297 123
rect -343 -123 -297 -112
rect -183 112 -137 123
rect -183 -123 -137 -112
rect -23 112 23 123
rect -23 -123 23 -112
rect 137 112 183 123
rect 137 -123 183 -112
rect 297 112 343 123
rect 297 -123 343 -112
rect 457 112 503 123
rect 457 -123 503 -112
rect 617 112 663 123
rect 617 -123 663 -112
rect -663 -274 -617 -263
rect -663 -509 -617 -498
rect -503 -274 -457 -263
rect -503 -509 -457 -498
rect -343 -274 -297 -263
rect -343 -509 -297 -498
rect -183 -274 -137 -263
rect -183 -509 -137 -498
rect -23 -274 23 -263
rect -23 -509 23 -498
rect 137 -274 183 -263
rect 137 -509 183 -498
rect 297 -274 343 -263
rect 297 -509 343 -498
rect 457 -274 503 -263
rect 457 -509 503 -498
rect 617 -274 663 -263
rect 617 -509 663 -498
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1.25 l 0.280 m 3 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
