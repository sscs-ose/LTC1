magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1175 1045 1175
<< metal1 >>
rect -45 169 45 175
rect -45 -169 -39 169
rect 39 -169 45 169
rect -45 -175 45 -169
<< via1 >>
rect -39 -169 39 169
<< metal2 >>
rect -45 169 45 175
rect -45 -169 -39 169
rect 39 -169 45 169
rect -45 -175 45 -169
<< end >>
