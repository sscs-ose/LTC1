* NGSPICE file created from CLK_div_4_mag_flat.ext - technology: gf180mcuC

.subckt CLK_div_4_mag_flat VDD VSS RST CLK Vdiv4
X0 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t47 VDD.t46 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_1.CLK VSS.t57 VSS.t56 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X2 a_4018_1378# VDD.t100 VSS.t44 VSS.t43 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X3 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_2_mag_1.JK_FF_mag_0.QB a_4178_1378# VSS.t4 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X4 CLK_div_2_mag_0.JK_FF_mag_0.QB CLK_div_2_mag_1.CLK a_2776_324# VSS.t55 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X5 a_4896_281# CLK_div_2_mag_1.RST a_4736_281# VSS.t6 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X6 VDD CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X7 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK.t0 VSS.t25 VSS.t24 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X8 a_4178_1378# CLK_div_2_mag_1.CLK a_4018_1378# VSS.t54 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X9 VDD CLK_div_2_mag_1.RST CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t13 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X10 CLK_div_2_mag_1.JK_FF_mag_0.QB CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t53 VDD.t52 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 a_764_280# VDD.t101 VSS.t42 VSS.t41 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X12 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_2_mag_0.JK_FF_mag_0.QB VDD.t3 VDD.t2 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 VDD CLK_div_2_mag_0.JK_FF_mag_0.QB CLK_div_2_mag_1.CLK VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X14 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t72 VDD.t71 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT Vdiv4.t3 a_4172_281# VSS.t2 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X16 VDD CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t28 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X17 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_4896_281# VSS.t28 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X18 a_4742_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t51 VSS.t50 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X19 Vdiv4 CLK_div_2_mag_1.JK_FF_mag_0.QB a_5870_1422# VSS.t3 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X20 a_924_280# CLK.t1 a_764_280# VSS.t7 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X21 a_1488_280# CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t9 VSS.t8 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X22 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_5306_1422# VSS.t23 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X23 a_5870_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t11 VSS.t10 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X24 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t51 VDD.t50 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X25 VDD Vdiv4.t4 CLK_div_2_mag_1.JK_FF_mag_0.QB VDD.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X26 a_6024_325# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t33 VSS.t32 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X27 VDD CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t25 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X28 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t58 VDD.t57 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X29 a_1648_280# CLK_div_2_mag_1.RST a_1488_280# VSS.t5 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X30 CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t24 VDD.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 VDD CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t54 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X32 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_1.CLK VDD.t99 VDD.t98 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2212_324# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X34 VDD CLK.t2 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t84 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t78 VDD.t77 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X36 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_1.CLK VDD.t97 VDD.t96 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_2_mag_0.JK_FF_mag_0.QB a_930_1377# VSS.t1 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X38 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t68 VDD.t70 VDD.t69 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X39 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK.t3 VDD.t49 VDD.t48 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X40 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t65 VDD.t67 VDD.t66 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X41 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t76 VDD.t75 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X42 CLK_div_2_mag_1.JK_FF_mag_0.QB Vdiv4.t5 a_6024_325# VSS.t29 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X43 a_5306_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t27 VSS.t26 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X44 VDD CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t41 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X45 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_1494_1421# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X46 a_4736_281# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t31 VSS.t30 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X47 a_5460_325# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t36 VSS.t35 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X48 a_1494_1421# CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t46 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X49 CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.QB a_2622_1421# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X50 VDD CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t93 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X51 CLK_div_2_mag_0.JK_FF_mag_0.QB CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t37 VDD.t36 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X52 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t62 VDD.t64 VDD.t63 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X53 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_2_mag_1.JK_FF_mag_0.QB VDD.t9 VDD.t8 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X54 VDD CLK_div_2_mag_1.JK_FF_mag_0.QB Vdiv4.t1 VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X55 VDD CLK_div_2_mag_1.RST CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t10 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X56 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t80 VDD.t79 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X57 VDD CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X58 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t59 VDD.t61 VDD.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X59 VDD CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X60 Vdiv4 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X61 a_930_1377# CLK.t4 a_770_1377# VSS.t14 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X62 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t32 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X63 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_1.CLK a_924_280# VSS.t53 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X64 a_770_1377# VDD.t102 VSS.t40 VSS.t39 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X65 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT Vdiv4.t6 VDD.t74 VDD.t73 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X66 a_4012_281# VDD.t103 VSS.t38 VSS.t37 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X67 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_5460_325# VSS.t22 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X68 VDD CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.QB VDD.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X69 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_1648_280# VSS.t49 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X70 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t20 VDD.t19 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X71 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t45 VDD.t44 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X72 a_2776_324# CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t21 VSS.t20 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X73 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2058_1421# VSS.t15 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X74 a_2622_1421# CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t13 VSS.t12 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X75 VDD CLK.t5 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X76 a_2058_1421# CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t48 VSS.t47 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X77 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_4742_1422# VSS.t34 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X78 a_2212_324# CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X79 a_4172_281# CLK_div_2_mag_1.CLK a_4012_281# VSS.t52 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
R0 VDD.t25 VDD.t23 961.905
R1 VDD.t2 VDD.t71 961.905
R2 VDD.t38 VDD.t21 765.152
R3 VDD.t46 VDD.t54 765.152
R4 VDD.t8 VDD.t79 765.152
R5 VDD.t28 VDD.t36 765.152
R6 VDD.t75 VDD.t31 765.152
R7 VDD.t98 VDD.t19 765.152
R8 VDD.t41 VDD.t52 765.152
R9 VDD.t44 VDD.t57 765.152
R10 VDD.t73 VDD.t50 765.152
R11 VDD.n79 VDD.t77 676.191
R12 VDD.n84 VDD.t66 485.714
R13 VDD VDD.n47 429.187
R14 VDD.t48 VDD.n84 426.44
R15 VDD.t84 VDD.t2 380.952
R16 VDD.t90 VDD.t8 303.031
R17 VDD.t13 VDD.t75 303.031
R18 VDD.t81 VDD.t98 303.031
R19 VDD.t10 VDD.t44 303.031
R20 VDD.t93 VDD.t73 303.031
R21 VDD.t33 VDD.n79 285.714
R22 VDD.n75 VDD.t0 242.857
R23 VDD.n77 VDD.t25 242.857
R24 VDD.n80 VDD.t33 242.857
R25 VDD.n83 VDD.t84 242.857
R26 VDD.n33 VDD.t5 193.183
R27 VDD.n34 VDD.t38 193.183
R28 VDD.n43 VDD.t54 193.183
R29 VDD.n44 VDD.t90 193.183
R30 VDD.n49 VDD.t87 193.183
R31 VDD.n51 VDD.t28 193.183
R32 VDD.n54 VDD.t13 193.183
R33 VDD.n57 VDD.t81 193.183
R34 VDD.n3 VDD.t16 193.183
R35 VDD.n5 VDD.t41 193.183
R36 VDD.n8 VDD.t10 193.183
R37 VDD.n11 VDD.t93 193.183
R38 VDD.t23 VDD.n75 138.095
R39 VDD.t77 VDD.n77 138.095
R40 VDD.t71 VDD.n80 138.095
R41 VDD.t66 VDD.n83 138.095
R42 VDD.t21 VDD.n33 109.849
R43 VDD.n34 VDD.t46 109.849
R44 VDD.t79 VDD.n43 109.849
R45 VDD.n44 VDD.t63 109.849
R46 VDD.t36 VDD.n49 109.849
R47 VDD.t31 VDD.n51 109.849
R48 VDD.t19 VDD.n54 109.849
R49 VDD.n57 VDD.t60 109.849
R50 VDD.t52 VDD.n3 109.849
R51 VDD.t57 VDD.n5 109.849
R52 VDD.t50 VDD.n8 109.849
R53 VDD.n11 VDD.t69 109.849
R54 VDD.n47 VDD.t96 59.702
R55 VDD.n58 VDD.t65 30.9379
R56 VDD.n60 VDD.t59 30.9379
R57 VDD.n12 VDD.t62 30.9379
R58 VDD.n14 VDD.t68 30.9379
R59 VDD.n58 VDD.t102 24.5101
R60 VDD.n60 VDD.t101 24.5101
R61 VDD.n12 VDD.t100 24.5101
R62 VDD.n14 VDD.t103 24.5101
R63 VDD VDD.t48 10.5649
R64 VDD.n63 VDD.n57 6.3005
R65 VDD.n66 VDD.n54 6.3005
R66 VDD.n69 VDD.n51 6.3005
R67 VDD.n72 VDD.n49 6.3005
R68 VDD.n86 VDD.n83 6.3005
R69 VDD.n89 VDD.n80 6.3005
R70 VDD.n92 VDD.n77 6.3005
R71 VDD.n95 VDD.n75 6.3005
R72 VDD.n17 VDD.n11 6.3005
R73 VDD.n20 VDD.n8 6.3005
R74 VDD.n23 VDD.n5 6.3005
R75 VDD.n26 VDD.n3 6.3005
R76 VDD.n33 VDD.n32 6.3005
R77 VDD.n35 VDD.n34 6.3005
R78 VDD.n43 VDD.n42 6.3005
R79 VDD.n45 VDD.n44 6.3005
R80 VDD.n62 VDD.t61 5.13287
R81 VDD.n65 VDD.t20 5.13287
R82 VDD.n68 VDD.t32 5.13287
R83 VDD.n70 VDD.n50 5.13287
R84 VDD.n71 VDD.t37 5.13287
R85 VDD.n73 VDD.n48 5.13287
R86 VDD.n16 VDD.t70 5.13287
R87 VDD.n19 VDD.t51 5.13287
R88 VDD.n22 VDD.t58 5.13287
R89 VDD.n24 VDD.n4 5.13287
R90 VDD.n25 VDD.t53 5.13287
R91 VDD.n27 VDD.n2 5.13287
R92 VDD VDD.t49 5.13124
R93 VDD.n85 VDD.t67 5.11708
R94 VDD.n88 VDD.t72 5.11708
R95 VDD.n90 VDD.n78 5.11708
R96 VDD.n91 VDD.t78 5.11708
R97 VDD.n93 VDD.n76 5.11708
R98 VDD.n94 VDD.t24 5.11708
R99 VDD.n96 VDD.n74 5.11708
R100 VDD.n46 VDD.t64 5.11708
R101 VDD.n41 VDD.t80 5.11708
R102 VDD.n37 VDD.n0 5.11708
R103 VDD.n36 VDD.t47 5.11708
R104 VDD.n30 VDD.n29 5.11708
R105 VDD.n31 VDD.t22 5.11708
R106 VDD.n28 VDD.n1 5.11708
R107 VDD.n98 VDD.t97 5.09407
R108 VDD VDD.n60 4.08487
R109 VDD VDD.n14 4.08487
R110 VDD.n59 VDD.n58 4.07684
R111 VDD.n13 VDD.n12 4.07684
R112 VDD.n61 VDD.n59 3.00126
R113 VDD.n15 VDD.n13 3.00126
R114 VDD.n61 VDD 2.87711
R115 VDD.n15 VDD 2.87711
R116 VDD.n64 VDD.n56 2.85787
R117 VDD.n67 VDD.n53 2.85787
R118 VDD.n18 VDD.n10 2.85787
R119 VDD.n21 VDD.n7 2.85787
R120 VDD.n87 VDD.n82 2.84208
R121 VDD.n40 VDD.n39 2.84208
R122 VDD.n62 VDD.n61 2.28069
R123 VDD.n16 VDD.n15 2.28069
R124 VDD.n82 VDD.t3 2.2755
R125 VDD.n82 VDD.n81 2.2755
R126 VDD.n56 VDD.t99 2.2755
R127 VDD.n56 VDD.n55 2.2755
R128 VDD.n53 VDD.t76 2.2755
R129 VDD.n53 VDD.n52 2.2755
R130 VDD.n39 VDD.t9 2.2755
R131 VDD.n39 VDD.n38 2.2755
R132 VDD.n10 VDD.t74 2.2755
R133 VDD.n10 VDD.n9 2.2755
R134 VDD.n7 VDD.t45 2.2755
R135 VDD.n7 VDD.n6 2.2755
R136 VDD.n28 VDD.n27 1.12142
R137 VDD.n97 VDD.n73 1.01882
R138 VDD.n68 VDD.n67 0.233919
R139 VDD.n65 VDD.n64 0.233919
R140 VDD.n22 VDD.n21 0.233919
R141 VDD.n19 VDD.n18 0.233919
R142 VDD.n98 VDD.n97 0.197054
R143 VDD VDD.n46 0.1472
R144 VDD.n85 VDD 0.14647
R145 VDD.n71 VDD.n70 0.141016
R146 VDD.n25 VDD.n24 0.141016
R147 VDD.n31 VDD.n30 0.1094
R148 VDD.n37 VDD.n36 0.1094
R149 VDD.n94 VDD.n93 0.108858
R150 VDD.n91 VDD.n90 0.108858
R151 VDD.n73 VDD.n72 0.107339
R152 VDD.n70 VDD.n69 0.107339
R153 VDD.n27 VDD.n26 0.107339
R154 VDD.n24 VDD.n23 0.107339
R155 VDD.n67 VDD 0.106177
R156 VDD.n64 VDD 0.106177
R157 VDD.n21 VDD 0.106177
R158 VDD.n18 VDD 0.106177
R159 VDD.n97 VDD.n96 0.10259
R160 VDD VDD.n40 0.0869
R161 VDD VDD.n87 0.0864701
R162 VDD.n32 VDD.n28 0.0833
R163 VDD.n42 VDD.n37 0.0833
R164 VDD.n96 VDD.n95 0.0828881
R165 VDD.n93 VDD.n92 0.0828881
R166 VDD.n90 VDD.n89 0.0828881
R167 VDD.n40 VDD 0.0824
R168 VDD.n87 VDD 0.0819925
R169 VDD.n66 VDD.n65 0.080629
R170 VDD.n63 VDD.n62 0.080629
R171 VDD.n20 VDD.n19 0.080629
R172 VDD.n17 VDD.n16 0.080629
R173 VDD VDD.n71 0.0794677
R174 VDD VDD.n68 0.0794677
R175 VDD VDD.n25 0.0794677
R176 VDD VDD.n22 0.0794677
R177 VDD.n46 VDD.n45 0.0626
R178 VDD.n86 VDD.n85 0.062291
R179 VDD VDD.n31 0.0617
R180 VDD.n36 VDD 0.0617
R181 VDD VDD.n41 0.0617
R182 VDD VDD.n94 0.0613955
R183 VDD VDD.n91 0.0613955
R184 VDD VDD.n88 0.0613955
R185 VDD.n35 VDD 0.0455
R186 VDD.n41 VDD 0.0455
R187 VDD.n88 VDD 0.0452761
R188 VDD.n30 VDD 0.0383
R189 VDD VDD.n98 0.03785
R190 VDD.n59 VDD 0.003875
R191 VDD.n13 VDD 0.003875
R192 VDD.n72 VDD 0.00166129
R193 VDD.n69 VDD 0.00166129
R194 VDD VDD.n66 0.00166129
R195 VDD VDD.n63 0.00166129
R196 VDD.n26 VDD 0.00166129
R197 VDD.n23 VDD 0.00166129
R198 VDD VDD.n20 0.00166129
R199 VDD VDD.n17 0.00166129
R200 VDD.n32 VDD 0.0014
R201 VDD VDD.n35 0.0014
R202 VDD.n42 VDD 0.0014
R203 VDD.n45 VDD 0.0014
R204 VDD.n95 VDD 0.00139552
R205 VDD.n92 VDD 0.00139552
R206 VDD.n89 VDD 0.00139552
R207 VDD VDD.n86 0.00139552
R208 VSS.t29 VSS.n1 9492.76
R209 VSS.t56 VSS.n29 4221.41
R210 VSS.t10 VSS.t23 2307.56
R211 VSS.t34 VSS.t26 2307.56
R212 VSS.t50 VSS.t4 2307.56
R213 VSS.t12 VSS.t15 2307.56
R214 VSS.t19 VSS.t47 2307.56
R215 VSS.t45 VSS.t1 2307.56
R216 VSS.n33 VSS.t37 2171.54
R217 VSS.n33 VSS.t55 2166.53
R218 VSS.t16 VSS.t20 2097.44
R219 VSS.t53 VSS.t8 2097.44
R220 VSS.t22 VSS.t32 2094.1
R221 VSS.t2 VSS.t30 2094.1
R222 VSS.n34 VSS.n33 1991.72
R223 VSS.n32 VSS.t43 1199.47
R224 VSS.n46 VSS.t39 1199.47
R225 VSS.t0 VSS.n34 1153.78
R226 VSS.t4 VSS.t54 913.885
R227 VSS.t1 VSS.t14 913.885
R228 VSS.n47 VSS.t24 874.567
R229 VSS.t5 VSS.t49 830.672
R230 VSS.t7 VSS.t53 830.672
R231 VSS.t6 VSS.t28 829.346
R232 VSS.t52 VSS.t2 829.346
R233 VSS.n31 VSS.t56 611.347
R234 VSS.n17 VSS.t3 548.331
R235 VSS.n22 VSS.t23 548.331
R236 VSS.n23 VSS.t34 548.331
R237 VSS.n28 VSS.t54 548.331
R238 VSS.n35 VSS.t0 548.331
R239 VSS.n40 VSS.t15 548.331
R240 VSS.n41 VSS.t19 548.331
R241 VSS.n45 VSS.t14 548.331
R242 VSS.t55 VSS.n12 498.404
R243 VSS.n13 VSS.t16 498.404
R244 VSS.n14 VSS.t5 498.404
R245 VSS.n15 VSS.t7 498.404
R246 VSS.n4 VSS.t29 497.608
R247 VSS.n5 VSS.t22 497.608
R248 VSS.n9 VSS.t6 497.608
R249 VSS.n10 VSS.t52 497.608
R250 VSS.n17 VSS.t10 365.555
R251 VSS.t26 VSS.n22 365.555
R252 VSS.n23 VSS.t50 365.555
R253 VSS.t43 VSS.n28 365.555
R254 VSS.n35 VSS.t12 365.555
R255 VSS.t47 VSS.n40 365.555
R256 VSS.n41 VSS.t45 365.555
R257 VSS.t39 VSS.n45 365.555
R258 VSS.t20 VSS.n12 332.269
R259 VSS.n13 VSS.t17 332.269
R260 VSS.t8 VSS.n14 332.269
R261 VSS.n15 VSS.t41 332.269
R262 VSS.t32 VSS.n4 331.738
R263 VSS.n5 VSS.t35 331.738
R264 VSS.t30 VSS.n9 331.738
R265 VSS.t37 VSS.n10 331.738
R266 VSS.n47 VSS.n46 28.2123
R267 VSS.n32 VSS.n31 19.7214
R268 VSS.n30 VSS.t57 9.3736
R269 VSS.n48 VSS.t25 9.3736
R270 VSS.n2 VSS.t33 7.19156
R271 VSS.n7 VSS.t36 7.19156
R272 VSS.n19 VSS.t11 7.19156
R273 VSS.n20 VSS.t27 7.19156
R274 VSS.n25 VSS.t51 7.19156
R275 VSS.n37 VSS.t13 7.19156
R276 VSS.n38 VSS.t48 7.19156
R277 VSS.n43 VSS.t46 7.19156
R278 VSS.n56 VSS.t21 7.18989
R279 VSS.n54 VSS.t18 7.18989
R280 VSS.n0 VSS.t31 5.91399
R281 VSS.n59 VSS.t38 5.91399
R282 VSS.n26 VSS.t44 5.91399
R283 VSS.n16 VSS.t40 5.91399
R284 VSS.n52 VSS.t9 5.91232
R285 VSS.n50 VSS.t42 5.91232
R286 VSS.n48 VSS.n47 5.2005
R287 VSS.n18 VSS.n17 5.2005
R288 VSS.n22 VSS.n21 5.2005
R289 VSS.n24 VSS.n23 5.2005
R290 VSS.n28 VSS.n27 5.2005
R291 VSS.n31 VSS.n30 5.2005
R292 VSS.n45 VSS.n44 5.2005
R293 VSS.n42 VSS.n41 5.2005
R294 VSS.n40 VSS.n39 5.2005
R295 VSS.n36 VSS.n35 5.2005
R296 VSS.n60 VSS.n10 5.2005
R297 VSS.n9 VSS.n8 5.2005
R298 VSS.n6 VSS.n5 5.2005
R299 VSS.n4 VSS.n3 5.2005
R300 VSS.n57 VSS.n12 5.2005
R301 VSS.n55 VSS.n13 5.2005
R302 VSS.n53 VSS.n14 5.2005
R303 VSS.n51 VSS.n15 5.2005
R304 VSS.n34 VSS.n32 3.94467
R305 VSS.n50 VSS.n49 0.941004
R306 VSS.n58 VSS.n11 0.845914
R307 VSS VSS.n19 0.343161
R308 VSS.n20 VSS 0.343161
R309 VSS VSS.n37 0.343161
R310 VSS.n38 VSS 0.343161
R311 VSS.n27 VSS 0.289491
R312 VSS.n44 VSS 0.289491
R313 VSS.n8 VSS.n7 0.245993
R314 VSS.n54 VSS.n53 0.245993
R315 VSS VSS.n25 0.191234
R316 VSS VSS.n43 0.191234
R317 VSS.n2 VSS 0.175852
R318 VSS.n56 VSS 0.175852
R319 VSS.n58 VSS 0.153458
R320 VSS VSS.n60 0.140359
R321 VSS VSS.n51 0.140359
R322 VSS VSS.n11 0.137685
R323 VSS.n49 VSS 0.137685
R324 VSS.n19 VSS.n18 0.118573
R325 VSS.n21 VSS.n20 0.118573
R326 VSS.n25 VSS.n24 0.118573
R327 VSS.n37 VSS.n36 0.118573
R328 VSS.n39 VSS.n38 0.118573
R329 VSS.n43 VSS.n42 0.118573
R330 VSS VSS.n26 0.115271
R331 VSS VSS.n16 0.115271
R332 VSS VSS.n0 0.106134
R333 VSS.n52 VSS 0.106134
R334 VSS.n26 VSS.n11 0.10206
R335 VSS.n49 VSS.n16 0.10206
R336 VSS.n59 VSS.n58 0.0964155
R337 VSS.n3 VSS.n2 0.0609225
R338 VSS.n7 VSS.n6 0.0609225
R339 VSS.n57 VSS.n56 0.0609225
R340 VSS.n55 VSS.n54 0.0609225
R341 VSS VSS.n0 0.0592324
R342 VSS VSS.n59 0.0592324
R343 VSS VSS.n52 0.0592324
R344 VSS VSS.n50 0.0592324
R345 VSS.n18 VSS 0.00545413
R346 VSS.n21 VSS 0.00545413
R347 VSS.n24 VSS 0.00545413
R348 VSS.n36 VSS 0.00545413
R349 VSS.n39 VSS 0.00545413
R350 VSS.n42 VSS 0.00545413
R351 VSS.n27 VSS 0.00380275
R352 VSS.n44 VSS 0.00380275
R353 VSS.n3 VSS 0.00303521
R354 VSS.n6 VSS 0.00303521
R355 VSS VSS.n57 0.00303521
R356 VSS VSS.n55 0.00303521
R357 VSS.n30 VSS 0.00219811
R358 VSS VSS.n48 0.00219811
R359 VSS.n8 VSS 0.00219014
R360 VSS.n60 VSS 0.00219014
R361 VSS.n53 VSS 0.00219014
R362 VSS.n51 VSS 0.00219014
R363 CLK.n9 CLK.t4 36.935
R364 CLK.n3 CLK.t1 36.935
R365 CLK.n14 CLK.t3 25.5361
R366 CLK.n9 CLK.t2 18.1962
R367 CLK.n3 CLK.t5 18.1962
R368 CLK.n14 CLK.t0 14.0734
R369 CLK.n5 CLK.n2 4.5005
R370 CLK.n5 CLK.n4 4.5005
R371 CLK.n8 CLK.n7 4.5005
R372 CLK.n10 CLK.n7 4.5005
R373 CLK.n16 CLK.n15 4.5005
R374 CLK.n17 CLK.n16 4.5005
R375 CLK.n12 CLK.n11 2.25107
R376 CLK.n13 CLK.n0 2.24235
R377 CLK.n4 CLK.n3 2.12175
R378 CLK.n10 CLK.n9 2.12075
R379 CLK.n7 CLK.n6 1.74297
R380 CLK.n6 CLK.n1 1.49778
R381 CLK.n15 CLK.n14 1.42775
R382 CLK.n13 CLK.n12 0.97145
R383 CLK CLK.n17 0.1605
R384 CLK.n8 CLK 0.0473512
R385 CLK.n2 CLK 0.0473512
R386 CLK.n11 CLK.n8 0.0361897
R387 CLK.n2 CLK.n1 0.0361897
R388 CLK.n17 CLK.n0 0.03175
R389 CLK.n16 CLK.n13 0.0246174
R390 CLK.n6 CLK.n5 0.0131772
R391 CLK.n12 CLK.n7 0.0122182
R392 CLK.n11 CLK.n10 0.00515517
R393 CLK.n4 CLK.n1 0.00515517
R394 CLK.n15 CLK.n0 0.00175
R395 Vdiv4.n5 Vdiv4.t3 36.935
R396 Vdiv4.n7 Vdiv4.t5 31.528
R397 Vdiv4.n5 Vdiv4.t6 18.1962
R398 Vdiv4.n7 Vdiv4.t4 15.3826
R399 Vdiv4.n3 Vdiv4.n0 7.09905
R400 Vdiv4.n8 Vdiv4.n7 6.86134
R401 Vdiv4.n9 Vdiv4.n6 5.01116
R402 Vdiv4.n3 Vdiv4.n2 3.25085
R403 Vdiv4.n10 Vdiv4.n4 2.33232
R404 Vdiv4.n2 Vdiv4.t1 2.2755
R405 Vdiv4.n2 Vdiv4.n1 2.2755
R406 Vdiv4.n6 Vdiv4.n5 2.13398
R407 Vdiv4.n10 Vdiv4.n9 1.35708
R408 Vdiv4.n9 Vdiv4.n8 1.12056
R409 Vdiv4 Vdiv4.n10 0.41675
R410 Vdiv4.n4 Vdiv4.n3 0.0919062
R411 Vdiv4.n8 Vdiv4 0.0857632
R412 Vdiv4.n6 Vdiv4 0.0810725
R413 Vdiv4.n4 Vdiv4 0.073625
C0 CLK_div_2_mag_1.CLK a_4012_281# 0.00165f
C1 a_5870_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C2 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C3 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_2058_1421# 4.52e-20
C4 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2212_324# 0.0036f
C5 CLK_div_2_mag_1.RST CLK_div_2_mag_0.JK_FF_mag_0.QB 0.204f
C6 a_4018_1378# VDD 0.00492f
C7 a_2622_1421# CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00372f
C8 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_924_280# 1.46e-19
C9 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_2776_324# 0.00372f
C10 CLK_div_2_mag_1.CLK a_1648_280# 0.0101f
C11 CLK_div_2_mag_1.CLK VDD 2.25f
C12 a_924_280# CLK 0.00164f
C13 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C14 a_770_1377# CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C15 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C16 VDD CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.23f
C17 CLK_div_2_mag_1.RST CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0816f
C18 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_4178_1378# 0.0732f
C19 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_764_280# 1.17e-20
C20 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_1.JK_FF_mag_0.QB 0.103f
C21 m2_175_583# CLK 6.19e-19
C22 RST VDD 0.00299f
C23 a_5870_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00372f
C24 a_5460_325# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C25 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT Vdiv4 0.0343f
C26 VDD m1_3423_584# 0.00266f
C27 a_2622_1421# CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C28 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_0.JK_FF_mag_0.QB 0.103f
C29 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C30 CLK_div_2_mag_1.CLK a_2058_1421# 3.95e-21
C31 a_4172_281# a_4012_281# 0.0504f
C32 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_1494_1421# 0.0697f
C33 CLK_div_2_mag_1.JK_FF_mag_0.QB a_4178_1378# 0.00392f
C34 a_4742_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C35 VDD CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.402f
C36 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.22f
C37 a_4736_281# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C38 a_5306_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C39 a_2212_324# CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C40 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_1.JK_FF_mag_0.QB 0.199f
C41 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C42 a_1488_280# a_1648_280# 0.0504f
C43 VDD a_2776_324# 3.14e-19
C44 a_6024_325# CLK_div_2_mag_1.JK_FF_mag_0.QB 0.0811f
C45 a_1488_280# VDD 2.21e-19
C46 VDD CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.758f
C47 a_770_1377# a_930_1377# 0.0504f
C48 CLK_div_2_mag_1.CLK Vdiv4 0.157f
C49 CLK_div_2_mag_1.CLK a_764_280# 0.00335f
C50 VDD CLK 1.06f
C51 a_5870_1422# CLK_div_2_mag_1.JK_FF_mag_0.QB 0.0114f
C52 VDD CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.402f
C53 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C54 Vdiv4 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0168f
C55 VDD m2_3423_584# 0.0206f
C56 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_4012_281# 0.0202f
C57 CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 9.71e-20
C58 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.RST 0.278f
C59 CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C60 a_770_1377# CLK 0.0101f
C61 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2058_1421# 0.011f
C62 VDD CLK_div_2_mag_1.JK_FF_mag_0.QB 0.908f
C63 CLK_div_2_mag_1.RST a_1494_1421# 3.11e-19
C64 a_5306_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C65 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD 0.747f
C66 a_2622_1421# VDD 3.6e-19
C67 CLK_div_2_mag_1.RST a_4742_1422# 3.11e-19
C68 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C69 a_4896_281# Vdiv4 0.0101f
C70 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 9.85e-22
C71 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_6024_325# 0.00372f
C72 CLK_div_2_mag_1.RST CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.253f
C73 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 Vdiv4 0.107f
C74 a_5460_325# CLK_div_2_mag_1.JK_FF_mag_0.QB 0.00964f
C75 a_2058_1421# CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C76 VDD CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C77 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_5870_1422# 4.52e-20
C78 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.QB 0.25f
C79 a_2212_324# VDD 3.14e-19
C80 a_4172_281# Vdiv4 0.00789f
C81 CLK_div_2_mag_0.JK_FF_mag_0.QB a_1494_1421# 3e-19
C82 Vdiv4 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C83 CLK_div_2_mag_1.RST CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00531f
C84 a_4896_281# a_4736_281# 0.0504f
C85 m2_175_583# VDD 0.0195f
C86 a_764_280# CLK 0.00117f
C87 a_4896_281# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C88 CLK_div_2_mag_1.RST a_4018_1378# 9.23e-19
C89 a_5306_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C90 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C91 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C92 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C93 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C94 CLK_div_2_mag_1.RST CLK_div_2_mag_1.CLK 0.164f
C95 a_6024_325# VDD 3.14e-19
C96 CLK_div_2_mag_0.JK_FF_mag_0.QB CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C97 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C98 CLK_div_2_mag_1.RST CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00463f
C99 a_5870_1422# VDD 3.6e-19
C100 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_5460_325# 0.069f
C101 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK 9.71e-20
C102 Vdiv4 CLK_div_2_mag_1.JK_FF_mag_0.QB 1.94f
C103 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT Vdiv4 0.338f
C104 a_4018_1378# CLK_div_2_mag_0.JK_FF_mag_0.QB 1.23e-20
C105 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C106 VDD a_4012_281# 0.00108f
C107 CLK_div_2_mag_1.RST RST 0.00399f
C108 CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.QB 1.96f
C109 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C110 CLK_div_2_mag_1.RST m1_3423_584# 0.00362f
C111 CLK_div_2_mag_1.RST a_930_1377# 7.69e-19
C112 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.QB 2.24e-19
C113 a_4736_281# CLK_div_2_mag_1.JK_FF_mag_0.QB 0.00695f
C114 a_5306_1422# CLK_div_2_mag_1.JK_FF_mag_0.QB 2.96e-19
C115 a_4736_281# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C116 CLK_div_2_mag_1.RST a_4896_281# 0.00153f
C117 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_1.JK_FF_mag_0.QB 0.0386f
C118 a_764_280# a_924_280# 0.0504f
C119 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.00165f
C120 CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C121 Vdiv4 a_4178_1378# 2.79e-20
C122 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_1.RST 0.0673f
C123 a_5460_325# VDD 3.14e-19
C124 CLK_div_2_mag_1.RST a_4172_281# 0.00188f
C125 CLK_div_2_mag_0.JK_FF_mag_0.QB m1_3423_584# 0.00478f
C126 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 Vdiv4 0.0635f
C127 CLK_div_2_mag_1.RST a_2776_324# 9.78e-19
C128 CLK_div_2_mag_1.RST a_1488_280# 0.0017f
C129 CLK_div_2_mag_1.RST CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00531f
C130 CLK_div_2_mag_0.JK_FF_mag_0.QB a_930_1377# 0.00392f
C131 VDD a_770_1377# 0.00492f
C132 a_6024_325# Vdiv4 0.0157f
C133 CLK_div_2_mag_1.RST CLK 0.0415f
C134 CLK_div_2_mag_1.RST CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00428f
C135 a_5870_1422# Vdiv4 0.069f
C136 VDD a_2058_1421# 3.18e-19
C137 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.QB 0.28f
C138 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_1494_1421# 0.0202f
C139 CLK_div_2_mag_1.RST m2_3423_584# 0.0408f
C140 Vdiv4 a_4012_281# 0.00335f
C141 CLK_div_2_mag_0.JK_FF_mag_0.QB a_2776_324# 0.0811f
C142 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_2_mag_0.JK_FF_mag_0.QB 2.97e-21
C143 a_1488_280# CLK_div_2_mag_0.JK_FF_mag_0.QB 0.00695f
C144 CLK_div_2_mag_0.JK_FF_mag_0.QB CLK 0.307f
C145 CLK_div_2_mag_1.RST CLK_div_2_mag_1.JK_FF_mag_0.QB 0.0996f
C146 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_0.JK_FF_mag_0.QB 0.0592f
C147 CLK_div_2_mag_1.RST CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0816f
C148 VDD Vdiv4 1.07f
C149 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00118f
C150 CLK_div_2_mag_1.RST a_2622_1421# 6.04e-19
C151 a_764_280# VDD 0.00108f
C152 a_4742_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C153 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_1488_280# 9.1e-19
C154 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C155 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK 0.235f
C156 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_1494_1421# 0.00378f
C157 a_5460_325# Vdiv4 0.00859f
C158 CLK_div_2_mag_1.RST CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0192f
C159 CLK_div_2_mag_1.RST a_2212_324# 9.57e-19
C160 CLK_div_2_mag_1.RST a_924_280# 0.00188f
C161 a_4736_281# VDD 2.21e-19
C162 a_5306_1422# VDD 3.18e-19
C163 a_2622_1421# CLK_div_2_mag_0.JK_FF_mag_0.QB 0.0114f
C164 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_1648_280# 8.64e-19
C165 VDD CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.656f
C166 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.CLK 0.0343f
C167 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.656f
C168 CLK_div_2_mag_1.RST m2_175_583# 0.0301f
C169 CLK_div_2_mag_1.RST a_4178_1378# 7.69e-19
C170 CLK_div_2_mag_1.CLK a_4742_1422# 6.43e-21
C171 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_1.RST 2.17e-19
C172 CLK_div_2_mag_0.JK_FF_mag_0.QB CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.199f
C173 a_2212_324# CLK_div_2_mag_0.JK_FF_mag_0.QB 0.00964f
C174 CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 6.64e-19
C175 a_4742_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C176 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C177 CLK_div_2_mag_0.JK_FF_mag_0.QB a_4178_1378# 9.82e-21
C178 CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C179 CLK_div_2_mag_1.RST a_4012_281# 0.00188f
C180 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_924_280# 0.0731f
C181 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_2058_1421# 0.0059f
C182 CLK_div_2_mag_1.CLK a_4018_1378# 0.0101f
C183 CLK_div_2_mag_1.RST a_1648_280# 0.00187f
C184 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C185 CLK_div_2_mag_1.RST VDD 0.741f
C186 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_1494_1421# 1.43e-19
C187 a_4736_281# Vdiv4 0.0102f
C188 a_4896_281# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C189 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_1488_280# 0.0203f
C190 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 Vdiv4 0.00335f
C191 CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.417f
C192 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK 6.64e-19
C193 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_930_1377# 0.0732f
C194 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C195 CLK a_1494_1421# 6.43e-21
C196 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C197 a_4742_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C198 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_4172_281# 1.5e-20
C199 CLK_div_2_mag_0.JK_FF_mag_0.QB a_1648_280# 0.00696f
C200 VDD CLK_div_2_mag_0.JK_FF_mag_0.QB 0.911f
C201 CLK_div_2_mag_1.RST a_770_1377# 9.23e-19
C202 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C203 CLK_div_2_mag_1.CLK m1_3423_584# 0.00833f
C204 a_5306_1422# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C205 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0889f
C206 CLK_div_2_mag_1.CLK a_930_1377# 2.79e-20
C207 CLK_div_2_mag_1.RST a_2058_1421# 6.04e-19
C208 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_1648_280# 2.88e-20
C209 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK 0.267f
C210 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD 0.747f
C211 CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 1.48e-20
C212 a_4018_1378# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C213 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_1.CLK 0.0177f
C214 a_4742_1422# CLK_div_2_mag_1.JK_FF_mag_0.QB 3e-19
C215 CLK_div_2_mag_1.CLK a_4172_281# 0.00202f
C216 CLK_div_2_mag_1.CLK a_2776_324# 0.0157f
C217 CLK_div_2_mag_1.CLK a_1488_280# 0.0102f
C218 CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.267f
C219 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C220 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_1.JK_FF_mag_0.QB 0.25f
C221 CLK_div_2_mag_1.RST Vdiv4 0.0427f
C222 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C223 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00191f
C224 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C225 CLK_div_2_mag_1.CLK CLK 0.149f
C226 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_2212_324# 0.00378f
C227 CLK_div_2_mag_1.RST a_764_280# 0.00188f
C228 a_4172_281# CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C229 a_2058_1421# CLK_div_2_mag_0.JK_FF_mag_0.QB 2.96e-19
C230 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_924_280# 1.5e-20
C231 CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C232 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0889f
C233 CLK_div_2_mag_1.CLK m2_3423_584# 0.0133f
C234 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C235 CLK_div_2_mag_1.RST a_4736_281# 0.0017f
C236 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_930_1377# 0.00119f
C237 RST CLK 4.42e-19
C238 Vdiv4 CLK_div_2_mag_0.JK_FF_mag_0.QB 1.03e-19
C239 CLK_div_2_mag_1.RST CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.152f
C240 CLK_div_2_mag_1.RST CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.188f
C241 CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.QB 0.307f
C242 CLK_div_2_mag_1.CLK CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C243 CLK_div_2_mag_1.CLK a_2622_1421# 0.069f
C244 CLK a_930_1377# 0.00939f
C245 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C246 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_1.JK_FF_mag_0.QB 0.28f
C247 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C248 m2_3423_584# m1_3423_584# 0.021f
C249 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT a_764_280# 0.0202f
C250 CLK_div_2_mag_1.CLK CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C251 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK 0.42f
C252 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_2_mag_0.JK_FF_mag_0.QB 0.0386f
C253 CLK_div_2_mag_1.CLK a_2212_324# 0.00859f
C254 CLK_div_2_mag_1.CLK a_924_280# 0.00789f
C255 a_4018_1378# a_4178_1378# 0.0504f
C256 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C257 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_1648_280# 0.0733f
C258 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.995f
C259 CLK_div_2_mag_1.CLK a_4178_1378# 0.00939f
C260 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_4012_281# 1.17e-20
C261 VDD a_1494_1421# 3.18e-19
C262 a_4896_281# CLK_div_2_mag_1.JK_FF_mag_0.QB 0.00696f
C263 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK 1.48e-20
C264 a_4742_1422# VDD 3.18e-19
C265 a_4896_281# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C266 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00165f
C267 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 a_4178_1378# 0.00119f
C268 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_2_mag_1.JK_FF_mag_0.QB 0.0592f
C269 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.995f
C270 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C271 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_2622_1421# 0.00118f
C272 m2_175_583# RST 0.0331f
C273 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_4172_281# 0.0731f
C274 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_2_mag_1.JK_FF_mag_0.QB 0.343f
C275 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C276 VDD CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.758f
C277 a_5460_325# CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C278 RST VSS 0.234f
C279 m2_3423_584# VSS 0.0503f $ **FLOATING
C280 m2_175_583# VSS 0.0631f $ **FLOATING
C281 m1_3423_584# VSS 0.139f $ **FLOATING
C282 a_6024_325# VSS 0.0675f
C283 a_5460_325# VSS 0.0676f
C284 a_4896_281# VSS 0.0343f
C285 a_4736_281# VSS 0.0881f
C286 a_4172_281# VSS 0.0343f
C287 a_4012_281# VSS 0.0881f
C288 a_2776_324# VSS 0.0676f
C289 a_2212_324# VSS 0.0677f
C290 a_1648_280# VSS 0.0345f
C291 a_1488_280# VSS 0.0883f
C292 a_924_280# VSS 0.0345f
C293 a_764_280# VSS 0.0883f
C294 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C295 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.54f
C296 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.416f
C297 CLK_div_2_mag_1.RST VSS 1.57f
C298 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.541f
C299 a_5870_1422# VSS 0.0676f
C300 a_5306_1422# VSS 0.0676f
C301 a_4742_1422# VSS 0.0676f
C302 a_4178_1378# VSS 0.0343f
C303 a_4018_1378# VSS 0.0881f
C304 a_2622_1421# VSS 0.0676f
C305 a_2058_1421# VSS 0.0676f
C306 a_1494_1421# VSS 0.0676f
C307 a_930_1377# VSS 0.0343f
C308 a_770_1377# VSS 0.0881f
C309 Vdiv4 VSS 1.64f
C310 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C311 CLK_div_2_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.934f
C312 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C313 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.81f
C314 CLK_div_2_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C315 CLK_div_2_mag_1.JK_FF_mag_0.QB VSS 0.918f
C316 CLK_div_2_mag_1.CLK VSS 2.39f
C317 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C318 CLK_div_2_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.936f
C319 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C320 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C321 CLK_div_2_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C322 CLK_div_2_mag_0.JK_FF_mag_0.QB VSS 0.897f
C323 CLK VSS 0.98f
C324 VDD VSS 27f
C325 VDD.t64 VSS 0.00225f
C326 VDD.t54 VSS 0.0298f
C327 VDD.n0 VSS 0.00225f
C328 VDD.t47 VSS 0.00225f
C329 VDD.t5 VSS 0.0294f
C330 VDD.n1 VSS 0.00225f
C331 VDD.n2 VSS 0.00226f
C332 VDD.t16 VSS 0.0294f
C333 VDD.n3 VSS 0.014f
C334 VDD.t53 VSS 0.00226f
C335 VDD.n4 VSS 0.00226f
C336 VDD.t52 VSS 0.0272f
C337 VDD.t41 VSS 0.0298f
C338 VDD.n5 VSS 0.014f
C339 VDD.t58 VSS 0.00226f
C340 VDD.t45 VSS 9.29e-19
C341 VDD.n6 VSS 9.29e-19
C342 VDD.n7 VSS 0.00203f
C343 VDD.t57 VSS 0.0272f
C344 VDD.t44 VSS 0.0332f
C345 VDD.t10 VSS 0.0154f
C346 VDD.n8 VSS 0.014f
C347 VDD.t51 VSS 0.00226f
C348 VDD.t74 VSS 9.29e-19
C349 VDD.n9 VSS 9.29e-19
C350 VDD.n10 VSS 0.00203f
C351 VDD.t50 VSS 0.0272f
C352 VDD.t73 VSS 0.0332f
C353 VDD.t93 VSS 0.0154f
C354 VDD.t69 VSS 0.0272f
C355 VDD.n11 VSS 0.014f
C356 VDD.t70 VSS 0.00226f
C357 VDD.t62 VSS 0.00194f
C358 VDD.t100 VSS 0.00147f
C359 VDD.n12 VSS 0.00381f
C360 VDD.n13 VSS 0.00367f
C361 VDD.t68 VSS 0.00194f
C362 VDD.t103 VSS 0.00147f
C363 VDD.n14 VSS 0.00381f
C364 VDD.n15 VSS 0.0171f
C365 VDD.n16 VSS 0.0105f
C366 VDD.n17 VSS 0.00701f
C367 VDD.n18 VSS 0.0129f
C368 VDD.n19 VSS 0.0132f
C369 VDD.n20 VSS 0.00701f
C370 VDD.n21 VSS 0.0129f
C371 VDD.n22 VSS 0.0132f
C372 VDD.n23 VSS 0.0078f
C373 VDD.n24 VSS 0.0112f
C374 VDD.n25 VSS 0.0104f
C375 VDD.n26 VSS 0.0078f
C376 VDD.n27 VSS 0.021f
C377 VDD.n28 VSS 0.0278f
C378 VDD.t22 VSS 0.00225f
C379 VDD.n29 VSS 0.00225f
C380 VDD.n30 VSS 0.011f
C381 VDD.n31 VSS 0.0122f
C382 VDD.n32 VSS 0.00874f
C383 VDD.n33 VSS 0.014f
C384 VDD.t21 VSS 0.0272f
C385 VDD.t38 VSS 0.0298f
C386 VDD.t46 VSS 0.0272f
C387 VDD.n34 VSS 0.014f
C388 VDD.n35 VSS 0.00686f
C389 VDD.n36 VSS 0.0122f
C390 VDD.n37 VSS 0.0132f
C391 VDD.t80 VSS 0.00225f
C392 VDD.t9 VSS 9.29e-19
C393 VDD.n38 VSS 9.29e-19
C394 VDD.n39 VSS 0.00201f
C395 VDD.n40 VSS 0.011f
C396 VDD.n41 VSS 0.00901f
C397 VDD.n42 VSS 0.00874f
C398 VDD.n43 VSS 0.014f
C399 VDD.t79 VSS 0.0272f
C400 VDD.t8 VSS 0.0332f
C401 VDD.t90 VSS 0.0154f
C402 VDD.t63 VSS 0.0154f
C403 VDD.n44 VSS 0.014f
C404 VDD.n45 VSS 0.00771f
C405 VDD.n46 VSS 0.0141f
C406 VDD.t96 VSS 0.0199f
C407 VDD.n47 VSS 0.021f
C408 VDD.t97 VSS 0.00225f
C409 VDD.n48 VSS 0.00226f
C410 VDD.t87 VSS 0.0294f
C411 VDD.n49 VSS 0.014f
C412 VDD.t37 VSS 0.00226f
C413 VDD.n50 VSS 0.00226f
C414 VDD.t36 VSS 0.0272f
C415 VDD.t28 VSS 0.0298f
C416 VDD.n51 VSS 0.014f
C417 VDD.t32 VSS 0.00226f
C418 VDD.t76 VSS 9.29e-19
C419 VDD.n52 VSS 9.29e-19
C420 VDD.n53 VSS 0.00203f
C421 VDD.t31 VSS 0.0272f
C422 VDD.t75 VSS 0.0332f
C423 VDD.t13 VSS 0.0154f
C424 VDD.n54 VSS 0.014f
C425 VDD.t20 VSS 0.00226f
C426 VDD.t99 VSS 9.29e-19
C427 VDD.n55 VSS 9.29e-19
C428 VDD.n56 VSS 0.00203f
C429 VDD.t19 VSS 0.0272f
C430 VDD.t98 VSS 0.0332f
C431 VDD.t81 VSS 0.0154f
C432 VDD.t60 VSS 0.0272f
C433 VDD.n57 VSS 0.014f
C434 VDD.t61 VSS 0.00226f
C435 VDD.t65 VSS 0.00194f
C436 VDD.t102 VSS 0.00147f
C437 VDD.n58 VSS 0.00381f
C438 VDD.n59 VSS 0.00367f
C439 VDD.t59 VSS 0.00194f
C440 VDD.t101 VSS 0.00147f
C441 VDD.n60 VSS 0.00381f
C442 VDD.n61 VSS 0.0171f
C443 VDD.n62 VSS 0.0105f
C444 VDD.n63 VSS 0.00701f
C445 VDD.n64 VSS 0.0129f
C446 VDD.n65 VSS 0.0132f
C447 VDD.n66 VSS 0.00701f
C448 VDD.n67 VSS 0.0129f
C449 VDD.n68 VSS 0.0132f
C450 VDD.n69 VSS 0.0078f
C451 VDD.n70 VSS 0.0112f
C452 VDD.n71 VSS 0.0104f
C453 VDD.n72 VSS 0.0078f
C454 VDD.n73 VSS 0.0195f
C455 VDD.n74 VSS 0.00225f
C456 VDD.t0 VSS 0.0237f
C457 VDD.n75 VSS 0.0121f
C458 VDD.t24 VSS 0.00225f
C459 VDD.n76 VSS 0.00225f
C460 VDD.t23 VSS 0.0217f
C461 VDD.t25 VSS 0.0237f
C462 VDD.n77 VSS 0.0121f
C463 VDD.t78 VSS 0.00225f
C464 VDD.n78 VSS 0.00225f
C465 VDD.t77 VSS 0.016f
C466 VDD.n79 VSS 0.0626f
C467 VDD.t33 VSS 0.0104f
C468 VDD.n80 VSS 0.0121f
C469 VDD.t72 VSS 0.00225f
C470 VDD.t3 VSS 9.29e-19
C471 VDD.n81 VSS 9.29e-19
C472 VDD.n82 VSS 0.00201f
C473 VDD.t71 VSS 0.0217f
C474 VDD.t2 VSS 0.0264f
C475 VDD.t84 VSS 0.0123f
C476 VDD.n83 VSS 0.0121f
C477 VDD.t67 VSS 0.00225f
C478 VDD.t66 VSS 0.0123f
C479 VDD.n84 VSS 0.0346f
C480 VDD.t48 VSS 0.0249f
C481 VDD.t49 VSS 0.00233f
C482 VDD.n85 VSS 0.0142f
C483 VDD.n86 VSS 0.00773f
C484 VDD.n87 VSS 0.011f
C485 VDD.n88 VSS 0.00904f
C486 VDD.n89 VSS 0.00876f
C487 VDD.n90 VSS 0.0133f
C488 VDD.n91 VSS 0.0122f
C489 VDD.n92 VSS 0.00876f
C490 VDD.n93 VSS 0.0133f
C491 VDD.n94 VSS 0.0122f
C492 VDD.n95 VSS 0.00876f
C493 VDD.n96 VSS 0.0129f
C494 VDD.n97 VSS 0.0243f
C495 VDD.n98 VSS 0.0158f
.ends

