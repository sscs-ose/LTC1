* NGSPICE file created from nand2_flat.ext - technology: gf180mcuC

.subckt nand2_flat VDD IN2 IN1 OUT VSS
X0 OUT IN2.t0 a_168_68# VSS.t2 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X1 OUT IN1.t0 VDD.t4 VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X2 a_168_68# IN1.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3 VDD IN2.t1 OUT.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
R0 IN2.n0 IN2.t0 31.528
R1 IN2.n0 IN2.t1 15.3826
R2 IN2 IN2.n0 8.86438
R3 OUT.n3 OUT.n2 7.16286
R4 OUT.n3 OUT.n1 3.21288
R5 OUT.n1 OUT.t1 2.2755
R6 OUT.n1 OUT.n0 2.2755
R7 OUT OUT.n3 0.0103182
R8 VSS.n0 VSS.t2 596.558
R9 VSS.n0 VSS.t0 397.707
R10 VSS VSS.t1 7.30881
R11 VSS VSS.n2 2.60133
R12 VSS.n2 VSS.n0 2.6005
R13 VSS.n2 VSS.n1 0.0904743
R14 IN1.n0 IN1.t0 30.9379
R15 IN1.n0 IN1.t1 21.6422
R16 IN1 IN1.n0 4.1052
R17 VDD.n1 VDD.t0 193.183
R18 VDD.n1 VDD.t3 109.849
R19 VDD.n2 VDD.n1 6.3005
R20 VDD VDD.n0 5.23506
R21 VDD.n2 VDD.t4 5.213
R22 VDD VDD.n2 0.00514516
C0 IN2 IN1 0.0466f
C1 VDD IN2 0.225f
C2 OUT IN1 0.0929f
C3 VDD OUT 0.201f
C4 VDD IN1 0.158f
C5 a_168_68# IN2 0.00348f
C6 a_168_68# OUT 0.069f
C7 a_168_68# IN1 0.00347f
C8 a_168_68# VDD 3.14e-19
C9 OUT IN2 0.191f
.ends

