magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 3032 71968
<< psubdiff >>
rect 0 69778 1000 69968
rect 0 13287 93 69778
rect 907 13287 1000 69778
rect 0 13097 1000 13287
<< metal1 >>
rect -32 69789 1032 69957
rect -32 13276 14 69789
rect 986 13276 1032 69789
rect -32 13108 1032 13276
<< metal2 >>
rect 56 65000 178 69660
rect 0 63600 178 65000
rect 56 50600 178 63600
rect 0 49200 178 50600
rect 56 13491 178 49200
rect 280 23600 356 68189
rect 656 14000 732 69589
rect 839 65000 915 69660
rect 839 63600 1000 65000
rect 839 50600 915 63600
rect 839 49200 1000 50600
rect 839 13494 915 49200
<< metal3 >>
rect 0 68400 1000 69678
rect 0 66800 1000 68200
rect 0 65200 1000 66600
rect 0 63600 1000 65000
rect 0 62000 1000 63400
rect 0 60400 1000 61800
rect 0 58800 1000 60200
rect 0 57200 1000 58600
rect 0 55600 1000 57000
rect 0 54000 1000 55400
rect 0 52400 1000 53800
rect 0 50800 1000 52200
rect 0 49200 1000 50600
rect 0 46000 1000 49000
rect 0 42800 1000 45800
rect 0 41200 1000 42600
rect 0 39600 1000 41000
rect 0 36400 1000 39400
rect 0 33200 1000 36200
rect 0 30000 1000 33000
rect 0 26800 1000 29800
rect 0 25200 1000 26600
rect 0 23600 1000 25000
rect 0 20400 1000 23400
rect 0 17200 1000 20200
rect 0 14000 1000 17000
use M1_PSUB_CDNS_690335831656  M1_PSUB_CDNS_690335831656_0
timestamp 1713338890
transform 1 0 952 0 1 41524
box -45 -28395 45 28395
use M1_PSUB_CDNS_690335831656  M1_PSUB_CDNS_690335831656_1
timestamp 1713338890
transform -1 0 48 0 1 41524
box -45 -28395 45 28395
use M1_PSUB_CDNS_6903358316578  M1_PSUB_CDNS_6903358316578_0
timestamp 1713338890
transform 1 0 500 0 -1 13192
box -345 -95 345 95
use M1_PSUB_CDNS_6903358316578  M1_PSUB_CDNS_6903358316578_1
timestamp 1713338890
transform 1 0 500 0 1 69873
box -345 -95 345 95
use M2_M1_CDNS_6903358316577  M2_M1_CDNS_6903358316577_0
timestamp 1713338890
transform 1 0 85 0 1 49900
box -38 -596 38 596
use M2_M1_CDNS_6903358316577  M2_M1_CDNS_6903358316577_1
timestamp 1713338890
transform 1 0 877 0 1 49900
box -38 -596 38 596
use M2_M1_CDNS_6903358316577  M2_M1_CDNS_6903358316577_2
timestamp 1713338890
transform 1 0 877 0 1 64300
box -38 -596 38 596
use M2_M1_CDNS_6903358316577  M2_M1_CDNS_6903358316577_3
timestamp 1713338890
transform 1 0 85 0 1 64300
box -38 -596 38 596
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_0
timestamp 1713338890
transform 1 0 694 0 1 15496
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_1
timestamp 1713338890
transform 1 0 694 0 1 18696
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_2
timestamp 1713338890
transform 1 0 694 0 1 21908
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_3
timestamp 1713338890
transform 1 0 318 0 1 28343
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_4
timestamp 1713338890
transform 1 0 318 0 1 31513
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_5
timestamp 1713338890
transform 1 0 318 0 1 34718
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_6
timestamp 1713338890
transform 1 0 318 0 1 37888
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_7
timestamp 1713338890
transform 1 0 318 0 1 44311
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316566  M3_M2_CDNS_6903358316566_8
timestamp 1713338890
transform 1 0 694 0 1 47528
box -38 -1292 38 1292
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_0
timestamp 1713338890
transform 1 0 318 0 1 24298
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_1
timestamp 1713338890
transform 1 0 694 0 1 25929
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_2
timestamp 1713338890
transform 1 0 318 0 1 41895
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_3
timestamp 1713338890
transform 1 0 694 0 1 40327
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_4
timestamp 1713338890
transform 1 0 510 0 1 51504
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_5
timestamp 1713338890
transform 1 0 318 0 1 53113
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_6
timestamp 1713338890
transform 1 0 318 0 1 54704
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_7
timestamp 1713338890
transform 1 0 318 0 1 56323
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_8
timestamp 1713338890
transform 1 0 318 0 1 59505
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_9
timestamp 1713338890
transform 1 0 694 0 1 57897
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_10
timestamp 1713338890
transform 1 0 694 0 1 61108
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_11
timestamp 1713338890
transform 1 0 510 0 1 62697
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_12
timestamp 1713338890
transform 1 0 318 0 1 67494
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_13
timestamp 1713338890
transform 1 0 694 0 1 65910
box -38 -566 38 566
use M3_M2_CDNS_6903358316567  M3_M2_CDNS_6903358316567_14
timestamp 1713338890
transform 1 0 694 0 1 69023
box -38 -566 38 566
use M3_M2_CDNS_6903358316576  M3_M2_CDNS_6903358316576_0
timestamp 1713338890
transform 1 0 85 0 1 49900
box -38 -596 38 596
use M3_M2_CDNS_6903358316576  M3_M2_CDNS_6903358316576_1
timestamp 1713338890
transform 1 0 877 0 1 49900
box -38 -596 38 596
use M3_M2_CDNS_6903358316576  M3_M2_CDNS_6903358316576_2
timestamp 1713338890
transform 1 0 877 0 1 64300
box -38 -596 38 596
use M3_M2_CDNS_6903358316576  M3_M2_CDNS_6903358316576_3
timestamp 1713338890
transform 1 0 85 0 1 64300
box -38 -596 38 596
use POLY_SUB_FILL  POLY_SUB_FILL_0
array 0 0 0 0 34 1600
timestamp 1713338890
transform 1 0 -806 0 1 13819
box 880 -349 1727 1343
<< labels >>
rlabel metal3 s 487 67458 487 67458 4 DVDD
port 1 nsew
rlabel metal3 s 487 59623 487 59623 4 DVDD
port 1 nsew
rlabel metal3 s 487 56423 487 56423 4 DVDD
port 1 nsew
rlabel metal3 s 487 54658 487 54658 4 DVDD
port 1 nsew
rlabel metal3 s 487 53223 487 53223 4 DVDD
port 1 nsew
rlabel metal3 s 487 44368 487 44368 4 DVDD
port 1 nsew
rlabel metal3 s 487 41977 487 41977 4 DVDD
port 1 nsew
rlabel metal3 s 487 37959 487 37959 4 DVDD
port 1 nsew
rlabel metal3 s 487 34723 487 34723 4 DVDD
port 1 nsew
rlabel metal3 s 487 31609 487 31609 4 DVDD
port 1 nsew
rlabel metal3 s 487 28394 487 28394 4 DVDD
port 1 nsew
rlabel metal3 s 487 24284 487 24284 4 DVDD
port 1 nsew
rlabel metal3 s 487 18921 487 18921 4 DVSS
port 2 nsew
rlabel metal3 s 487 15750 487 15750 4 DVSS
port 2 nsew
rlabel metal3 s 487 21907 487 21907 4 DVSS
port 2 nsew
rlabel metal3 s 487 26100 487 26100 4 DVSS
port 2 nsew
rlabel metal3 s 487 40342 487 40342 4 DVSS
port 2 nsew
rlabel metal3 s 487 47595 487 47595 4 DVSS
port 2 nsew
rlabel metal3 s 487 57858 487 57858 4 DVSS
port 2 nsew
rlabel metal3 s 487 61058 487 61058 4 DVSS
port 2 nsew
rlabel metal3 s 487 66023 487 66023 4 DVSS
port 2 nsew
rlabel metal3 s 487 69049 487 69049 4 DVSS
port 2 nsew
rlabel metal3 s 487 51458 487 51458 4 VDD
port 3 nsew
rlabel metal3 s 487 62823 487 62823 4 VDD
port 3 nsew
rlabel metal3 s 487 64258 487 64258 4 VSS
port 4 nsew
rlabel metal3 s 487 50023 487 50023 4 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1000 70000
<< end >>
