magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1046 -1775 1046 1775
<< metal1 >>
rect -46 769 46 775
rect -46 743 -40 769
rect -14 743 14 769
rect 40 743 46 769
rect -46 715 46 743
rect -46 689 -40 715
rect -14 689 14 715
rect 40 689 46 715
rect -46 661 46 689
rect -46 635 -40 661
rect -14 635 14 661
rect 40 635 46 661
rect -46 607 46 635
rect -46 581 -40 607
rect -14 581 14 607
rect 40 581 46 607
rect -46 553 46 581
rect -46 527 -40 553
rect -14 527 14 553
rect 40 527 46 553
rect -46 499 46 527
rect -46 473 -40 499
rect -14 473 14 499
rect 40 473 46 499
rect -46 445 46 473
rect -46 419 -40 445
rect -14 419 14 445
rect 40 419 46 445
rect -46 391 46 419
rect -46 365 -40 391
rect -14 365 14 391
rect 40 365 46 391
rect -46 337 46 365
rect -46 311 -40 337
rect -14 311 14 337
rect 40 311 46 337
rect -46 283 46 311
rect -46 257 -40 283
rect -14 257 14 283
rect 40 257 46 283
rect -46 229 46 257
rect -46 203 -40 229
rect -14 203 14 229
rect 40 203 46 229
rect -46 175 46 203
rect -46 149 -40 175
rect -14 149 14 175
rect 40 149 46 175
rect -46 121 46 149
rect -46 95 -40 121
rect -14 95 14 121
rect 40 95 46 121
rect -46 67 46 95
rect -46 41 -40 67
rect -14 41 14 67
rect 40 41 46 67
rect -46 13 46 41
rect -46 -13 -40 13
rect -14 -13 14 13
rect 40 -13 46 13
rect -46 -41 46 -13
rect -46 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 46 -41
rect -46 -95 46 -67
rect -46 -121 -40 -95
rect -14 -121 14 -95
rect 40 -121 46 -95
rect -46 -149 46 -121
rect -46 -175 -40 -149
rect -14 -175 14 -149
rect 40 -175 46 -149
rect -46 -203 46 -175
rect -46 -229 -40 -203
rect -14 -229 14 -203
rect 40 -229 46 -203
rect -46 -257 46 -229
rect -46 -283 -40 -257
rect -14 -283 14 -257
rect 40 -283 46 -257
rect -46 -311 46 -283
rect -46 -337 -40 -311
rect -14 -337 14 -311
rect 40 -337 46 -311
rect -46 -365 46 -337
rect -46 -391 -40 -365
rect -14 -391 14 -365
rect 40 -391 46 -365
rect -46 -419 46 -391
rect -46 -445 -40 -419
rect -14 -445 14 -419
rect 40 -445 46 -419
rect -46 -473 46 -445
rect -46 -499 -40 -473
rect -14 -499 14 -473
rect 40 -499 46 -473
rect -46 -527 46 -499
rect -46 -553 -40 -527
rect -14 -553 14 -527
rect 40 -553 46 -527
rect -46 -581 46 -553
rect -46 -607 -40 -581
rect -14 -607 14 -581
rect 40 -607 46 -581
rect -46 -635 46 -607
rect -46 -661 -40 -635
rect -14 -661 14 -635
rect 40 -661 46 -635
rect -46 -689 46 -661
rect -46 -715 -40 -689
rect -14 -715 14 -689
rect 40 -715 46 -689
rect -46 -743 46 -715
rect -46 -769 -40 -743
rect -14 -769 14 -743
rect 40 -769 46 -743
rect -46 -775 46 -769
<< via1 >>
rect -40 743 -14 769
rect 14 743 40 769
rect -40 689 -14 715
rect 14 689 40 715
rect -40 635 -14 661
rect 14 635 40 661
rect -40 581 -14 607
rect 14 581 40 607
rect -40 527 -14 553
rect 14 527 40 553
rect -40 473 -14 499
rect 14 473 40 499
rect -40 419 -14 445
rect 14 419 40 445
rect -40 365 -14 391
rect 14 365 40 391
rect -40 311 -14 337
rect 14 311 40 337
rect -40 257 -14 283
rect 14 257 40 283
rect -40 203 -14 229
rect 14 203 40 229
rect -40 149 -14 175
rect 14 149 40 175
rect -40 95 -14 121
rect 14 95 40 121
rect -40 41 -14 67
rect 14 41 40 67
rect -40 -13 -14 13
rect 14 -13 40 13
rect -40 -67 -14 -41
rect 14 -67 40 -41
rect -40 -121 -14 -95
rect 14 -121 40 -95
rect -40 -175 -14 -149
rect 14 -175 40 -149
rect -40 -229 -14 -203
rect 14 -229 40 -203
rect -40 -283 -14 -257
rect 14 -283 40 -257
rect -40 -337 -14 -311
rect 14 -337 40 -311
rect -40 -391 -14 -365
rect 14 -391 40 -365
rect -40 -445 -14 -419
rect 14 -445 40 -419
rect -40 -499 -14 -473
rect 14 -499 40 -473
rect -40 -553 -14 -527
rect 14 -553 40 -527
rect -40 -607 -14 -581
rect 14 -607 40 -581
rect -40 -661 -14 -635
rect 14 -661 40 -635
rect -40 -715 -14 -689
rect 14 -715 40 -689
rect -40 -769 -14 -743
rect 14 -769 40 -743
<< metal2 >>
rect -46 769 46 775
rect -46 743 -40 769
rect -14 743 14 769
rect 40 743 46 769
rect -46 715 46 743
rect -46 689 -40 715
rect -14 689 14 715
rect 40 689 46 715
rect -46 661 46 689
rect -46 635 -40 661
rect -14 635 14 661
rect 40 635 46 661
rect -46 607 46 635
rect -46 581 -40 607
rect -14 581 14 607
rect 40 581 46 607
rect -46 553 46 581
rect -46 527 -40 553
rect -14 527 14 553
rect 40 527 46 553
rect -46 499 46 527
rect -46 473 -40 499
rect -14 473 14 499
rect 40 473 46 499
rect -46 445 46 473
rect -46 419 -40 445
rect -14 419 14 445
rect 40 419 46 445
rect -46 391 46 419
rect -46 365 -40 391
rect -14 365 14 391
rect 40 365 46 391
rect -46 337 46 365
rect -46 311 -40 337
rect -14 311 14 337
rect 40 311 46 337
rect -46 283 46 311
rect -46 257 -40 283
rect -14 257 14 283
rect 40 257 46 283
rect -46 229 46 257
rect -46 203 -40 229
rect -14 203 14 229
rect 40 203 46 229
rect -46 175 46 203
rect -46 149 -40 175
rect -14 149 14 175
rect 40 149 46 175
rect -46 121 46 149
rect -46 95 -40 121
rect -14 95 14 121
rect 40 95 46 121
rect -46 67 46 95
rect -46 41 -40 67
rect -14 41 14 67
rect 40 41 46 67
rect -46 13 46 41
rect -46 -13 -40 13
rect -14 -13 14 13
rect 40 -13 46 13
rect -46 -41 46 -13
rect -46 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 46 -41
rect -46 -95 46 -67
rect -46 -121 -40 -95
rect -14 -121 14 -95
rect 40 -121 46 -95
rect -46 -149 46 -121
rect -46 -175 -40 -149
rect -14 -175 14 -149
rect 40 -175 46 -149
rect -46 -203 46 -175
rect -46 -229 -40 -203
rect -14 -229 14 -203
rect 40 -229 46 -203
rect -46 -257 46 -229
rect -46 -283 -40 -257
rect -14 -283 14 -257
rect 40 -283 46 -257
rect -46 -311 46 -283
rect -46 -337 -40 -311
rect -14 -337 14 -311
rect 40 -337 46 -311
rect -46 -365 46 -337
rect -46 -391 -40 -365
rect -14 -391 14 -365
rect 40 -391 46 -365
rect -46 -419 46 -391
rect -46 -445 -40 -419
rect -14 -445 14 -419
rect 40 -445 46 -419
rect -46 -473 46 -445
rect -46 -499 -40 -473
rect -14 -499 14 -473
rect 40 -499 46 -473
rect -46 -527 46 -499
rect -46 -553 -40 -527
rect -14 -553 14 -527
rect 40 -553 46 -527
rect -46 -581 46 -553
rect -46 -607 -40 -581
rect -14 -607 14 -581
rect 40 -607 46 -581
rect -46 -635 46 -607
rect -46 -661 -40 -635
rect -14 -661 14 -635
rect 40 -661 46 -635
rect -46 -689 46 -661
rect -46 -715 -40 -689
rect -14 -715 14 -689
rect 40 -715 46 -689
rect -46 -743 46 -715
rect -46 -769 -40 -743
rect -14 -769 14 -743
rect 40 -769 46 -743
rect -46 -775 46 -769
<< end >>
