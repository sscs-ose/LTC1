magic
tech gf180mcuC
magscale 1 10
timestamp 1691396512
<< pwell >>
rect -460 -736 460 736
<< nmos >>
rect -348 68 -292 668
rect -188 68 -132 668
rect -28 68 28 668
rect 132 68 188 668
rect 292 68 348 668
rect -348 -668 -292 -68
rect -188 -668 -132 -68
rect -28 -668 28 -68
rect 132 -668 188 -68
rect 292 -668 348 -68
<< ndiff >>
rect -436 655 -348 668
rect -436 81 -423 655
rect -377 81 -348 655
rect -436 68 -348 81
rect -292 655 -188 668
rect -292 81 -263 655
rect -217 81 -188 655
rect -292 68 -188 81
rect -132 655 -28 668
rect -132 81 -103 655
rect -57 81 -28 655
rect -132 68 -28 81
rect 28 655 132 668
rect 28 81 57 655
rect 103 81 132 655
rect 28 68 132 81
rect 188 655 292 668
rect 188 81 217 655
rect 263 81 292 655
rect 188 68 292 81
rect 348 655 436 668
rect 348 81 377 655
rect 423 81 436 655
rect 348 68 436 81
rect -436 -81 -348 -68
rect -436 -655 -423 -81
rect -377 -655 -348 -81
rect -436 -668 -348 -655
rect -292 -81 -188 -68
rect -292 -655 -263 -81
rect -217 -655 -188 -81
rect -292 -668 -188 -655
rect -132 -81 -28 -68
rect -132 -655 -103 -81
rect -57 -655 -28 -81
rect -132 -668 -28 -655
rect 28 -81 132 -68
rect 28 -655 57 -81
rect 103 -655 132 -81
rect 28 -668 132 -655
rect 188 -81 292 -68
rect 188 -655 217 -81
rect 263 -655 292 -81
rect 188 -668 292 -655
rect 348 -81 436 -68
rect 348 -655 377 -81
rect 423 -655 436 -81
rect 348 -668 436 -655
<< ndiffc >>
rect -423 81 -377 655
rect -263 81 -217 655
rect -103 81 -57 655
rect 57 81 103 655
rect 217 81 263 655
rect 377 81 423 655
rect -423 -655 -377 -81
rect -263 -655 -217 -81
rect -103 -655 -57 -81
rect 57 -655 103 -81
rect 217 -655 263 -81
rect 377 -655 423 -81
<< polysilicon >>
rect -348 668 -292 712
rect -188 668 -132 712
rect -28 668 28 712
rect 132 668 188 712
rect 292 668 348 712
rect -348 24 -292 68
rect -188 24 -132 68
rect -28 24 28 68
rect 132 24 188 68
rect 292 24 348 68
rect -348 -68 -292 -24
rect -188 -68 -132 -24
rect -28 -68 28 -24
rect 132 -68 188 -24
rect 292 -68 348 -24
rect -348 -712 -292 -668
rect -188 -712 -132 -668
rect -28 -712 28 -668
rect 132 -712 188 -668
rect 292 -712 348 -668
<< metal1 >>
rect -423 655 -377 666
rect -423 70 -377 81
rect -263 655 -217 666
rect -263 70 -217 81
rect -103 655 -57 666
rect -103 70 -57 81
rect 57 655 103 666
rect 57 70 103 81
rect 217 655 263 666
rect 217 70 263 81
rect 377 655 423 666
rect 377 70 423 81
rect -423 -81 -377 -70
rect -423 -666 -377 -655
rect -263 -81 -217 -70
rect -263 -666 -217 -655
rect -103 -81 -57 -70
rect -103 -666 -57 -655
rect 57 -81 103 -70
rect 57 -666 103 -655
rect 217 -81 263 -70
rect 217 -666 263 -655
rect 377 -81 423 -70
rect 377 -666 423 -655
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 2 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
