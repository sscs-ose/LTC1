** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/pex_LSBs_magic_TG_TB.sch
**.subckt pex_LSBs_magic_TG_TB
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
V6 B4 VSS pulse(0 3.3 0 10p 10p 400n 800n)
.save i(v6)
V7 B5 VSS pulse(0 3.3 0 10p 10p 800n 1.6u)
.save i(v7)
V8 B6 VSS pulse(0 3.3 0 10p 10p 1.6u 3.2u)
.save i(v8)
V10 B3 VSS pulse(0 3.3 0 10p 10p 200n 400n)
.save i(v10)
V11 B2 VSS pulse(0 3.3 0 10p 10p 100n 200n)
.save i(v11)
V12 B1 VSS pulse(0 3.3 0 10p 10p 50n 100n)
.save i(v12)
I0 VDD ITAIL 2.5u
R1 VDD OUT+ 5k m=1
R2 VDD OUT- 5k m=1
V9 SEL_L VSS 3.3
.save i(v9)
x1 VDD VSS B1 B2 B3 B4 B5 B6 ITAIL OUT+ OUT- net2 net3 net4 net5 net6 net7 SEL_L C32_D C32_U
+ pex_LSBs_magic_TG
XM1 V_ext C32_U net1 VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net1 C32_D VSS VSS nfet_03v3 L=0.5u W=19.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
R3 V_ext VDD 5k m=1
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_LSBs_magic_TG.spice
.option savecurrents
.control
save all
op

tran 10n 3.2u
plot v(OUT+) v(OUT-)
write pex_LSBs_magic_TG_TB.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
