magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -3133 -3188 4101 3774
<< nwell >>
rect -928 972 1872 1345
rect -460 903 4 972
rect 1593 882 1595 951
rect 178 607 273 610
rect 277 607 290 610
rect 197 558 199 607
rect 659 552 663 630
rect 1207 544 1212 628
rect 197 226 199 308
rect 646 303 663 307
rect 666 303 758 307
rect 178 -22 290 -21
rect 1207 -96 1212 -17
rect 1675 -97 1679 -22
rect -717 -102 -671 -101
<< pwell >>
rect -227 -516 1567 -507
rect -746 -564 1567 -516
rect -746 -908 1582 -564
<< psubdiff >>
rect -836 -1066 1675 -1044
rect -836 -1112 -803 -1066
rect -757 -1112 -603 -1066
rect -557 -1112 -403 -1066
rect -357 -1112 -203 -1066
rect -157 -1112 -3 -1066
rect 43 -1112 197 -1066
rect 243 -1112 397 -1066
rect 443 -1112 597 -1066
rect 643 -1112 797 -1066
rect 843 -1112 997 -1066
rect 1043 -1112 1197 -1066
rect 1243 -1112 1397 -1066
rect 1443 -1112 1597 -1066
rect 1643 -1112 1675 -1066
rect -836 -1134 1675 -1112
<< nsubdiff >>
rect -868 1290 -757 1292
rect -868 1270 1815 1290
rect -868 1224 -837 1270
rect -791 1268 1815 1270
rect -791 1224 -665 1268
rect -868 1222 -665 1224
rect -619 1222 -465 1268
rect -419 1222 -265 1268
rect -219 1222 -65 1268
rect -19 1222 135 1268
rect 181 1222 335 1268
rect 381 1222 535 1268
rect 581 1222 735 1268
rect 781 1222 935 1268
rect 981 1222 1135 1268
rect 1181 1222 1335 1268
rect 1381 1222 1535 1268
rect 1581 1222 1735 1268
rect 1781 1222 1815 1268
rect -868 1200 1815 1222
<< psubdiffcont >>
rect -803 -1112 -757 -1066
rect -603 -1112 -557 -1066
rect -403 -1112 -357 -1066
rect -203 -1112 -157 -1066
rect -3 -1112 43 -1066
rect 197 -1112 243 -1066
rect 397 -1112 443 -1066
rect 597 -1112 643 -1066
rect 797 -1112 843 -1066
rect 997 -1112 1043 -1066
rect 1197 -1112 1243 -1066
rect 1397 -1112 1443 -1066
rect 1597 -1112 1643 -1066
<< nsubdiffcont >>
rect -837 1224 -791 1270
rect -665 1222 -619 1268
rect -465 1222 -419 1268
rect -265 1222 -219 1268
rect -65 1222 -19 1268
rect 135 1222 181 1268
rect 335 1222 381 1268
rect 535 1222 581 1268
rect 735 1222 781 1268
rect 935 1222 981 1268
rect 1135 1222 1181 1268
rect 1335 1222 1381 1268
rect 1535 1222 1581 1268
rect 1735 1222 1781 1268
<< polysilicon >>
rect 646 943 758 963
rect -750 919 -637 934
rect -750 882 -717 919
rect -671 882 -637 919
rect 177 923 290 941
rect 177 882 218 923
rect 264 882 290 923
rect 646 897 682 943
rect 728 897 758 943
rect 646 882 758 897
rect 1114 940 1226 957
rect 1114 894 1145 940
rect 1191 894 1226 940
rect 1114 882 1226 894
rect 1582 937 1694 951
rect 1582 891 1612 937
rect 1658 891 1694 937
rect 1582 882 1694 891
rect -286 853 -174 868
rect -286 818 -259 853
rect -213 818 -174 853
rect 646 614 758 630
rect -750 593 -638 607
rect -750 558 -717 593
rect -671 558 -638 593
rect 178 596 290 610
rect -286 542 -174 590
rect 178 558 212 596
rect 258 558 290 596
rect 646 568 678 614
rect 724 568 758 614
rect 646 558 758 568
rect 1114 614 1226 631
rect 1114 568 1148 614
rect 1194 568 1226 614
rect 1114 558 1226 568
rect 1582 615 1694 629
rect 1582 569 1616 615
rect 1662 569 1694 615
rect 1582 558 1694 569
rect 659 552 663 558
rect 1207 544 1212 558
rect -750 270 -638 285
rect -750 234 -717 270
rect -671 234 -638 270
rect -286 266 -174 314
rect 178 291 290 308
rect 178 245 212 291
rect 258 245 290 291
rect 178 234 290 245
rect 646 291 758 307
rect 646 245 680 291
rect 726 245 758 291
rect 646 234 758 245
rect 1114 291 1226 309
rect 1114 245 1143 291
rect 1189 245 1226 291
rect 1114 234 1226 245
rect 1582 292 1694 306
rect 1582 246 1616 292
rect 1662 246 1694 292
rect 1582 234 1694 246
rect 178 233 273 234
rect 278 233 290 234
rect 191 226 199 233
rect 1675 227 1679 234
rect -286 -10 -174 38
rect -750 -55 -638 -29
rect -750 -90 -717 -55
rect -671 -90 -638 -55
rect 178 -35 290 -21
rect 178 -81 211 -35
rect 257 -81 290 -35
rect 178 -90 290 -81
rect 646 -35 758 -21
rect 646 -81 678 -35
rect 724 -81 758 -35
rect 646 -90 758 -81
rect 1114 -33 1226 -15
rect 1114 -79 1145 -33
rect 1191 -79 1226 -33
rect 1114 -90 1226 -79
rect 1582 -34 1694 -14
rect 1582 -80 1612 -34
rect 1658 -80 1694 -34
rect 1582 -90 1694 -80
rect 1207 -96 1212 -90
rect 1675 -97 1679 -90
rect -717 -102 -671 -101
rect -711 -134 -702 -102
rect -630 -503 -518 -475
rect -630 -544 -600 -503
rect -601 -549 -600 -544
rect -554 -544 -518 -503
rect -554 -549 -553 -544
rect -601 -551 -553 -549
rect 58 -679 282 -669
rect -278 -686 282 -679
rect -630 -736 -518 -688
rect -278 -732 206 -686
rect 252 -732 282 -686
rect -278 -735 282 -732
rect 394 -689 1084 -678
rect 394 -735 425 -689
rect 471 -734 1084 -689
rect 1324 -684 1436 -675
rect 1324 -730 1362 -684
rect 1408 -730 1436 -684
rect 1324 -731 1436 -730
rect 1358 -734 1412 -731
rect 471 -735 748 -734
rect 421 -739 475 -735
rect 505 -741 748 -735
<< polycontact >>
rect -717 873 -671 919
rect 218 877 264 923
rect 682 897 728 943
rect 1145 894 1191 940
rect 1612 891 1658 937
rect -259 807 -213 853
rect -717 547 -671 593
rect 212 550 258 596
rect 678 568 724 614
rect 1148 568 1194 614
rect 1616 569 1662 615
rect -717 224 -671 270
rect 212 245 258 291
rect 680 245 726 291
rect 1143 245 1189 291
rect 1616 246 1662 292
rect -717 -101 -671 -55
rect 211 -81 257 -35
rect 678 -81 724 -35
rect 1145 -79 1191 -33
rect 1612 -80 1658 -34
rect -600 -549 -554 -503
rect 206 -732 252 -686
rect 425 -735 471 -689
rect 1362 -730 1408 -684
<< metal1 >>
rect -61 1749 145 1774
rect -61 1697 78 1749
rect 130 1697 145 1749
rect -61 1676 145 1697
rect 54 1675 145 1676
rect -928 1270 1872 1345
rect -928 1224 -837 1270
rect -791 1268 1872 1270
rect -791 1224 -665 1268
rect -928 1222 -665 1224
rect -619 1222 -465 1268
rect -419 1222 -265 1268
rect -219 1222 -65 1268
rect -19 1222 135 1268
rect 181 1222 335 1268
rect 381 1222 535 1268
rect 581 1222 735 1268
rect 781 1222 935 1268
rect 981 1222 1135 1268
rect 1181 1222 1335 1268
rect 1381 1222 1535 1268
rect 1581 1222 1735 1268
rect 1781 1222 1872 1268
rect -928 1214 1872 1222
rect -928 1204 1736 1214
rect -928 1152 81 1204
rect 133 1162 1736 1204
rect 1788 1162 1872 1214
rect 133 1152 1872 1162
rect -928 1147 1872 1152
rect -840 -185 -772 1147
rect -724 919 -666 931
rect -724 873 -717 919
rect -671 873 -666 919
rect -724 593 -666 873
rect -494 926 -199 994
rect -724 547 -717 593
rect -671 547 -666 593
rect -724 270 -666 547
rect -724 224 -717 270
rect -671 224 -666 270
rect -724 -55 -666 224
rect -724 -101 -717 -55
rect -671 -101 -666 -55
rect -724 -307 -666 -101
rect -616 726 -548 833
rect -494 726 -426 926
rect -270 853 -199 926
rect -270 807 -259 853
rect -213 807 -199 853
rect -270 789 -199 807
rect -616 658 -426 726
rect -616 -138 -548 658
rect -616 -184 -439 -138
rect -616 -185 -614 -184
rect -724 -309 -541 -307
rect -881 -355 -541 -309
rect -612 -503 -541 -355
rect -612 -549 -600 -503
rect -554 -549 -541 -503
rect -612 -562 -541 -549
rect -899 -580 -809 -574
rect -1133 -599 -809 -580
rect -1133 -651 -879 -599
rect -827 -651 -809 -599
rect -1133 -664 -809 -651
rect -899 -673 -809 -664
rect -709 -990 -663 -576
rect -485 -831 -439 -184
rect -362 -304 -315 772
rect -145 -192 -99 1147
rect -23 1043 1906 1094
rect -23 838 28 1043
rect 199 937 275 950
rect 199 885 212 937
rect 199 877 218 885
rect 264 877 275 937
rect 667 946 746 960
rect 667 894 680 946
rect 732 894 746 946
rect 667 882 746 894
rect 199 876 275 877
rect 199 871 273 876
rect -23 787 161 838
rect 311 787 489 833
rect -23 185 28 787
rect 197 600 271 634
rect 197 548 210 600
rect 262 548 271 600
rect 197 534 271 548
rect 75 509 149 521
rect 75 457 84 509
rect 136 457 149 509
rect 75 441 149 457
rect 316 507 395 522
rect 316 455 334 507
rect 386 455 395 507
rect 316 442 395 455
rect 443 509 489 787
rect 542 830 619 846
rect 542 778 555 830
rect 607 778 619 830
rect 781 790 954 836
rect 542 762 619 778
rect 666 617 745 641
rect 666 565 676 617
rect 728 565 745 617
rect 666 555 745 565
rect 780 509 860 521
rect 443 463 625 509
rect 191 293 273 308
rect 191 241 209 293
rect 261 241 273 293
rect 191 226 273 241
rect 443 185 489 463
rect 780 457 805 509
rect 857 457 860 509
rect 780 437 860 457
rect 908 512 954 790
rect 1004 731 1083 1043
rect 1129 944 1207 955
rect 1129 892 1142 944
rect 1194 892 1207 944
rect 1596 942 1675 959
rect 1596 897 1608 942
rect 1129 878 1207 892
rect 1600 890 1608 897
rect 1660 890 1675 942
rect 1600 874 1675 890
rect 1252 831 1425 834
rect 1251 788 1425 831
rect 1004 679 1015 731
rect 1067 679 1083 731
rect 1004 666 1083 679
rect 1133 618 1212 626
rect 1133 566 1146 618
rect 1198 566 1212 618
rect 1133 547 1212 566
rect 908 466 1095 512
rect 1248 508 1329 516
rect 666 295 743 308
rect 666 243 677 295
rect 729 243 743 295
rect 666 230 743 243
rect -23 139 145 185
rect -23 -304 24 139
rect 312 138 489 185
rect 199 -31 273 -18
rect 199 -83 208 -31
rect 260 -83 273 -31
rect 199 -97 273 -83
rect 70 -139 146 -127
rect 70 -191 84 -139
rect 136 -191 146 -139
rect 70 -207 146 -191
rect 312 -141 394 -127
rect 312 -193 334 -141
rect 386 -193 394 -141
rect 312 -208 394 -193
rect 443 -143 489 138
rect 541 183 620 196
rect 908 188 955 466
rect 1248 456 1265 508
rect 1317 456 1329 508
rect 1248 437 1329 456
rect 1379 510 1425 788
rect 1478 828 1554 841
rect 1478 776 1490 828
rect 1542 776 1554 828
rect 1478 767 1554 776
rect 1716 831 1790 845
rect 1716 779 1733 831
rect 1785 779 1790 831
rect 1716 764 1790 779
rect 1601 618 1675 632
rect 1601 566 1614 618
rect 1666 566 1675 618
rect 1601 547 1675 566
rect 1379 464 1560 510
rect 1853 509 1906 1043
rect 1128 295 1207 307
rect 1128 243 1140 295
rect 1192 243 1207 295
rect 1128 230 1207 243
rect 541 131 555 183
rect 607 131 620 183
rect 782 141 955 188
rect 541 115 620 131
rect 666 -31 742 -19
rect 666 -83 676 -31
rect 728 -83 742 -31
rect 666 -97 742 -83
rect 791 -120 862 -107
rect 443 -189 624 -143
rect 791 -172 805 -120
rect 857 -172 862 -120
rect 443 -257 489 -189
rect 791 -194 862 -172
rect 908 -140 955 141
rect 1003 185 1092 191
rect 1379 186 1426 464
rect 1495 463 1506 464
rect 1552 463 1560 464
rect 1716 463 1906 509
rect 1601 293 1675 307
rect 1601 241 1614 293
rect 1666 241 1675 293
rect 1601 227 1675 241
rect 1003 133 1015 185
rect 1067 133 1092 185
rect 1253 183 1426 186
rect 1251 139 1426 183
rect 1003 119 1092 133
rect 1128 -29 1208 -22
rect 1128 -81 1144 -29
rect 1196 -81 1208 -29
rect 1128 -96 1208 -81
rect 1010 -140 1086 -135
rect 1248 -140 1329 -127
rect 908 -141 1094 -140
rect 908 -186 1022 -141
rect 1010 -193 1022 -186
rect 1074 -186 1094 -141
rect 1074 -193 1086 -186
rect 1010 -211 1086 -193
rect 1248 -192 1265 -140
rect 1317 -192 1329 -140
rect 1248 -210 1329 -192
rect 1379 -142 1426 139
rect 1478 184 1554 197
rect 1478 132 1490 184
rect 1542 132 1554 184
rect 1478 120 1554 132
rect 1716 183 1790 198
rect 1716 131 1733 183
rect 1785 131 1790 183
rect 1716 118 1790 131
rect 1596 -32 1675 -22
rect 1596 -84 1609 -32
rect 1661 -84 1675 -32
rect 1596 -97 1675 -84
rect 1860 -138 1906 463
rect 1495 -142 1506 -141
rect 1379 -188 1548 -142
rect 1379 -242 1441 -188
rect 1716 -191 1906 -138
rect 1379 -257 1665 -242
rect 443 -304 1665 -257
rect -362 -351 24 -304
rect 1603 -348 1665 -304
rect 315 -445 1518 -399
rect 1603 -410 2101 -348
rect -358 -512 19 -466
rect -358 -990 -311 -512
rect -27 -584 19 -512
rect -133 -897 -87 -584
rect -27 -630 137 -584
rect 315 -630 361 -445
rect 669 -537 1163 -491
rect 421 -574 593 -561
rect 421 -626 529 -574
rect 581 -584 593 -574
rect 581 -626 596 -584
rect 421 -630 596 -626
rect -27 -784 19 -630
rect 421 -637 593 -630
rect 193 -683 266 -657
rect 421 -674 486 -637
rect 193 -735 204 -683
rect 256 -735 266 -683
rect 193 -749 266 -735
rect 410 -689 486 -674
rect 669 -683 715 -537
rect 895 -680 941 -583
rect 1117 -680 1163 -537
rect 1223 -570 1411 -557
rect 1223 -622 1235 -570
rect 1287 -622 1411 -570
rect 1223 -634 1411 -622
rect 1469 -580 1518 -445
rect 1727 -572 1939 -543
rect 1469 -626 1642 -580
rect 1356 -669 1411 -634
rect 410 -735 425 -689
rect 471 -735 486 -689
rect 410 -752 486 -735
rect 539 -729 715 -683
rect 778 -726 1056 -680
rect 1117 -726 1289 -680
rect -27 -830 137 -784
rect 315 -897 361 -784
rect 539 -830 585 -729
rect 649 -784 723 -775
rect 649 -788 729 -784
rect 649 -840 659 -788
rect 711 -840 729 -788
rect 649 -851 729 -840
rect 778 -897 824 -726
rect -133 -943 824 -897
rect 890 -990 939 -783
rect 1010 -895 1056 -726
rect 1234 -762 1289 -726
rect 1356 -684 1423 -669
rect 1356 -730 1362 -684
rect 1408 -730 1423 -684
rect 1356 -745 1423 -730
rect 1107 -784 1183 -772
rect 1107 -836 1119 -784
rect 1171 -836 1183 -784
rect 1107 -848 1183 -836
rect 1234 -775 1310 -762
rect 1234 -827 1247 -775
rect 1299 -827 1310 -775
rect 1234 -839 1310 -827
rect 1468 -895 1519 -780
rect 1010 -941 1519 -895
rect 1596 -990 1642 -626
rect 1727 -624 1749 -572
rect 1801 -624 1939 -572
rect 1727 -653 1939 -624
rect 1752 -766 1954 -743
rect 2039 -766 2101 -410
rect 1752 -775 2101 -766
rect 1752 -827 1772 -775
rect 1824 -827 2101 -775
rect 1752 -828 2101 -827
rect 1752 -853 1954 -828
rect -928 -1066 1872 -990
rect -928 -1112 -803 -1066
rect -757 -1112 -603 -1066
rect -557 -1112 -403 -1066
rect -357 -1112 -203 -1066
rect -157 -1112 -3 -1066
rect 43 -1112 197 -1066
rect 243 -1112 397 -1066
rect 443 -1112 597 -1066
rect 643 -1112 797 -1066
rect 843 -1112 997 -1066
rect 1043 -1112 1197 -1066
rect 1243 -1112 1397 -1066
rect 1443 -1112 1597 -1066
rect 1643 -1112 1872 -1066
rect -928 -1188 1872 -1112
<< via1 >>
rect 78 1697 130 1749
rect 81 1152 133 1204
rect 1736 1162 1788 1214
rect -879 -651 -827 -599
rect 212 923 264 937
rect 212 885 218 923
rect 218 885 264 923
rect 680 943 732 946
rect 680 897 682 943
rect 682 897 728 943
rect 728 897 732 943
rect 680 894 732 897
rect 210 596 262 600
rect 210 550 212 596
rect 212 550 258 596
rect 258 550 262 596
rect 210 548 262 550
rect 84 457 136 509
rect 334 455 386 507
rect 555 778 607 830
rect 676 614 728 617
rect 676 568 678 614
rect 678 568 724 614
rect 724 568 728 614
rect 676 565 728 568
rect 209 291 261 293
rect 209 245 212 291
rect 212 245 258 291
rect 258 245 261 291
rect 209 241 261 245
rect 805 457 857 509
rect 1142 940 1194 944
rect 1142 894 1145 940
rect 1145 894 1191 940
rect 1191 894 1194 940
rect 1142 892 1194 894
rect 1608 937 1660 942
rect 1608 891 1612 937
rect 1612 891 1658 937
rect 1658 891 1660 937
rect 1608 890 1660 891
rect 1015 679 1067 731
rect 1146 614 1198 618
rect 1146 568 1148 614
rect 1148 568 1194 614
rect 1194 568 1198 614
rect 1146 566 1198 568
rect 677 291 729 295
rect 677 245 680 291
rect 680 245 726 291
rect 726 245 729 291
rect 677 243 729 245
rect 208 -35 260 -31
rect 208 -81 211 -35
rect 211 -81 257 -35
rect 257 -81 260 -35
rect 208 -83 260 -81
rect 84 -191 136 -139
rect 334 -193 386 -141
rect 1265 456 1317 508
rect 1490 776 1542 828
rect 1733 779 1785 831
rect 1614 615 1666 618
rect 1614 569 1616 615
rect 1616 569 1662 615
rect 1662 569 1666 615
rect 1614 566 1666 569
rect 1140 291 1192 295
rect 1140 245 1143 291
rect 1143 245 1189 291
rect 1189 245 1192 291
rect 1140 243 1192 245
rect 555 131 607 183
rect 676 -35 728 -31
rect 676 -81 678 -35
rect 678 -81 724 -35
rect 724 -81 728 -35
rect 676 -83 728 -81
rect 805 -172 857 -120
rect 1614 292 1666 293
rect 1614 246 1616 292
rect 1616 246 1662 292
rect 1662 246 1666 292
rect 1614 241 1666 246
rect 1015 133 1067 185
rect 1144 -33 1196 -29
rect 1144 -79 1145 -33
rect 1145 -79 1191 -33
rect 1191 -79 1196 -33
rect 1144 -81 1196 -79
rect 1022 -193 1074 -141
rect 1265 -192 1317 -140
rect 1490 132 1542 184
rect 1733 131 1785 183
rect 1609 -34 1661 -32
rect 1609 -80 1612 -34
rect 1612 -80 1658 -34
rect 1658 -80 1661 -34
rect 1609 -84 1661 -80
rect 529 -626 581 -574
rect 204 -686 256 -683
rect 204 -732 206 -686
rect 206 -732 252 -686
rect 252 -732 256 -686
rect 204 -735 256 -732
rect 1235 -622 1287 -570
rect 659 -840 711 -788
rect 1119 -836 1171 -784
rect 1247 -827 1299 -775
rect 1749 -624 1801 -572
rect 1772 -827 1824 -775
<< metal2 >>
rect 54 1759 145 1774
rect 54 1758 275 1759
rect 54 1749 480 1758
rect 54 1697 78 1749
rect 130 1697 480 1749
rect 54 1686 480 1697
rect 54 1675 145 1686
rect 73 1204 142 1214
rect 73 1152 81 1204
rect 133 1152 142 1204
rect 73 509 142 1152
rect 408 974 480 1686
rect 1721 1214 1806 1222
rect 1721 1162 1736 1214
rect 1788 1162 1806 1214
rect 1721 1155 1806 1162
rect 73 457 84 509
rect 136 457 142 509
rect 73 -139 142 457
rect 199 946 1675 974
rect 199 937 680 946
rect 199 885 212 937
rect 264 902 680 937
rect 264 885 275 902
rect 199 875 275 885
rect 666 894 680 902
rect 732 944 1675 946
rect 732 897 1142 944
rect 732 894 746 897
rect 199 600 273 875
rect 199 548 210 600
rect 262 548 273 600
rect 199 293 273 548
rect 552 830 610 845
rect 552 778 555 830
rect 607 778 610 830
rect 331 507 389 523
rect 331 455 334 507
rect 386 455 389 507
rect 331 315 389 455
rect 552 315 610 778
rect 199 241 209 293
rect 261 241 273 293
rect 330 249 610 315
rect 199 104 273 241
rect 331 104 389 249
rect 552 183 610 249
rect 552 131 555 183
rect 607 131 610 183
rect 552 118 610 131
rect 666 617 746 894
rect 1128 892 1142 897
rect 1194 942 1675 944
rect 1194 897 1608 942
rect 1194 892 1207 897
rect 666 565 676 617
rect 728 565 746 617
rect 666 295 746 565
rect 1004 731 1069 746
rect 1004 679 1015 731
rect 1067 679 1069 731
rect 666 243 677 295
rect 729 243 746 295
rect 199 29 389 104
rect 199 -31 273 29
rect 199 -83 208 -31
rect 260 -83 273 -31
rect 199 -97 273 -83
rect 73 -191 84 -139
rect 136 -191 142 -139
rect 73 -382 142 -191
rect 331 -141 389 29
rect 666 -18 746 243
rect 803 509 873 521
rect 803 457 805 509
rect 857 457 873 509
rect 803 308 873 457
rect 1004 308 1069 679
rect 803 241 1069 308
rect 666 -31 747 -18
rect 666 -83 676 -31
rect 728 -83 747 -31
rect 666 -97 747 -83
rect 331 -193 334 -141
rect 386 -193 389 -141
rect 803 -120 873 241
rect 1004 185 1069 241
rect 1004 133 1015 185
rect 1067 133 1069 185
rect 1004 121 1069 133
rect 1128 618 1207 892
rect 1600 890 1608 897
rect 1660 890 1675 942
rect 1128 566 1146 618
rect 1198 566 1207 618
rect 1128 295 1207 566
rect 1488 828 1544 841
rect 1488 776 1490 828
rect 1542 776 1544 828
rect 1128 243 1140 295
rect 1192 243 1207 295
rect 1128 -29 1207 243
rect 1128 -81 1144 -29
rect 1196 -81 1207 -29
rect 1128 -96 1207 -81
rect 1263 508 1319 521
rect 1263 456 1265 508
rect 1317 456 1319 508
rect 1263 312 1319 456
rect 1488 312 1544 776
rect 1263 241 1544 312
rect 803 -172 805 -120
rect 857 -172 873 -120
rect 803 -186 873 -172
rect 992 -141 1077 -128
rect 992 -143 1022 -141
rect 331 -268 389 -193
rect 992 -199 1008 -143
rect 1074 -193 1077 -141
rect 1064 -199 1077 -193
rect 992 -211 1077 -199
rect 1263 -140 1319 241
rect 1488 184 1544 241
rect 1488 132 1490 184
rect 1542 132 1544 184
rect 1488 119 1544 132
rect 1600 618 1675 890
rect 1600 566 1614 618
rect 1666 566 1675 618
rect 1600 293 1675 566
rect 1600 241 1614 293
rect 1666 241 1675 293
rect 1600 -32 1675 241
rect 1600 -84 1609 -32
rect 1661 -84 1675 -32
rect 1600 -97 1675 -84
rect 1731 831 1790 1155
rect 1731 779 1733 831
rect 1785 779 1790 831
rect 1731 199 1790 779
rect 1731 187 1811 199
rect 1731 183 1744 187
rect 1731 131 1733 183
rect 1800 131 1811 187
rect 1731 116 1811 131
rect 1263 -192 1265 -140
rect 1317 -192 1319 -140
rect 1263 -268 1319 -192
rect 331 -326 1319 -268
rect 1731 -382 1790 116
rect 73 -451 1790 -382
rect 1727 -557 1833 -543
rect 517 -570 1833 -557
rect 517 -574 1235 -570
rect -899 -588 -809 -574
rect -899 -599 266 -588
rect -899 -651 -879 -599
rect -827 -651 266 -599
rect 517 -626 529 -574
rect 581 -622 1235 -574
rect 1287 -572 1833 -570
rect 1287 -622 1749 -572
rect 581 -624 1749 -622
rect 1801 -624 1833 -572
rect 581 -626 1833 -624
rect 517 -637 1833 -626
rect 593 -638 1833 -637
rect -899 -661 266 -651
rect -899 -673 -809 -661
rect 193 -683 266 -661
rect 193 -735 204 -683
rect 256 -735 266 -683
rect 193 -749 266 -735
rect 803 -771 860 -638
rect 1727 -653 1833 -638
rect 1752 -762 1853 -743
rect 648 -784 1183 -771
rect 648 -788 1119 -784
rect 648 -840 659 -788
rect 711 -836 1119 -788
rect 1171 -836 1183 -784
rect 711 -840 1183 -836
rect 1239 -775 1853 -762
rect 1239 -827 1247 -775
rect 1299 -827 1772 -775
rect 1824 -827 1853 -775
rect 1239 -839 1853 -827
rect 648 -851 1183 -840
rect 1752 -853 1853 -839
<< via2 >>
rect 1008 -193 1022 -143
rect 1022 -193 1064 -143
rect 1008 -199 1064 -193
rect 1744 183 1800 187
rect 1744 131 1785 183
rect 1785 131 1800 183
<< metal3 >>
rect 1734 187 1811 199
rect 1734 131 1744 187
rect 1800 131 1811 187
rect 992 -129 1077 -128
rect 1734 -129 1811 131
rect 992 -143 1811 -129
rect 992 -199 1008 -143
rect 1064 -199 1811 -143
rect 992 -211 1811 -199
rect 1076 -212 1811 -211
use nmos_3p3_FYTGVN  nmos_3p3_FYTGVN_0
timestamp 1713185578
transform 1 0 1380 0 1 -803
box -172 -100 172 100
use nmos_3p3_FYTGVN  nmos_3p3_FYTGVN_1
timestamp 1713185578
transform 1 0 450 0 1 -807
box -172 -100 172 100
use nmos_3p3_FYTGVN  nmos_3p3_FYTGVN_2
timestamp 1713185578
transform 1 0 226 0 1 -807
box -172 -100 172 100
use nmos_3p3_FYTGVN  nmos_3p3_FYTGVN_4
timestamp 1713185578
transform 1 0 450 0 1 -607
box -172 -100 172 100
use nmos_3p3_FYTGVN  nmos_3p3_FYTGVN_7
timestamp 1713185578
transform 1 0 1380 0 1 -603
box -172 -100 172 100
use nmos_3p3_GYTGVN  nmos_3p3_GYTGVN_0
timestamp 1713185578
transform 1 0 916 0 1 -806
box -284 -100 284 100
use nmos_3p3_GYTGVN  nmos_3p3_GYTGVN_1
timestamp 1713185578
transform 1 0 916 0 1 -606
box -284 -100 284 100
use nmos_3p3_GYTGVN  nmos_3p3_GYTGVN_2
timestamp 1713185578
transform 1 0 -110 0 1 -807
box -284 -100 284 100
use nmos_3p3_GYTGVN  nmos_3p3_GYTGVN_3
timestamp 1713185578
transform 1 0 -110 0 1 -607
box -284 -100 284 100
use nmos_3p3_XYTGVN  nmos_3p3_XYTGVN_0
timestamp 1713185578
transform 1 0 -574 0 1 -712
box -172 -196 172 196
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_0
timestamp 1713185578
transform 1 0 234 0 1 486
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_1
timestamp 1713185578
transform 1 0 234 0 1 -162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_2
timestamp 1713185578
transform 1 0 702 0 1 -162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_3
timestamp 1713185578
transform 1 0 1170 0 1 -162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_4
timestamp 1713185578
transform 1 0 1638 0 1 -162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_5
timestamp 1713185578
transform 1 0 702 0 1 486
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_6
timestamp 1713185578
transform 1 0 1170 0 1 486
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_7
timestamp 1713185578
transform 1 0 1638 0 1 486
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_8
timestamp 1713185578
transform 1 0 234 0 1 810
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_9
timestamp 1713185578
transform 1 0 702 0 1 810
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_10
timestamp 1713185578
transform 1 0 1170 0 1 810
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_11
timestamp 1713185578
transform 1 0 1638 0 1 810
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_12
timestamp 1713185578
transform 1 0 1638 0 1 162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_13
timestamp 1713185578
transform 1 0 1170 0 1 162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_14
timestamp 1713185578
transform 1 0 702 0 1 162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_15
timestamp 1713185578
transform 1 0 234 0 1 162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_16
timestamp 1713185578
transform 1 0 -694 0 1 162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_17
timestamp 1713185578
transform 1 0 -694 0 1 -162
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_18
timestamp 1713185578
transform 1 0 -694 0 1 810
box -234 -162 234 162
use pmos_3p3_MDK7F7  pmos_3p3_MDK7F7_19
timestamp 1713185578
transform 1 0 -694 0 1 486
box -234 -162 234 162
use pmos_3p3_RL7FD7  pmos_3p3_RL7FD7_0
timestamp 1713185578
transform 1 0 -230 0 1 290
box -230 -614 230 614
<< labels >>
flabel nsubdiffcont 555 1244 555 1244 0 FreeSans 2500 0 0 0 VDD
flabel psubdiffcont 620 -1089 620 -1089 0 FreeSans 750 0 0 0 VSS
flabel metal1 s -870 -339 -870 -339 0 FreeSans 2500 0 0 0 UP
port 1 nsew
flabel metal1 s -1089 -626 -1089 -626 0 FreeSans 2500 0 0 0 down
port 2 nsew
flabel metal1 s 1928 -809 1928 -809 0 FreeSans 2500 0 0 0 VCTRL
port 3 nsew
flabel metal1 s 1909 -590 1909 -590 0 FreeSans 2500 0 0 0 ITAIL1
port 4 nsew
flabel metal1 s -43 1710 -43 1710 0 FreeSans 2500 0 0 0 ITAIL
port 5 nsew
<< end >>
