** sch_path: /home/shahid/GF180Projects/Divider/Xschem/DIFF_CLK_div_4_TB.sch
**.subckt DIFF_CLK_div_4_TB
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 CLK VSS pulse(3.3 0 0 100p 100p 2.50n 5n)
.save i(v3)
C1 Vdiv4 VSS 1p m=1
C2 Vdiv4B VSS 1p m=1
V5 RST VSS PWL( 0 0 10n 0 10.001n 3)
.save i(v5)
V4 CLKB VSS pulse(0 3.3 0 100p 100p 2.50n 5n)
.save i(v4)
x1 VSS VDD RST Vdiv4 Vdiv4B CLKB CLK DIFFER_CLK_div_4
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical




.control
save all
tran 50p 100n
plot v(CLK) v(Vdiv4)+3.5 v(Vdiv4B)+7 v(RST)+10.5
write DIFF_CLK_div_4_TB.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  DIFFER_CLK_div_4.sym # of pins=7
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/DIFFER_CLK_div_4.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/DIFFER_CLK_div_4.sch
.subckt DIFFER_CLK_div_4 VSS VDD RST Vdiv4 Vdiv4B CLKB CLK
*.ipin CLK
*.iopin VSS
*.iopin VDD
*.ipin RST
*.opin Vdiv4
*.opin Vdiv4B
*.ipin CLKB
x1 VSS VDD net1 Vdiv4B RST CLKB Diff_CLK_div_4
x2 VSS VDD net2 Vdiv4 RST CLK CLK_div_4
.ends


* expanding   symbol:  Diff_CLK_div_4.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/Diff_CLK_div_4.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/Diff_CLK_div_4.sch
.subckt Diff_CLK_div_4 VSS VDD Q0 Q1 RST CLK
*.ipin CLK
*.iopin VSS
*.iopin VDD
*.opin Q0
*.opin Q1
*.ipin RST
x1 CLK VSS VDD net1 VDD net4 RST VDD Diff_JK_flipflop
x2 Q0 VSS VDD net2 VDD net5 RST VDD Diff_JK_flipflop
x3 VSS VDD Q0 net1 GF_INV
x4 VSS VDD net3 net2 GF_INV
x5 VSS net3 Q1 VDD Load_BUFF
.ends


* expanding   symbol:  CLK_div_4.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/CLK_div_4.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/CLK_div_4.sch
.subckt CLK_div_4 VSS VDD Q0 Q1 RST CLK
*.ipin CLK
*.iopin VSS
*.iopin VDD
*.opin Q0
*.opin Q1
*.ipin RST
x1 CLK VSS VDD Q0 VDD net2 RST VDD JK_flipflop
x2 Q0 VSS VDD net1 VDD net3 RST VDD JK_flipflop
x3 VSS net1 Q1 VDD Load_BUFF
.ends


* expanding   symbol:  Diff_JK_flipflop.sym # of pins=8
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/Diff_JK_flipflop.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/Diff_JK_flipflop.sch
.subckt Diff_JK_flipflop CLK VSS VDD Q J Qb RST K
*.ipin K
*.ipin CLK
*.iopin VSS
*.iopin VDD
*.opin Q
*.ipin J
*.opin Qb
*.ipin RST
x1 J VSS VDD net5 Qb CLK_b nand_3
x2 CLK_b VSS VDD net6 Q K nand_3
x9 VSS VDD CLK_b CLK GF_INV
x3 net5 VSS VDD net1 net2 NAND
x5 CLK VSS VDD net3 net2 NAND
x6 net1 VSS VDD net4 CLK NAND
x7 net4 VSS VDD Q Qb NAND
x8 net3 VSS VDD Qb Q NAND
x4 net6 VSS VDD net2 net1 RST nand_3
.ends


* expanding   symbol:  GF_INV.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/GF_INV.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/GF_INV.sch
.subckt GF_INV VSS VDD OUT IN
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  Load_BUFF.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/Load_BUFF.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/Load_BUFF.sch
.subckt Load_BUFF VSS IN OUT VDD
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
x3 VSS VDD net1 IN INV_BUFF
x1 VSS VDD OUT net1 INV_BUFF
.ends


* expanding   symbol:  JK_flipflop.sym # of pins=8
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/JK_flipflop.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/JK_flipflop.sch
.subckt JK_flipflop CLK VSS VDD Q J Qb RST K
*.ipin K
*.ipin CLK
*.iopin VSS
*.iopin VDD
*.opin Q
*.ipin J
*.opin Qb
*.ipin RST
x1 J VSS VDD net5 Qb CLK nand_3
x2 CLK VSS VDD net6 Q K nand_3
x4 net6 VSS VDD net2 net1 RST nand_3
x9 VSS VDD CLK_b CLK GF_INV
x3 net5 VSS VDD net1 net2 NAND
x5 CLK_b VSS VDD net3 net2 NAND
x6 net1 VSS VDD net4 CLK_b NAND
x7 net4 VSS VDD Q Qb NAND
x8 net3 VSS VDD Qb Q NAND
.ends


* expanding   symbol:  nand_3.sym # of pins=6
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/nand_3.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/nand_3.sch
.subckt nand_3 IN1 VSS VDD OUT IN3 IN2
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin OUT
*.ipin IN3
XM3 net1 IN3 VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=3
XM4 OUT IN1 net2 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=3
XM1 OUT IN3 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN1 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM7 net2 IN2 net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=3
XM8 OUT IN2 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  NAND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/NAND.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/NAND.sch
.subckt NAND IN1 VSS VDD OUT IN2
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin OUT
XM3 net1 IN2 VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM4 OUT IN1 net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM5 OUT IN1 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN2 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  INV_BUFF.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/Divider/Xschem/INV_BUFF.sym
** sch_path: /home/shahid/GF180Projects/Divider/Xschem/INV_BUFF.sch
.subckt INV_BUFF VSS VDD OUT IN
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=14.08u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=51.2u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
