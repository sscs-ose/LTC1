magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1085 -1646 1085 1646
<< metal1 >>
rect -85 640 85 646
rect -85 614 -79 640
rect -53 614 -13 640
rect 13 614 53 640
rect 79 614 85 640
rect -85 574 85 614
rect -85 548 -79 574
rect -53 548 -13 574
rect 13 548 53 574
rect 79 548 85 574
rect -85 508 85 548
rect -85 482 -79 508
rect -53 482 -13 508
rect 13 482 53 508
rect 79 482 85 508
rect -85 442 85 482
rect -85 416 -79 442
rect -53 416 -13 442
rect 13 416 53 442
rect 79 416 85 442
rect -85 376 85 416
rect -85 350 -79 376
rect -53 350 -13 376
rect 13 350 53 376
rect 79 350 85 376
rect -85 310 85 350
rect -85 284 -79 310
rect -53 284 -13 310
rect 13 284 53 310
rect 79 284 85 310
rect -85 244 85 284
rect -85 218 -79 244
rect -53 218 -13 244
rect 13 218 53 244
rect 79 218 85 244
rect -85 178 85 218
rect -85 152 -79 178
rect -53 152 -13 178
rect 13 152 53 178
rect 79 152 85 178
rect -85 112 85 152
rect -85 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 85 112
rect -85 46 85 86
rect -85 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 85 46
rect -85 -20 85 20
rect -85 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 85 -20
rect -85 -86 85 -46
rect -85 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 85 -86
rect -85 -152 85 -112
rect -85 -178 -79 -152
rect -53 -178 -13 -152
rect 13 -178 53 -152
rect 79 -178 85 -152
rect -85 -218 85 -178
rect -85 -244 -79 -218
rect -53 -244 -13 -218
rect 13 -244 53 -218
rect 79 -244 85 -218
rect -85 -284 85 -244
rect -85 -310 -79 -284
rect -53 -310 -13 -284
rect 13 -310 53 -284
rect 79 -310 85 -284
rect -85 -350 85 -310
rect -85 -376 -79 -350
rect -53 -376 -13 -350
rect 13 -376 53 -350
rect 79 -376 85 -350
rect -85 -416 85 -376
rect -85 -442 -79 -416
rect -53 -442 -13 -416
rect 13 -442 53 -416
rect 79 -442 85 -416
rect -85 -482 85 -442
rect -85 -508 -79 -482
rect -53 -508 -13 -482
rect 13 -508 53 -482
rect 79 -508 85 -482
rect -85 -548 85 -508
rect -85 -574 -79 -548
rect -53 -574 -13 -548
rect 13 -574 53 -548
rect 79 -574 85 -548
rect -85 -614 85 -574
rect -85 -640 -79 -614
rect -53 -640 -13 -614
rect 13 -640 53 -614
rect 79 -640 85 -614
rect -85 -646 85 -640
<< via1 >>
rect -79 614 -53 640
rect -13 614 13 640
rect 53 614 79 640
rect -79 548 -53 574
rect -13 548 13 574
rect 53 548 79 574
rect -79 482 -53 508
rect -13 482 13 508
rect 53 482 79 508
rect -79 416 -53 442
rect -13 416 13 442
rect 53 416 79 442
rect -79 350 -53 376
rect -13 350 13 376
rect 53 350 79 376
rect -79 284 -53 310
rect -13 284 13 310
rect 53 284 79 310
rect -79 218 -53 244
rect -13 218 13 244
rect 53 218 79 244
rect -79 152 -53 178
rect -13 152 13 178
rect 53 152 79 178
rect -79 86 -53 112
rect -13 86 13 112
rect 53 86 79 112
rect -79 20 -53 46
rect -13 20 13 46
rect 53 20 79 46
rect -79 -46 -53 -20
rect -13 -46 13 -20
rect 53 -46 79 -20
rect -79 -112 -53 -86
rect -13 -112 13 -86
rect 53 -112 79 -86
rect -79 -178 -53 -152
rect -13 -178 13 -152
rect 53 -178 79 -152
rect -79 -244 -53 -218
rect -13 -244 13 -218
rect 53 -244 79 -218
rect -79 -310 -53 -284
rect -13 -310 13 -284
rect 53 -310 79 -284
rect -79 -376 -53 -350
rect -13 -376 13 -350
rect 53 -376 79 -350
rect -79 -442 -53 -416
rect -13 -442 13 -416
rect 53 -442 79 -416
rect -79 -508 -53 -482
rect -13 -508 13 -482
rect 53 -508 79 -482
rect -79 -574 -53 -548
rect -13 -574 13 -548
rect 53 -574 79 -548
rect -79 -640 -53 -614
rect -13 -640 13 -614
rect 53 -640 79 -614
<< metal2 >>
rect -85 640 85 646
rect -85 614 -79 640
rect -53 614 -13 640
rect 13 614 53 640
rect 79 614 85 640
rect -85 574 85 614
rect -85 548 -79 574
rect -53 548 -13 574
rect 13 548 53 574
rect 79 548 85 574
rect -85 508 85 548
rect -85 482 -79 508
rect -53 482 -13 508
rect 13 482 53 508
rect 79 482 85 508
rect -85 442 85 482
rect -85 416 -79 442
rect -53 416 -13 442
rect 13 416 53 442
rect 79 416 85 442
rect -85 376 85 416
rect -85 350 -79 376
rect -53 350 -13 376
rect 13 350 53 376
rect 79 350 85 376
rect -85 310 85 350
rect -85 284 -79 310
rect -53 284 -13 310
rect 13 284 53 310
rect 79 284 85 310
rect -85 244 85 284
rect -85 218 -79 244
rect -53 218 -13 244
rect 13 218 53 244
rect 79 218 85 244
rect -85 178 85 218
rect -85 152 -79 178
rect -53 152 -13 178
rect 13 152 53 178
rect 79 152 85 178
rect -85 112 85 152
rect -85 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 85 112
rect -85 46 85 86
rect -85 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 85 46
rect -85 -20 85 20
rect -85 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 85 -20
rect -85 -86 85 -46
rect -85 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 85 -86
rect -85 -152 85 -112
rect -85 -178 -79 -152
rect -53 -178 -13 -152
rect 13 -178 53 -152
rect 79 -178 85 -152
rect -85 -218 85 -178
rect -85 -244 -79 -218
rect -53 -244 -13 -218
rect 13 -244 53 -218
rect 79 -244 85 -218
rect -85 -284 85 -244
rect -85 -310 -79 -284
rect -53 -310 -13 -284
rect 13 -310 53 -284
rect 79 -310 85 -284
rect -85 -350 85 -310
rect -85 -376 -79 -350
rect -53 -376 -13 -350
rect 13 -376 53 -350
rect 79 -376 85 -350
rect -85 -416 85 -376
rect -85 -442 -79 -416
rect -53 -442 -13 -416
rect 13 -442 53 -416
rect 79 -442 85 -416
rect -85 -482 85 -442
rect -85 -508 -79 -482
rect -53 -508 -13 -482
rect 13 -508 53 -482
rect 79 -508 85 -482
rect -85 -548 85 -508
rect -85 -574 -79 -548
rect -53 -574 -13 -548
rect 13 -574 53 -548
rect 79 -574 85 -548
rect -85 -614 85 -574
rect -85 -640 -79 -614
rect -53 -640 -13 -614
rect 13 -640 53 -614
rect 79 -640 85 -614
rect -85 -646 85 -640
<< end >>
