magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1046 -1208 1046 1208
<< metal1 >>
rect -46 202 46 208
rect -46 176 -40 202
rect -14 176 14 202
rect 40 176 46 202
rect -46 148 46 176
rect -46 122 -40 148
rect -14 122 14 148
rect 40 122 46 148
rect -46 94 46 122
rect -46 68 -40 94
rect -14 68 14 94
rect 40 68 46 94
rect -46 40 46 68
rect -46 14 -40 40
rect -14 14 14 40
rect 40 14 46 40
rect -46 -14 46 14
rect -46 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 46 -14
rect -46 -68 46 -40
rect -46 -94 -40 -68
rect -14 -94 14 -68
rect 40 -94 46 -68
rect -46 -122 46 -94
rect -46 -148 -40 -122
rect -14 -148 14 -122
rect 40 -148 46 -122
rect -46 -176 46 -148
rect -46 -202 -40 -176
rect -14 -202 14 -176
rect 40 -202 46 -176
rect -46 -208 46 -202
<< via1 >>
rect -40 176 -14 202
rect 14 176 40 202
rect -40 122 -14 148
rect 14 122 40 148
rect -40 68 -14 94
rect 14 68 40 94
rect -40 14 -14 40
rect 14 14 40 40
rect -40 -40 -14 -14
rect 14 -40 40 -14
rect -40 -94 -14 -68
rect 14 -94 40 -68
rect -40 -148 -14 -122
rect 14 -148 40 -122
rect -40 -202 -14 -176
rect 14 -202 40 -176
<< metal2 >>
rect -46 202 46 208
rect -46 176 -40 202
rect -14 176 14 202
rect 40 176 46 202
rect -46 148 46 176
rect -46 122 -40 148
rect -14 122 14 148
rect 40 122 46 148
rect -46 94 46 122
rect -46 68 -40 94
rect -14 68 14 94
rect 40 68 46 94
rect -46 40 46 68
rect -46 14 -40 40
rect -14 14 14 40
rect 40 14 46 40
rect -46 -14 46 14
rect -46 -40 -40 -14
rect -14 -40 14 -14
rect 40 -40 46 -14
rect -46 -68 46 -40
rect -46 -94 -40 -68
rect -14 -94 14 -68
rect 40 -94 46 -68
rect -46 -122 46 -94
rect -46 -148 -40 -122
rect -14 -148 14 -122
rect 40 -148 46 -122
rect -46 -176 46 -148
rect -46 -202 -40 -176
rect -14 -202 14 -176
rect 40 -202 46 -176
rect -46 -208 46 -202
<< end >>
