magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3408 -2045 3408 2045
<< psubdiff >>
rect -1408 23 1408 45
rect -1408 -23 -1386 23
rect 1386 -23 1408 23
rect -1408 -45 1408 -23
<< psubdiffcont >>
rect -1386 -23 1386 23
<< metal1 >>
rect -1397 23 1397 34
rect -1397 -23 -1386 23
rect 1386 -23 1397 23
rect -1397 -34 1397 -23
<< end >>
