magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1205 -1329 1205 1329
<< metal2 >>
rect -205 324 205 329
rect -205 296 -200 324
rect -172 296 -138 324
rect -110 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 110 324
rect 138 296 172 324
rect 200 296 205 324
rect -205 262 205 296
rect -205 234 -200 262
rect -172 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 172 262
rect 200 234 205 262
rect -205 200 205 234
rect -205 172 -200 200
rect -172 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 172 200
rect 200 172 205 200
rect -205 138 205 172
rect -205 110 -200 138
rect -172 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 172 138
rect 200 110 205 138
rect -205 76 205 110
rect -205 48 -200 76
rect -172 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 172 76
rect 200 48 205 76
rect -205 14 205 48
rect -205 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 205 14
rect -205 -48 205 -14
rect -205 -76 -200 -48
rect -172 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 172 -48
rect 200 -76 205 -48
rect -205 -110 205 -76
rect -205 -138 -200 -110
rect -172 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 172 -110
rect 200 -138 205 -110
rect -205 -172 205 -138
rect -205 -200 -200 -172
rect -172 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 172 -172
rect 200 -200 205 -172
rect -205 -234 205 -200
rect -205 -262 -200 -234
rect -172 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 172 -234
rect 200 -262 205 -234
rect -205 -296 205 -262
rect -205 -324 -200 -296
rect -172 -324 -138 -296
rect -110 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 110 -296
rect 138 -324 172 -296
rect 200 -324 205 -296
rect -205 -329 205 -324
<< via2 >>
rect -200 296 -172 324
rect -138 296 -110 324
rect -76 296 -48 324
rect -14 296 14 324
rect 48 296 76 324
rect 110 296 138 324
rect 172 296 200 324
rect -200 234 -172 262
rect -138 234 -110 262
rect -76 234 -48 262
rect -14 234 14 262
rect 48 234 76 262
rect 110 234 138 262
rect 172 234 200 262
rect -200 172 -172 200
rect -138 172 -110 200
rect -76 172 -48 200
rect -14 172 14 200
rect 48 172 76 200
rect 110 172 138 200
rect 172 172 200 200
rect -200 110 -172 138
rect -138 110 -110 138
rect -76 110 -48 138
rect -14 110 14 138
rect 48 110 76 138
rect 110 110 138 138
rect 172 110 200 138
rect -200 48 -172 76
rect -138 48 -110 76
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect 110 48 138 76
rect 172 48 200 76
rect -200 -14 -172 14
rect -138 -14 -110 14
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect 110 -14 138 14
rect 172 -14 200 14
rect -200 -76 -172 -48
rect -138 -76 -110 -48
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect 110 -76 138 -48
rect 172 -76 200 -48
rect -200 -138 -172 -110
rect -138 -138 -110 -110
rect -76 -138 -48 -110
rect -14 -138 14 -110
rect 48 -138 76 -110
rect 110 -138 138 -110
rect 172 -138 200 -110
rect -200 -200 -172 -172
rect -138 -200 -110 -172
rect -76 -200 -48 -172
rect -14 -200 14 -172
rect 48 -200 76 -172
rect 110 -200 138 -172
rect 172 -200 200 -172
rect -200 -262 -172 -234
rect -138 -262 -110 -234
rect -76 -262 -48 -234
rect -14 -262 14 -234
rect 48 -262 76 -234
rect 110 -262 138 -234
rect 172 -262 200 -234
rect -200 -324 -172 -296
rect -138 -324 -110 -296
rect -76 -324 -48 -296
rect -14 -324 14 -296
rect 48 -324 76 -296
rect 110 -324 138 -296
rect 172 -324 200 -296
<< metal3 >>
rect -205 324 205 329
rect -205 296 -200 324
rect -172 296 -138 324
rect -110 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 110 324
rect 138 296 172 324
rect 200 296 205 324
rect -205 262 205 296
rect -205 234 -200 262
rect -172 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 172 262
rect 200 234 205 262
rect -205 200 205 234
rect -205 172 -200 200
rect -172 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 172 200
rect 200 172 205 200
rect -205 138 205 172
rect -205 110 -200 138
rect -172 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 172 138
rect 200 110 205 138
rect -205 76 205 110
rect -205 48 -200 76
rect -172 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 172 76
rect 200 48 205 76
rect -205 14 205 48
rect -205 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 205 14
rect -205 -48 205 -14
rect -205 -76 -200 -48
rect -172 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 172 -48
rect 200 -76 205 -48
rect -205 -110 205 -76
rect -205 -138 -200 -110
rect -172 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 172 -110
rect 200 -138 205 -110
rect -205 -172 205 -138
rect -205 -200 -200 -172
rect -172 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 172 -172
rect 200 -200 205 -172
rect -205 -234 205 -200
rect -205 -262 -200 -234
rect -172 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 172 -234
rect 200 -262 205 -234
rect -205 -296 205 -262
rect -205 -324 -200 -296
rect -172 -324 -138 -296
rect -110 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 110 -296
rect 138 -324 172 -296
rect 200 -324 205 -296
rect -205 -329 205 -324
<< end >>
