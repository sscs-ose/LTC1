magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1247 -1665 1247 1665
<< metal2 >>
rect -247 660 247 665
rect -247 632 -242 660
rect -214 632 -166 660
rect -138 632 -90 660
rect -62 632 -14 660
rect 14 632 62 660
rect 90 632 138 660
rect 166 632 214 660
rect 242 632 247 660
rect -247 584 247 632
rect -247 556 -242 584
rect -214 556 -166 584
rect -138 556 -90 584
rect -62 556 -14 584
rect 14 556 62 584
rect 90 556 138 584
rect 166 556 214 584
rect 242 556 247 584
rect -247 508 247 556
rect -247 480 -242 508
rect -214 480 -166 508
rect -138 480 -90 508
rect -62 480 -14 508
rect 14 480 62 508
rect 90 480 138 508
rect 166 480 214 508
rect 242 480 247 508
rect -247 432 247 480
rect -247 404 -242 432
rect -214 404 -166 432
rect -138 404 -90 432
rect -62 404 -14 432
rect 14 404 62 432
rect 90 404 138 432
rect 166 404 214 432
rect 242 404 247 432
rect -247 356 247 404
rect -247 328 -242 356
rect -214 328 -166 356
rect -138 328 -90 356
rect -62 328 -14 356
rect 14 328 62 356
rect 90 328 138 356
rect 166 328 214 356
rect 242 328 247 356
rect -247 280 247 328
rect -247 252 -242 280
rect -214 252 -166 280
rect -138 252 -90 280
rect -62 252 -14 280
rect 14 252 62 280
rect 90 252 138 280
rect 166 252 214 280
rect 242 252 247 280
rect -247 204 247 252
rect -247 176 -242 204
rect -214 176 -166 204
rect -138 176 -90 204
rect -62 176 -14 204
rect 14 176 62 204
rect 90 176 138 204
rect 166 176 214 204
rect 242 176 247 204
rect -247 128 247 176
rect -247 100 -242 128
rect -214 100 -166 128
rect -138 100 -90 128
rect -62 100 -14 128
rect 14 100 62 128
rect 90 100 138 128
rect 166 100 214 128
rect 242 100 247 128
rect -247 52 247 100
rect -247 24 -242 52
rect -214 24 -166 52
rect -138 24 -90 52
rect -62 24 -14 52
rect 14 24 62 52
rect 90 24 138 52
rect 166 24 214 52
rect 242 24 247 52
rect -247 -24 247 24
rect -247 -52 -242 -24
rect -214 -52 -166 -24
rect -138 -52 -90 -24
rect -62 -52 -14 -24
rect 14 -52 62 -24
rect 90 -52 138 -24
rect 166 -52 214 -24
rect 242 -52 247 -24
rect -247 -100 247 -52
rect -247 -128 -242 -100
rect -214 -128 -166 -100
rect -138 -128 -90 -100
rect -62 -128 -14 -100
rect 14 -128 62 -100
rect 90 -128 138 -100
rect 166 -128 214 -100
rect 242 -128 247 -100
rect -247 -176 247 -128
rect -247 -204 -242 -176
rect -214 -204 -166 -176
rect -138 -204 -90 -176
rect -62 -204 -14 -176
rect 14 -204 62 -176
rect 90 -204 138 -176
rect 166 -204 214 -176
rect 242 -204 247 -176
rect -247 -252 247 -204
rect -247 -280 -242 -252
rect -214 -280 -166 -252
rect -138 -280 -90 -252
rect -62 -280 -14 -252
rect 14 -280 62 -252
rect 90 -280 138 -252
rect 166 -280 214 -252
rect 242 -280 247 -252
rect -247 -328 247 -280
rect -247 -356 -242 -328
rect -214 -356 -166 -328
rect -138 -356 -90 -328
rect -62 -356 -14 -328
rect 14 -356 62 -328
rect 90 -356 138 -328
rect 166 -356 214 -328
rect 242 -356 247 -328
rect -247 -404 247 -356
rect -247 -432 -242 -404
rect -214 -432 -166 -404
rect -138 -432 -90 -404
rect -62 -432 -14 -404
rect 14 -432 62 -404
rect 90 -432 138 -404
rect 166 -432 214 -404
rect 242 -432 247 -404
rect -247 -480 247 -432
rect -247 -508 -242 -480
rect -214 -508 -166 -480
rect -138 -508 -90 -480
rect -62 -508 -14 -480
rect 14 -508 62 -480
rect 90 -508 138 -480
rect 166 -508 214 -480
rect 242 -508 247 -480
rect -247 -556 247 -508
rect -247 -584 -242 -556
rect -214 -584 -166 -556
rect -138 -584 -90 -556
rect -62 -584 -14 -556
rect 14 -584 62 -556
rect 90 -584 138 -556
rect 166 -584 214 -556
rect 242 -584 247 -556
rect -247 -632 247 -584
rect -247 -660 -242 -632
rect -214 -660 -166 -632
rect -138 -660 -90 -632
rect -62 -660 -14 -632
rect 14 -660 62 -632
rect 90 -660 138 -632
rect 166 -660 214 -632
rect 242 -660 247 -632
rect -247 -665 247 -660
<< via2 >>
rect -242 632 -214 660
rect -166 632 -138 660
rect -90 632 -62 660
rect -14 632 14 660
rect 62 632 90 660
rect 138 632 166 660
rect 214 632 242 660
rect -242 556 -214 584
rect -166 556 -138 584
rect -90 556 -62 584
rect -14 556 14 584
rect 62 556 90 584
rect 138 556 166 584
rect 214 556 242 584
rect -242 480 -214 508
rect -166 480 -138 508
rect -90 480 -62 508
rect -14 480 14 508
rect 62 480 90 508
rect 138 480 166 508
rect 214 480 242 508
rect -242 404 -214 432
rect -166 404 -138 432
rect -90 404 -62 432
rect -14 404 14 432
rect 62 404 90 432
rect 138 404 166 432
rect 214 404 242 432
rect -242 328 -214 356
rect -166 328 -138 356
rect -90 328 -62 356
rect -14 328 14 356
rect 62 328 90 356
rect 138 328 166 356
rect 214 328 242 356
rect -242 252 -214 280
rect -166 252 -138 280
rect -90 252 -62 280
rect -14 252 14 280
rect 62 252 90 280
rect 138 252 166 280
rect 214 252 242 280
rect -242 176 -214 204
rect -166 176 -138 204
rect -90 176 -62 204
rect -14 176 14 204
rect 62 176 90 204
rect 138 176 166 204
rect 214 176 242 204
rect -242 100 -214 128
rect -166 100 -138 128
rect -90 100 -62 128
rect -14 100 14 128
rect 62 100 90 128
rect 138 100 166 128
rect 214 100 242 128
rect -242 24 -214 52
rect -166 24 -138 52
rect -90 24 -62 52
rect -14 24 14 52
rect 62 24 90 52
rect 138 24 166 52
rect 214 24 242 52
rect -242 -52 -214 -24
rect -166 -52 -138 -24
rect -90 -52 -62 -24
rect -14 -52 14 -24
rect 62 -52 90 -24
rect 138 -52 166 -24
rect 214 -52 242 -24
rect -242 -128 -214 -100
rect -166 -128 -138 -100
rect -90 -128 -62 -100
rect -14 -128 14 -100
rect 62 -128 90 -100
rect 138 -128 166 -100
rect 214 -128 242 -100
rect -242 -204 -214 -176
rect -166 -204 -138 -176
rect -90 -204 -62 -176
rect -14 -204 14 -176
rect 62 -204 90 -176
rect 138 -204 166 -176
rect 214 -204 242 -176
rect -242 -280 -214 -252
rect -166 -280 -138 -252
rect -90 -280 -62 -252
rect -14 -280 14 -252
rect 62 -280 90 -252
rect 138 -280 166 -252
rect 214 -280 242 -252
rect -242 -356 -214 -328
rect -166 -356 -138 -328
rect -90 -356 -62 -328
rect -14 -356 14 -328
rect 62 -356 90 -328
rect 138 -356 166 -328
rect 214 -356 242 -328
rect -242 -432 -214 -404
rect -166 -432 -138 -404
rect -90 -432 -62 -404
rect -14 -432 14 -404
rect 62 -432 90 -404
rect 138 -432 166 -404
rect 214 -432 242 -404
rect -242 -508 -214 -480
rect -166 -508 -138 -480
rect -90 -508 -62 -480
rect -14 -508 14 -480
rect 62 -508 90 -480
rect 138 -508 166 -480
rect 214 -508 242 -480
rect -242 -584 -214 -556
rect -166 -584 -138 -556
rect -90 -584 -62 -556
rect -14 -584 14 -556
rect 62 -584 90 -556
rect 138 -584 166 -556
rect 214 -584 242 -556
rect -242 -660 -214 -632
rect -166 -660 -138 -632
rect -90 -660 -62 -632
rect -14 -660 14 -632
rect 62 -660 90 -632
rect 138 -660 166 -632
rect 214 -660 242 -632
<< metal3 >>
rect -247 660 247 665
rect -247 632 -242 660
rect -214 632 -166 660
rect -138 632 -90 660
rect -62 632 -14 660
rect 14 632 62 660
rect 90 632 138 660
rect 166 632 214 660
rect 242 632 247 660
rect -247 584 247 632
rect -247 556 -242 584
rect -214 556 -166 584
rect -138 556 -90 584
rect -62 556 -14 584
rect 14 556 62 584
rect 90 556 138 584
rect 166 556 214 584
rect 242 556 247 584
rect -247 508 247 556
rect -247 480 -242 508
rect -214 480 -166 508
rect -138 480 -90 508
rect -62 480 -14 508
rect 14 480 62 508
rect 90 480 138 508
rect 166 480 214 508
rect 242 480 247 508
rect -247 432 247 480
rect -247 404 -242 432
rect -214 404 -166 432
rect -138 404 -90 432
rect -62 404 -14 432
rect 14 404 62 432
rect 90 404 138 432
rect 166 404 214 432
rect 242 404 247 432
rect -247 356 247 404
rect -247 328 -242 356
rect -214 328 -166 356
rect -138 328 -90 356
rect -62 328 -14 356
rect 14 328 62 356
rect 90 328 138 356
rect 166 328 214 356
rect 242 328 247 356
rect -247 280 247 328
rect -247 252 -242 280
rect -214 252 -166 280
rect -138 252 -90 280
rect -62 252 -14 280
rect 14 252 62 280
rect 90 252 138 280
rect 166 252 214 280
rect 242 252 247 280
rect -247 204 247 252
rect -247 176 -242 204
rect -214 176 -166 204
rect -138 176 -90 204
rect -62 176 -14 204
rect 14 176 62 204
rect 90 176 138 204
rect 166 176 214 204
rect 242 176 247 204
rect -247 128 247 176
rect -247 100 -242 128
rect -214 100 -166 128
rect -138 100 -90 128
rect -62 100 -14 128
rect 14 100 62 128
rect 90 100 138 128
rect 166 100 214 128
rect 242 100 247 128
rect -247 52 247 100
rect -247 24 -242 52
rect -214 24 -166 52
rect -138 24 -90 52
rect -62 24 -14 52
rect 14 24 62 52
rect 90 24 138 52
rect 166 24 214 52
rect 242 24 247 52
rect -247 -24 247 24
rect -247 -52 -242 -24
rect -214 -52 -166 -24
rect -138 -52 -90 -24
rect -62 -52 -14 -24
rect 14 -52 62 -24
rect 90 -52 138 -24
rect 166 -52 214 -24
rect 242 -52 247 -24
rect -247 -100 247 -52
rect -247 -128 -242 -100
rect -214 -128 -166 -100
rect -138 -128 -90 -100
rect -62 -128 -14 -100
rect 14 -128 62 -100
rect 90 -128 138 -100
rect 166 -128 214 -100
rect 242 -128 247 -100
rect -247 -176 247 -128
rect -247 -204 -242 -176
rect -214 -204 -166 -176
rect -138 -204 -90 -176
rect -62 -204 -14 -176
rect 14 -204 62 -176
rect 90 -204 138 -176
rect 166 -204 214 -176
rect 242 -204 247 -176
rect -247 -252 247 -204
rect -247 -280 -242 -252
rect -214 -280 -166 -252
rect -138 -280 -90 -252
rect -62 -280 -14 -252
rect 14 -280 62 -252
rect 90 -280 138 -252
rect 166 -280 214 -252
rect 242 -280 247 -252
rect -247 -328 247 -280
rect -247 -356 -242 -328
rect -214 -356 -166 -328
rect -138 -356 -90 -328
rect -62 -356 -14 -328
rect 14 -356 62 -328
rect 90 -356 138 -328
rect 166 -356 214 -328
rect 242 -356 247 -328
rect -247 -404 247 -356
rect -247 -432 -242 -404
rect -214 -432 -166 -404
rect -138 -432 -90 -404
rect -62 -432 -14 -404
rect 14 -432 62 -404
rect 90 -432 138 -404
rect 166 -432 214 -404
rect 242 -432 247 -404
rect -247 -480 247 -432
rect -247 -508 -242 -480
rect -214 -508 -166 -480
rect -138 -508 -90 -480
rect -62 -508 -14 -480
rect 14 -508 62 -480
rect 90 -508 138 -480
rect 166 -508 214 -480
rect 242 -508 247 -480
rect -247 -556 247 -508
rect -247 -584 -242 -556
rect -214 -584 -166 -556
rect -138 -584 -90 -556
rect -62 -584 -14 -556
rect 14 -584 62 -556
rect 90 -584 138 -556
rect 166 -584 214 -556
rect 242 -584 247 -556
rect -247 -632 247 -584
rect -247 -660 -242 -632
rect -214 -660 -166 -632
rect -138 -660 -90 -632
rect -62 -660 -14 -632
rect 14 -660 62 -632
rect 90 -660 138 -632
rect 166 -660 214 -632
rect 242 -660 247 -632
rect -247 -665 247 -660
<< end >>
