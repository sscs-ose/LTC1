magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1437 -1019 1437 1019
<< metal2 >>
rect -437 14 437 19
rect -437 -14 -432 14
rect -404 -14 -356 14
rect -328 -14 -280 14
rect -252 -14 -204 14
rect -176 -14 -128 14
rect -100 -14 -52 14
rect -24 -14 24 14
rect 52 -14 100 14
rect 128 -14 176 14
rect 204 -14 252 14
rect 280 -14 328 14
rect 356 -14 404 14
rect 432 -14 437 14
rect -437 -19 437 -14
<< via2 >>
rect -432 -14 -404 14
rect -356 -14 -328 14
rect -280 -14 -252 14
rect -204 -14 -176 14
rect -128 -14 -100 14
rect -52 -14 -24 14
rect 24 -14 52 14
rect 100 -14 128 14
rect 176 -14 204 14
rect 252 -14 280 14
rect 328 -14 356 14
rect 404 -14 432 14
<< metal3 >>
rect -437 14 437 19
rect -437 -14 -432 14
rect -404 -14 -356 14
rect -328 -14 -280 14
rect -252 -14 -204 14
rect -176 -14 -128 14
rect -100 -14 -52 14
rect -24 -14 24 14
rect 52 -14 100 14
rect 128 -14 176 14
rect 204 -14 252 14
rect 280 -14 328 14
rect 356 -14 404 14
rect 432 -14 437 14
rect -437 -19 437 -14
<< end >>
