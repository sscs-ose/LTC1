** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/untitled-15.sch
**.subckt untitled-15
I0 VDD ITAIL 2.5u
V1 VSS GND 0
.save i(v1)
V2 VDD GND 3.3
.save i(v2)
R1 VDD OUT1 2k m=1
x1 OUT1 ITAIL VSS net1 net2 net3 net4 pex_CM_LSB
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_CM_LSB.spice
.option savecurrents
.control
save all
op

tran 10n 3.2u
plot v(OUT1)
write LSB_TB.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
