magic
tech gf180mcuC
magscale 1 10
timestamp 1714126786
<< metal1 >>
rect -20077 6778 -19597 6870
rect -20077 6588 -19961 6778
rect -19741 6588 -19597 6778
rect -20077 6500 -19597 6588
rect -12620 -38786 -12140 -38694
rect -12620 -38976 -12504 -38786
rect -12284 -38976 -12140 -38786
rect -12620 -39064 -12140 -38976
<< via1 >>
rect -19961 6588 -19741 6778
rect -12504 -38976 -12284 -38786
<< metal2 >>
rect -20077 6782 -19597 6870
rect -20077 6578 -19990 6782
rect -19729 6578 -19597 6782
rect -20077 6500 -19597 6578
rect -12620 -38782 -12140 -38694
rect -12620 -38986 -12533 -38782
rect -12272 -38986 -12140 -38782
rect -12620 -39064 -12140 -38986
<< via2 >>
rect -19990 6778 -19729 6782
rect -19990 6588 -19961 6778
rect -19961 6588 -19741 6778
rect -19741 6588 -19729 6778
rect -19990 6578 -19729 6588
rect -12533 -38786 -12272 -38782
rect -12533 -38976 -12504 -38786
rect -12504 -38976 -12284 -38786
rect -12284 -38976 -12272 -38786
rect -12533 -38986 -12272 -38976
<< metal3 >>
rect -20077 6816 -19597 6870
rect -20077 6542 -20020 6816
rect -19666 6542 -19597 6816
rect -20077 6500 -19597 6542
rect -12620 -38748 -12140 -38694
rect -12620 -39022 -12563 -38748
rect -12209 -39022 -12140 -38748
rect -12620 -39064 -12140 -39022
<< via3 >>
rect -20020 6782 -19666 6816
rect -20020 6578 -19990 6782
rect -19990 6578 -19729 6782
rect -19729 6578 -19666 6782
rect -20020 6542 -19666 6578
rect -12563 -38782 -12209 -38748
rect -12563 -38986 -12533 -38782
rect -12533 -38986 -12272 -38782
rect -12272 -38986 -12209 -38782
rect -12563 -39022 -12209 -38986
<< metal4 >>
rect -20077 6845 -19597 6870
rect -20077 6527 -20038 6845
rect -19642 6527 -19597 6845
rect -20077 6500 -19597 6527
rect -12620 -38719 -12140 -38694
rect -12620 -39037 -12581 -38719
rect -12185 -39037 -12140 -38719
rect -12620 -39064 -12140 -39037
<< via4 >>
rect -20038 6816 -19642 6845
rect -20038 6542 -20020 6816
rect -20020 6542 -19666 6816
rect -19666 6542 -19642 6816
rect -20038 6527 -19642 6542
rect -12581 -38748 -12185 -38719
rect -12581 -39022 -12563 -38748
rect -12563 -39022 -12209 -38748
rect -12209 -39022 -12185 -38748
rect -12581 -39037 -12185 -39022
<< metal5 >>
rect -20077 6845 -19597 6870
rect -20077 6527 -20038 6845
rect -19642 6527 -19597 6845
rect -20077 6500 -19597 6527
rect -20011 5766 -19639 6500
rect -36784 5606 2723 5766
rect -36784 5394 2726 5606
rect -36784 5088 -36572 5394
rect -31170 5088 -30958 5394
rect -25556 5088 -25344 5394
rect -19942 5088 -19730 5394
rect -14328 5088 -14116 5394
rect -8714 5088 -8502 5394
rect -3100 5088 -2888 5394
rect 2514 5088 2726 5394
rect -34030 -37845 -33818 -37423
rect -28331 -37497 -28204 -37453
rect -28413 -37845 -28204 -37497
rect -22802 -37845 -22593 -37575
rect -17187 -37845 -16978 -37565
rect -12507 -37845 -12298 -37844
rect -11574 -37845 -11365 -37568
rect -5959 -37845 -5750 -37560
rect -346 -37845 -137 -37562
rect 5270 -37845 5479 -37571
rect -34030 -38054 5479 -37845
rect -34030 -38177 5457 -38054
rect -12507 -38694 -12298 -38177
rect -12620 -38719 -12140 -38694
rect -12620 -39037 -12581 -38719
rect -12185 -39037 -12140 -38719
rect -12620 -39064 -12140 -39037
use mim_2p0fF_Q67PCK  mim_2p0fF_Q67PCK_0
timestamp 1714046564
transform 1 0 -16909 0 1 -16140
box -22389 -21440 22389 21440
<< labels >>
flabel via4 -12407 -38891 -12407 -38891 0 FreeSans 1280 0 0 0 N
port 1 nsew
flabel via4 -19855 6679 -19855 6679 0 FreeSans 1280 0 0 0 P
port 0 nsew
<< end >>
