magic
tech gf180mcuC
magscale 1 10
timestamp 1692680230
<< pwell >>
rect -700 -1340 700 1340
<< nmos >>
rect -588 872 -532 1272
rect -428 872 -372 1272
rect -268 872 -212 1272
rect -108 872 -52 1272
rect 52 872 108 1272
rect 212 872 268 1272
rect 372 872 428 1272
rect 532 872 588 1272
rect -588 336 -532 736
rect -428 336 -372 736
rect -268 336 -212 736
rect -108 336 -52 736
rect 52 336 108 736
rect 212 336 268 736
rect 372 336 428 736
rect 532 336 588 736
rect -588 -200 -532 200
rect -428 -200 -372 200
rect -268 -200 -212 200
rect -108 -200 -52 200
rect 52 -200 108 200
rect 212 -200 268 200
rect 372 -200 428 200
rect 532 -200 588 200
rect -588 -736 -532 -336
rect -428 -736 -372 -336
rect -268 -736 -212 -336
rect -108 -736 -52 -336
rect 52 -736 108 -336
rect 212 -736 268 -336
rect 372 -736 428 -336
rect 532 -736 588 -336
rect -588 -1272 -532 -872
rect -428 -1272 -372 -872
rect -268 -1272 -212 -872
rect -108 -1272 -52 -872
rect 52 -1272 108 -872
rect 212 -1272 268 -872
rect 372 -1272 428 -872
rect 532 -1272 588 -872
<< ndiff >>
rect -676 1259 -588 1272
rect -676 885 -663 1259
rect -617 885 -588 1259
rect -676 872 -588 885
rect -532 1259 -428 1272
rect -532 885 -503 1259
rect -457 885 -428 1259
rect -532 872 -428 885
rect -372 1259 -268 1272
rect -372 885 -343 1259
rect -297 885 -268 1259
rect -372 872 -268 885
rect -212 1259 -108 1272
rect -212 885 -183 1259
rect -137 885 -108 1259
rect -212 872 -108 885
rect -52 1259 52 1272
rect -52 885 -23 1259
rect 23 885 52 1259
rect -52 872 52 885
rect 108 1259 212 1272
rect 108 885 137 1259
rect 183 885 212 1259
rect 108 872 212 885
rect 268 1259 372 1272
rect 268 885 297 1259
rect 343 885 372 1259
rect 268 872 372 885
rect 428 1259 532 1272
rect 428 885 457 1259
rect 503 885 532 1259
rect 428 872 532 885
rect 588 1259 676 1272
rect 588 885 617 1259
rect 663 885 676 1259
rect 588 872 676 885
rect -676 723 -588 736
rect -676 349 -663 723
rect -617 349 -588 723
rect -676 336 -588 349
rect -532 723 -428 736
rect -532 349 -503 723
rect -457 349 -428 723
rect -532 336 -428 349
rect -372 723 -268 736
rect -372 349 -343 723
rect -297 349 -268 723
rect -372 336 -268 349
rect -212 723 -108 736
rect -212 349 -183 723
rect -137 349 -108 723
rect -212 336 -108 349
rect -52 723 52 736
rect -52 349 -23 723
rect 23 349 52 723
rect -52 336 52 349
rect 108 723 212 736
rect 108 349 137 723
rect 183 349 212 723
rect 108 336 212 349
rect 268 723 372 736
rect 268 349 297 723
rect 343 349 372 723
rect 268 336 372 349
rect 428 723 532 736
rect 428 349 457 723
rect 503 349 532 723
rect 428 336 532 349
rect 588 723 676 736
rect 588 349 617 723
rect 663 349 676 723
rect 588 336 676 349
rect -676 187 -588 200
rect -676 -187 -663 187
rect -617 -187 -588 187
rect -676 -200 -588 -187
rect -532 187 -428 200
rect -532 -187 -503 187
rect -457 -187 -428 187
rect -532 -200 -428 -187
rect -372 187 -268 200
rect -372 -187 -343 187
rect -297 -187 -268 187
rect -372 -200 -268 -187
rect -212 187 -108 200
rect -212 -187 -183 187
rect -137 -187 -108 187
rect -212 -200 -108 -187
rect -52 187 52 200
rect -52 -187 -23 187
rect 23 -187 52 187
rect -52 -200 52 -187
rect 108 187 212 200
rect 108 -187 137 187
rect 183 -187 212 187
rect 108 -200 212 -187
rect 268 187 372 200
rect 268 -187 297 187
rect 343 -187 372 187
rect 268 -200 372 -187
rect 428 187 532 200
rect 428 -187 457 187
rect 503 -187 532 187
rect 428 -200 532 -187
rect 588 187 676 200
rect 588 -187 617 187
rect 663 -187 676 187
rect 588 -200 676 -187
rect -676 -349 -588 -336
rect -676 -723 -663 -349
rect -617 -723 -588 -349
rect -676 -736 -588 -723
rect -532 -349 -428 -336
rect -532 -723 -503 -349
rect -457 -723 -428 -349
rect -532 -736 -428 -723
rect -372 -349 -268 -336
rect -372 -723 -343 -349
rect -297 -723 -268 -349
rect -372 -736 -268 -723
rect -212 -349 -108 -336
rect -212 -723 -183 -349
rect -137 -723 -108 -349
rect -212 -736 -108 -723
rect -52 -349 52 -336
rect -52 -723 -23 -349
rect 23 -723 52 -349
rect -52 -736 52 -723
rect 108 -349 212 -336
rect 108 -723 137 -349
rect 183 -723 212 -349
rect 108 -736 212 -723
rect 268 -349 372 -336
rect 268 -723 297 -349
rect 343 -723 372 -349
rect 268 -736 372 -723
rect 428 -349 532 -336
rect 428 -723 457 -349
rect 503 -723 532 -349
rect 428 -736 532 -723
rect 588 -349 676 -336
rect 588 -723 617 -349
rect 663 -723 676 -349
rect 588 -736 676 -723
rect -676 -885 -588 -872
rect -676 -1259 -663 -885
rect -617 -1259 -588 -885
rect -676 -1272 -588 -1259
rect -532 -885 -428 -872
rect -532 -1259 -503 -885
rect -457 -1259 -428 -885
rect -532 -1272 -428 -1259
rect -372 -885 -268 -872
rect -372 -1259 -343 -885
rect -297 -1259 -268 -885
rect -372 -1272 -268 -1259
rect -212 -885 -108 -872
rect -212 -1259 -183 -885
rect -137 -1259 -108 -885
rect -212 -1272 -108 -1259
rect -52 -885 52 -872
rect -52 -1259 -23 -885
rect 23 -1259 52 -885
rect -52 -1272 52 -1259
rect 108 -885 212 -872
rect 108 -1259 137 -885
rect 183 -1259 212 -885
rect 108 -1272 212 -1259
rect 268 -885 372 -872
rect 268 -1259 297 -885
rect 343 -1259 372 -885
rect 268 -1272 372 -1259
rect 428 -885 532 -872
rect 428 -1259 457 -885
rect 503 -1259 532 -885
rect 428 -1272 532 -1259
rect 588 -885 676 -872
rect 588 -1259 617 -885
rect 663 -1259 676 -885
rect 588 -1272 676 -1259
<< ndiffc >>
rect -663 885 -617 1259
rect -503 885 -457 1259
rect -343 885 -297 1259
rect -183 885 -137 1259
rect -23 885 23 1259
rect 137 885 183 1259
rect 297 885 343 1259
rect 457 885 503 1259
rect 617 885 663 1259
rect -663 349 -617 723
rect -503 349 -457 723
rect -343 349 -297 723
rect -183 349 -137 723
rect -23 349 23 723
rect 137 349 183 723
rect 297 349 343 723
rect 457 349 503 723
rect 617 349 663 723
rect -663 -187 -617 187
rect -503 -187 -457 187
rect -343 -187 -297 187
rect -183 -187 -137 187
rect -23 -187 23 187
rect 137 -187 183 187
rect 297 -187 343 187
rect 457 -187 503 187
rect 617 -187 663 187
rect -663 -723 -617 -349
rect -503 -723 -457 -349
rect -343 -723 -297 -349
rect -183 -723 -137 -349
rect -23 -723 23 -349
rect 137 -723 183 -349
rect 297 -723 343 -349
rect 457 -723 503 -349
rect 617 -723 663 -349
rect -663 -1259 -617 -885
rect -503 -1259 -457 -885
rect -343 -1259 -297 -885
rect -183 -1259 -137 -885
rect -23 -1259 23 -885
rect 137 -1259 183 -885
rect 297 -1259 343 -885
rect 457 -1259 503 -885
rect 617 -1259 663 -885
<< polysilicon >>
rect -588 1272 -532 1316
rect -428 1272 -372 1316
rect -268 1272 -212 1316
rect -108 1272 -52 1316
rect 52 1272 108 1316
rect 212 1272 268 1316
rect 372 1272 428 1316
rect 532 1272 588 1316
rect -588 828 -532 872
rect -428 828 -372 872
rect -268 828 -212 872
rect -108 828 -52 872
rect 52 828 108 872
rect 212 828 268 872
rect 372 828 428 872
rect 532 828 588 872
rect -588 736 -532 780
rect -428 736 -372 780
rect -268 736 -212 780
rect -108 736 -52 780
rect 52 736 108 780
rect 212 736 268 780
rect 372 736 428 780
rect 532 736 588 780
rect -588 292 -532 336
rect -428 292 -372 336
rect -268 292 -212 336
rect -108 292 -52 336
rect 52 292 108 336
rect 212 292 268 336
rect 372 292 428 336
rect 532 292 588 336
rect -588 200 -532 244
rect -428 200 -372 244
rect -268 200 -212 244
rect -108 200 -52 244
rect 52 200 108 244
rect 212 200 268 244
rect 372 200 428 244
rect 532 200 588 244
rect -588 -244 -532 -200
rect -428 -244 -372 -200
rect -268 -244 -212 -200
rect -108 -244 -52 -200
rect 52 -244 108 -200
rect 212 -244 268 -200
rect 372 -244 428 -200
rect 532 -244 588 -200
rect -588 -336 -532 -292
rect -428 -336 -372 -292
rect -268 -336 -212 -292
rect -108 -336 -52 -292
rect 52 -336 108 -292
rect 212 -336 268 -292
rect 372 -336 428 -292
rect 532 -336 588 -292
rect -588 -780 -532 -736
rect -428 -780 -372 -736
rect -268 -780 -212 -736
rect -108 -780 -52 -736
rect 52 -780 108 -736
rect 212 -780 268 -736
rect 372 -780 428 -736
rect 532 -780 588 -736
rect -588 -872 -532 -828
rect -428 -872 -372 -828
rect -268 -872 -212 -828
rect -108 -872 -52 -828
rect 52 -872 108 -828
rect 212 -872 268 -828
rect 372 -872 428 -828
rect 532 -872 588 -828
rect -588 -1316 -532 -1272
rect -428 -1316 -372 -1272
rect -268 -1316 -212 -1272
rect -108 -1316 -52 -1272
rect 52 -1316 108 -1272
rect 212 -1316 268 -1272
rect 372 -1316 428 -1272
rect 532 -1316 588 -1272
<< metal1 >>
rect -663 1259 -617 1270
rect -663 874 -617 885
rect -503 1259 -457 1270
rect -503 874 -457 885
rect -343 1259 -297 1270
rect -343 874 -297 885
rect -183 1259 -137 1270
rect -183 874 -137 885
rect -23 1259 23 1270
rect -23 874 23 885
rect 137 1259 183 1270
rect 137 874 183 885
rect 297 1259 343 1270
rect 297 874 343 885
rect 457 1259 503 1270
rect 457 874 503 885
rect 617 1259 663 1270
rect 617 874 663 885
rect -663 723 -617 734
rect -663 338 -617 349
rect -503 723 -457 734
rect -503 338 -457 349
rect -343 723 -297 734
rect -343 338 -297 349
rect -183 723 -137 734
rect -183 338 -137 349
rect -23 723 23 734
rect -23 338 23 349
rect 137 723 183 734
rect 137 338 183 349
rect 297 723 343 734
rect 297 338 343 349
rect 457 723 503 734
rect 457 338 503 349
rect 617 723 663 734
rect 617 338 663 349
rect -663 187 -617 198
rect -663 -198 -617 -187
rect -503 187 -457 198
rect -503 -198 -457 -187
rect -343 187 -297 198
rect -343 -198 -297 -187
rect -183 187 -137 198
rect -183 -198 -137 -187
rect -23 187 23 198
rect -23 -198 23 -187
rect 137 187 183 198
rect 137 -198 183 -187
rect 297 187 343 198
rect 297 -198 343 -187
rect 457 187 503 198
rect 457 -198 503 -187
rect 617 187 663 198
rect 617 -198 663 -187
rect -663 -349 -617 -338
rect -663 -734 -617 -723
rect -503 -349 -457 -338
rect -503 -734 -457 -723
rect -343 -349 -297 -338
rect -343 -734 -297 -723
rect -183 -349 -137 -338
rect -183 -734 -137 -723
rect -23 -349 23 -338
rect -23 -734 23 -723
rect 137 -349 183 -338
rect 137 -734 183 -723
rect 297 -349 343 -338
rect 297 -734 343 -723
rect 457 -349 503 -338
rect 457 -734 503 -723
rect 617 -349 663 -338
rect 617 -734 663 -723
rect -663 -885 -617 -874
rect -663 -1270 -617 -1259
rect -503 -885 -457 -874
rect -503 -1270 -457 -1259
rect -343 -885 -297 -874
rect -343 -1270 -297 -1259
rect -183 -885 -137 -874
rect -183 -1270 -137 -1259
rect -23 -885 23 -874
rect -23 -1270 23 -1259
rect 137 -885 183 -874
rect 137 -1270 183 -1259
rect 297 -885 343 -874
rect 297 -1270 343 -1259
rect 457 -885 503 -874
rect 457 -1270 503 -1259
rect 617 -885 663 -874
rect 617 -1270 663 -1259
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 2.0 l 0.280 m 5 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
