magic
tech gf180mcuC
magscale 1 10
timestamp 1690963719
<< pwell >>
rect -860 -504 860 504
<< nmos >>
rect -748 236 -692 436
rect -588 236 -532 436
rect -428 236 -372 436
rect -268 236 -212 436
rect -108 236 -52 436
rect 52 236 108 436
rect 212 236 268 436
rect 372 236 428 436
rect 532 236 588 436
rect 692 236 748 436
rect -748 -100 -692 100
rect -588 -100 -532 100
rect -428 -100 -372 100
rect -268 -100 -212 100
rect -108 -100 -52 100
rect 52 -100 108 100
rect 212 -100 268 100
rect 372 -100 428 100
rect 532 -100 588 100
rect 692 -100 748 100
rect -748 -436 -692 -236
rect -588 -436 -532 -236
rect -428 -436 -372 -236
rect -268 -436 -212 -236
rect -108 -436 -52 -236
rect 52 -436 108 -236
rect 212 -436 268 -236
rect 372 -436 428 -236
rect 532 -436 588 -236
rect 692 -436 748 -236
<< ndiff >>
rect -836 423 -748 436
rect -836 249 -823 423
rect -777 249 -748 423
rect -836 236 -748 249
rect -692 423 -588 436
rect -692 249 -663 423
rect -617 249 -588 423
rect -692 236 -588 249
rect -532 423 -428 436
rect -532 249 -503 423
rect -457 249 -428 423
rect -532 236 -428 249
rect -372 423 -268 436
rect -372 249 -343 423
rect -297 249 -268 423
rect -372 236 -268 249
rect -212 423 -108 436
rect -212 249 -183 423
rect -137 249 -108 423
rect -212 236 -108 249
rect -52 423 52 436
rect -52 249 -23 423
rect 23 249 52 423
rect -52 236 52 249
rect 108 423 212 436
rect 108 249 137 423
rect 183 249 212 423
rect 108 236 212 249
rect 268 423 372 436
rect 268 249 297 423
rect 343 249 372 423
rect 268 236 372 249
rect 428 423 532 436
rect 428 249 457 423
rect 503 249 532 423
rect 428 236 532 249
rect 588 423 692 436
rect 588 249 617 423
rect 663 249 692 423
rect 588 236 692 249
rect 748 423 836 436
rect 748 249 777 423
rect 823 249 836 423
rect 748 236 836 249
rect -836 87 -748 100
rect -836 -87 -823 87
rect -777 -87 -748 87
rect -836 -100 -748 -87
rect -692 87 -588 100
rect -692 -87 -663 87
rect -617 -87 -588 87
rect -692 -100 -588 -87
rect -532 87 -428 100
rect -532 -87 -503 87
rect -457 -87 -428 87
rect -532 -100 -428 -87
rect -372 87 -268 100
rect -372 -87 -343 87
rect -297 -87 -268 87
rect -372 -100 -268 -87
rect -212 87 -108 100
rect -212 -87 -183 87
rect -137 -87 -108 87
rect -212 -100 -108 -87
rect -52 87 52 100
rect -52 -87 -23 87
rect 23 -87 52 87
rect -52 -100 52 -87
rect 108 87 212 100
rect 108 -87 137 87
rect 183 -87 212 87
rect 108 -100 212 -87
rect 268 87 372 100
rect 268 -87 297 87
rect 343 -87 372 87
rect 268 -100 372 -87
rect 428 87 532 100
rect 428 -87 457 87
rect 503 -87 532 87
rect 428 -100 532 -87
rect 588 87 692 100
rect 588 -87 617 87
rect 663 -87 692 87
rect 588 -100 692 -87
rect 748 87 836 100
rect 748 -87 777 87
rect 823 -87 836 87
rect 748 -100 836 -87
rect -836 -249 -748 -236
rect -836 -423 -823 -249
rect -777 -423 -748 -249
rect -836 -436 -748 -423
rect -692 -249 -588 -236
rect -692 -423 -663 -249
rect -617 -423 -588 -249
rect -692 -436 -588 -423
rect -532 -249 -428 -236
rect -532 -423 -503 -249
rect -457 -423 -428 -249
rect -532 -436 -428 -423
rect -372 -249 -268 -236
rect -372 -423 -343 -249
rect -297 -423 -268 -249
rect -372 -436 -268 -423
rect -212 -249 -108 -236
rect -212 -423 -183 -249
rect -137 -423 -108 -249
rect -212 -436 -108 -423
rect -52 -249 52 -236
rect -52 -423 -23 -249
rect 23 -423 52 -249
rect -52 -436 52 -423
rect 108 -249 212 -236
rect 108 -423 137 -249
rect 183 -423 212 -249
rect 108 -436 212 -423
rect 268 -249 372 -236
rect 268 -423 297 -249
rect 343 -423 372 -249
rect 268 -436 372 -423
rect 428 -249 532 -236
rect 428 -423 457 -249
rect 503 -423 532 -249
rect 428 -436 532 -423
rect 588 -249 692 -236
rect 588 -423 617 -249
rect 663 -423 692 -249
rect 588 -436 692 -423
rect 748 -249 836 -236
rect 748 -423 777 -249
rect 823 -423 836 -249
rect 748 -436 836 -423
<< ndiffc >>
rect -823 249 -777 423
rect -663 249 -617 423
rect -503 249 -457 423
rect -343 249 -297 423
rect -183 249 -137 423
rect -23 249 23 423
rect 137 249 183 423
rect 297 249 343 423
rect 457 249 503 423
rect 617 249 663 423
rect 777 249 823 423
rect -823 -87 -777 87
rect -663 -87 -617 87
rect -503 -87 -457 87
rect -343 -87 -297 87
rect -183 -87 -137 87
rect -23 -87 23 87
rect 137 -87 183 87
rect 297 -87 343 87
rect 457 -87 503 87
rect 617 -87 663 87
rect 777 -87 823 87
rect -823 -423 -777 -249
rect -663 -423 -617 -249
rect -503 -423 -457 -249
rect -343 -423 -297 -249
rect -183 -423 -137 -249
rect -23 -423 23 -249
rect 137 -423 183 -249
rect 297 -423 343 -249
rect 457 -423 503 -249
rect 617 -423 663 -249
rect 777 -423 823 -249
<< polysilicon >>
rect -748 436 -692 480
rect -588 436 -532 480
rect -428 436 -372 480
rect -268 436 -212 480
rect -108 436 -52 480
rect 52 436 108 480
rect 212 436 268 480
rect 372 436 428 480
rect 532 436 588 480
rect 692 436 748 480
rect -748 192 -692 236
rect -588 192 -532 236
rect -428 192 -372 236
rect -268 192 -212 236
rect -108 192 -52 236
rect 52 192 108 236
rect 212 192 268 236
rect 372 192 428 236
rect 532 192 588 236
rect 692 192 748 236
rect -748 100 -692 144
rect -588 100 -532 144
rect -428 100 -372 144
rect -268 100 -212 144
rect -108 100 -52 144
rect 52 100 108 144
rect 212 100 268 144
rect 372 100 428 144
rect 532 100 588 144
rect 692 100 748 144
rect -748 -144 -692 -100
rect -588 -144 -532 -100
rect -428 -144 -372 -100
rect -268 -144 -212 -100
rect -108 -144 -52 -100
rect 52 -144 108 -100
rect 212 -144 268 -100
rect 372 -144 428 -100
rect 532 -144 588 -100
rect 692 -144 748 -100
rect -748 -236 -692 -192
rect -588 -236 -532 -192
rect -428 -236 -372 -192
rect -268 -236 -212 -192
rect -108 -236 -52 -192
rect 52 -236 108 -192
rect 212 -236 268 -192
rect 372 -236 428 -192
rect 532 -236 588 -192
rect 692 -236 748 -192
rect -748 -480 -692 -436
rect -588 -480 -532 -436
rect -428 -480 -372 -436
rect -268 -480 -212 -436
rect -108 -480 -52 -436
rect 52 -480 108 -436
rect 212 -480 268 -436
rect 372 -480 428 -436
rect 532 -480 588 -436
rect 692 -480 748 -436
<< metal1 >>
rect -823 423 -777 434
rect -823 238 -777 249
rect -663 423 -617 434
rect -663 238 -617 249
rect -503 423 -457 434
rect -503 238 -457 249
rect -343 423 -297 434
rect -343 238 -297 249
rect -183 423 -137 434
rect -183 238 -137 249
rect -23 423 23 434
rect -23 238 23 249
rect 137 423 183 434
rect 137 238 183 249
rect 297 423 343 434
rect 297 238 343 249
rect 457 423 503 434
rect 457 238 503 249
rect 617 423 663 434
rect 617 238 663 249
rect 777 423 823 434
rect 777 238 823 249
rect -823 87 -777 98
rect -823 -98 -777 -87
rect -663 87 -617 98
rect -663 -98 -617 -87
rect -503 87 -457 98
rect -503 -98 -457 -87
rect -343 87 -297 98
rect -343 -98 -297 -87
rect -183 87 -137 98
rect -183 -98 -137 -87
rect -23 87 23 98
rect -23 -98 23 -87
rect 137 87 183 98
rect 137 -98 183 -87
rect 297 87 343 98
rect 297 -98 343 -87
rect 457 87 503 98
rect 457 -98 503 -87
rect 617 87 663 98
rect 617 -98 663 -87
rect 777 87 823 98
rect 777 -98 823 -87
rect -823 -249 -777 -238
rect -823 -434 -777 -423
rect -663 -249 -617 -238
rect -663 -434 -617 -423
rect -503 -249 -457 -238
rect -503 -434 -457 -423
rect -343 -249 -297 -238
rect -343 -434 -297 -423
rect -183 -249 -137 -238
rect -183 -434 -137 -423
rect -23 -249 23 -238
rect -23 -434 23 -423
rect 137 -249 183 -238
rect 137 -434 183 -423
rect 297 -249 343 -238
rect 297 -434 343 -423
rect 457 -249 503 -238
rect 457 -434 503 -423
rect 617 -249 663 -238
rect 617 -434 663 -423
rect 777 -249 823 -238
rect 777 -434 823 -423
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1 l 0.280 m 3 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
