magic
tech gf180mcuC
magscale 1 10
timestamp 1692688075
<< nwell >>
rect -1270 60 5529 271
rect -2639 5 5529 60
rect -2374 -36 -2311 5
rect -2174 -36 -2111 5
rect -1974 -36 -1911 5
rect -1774 -36 -1711 5
rect -1574 -36 -1511 5
rect -1374 -36 -1311 5
rect -1270 -72 5529 5
<< pwell >>
rect -1498 -993 -517 -680
rect 4061 -993 5664 -680
rect -2620 -1529 5664 -993
<< psubdiff >>
rect -2544 -1240 -2437 -1226
rect -2544 -1324 -2531 -1240
rect -2450 -1244 -2437 -1240
rect -2344 -1240 -2237 -1226
rect -2344 -1244 -2331 -1240
rect -2450 -1322 -2331 -1244
rect -2450 -1324 -2437 -1322
rect -2544 -1339 -2437 -1324
rect -2344 -1324 -2331 -1322
rect -2250 -1244 -2237 -1240
rect -2144 -1240 -2037 -1226
rect -2144 -1244 -2131 -1240
rect -2250 -1322 -2131 -1244
rect -2250 -1324 -2237 -1322
rect -2344 -1339 -2237 -1324
rect -2144 -1324 -2131 -1322
rect -2050 -1244 -2037 -1240
rect -1944 -1240 -1837 -1226
rect -1944 -1244 -1931 -1240
rect -2050 -1322 -1931 -1244
rect -2050 -1324 -2037 -1322
rect -2144 -1339 -2037 -1324
rect -1944 -1324 -1931 -1322
rect -1850 -1244 -1837 -1240
rect -1744 -1240 -1637 -1226
rect -1744 -1244 -1731 -1240
rect -1850 -1322 -1731 -1244
rect -1850 -1324 -1837 -1322
rect -1944 -1339 -1837 -1324
rect -1744 -1324 -1731 -1322
rect -1650 -1244 -1637 -1240
rect -1544 -1240 -1437 -1226
rect -1544 -1244 -1531 -1240
rect -1650 -1322 -1531 -1244
rect -1650 -1324 -1637 -1322
rect -1744 -1339 -1637 -1324
rect -1544 -1324 -1531 -1322
rect -1450 -1244 -1437 -1240
rect -1344 -1240 -1237 -1226
rect -1344 -1244 -1331 -1240
rect -1450 -1322 -1331 -1244
rect -1450 -1324 -1437 -1322
rect -1544 -1339 -1437 -1324
rect -1344 -1324 -1331 -1322
rect -1250 -1324 -1237 -1240
rect -1344 -1339 -1237 -1324
rect -1170 -1400 -1063 -1386
rect -1170 -1484 -1157 -1400
rect -1076 -1406 -1063 -1400
rect -970 -1400 -863 -1386
rect -970 -1406 -957 -1400
rect -1076 -1484 -957 -1406
rect -876 -1406 -863 -1400
rect -770 -1400 -663 -1386
rect -770 -1406 -757 -1400
rect -876 -1484 -757 -1406
rect -676 -1406 -663 -1400
rect -570 -1400 -463 -1386
rect -570 -1406 -557 -1400
rect -676 -1484 -557 -1406
rect -476 -1406 -463 -1400
rect -370 -1400 -263 -1386
rect -370 -1406 -357 -1400
rect -476 -1484 -357 -1406
rect -276 -1406 -263 -1400
rect -170 -1400 -63 -1386
rect -170 -1406 -157 -1400
rect -276 -1484 -157 -1406
rect -76 -1406 -63 -1400
rect 30 -1400 137 -1386
rect 30 -1406 43 -1400
rect -76 -1484 43 -1406
rect 124 -1484 137 -1400
rect -1170 -1499 -1063 -1484
rect -970 -1499 -863 -1484
rect -770 -1499 -663 -1484
rect -570 -1499 -463 -1484
rect -370 -1499 -263 -1484
rect -170 -1499 -63 -1484
rect 30 -1499 137 -1484
rect 255 -1400 362 -1386
rect 255 -1484 268 -1400
rect 349 -1404 362 -1400
rect 455 -1400 562 -1386
rect 455 -1404 468 -1400
rect 349 -1482 468 -1404
rect 349 -1484 362 -1482
rect 255 -1499 362 -1484
rect 455 -1484 468 -1482
rect 549 -1404 562 -1400
rect 655 -1400 762 -1386
rect 655 -1404 668 -1400
rect 549 -1482 668 -1404
rect 549 -1484 562 -1482
rect 455 -1499 562 -1484
rect 655 -1484 668 -1482
rect 749 -1404 762 -1400
rect 855 -1400 962 -1386
rect 855 -1404 868 -1400
rect 749 -1482 868 -1404
rect 749 -1484 762 -1482
rect 655 -1499 762 -1484
rect 855 -1484 868 -1482
rect 949 -1404 962 -1400
rect 1055 -1400 1162 -1386
rect 1055 -1404 1068 -1400
rect 949 -1482 1068 -1404
rect 949 -1484 962 -1482
rect 855 -1499 962 -1484
rect 1055 -1484 1068 -1482
rect 1149 -1404 1162 -1400
rect 1255 -1400 1362 -1386
rect 1255 -1404 1268 -1400
rect 1149 -1482 1268 -1404
rect 1149 -1484 1162 -1482
rect 1055 -1499 1162 -1484
rect 1255 -1484 1268 -1482
rect 1349 -1404 1362 -1400
rect 1455 -1400 1562 -1386
rect 1455 -1404 1468 -1400
rect 1349 -1482 1468 -1404
rect 1349 -1484 1362 -1482
rect 1255 -1499 1362 -1484
rect 1455 -1484 1468 -1482
rect 1549 -1484 1562 -1400
rect 1455 -1499 1562 -1484
rect 1680 -1400 1787 -1386
rect 1880 -1400 1987 -1386
rect 2080 -1400 2187 -1386
rect 2280 -1400 2387 -1386
rect 2480 -1400 2587 -1386
rect 2680 -1400 2787 -1386
rect 2880 -1400 2987 -1386
rect 1680 -1484 1693 -1400
rect 1774 -1478 1893 -1400
rect 1774 -1484 1787 -1478
rect 1680 -1499 1787 -1484
rect 1880 -1484 1893 -1478
rect 1974 -1478 2093 -1400
rect 1974 -1484 1987 -1478
rect 1880 -1499 1987 -1484
rect 2080 -1484 2093 -1478
rect 2174 -1478 2293 -1400
rect 2174 -1484 2187 -1478
rect 2080 -1499 2187 -1484
rect 2280 -1484 2293 -1478
rect 2374 -1478 2493 -1400
rect 2374 -1484 2387 -1478
rect 2280 -1499 2387 -1484
rect 2480 -1484 2493 -1478
rect 2574 -1478 2693 -1400
rect 2574 -1484 2587 -1478
rect 2480 -1499 2587 -1484
rect 2680 -1484 2693 -1478
rect 2774 -1478 2893 -1400
rect 2774 -1484 2787 -1478
rect 2680 -1499 2787 -1484
rect 2880 -1484 2893 -1478
rect 2974 -1484 2987 -1400
rect 2880 -1499 2987 -1484
rect 3105 -1400 3212 -1386
rect 3105 -1484 3118 -1400
rect 3199 -1408 3212 -1400
rect 3305 -1400 3412 -1386
rect 3305 -1408 3318 -1400
rect 3199 -1484 3318 -1408
rect 3399 -1408 3412 -1400
rect 3505 -1400 3612 -1386
rect 3505 -1408 3518 -1400
rect 3399 -1484 3518 -1408
rect 3599 -1408 3612 -1400
rect 3705 -1400 3812 -1386
rect 3705 -1408 3718 -1400
rect 3599 -1484 3718 -1408
rect 3799 -1408 3812 -1400
rect 3905 -1400 4012 -1386
rect 3905 -1408 3918 -1400
rect 3799 -1484 3918 -1408
rect 3999 -1408 4012 -1400
rect 4105 -1400 4212 -1386
rect 4105 -1408 4118 -1400
rect 3999 -1484 4118 -1408
rect 4199 -1408 4212 -1400
rect 4305 -1400 4412 -1386
rect 4305 -1408 4318 -1400
rect 4199 -1484 4318 -1408
rect 4399 -1404 4412 -1400
rect 4530 -1400 4637 -1386
rect 4530 -1404 4543 -1400
rect 4399 -1482 4543 -1404
rect 4399 -1484 4412 -1482
rect 3105 -1486 4412 -1484
rect 3105 -1499 3212 -1486
rect 3305 -1499 3412 -1486
rect 3505 -1499 3612 -1486
rect 3705 -1499 3812 -1486
rect 3905 -1499 4012 -1486
rect 4105 -1499 4212 -1486
rect 4305 -1499 4412 -1486
rect 4530 -1484 4543 -1482
rect 4624 -1404 4637 -1400
rect 4730 -1400 4837 -1386
rect 4730 -1404 4743 -1400
rect 4624 -1482 4743 -1404
rect 4624 -1484 4637 -1482
rect 4530 -1499 4637 -1484
rect 4730 -1484 4743 -1482
rect 4824 -1404 4837 -1400
rect 4930 -1400 5037 -1386
rect 4930 -1404 4943 -1400
rect 4824 -1482 4943 -1404
rect 4824 -1484 4837 -1482
rect 4730 -1499 4837 -1484
rect 4930 -1484 4943 -1482
rect 5024 -1404 5037 -1400
rect 5130 -1400 5237 -1386
rect 5130 -1404 5143 -1400
rect 5024 -1482 5143 -1404
rect 5024 -1484 5037 -1482
rect 4930 -1499 5037 -1484
rect 5130 -1484 5143 -1482
rect 5224 -1404 5237 -1400
rect 5330 -1400 5437 -1386
rect 5330 -1404 5343 -1400
rect 5224 -1482 5343 -1404
rect 5224 -1484 5237 -1482
rect 5130 -1499 5237 -1484
rect 5330 -1484 5343 -1482
rect 5424 -1404 5437 -1400
rect 5530 -1400 5637 -1386
rect 5530 -1404 5543 -1400
rect 5424 -1482 5543 -1404
rect 5424 -1484 5437 -1482
rect 5330 -1499 5437 -1484
rect 5530 -1484 5543 -1482
rect 5624 -1484 5637 -1400
rect 5530 -1499 5637 -1484
<< nsubdiff >>
rect -1230 233 119 247
rect -1230 175 -1205 233
rect -1142 175 -1005 233
rect -942 175 -805 233
rect -742 175 -605 233
rect -542 175 -405 233
rect -342 175 -205 233
rect -142 175 -5 233
rect 58 175 119 233
rect -1230 159 119 175
rect 195 233 1544 247
rect 195 175 220 233
rect 283 175 420 233
rect 483 175 620 233
rect 683 175 820 233
rect 883 175 1020 233
rect 1083 175 1220 233
rect 1283 175 1420 233
rect 1483 175 1544 233
rect 195 159 1544 175
rect 1620 233 2969 247
rect 1620 175 1645 233
rect 1708 175 1845 233
rect 1908 175 2045 233
rect 2108 175 2245 233
rect 2308 175 2445 233
rect 2508 175 2645 233
rect 2708 175 2845 233
rect 2908 175 2969 233
rect 1620 159 2969 175
rect 3045 233 4394 247
rect 3045 175 3070 233
rect 3133 175 3270 233
rect 3333 175 3470 233
rect 3533 175 3670 233
rect 3733 175 3870 233
rect 3933 175 4070 233
rect 4133 175 4270 233
rect 4333 175 4394 233
rect 3045 159 4394 175
rect 4470 233 5458 247
rect 4470 175 4495 233
rect 4558 175 4695 233
rect 4758 175 4895 233
rect 4958 175 5095 233
rect 5158 175 5295 233
rect 5358 175 5458 233
rect 4470 159 5458 175
rect -2599 22 -1250 36
rect -2599 -36 -2574 22
rect -2511 -36 -2374 22
rect -2311 -36 -2174 22
rect -2111 -36 -1974 22
rect -1911 -36 -1774 22
rect -1711 -36 -1574 22
rect -1511 -36 -1374 22
rect -1311 -36 -1250 22
rect -2599 -52 -1250 -36
<< psubdiffcont >>
rect -2531 -1324 -2450 -1240
rect -2331 -1324 -2250 -1240
rect -2131 -1324 -2050 -1240
rect -1931 -1324 -1850 -1240
rect -1731 -1324 -1650 -1240
rect -1531 -1324 -1450 -1240
rect -1331 -1324 -1250 -1240
rect -1157 -1484 -1076 -1400
rect -957 -1484 -876 -1400
rect -757 -1484 -676 -1400
rect -557 -1484 -476 -1400
rect -357 -1484 -276 -1400
rect -157 -1484 -76 -1400
rect 43 -1484 124 -1400
rect 268 -1484 349 -1400
rect 468 -1484 549 -1400
rect 668 -1484 749 -1400
rect 868 -1484 949 -1400
rect 1068 -1484 1149 -1400
rect 1268 -1484 1349 -1400
rect 1468 -1484 1549 -1400
rect 1693 -1484 1774 -1400
rect 1893 -1484 1974 -1400
rect 2093 -1484 2174 -1400
rect 2293 -1484 2374 -1400
rect 2493 -1484 2574 -1400
rect 2693 -1484 2774 -1400
rect 2893 -1484 2974 -1400
rect 3118 -1484 3199 -1400
rect 3318 -1484 3399 -1400
rect 3518 -1484 3599 -1400
rect 3718 -1484 3799 -1400
rect 3918 -1484 3999 -1400
rect 4118 -1484 4199 -1400
rect 4318 -1484 4399 -1400
rect 4543 -1484 4624 -1400
rect 4743 -1484 4824 -1400
rect 4943 -1484 5024 -1400
rect 5143 -1484 5224 -1400
rect 5343 -1484 5424 -1400
rect 5543 -1484 5624 -1400
<< nsubdiffcont >>
rect -1205 175 -1142 233
rect -1005 175 -942 233
rect -805 175 -742 233
rect -605 175 -542 233
rect -405 175 -342 233
rect -205 175 -142 233
rect -5 175 58 233
rect 220 175 283 233
rect 420 175 483 233
rect 620 175 683 233
rect 820 175 883 233
rect 1020 175 1083 233
rect 1220 175 1283 233
rect 1420 175 1483 233
rect 1645 175 1708 233
rect 1845 175 1908 233
rect 2045 175 2108 233
rect 2245 175 2308 233
rect 2445 175 2508 233
rect 2645 175 2708 233
rect 2845 175 2908 233
rect 3070 175 3133 233
rect 3270 175 3333 233
rect 3470 175 3533 233
rect 3670 175 3733 233
rect 3870 175 3933 233
rect 4070 175 4133 233
rect 4270 175 4333 233
rect 4495 175 4558 233
rect 4695 175 4758 233
rect 4895 175 4958 233
rect 5095 175 5158 233
rect 5295 175 5358 233
rect -2574 -36 -2511 22
rect -2374 -36 -2311 22
rect -2174 -36 -2111 22
rect -1974 -36 -1911 22
rect -1774 -36 -1711 22
rect -1574 -36 -1511 22
rect -1374 -36 -1311 22
<< polysilicon >>
rect -941 -101 5355 -48
rect -941 -129 -888 -101
rect -2631 -626 -2544 -613
rect -2631 -678 -2616 -626
rect -2564 -629 -2544 -626
rect -2465 -616 -1289 -560
rect -2465 -629 -2409 -616
rect -2564 -678 -2409 -629
rect -2631 -685 -2409 -678
rect -2631 -696 -2544 -685
rect -2145 -704 -2089 -616
rect -1985 -704 -1929 -616
rect -1825 -704 -1769 -616
rect -1665 -704 -1609 -616
rect -1195 -619 -885 -563
rect -1428 -676 -1346 -667
rect -1195 -676 -1139 -619
rect -1428 -680 -1139 -676
rect -1428 -731 -1415 -680
rect -1362 -731 -1139 -680
rect -1428 -732 -1139 -731
rect -1428 -745 -1346 -732
rect -1302 -1051 -1197 -1037
rect -1302 -1058 -1093 -1051
rect -1302 -1106 -1281 -1058
rect -1223 -1106 -1093 -1058
rect -1302 -1107 -1093 -1106
rect -1302 -1137 -1197 -1107
rect -1149 -1182 -1093 -1107
rect -941 -1182 -886 -1142
rect -1149 -1183 -885 -1182
rect -1149 -1238 5355 -1183
<< polycontact >>
rect -2616 -678 -2564 -626
rect -1415 -731 -1362 -680
rect -1281 -1106 -1223 -1058
<< metal1 >>
rect -1311 233 5529 271
rect -1311 175 -1205 233
rect -1142 175 -1005 233
rect -942 175 -805 233
rect -742 175 -605 233
rect -542 175 -405 233
rect -342 175 -205 233
rect -142 175 -5 233
rect 58 175 220 233
rect 283 175 420 233
rect 483 175 620 233
rect 683 175 820 233
rect 883 175 1020 233
rect 1083 175 1220 233
rect 1283 175 1420 233
rect 1483 175 1645 233
rect 1708 175 1845 233
rect 1908 175 2045 233
rect 2108 175 2245 233
rect 2308 175 2445 233
rect 2508 175 2645 233
rect 2708 175 2845 233
rect 2908 175 3070 233
rect 3133 175 3270 233
rect 3333 175 3470 233
rect 3533 175 3670 233
rect 3733 175 3870 233
rect 3933 175 4070 233
rect 4133 175 4270 233
rect 4333 175 4495 233
rect 4558 175 4695 233
rect 4758 175 4895 233
rect 4958 175 5095 233
rect 5158 175 5295 233
rect 5358 175 5529 233
rect -1311 130 5529 175
rect -1311 60 -1214 130
rect 5458 117 5529 130
rect -2639 22 -1214 60
rect -2639 -36 -2574 22
rect -2511 -36 -2374 22
rect -2311 -36 -2174 22
rect -2111 -36 -1974 22
rect -1911 -36 -1774 22
rect -1711 -36 -1574 22
rect -1511 -36 -1374 22
rect -1311 -36 -1214 22
rect -2639 -81 -1214 -36
rect -2540 -149 -2494 -81
rect -2220 -127 -2174 -81
rect -1900 -127 -1854 -81
rect -1580 -127 -1534 -81
rect -1260 -131 -1214 -81
rect -1075 -79 5430 60
rect -2380 -580 -2334 -522
rect -2060 -580 -2014 -522
rect -1740 -580 -1694 -523
rect -1420 -580 -1374 -523
rect -2631 -626 -2544 -613
rect -2380 -626 -1374 -580
rect -2631 -678 -2616 -626
rect -2564 -649 -2544 -626
rect -2564 -678 -2420 -649
rect -2631 -695 -2420 -678
rect -2631 -696 -2544 -695
rect -2664 -804 -2518 -774
rect -2664 -885 -2638 -804
rect -2542 -885 -2518 -804
rect -2664 -911 -2518 -885
rect -2466 -1059 -2420 -695
rect -2060 -750 -2014 -626
rect -1740 -755 -1694 -626
rect -1428 -667 -1374 -626
rect -1428 -680 -1346 -667
rect -1428 -731 -1415 -680
rect -1362 -731 -1346 -680
rect -1428 -745 -1346 -731
rect -1075 -779 -970 -79
rect -856 -750 -810 -489
rect -696 -750 -650 -79
rect -1246 -798 -970 -779
rect -1246 -874 -1224 -798
rect -1130 -874 -970 -798
rect -1246 -911 -970 -874
rect -1246 -917 -1103 -911
rect -1302 -1058 -1197 -1037
rect -2486 -1071 -2404 -1059
rect -2486 -1125 -2470 -1071
rect -2416 -1125 -2404 -1071
rect -2486 -1137 -2404 -1125
rect -1302 -1070 -1281 -1058
rect -1302 -1126 -1285 -1070
rect -1223 -1106 -1197 -1058
rect -1229 -1126 -1197 -1106
rect -1302 -1137 -1197 -1126
rect -2220 -1212 -2174 -1143
rect -1900 -1212 -1854 -1145
rect -1580 -1212 -1534 -1146
rect -856 -1205 -810 -1146
rect -536 -1205 -490 -489
rect -376 -750 -330 -79
rect -216 -1205 -170 -489
rect -56 -750 -10 -79
rect 104 -1205 150 -478
rect 264 -750 310 -79
rect 424 -1205 470 -478
rect 584 -750 630 -79
rect 744 -1205 790 -478
rect 904 -750 950 -79
rect 1064 -1205 1110 -478
rect 1224 -750 1270 -79
rect 1384 -1205 1430 -478
rect 1544 -750 1590 -79
rect 1704 -1205 1750 -478
rect 1864 -750 1910 -79
rect 2024 -1205 2070 -478
rect 2184 -750 2230 -79
rect 2344 -1205 2390 -478
rect 2504 -750 2550 -79
rect 2664 -1205 2710 -478
rect 2824 -750 2870 -79
rect 2984 -1205 3030 -478
rect 3144 -750 3190 -79
rect 3304 -1205 3350 -478
rect 3464 -750 3510 -79
rect 3624 -1205 3670 -478
rect 3784 -750 3830 -79
rect 3944 -1205 3990 -478
rect 4104 -750 4150 -79
rect 4264 -1205 4310 -478
rect 4424 -750 4470 -79
rect 4584 -1205 4630 -478
rect 4744 -750 4790 -79
rect 4904 -1205 4950 -478
rect 5064 -750 5110 -79
rect 5384 -127 5430 -79
rect 5224 -1205 5270 -478
rect 5384 -750 5430 -478
rect -2612 -1240 -1187 -1212
rect -2612 -1324 -2531 -1240
rect -2450 -1324 -2331 -1240
rect -2250 -1324 -2131 -1240
rect -2050 -1324 -1931 -1240
rect -1850 -1324 -1731 -1240
rect -1650 -1324 -1531 -1240
rect -1450 -1324 -1331 -1240
rect -1250 -1324 -1187 -1240
rect -2612 -1339 -1187 -1324
rect -856 -1332 5711 -1205
rect -1333 -1378 -1187 -1339
rect -1333 -1400 5702 -1378
rect -1333 -1484 -1157 -1400
rect -1076 -1484 -957 -1400
rect -876 -1484 -757 -1400
rect -676 -1484 -557 -1400
rect -476 -1484 -357 -1400
rect -276 -1484 -157 -1400
rect -76 -1484 43 -1400
rect 124 -1484 268 -1400
rect 349 -1484 468 -1400
rect 549 -1484 668 -1400
rect 749 -1484 868 -1400
rect 949 -1484 1068 -1400
rect 1149 -1484 1268 -1400
rect 1349 -1484 1468 -1400
rect 1549 -1484 1693 -1400
rect 1774 -1484 1893 -1400
rect 1974 -1484 2093 -1400
rect 2174 -1484 2293 -1400
rect 2374 -1484 2493 -1400
rect 2574 -1484 2693 -1400
rect 2774 -1484 2893 -1400
rect 2974 -1484 3118 -1400
rect 3199 -1484 3318 -1400
rect 3399 -1484 3518 -1400
rect 3599 -1484 3718 -1400
rect 3799 -1484 3918 -1400
rect 3999 -1484 4118 -1400
rect 4199 -1484 4318 -1400
rect 4399 -1484 4543 -1400
rect 4624 -1484 4743 -1400
rect 4824 -1484 4943 -1400
rect 5024 -1484 5143 -1400
rect 5224 -1484 5343 -1400
rect 5424 -1484 5543 -1400
rect 5624 -1484 5702 -1400
rect -1333 -1499 5702 -1484
<< via1 >>
rect -2638 -885 -2542 -804
rect -1224 -874 -1130 -798
rect -2470 -1125 -2416 -1071
rect -1285 -1106 -1281 -1070
rect -1281 -1106 -1229 -1070
rect -1285 -1126 -1229 -1106
<< metal2 >>
rect -2664 -798 -1103 -774
rect -2664 -804 -1224 -798
rect -2664 -885 -2638 -804
rect -2542 -874 -1224 -804
rect -1130 -847 -1103 -798
rect -1130 -874 -1101 -847
rect -2542 -885 -1101 -874
rect -2664 -911 -1101 -885
rect -1246 -917 -1103 -911
rect -2486 -1070 -2404 -1059
rect -1302 -1070 -1197 -1037
rect -2486 -1071 -1285 -1070
rect -2486 -1125 -2470 -1071
rect -2416 -1125 -1285 -1071
rect -2486 -1126 -1285 -1125
rect -1229 -1126 -1197 -1070
rect -2486 -1137 -2404 -1126
rect -1302 -1137 -1197 -1126
use nmos_3p3_AEBEG7  nmos_3p3_AEBEG7_0
timestamp 1692680230
transform 1 0 2207 0 1 -948
box -3260 -268 3260 268
use nmos_3p3_ECASTA  nmos_3p3_ECASTA_0
timestamp 1692680230
transform 1 0 -1877 0 1 -948
box -380 -268 380 268
use pmos_3p3_MLZUAR  pmos_3p3_MLZUAR_0
timestamp 1692680230
transform 1 0 -1877 0 1 -325
box -762 -330 762 330
use pmos_3p3_Q3Y3KU  pmos_3p3_Q3Y3KU_0
timestamp 1692680230
transform 1 0 2207 0 1 -325
box -3322 -330 3322 330
<< labels >>
flabel metal1 -2050 -19 -2050 -19 0 FreeSans 480 0 0 0 VDD
port 0 nsew
flabel metal1 -1995 -1290 -1995 -1290 0 FreeSans 480 0 0 0 VSS
port 1 nsew
flabel polycontact -2595 -658 -2595 -658 0 FreeSans 480 0 0 0 SEL
port 2 nsew
flabel metal1 5624 -1262 5624 -1262 0 FreeSans 480 0 0 0 OUT
port 4 nsew
flabel via1 -2601 -841 -2601 -841 0 FreeSans 480 0 0 0 IN
port 3 nsew
<< end >>
