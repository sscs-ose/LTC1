* NGSPICE file created from NAND_flat.ext - technology: gf180mcuC

.subckt pex_NAND VDD VSS A B OUT
X0 OUT A.t0 a_230_68# VSS.t2 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X1 VDD A.t1 OUT.t0 VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X2 a_230_68# B.t0 VSS.t1 VSS.t0 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X3 OUT B.t1 VDD.t4 VDD.t3 pfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 A.n0 A.t1 26.4688
R1 A.n0 A.t0 15.0091
R2 A A.n0 4.94817
R3 OUT.n1 OUT.n0 6.94485
R4 OUT.n3 OUT.n2 6.89411
R5 OUT.n1 OUT.t0 6.2405
R6 OUT.n3 OUT.n1 0.466152
R7 OUT OUT.n3 0.158978
R8 VSS.n1 VSS.t2 1692.54
R9 VSS.n1 VSS.t0 1517.73
R10 VSS VSS.t1 6.99468
R11 VSS.n2 VSS.n1 2.6005
R12 VSS VSS.n2 2.6005
R13 VSS.n2 VSS.n0 0.0188246
R14 VDD.n2 VDD.t3 445.175
R15 VDD.n2 VDD.t0 440.789
R16 VDD.n4 VDD.t4 6.82193
R17 VDD VDD.n0 6.81846
R18 VDD.n4 VDD.n3 3.1505
R19 VDD.n3 VDD.n2 3.1505
R20 VDD.n3 VDD.n1 0.158
R21 VDD VDD.n4 0.00223077
R22 B.n0 B.t0 25.5505
R23 B.n2 B.n0 19.4523
R24 B.n0 B.t1 14.4701
R25 B B.n2 4.00297
R26 B.n2 B.n1 0.2005
C0 A a_230_68# 0.235f
C1 A VDD 0.181f
C2 OUT A 0.212f
C3 B a_230_68# 8.64e-19
C4 B VDD 0.208f
C5 OUT B 0.014f
C6 OUT a_230_68# 0.038f
C7 OUT VDD 0.493f
C8 B A 0.121f
.ends

