magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 4032 71968
<< metal5 >>
rect 0 68400 2000 69678
rect 0 66800 2000 68200
rect 0 65200 2000 66600
rect 0 63600 2000 65000
rect 0 62000 2000 63400
rect 0 60400 2000 61800
rect 0 58800 2000 60200
rect 0 57200 2000 58600
rect 0 55600 2000 57000
rect 0 54000 2000 55400
rect 0 52400 2000 53800
rect 0 50800 2000 52200
rect 0 49200 2000 50600
rect 0 46000 2000 49000
rect 0 42800 2000 45800
rect 0 41200 2000 42600
rect 0 39600 2000 41000
rect 0 36400 2000 39400
rect 0 33200 2000 36200
rect 0 30000 2000 33000
rect 0 26800 2000 29800
rect 0 25200 2000 26600
rect 0 23600 2000 25000
rect 0 20400 2000 23400
rect 0 17200 2000 20200
rect 0 14000 2000 17000
use GF_NI_FILL10_0  GF_NI_FILL10_0_0
timestamp 1713338890
transform 1 0 0 0 1 0
box -32 13097 2032 69968
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_0
timestamp 1713338890
transform 1 0 1010 0 1 24302
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_1
timestamp 1713338890
transform 1 0 1010 0 1 25915
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_2
timestamp 1713338890
transform 1 0 1010 0 1 40305
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_3
timestamp 1713338890
transform 1 0 1010 0 1 41901
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_4
timestamp 1713338890
transform 1 0 1010 0 1 49894
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_5
timestamp 1713338890
transform 1 0 1010 0 1 51514
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_6
timestamp 1713338890
transform 1 0 1010 0 1 54694
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_7
timestamp 1713338890
transform 1 0 1010 0 1 53121
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_8
timestamp 1713338890
transform 1 0 1010 0 1 57899
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_9
timestamp 1713338890
transform 1 0 1010 0 1 56303
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_10
timestamp 1713338890
transform 1 0 1010 0 1 59504
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_11
timestamp 1713338890
transform 1 0 1010 0 1 62709
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_12
timestamp 1713338890
transform 1 0 1010 0 1 61109
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_13
timestamp 1713338890
transform 1 0 1010 0 1 65898
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_14
timestamp 1713338890
transform 1 0 1010 0 1 64300
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_15
timestamp 1713338890
transform 1 0 1010 0 1 67508
box -912 -602 912 602
use M5_M4_CDNS_6903358316562  M5_M4_CDNS_6903358316562_16
timestamp 1713338890
transform 1 0 1010 0 1 69038
box -912 -602 912 602
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_0
timestamp 1713338890
transform 1 0 1010 0 1 15522
box -912 -1346 912 1346
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_1
timestamp 1713338890
transform 1 0 1010 0 1 18693
box -912 -1346 912 1346
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_2
timestamp 1713338890
transform 1 0 1010 0 1 21904
box -912 -1346 912 1346
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_3
timestamp 1713338890
transform 1 0 1010 0 1 28313
box -912 -1346 912 1346
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_4
timestamp 1713338890
transform 1 0 1010 0 1 31514
box -912 -1346 912 1346
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_5
timestamp 1713338890
transform 1 0 1010 0 1 34729
box -912 -1346 912 1346
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_6
timestamp 1713338890
transform 1 0 1010 0 1 37914
box -912 -1346 912 1346
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_7
timestamp 1713338890
transform 1 0 1010 0 1 44322
box -912 -1346 912 1346
use M5_M4_CDNS_6903358316563  M5_M4_CDNS_6903358316563_8
timestamp 1713338890
transform 1 0 1010 0 1 47511
box -912 -1346 912 1346
<< labels >>
rlabel metal5 s 1018 18921 1018 18921 4 DVSS
port 1 nsew
rlabel metal5 s 1018 15750 1018 15750 4 DVSS
port 1 nsew
rlabel metal5 s 1018 21907 1018 21907 4 DVSS
port 1 nsew
rlabel metal5 s 1018 26100 1018 26100 4 DVSS
port 1 nsew
rlabel metal5 s 1018 40342 1018 40342 4 DVSS
port 1 nsew
rlabel metal5 s 1018 47595 1018 47595 4 DVSS
port 1 nsew
rlabel metal5 s 1018 57858 1018 57858 4 DVSS
port 1 nsew
rlabel metal5 s 1018 61058 1018 61058 4 DVSS
port 1 nsew
rlabel metal5 s 1018 66023 1018 66023 4 DVSS
port 1 nsew
rlabel metal5 s 1018 69049 1018 69049 4 DVSS
port 1 nsew
rlabel metal4 s 1018 69049 1018 69049 4 DVSS
port 1 nsew
rlabel metal4 s 1018 66023 1018 66023 4 DVSS
port 1 nsew
rlabel metal4 s 1018 61058 1018 61058 4 DVSS
port 1 nsew
rlabel metal4 s 1018 57858 1018 57858 4 DVSS
port 1 nsew
rlabel metal4 s 1018 47595 1018 47595 4 DVSS
port 1 nsew
rlabel metal4 s 1018 40342 1018 40342 4 DVSS
port 1 nsew
rlabel metal4 s 1018 26100 1018 26100 4 DVSS
port 1 nsew
rlabel metal4 s 1018 21907 1018 21907 4 DVSS
port 1 nsew
rlabel metal4 s 1018 15750 1018 15750 4 DVSS
port 1 nsew
rlabel metal4 s 1018 18921 1018 18921 4 DVSS
port 1 nsew
rlabel metal3 s 1018 66023 1018 66023 4 DVSS
port 1 nsew
rlabel metal3 s 1018 47595 1018 47595 4 DVSS
port 1 nsew
rlabel metal3 s 1018 57858 1018 57858 4 DVSS
port 1 nsew
rlabel metal3 s 1018 61058 1018 61058 4 DVSS
port 1 nsew
rlabel metal3 s 1018 15750 1018 15750 4 DVSS
port 1 nsew
rlabel metal3 s 1018 18921 1018 18921 4 DVSS
port 1 nsew
rlabel metal3 s 1018 21907 1018 21907 4 DVSS
port 1 nsew
rlabel metal3 s 1018 26100 1018 26100 4 DVSS
port 1 nsew
rlabel metal3 s 1018 40342 1018 40342 4 DVSS
port 1 nsew
rlabel metal3 s 1018 69049 1018 69049 4 DVSS
port 1 nsew
rlabel metal5 s 1018 31609 1018 31609 4 DVDD
port 2 nsew
rlabel metal5 s 1018 28394 1018 28394 4 DVDD
port 2 nsew
rlabel metal5 s 1018 24284 1018 24284 4 DVDD
port 2 nsew
rlabel metal5 s 1018 59623 1018 59623 4 DVDD
port 2 nsew
rlabel metal5 s 1018 56423 1018 56423 4 DVDD
port 2 nsew
rlabel metal5 s 1018 54658 1018 54658 4 DVDD
port 2 nsew
rlabel metal5 s 1018 53223 1018 53223 4 DVDD
port 2 nsew
rlabel metal5 s 1018 44368 1018 44368 4 DVDD
port 2 nsew
rlabel metal5 s 1018 41977 1018 41977 4 DVDD
port 2 nsew
rlabel metal5 s 1018 37959 1018 37959 4 DVDD
port 2 nsew
rlabel metal5 s 1018 34723 1018 34723 4 DVDD
port 2 nsew
rlabel metal5 s 1018 67458 1018 67458 4 DVDD
port 2 nsew
rlabel metal4 s 1018 67458 1018 67458 4 DVDD
port 2 nsew
rlabel metal4 s 1018 34723 1018 34723 4 DVDD
port 2 nsew
rlabel metal4 s 1018 37959 1018 37959 4 DVDD
port 2 nsew
rlabel metal4 s 1018 41977 1018 41977 4 DVDD
port 2 nsew
rlabel metal4 s 1018 44368 1018 44368 4 DVDD
port 2 nsew
rlabel metal4 s 1018 53223 1018 53223 4 DVDD
port 2 nsew
rlabel metal4 s 1018 54658 1018 54658 4 DVDD
port 2 nsew
rlabel metal4 s 1018 56423 1018 56423 4 DVDD
port 2 nsew
rlabel metal4 s 1018 59623 1018 59623 4 DVDD
port 2 nsew
rlabel metal4 s 1018 24284 1018 24284 4 DVDD
port 2 nsew
rlabel metal4 s 1018 28394 1018 28394 4 DVDD
port 2 nsew
rlabel metal4 s 1018 31609 1018 31609 4 DVDD
port 2 nsew
rlabel metal3 s 1018 67458 1018 67458 4 DVDD
port 2 nsew
rlabel metal3 s 1018 44368 1018 44368 4 DVDD
port 2 nsew
rlabel metal3 s 1018 53223 1018 53223 4 DVDD
port 2 nsew
rlabel metal3 s 1018 54658 1018 54658 4 DVDD
port 2 nsew
rlabel metal3 s 1018 56423 1018 56423 4 DVDD
port 2 nsew
rlabel metal3 s 1018 59623 1018 59623 4 DVDD
port 2 nsew
rlabel metal3 s 1018 24284 1018 24284 4 DVDD
port 2 nsew
rlabel metal3 s 1018 28394 1018 28394 4 DVDD
port 2 nsew
rlabel metal3 s 1018 31609 1018 31609 4 DVDD
port 2 nsew
rlabel metal3 s 1018 34723 1018 34723 4 DVDD
port 2 nsew
rlabel metal3 s 1018 37959 1018 37959 4 DVDD
port 2 nsew
rlabel metal3 s 1018 41977 1018 41977 4 DVDD
port 2 nsew
rlabel metal5 s 1018 51458 1018 51458 4 VDD
port 3 nsew
rlabel metal5 s 1018 62823 1018 62823 4 VDD
port 3 nsew
rlabel metal4 s 1018 62823 1018 62823 4 VDD
port 3 nsew
rlabel metal4 s 1018 51458 1018 51458 4 VDD
port 3 nsew
rlabel metal3 s 1018 62823 1018 62823 4 VDD
port 3 nsew
rlabel metal3 s 1018 51458 1018 51458 4 VDD
port 3 nsew
rlabel metal5 s 1018 64258 1018 64258 4 VSS
port 4 nsew
rlabel metal5 s 1018 50023 1018 50023 4 VSS
port 4 nsew
rlabel metal4 s 1018 50023 1018 50023 4 VSS
port 4 nsew
rlabel metal4 s 1018 64258 1018 64258 4 VSS
port 4 nsew
rlabel metal3 s 1018 64258 1018 64258 4 VSS
port 4 nsew
rlabel metal3 s 1018 50023 1018 50023 4 VSS
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2000 70000
<< end >>
