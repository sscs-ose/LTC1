magic
tech gf180mcuC
magscale 1 10
timestamp 1692680230
<< nwell >>
rect -3322 -330 3322 330
<< pmos >>
rect -3148 -200 -3092 200
rect -2988 -200 -2932 200
rect -2828 -200 -2772 200
rect -2668 -200 -2612 200
rect -2508 -200 -2452 200
rect -2348 -200 -2292 200
rect -2188 -200 -2132 200
rect -2028 -200 -1972 200
rect -1868 -200 -1812 200
rect -1708 -200 -1652 200
rect -1548 -200 -1492 200
rect -1388 -200 -1332 200
rect -1228 -200 -1172 200
rect -1068 -200 -1012 200
rect -908 -200 -852 200
rect -748 -200 -692 200
rect -588 -200 -532 200
rect -428 -200 -372 200
rect -268 -200 -212 200
rect -108 -200 -52 200
rect 52 -200 108 200
rect 212 -200 268 200
rect 372 -200 428 200
rect 532 -200 588 200
rect 692 -200 748 200
rect 852 -200 908 200
rect 1012 -200 1068 200
rect 1172 -200 1228 200
rect 1332 -200 1388 200
rect 1492 -200 1548 200
rect 1652 -200 1708 200
rect 1812 -200 1868 200
rect 1972 -200 2028 200
rect 2132 -200 2188 200
rect 2292 -200 2348 200
rect 2452 -200 2508 200
rect 2612 -200 2668 200
rect 2772 -200 2828 200
rect 2932 -200 2988 200
rect 3092 -200 3148 200
<< pdiff >>
rect -3236 187 -3148 200
rect -3236 -187 -3223 187
rect -3177 -187 -3148 187
rect -3236 -200 -3148 -187
rect -3092 187 -2988 200
rect -3092 -187 -3063 187
rect -3017 -187 -2988 187
rect -3092 -200 -2988 -187
rect -2932 187 -2828 200
rect -2932 -187 -2903 187
rect -2857 -187 -2828 187
rect -2932 -200 -2828 -187
rect -2772 187 -2668 200
rect -2772 -187 -2743 187
rect -2697 -187 -2668 187
rect -2772 -200 -2668 -187
rect -2612 187 -2508 200
rect -2612 -187 -2583 187
rect -2537 -187 -2508 187
rect -2612 -200 -2508 -187
rect -2452 187 -2348 200
rect -2452 -187 -2423 187
rect -2377 -187 -2348 187
rect -2452 -200 -2348 -187
rect -2292 187 -2188 200
rect -2292 -187 -2263 187
rect -2217 -187 -2188 187
rect -2292 -200 -2188 -187
rect -2132 187 -2028 200
rect -2132 -187 -2103 187
rect -2057 -187 -2028 187
rect -2132 -200 -2028 -187
rect -1972 187 -1868 200
rect -1972 -187 -1943 187
rect -1897 -187 -1868 187
rect -1972 -200 -1868 -187
rect -1812 187 -1708 200
rect -1812 -187 -1783 187
rect -1737 -187 -1708 187
rect -1812 -200 -1708 -187
rect -1652 187 -1548 200
rect -1652 -187 -1623 187
rect -1577 -187 -1548 187
rect -1652 -200 -1548 -187
rect -1492 187 -1388 200
rect -1492 -187 -1463 187
rect -1417 -187 -1388 187
rect -1492 -200 -1388 -187
rect -1332 187 -1228 200
rect -1332 -187 -1303 187
rect -1257 -187 -1228 187
rect -1332 -200 -1228 -187
rect -1172 187 -1068 200
rect -1172 -187 -1143 187
rect -1097 -187 -1068 187
rect -1172 -200 -1068 -187
rect -1012 187 -908 200
rect -1012 -187 -983 187
rect -937 -187 -908 187
rect -1012 -200 -908 -187
rect -852 187 -748 200
rect -852 -187 -823 187
rect -777 -187 -748 187
rect -852 -200 -748 -187
rect -692 187 -588 200
rect -692 -187 -663 187
rect -617 -187 -588 187
rect -692 -200 -588 -187
rect -532 187 -428 200
rect -532 -187 -503 187
rect -457 -187 -428 187
rect -532 -200 -428 -187
rect -372 187 -268 200
rect -372 -187 -343 187
rect -297 -187 -268 187
rect -372 -200 -268 -187
rect -212 187 -108 200
rect -212 -187 -183 187
rect -137 -187 -108 187
rect -212 -200 -108 -187
rect -52 187 52 200
rect -52 -187 -23 187
rect 23 -187 52 187
rect -52 -200 52 -187
rect 108 187 212 200
rect 108 -187 137 187
rect 183 -187 212 187
rect 108 -200 212 -187
rect 268 187 372 200
rect 268 -187 297 187
rect 343 -187 372 187
rect 268 -200 372 -187
rect 428 187 532 200
rect 428 -187 457 187
rect 503 -187 532 187
rect 428 -200 532 -187
rect 588 187 692 200
rect 588 -187 617 187
rect 663 -187 692 187
rect 588 -200 692 -187
rect 748 187 852 200
rect 748 -187 777 187
rect 823 -187 852 187
rect 748 -200 852 -187
rect 908 187 1012 200
rect 908 -187 937 187
rect 983 -187 1012 187
rect 908 -200 1012 -187
rect 1068 187 1172 200
rect 1068 -187 1097 187
rect 1143 -187 1172 187
rect 1068 -200 1172 -187
rect 1228 187 1332 200
rect 1228 -187 1257 187
rect 1303 -187 1332 187
rect 1228 -200 1332 -187
rect 1388 187 1492 200
rect 1388 -187 1417 187
rect 1463 -187 1492 187
rect 1388 -200 1492 -187
rect 1548 187 1652 200
rect 1548 -187 1577 187
rect 1623 -187 1652 187
rect 1548 -200 1652 -187
rect 1708 187 1812 200
rect 1708 -187 1737 187
rect 1783 -187 1812 187
rect 1708 -200 1812 -187
rect 1868 187 1972 200
rect 1868 -187 1897 187
rect 1943 -187 1972 187
rect 1868 -200 1972 -187
rect 2028 187 2132 200
rect 2028 -187 2057 187
rect 2103 -187 2132 187
rect 2028 -200 2132 -187
rect 2188 187 2292 200
rect 2188 -187 2217 187
rect 2263 -187 2292 187
rect 2188 -200 2292 -187
rect 2348 187 2452 200
rect 2348 -187 2377 187
rect 2423 -187 2452 187
rect 2348 -200 2452 -187
rect 2508 187 2612 200
rect 2508 -187 2537 187
rect 2583 -187 2612 187
rect 2508 -200 2612 -187
rect 2668 187 2772 200
rect 2668 -187 2697 187
rect 2743 -187 2772 187
rect 2668 -200 2772 -187
rect 2828 187 2932 200
rect 2828 -187 2857 187
rect 2903 -187 2932 187
rect 2828 -200 2932 -187
rect 2988 187 3092 200
rect 2988 -187 3017 187
rect 3063 -187 3092 187
rect 2988 -200 3092 -187
rect 3148 187 3236 200
rect 3148 -187 3177 187
rect 3223 -187 3236 187
rect 3148 -200 3236 -187
<< pdiffc >>
rect -3223 -187 -3177 187
rect -3063 -187 -3017 187
rect -2903 -187 -2857 187
rect -2743 -187 -2697 187
rect -2583 -187 -2537 187
rect -2423 -187 -2377 187
rect -2263 -187 -2217 187
rect -2103 -187 -2057 187
rect -1943 -187 -1897 187
rect -1783 -187 -1737 187
rect -1623 -187 -1577 187
rect -1463 -187 -1417 187
rect -1303 -187 -1257 187
rect -1143 -187 -1097 187
rect -983 -187 -937 187
rect -823 -187 -777 187
rect -663 -187 -617 187
rect -503 -187 -457 187
rect -343 -187 -297 187
rect -183 -187 -137 187
rect -23 -187 23 187
rect 137 -187 183 187
rect 297 -187 343 187
rect 457 -187 503 187
rect 617 -187 663 187
rect 777 -187 823 187
rect 937 -187 983 187
rect 1097 -187 1143 187
rect 1257 -187 1303 187
rect 1417 -187 1463 187
rect 1577 -187 1623 187
rect 1737 -187 1783 187
rect 1897 -187 1943 187
rect 2057 -187 2103 187
rect 2217 -187 2263 187
rect 2377 -187 2423 187
rect 2537 -187 2583 187
rect 2697 -187 2743 187
rect 2857 -187 2903 187
rect 3017 -187 3063 187
rect 3177 -187 3223 187
<< polysilicon >>
rect -3148 200 -3092 244
rect -2988 200 -2932 244
rect -2828 200 -2772 244
rect -2668 200 -2612 244
rect -2508 200 -2452 244
rect -2348 200 -2292 244
rect -2188 200 -2132 244
rect -2028 200 -1972 244
rect -1868 200 -1812 244
rect -1708 200 -1652 244
rect -1548 200 -1492 244
rect -1388 200 -1332 244
rect -1228 200 -1172 244
rect -1068 200 -1012 244
rect -908 200 -852 244
rect -748 200 -692 244
rect -588 200 -532 244
rect -428 200 -372 244
rect -268 200 -212 244
rect -108 200 -52 244
rect 52 200 108 244
rect 212 200 268 244
rect 372 200 428 244
rect 532 200 588 244
rect 692 200 748 244
rect 852 200 908 244
rect 1012 200 1068 244
rect 1172 200 1228 244
rect 1332 200 1388 244
rect 1492 200 1548 244
rect 1652 200 1708 244
rect 1812 200 1868 244
rect 1972 200 2028 244
rect 2132 200 2188 244
rect 2292 200 2348 244
rect 2452 200 2508 244
rect 2612 200 2668 244
rect 2772 200 2828 244
rect 2932 200 2988 244
rect 3092 200 3148 244
rect -3148 -244 -3092 -200
rect -2988 -244 -2932 -200
rect -2828 -244 -2772 -200
rect -2668 -244 -2612 -200
rect -2508 -244 -2452 -200
rect -2348 -244 -2292 -200
rect -2188 -244 -2132 -200
rect -2028 -244 -1972 -200
rect -1868 -244 -1812 -200
rect -1708 -244 -1652 -200
rect -1548 -244 -1492 -200
rect -1388 -244 -1332 -200
rect -1228 -244 -1172 -200
rect -1068 -244 -1012 -200
rect -908 -244 -852 -200
rect -748 -244 -692 -200
rect -588 -244 -532 -200
rect -428 -244 -372 -200
rect -268 -244 -212 -200
rect -108 -244 -52 -200
rect 52 -244 108 -200
rect 212 -244 268 -200
rect 372 -244 428 -200
rect 532 -244 588 -200
rect 692 -244 748 -200
rect 852 -244 908 -200
rect 1012 -244 1068 -200
rect 1172 -244 1228 -200
rect 1332 -244 1388 -200
rect 1492 -244 1548 -200
rect 1652 -244 1708 -200
rect 1812 -244 1868 -200
rect 1972 -244 2028 -200
rect 2132 -244 2188 -200
rect 2292 -244 2348 -200
rect 2452 -244 2508 -200
rect 2612 -244 2668 -200
rect 2772 -244 2828 -200
rect 2932 -244 2988 -200
rect 3092 -244 3148 -200
<< metal1 >>
rect -3223 187 -3177 198
rect -3223 -198 -3177 -187
rect -3063 187 -3017 198
rect -3063 -198 -3017 -187
rect -2903 187 -2857 198
rect -2903 -198 -2857 -187
rect -2743 187 -2697 198
rect -2743 -198 -2697 -187
rect -2583 187 -2537 198
rect -2583 -198 -2537 -187
rect -2423 187 -2377 198
rect -2423 -198 -2377 -187
rect -2263 187 -2217 198
rect -2263 -198 -2217 -187
rect -2103 187 -2057 198
rect -2103 -198 -2057 -187
rect -1943 187 -1897 198
rect -1943 -198 -1897 -187
rect -1783 187 -1737 198
rect -1783 -198 -1737 -187
rect -1623 187 -1577 198
rect -1623 -198 -1577 -187
rect -1463 187 -1417 198
rect -1463 -198 -1417 -187
rect -1303 187 -1257 198
rect -1303 -198 -1257 -187
rect -1143 187 -1097 198
rect -1143 -198 -1097 -187
rect -983 187 -937 198
rect -983 -198 -937 -187
rect -823 187 -777 198
rect -823 -198 -777 -187
rect -663 187 -617 198
rect -663 -198 -617 -187
rect -503 187 -457 198
rect -503 -198 -457 -187
rect -343 187 -297 198
rect -343 -198 -297 -187
rect -183 187 -137 198
rect -183 -198 -137 -187
rect -23 187 23 198
rect -23 -198 23 -187
rect 137 187 183 198
rect 137 -198 183 -187
rect 297 187 343 198
rect 297 -198 343 -187
rect 457 187 503 198
rect 457 -198 503 -187
rect 617 187 663 198
rect 617 -198 663 -187
rect 777 187 823 198
rect 777 -198 823 -187
rect 937 187 983 198
rect 937 -198 983 -187
rect 1097 187 1143 198
rect 1097 -198 1143 -187
rect 1257 187 1303 198
rect 1257 -198 1303 -187
rect 1417 187 1463 198
rect 1417 -198 1463 -187
rect 1577 187 1623 198
rect 1577 -198 1623 -187
rect 1737 187 1783 198
rect 1737 -198 1783 -187
rect 1897 187 1943 198
rect 1897 -198 1943 -187
rect 2057 187 2103 198
rect 2057 -198 2103 -187
rect 2217 187 2263 198
rect 2217 -198 2263 -187
rect 2377 187 2423 198
rect 2377 -198 2423 -187
rect 2537 187 2583 198
rect 2537 -198 2583 -187
rect 2697 187 2743 198
rect 2697 -198 2743 -187
rect 2857 187 2903 198
rect 2857 -198 2903 -187
rect 3017 187 3063 198
rect 3017 -198 3063 -187
rect 3177 187 3223 198
rect 3177 -198 3223 -187
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2 l 0.280 m 1 nf 40 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
