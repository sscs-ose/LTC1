magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1669 1019 1669
<< metal1 >>
rect -19 663 19 669
rect -19 -663 -13 663
rect 13 -663 19 663
rect -19 -669 19 -663
<< via1 >>
rect -13 -663 13 663
<< metal2 >>
rect -19 663 19 669
rect -19 -663 -13 663
rect 13 -663 19 663
rect -19 -669 19 -663
<< end >>
