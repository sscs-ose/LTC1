magic
tech gf180mcuC
magscale 1 10
timestamp 1695206022
<< nwell >>
rect 10248 3042 10374 3094
rect 10247 3041 10374 3042
rect 11287 3041 11348 3094
rect 10247 2717 10321 3041
rect 11252 2681 11501 2708
rect 11252 2679 11504 2681
rect 11269 2671 11504 2679
rect 11252 2661 11487 2664
rect 11252 2652 11503 2661
rect 11251 2635 11502 2652
rect 11874 2639 11887 2644
rect 6789 2003 6846 2079
rect 9416 1947 9464 1949
rect 3150 1861 3207 1946
rect 9184 1863 9241 1895
rect 9461 1892 9465 1947
rect 9586 1944 9642 1945
rect 9384 1891 9472 1892
rect 9585 1887 9642 1889
rect 1475 608 1482 618
rect 1475 554 1485 608
rect 1529 558 1541 620
rect 4477 618 4552 626
rect 1537 554 1540 558
rect 1475 550 1540 554
rect 4477 555 4565 618
rect 4477 553 4552 555
rect 1482 523 1540 550
rect 10473 549 10523 625
<< pwell >>
rect 2796 1558 3167 1591
<< nsubdiff >>
rect 6789 2003 6846 2079
<< polysilicon >>
rect 9593 1594 9657 1605
<< metal1 >>
rect 11213 3407 11430 3419
rect 11213 3346 11479 3407
rect 11213 3300 11435 3346
rect 7141 3096 7491 3245
rect 7141 3090 7349 3096
rect 2963 1983 3024 2089
rect 5978 1983 6038 2089
rect 6789 2003 6846 2079
rect 7141 1999 7290 3090
rect 10191 3080 10457 3186
rect 10348 3071 10457 3080
rect 11213 3072 11304 3300
rect 11213 3071 11302 3072
rect 11219 3070 11302 3071
rect 10160 2663 10248 2709
rect 11252 2681 11501 2708
rect 11252 2673 11504 2681
rect 10101 2591 10424 2663
rect 11252 2653 11505 2673
rect 11252 2652 11503 2653
rect 11251 2635 11502 2652
rect 11978 2576 12021 2610
rect 8310 2380 8423 2486
rect 9279 2380 9392 2486
rect 10236 2467 10349 2486
rect 10185 2404 10350 2467
rect 10236 2380 10349 2404
rect 11298 2195 11359 2394
rect 11831 2197 12197 2302
rect 8767 2004 8897 2060
rect 8997 2036 9055 2089
rect 8996 1983 9104 2036
rect 9 1602 38 1639
rect 481 1569 507 1601
rect 9593 1597 9657 1605
rect 9593 1594 9597 1597
rect 2803 1544 2828 1585
rect 5824 1540 5846 1584
rect 8835 1548 8864 1584
rect 9652 1594 9657 1597
rect 11862 1543 11885 1589
rect 1539 551 1549 598
rect 1555 551 1569 591
rect 476 472 505 508
rect 9543 506 9600 716
rect 9543 467 9592 506
rect 11942 455 12012 481
rect 12092 109 12197 2197
rect 2856 0 3301 109
rect 5873 0 6332 109
rect 8890 0 9395 109
rect 11907 0 12197 109
<< via1 >>
rect 7729 2743 7781 2795
rect 7471 2648 7523 2700
rect 8248 2692 8300 2744
rect 8711 2743 8763 2795
rect 9665 2742 9717 2794
rect 8454 2637 8506 2689
rect 9216 2686 9268 2738
rect 9418 2637 9470 2689
rect 11671 2656 11723 2708
rect 11817 2640 11869 2692
rect 543 1539 595 1591
rect 3563 1540 3615 1592
rect 6575 1539 6627 1591
rect 9597 1545 9649 1597
rect 1485 553 1537 605
rect 4503 549 4555 601
rect 7519 550 7571 602
rect 10536 550 10588 602
rect 542 453 594 505
rect 3541 454 3593 506
rect 6575 453 6627 505
rect 9592 454 9644 506
<< metal2 >>
rect 8246 2863 11725 2919
rect 7727 2795 7783 2807
rect 7727 2743 7729 2795
rect 7781 2743 7783 2795
rect 7467 2700 7526 2712
rect 7467 2648 7471 2700
rect 7523 2648 7526 2700
rect 6789 2069 6846 2079
rect 6845 2060 6846 2069
rect 7467 2060 7526 2648
rect 7727 2173 7783 2743
rect 8246 2744 8302 2863
rect 8246 2692 8248 2744
rect 8300 2692 8302 2744
rect 8709 2795 8765 2807
rect 8709 2743 8711 2795
rect 8763 2743 8765 2795
rect 9660 2794 9721 2806
rect 8246 2680 8302 2692
rect 8452 2689 8508 2701
rect 8452 2637 8454 2689
rect 8506 2637 8508 2689
rect 8452 2173 8508 2637
rect 7727 2117 8587 2173
rect 8643 2117 8653 2173
rect 8709 2060 8765 2743
rect 9214 2738 9270 2750
rect 9214 2686 9216 2738
rect 9268 2686 9270 2738
rect 9660 2742 9665 2794
rect 9717 2742 9721 2794
rect 9214 2174 9270 2686
rect 9416 2689 9472 2701
rect 9416 2637 9418 2689
rect 9470 2637 9472 2689
rect 9416 2296 9472 2637
rect 9416 2230 9472 2240
rect 9214 2173 9604 2174
rect 9214 2117 9538 2173
rect 9594 2117 9604 2173
rect 9214 2116 9604 2117
rect 9660 2060 9721 2742
rect 11669 2708 11725 2863
rect 11669 2656 11671 2708
rect 11723 2656 11725 2708
rect 11669 2644 11725 2656
rect 11815 2692 11871 2704
rect 6845 2013 8765 2060
rect 6789 2004 8765 2013
rect 8821 2004 8831 2060
rect 8887 2004 9721 2060
rect 11815 2640 11817 2692
rect 11869 2640 11871 2692
rect 6789 2003 6846 2004
rect 3150 1891 9406 1947
rect 9462 1891 9472 1947
rect 3150 1890 9472 1891
rect 537 1591 597 1603
rect 3150 1591 3207 1890
rect 9184 1664 9241 1890
rect 537 1539 543 1591
rect 595 1539 597 1591
rect 2796 1564 3207 1591
rect 2787 1551 3207 1564
rect 537 505 597 1539
rect 2796 1535 3207 1551
rect 3561 1592 3617 1604
rect 3561 1540 3563 1592
rect 3615 1540 3617 1592
rect 6569 1591 6629 1603
rect 9583 1598 9658 1608
rect 9583 1597 9598 1598
rect 3561 741 3617 1540
rect 5810 1535 6236 1591
rect 6569 1539 6575 1591
rect 6627 1539 6629 1591
rect 3561 740 3717 741
rect 3561 684 3651 740
rect 3707 684 3717 740
rect 1465 616 1541 618
rect 1465 560 1475 616
rect 1531 605 1541 616
rect 1465 553 1485 560
rect 1537 558 1541 605
rect 4477 616 4557 626
rect 4477 560 4492 616
rect 4548 601 4557 616
rect 1537 553 1540 558
rect 1465 519 1540 553
rect 4477 549 4503 560
rect 4555 549 4557 601
rect 4477 519 4557 549
rect 537 453 542 505
rect 594 453 597 505
rect 537 447 597 453
rect 3529 506 3605 508
rect 3529 454 3541 506
rect 3593 454 3605 506
rect 3529 451 3605 454
rect 6569 505 6629 1539
rect 9583 1545 9597 1597
rect 9583 1542 9598 1545
rect 9654 1542 9658 1598
rect 11815 1588 11871 2640
rect 11838 1567 11871 1588
rect 11848 1566 11871 1567
rect 11850 1552 11871 1566
rect 9583 1503 9658 1542
rect 11851 1535 11871 1552
rect 7494 616 7574 626
rect 7494 560 7509 616
rect 7565 602 7574 616
rect 7494 550 7519 560
rect 7571 550 7574 602
rect 7494 519 7574 550
rect 10511 616 10590 626
rect 10511 560 10526 616
rect 10582 602 10590 616
rect 10511 550 10536 560
rect 10588 550 10590 602
rect 10511 519 10590 550
rect 6569 453 6575 505
rect 6627 453 6629 505
rect 537 441 596 447
rect 539 154 596 441
rect 3529 154 3585 451
rect 6569 154 6629 453
rect 9586 506 9646 518
rect 9586 454 9592 506
rect 9644 454 9646 506
rect 9586 154 9646 454
rect 539 98 9646 154
<< via2 >>
rect 6789 2013 6845 2069
rect 8587 2117 8643 2173
rect 9416 2240 9472 2296
rect 9538 2117 9594 2173
rect 8831 2004 8887 2060
rect 9406 1891 9462 1947
rect 6790 1654 6846 1710
rect 9598 1597 9654 1598
rect 3651 684 3707 740
rect 1475 605 1531 616
rect 1475 560 1485 605
rect 1485 560 1531 605
rect 4492 601 4548 616
rect 4492 560 4503 601
rect 4503 560 4548 601
rect 8768 1535 8824 1591
rect 9598 1545 9649 1597
rect 9649 1545 9654 1597
rect 9598 1542 9654 1545
rect 10105 684 10161 740
rect 7509 602 7565 616
rect 7509 560 7519 602
rect 7519 560 7565 602
rect 10526 602 10582 616
rect 10526 560 10536 602
rect 10536 560 10582 602
<< metal3 >>
rect 9416 2296 9472 2306
rect 8577 2117 8587 2173
rect 8643 2117 8824 2173
rect 6789 2069 6846 2079
rect 6845 2013 6846 2069
rect 6789 1710 6846 2013
rect 6789 1654 6790 1710
rect 6789 1643 6846 1654
rect 8768 2060 8824 2117
rect 8768 2004 8831 2060
rect 8887 2004 8897 2060
rect 8768 1591 8824 2004
rect 9416 1947 9472 2240
rect 9528 2173 9642 2174
rect 9528 2117 9538 2173
rect 9594 2117 9642 2173
rect 9528 2116 9642 2117
rect 9384 1891 9406 1947
rect 9462 1891 9472 1947
rect 8768 1525 8824 1535
rect 9583 1608 9642 2116
rect 9583 1598 9671 1608
rect 9583 1542 9598 1598
rect 9654 1542 9671 1598
rect 9583 1533 9671 1542
rect 3641 740 10070 741
rect 3641 684 3651 740
rect 3707 684 10105 740
rect 10161 684 10171 740
rect 1472 616 10599 626
rect 1472 560 1475 616
rect 1531 560 4492 616
rect 4548 560 7509 616
rect 7565 560 10526 616
rect 10582 560 10599 616
rect 1472 549 10599 560
use and2_mag  and2_mag_0
timestamp 1695127730
transform 1 0 7406 0 1 2382
box -70 -188 1009 863
use and2_mag  and2_mag_1
timestamp 1695127730
transform 1 0 9342 0 1 2382
box -70 -188 1009 863
use and2_mag  and2_mag_2
timestamp 1695127730
transform 1 0 8374 0 1 2382
box -70 -188 1009 863
use Buffer_delayed_mag  Buffer_delayed_mag_0
timestamp 1694693600
transform 1 0 10470 0 1 2463
box -218 -175 878 631
use JK_FF_mag  JK_FF_mag_0
timestamp 1695127730
transform 1 0 9441 0 1 0
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_1
timestamp 1695127730
transform 1 0 390 0 1 0
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_2
timestamp 1695127730
transform 1 0 3407 0 1 0
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_3
timestamp 1695127730
transform 1 0 6424 0 1 0
box -390 0 2603 2148
use nor_3_mag  nor_3_mag_0
timestamp 1695119997
transform 1 0 11018 0 1 1755
box 329 440 1054 1778
<< labels >>
flabel metal3 1544 593 1544 593 0 FreeSans 320 0 0 0 RST
port 0 nsew
flabel metal1 22 1615 22 1615 0 FreeSans 320 0 0 0 CLK
port 1 nsew
flabel metal1 3049 74 3049 74 0 FreeSans 320 0 0 0 VSS
port 2 nsew
flabel metal1 2984 2031 2984 2031 0 FreeSans 320 0 0 0 VDD
port 3 nsew
flabel metal2 2817 1562 2817 1562 0 FreeSans 320 0 0 0 Q0
port 4 nsew
flabel metal2 5836 1565 5836 1565 0 FreeSans 320 0 0 0 Q1
port 5 nsew
flabel metal1 8847 1567 8847 1567 0 FreeSans 320 0 0 0 Q2
port 6 nsew
flabel metal1 11875 1567 11875 1567 0 FreeSans 320 0 0 0 Q3
port 7 nsew
flabel metal1 11998 2594 11998 2594 0 FreeSans 320 0 0 0 Vdiv10
port 8 nsew
<< end >>
