* NGSPICE file created from PGA_Dec_Layout_flat.ext - technology: gf180mcuC

.subckt PGA_Decoder_PEX S2 S3 S1 VDD A S6 B S4 C VSS S5
X0 a_3328_375# C.t0 a_3184_375# VSS.t14 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X1 a_945_n363# B.t0 a_1425_n363# VSS.t28 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 VDD C.t1 a_801_n1645# VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_3808_375# B.t1 a_3328_375# VSS.t11 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X4 VDD C.t2 OR_2_In_Layout_0.B VDD.t31 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X5 VDD OR_2_In_Layout_0.B a_801_n363# VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 a_3184_n363# OR_2_In_Layout_0.A VDD.t65 VDD.t64 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 S3 a_3184_n363# VDD.t3 VDD.t2 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X8 VSS C.t3 a_1425_375# VSS.t17 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X9 S4 a_801_n1645# VSS.t84 VSS.t83 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X10 VDD A.t0 a_801_375# VDD.t44 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X11 S6 a_801_375# VDD.t21 VDD.t20 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X12 a_801_375# A.t1 a_945_375# VSS.t7 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X13 a_801_n363# B.t2 VDD.t57 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X14 a_1425_n1645# OR_2_In_Layout_0.A a_945_n1645# VSS.t80 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X15 AND_2_In_Layout_0.A a_3303_n1718# VSS.t41 VSS.t40 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X16 a_945_375# B.t3 a_1425_375# VSS.t28 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X17 VSS C.t4 a_1425_n1645# VSS.t56 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X18 S1 a_4292_n1650# VDD.t37 VDD.t36 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X19 S2 a_3184_375# VDD.t70 VDD.t69 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X20 a_3808_n363# OR_2_In_Layout_0.A a_3328_n363# VSS.t11 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X21 a_3808_n363# OR_2_In_Layout_0.A a_3328_n363# VSS.t79 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X22 VDD A.t2 AND_3_In_Layout_1.C VDD.t66 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X23 a_945_n1645# A.t3 a_801_n1645# VSS.t29 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X24 VSS C.t5 a_1425_n1645# VSS.t53 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X25 a_1425_375# B.t4 a_945_375# VSS.t39 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X26 a_1425_n363# B.t5 a_945_n363# VSS.t74 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X27 VSS B.t6 OR_2_In_Layout_0.A VSS.t34 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X28 a_945_n363# A.t4 a_801_n363# VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X29 VDD OR_2_In_Layout_0.B a_3184_n363# VDD.t14 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X30 VDD A.t5 a_3184_n363# VDD.t4 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X31 a_3303_n1718# OR_2_In_Layout_0.B a_2999_n1346# VDD.t13 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X32 S3 a_3184_n363# VSS.t3 VSS.t2 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X33 VDD a_3303_n1718# AND_2_In_Layout_0.A VDD.t22 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X34 VDD AND_3_In_Layout_1.C a_4292_n1650# VDD.t40 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X35 a_1425_n1645# OR_2_In_Layout_0.A a_945_n1645# VSS.t78 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X36 a_3808_375# B.t7 a_3328_375# VSS.t79 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X37 VSS AND_3_In_Layout_1.C a_3808_375# VSS.t8 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X38 VDD A.t6 a_801_n363# VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X39 VDD C.t6 a_3184_375# VDD.t28 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X40 S5 a_801_n363# VSS.t6 VSS.t5 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X41 VSS C.t7 OR_2_In_Layout_0.B VSS.t50 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X42 a_3184_375# C.t8 a_3328_375# VSS.t26 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X43 a_3328_375# B.t8 a_3808_375# VSS.t4 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X44 S6 a_801_375# VSS.t33 VSS.t5 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X45 a_4292_n1650# AND_2_In_Layout_0.A a_4148_n1650# VSS.t1 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X46 a_3328_n363# OR_2_In_Layout_0.B a_3184_n363# VSS.t27 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X47 a_4148_n1650# AND_3_In_Layout_1.C VSS.t71 VSS.t70 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X48 a_801_375# B.t9 VDD.t55 VDD.t54 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X49 a_945_375# A.t7 a_801_375# VSS.t12 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X50 a_2999_n1346# OR_2_In_Layout_0.A VDD.t63 VDD.t62 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X51 a_3184_n363# OR_2_In_Layout_0.B a_3328_n363# VSS.t26 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X52 a_801_n1645# OR_2_In_Layout_0.A VDD.t61 VDD.t56 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X53 a_4292_n1650# AND_2_In_Layout_0.A VDD.t1 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X54 a_945_375# A.t8 a_801_375# VSS.t13 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X55 a_3328_375# C.t9 a_3184_375# VSS.t27 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X56 VDD B.t10 OR_2_In_Layout_0.A VDD.t51 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X57 a_801_n363# A.t9 a_945_n363# VSS.t7 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X58 VSS A.t10 a_3808_n363# VSS.t8 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X59 VSS OR_2_In_Layout_0.B a_1425_n363# VSS.t23 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X60 a_945_n1645# A.t11 a_801_n1645# VSS.t38 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X61 VSS OR_2_In_Layout_0.B a_3303_n1718# VSS.t20 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X62 VDD C.t10 a_801_375# VDD.t25 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X63 a_1425_375# B.t11 a_945_375# VSS.t74 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X64 VSS OR_2_In_Layout_0.B a_1425_n363# VSS.t17 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X65 VSS AND_3_In_Layout_1.C a_4148_n1650# VSS.t67 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X66 S1 a_4292_n1650# VSS.t62 VSS.t61 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X67 VSS C.t11 a_1425_375# VSS.t23 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X68 a_1425_n363# OR_2_In_Layout_0.B VSS.t16 VSS.t15 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X69 VDD AND_3_In_Layout_1.C a_3184_375# VDD.t38 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X70 S5 a_801_n363# VDD.t8 VDD.t7 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X71 VDD OR_2_In_Layout_0.A a_2999_n1346# VDD.t58 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X72 VSS AND_3_In_Layout_1.C a_3808_375# VSS.t42 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X73 VDD A.t12 a_801_n1645# VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X74 a_2999_n1346# OR_2_In_Layout_0.B a_3303_n1718# VDD.t12 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X75 S2 a_3184_375# VSS.t81 VSS.t2 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X76 S4 a_801_n1645# VDD.t71 VDD.t7 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X77 a_1425_n1645# C.t12 VSS.t47 VSS.t46 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X78 a_3184_375# B.t12 VDD.t50 VDD.t49 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X79 a_3328_n363# OR_2_In_Layout_0.B a_3184_n363# VSS.t14 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X80 VSS A.t13 AND_3_In_Layout_1.C VSS.t30 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
X81 a_1425_375# C.t13 VSS.t45 VSS.t15 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X82 a_801_n1645# A.t14 a_945_n1645# VSS.t37 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X83 a_3303_n1718# OR_2_In_Layout_0.A VSS.t77 VSS.t76 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X84 a_3808_n363# A.t15 VSS.t82 VSS.t63 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X85 a_945_n1645# OR_2_In_Layout_0.A a_1425_n1645# VSS.t75 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X86 a_4148_n1650# AND_2_In_Layout_0.A a_4292_n1650# VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X87 a_3808_375# AND_3_In_Layout_1.C VSS.t64 VSS.t63 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X88 a_945_n363# A.t16 a_801_n363# VSS.t13 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X89 a_3328_n363# OR_2_In_Layout_0.A a_3808_n363# VSS.t4 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X90 VSS A.t17 a_3808_n363# VSS.t42 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X91 a_1425_n363# B.t13 a_945_n363# VSS.t39 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
R0 C.t11 C.t10 68.5684
R1 C.t4 C.t1 68.5684
R2 C.n1 C.t6 39.6291
R3 C C.n4 37.2709
R4 C C.n10 37.2709
R5 C.n6 C.t2 34.6755
R6 C.n0 C.t0 29.9826
R7 C.t9 C.n0 29.9826
R8 C.n3 C.t11 29.9826
R9 C.n9 C.t4 29.9826
R10 C.n1 C.t9 28.9398
R11 C C.n1 21.7803
R12 C.n4 C.n3 20.8576
R13 C.n10 C.n9 20.8576
R14 C.n7 C.n6 15.6818
R15 C.n6 C.t7 13.0362
R16 C.n0 C.t8 9.1255
R17 C.n4 C.t3 9.1255
R18 C.n3 C.t13 9.1255
R19 C.n10 C.t5 9.1255
R20 C.n9 C.t12 9.1255
R21 C.n8 C.n7 8.94075
R22 C.n2 C 7.52298
R23 C C.n8 3.42211
R24 C.n2 C 3.3252
R25 C.n5 C 2.46264
R26 C.n8 C.n5 2.2178
R27 C.n5 C.n2 0.687246
R28 C.n7 C 0.0956588
R29 VSS.n32 VSS.n31 3733.93
R30 VSS.n142 VSS.n141 2883.68
R31 VSS.n175 VSS.t30 921.495
R32 VSS.n175 VSS.t34 921.495
R33 VSS.n247 VSS.t20 277.728
R34 VSS.n88 VSS.n87 272.283
R35 VSS.n264 VSS.t0 241.91
R36 VSS.n210 VSS.t78 177.369
R37 VSS.n208 VSS.t75 166.935
R38 VSS.n165 VSS.t37 150.829
R39 VSS.n185 VSS.n184 140.055
R40 VSS.n94 VSS.t8 127.451
R41 VSS.n226 VSS.t53 125.329
R42 VSS.n195 VSS.t38 125.201
R43 VSS.n40 VSS.t7 121.659
R44 VSS.n161 VSS.t46 114.767
R45 VSS.n33 VSS.n32 112.969
R46 VSS.n251 VSS.t40 112.273
R47 VSS.n241 VSS.t76 112.273
R48 VSS.n267 VSS.t67 105.178
R49 VSS.n58 VSS.t39 98.4853
R50 VSS.n111 VSS.t79 98.4853
R51 VSS.n258 VSS.t1 94.6607
R52 VSS.n56 VSS.t28 92.6921
R53 VSS.n113 VSS.t4 92.6921
R54 VSS.n143 VSS.n142 80.9189
R55 VSS.n43 VSS.t12 69.5192
R56 VSS.n126 VSS.t27 69.5192
R57 VSS.n25 VSS.t15 63.726
R58 VSS.n97 VSS.t63 63.726
R59 VSS.n153 VSS.t17 58.3678
R60 VSS.n25 VSS.n24 57.9328
R61 VSS.n129 VSS.t26 55.7148
R62 VSS.n126 VSS.n125 52.1395
R63 VSS.n188 VSS.t29 50.2767
R64 VSS.n85 VSS.t2 46.3463
R65 VSS.n233 VSS.t83 45.5746
R66 VSS.n3 VSS.t61 42.0717
R67 VSS.n13 VSS.t70 42.0717
R68 VSS.n34 VSS.t13 40.5531
R69 VSS.n216 VSS.t56 31.3007
R70 VSS.n146 VSS.t5 21.225
R71 VSS.n201 VSS.t80 20.8673
R72 VSS.n135 VSS.t14 18.5719
R73 VSS.n64 VSS.t23 17.3802
R74 VSS.n104 VSS.t42 17.3802
R75 VSS.n49 VSS.t74 11.587
R76 VSS.n119 VSS.t11 11.587
R77 VSS.n181 VSS.n168 9.13939
R78 VSS.n181 VSS.n180 9.13939
R79 VSS.n248 VSS.n246 9.13939
R80 VSS.n6 VSS.t62 7.04085
R81 VSS.n239 VSS.t77 6.9078
R82 VSS.n173 VSS.n171 6.68085
R83 VSS.n173 VSS.n172 6.68085
R84 VSS.n182 VSS.n169 6.67693
R85 VSS.n178 VSS.n177 6.36078
R86 VSS VSS.n112 4.66717
R87 VSS.n211 VSS 4.66717
R88 VSS.n59 VSS 4.66717
R89 VSS.n114 VSS 4.47272
R90 VSS VSS.n209 4.47272
R91 VSS VSS.n57 4.47272
R92 VSS.n89 VSS.n88 4.29799
R93 VSS.n5 VSS.n2 4.29732
R94 VSS.n36 VSS.n33 4.29732
R95 VSS.n177 VSS.n176 4.25879
R96 VSS.n16 VSS.n1 3.76485
R97 VSS.n90 VSS.n82 3.76289
R98 VSS.n90 VSS.n84 3.76289
R99 VSS.n103 VSS.n78 3.76289
R100 VSS.n103 VSS.n80 3.76289
R101 VSS.n149 VSS.n74 3.76289
R102 VSS.n149 VSS.n76 3.76289
R103 VSS.n67 VSS.n28 3.76289
R104 VSS.n67 VSS.n30 3.76289
R105 VSS.n232 VSS.n23 3.76289
R106 VSS.n219 VSS.n164 3.76289
R107 VSS.n250 VSS.n20 3.6318
R108 VSS.n84 VSS.t3 3.2765
R109 VSS.n84 VSS.n83 3.2765
R110 VSS.n82 VSS.t81 3.2765
R111 VSS.n82 VSS.n81 3.2765
R112 VSS.n80 VSS.t82 3.2765
R113 VSS.n80 VSS.n79 3.2765
R114 VSS.n78 VSS.t64 3.2765
R115 VSS.n78 VSS.n77 3.2765
R116 VSS.n76 VSS.t6 3.2765
R117 VSS.n76 VSS.n75 3.2765
R118 VSS.n74 VSS.t33 3.2765
R119 VSS.n74 VSS.n73 3.2765
R120 VSS.n30 VSS.t16 3.2765
R121 VSS.n30 VSS.n29 3.2765
R122 VSS.n28 VSS.t45 3.2765
R123 VSS.n28 VSS.n27 3.2765
R124 VSS.n23 VSS.t84 3.2765
R125 VSS.n23 VSS.n22 3.2765
R126 VSS.n164 VSS.t47 3.2765
R127 VSS.n164 VSS.n163 3.2765
R128 VSS.n1 VSS.t71 3.2765
R129 VSS.n1 VSS.n0 3.2765
R130 VSS.n20 VSS.t41 3.2765
R131 VSS.n20 VSS.n19 3.2765
R132 VSS.n174 VSS.n173 2.61175
R133 VSS.n66 VSS.n65 2.6005
R134 VSS.n65 VSS.n64 2.6005
R135 VSS.n63 VSS.n62 2.6005
R136 VSS.n62 VSS.n61 2.6005
R137 VSS.n60 VSS.n59 2.6005
R138 VSS.n59 VSS.n58 2.6005
R139 VSS.n57 VSS.n55 2.6005
R140 VSS.n57 VSS.n56 2.6005
R141 VSS.n54 VSS.n53 2.6005
R142 VSS.n53 VSS.n52 2.6005
R143 VSS.n51 VSS.n50 2.6005
R144 VSS.n50 VSS.n49 2.6005
R145 VSS.n48 VSS.n47 2.6005
R146 VSS.n47 VSS.n46 2.6005
R147 VSS.n45 VSS.n44 2.6005
R148 VSS.n44 VSS.n43 2.6005
R149 VSS.n42 VSS.n41 2.6005
R150 VSS.n41 VSS.n40 2.6005
R151 VSS.n39 VSS.n38 2.6005
R152 VSS.n38 VSS.n37 2.6005
R153 VSS.n35 VSS.n34 2.6005
R154 VSS.n70 VSS.n69 2.6005
R155 VSS.n69 VSS.n68 2.6005
R156 VSS.n170 VSS 2.6005
R157 VSS.n175 VSS.n174 2.6005
R158 VSS.n194 VSS.n166 2.6005
R159 VSS.n166 VSS.n165 2.6005
R160 VSS.n193 VSS.n192 2.6005
R161 VSS.n192 VSS.n191 2.6005
R162 VSS.n190 VSS.n189 2.6005
R163 VSS.n189 VSS.n188 2.6005
R164 VSS.n187 VSS.n186 2.6005
R165 VSS.n186 VSS.n185 2.6005
R166 VSS.n183 VSS.n168 2.6005
R167 VSS.n168 VSS.n167 2.6005
R168 VSS VSS.n181 2.6005
R169 VSS.n181 VSS.t50 2.6005
R170 VSS.n180 VSS.n178 2.6005
R171 VSS.n180 VSS.n179 2.6005
R172 VSS.n222 VSS.n221 2.6005
R173 VSS.n221 VSS.n220 2.6005
R174 VSS.n218 VSS.n217 2.6005
R175 VSS.n217 VSS.n216 2.6005
R176 VSS.n215 VSS.n214 2.6005
R177 VSS.n214 VSS.n213 2.6005
R178 VSS.n212 VSS.n211 2.6005
R179 VSS.n211 VSS.n210 2.6005
R180 VSS.n209 VSS.n207 2.6005
R181 VSS.n209 VSS.n208 2.6005
R182 VSS.n206 VSS.n205 2.6005
R183 VSS.n205 VSS.n204 2.6005
R184 VSS.n203 VSS.n202 2.6005
R185 VSS.n202 VSS.n201 2.6005
R186 VSS.n200 VSS.n199 2.6005
R187 VSS.n199 VSS.n198 2.6005
R188 VSS.n197 VSS.n196 2.6005
R189 VSS.n196 VSS.n195 2.6005
R190 VSS.n238 VSS.n237 2.6005
R191 VSS.n237 VSS.n236 2.6005
R192 VSS.n235 VSS.n234 2.6005
R193 VSS.n234 VSS.n233 2.6005
R194 VSS.n231 VSS.n230 2.6005
R195 VSS.n230 VSS.n229 2.6005
R196 VSS.n228 VSS.n227 2.6005
R197 VSS.n227 VSS.n226 2.6005
R198 VSS.n131 VSS.n130 2.6005
R199 VSS.n130 VSS.n129 2.6005
R200 VSS.n134 VSS.n133 2.6005
R201 VSS.n133 VSS.n132 2.6005
R202 VSS.n137 VSS.n136 2.6005
R203 VSS.n136 VSS.n135 2.6005
R204 VSS.n140 VSS.n139 2.6005
R205 VSS.n139 VSS.n138 2.6005
R206 VSS.n145 VSS.n144 2.6005
R207 VSS.n144 VSS.n143 2.6005
R208 VSS.n148 VSS.n147 2.6005
R209 VSS.n147 VSS.n146 2.6005
R210 VSS.n152 VSS.n151 2.6005
R211 VSS.n151 VSS.n150 2.6005
R212 VSS.n155 VSS.n154 2.6005
R213 VSS.n154 VSS.n153 2.6005
R214 VSS.n86 VSS.n85 2.6005
R215 VSS.n93 VSS.n92 2.6005
R216 VSS.n92 VSS.n91 2.6005
R217 VSS.n96 VSS.n95 2.6005
R218 VSS.n95 VSS.n94 2.6005
R219 VSS.n99 VSS.n98 2.6005
R220 VSS.n98 VSS.n97 2.6005
R221 VSS.n102 VSS.n101 2.6005
R222 VSS.n101 VSS.n100 2.6005
R223 VSS.n106 VSS.n105 2.6005
R224 VSS.n105 VSS.n104 2.6005
R225 VSS.n109 VSS.n108 2.6005
R226 VSS.n108 VSS.n107 2.6005
R227 VSS.n112 VSS.n110 2.6005
R228 VSS.n112 VSS.n111 2.6005
R229 VSS.n115 VSS.n114 2.6005
R230 VSS.n114 VSS.n113 2.6005
R231 VSS.n118 VSS.n117 2.6005
R232 VSS.n117 VSS.n116 2.6005
R233 VSS.n121 VSS.n120 2.6005
R234 VSS.n120 VSS.n119 2.6005
R235 VSS.n124 VSS.n123 2.6005
R236 VSS.n123 VSS.n122 2.6005
R237 VSS.n128 VSS.n127 2.6005
R238 VSS.n127 VSS.n126 2.6005
R239 VSS.n240 VSS.n21 2.6005
R240 VSS.n141 VSS.n21 2.6005
R241 VSS.n253 VSS.n252 2.6005
R242 VSS.n252 VSS.n251 2.6005
R243 VSS.n249 VSS.n248 2.6005
R244 VSS.n248 VSS.n247 2.6005
R245 VSS.n246 VSS.n244 2.6005
R246 VSS.n246 VSS.n245 2.6005
R247 VSS.n243 VSS.n242 2.6005
R248 VSS.n242 VSS.n241 2.6005
R249 VSS.n256 VSS.n255 2.6005
R250 VSS.n255 VSS.n254 2.6005
R251 VSS.n257 VSS.n18 2.6005
R252 VSS.n18 VSS.n17 2.6005
R253 VSS.n4 VSS.n3 2.6005
R254 VSS.n9 VSS.n8 2.6005
R255 VSS.n8 VSS.n7 2.6005
R256 VSS.n12 VSS.n11 2.6005
R257 VSS.n11 VSS.n10 2.6005
R258 VSS.n15 VSS.n14 2.6005
R259 VSS.n14 VSS.n13 2.6005
R260 VSS VSS.n271 2.6005
R261 VSS.n271 VSS.n270 2.6005
R262 VSS.n269 VSS.n268 2.6005
R263 VSS.n268 VSS.n267 2.6005
R264 VSS.n266 VSS.n265 2.6005
R265 VSS.n265 VSS.n264 2.6005
R266 VSS.n263 VSS.n262 2.6005
R267 VSS.n262 VSS.n261 2.6005
R268 VSS.n260 VSS.n259 2.6005
R269 VSS.n259 VSS.n258 2.6005
R270 VSS.n72 VSS.n26 2.41287
R271 VSS.n26 VSS.n25 2.41287
R272 VSS.n224 VSS.n162 2.41287
R273 VSS.n162 VSS.n161 2.41287
R274 VSS.n157 VSS.n156 2.24619
R275 VSS.n176 VSS.n170 1.65822
R276 VSS.n89 VSS.n86 1.64953
R277 VSS.n36 VSS.n35 1.64943
R278 VSS.n5 VSS.n4 1.64943
R279 VSS.n159 VSS.n158 1.59484
R280 VSS.n225 VSS.n160 1.49673
R281 VSS.n145 VSS.n140 0.631304
R282 VSS.n187 VSS.n183 0.595946
R283 VSS.n39 VSS.n36 0.559135
R284 VSS.n6 VSS.n5 0.541457
R285 VSS.n90 VSS.n89 0.535268
R286 VSS VSS.n238 0.489511
R287 VSS.n176 VSS.n175 0.472687
R288 VSS.n257 VSS.n256 0.41675
R289 VSS.n239 VSS 0.15145
R290 VSS.n96 VSS.n93 0.0760357
R291 VSS.n99 VSS.n96 0.0760357
R292 VSS.n102 VSS.n99 0.0760357
R293 VSS.n109 VSS.n106 0.0760357
R294 VSS.n110 VSS.n109 0.0760357
R295 VSS.n115 VSS.n110 0.0760357
R296 VSS.n118 VSS.n115 0.0760357
R297 VSS.n121 VSS.n118 0.0760357
R298 VSS.n124 VSS.n121 0.0760357
R299 VSS.n128 VSS.n124 0.0760357
R300 VSS.n131 VSS.n128 0.0760357
R301 VSS.n134 VSS.n131 0.0760357
R302 VSS.n137 VSS.n134 0.0760357
R303 VSS.n140 VSS.n137 0.0760357
R304 VSS.n148 VSS.n145 0.0760357
R305 VSS.n155 VSS.n152 0.0760357
R306 VSS.n66 VSS.n63 0.0760357
R307 VSS.n63 VSS.n60 0.0760357
R308 VSS.n60 VSS.n55 0.0760357
R309 VSS.n55 VSS.n54 0.0760357
R310 VSS.n54 VSS.n51 0.0760357
R311 VSS.n51 VSS.n48 0.0760357
R312 VSS.n48 VSS.n45 0.0760357
R313 VSS.n45 VSS.n42 0.0760357
R314 VSS.n42 VSS.n39 0.0760357
R315 VSS.n177 VSS 0.0760357
R316 VSS.n238 VSS.n235 0.0760357
R317 VSS.n231 VSS.n228 0.0760357
R318 VSS.n218 VSS.n215 0.0760357
R319 VSS.n215 VSS.n212 0.0760357
R320 VSS.n212 VSS.n207 0.0760357
R321 VSS.n207 VSS.n206 0.0760357
R322 VSS.n206 VSS.n203 0.0760357
R323 VSS.n203 VSS.n200 0.0760357
R324 VSS.n200 VSS.n197 0.0760357
R325 VSS.n197 VSS.n194 0.0760357
R326 VSS.n194 VSS.n193 0.0760357
R327 VSS.n193 VSS.n190 0.0760357
R328 VSS.n190 VSS.n187 0.0760357
R329 VSS.n12 VSS.n9 0.0760357
R330 VSS.n15 VSS.n12 0.0760357
R331 VSS VSS.n269 0.0760357
R332 VSS.n269 VSS.n266 0.0760357
R333 VSS.n266 VSS.n263 0.0760357
R334 VSS.n263 VSS.n260 0.0760357
R335 VSS.n260 VSS.n257 0.0760357
R336 VSS.n256 VSS.n253 0.0760357
R337 VSS.n244 VSS.n243 0.0760357
R338 VSS.n243 VSS.n240 0.0760357
R339 VSS VSS.n178 0.0747105
R340 VSS.n16 VSS.n15 0.0712143
R341 VSS.n228 VSS.n225 0.0700705
R342 VSS.n106 VSS.n103 0.0696071
R343 VSS.n67 VSS.n66 0.0696071
R344 VSS.n219 VSS.n218 0.0696071
R345 VSS.n156 VSS.n155 0.0668722
R346 VSS.n71 VSS.n70 0.0664687
R347 VSS.n223 VSS.n222 0.0664464
R348 VSS.n173 VSS 0.0647857
R349 VSS.n182 VSS 0.0636579
R350 VSS.n149 VSS.n148 0.0519286
R351 VSS.n235 VSS.n232 0.0519286
R352 VSS.n253 VSS.n250 0.0495179
R353 VSS.n244 VSS 0.0446964
R354 VSS.n249 VSS 0.0318393
R355 VSS.n250 VSS.n249 0.0270179
R356 VSS.n93 VSS.n90 0.0246071
R357 VSS.n152 VSS.n149 0.0246071
R358 VSS.n232 VSS.n231 0.0246071
R359 VSS.n160 VSS.n159 0.0197857
R360 VSS.n9 VSS.n6 0.0181786
R361 VSS.n183 VSS.n182 0.0115526
R362 VSS.n224 VSS.n223 0.0110446
R363 VSS.n158 VSS.n157 0.0110437
R364 VSS.n72 VSS.n71 0.0110223
R365 VSS.n156 VSS.n72 0.0106222
R366 VSS.n225 VSS.n224 0.00741026
R367 VSS.n103 VSS.n102 0.00692857
R368 VSS.n70 VSS.n67 0.00692857
R369 VSS.n222 VSS.n219 0.00692857
R370 VSS VSS.n16 0.00532143
R371 VSS.n240 VSS.n239 0.00451786
R372 B.t8 B.t12 55.0112
R373 B.t3 B.t9 55.0112
R374 B.t0 B.t2 55.0112
R375 B.n2 B.t10 34.6755
R376 B.n5 B.t7 29.9826
R377 B.n3 B.t4 29.9826
R378 B.n0 B.t13 29.9826
R379 B B.n4 27.1952
R380 B B.n1 27.1952
R381 B.n7 B.n6 25.905
R382 B.n6 B.t1 22.5523
R383 B.n4 B.t11 22.5523
R384 B.n1 B.t5 22.5523
R385 B B.n2 17.6692
R386 B.n2 B.t6 13.0362
R387 B.n5 B.t8 9.1255
R388 B.n3 B.t3 9.1255
R389 B.n0 B.t0 9.1255
R390 B.n8 B.n7 9.08249
R391 B.n6 B.n5 7.43086
R392 B.n4 B.n3 7.43086
R393 B.n1 B.n0 7.43086
R394 B.n9 B 4.35984
R395 B.n9 B.n8 3.06371
R396 B.n10 B.n9 2.6555
R397 B B.n10 1.07086
R398 B.n8 B 0.2255
R399 B.n7 B 0.171539
R400 B.n10 B 0.0771537
R401 VDD.n67 VDD.n66 1387.55
R402 VDD.n65 VDD.n47 804.168
R403 VDD.n66 VDD.n65 791.668
R404 VDD.n128 VDD.t66 611.386
R405 VDD.n138 VDD.t51 611.386
R406 VDD.n138 VDD.t31 611.386
R407 VDD.n160 VDD.n159 181.468
R408 VDD.n150 VDD.n125 181.468
R409 VDD.t40 VDD.n55 179.732
R410 VDD.t40 VDD.n56 179.732
R411 VDD.n86 VDD.n85 159.053
R412 VDD.n94 VDD.n31 159.053
R413 VDD.t25 VDD.n158 154.44
R414 VDD.n158 VDD.t54 154.44
R415 VDD.n87 VDD.t13 145.517
R416 VDD.n47 VDD.t0 129.167
R417 VDD.n55 VDD.t36 126.195
R418 VDD.n87 VDD.t62 125.213
R419 VDD.n66 VDD.t2 120.834
R420 VDD.n114 VDD.n101 104.677
R421 VDD.n112 VDD.n102 104.677
R422 VDD.n160 VDD.t20 100.386
R423 VDD.n150 VDD.t44 100.386
R424 VDD.n79 VDD.n78 96.8079
R425 VDD.t17 VDD.n113 89.0874
R426 VDD.n113 VDD.t56 89.0874
R427 VDD.n4 VDD.t69 85.6385
R428 VDD.n95 VDD.t58 84.1628
R429 VDD.t20 VDD.n11 84.0493
R430 VDD.t44 VDD.n149 84.0493
R431 VDD.n166 VDD.t28 84.0493
R432 VDD.n46 VDD.t64 82.3898
R433 VDD.n85 VDD.t12 80.2579
R434 VDD.t58 VDD.n94 77.8347
R435 VDD.n66 VDD.n46 66.9418
R436 VDD.t36 VDD.n54 58.0938
R437 VDD.n101 VDD.t7 57.907
R438 VDD.t9 VDD.n102 57.907
R439 VDD.t14 VDD.n77 53.5535
R440 VDD.n56 VDD.n47 53.5378
R441 VDD.n77 VDD.t22 52.5237
R442 VDD.n108 VDD.t9 51.2582
R443 VDD.n78 VDD.t12 50.4639
R444 VDD.t7 VDD.n100 49.621
R445 VDD.t22 VDD.n76 44.2847
R446 VDD.n79 VDD.t14 43.2549
R447 VDD.t62 VDD.n31 33.8415
R448 VDD.n159 VDD.t25 27.0275
R449 VDD.n125 VDD.t54 27.0275
R450 VDD.n6 VDD.t38 27.0275
R451 VDD.n173 VDD.t49 27.0275
R452 VDD.n114 VDD.t17 15.5907
R453 VDD.t56 VDD.n112 15.5907
R454 VDD.n76 VDD.t64 14.4186
R455 VDD.n66 VDD.t4 14.3978
R456 VDD.t13 VDD.n86 13.5369
R457 VDD.n164 VDD.n11 10.8994
R458 VDD.n149 VDD.n148 10.8986
R459 VDD.n96 VDD.n95 10.837
R460 VDD.n100 VDD.n99 10.5918
R461 VDD.n84 VDD.n37 9.363
R462 VDD.n144 VDD.n143 8.2255
R463 VDD.n162 VDD.n161 8.2255
R464 VDD.n161 VDD.n13 8.2255
R465 VDD.n157 VDD.n13 8.2255
R466 VDD.n157 VDD.n14 8.2255
R467 VDD.n151 VDD.n14 8.2255
R468 VDD.n151 VDD.n124 8.2255
R469 VDD.n132 VDD.n131 8.2255
R470 VDD.n28 VDD.n26 8.2255
R471 VDD.n115 VDD.n26 8.2255
R472 VDD.n115 VDD.n27 8.2255
R473 VDD.n111 VDD.n27 8.2255
R474 VDD.n111 VDD.n103 8.2255
R475 VDD.n57 VDD.n53 8.2255
R476 VDD.n57 VDD.n49 8.2255
R477 VDD.n63 VDD.n49 8.2255
R478 VDD.n48 VDD.n45 8.2255
R479 VDD.n68 VDD.n40 8.2255
R480 VDD.n75 VDD.n40 8.2255
R481 VDD.n75 VDD.n39 8.2255
R482 VDD.n80 VDD.n39 8.2255
R483 VDD.n80 VDD.n37 8.2255
R484 VDD.n84 VDD.n36 8.2255
R485 VDD.n88 VDD.n36 8.2255
R486 VDD.n88 VDD.n32 8.2255
R487 VDD.n93 VDD.n32 8.2255
R488 VDD.n93 VDD.n30 8.2255
R489 VDD.n141 VDD.n140 6.01764
R490 VDD.n137 VDD.n136 4.98375
R491 VDD.n141 VDD.n129 4.93474
R492 VDD.n140 VDD.n139 4.93474
R493 VDD.n147 VDD.n126 4.93474
R494 VDD.n70 VDD.n41 4.88224
R495 VDD.n136 VDD.n133 4.7942
R496 VDD.n136 VDD.n134 4.7942
R497 VDD.n146 VDD.n127 4.7942
R498 VDD.n61 VDD.t1 4.7492
R499 VDD.n155 VDD.n19 4.5005
R500 VDD.n156 VDD.n155 4.5005
R501 VDD.n135 VDD.n132 3.1505
R502 VDD.n131 VDD.n130 3.1505
R503 VDD.n55 VDD.n53 3.1505
R504 VDD VDD.n57 3.1505
R505 VDD.n57 VDD.t40 3.1505
R506 VDD.n58 VDD.n49 3.1505
R507 VDD.n56 VDD.n49 3.1505
R508 VDD.n63 VDD.n62 3.1505
R509 VDD.n60 VDD.n48 3.1505
R510 VDD.n59 VDD.n45 3.1505
R511 VDD.n69 VDD.n68 3.1505
R512 VDD VDD.n40 3.1505
R513 VDD.n46 VDD.n40 3.1505
R514 VDD.n75 VDD.n74 3.1505
R515 VDD.n76 VDD.n75 3.1505
R516 VDD.n39 VDD.n38 3.1505
R517 VDD.n77 VDD.n39 3.1505
R518 VDD.n81 VDD.n80 3.1505
R519 VDD.n80 VDD.n79 3.1505
R520 VDD.n82 VDD.n37 3.1505
R521 VDD.n78 VDD.n37 3.1505
R522 VDD.n84 VDD.n83 3.1505
R523 VDD.n85 VDD.n84 3.1505
R524 VDD.n36 VDD.n35 3.1505
R525 VDD.n86 VDD.n36 3.1505
R526 VDD.n89 VDD.n88 3.1505
R527 VDD.n88 VDD.n87 3.1505
R528 VDD.n90 VDD.n32 3.1505
R529 VDD.n32 VDD.n31 3.1505
R530 VDD.n93 VDD.n92 3.1505
R531 VDD.n94 VDD.n93 3.1505
R532 VDD.n30 VDD.n29 3.1505
R533 VDD.n103 VDD.n102 3.1505
R534 VDD.n98 VDD.n28 3.1505
R535 VDD.n97 VDD.n26 3.1505
R536 VDD.n101 VDD.n26 3.1505
R537 VDD.n116 VDD.n115 3.1505
R538 VDD.n115 VDD.n114 3.1505
R539 VDD.n111 VDD.n110 3.1505
R540 VDD.n112 VDD.n111 3.1505
R541 VDD.n3 VDD.n2 3.1505
R542 VDD.n8 VDD.n7 3.1505
R543 VDD.n7 VDD.n6 3.1505
R544 VDD VDD.n177 3.1505
R545 VDD.n177 VDD.n176 3.1505
R546 VDD.n175 VDD.n174 3.1505
R547 VDD.n174 VDD.n173 3.1505
R548 VDD.n171 VDD.n170 3.1505
R549 VDD.n170 VDD.n169 3.1505
R550 VDD.n168 VDD.n167 3.1505
R551 VDD.n163 VDD.n162 3.1505
R552 VDD.n161 VDD.n12 3.1505
R553 VDD.n161 VDD.n160 3.1505
R554 VDD.n18 VDD.n13 3.1505
R555 VDD.n159 VDD.n13 3.1505
R556 VDD.n154 VDD.n14 3.1505
R557 VDD.n125 VDD.n14 3.1505
R558 VDD.n152 VDD.n151 3.1505
R559 VDD.n151 VDD.n150 3.1505
R560 VDD.n124 VDD.n123 3.1505
R561 VDD.n145 VDD.n144 3.1505
R562 VDD.n143 VDD.n142 3.1505
R563 VDD.n91 VDD.n34 3.06224
R564 VDD.n52 VDD.n51 2.9292
R565 VDD.n44 VDD.n43 2.91941
R566 VDD.n25 VDD.n22 2.91941
R567 VDD.n25 VDD.n24 2.91941
R568 VDD.n17 VDD.n16 2.91941
R569 VDD.n5 VDD.n1 2.91941
R570 VDD.n73 VDD.n72 2.91705
R571 VDD.n109 VDD.n107 2.91705
R572 VDD.n109 VDD.n105 2.91705
R573 VDD.n153 VDD.n122 2.91705
R574 VDD.n172 VDD.n10 2.91705
R575 VDD.n27 VDD 2.6255
R576 VDD.n113 VDD.n27 2.6255
R577 VDD.n157 VDD 2.6255
R578 VDD.n158 VDD.n157 2.6255
R579 VDD.n119 VDD 2.2512
R580 VDD.n118 VDD.n117 2.24619
R581 VDD.n118 VDD.n20 2.24599
R582 VDD.n108 VDD.n103 1.87673
R583 VDD.n54 VDD.n53 1.87118
R584 VDD.n4 VDD.n3 1.8711
R585 VDD.n43 VDD.t3 1.8205
R586 VDD.n43 VDD.n42 1.8205
R587 VDD.n72 VDD.t65 1.8205
R588 VDD.n72 VDD.n71 1.8205
R589 VDD.n24 VDD.t71 1.8205
R590 VDD.n24 VDD.n23 1.8205
R591 VDD.n22 VDD.t8 1.8205
R592 VDD.n22 VDD.n21 1.8205
R593 VDD.n107 VDD.t61 1.8205
R594 VDD.n107 VDD.n106 1.8205
R595 VDD.n105 VDD.t57 1.8205
R596 VDD.n105 VDD.n104 1.8205
R597 VDD.n34 VDD.t63 1.8205
R598 VDD.n34 VDD.n33 1.8205
R599 VDD.n51 VDD.t37 1.8205
R600 VDD.n51 VDD.n50 1.8205
R601 VDD.n122 VDD.t55 1.8205
R602 VDD.n122 VDD.n121 1.8205
R603 VDD.n16 VDD.t21 1.8205
R604 VDD.n16 VDD.n15 1.8205
R605 VDD.n10 VDD.t50 1.8205
R606 VDD.n10 VDD.n9 1.8205
R607 VDD.n1 VDD.t70 1.8205
R608 VDD.n1 VDD.n0 1.8205
R609 VDD.n64 VDD.n63 1.7854
R610 VDD.n67 VDD.n45 1.7854
R611 VDD.n64 VDD.n48 1.78487
R612 VDD.n68 VDD.n67 1.78487
R613 VDD.n144 VDD.n126 1.78473
R614 VDD.n137 VDD.n132 1.78473
R615 VDD.n139 VDD.n131 1.78473
R616 VDD.n143 VDD.n129 1.78473
R617 VDD.n120 VDD.n119 1.61133
R618 VDD VDD.n120 1.12363
R619 VDD VDD.n164 0.961571
R620 VDD.n99 VDD.n96 0.771929
R621 VDD.n65 VDD.n64 0.684371
R622 VDD.n138 VDD.n137 0.684132
R623 VDD.n139 VDD.n138 0.684132
R624 VDD.n128 VDD.n126 0.684132
R625 VDD.n129 VDD.n128 0.684132
R626 VDD.n148 VDD.n147 0.615232
R627 VDD.n5 VDD.n4 0.590232
R628 VDD.n109 VDD.n108 0.582082
R629 VDD.n54 VDD.n52 0.578894
R630 VDD.n165 VDD 0.350054
R631 VDD.n100 VDD.n28 0.21859
R632 VDD.n95 VDD.n30 0.150263
R633 VDD.n162 VDD.n11 0.133436
R634 VDD.n167 VDD.n166 0.133193
R635 VDD.n149 VDD.n124 0.133193
R636 VDD.n83 VDD.n82 0.0864821
R637 VDD.n140 VDD.n130 0.0760357
R638 VDD.n58 VDD 0.0760357
R639 VDD.n62 VDD.n58 0.0760357
R640 VDD.n60 VDD.n59 0.0760357
R641 VDD VDD.n69 0.0760357
R642 VDD.n81 VDD.n38 0.0760357
R643 VDD.n82 VDD.n81 0.0760357
R644 VDD.n89 VDD.n35 0.0760357
R645 VDD.n90 VDD.n89 0.0760357
R646 VDD.n92 VDD.n29 0.0760357
R647 VDD.n96 VDD.n29 0.0760357
R648 VDD.n99 VDD.n98 0.0760357
R649 VDD.n98 VDD.n97 0.0760357
R650 VDD VDD.n8 0.0760357
R651 VDD VDD.n175 0.0760357
R652 VDD.n171 VDD.n168 0.0760357
R653 VDD.n168 VDD.n165 0.0760357
R654 VDD.n164 VDD.n163 0.0760357
R655 VDD.n163 VDD.n12 0.0760357
R656 VDD.n152 VDD.n123 0.0760357
R657 VDD.n148 VDD.n123 0.0760357
R658 VDD.n142 VDD.n141 0.0760357
R659 VDD.n117 VDD.n116 0.0668722
R660 VDD.n110 VDD.n20 0.0664687
R661 VDD VDD.n52 0.0647857
R662 VDD.n19 VDD.n18 0.05675
R663 VDD.n156 VDD.n154 0.0559464
R664 VDD.n74 VDD.n73 0.0551429
R665 VDD.n110 VDD.n109 0.0551429
R666 VDD.n175 VDD.n172 0.0551429
R667 VDD.n154 VDD.n153 0.0551429
R668 VDD.n69 VDD.n44 0.0535357
R669 VDD.n116 VDD.n25 0.0535357
R670 VDD.n8 VDD.n5 0.0535357
R671 VDD.n18 VDD.n17 0.0535357
R672 VDD.n147 VDD.n146 0.0495179
R673 VDD.n91 VDD.n90 0.0487143
R674 VDD.n70 VDD 0.0463036
R675 VDD.n62 VDD.n61 0.0422857
R676 VDD.n135 VDD 0.0382679
R677 VDD VDD.n130 0.0382679
R678 VDD.n83 VDD 0.0382679
R679 VDD VDD.n35 0.0382679
R680 VDD.n145 VDD 0.0382679
R681 VDD.n142 VDD 0.0382679
R682 VDD.n61 VDD.n60 0.03425
R683 VDD.n74 VDD.n70 0.0302321
R684 VDD.n92 VDD.n91 0.0278214
R685 VDD.n136 VDD.n135 0.0270179
R686 VDD.n146 VDD.n145 0.0270179
R687 VDD.n59 VDD.n44 0.023
R688 VDD.n97 VDD.n25 0.023
R689 VDD.n17 VDD.n12 0.023
R690 VDD.n73 VDD.n38 0.0213929
R691 VDD.n172 VDD.n171 0.0213929
R692 VDD.n153 VDD.n152 0.0213929
R693 VDD VDD.n156 0.0205893
R694 VDD VDD.n19 0.0197857
R695 VDD.n20 VDD 0.0110223
R696 VDD.n119 VDD.n118 0.0106437
R697 VDD.n117 VDD 0.0106222
R698 VDD.n155 VDD.n120 0.00663296
R699 S3.n2 S3.n0 7.06041
R700 S3.n2 S3.n1 5.46137
R701 S3 S3.n2 0.196152
R702 S4.n2 S4.n0 7.06041
R703 S4.n2 S4.n1 5.46137
R704 S4 S4.n2 0.17869
R705 A.t17 A.t5 68.5684
R706 A.n3 A.t0 39.6291
R707 A.n12 A.t6 39.6291
R708 A.n1 A.t12 39.6291
R709 A.n9 A.n8 35.9467
R710 A.n5 A.t2 34.6755
R711 A.n2 A.t8 29.9826
R712 A.t7 A.n2 29.9826
R713 A.n7 A.t17 29.9826
R714 A.n11 A.t16 29.9826
R715 A.t4 A.n11 29.9826
R716 A.n0 A.t3 29.9826
R717 A.t11 A.n0 29.9826
R718 A.n3 A.t7 28.9398
R719 A.n12 A.t4 28.9398
R720 A.n1 A.t11 28.9398
R721 A A.n3 21.7803
R722 A A.n12 21.7803
R723 A A.n1 21.7803
R724 A.n8 A.n7 20.8576
R725 A A.n5 17.6692
R726 A.n5 A.t13 13.0362
R727 A.n10 A.n9 11.7535
R728 A.n2 A.t1 9.1255
R729 A.n8 A.t10 9.1255
R730 A.n7 A.t15 9.1255
R731 A.n11 A.t9 9.1255
R732 A.n0 A.t14 9.1255
R733 A.n4 A 4.02486
R734 A A.n13 3.8705
R735 A.n4 A 2.66023
R736 A.n13 A 2.65229
R737 A.n6 A 2.58311
R738 A.n10 A.n6 0.996929
R739 A.n13 A.n10 0.689964
R740 A.n6 A.n4 0.194964
R741 A.n9 A 0.194521
R742 S6.n3 S6.n0 7.06041
R743 S6.n2 S6 6.56414
R744 S6.n2 S6.n1 5.18354
R745 S6.n3 S6.n2 0.21963
R746 S6 S6.n3 0.196152
R747 S1.n2 S1.n0 7.06041
R748 S1.n2 S1.n1 5.10528
R749 S1 S1.n2 0.0533261
R750 S2.n2 S2.n0 7.06041
R751 S2.n2 S2.n1 5.46137
R752 S2 S2.n2 0.196152
R753 S5.n2 S5 8.45295
R754 S5.n3 S5.n0 7.03107
R755 S5.n2 S5.n1 5.4242
R756 S5 S5.n3 0.169894
R757 S5.n3 S5.n2 0.00523684
C0 VDD S4 0.357f
C1 a_3303_n1718# AND_3_In_Layout_1.C 0.00246f
C2 A VDD 1.32f
C3 OR_2_In_Layout_0.B S5 0.0819f
C4 a_801_375# S4 8.72e-19
C5 a_801_375# A 0.387f
C6 B a_3184_375# 0.0405f
C7 C a_2999_n1346# 0.00286f
C8 B a_801_n1645# 2.21e-19
C9 S4 a_3303_n1718# 0.00472f
C10 B a_801_n363# 0.0623f
C11 S3 a_3184_n363# 0.259f
C12 a_3328_375# a_3184_375# 0.343f
C13 a_945_n1645# a_1425_n1645# 0.248f
C14 A a_3303_n1718# 0.00339f
C15 AND_2_In_Layout_0.A OR_2_In_Layout_0.A 0.00426f
C16 A a_1425_n363# 0.00379f
C17 AND_2_In_Layout_0.A AND_3_In_Layout_1.C 0.0481f
C18 OR_2_In_Layout_0.A AND_3_In_Layout_1.C 0.0466f
C19 B a_945_n1645# 3.19e-20
C20 B OR_2_In_Layout_0.B 0.0696f
C21 VDD S2 0.147f
C22 VDD S5 0.319f
C23 A AND_2_In_Layout_0.A 0.00443f
C24 VDD a_945_375# 0.0453f
C25 OR_2_In_Layout_0.B a_3328_375# 3.07e-19
C26 S4 OR_2_In_Layout_0.A 0.0415f
C27 A OR_2_In_Layout_0.A 1.22f
C28 S3 a_3808_n363# 0.0155f
C29 C a_1425_375# 0.0543f
C30 a_801_375# S5 0.0114f
C31 a_3184_n363# a_801_n363# 2.33e-19
C32 a_801_375# a_945_375# 0.343f
C33 S4 AND_3_In_Layout_1.C 0.0324f
C34 VDD a_1425_n1645# 0.0054f
C35 A AND_3_In_Layout_1.C 0.321f
C36 VDD a_3808_375# 0.00487f
C37 a_1425_375# S6 0.0155f
C38 a_1425_n363# S5 0.0172f
C39 S3 a_4292_n1650# 7.29e-19
C40 A S4 0.0223f
C41 B VDD 0.838f
C42 a_3184_n363# OR_2_In_Layout_0.B 0.294f
C43 C a_3184_375# 0.299f
C44 C a_801_n1645# 0.154f
C45 VDD a_3328_375# 6.85e-19
C46 a_801_375# B 0.0705f
C47 C a_801_n363# 0.00124f
C48 S1 a_4148_n1650# 0.0273f
C49 a_3184_375# S6 0.0162f
C50 a_801_375# a_3328_375# 7.18e-20
C51 a_945_n363# a_801_n363# 0.343f
C52 S5 OR_2_In_Layout_0.A 0.035f
C53 B a_1425_n363# 0.0405f
C54 a_801_n363# S6 3.82e-19
C55 S2 AND_3_In_Layout_1.C 0.0889f
C56 S5 AND_3_In_Layout_1.C 0.0391f
C57 a_945_375# AND_3_In_Layout_1.C 0.00869f
C58 a_1425_n1645# OR_2_In_Layout_0.A 0.0513f
C59 C a_945_n1645# 0.01f
C60 C OR_2_In_Layout_0.B 1.86f
C61 a_3328_n363# a_801_n363# 7.18e-20
C62 OR_2_In_Layout_0.B a_3808_n363# 0.00131f
C63 VDD a_3184_n363# 0.711f
C64 a_3808_375# AND_3_In_Layout_1.C 0.0723f
C65 VDD a_4148_n1650# 0.0116f
C66 OR_2_In_Layout_0.B a_945_n363# 0.0035f
C67 OR_2_In_Layout_0.B S6 1.68e-19
C68 S4 S5 1.1f
C69 A S2 0.00246f
C70 B AND_2_In_Layout_0.A 1.75e-19
C71 A S5 0.0264f
C72 A a_945_375# 0.0604f
C73 a_801_n1645# a_2999_n1346# 2.96e-19
C74 B OR_2_In_Layout_0.A 0.115f
C75 S4 a_1425_n1645# 0.0155f
C76 a_4292_n1650# OR_2_In_Layout_0.B 2.25e-21
C77 a_3303_n1718# a_3184_n363# 2.98e-19
C78 A a_1425_n1645# 0.00131f
C79 OR_2_In_Layout_0.A a_3328_375# 7.68e-20
C80 B AND_3_In_Layout_1.C 0.534f
C81 A a_3808_375# 0.00663f
C82 a_3328_n363# OR_2_In_Layout_0.B 0.0502f
C83 a_3303_n1718# a_4148_n1650# 7.19e-19
C84 a_3328_375# AND_3_In_Layout_1.C 0.0143f
C85 a_4292_n1650# S1 0.0558f
C86 C VDD 2.8f
C87 VDD a_3808_n363# 0.00487f
C88 OR_2_In_Layout_0.B a_2999_n1346# 0.0408f
C89 B S4 0.0286f
C90 B A 1.67f
C91 VDD a_945_n363# 0.0473f
C92 VDD S6 0.332f
C93 a_801_375# C 0.114f
C94 S4 a_3328_375# 1.33e-19
C95 A a_3328_375# 0.00285f
C96 a_3184_n363# AND_2_In_Layout_0.A 0.00416f
C97 AND_2_In_Layout_0.A a_4148_n1650# 0.101f
C98 a_3184_n363# OR_2_In_Layout_0.A 0.0737f
C99 C a_3303_n1718# 8.7e-19
C100 a_801_375# S6 0.266f
C101 a_4148_n1650# OR_2_In_Layout_0.A 7.87e-19
C102 C a_1425_n363# 1.37e-19
C103 a_3303_n1718# a_3808_n363# 1.57e-19
C104 VDD a_4292_n1650# 0.537f
C105 VDD a_3328_n363# 6.85e-19
C106 a_3184_n363# AND_3_In_Layout_1.C 0.0129f
C107 a_4148_n1650# AND_3_In_Layout_1.C 0.055f
C108 a_1425_n363# a_945_n363# 0.248f
C109 a_3808_375# S2 0.0155f
C110 VDD a_2999_n1346# 0.792f
C111 a_4292_n1650# a_3303_n1718# 0.00149f
C112 S4 a_3184_n363# 3.37e-19
C113 A a_3184_n363# 0.133f
C114 OR_2_In_Layout_0.B a_1425_375# 1.37e-19
C115 C AND_2_In_Layout_0.A 2.89e-19
C116 A a_4148_n1650# 0.00194f
C117 C OR_2_In_Layout_0.A 0.292f
C118 B S2 1.47e-19
C119 B S5 0.036f
C120 B a_945_375# 0.44f
C121 a_801_n1645# a_801_n363# 0.0152f
C122 a_3808_n363# OR_2_In_Layout_0.A 0.0423f
C123 S3 S1 0.0314f
C124 S5 a_3328_375# 1.01e-19
C125 a_945_n363# OR_2_In_Layout_0.A 0.0319f
C126 C AND_3_In_Layout_1.C 0.0965f
C127 a_3303_n1718# a_2999_n1346# 0.293f
C128 OR_2_In_Layout_0.A S6 8.71e-20
C129 a_3808_n363# AND_3_In_Layout_1.C 0.00324f
C130 B a_1425_n1645# 9.88e-20
C131 B a_3808_375# 0.0405f
C132 S6 AND_3_In_Layout_1.C 0.0269f
C133 a_4292_n1650# AND_2_In_Layout_0.A 0.135f
C134 a_3808_375# a_3328_375# 0.248f
C135 a_4292_n1650# OR_2_In_Layout_0.A 8.96e-19
C136 a_945_n1645# a_801_n1645# 0.343f
C137 OR_2_In_Layout_0.B a_3184_375# 6.34e-20
C138 OR_2_In_Layout_0.B a_801_n1645# 0.0148f
C139 a_3328_n363# OR_2_In_Layout_0.A 0.42f
C140 C S4 1.28f
C141 C A 0.158f
C142 A a_3808_n363# 0.0679f
C143 OR_2_In_Layout_0.B a_801_n363# 0.128f
C144 VDD S3 0.244f
C145 a_4292_n1650# AND_3_In_Layout_1.C 0.0885f
C146 a_3328_n363# AND_3_In_Layout_1.C 0.00109f
C147 VDD a_1425_375# 0.0552f
C148 A a_945_n363# 0.0656f
C149 S4 S6 0.0231f
C150 A S6 0.0101f
C151 AND_2_In_Layout_0.A a_2999_n1346# 0.121f
C152 B a_3328_375# 0.206f
C153 a_3184_n363# S5 0.016f
C154 a_2999_n1346# OR_2_In_Layout_0.A 0.235f
C155 a_801_375# a_1425_375# 0.429f
C156 a_2999_n1346# AND_3_In_Layout_1.C 5.08e-19
C157 A a_4292_n1650# 0.00422f
C158 S4 a_3328_n363# 1.33e-19
C159 A a_3328_n363# 0.0185f
C160 VDD a_3184_375# 0.693f
C161 VDD a_801_n1645# 0.703f
C162 S4 a_2999_n1346# 0.0217f
C163 A a_2999_n1346# 0.00406f
C164 VDD a_801_n363# 0.806f
C165 B a_3184_n363# 3.97e-19
C166 C S2 1.38e-19
C167 a_801_375# a_3184_375# 2.33e-19
C168 C S5 0.086f
C169 C a_945_375# 0.002f
C170 S3 AND_2_In_Layout_0.A 3.8e-19
C171 a_3303_n1718# a_801_n1645# 4.47e-20
C172 S5 S6 0.693f
C173 S3 OR_2_In_Layout_0.A 6.27e-19
C174 C a_1425_n1645# 0.0637f
C175 C a_3808_375# 0.00222f
C176 a_1425_n363# a_801_n363# 0.429f
C177 VDD a_945_n1645# 0.00185f
C178 S3 AND_3_In_Layout_1.C 0.055f
C179 VDD OR_2_In_Layout_0.B 0.996f
C180 a_1425_375# AND_3_In_Layout_1.C 0.0134f
C181 a_3328_n363# S5 1.09e-19
C182 VDD S1 0.149f
C183 C B 0.425f
C184 A S3 0.0494f
C185 a_801_n1645# AND_2_In_Layout_0.A 2.64e-20
C186 a_3303_n1718# OR_2_In_Layout_0.B 0.108f
C187 a_1425_n363# OR_2_In_Layout_0.B 0.0587f
C188 A a_1425_375# 0.00234f
C189 C a_3328_375# 0.0526f
C190 a_3184_n363# a_4148_n1650# 2.4e-19
C191 B a_945_n363# 0.413f
C192 B S6 0.00132f
C193 a_801_n1645# OR_2_In_Layout_0.A 0.0448f
C194 a_801_n363# OR_2_In_Layout_0.A 0.0302f
C195 a_3328_375# S6 8.24e-21
C196 a_3303_n1718# S1 4.29e-20
C197 a_3184_375# AND_3_In_Layout_1.C 0.165f
C198 B a_3328_n363# 8.97e-19
C199 OR_2_In_Layout_0.B AND_2_In_Layout_0.A 0.00473f
C200 a_801_375# VDD 0.79f
C201 S4 a_3184_375# 3.42e-19
C202 S4 a_801_n1645# 0.259f
C203 A a_3184_375# 0.0018f
C204 a_945_n1645# OR_2_In_Layout_0.A 0.203f
C205 A a_801_n1645# 0.299f
C206 OR_2_In_Layout_0.B OR_2_In_Layout_0.A 1.3f
C207 C a_3184_n363# 5.7e-19
C208 S4 a_801_n363# 0.00164f
C209 A a_801_n363# 0.314f
C210 a_3184_n363# a_3808_n363# 0.429f
C211 VDD a_3303_n1718# 0.189f
C212 AND_2_In_Layout_0.A S1 2.75e-19
C213 VDD a_1425_n363# 0.0527f
C214 OR_2_In_Layout_0.B AND_3_In_Layout_1.C 0.00284f
C215 S3 S2 0.00677f
C216 a_1425_375# S5 0.00586f
C217 a_1425_375# a_945_375# 0.248f
C218 S1 AND_3_In_Layout_1.C 0.0853f
C219 S4 OR_2_In_Layout_0.B 0.0626f
C220 a_4292_n1650# a_3184_n363# 0.00209f
C221 A a_945_n1645# 0.0499f
C222 A OR_2_In_Layout_0.B 0.108f
C223 a_3328_n363# a_3184_n363# 0.343f
C224 a_4292_n1650# a_4148_n1650# 0.361f
C225 VDD AND_2_In_Layout_0.A 0.372f
C226 VDD OR_2_In_Layout_0.A 0.933f
C227 A S1 0.00105f
C228 C S6 0.105f
C229 S2 a_3184_375# 0.259f
C230 S5 a_3184_375# 1.14e-20
C231 a_801_n1645# S5 7.66e-19
C232 VDD AND_3_In_Layout_1.C 0.71f
C233 B a_1425_375# 0.0525f
C234 S5 a_801_n363# 0.267f
C235 a_3303_n1718# AND_2_In_Layout_0.A 0.127f
C236 a_801_375# AND_3_In_Layout_1.C 0.0531f
C237 a_3303_n1718# OR_2_In_Layout_0.A 0.0325f
C238 a_1425_n1645# a_801_n1645# 0.429f
C239 a_3808_375# a_3184_375# 0.429f
C240 a_1425_n363# OR_2_In_Layout_0.A 0.0125f
C241 C a_3328_n363# 4.96e-19
C242 a_3328_n363# a_3808_n363# 0.248f
C243 a_4148_n1650# VSS 0.468f
C244 a_1425_n1645# VSS 0.37f
C245 a_945_n1645# VSS 0.248f
C246 S1 VSS 0.33f
C247 a_2999_n1346# VSS 0.102f
C248 a_3303_n1718# VSS 0.563f
C249 a_4292_n1650# VSS 0.383f
C250 AND_2_In_Layout_0.A VSS 0.567f
C251 S4 VSS 0.613f
C252 a_801_n1645# VSS 0.708f
C253 S3 VSS 0.422f
C254 a_3808_n363# VSS 0.316f
C255 a_3328_n363# VSS 0.16f
C256 S5 VSS 0.678f
C257 a_1425_n363# VSS 0.367f
C258 a_945_n363# VSS 0.152f
C259 a_3184_n363# VSS 0.615f
C260 a_801_n363# VSS 0.645f
C261 OR_2_In_Layout_0.B VSS 3.62f
C262 OR_2_In_Layout_0.A VSS 3.9f
C263 a_3808_375# VSS 0.316f
C264 a_3328_375# VSS 0.242f
C265 a_1425_375# VSS 0.318f
C266 a_945_375# VSS 0.16f
C267 S2 VSS 0.509f
C268 S6 VSS 0.554f
C269 a_3184_375# VSS 0.664f
C270 AND_3_In_Layout_1.C VSS 3.72f
C271 a_801_375# VSS 0.622f
C272 C VSS 5.44f
C273 B VSS 4.48f
C274 A VSS 4.66f
C275 VDD VSS 14f
C276 VDD.t70 VSS 0.0024f
C277 VDD.n0 VSS 0.0024f
C278 VDD.n1 VSS 0.00521f
C279 VDD.n2 VSS 0.0174f
C280 VDD.n3 VSS 0.00313f
C281 VDD.t69 VSS 0.0123f
C282 VDD.n4 VSS 0.0296f
C283 VDD.n5 VSS 0.0398f
C284 VDD.t38 VSS 0.0112f
C285 VDD.n6 VSS 0.0129f
C286 VDD.n7 VSS 0.00312f
C287 VDD.n8 VSS 0.00413f
C288 VDD.t50 VSS 0.0024f
C289 VDD.n9 VSS 0.0024f
C290 VDD.n10 VSS 0.00521f
C291 VDD.n11 VSS 0.0246f
C292 VDD.n12 VSS 0.00315f
C293 VDD.n13 VSS 0.00312f
C294 VDD.t20 VSS 0.0118f
C295 VDD.t54 VSS 0.0112f
C296 VDD.n14 VSS 0.00312f
C297 VDD.t21 VSS 0.0024f
C298 VDD.n15 VSS 0.0024f
C299 VDD.n16 VSS 0.00521f
C300 VDD.n17 VSS 0.00754f
C301 VDD.n18 VSS 0.00351f
C302 VDD.n19 VSS 0.00243f
C303 VDD.n20 VSS 0.00204f
C304 VDD.t8 VSS 0.0024f
C305 VDD.n21 VSS 0.0024f
C306 VDD.n22 VSS 0.00521f
C307 VDD.t71 VSS 0.0024f
C308 VDD.n23 VSS 0.0024f
C309 VDD.n24 VSS 0.00521f
C310 VDD.n25 VSS 0.0127f
C311 VDD.n26 VSS 0.00312f
C312 VDD.n27 VSS 0.00312f
C313 VDD.n28 VSS 0.00312f
C314 VDD.n29 VSS 0.00485f
C315 VDD.n30 VSS 0.00312f
C316 VDD.n31 VSS 0.0155f
C317 VDD.n32 VSS 0.00312f
C318 VDD.t63 VSS 0.0024f
C319 VDD.n33 VSS 0.0024f
C320 VDD.n34 VSS 0.00548f
C321 VDD.n35 VSS 0.00364f
C322 VDD.n36 VSS 0.00312f
C323 VDD.t12 VSS 0.0226f
C324 VDD.n37 VSS 0.00334f
C325 VDD.n38 VSS 0.0031f
C326 VDD.n39 VSS 0.00312f
C327 VDD.t64 VSS 0.021f
C328 VDD.n40 VSS 0.00312f
C329 VDD.n41 VSS 0.00641f
C330 VDD.t3 VSS 0.0024f
C331 VDD.n42 VSS 0.0024f
C332 VDD.n43 VSS 0.00521f
C333 VDD.n44 VSS 0.00754f
C334 VDD.n45 VSS 0.00312f
C335 VDD.n46 VSS 0.0324f
C336 VDD.t4 VSS 0.0121f
C337 VDD.t2 VSS 0.027f
C338 VDD.t0 VSS 0.0272f
C339 VDD.n47 VSS 0.0158f
C340 VDD.n48 VSS 0.00312f
C341 VDD.n49 VSS 0.00312f
C342 VDD.t37 VSS 0.0024f
C343 VDD.n50 VSS 0.0024f
C344 VDD.n51 VSS 0.00523f
C345 VDD.n52 VSS 0.0432f
C346 VDD.n53 VSS 0.00313f
C347 VDD.n54 VSS 0.0282f
C348 VDD.t36 VSS 0.0129f
C349 VDD.n55 VSS 0.0193f
C350 VDD.n56 VSS 0.0147f
C351 VDD.t40 VSS 0.0227f
C352 VDD.n57 VSS 0.00312f
C353 VDD.n58 VSS 0.00485f
C354 VDD.t1 VSS 0.00619f
C355 VDD.n59 VSS 0.00315f
C356 VDD.n60 VSS 0.00351f
C357 VDD.n61 VSS 0.00999f
C358 VDD.n62 VSS 0.00377f
C359 VDD.n63 VSS 0.00312f
C360 VDD.n65 VSS 0.0212f
C361 VDD.n66 VSS 0.0369f
C362 VDD.n67 VSS 0.0104f
C363 VDD.n68 VSS 0.00312f
C364 VDD.n69 VSS 0.00413f
C365 VDD.n70 VSS 0.0112f
C366 VDD.t65 VSS 0.0024f
C367 VDD.n71 VSS 0.0024f
C368 VDD.n72 VSS 0.00521f
C369 VDD.n73 VSS 0.00757f
C370 VDD.n74 VSS 0.00271f
C371 VDD.n75 VSS 0.00312f
C372 VDD.n76 VSS 0.0128f
C373 VDD.t22 VSS 0.021f
C374 VDD.n77 VSS 0.023f
C375 VDD.t14 VSS 0.021f
C376 VDD.n78 VSS 0.032f
C377 VDD.n79 VSS 0.0304f
C378 VDD.n80 VSS 0.00312f
C379 VDD.n81 VSS 0.00485f
C380 VDD.n82 VSS 0.00519f
C381 VDD.n83 VSS 0.00397f
C382 VDD.n84 VSS 0.00334f
C383 VDD.n85 VSS 0.02f
C384 VDD.n86 VSS 0.0139f
C385 VDD.t13 VSS 0.0128f
C386 VDD.t62 VSS 0.0128f
C387 VDD.n87 VSS 0.0218f
C388 VDD.n88 VSS 0.00312f
C389 VDD.n89 VSS 0.00485f
C390 VDD.n90 VSS 0.00397f
C391 VDD.n91 VSS 0.00882f
C392 VDD.n92 VSS 0.0033f
C393 VDD.n93 VSS 0.00312f
C394 VDD.n94 VSS 0.0191f
C395 VDD.t58 VSS 0.0135f
C396 VDD.n95 VSS 0.0283f
C397 VDD.n96 VSS 0.0494f
C398 VDD.n97 VSS 0.00315f
C399 VDD.n98 VSS 0.00485f
C400 VDD.n99 VSS 0.061f
C401 VDD.n100 VSS 0.0421f
C402 VDD.t7 VSS 0.0211f
C403 VDD.n101 VSS 0.0302f
C404 VDD.n102 VSS 0.0302f
C405 VDD.n103 VSS 0.00314f
C406 VDD.t57 VSS 0.0024f
C407 VDD.n104 VSS 0.0024f
C408 VDD.n105 VSS 0.00521f
C409 VDD.t61 VSS 0.0024f
C410 VDD.n106 VSS 0.0024f
C411 VDD.n107 VSS 0.00521f
C412 VDD.t9 VSS 0.0226f
C413 VDD.n108 VSS 0.047f
C414 VDD.n109 VSS 0.057f
C415 VDD.n110 VSS 0.00392f
C416 VDD.n111 VSS 0.00312f
C417 VDD.n112 VSS 0.0224f
C418 VDD.t56 VSS 0.0195f
C419 VDD.n113 VSS 0.0331f
C420 VDD.t17 VSS 0.0195f
C421 VDD.n114 VSS 0.0224f
C422 VDD.n115 VSS 0.00312f
C423 VDD.n116 VSS 0.00388f
C424 VDD.n117 VSS 0.00206f
C425 VDD.n118 VSS 0.0035f
C426 VDD.n119 VSS 0.0517f
C427 VDD.n120 VSS 0.0513f
C428 VDD.t55 VSS 0.0024f
C429 VDD.n121 VSS 0.0024f
C430 VDD.n122 VSS 0.00521f
C431 VDD.n123 VSS 0.00485f
C432 VDD.n124 VSS 0.00312f
C433 VDD.n125 VSS 0.0129f
C434 VDD.n126 VSS 0.00176f
C435 VDD.n127 VSS 0.00626f
C436 VDD.t66 VSS 0.0658f
C437 VDD.n128 VSS 0.0358f
C438 VDD.n129 VSS 0.00176f
C439 VDD.n130 VSS 0.00364f
C440 VDD.n131 VSS 0.00312f
C441 VDD.t51 VSS 0.0658f
C442 VDD.t31 VSS 0.0658f
C443 VDD.n132 VSS 0.00312f
C444 VDD.n133 VSS 0.00626f
C445 VDD.n134 VSS 0.00626f
C446 VDD.n135 VSS 0.00206f
C447 VDD.n136 VSS 0.024f
C448 VDD.n137 VSS 0.00181f
C449 VDD.n138 VSS 0.046f
C450 VDD.n139 VSS 0.00176f
C451 VDD.n140 VSS 0.0579f
C452 VDD.n141 VSS 0.0579f
C453 VDD.n142 VSS 0.00364f
C454 VDD.n143 VSS 0.00312f
C455 VDD.n144 VSS 0.00312f
C456 VDD.n145 VSS 0.00206f
C457 VDD.n146 VSS 0.0104f
C458 VDD.n147 VSS 0.0223f
C459 VDD.n148 VSS 0.043f
C460 VDD.n149 VSS 0.0246f
C461 VDD.t44 VSS 0.0118f
C462 VDD.n150 VSS 0.0174f
C463 VDD.n151 VSS 0.00312f
C464 VDD.n152 VSS 0.0031f
C465 VDD.n153 VSS 0.00757f
C466 VDD.n154 VSS 0.00354f
C467 VDD.n155 VSS 0.00353f
C468 VDD.n156 VSS 0.00243f
C469 VDD.n157 VSS 0.00312f
C470 VDD.n158 VSS 0.0191f
C471 VDD.t25 VSS 0.0112f
C472 VDD.n159 VSS 0.0129f
C473 VDD.n160 VSS 0.0174f
C474 VDD.n161 VSS 0.00312f
C475 VDD.n162 VSS 0.00312f
C476 VDD.n163 VSS 0.00485f
C477 VDD.n164 VSS 0.0541f
C478 VDD.n165 VSS 0.0345f
C479 VDD.t28 VSS 0.0118f
C480 VDD.n166 VSS 0.0246f
C481 VDD.n167 VSS 0.00312f
C482 VDD.n168 VSS 0.00485f
C483 VDD.n169 VSS 0.0174f
C484 VDD.n170 VSS 0.00312f
C485 VDD.n171 VSS 0.0031f
C486 VDD.n172 VSS 0.00757f
C487 VDD.t49 VSS 0.0112f
C488 VDD.n173 VSS 0.0129f
C489 VDD.n174 VSS 0.00312f
C490 VDD.n175 VSS 0.00418f
C491 VDD.n176 VSS 0.0191f
C492 VDD.n177 VSS 0.00312f
C493 C.t8 VSS 0.00777f
C494 C.t0 VSS 0.0266f
C495 C.n0 VSS 0.0535f
C496 C.t9 VSS 0.0465f
C497 C.t6 VSS 0.0422f
C498 C.n1 VSS 0.0707f
C499 C.n2 VSS 0.296f
C500 C.t3 VSS 0.00777f
C501 C.t13 VSS 0.00777f
C502 C.t10 VSS 0.065f
C503 C.t11 VSS 0.0815f
C504 C.n3 VSS 0.0452f
C505 C.n4 VSS 0.0601f
C506 C.n5 VSS 0.185f
C507 C.t2 VSS 0.0358f
C508 C.t7 VSS 0.0106f
C509 C.n6 VSS 0.0533f
C510 C.n7 VSS 0.261f
C511 C.n8 VSS 0.499f
C512 C.t5 VSS 0.00777f
C513 C.t12 VSS 0.00777f
C514 C.t1 VSS 0.065f
C515 C.t4 VSS 0.0815f
C516 C.n9 VSS 0.0452f
C517 C.n10 VSS 0.0601f
.ends

