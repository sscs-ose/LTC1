magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2186 -2045 2186 2045
<< psubdiff >>
rect -186 23 186 45
rect -186 -23 -164 23
rect 164 -23 186 23
rect -186 -45 186 -23
<< psubdiffcont >>
rect -164 -23 164 23
<< metal1 >>
rect -175 23 175 34
rect -175 -23 -164 23
rect 164 -23 175 23
rect -175 -34 175 -23
<< end >>
