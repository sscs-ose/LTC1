magic
tech gf180mcuC
magscale 1 10
timestamp 1691493578
<< nwell >>
rect -522 -230 522 230
<< pmos >>
rect -348 -100 -292 100
rect -188 -100 -132 100
rect -28 -100 28 100
rect 132 -100 188 100
rect 292 -100 348 100
<< pdiff >>
rect -436 87 -348 100
rect -436 -87 -423 87
rect -377 -87 -348 87
rect -436 -100 -348 -87
rect -292 87 -188 100
rect -292 -87 -263 87
rect -217 -87 -188 87
rect -292 -100 -188 -87
rect -132 87 -28 100
rect -132 -87 -103 87
rect -57 -87 -28 87
rect -132 -100 -28 -87
rect 28 87 132 100
rect 28 -87 57 87
rect 103 -87 132 87
rect 28 -100 132 -87
rect 188 87 292 100
rect 188 -87 217 87
rect 263 -87 292 87
rect 188 -100 292 -87
rect 348 87 436 100
rect 348 -87 377 87
rect 423 -87 436 87
rect 348 -100 436 -87
<< pdiffc >>
rect -423 -87 -377 87
rect -263 -87 -217 87
rect -103 -87 -57 87
rect 57 -87 103 87
rect 217 -87 263 87
rect 377 -87 423 87
<< polysilicon >>
rect -348 100 -292 144
rect -188 100 -132 144
rect -28 100 28 144
rect 132 100 188 144
rect 292 100 348 144
rect -348 -144 -292 -100
rect -188 -144 -132 -100
rect -28 -144 28 -100
rect 132 -144 188 -100
rect 292 -144 348 -100
<< metal1 >>
rect -423 87 -377 98
rect -423 -98 -377 -87
rect -263 87 -217 98
rect -263 -98 -217 -87
rect -103 87 -57 98
rect -103 -98 -57 -87
rect 57 87 103 98
rect 57 -98 103 -87
rect 217 87 263 98
rect 217 -98 263 -87
rect 377 87 423 98
rect 377 -98 423 -87
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 1 l 0.280 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
