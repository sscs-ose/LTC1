magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2000 -2000 14876 23798
<< metal1 >>
rect 124 3386 12876 3586
rect 0 106 6716 306
rect 6892 106 12876 306
<< metal2 >>
rect 0 0 1102 20299
rect 1438 0 3266 16554
rect 3366 0 5194 21210
rect 5294 0 6388 21798
rect 6488 0 7582 17815
rect 7682 0 9510 19430
rect 9610 0 11438 17818
rect 11774 0 12876 19431
use M2_M1_CDNS_69033583165352  M2_M1_CDNS_69033583165352_0
timestamp 1713338890
transform 1 0 5841 0 1 206
box -524 -92 524 92
use M2_M1_CDNS_69033583165352  M2_M1_CDNS_69033583165352_1
timestamp 1713338890
transform 1 0 7035 0 1 3486
box -524 -92 524 92
use M2_M1_CDNS_69033583165352  M2_M1_CDNS_69033583165352_2
timestamp 1713338890
transform 1 0 12325 0 1 206
box -524 -92 524 92
use M2_M1_CDNS_69033583165352  M2_M1_CDNS_69033583165352_3
timestamp 1713338890
transform 1 0 5841 0 1 3954
box -524 -92 524 92
use M2_M1_CDNS_69033583165352  M2_M1_CDNS_69033583165352_4
timestamp 1713338890
transform 1 0 5841 0 1 16038
box -524 -92 524 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_0
timestamp 1713338890
transform 1 0 2352 0 1 206
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_1
timestamp 1713338890
transform 1 0 4280 0 1 3486
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_2
timestamp 1713338890
transform 1 0 10524 0 1 3486
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_3
timestamp 1713338890
transform 1 0 2352 0 1 3954
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_4
timestamp 1713338890
transform 1 0 8596 0 1 3954
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_5
timestamp 1713338890
transform 1 0 2352 0 1 16038
box -902 -92 902 92
use M2_M1_CDNS_69033583165353  M2_M1_CDNS_69033583165353_6
timestamp 1713338890
transform 1 0 8596 0 1 16038
box -902 -92 902 92
use M2_M1_CDNS_69033583165365  M2_M1_CDNS_69033583165365_0
timestamp 1713338890
transform 1 0 8686 0 1 206
box -794 -92 794 92
use M2_M1_CDNS_69033583165366  M2_M1_CDNS_69033583165366_0
timestamp 1713338890
transform 1 0 5841 0 1 10045
box -534 -348 534 348
use M2_M1_CDNS_69033583165367  M2_M1_CDNS_69033583165367_0
timestamp 1713338890
transform 1 0 2352 0 1 10045
box -906 -348 906 348
use M2_M1_CDNS_69033583165367  M2_M1_CDNS_69033583165367_1
timestamp 1713338890
transform 1 0 8596 0 1 10045
box -906 -348 906 348
use M2_M1_CDNS_69033583165368  M2_M1_CDNS_69033583165368_0
timestamp 1713338890
transform 1 0 608 0 1 3486
box -470 -92 470 92
use M2_M1_CDNS_69033583165369  M2_M1_CDNS_69033583165369_0
timestamp 1713338890
transform 1 0 607 0 1 16529
box -416 -38 416 38
<< end >>
