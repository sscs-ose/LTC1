magic
tech gf180mcuC
magscale 1 10
timestamp 1691568605
<< nwell >>
rect -296 -330 296 330
<< pmos >>
rect -122 -200 -52 200
rect 52 -200 122 200
<< pdiff >>
rect -210 187 -122 200
rect -210 -187 -197 187
rect -151 -187 -122 187
rect -210 -200 -122 -187
rect -52 187 52 200
rect -52 -187 -23 187
rect 23 -187 52 187
rect -52 -200 52 -187
rect 122 187 210 200
rect 122 -187 151 187
rect 197 -187 210 187
rect 122 -200 210 -187
<< pdiffc >>
rect -197 -187 -151 187
rect -23 -187 23 187
rect 151 -187 197 187
<< polysilicon >>
rect -122 200 -52 244
rect 52 200 122 244
rect -122 -244 -52 -200
rect 52 -244 122 -200
<< metal1 >>
rect -197 187 -151 198
rect -197 -198 -151 -187
rect -23 187 23 198
rect -23 -198 23 -187
rect 151 187 197 198
rect 151 -198 197 -187
<< properties >>
string gencell pmos_3p3
string library gf180mcu
string parameters w 2 l 0.35 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {pmos_3p3 pmos_6p0}
<< end >>
