** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/GF_INV_PEX_TB.sym
**.subckt GF_INV_PEX_TB
C1 OUT VSS 50f m=1
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
V3 IN VSS pulse(0 3.3 0 100p 100p 100n 200n)
.save i(v3)
x1 VSS VDD OUT IN GF_INV_PEX
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_GF_INV_MAG.spice
.control
save all
dc v3 0 3.3 0.1
plot v(IN) v(OUT)

tran 10p 1u
plot v(IN) v(OUT)
*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
