magic
tech gf180mcuD
magscale 1 10
timestamp 1713971633
<< checkpaint >>
rect -4075 -2823 7510 3762
<< nwell >>
rect 1083 1624 2885 1631
rect 126 1530 1112 1538
rect 1990 1069 2885 1624
rect 1990 1043 2353 1069
rect 2606 1043 2885 1069
rect 1083 -739 1128 -159
rect 2199 -177 2400 -151
rect 2199 -642 2352 -177
rect 2107 -715 2444 -642
rect 2199 -739 2352 -715
<< pwell >>
rect -1173 649 -919 1009
rect 1021 971 2353 1016
rect 2606 984 5127 1016
rect 2714 983 5127 984
rect 2606 971 5127 983
rect 1021 647 5127 971
rect 1136 -87 4626 236
rect 1136 -96 4296 -87
rect 4350 -96 4626 -87
rect 1136 -116 4626 -96
<< psubdiff >>
rect -959 538 -801 556
rect -959 492 -906 538
rect -860 492 -801 538
rect -959 475 -801 492
<< nsubdiff >>
rect 2107 -655 2444 -642
rect 2107 -701 2232 -655
rect 2278 -701 2444 -655
rect 2107 -715 2444 -701
<< psubdiffcont >>
rect -906 492 -860 538
<< nsubdiffcont >>
rect 2232 -701 2278 -655
<< metal1 >>
rect -1048 1750 -971 1762
rect -1048 1731 -1036 1750
rect -2075 1698 -1036 1731
rect -984 1731 -971 1750
rect -853 1750 -776 1762
rect -853 1731 -841 1750
rect -984 1698 -841 1731
rect -789 1731 -776 1750
rect 5427 1736 5505 1752
rect 5427 1731 5440 1736
rect -789 1698 5440 1731
rect -2075 1685 5440 1698
rect -2075 1035 -2029 1685
rect 5421 1684 5440 1685
rect 5492 1684 5505 1736
rect 5421 1670 5505 1684
rect 126 1622 2087 1624
rect -1940 1566 2087 1622
rect -1940 1514 -1902 1566
rect -1850 1538 2087 1566
rect -1850 1514 126 1538
rect 1112 1530 2087 1538
rect 2375 1584 5357 1630
rect 2375 1583 5287 1584
rect 2375 1579 5087 1583
rect 2375 1534 4393 1579
rect 4392 1527 4393 1534
rect 4445 1578 5087 1579
rect 4445 1534 4585 1578
rect 4445 1527 4446 1534
rect 4392 1524 4446 1527
rect 4584 1526 4585 1534
rect 4637 1534 5087 1578
rect 4637 1526 4638 1534
rect 5086 1531 5087 1534
rect 5139 1534 5287 1583
rect 5139 1531 5140 1534
rect 5086 1528 5140 1531
rect 5273 1532 5287 1534
rect 5339 1534 5357 1584
rect 5421 1587 5467 1670
rect 5421 1571 5507 1587
rect 5339 1532 5352 1534
rect 4584 1523 4638 1526
rect 5273 1523 5352 1532
rect -1940 1504 126 1514
rect 5421 1519 5442 1571
rect 5494 1519 5507 1571
rect 5421 1504 5507 1519
rect -1911 1503 -1213 1504
rect -958 1503 -812 1504
rect 5421 1479 5467 1504
rect -1140 1081 -1084 1128
rect -1140 1042 -1050 1081
rect -2075 989 -1738 1035
rect -1140 990 -1117 1042
rect -1065 990 -1050 1042
rect -1140 984 -1050 990
rect -837 1048 -760 1060
rect -837 996 -825 1048
rect -773 1036 -760 1048
rect -773 996 -566 1036
rect -837 989 -566 996
rect 1082 1035 1127 1055
rect 1906 1049 1953 1128
rect 5197 1089 5510 1135
rect 1082 989 1364 1035
rect 1906 1002 2219 1049
rect -837 983 -760 989
rect 1157 771 1213 989
rect 1145 755 1227 771
rect 1145 703 1160 755
rect 1212 703 1227 755
rect 1145 688 1227 703
rect 86 620 168 666
rect 2172 660 2219 1002
rect 2288 1043 2511 1053
rect 2288 1039 2539 1043
rect 2288 987 2302 1039
rect 2354 987 2412 1039
rect 2464 1034 2539 1039
rect 4291 1042 4343 1055
rect 4291 1041 4558 1042
rect 2606 1034 2763 1035
rect 2464 988 2763 1034
rect 4291 1003 4580 1041
rect 2464 987 2539 988
rect 2288 983 2539 987
rect 2606 984 2763 988
rect 2714 983 2763 984
rect 2288 973 2511 983
rect 2711 945 2763 983
rect 4294 996 4580 1003
rect 3294 673 3416 690
rect 2156 647 2235 660
rect 2156 595 2169 647
rect 2221 595 2235 647
rect 3294 621 3312 673
rect 3364 666 3416 673
rect 3364 621 3551 666
rect 3294 609 3551 621
rect 3294 603 3416 609
rect 2156 583 2235 595
rect -936 538 -816 556
rect -936 492 -906 538
rect -860 492 -816 538
rect -936 475 -816 492
rect 1033 475 1153 556
rect 2004 542 2081 554
rect 1999 540 2081 542
rect 1999 488 2002 540
rect 2054 488 2081 540
rect 1999 486 2081 488
rect -985 409 -907 424
rect -985 357 -972 409
rect -920 357 -907 409
rect -985 342 -907 357
rect -965 -116 -919 342
rect 1034 337 1163 410
rect 2004 331 2081 486
rect -5 269 85 287
rect -5 217 15 269
rect 67 217 85 269
rect -5 198 85 217
rect 935 72 1011 86
rect 935 20 947 72
rect 999 71 1011 72
rect 999 25 1332 71
rect 999 20 1011 25
rect 935 8 1011 20
rect 855 -90 942 -77
rect -965 -162 -887 -116
rect 855 -142 873 -90
rect 925 -142 942 -90
rect 855 -154 942 -142
rect 1286 -240 1332 25
rect 2172 -104 2219 583
rect 4067 551 4153 553
rect 4051 543 4153 551
rect 2542 535 2600 536
rect 2410 532 2468 533
rect 2410 480 2413 532
rect 2465 480 2468 532
rect 2542 483 2545 535
rect 2597 483 2600 535
rect 2542 482 2600 483
rect 3046 533 3104 534
rect 3046 481 3049 533
rect 3101 481 3104 533
rect 3046 480 3104 481
rect 2410 479 2468 480
rect 3232 375 3300 531
rect 4051 491 4083 543
rect 4135 491 4153 543
rect 4051 481 4153 491
rect 4051 379 4125 481
rect 2292 263 2381 272
rect 2292 211 2309 263
rect 2361 211 2381 263
rect 2292 210 2381 211
rect 2294 208 2381 210
rect 3194 268 3280 281
rect 4294 278 4343 996
rect 4390 543 4471 559
rect 4606 549 5094 563
rect 4606 546 5017 549
rect 4390 491 4404 543
rect 4456 540 4471 543
rect 4585 542 5017 546
rect 4456 491 4534 540
rect 4390 474 4534 491
rect 4585 490 4587 542
rect 4639 497 5017 542
rect 5069 497 5094 549
rect 4639 490 5094 497
rect 4585 486 5094 490
rect 4606 482 5094 486
rect 4453 329 4534 474
rect 4658 329 4739 482
rect 5235 340 5302 543
rect 3194 216 3211 268
rect 3263 216 3280 268
rect 1888 -150 2219 -104
rect 2302 -163 2369 208
rect 3194 204 3280 216
rect 4266 266 4350 278
rect 4266 214 4282 266
rect 4334 214 4350 266
rect 4266 202 4350 214
rect 4174 82 4256 96
rect 4174 30 4189 82
rect 4241 80 4256 82
rect 4241 34 4506 80
rect 4241 30 4256 34
rect 4174 18 4256 30
rect 4287 -96 4365 -85
rect 4119 -97 4365 -96
rect 4119 -142 4300 -97
rect 4287 -149 4300 -142
rect 4352 -149 4365 -97
rect 4287 -161 4365 -149
rect 4460 -197 4506 34
rect 5464 -105 5510 1089
rect 5195 -107 5510 -105
rect 5127 -151 5510 -107
rect 4460 -243 4574 -197
rect -720 -684 -631 -679
rect -720 -736 -701 -684
rect -649 -736 -631 -684
rect 975 -692 1312 -641
rect 2107 -655 2444 -642
rect 2107 -701 2232 -655
rect 2278 -701 2444 -655
rect 4187 -687 4453 -617
rect 5174 -633 5229 -632
rect 5174 -685 5175 -633
rect 5227 -685 5229 -633
rect 5174 -686 5229 -685
rect 5292 -633 5347 -632
rect 5292 -685 5293 -633
rect 5345 -685 5347 -633
rect 5292 -686 5347 -685
rect 2107 -721 2444 -701
rect -720 -757 -631 -736
<< via1 >>
rect -1036 1698 -984 1750
rect -841 1698 -789 1750
rect 5440 1684 5492 1736
rect -1902 1514 -1850 1566
rect 4393 1527 4445 1579
rect 4585 1526 4637 1578
rect 5087 1531 5139 1583
rect 5287 1532 5339 1584
rect 5442 1519 5494 1571
rect -1117 990 -1065 1042
rect -825 996 -773 1048
rect 1160 703 1212 755
rect 2302 987 2354 1039
rect 2412 987 2464 1039
rect 2169 595 2221 647
rect 3312 621 3364 673
rect 2002 488 2054 540
rect -972 357 -920 409
rect 15 217 67 269
rect 947 20 999 72
rect 873 -142 925 -90
rect 2413 480 2465 532
rect 2545 483 2597 535
rect 3049 481 3101 533
rect 4083 491 4135 543
rect 2309 211 2361 263
rect 4404 491 4456 543
rect 4587 490 4639 542
rect 5017 497 5069 549
rect 3211 216 3263 268
rect 4282 214 4334 266
rect 4189 30 4241 82
rect 4300 -149 4352 -97
rect -701 -736 -649 -684
rect 5175 -685 5227 -633
rect 5293 -685 5345 -633
<< metal2 >>
rect -1048 1755 -971 1762
rect -853 1755 -776 1762
rect -1055 1750 -776 1755
rect -1055 1698 -1036 1750
rect -984 1698 -841 1750
rect -789 1698 -776 1750
rect -1055 1695 -776 1698
rect -2014 1566 -1833 1580
rect -2014 1514 -1902 1566
rect -1850 1514 -1833 1566
rect -2014 1500 -1833 1514
rect -1758 1576 -1658 1580
rect -1566 1576 -1503 1582
rect -1273 1579 -1210 1588
rect -1338 1577 -1210 1579
rect -2014 -756 -1845 1500
rect -1758 -756 -1503 1576
rect -1400 -756 -1210 1577
rect -1055 1446 -995 1695
rect -853 1693 -776 1695
rect 5427 1736 5505 1752
rect 5427 1684 5440 1736
rect 5492 1684 5505 1736
rect 5427 1670 5505 1684
rect 5273 1589 5357 1607
rect 4375 1584 5357 1589
rect 5440 1587 5496 1670
rect 4375 1583 5287 1584
rect 4375 1579 5087 1583
rect 4375 1527 4393 1579
rect 4445 1578 5087 1579
rect 4445 1527 4585 1578
rect 4375 1526 4585 1527
rect 4637 1531 5087 1578
rect 5139 1532 5287 1583
rect 5339 1532 5357 1584
rect 5139 1531 5357 1532
rect 4637 1526 5357 1531
rect 4375 1523 5357 1526
rect 5431 1571 5507 1587
rect 4375 1520 4704 1523
rect -1055 1386 -772 1446
rect -832 1060 -772 1386
rect -1140 1042 -1050 1055
rect -1140 990 -1117 1042
rect -1065 990 -1050 1042
rect -1140 984 -1050 990
rect -837 1050 -760 1060
rect -837 1048 -587 1050
rect -837 996 -825 1048
rect -773 996 -587 1048
rect 2288 1043 2511 1053
rect 2288 1042 2539 1043
rect -837 990 -587 996
rect 910 1039 2539 1042
rect -1121 811 -1062 984
rect -837 983 -760 990
rect 910 987 2302 1039
rect 2354 987 2412 1039
rect 2464 987 2539 1039
rect 910 983 2539 987
rect 910 811 969 983
rect 2288 973 2511 983
rect -1121 752 969 811
rect 1145 755 1227 771
rect -1121 -495 -1062 752
rect 1145 703 1160 755
rect 1212 703 1227 755
rect 1145 688 1227 703
rect 1145 635 1209 688
rect 3294 673 3416 690
rect 3294 670 3312 673
rect 2200 660 3312 670
rect 1095 577 1209 635
rect 2156 647 3312 660
rect 2156 595 2169 647
rect 2221 621 3312 647
rect 3364 670 3416 673
rect 3364 621 3491 670
rect 2221 596 3491 621
rect 2221 595 2235 596
rect 2156 583 2235 595
rect -985 418 -907 424
rect 1095 418 1153 577
rect 1987 540 2072 556
rect 4390 553 5100 559
rect 1987 488 2002 540
rect 2054 517 2072 540
rect 4067 549 5100 553
rect 4067 543 5017 549
rect 2383 535 3150 539
rect 2383 532 2545 535
rect 2383 517 2413 532
rect 2054 488 2413 517
rect 1987 480 2413 488
rect 2465 483 2545 532
rect 2597 533 3150 535
rect 2597 483 3049 533
rect 2465 481 3049 483
rect 3101 481 3150 533
rect 4067 491 4083 543
rect 4135 491 4404 543
rect 4456 542 5017 543
rect 4456 491 4587 542
rect 4067 490 4587 491
rect 4639 497 5017 542
rect 5069 497 5100 549
rect 4639 490 5100 497
rect 4067 483 5100 490
rect 4067 481 4153 483
rect 2465 480 3150 481
rect 1987 475 3150 480
rect 1987 473 2481 475
rect 4390 474 4471 483
rect 2000 460 2481 473
rect 2000 459 2244 460
rect 2000 445 2058 459
rect -985 409 1157 418
rect -985 357 -972 409
rect -920 360 1157 409
rect -920 357 -907 360
rect -985 342 -907 357
rect 2300 337 4344 404
rect -5 271 85 287
rect 2300 272 2367 337
rect 3194 274 3280 281
rect 4277 278 4344 337
rect -17 269 266 271
rect -17 217 15 269
rect 67 217 266 269
rect -17 207 266 217
rect 2292 263 2381 272
rect 2292 211 2309 263
rect 2361 211 2381 263
rect 2292 210 2381 211
rect 2294 208 2381 210
rect 3194 268 3580 274
rect 3194 216 3211 268
rect 3263 216 3580 268
rect 3194 211 3580 216
rect -5 198 85 207
rect 202 79 266 207
rect 3194 204 3280 211
rect 3517 91 3580 211
rect 4266 266 4350 278
rect 4266 214 4282 266
rect 4334 214 4350 266
rect 4266 202 4350 214
rect 4174 91 4256 96
rect 935 79 1011 86
rect 202 72 1011 79
rect 202 20 947 72
rect 999 20 1011 72
rect 3517 82 4256 91
rect 3517 30 4189 82
rect 4241 30 4256 82
rect 3517 28 4256 30
rect 4125 26 4256 28
rect 202 15 1011 20
rect 4174 18 4256 26
rect 935 8 1011 15
rect 886 -77 945 -71
rect 855 -90 945 -77
rect 4287 -88 4365 -85
rect 855 -142 873 -90
rect 925 -142 945 -90
rect 855 -154 945 -142
rect 4261 -97 4408 -88
rect 4261 -144 4300 -97
rect 886 -388 945 -154
rect 4287 -149 4300 -144
rect 4352 -149 4408 -97
rect 4287 -161 4408 -149
rect 886 -495 949 -388
rect -1121 -554 949 -495
rect -720 -684 -631 -679
rect -720 -736 -701 -684
rect -649 -736 -631 -684
rect -720 -756 -631 -736
rect -2014 -819 -631 -756
rect 4352 -767 4408 -161
rect 5290 -619 5356 1523
rect 5431 1519 5442 1571
rect 5494 1519 5507 1571
rect 5431 1504 5507 1519
rect 5280 -625 5360 -619
rect 5162 -633 5360 -625
rect 5162 -685 5175 -633
rect 5227 -685 5293 -633
rect 5345 -685 5360 -633
rect 5162 -691 5360 -685
rect 5280 -698 5360 -691
rect 5440 -767 5496 1504
rect 4352 -823 5496 -767
use inverter_magic  inverter_magic_2
timestamp 1713185578
transform 1 0 4297 0 1 1051
box 0 -569 1108 580
use inverter_magic  inverter_magic_3
timestamp 1713185578
transform -1 0 5456 0 -1 -159
box 0 -569 1108 580
use inverter_magic  inverter_magic_4
timestamp 1713185578
transform -1 0 2199 0 -1 -159
box 0 -569 1108 580
use inverter_magic  inverter_magic_5
timestamp 1713185578
transform 1 0 -2001 0 1 1044
box 0 -569 1108 580
use inverter_magic  inverter_magic_6
timestamp 1713185578
transform 1 0 1034 0 1 1044
box 0 -569 1108 580
use tg_magic  tg_magic_0
timestamp 1713185578
transform -1 0 1134 0 -1 378
box -2 -52 2031 1117
use tg_magic  tg_magic_1
timestamp 1713185578
transform 1 0 2297 0 1 514
box -2 -52 2031 1117
use tg_magic  tg_magic_2
timestamp 1713185578
transform -1 0 4348 0 -1 378
box -2 -52 2031 1117
use tg_magic  tg_magic_3
timestamp 1713185578
transform 1 0 -917 0 1 515
box -2 -52 2031 1117
<< labels >>
flabel psubdiffcont -883 516 -883 516 0 FreeSans 750 0 0 0 VSS
flabel nsubdiffcont 2255 -678 2255 -678 0 FreeSans 750 0 0 0 VDD
flabel metal1 s -1848 1012 -1848 1012 0 FreeSans 750 0 0 0 CLK
port 1 nsew
flabel metal1 s 106 642 106 642 0 FreeSans 750 0 0 0 D
port 2 nsew
flabel metal1 s 5488 450 5488 450 0 FreeSans 750 0 0 0 Q
port 3 nsew
<< end >>
