magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1127 -1019 1127 1019
<< metal1 >>
rect -127 13 127 19
rect -127 -13 -121 13
rect -95 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 95 13
rect 121 -13 127 13
rect -127 -19 127 -13
<< via1 >>
rect -121 -13 -95 13
rect -67 -13 -41 13
rect -13 -13 13 13
rect 41 -13 67 13
rect 95 -13 121 13
<< metal2 >>
rect -127 13 127 19
rect -127 -13 -121 13
rect -95 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 95 13
rect 121 -13 127 13
rect -127 -19 127 -13
<< end >>
