magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1073 -1127 1073 1127
<< metal1 >>
rect -73 121 73 127
rect -73 95 -67 121
rect -41 95 -13 121
rect 13 95 41 121
rect 67 95 73 121
rect -73 67 73 95
rect -73 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 73 67
rect -73 13 73 41
rect -73 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 73 13
rect -73 -41 73 -13
rect -73 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 73 -41
rect -73 -95 73 -67
rect -73 -121 -67 -95
rect -41 -121 -13 -95
rect 13 -121 41 -95
rect 67 -121 73 -95
rect -73 -127 73 -121
<< via1 >>
rect -67 95 -41 121
rect -13 95 13 121
rect 41 95 67 121
rect -67 41 -41 67
rect -13 41 13 67
rect 41 41 67 67
rect -67 -13 -41 13
rect -13 -13 13 13
rect 41 -13 67 13
rect -67 -67 -41 -41
rect -13 -67 13 -41
rect 41 -67 67 -41
rect -67 -121 -41 -95
rect -13 -121 13 -95
rect 41 -121 67 -95
<< metal2 >>
rect -73 121 73 127
rect -73 95 -67 121
rect -41 95 -13 121
rect 13 95 41 121
rect 67 95 73 121
rect -73 67 73 95
rect -73 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 73 67
rect -73 13 73 41
rect -73 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 73 13
rect -73 -41 73 -13
rect -73 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 73 -41
rect -73 -95 73 -67
rect -73 -121 -67 -95
rect -41 -121 -13 -95
rect 13 -121 41 -95
rect 67 -121 73 -95
rect -73 -127 73 -121
<< end >>
