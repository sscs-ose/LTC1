magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1208 -1704 1208 1704
<< metal4 >>
rect -205 696 205 701
rect -205 668 -200 696
rect -172 668 -138 696
rect -110 668 -76 696
rect -48 668 -14 696
rect 14 668 48 696
rect 76 668 110 696
rect 138 668 172 696
rect 200 668 205 696
rect -205 634 205 668
rect -205 606 -200 634
rect -172 606 -138 634
rect -110 606 -76 634
rect -48 606 -14 634
rect 14 606 48 634
rect 76 606 110 634
rect 138 606 172 634
rect 200 606 205 634
rect -205 572 205 606
rect -205 544 -200 572
rect -172 544 -138 572
rect -110 544 -76 572
rect -48 544 -14 572
rect 14 544 48 572
rect 76 544 110 572
rect 138 544 172 572
rect 200 544 205 572
rect -205 510 205 544
rect -205 482 -200 510
rect -172 482 -138 510
rect -110 482 -76 510
rect -48 482 -14 510
rect 14 482 48 510
rect 76 482 110 510
rect 138 482 172 510
rect 200 482 205 510
rect -205 448 205 482
rect -205 420 -200 448
rect -172 420 -138 448
rect -110 420 -76 448
rect -48 420 -14 448
rect 14 420 48 448
rect 76 420 110 448
rect 138 420 172 448
rect 200 420 205 448
rect -205 386 205 420
rect -205 358 -200 386
rect -172 358 -138 386
rect -110 358 -76 386
rect -48 358 -14 386
rect 14 358 48 386
rect 76 358 110 386
rect 138 358 172 386
rect 200 358 205 386
rect -205 324 205 358
rect -205 296 -200 324
rect -172 296 -138 324
rect -110 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 110 324
rect 138 296 172 324
rect 200 296 205 324
rect -205 262 205 296
rect -205 234 -200 262
rect -172 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 172 262
rect 200 234 205 262
rect -205 200 205 234
rect -205 172 -200 200
rect -172 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 172 200
rect 200 172 205 200
rect -205 138 205 172
rect -205 110 -200 138
rect -172 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 172 138
rect 200 110 205 138
rect -205 76 205 110
rect -205 48 -200 76
rect -172 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 172 76
rect 200 48 205 76
rect -205 14 205 48
rect -205 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 205 14
rect -205 -48 205 -14
rect -205 -76 -200 -48
rect -172 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 172 -48
rect 200 -76 205 -48
rect -205 -110 205 -76
rect -205 -138 -200 -110
rect -172 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 172 -110
rect 200 -138 205 -110
rect -205 -172 205 -138
rect -205 -200 -200 -172
rect -172 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 172 -172
rect 200 -200 205 -172
rect -205 -234 205 -200
rect -205 -262 -200 -234
rect -172 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 172 -234
rect 200 -262 205 -234
rect -205 -296 205 -262
rect -205 -324 -200 -296
rect -172 -324 -138 -296
rect -110 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 110 -296
rect 138 -324 172 -296
rect 200 -324 205 -296
rect -205 -358 205 -324
rect -205 -386 -200 -358
rect -172 -386 -138 -358
rect -110 -386 -76 -358
rect -48 -386 -14 -358
rect 14 -386 48 -358
rect 76 -386 110 -358
rect 138 -386 172 -358
rect 200 -386 205 -358
rect -205 -420 205 -386
rect -205 -448 -200 -420
rect -172 -448 -138 -420
rect -110 -448 -76 -420
rect -48 -448 -14 -420
rect 14 -448 48 -420
rect 76 -448 110 -420
rect 138 -448 172 -420
rect 200 -448 205 -420
rect -205 -482 205 -448
rect -205 -510 -200 -482
rect -172 -510 -138 -482
rect -110 -510 -76 -482
rect -48 -510 -14 -482
rect 14 -510 48 -482
rect 76 -510 110 -482
rect 138 -510 172 -482
rect 200 -510 205 -482
rect -205 -544 205 -510
rect -205 -572 -200 -544
rect -172 -572 -138 -544
rect -110 -572 -76 -544
rect -48 -572 -14 -544
rect 14 -572 48 -544
rect 76 -572 110 -544
rect 138 -572 172 -544
rect 200 -572 205 -544
rect -205 -606 205 -572
rect -205 -634 -200 -606
rect -172 -634 -138 -606
rect -110 -634 -76 -606
rect -48 -634 -14 -606
rect 14 -634 48 -606
rect 76 -634 110 -606
rect 138 -634 172 -606
rect 200 -634 205 -606
rect -205 -668 205 -634
rect -205 -696 -200 -668
rect -172 -696 -138 -668
rect -110 -696 -76 -668
rect -48 -696 -14 -668
rect 14 -696 48 -668
rect 76 -696 110 -668
rect 138 -696 172 -668
rect 200 -696 205 -668
rect -205 -701 205 -696
<< via4 >>
rect -200 668 -172 696
rect -138 668 -110 696
rect -76 668 -48 696
rect -14 668 14 696
rect 48 668 76 696
rect 110 668 138 696
rect 172 668 200 696
rect -200 606 -172 634
rect -138 606 -110 634
rect -76 606 -48 634
rect -14 606 14 634
rect 48 606 76 634
rect 110 606 138 634
rect 172 606 200 634
rect -200 544 -172 572
rect -138 544 -110 572
rect -76 544 -48 572
rect -14 544 14 572
rect 48 544 76 572
rect 110 544 138 572
rect 172 544 200 572
rect -200 482 -172 510
rect -138 482 -110 510
rect -76 482 -48 510
rect -14 482 14 510
rect 48 482 76 510
rect 110 482 138 510
rect 172 482 200 510
rect -200 420 -172 448
rect -138 420 -110 448
rect -76 420 -48 448
rect -14 420 14 448
rect 48 420 76 448
rect 110 420 138 448
rect 172 420 200 448
rect -200 358 -172 386
rect -138 358 -110 386
rect -76 358 -48 386
rect -14 358 14 386
rect 48 358 76 386
rect 110 358 138 386
rect 172 358 200 386
rect -200 296 -172 324
rect -138 296 -110 324
rect -76 296 -48 324
rect -14 296 14 324
rect 48 296 76 324
rect 110 296 138 324
rect 172 296 200 324
rect -200 234 -172 262
rect -138 234 -110 262
rect -76 234 -48 262
rect -14 234 14 262
rect 48 234 76 262
rect 110 234 138 262
rect 172 234 200 262
rect -200 172 -172 200
rect -138 172 -110 200
rect -76 172 -48 200
rect -14 172 14 200
rect 48 172 76 200
rect 110 172 138 200
rect 172 172 200 200
rect -200 110 -172 138
rect -138 110 -110 138
rect -76 110 -48 138
rect -14 110 14 138
rect 48 110 76 138
rect 110 110 138 138
rect 172 110 200 138
rect -200 48 -172 76
rect -138 48 -110 76
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect 110 48 138 76
rect 172 48 200 76
rect -200 -14 -172 14
rect -138 -14 -110 14
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect 110 -14 138 14
rect 172 -14 200 14
rect -200 -76 -172 -48
rect -138 -76 -110 -48
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect 110 -76 138 -48
rect 172 -76 200 -48
rect -200 -138 -172 -110
rect -138 -138 -110 -110
rect -76 -138 -48 -110
rect -14 -138 14 -110
rect 48 -138 76 -110
rect 110 -138 138 -110
rect 172 -138 200 -110
rect -200 -200 -172 -172
rect -138 -200 -110 -172
rect -76 -200 -48 -172
rect -14 -200 14 -172
rect 48 -200 76 -172
rect 110 -200 138 -172
rect 172 -200 200 -172
rect -200 -262 -172 -234
rect -138 -262 -110 -234
rect -76 -262 -48 -234
rect -14 -262 14 -234
rect 48 -262 76 -234
rect 110 -262 138 -234
rect 172 -262 200 -234
rect -200 -324 -172 -296
rect -138 -324 -110 -296
rect -76 -324 -48 -296
rect -14 -324 14 -296
rect 48 -324 76 -296
rect 110 -324 138 -296
rect 172 -324 200 -296
rect -200 -386 -172 -358
rect -138 -386 -110 -358
rect -76 -386 -48 -358
rect -14 -386 14 -358
rect 48 -386 76 -358
rect 110 -386 138 -358
rect 172 -386 200 -358
rect -200 -448 -172 -420
rect -138 -448 -110 -420
rect -76 -448 -48 -420
rect -14 -448 14 -420
rect 48 -448 76 -420
rect 110 -448 138 -420
rect 172 -448 200 -420
rect -200 -510 -172 -482
rect -138 -510 -110 -482
rect -76 -510 -48 -482
rect -14 -510 14 -482
rect 48 -510 76 -482
rect 110 -510 138 -482
rect 172 -510 200 -482
rect -200 -572 -172 -544
rect -138 -572 -110 -544
rect -76 -572 -48 -544
rect -14 -572 14 -544
rect 48 -572 76 -544
rect 110 -572 138 -544
rect 172 -572 200 -544
rect -200 -634 -172 -606
rect -138 -634 -110 -606
rect -76 -634 -48 -606
rect -14 -634 14 -606
rect 48 -634 76 -606
rect 110 -634 138 -606
rect 172 -634 200 -606
rect -200 -696 -172 -668
rect -138 -696 -110 -668
rect -76 -696 -48 -668
rect -14 -696 14 -668
rect 48 -696 76 -668
rect 110 -696 138 -668
rect 172 -696 200 -668
<< metal5 >>
rect -208 696 208 704
rect -208 668 -200 696
rect -172 668 -138 696
rect -110 668 -76 696
rect -48 668 -14 696
rect 14 668 48 696
rect 76 668 110 696
rect 138 668 172 696
rect 200 668 208 696
rect -208 634 208 668
rect -208 606 -200 634
rect -172 606 -138 634
rect -110 606 -76 634
rect -48 606 -14 634
rect 14 606 48 634
rect 76 606 110 634
rect 138 606 172 634
rect 200 606 208 634
rect -208 572 208 606
rect -208 544 -200 572
rect -172 544 -138 572
rect -110 544 -76 572
rect -48 544 -14 572
rect 14 544 48 572
rect 76 544 110 572
rect 138 544 172 572
rect 200 544 208 572
rect -208 510 208 544
rect -208 482 -200 510
rect -172 482 -138 510
rect -110 482 -76 510
rect -48 482 -14 510
rect 14 482 48 510
rect 76 482 110 510
rect 138 482 172 510
rect 200 482 208 510
rect -208 448 208 482
rect -208 420 -200 448
rect -172 420 -138 448
rect -110 420 -76 448
rect -48 420 -14 448
rect 14 420 48 448
rect 76 420 110 448
rect 138 420 172 448
rect 200 420 208 448
rect -208 386 208 420
rect -208 358 -200 386
rect -172 358 -138 386
rect -110 358 -76 386
rect -48 358 -14 386
rect 14 358 48 386
rect 76 358 110 386
rect 138 358 172 386
rect 200 358 208 386
rect -208 324 208 358
rect -208 296 -200 324
rect -172 296 -138 324
rect -110 296 -76 324
rect -48 296 -14 324
rect 14 296 48 324
rect 76 296 110 324
rect 138 296 172 324
rect 200 296 208 324
rect -208 262 208 296
rect -208 234 -200 262
rect -172 234 -138 262
rect -110 234 -76 262
rect -48 234 -14 262
rect 14 234 48 262
rect 76 234 110 262
rect 138 234 172 262
rect 200 234 208 262
rect -208 200 208 234
rect -208 172 -200 200
rect -172 172 -138 200
rect -110 172 -76 200
rect -48 172 -14 200
rect 14 172 48 200
rect 76 172 110 200
rect 138 172 172 200
rect 200 172 208 200
rect -208 138 208 172
rect -208 110 -200 138
rect -172 110 -138 138
rect -110 110 -76 138
rect -48 110 -14 138
rect 14 110 48 138
rect 76 110 110 138
rect 138 110 172 138
rect 200 110 208 138
rect -208 76 208 110
rect -208 48 -200 76
rect -172 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 172 76
rect 200 48 208 76
rect -208 14 208 48
rect -208 -14 -200 14
rect -172 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 172 14
rect 200 -14 208 14
rect -208 -48 208 -14
rect -208 -76 -200 -48
rect -172 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 172 -48
rect 200 -76 208 -48
rect -208 -110 208 -76
rect -208 -138 -200 -110
rect -172 -138 -138 -110
rect -110 -138 -76 -110
rect -48 -138 -14 -110
rect 14 -138 48 -110
rect 76 -138 110 -110
rect 138 -138 172 -110
rect 200 -138 208 -110
rect -208 -172 208 -138
rect -208 -200 -200 -172
rect -172 -200 -138 -172
rect -110 -200 -76 -172
rect -48 -200 -14 -172
rect 14 -200 48 -172
rect 76 -200 110 -172
rect 138 -200 172 -172
rect 200 -200 208 -172
rect -208 -234 208 -200
rect -208 -262 -200 -234
rect -172 -262 -138 -234
rect -110 -262 -76 -234
rect -48 -262 -14 -234
rect 14 -262 48 -234
rect 76 -262 110 -234
rect 138 -262 172 -234
rect 200 -262 208 -234
rect -208 -296 208 -262
rect -208 -324 -200 -296
rect -172 -324 -138 -296
rect -110 -324 -76 -296
rect -48 -324 -14 -296
rect 14 -324 48 -296
rect 76 -324 110 -296
rect 138 -324 172 -296
rect 200 -324 208 -296
rect -208 -358 208 -324
rect -208 -386 -200 -358
rect -172 -386 -138 -358
rect -110 -386 -76 -358
rect -48 -386 -14 -358
rect 14 -386 48 -358
rect 76 -386 110 -358
rect 138 -386 172 -358
rect 200 -386 208 -358
rect -208 -420 208 -386
rect -208 -448 -200 -420
rect -172 -448 -138 -420
rect -110 -448 -76 -420
rect -48 -448 -14 -420
rect 14 -448 48 -420
rect 76 -448 110 -420
rect 138 -448 172 -420
rect 200 -448 208 -420
rect -208 -482 208 -448
rect -208 -510 -200 -482
rect -172 -510 -138 -482
rect -110 -510 -76 -482
rect -48 -510 -14 -482
rect 14 -510 48 -482
rect 76 -510 110 -482
rect 138 -510 172 -482
rect 200 -510 208 -482
rect -208 -544 208 -510
rect -208 -572 -200 -544
rect -172 -572 -138 -544
rect -110 -572 -76 -544
rect -48 -572 -14 -544
rect 14 -572 48 -544
rect 76 -572 110 -544
rect 138 -572 172 -544
rect 200 -572 208 -544
rect -208 -606 208 -572
rect -208 -634 -200 -606
rect -172 -634 -138 -606
rect -110 -634 -76 -606
rect -48 -634 -14 -606
rect 14 -634 48 -606
rect 76 -634 110 -606
rect 138 -634 172 -606
rect 200 -634 208 -606
rect -208 -668 208 -634
rect -208 -696 -200 -668
rect -172 -696 -138 -668
rect -110 -696 -76 -668
rect -48 -696 -14 -668
rect 14 -696 48 -668
rect 76 -696 110 -668
rect 138 -696 172 -668
rect 200 -696 208 -668
rect -208 -704 208 -696
<< end >>
