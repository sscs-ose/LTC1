magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2366 -2118 2366 2118
<< pwell >>
rect -366 -118 366 118
<< nmos >>
rect -254 -50 -154 50
rect -50 -50 50 50
rect 154 -50 254 50
<< ndiff >>
rect -342 23 -254 50
rect -342 -23 -329 23
rect -283 -23 -254 23
rect -342 -50 -254 -23
rect -154 23 -50 50
rect -154 -23 -125 23
rect -79 -23 -50 23
rect -154 -50 -50 -23
rect 50 23 154 50
rect 50 -23 79 23
rect 125 -23 154 23
rect 50 -50 154 -23
rect 254 23 342 50
rect 254 -23 283 23
rect 329 -23 342 23
rect 254 -50 342 -23
<< ndiffc >>
rect -329 -23 -283 23
rect -125 -23 -79 23
rect 79 -23 125 23
rect 283 -23 329 23
<< polysilicon >>
rect -254 50 -154 94
rect -50 50 50 94
rect 154 50 254 94
rect -254 -94 -154 -50
rect -50 -94 50 -50
rect 154 -94 254 -50
<< metal1 >>
rect -329 23 -283 48
rect -329 -48 -283 -23
rect -125 23 -79 48
rect -125 -48 -79 -23
rect 79 23 125 48
rect 79 -48 125 -23
rect 283 23 329 48
rect 283 -48 329 -23
<< end >>
