* NGSPICE file created from AND_flat.ext - technology: gf180mcuC

.subckt AND_flat A B OUT VDD VSS
X0 a_176_156# A.t0 a_28_145# VSS.t3 nfet_03v3 ad=89.8f pd=0.92u as=0.155p ps=1.64u w=0.25u l=0.28u
X1 VDD B.t0 a_176_156# VDD.t2 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 a_28_145# B.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.155p pd=1.64u as=89.8f ps=0.92u w=0.25u l=0.28u
X3 VSS B.t2 a_28_145# VSS.t6 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X4 OUT a_176_156# VDD.t6 VDD.t5 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X5 a_28_145# A.t1 a_176_156# VSS.t2 nfet_03v3 ad=89.8f pd=0.92u as=89.8f ps=0.92u w=0.25u l=0.28u
X6 a_176_156# A.t2 VDD.t1 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X7 OUT a_176_156# VSS.t5 VSS.t4 nfet_03v3 ad=0.155p pd=1.64u as=0.155p ps=1.64u w=0.25u l=0.28u
R0 A.n0 A.t2 32.0684
R1 A.n1 A.n0 18.3194
R2 A.n1 A.t0 12.0032
R3 A.n0 A.t1 10.8201
R4 A A.n1 4.14206
R5 VSS.n5 VSS.t6 745.903
R6 VSS.n5 VSS.t0 372.952
R7 VSS.n2 VSS.t4 338.298
R8 VSS.n8 VSS.t2 319.673
R9 VSS.n9 VSS.t3 198.53
R10 VSS.n2 VSS.t5 9.13659
R11 VSS.n1 VSS.n0 5.6705
R12 VSS.n1 VSS.t1 5.6705
R13 VSS.n9 VSS.n8 5.2005
R14 VSS.n6 VSS.n5 5.2005
R15 VSS.n4 VSS.n3 5.2005
R16 VSS.n7 VSS.n1 3.46659
R17 VSS.n6 VSS.n4 0.1955
R18 VSS VSS.n9 0.0944474
R19 VSS.n4 VSS.n2 0.0715526
R20 VSS VSS.n7 0.0676053
R21 VSS.n7 VSS.n6 0.0226053
R22 B B.t0 75.0339
R23 B.t0 B.n0 40.4981
R24 B.n0 B.t1 30.7213
R25 B.n0 B.t2 13.688
R26 VDD.n7 VDD.t0 170.888
R27 VDD.n2 VDD.t5 147.74
R28 VDD.n7 VDD.t1 6.74137
R29 VDD.n1 VDD.t6 3.6405
R30 VDD.n1 VDD.n0 3.6405
R31 VDD.n6 VDD.n5 3.1505
R32 VDD.n5 VDD.n4 3.1505
R33 VDD.n2 VDD.n1 3.10137
R34 VDD.n5 VDD.n3 2.17828
R35 VDD.n4 VDD.t2 1.78941
R36 VDD VDD.n7 0.15489
R37 VDD.n6 VDD.n2 0.0597683
R38 VDD VDD.n6 0.0209878
R39 OUT.n2 OUT.n0 9.37773
R40 OUT.n2 OUT.n1 7.06778
R41 OUT OUT.n2 0.0502872
C0 VDD OUT 0.0845f
C1 a_28_145# OUT 0.0315f
C2 VDD a_176_156# 0.403f
C3 a_28_145# a_176_156# 0.319f
C4 VDD A 0.119f
C5 A a_28_145# 0.109f
C6 a_176_156# OUT 0.0738f
C7 A OUT 2.31e-19
C8 VDD B 0.489f
C9 B a_28_145# 0.0441f
C10 A a_176_156# 0.122f
C11 B OUT 0.00142f
C12 B a_176_156# 0.0859f
C13 B A 0.0797f
C14 VDD a_28_145# 0.0109f
.ends

