magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2032 11097 17032 71968
use gf180mcu_fd_io__fill5  gf180mcu_fd_io__fill5_0
array 0 14 1000 0 0 70000
timestamp 1713338890
transform 1 0 0 0 1 0
box -32 13097 1032 69968
<< end >>
