magic
tech gf180mcuD
magscale 1 10
timestamp 1713971188
<< checkpaint >>
rect -3158 -3186 4262 2549
<< nwell >>
rect -38 542 1117 549
rect -38 538 1139 542
rect -38 521 1157 538
rect -136 477 1157 521
rect -136 461 149 477
rect -138 445 149 461
rect 963 458 1157 477
rect 974 449 1157 458
rect 982 445 1138 449
rect -138 434 100 445
rect 1104 443 1125 445
rect -138 425 88 434
rect -38 -31 25 425
rect 174 36 502 106
rect 605 25 933 95
rect 1108 -31 1117 443
<< psubdiff >>
rect 490 -962 811 -935
rect 490 -1008 526 -962
rect 572 -1008 675 -962
rect 721 -1008 811 -962
rect 490 -1029 811 -1008
<< nsubdiff >>
rect -136 502 57 521
rect -136 456 -119 502
rect 21 456 57 502
rect -136 441 57 456
<< psubdiffcont >>
rect 526 -1008 572 -962
rect 675 -1008 721 -962
<< nsubdiffcont >>
rect -119 456 21 502
<< polysilicon >>
rect 174 95 502 106
rect 822 95 934 110
rect 174 49 206 95
rect 252 49 502 95
rect 174 36 502 49
rect 605 70 934 95
rect 605 53 947 70
rect 605 25 884 53
rect 822 7 884 25
rect 930 7 947 53
rect 822 -7 947 7
rect 174 -97 502 -61
rect 606 -97 934 -61
rect 174 -448 286 -379
rect 169 -460 286 -448
rect 169 -506 183 -460
rect 229 -506 286 -460
rect 169 -533 286 -506
rect 174 -555 286 -533
rect 390 -466 502 -449
rect 390 -512 423 -466
rect 469 -512 502 -466
rect 390 -544 502 -512
rect 606 -474 718 -378
rect 606 -520 651 -474
rect 697 -520 718 -474
rect 606 -562 718 -520
rect 1078 -822 1203 -803
rect 1078 -834 1131 -822
rect 821 -868 1131 -834
rect 1177 -868 1203 -822
rect 821 -895 1203 -868
<< polycontact >>
rect 206 49 252 95
rect 884 7 930 53
rect 183 -506 229 -460
rect 423 -512 469 -466
rect 651 -520 697 -474
rect 1131 -868 1177 -822
<< metal1 >>
rect 1062 543 2160 544
rect -1068 502 2160 543
rect -1068 456 -119 502
rect 21 456 2160 502
rect -1068 445 2160 456
rect -233 425 158 445
rect 99 255 145 352
rect 78 243 145 255
rect 78 191 90 243
rect 142 191 145 243
rect 78 179 145 191
rect 99 132 145 179
rect 195 95 264 106
rect -286 24 -240 53
rect 195 49 206 95
rect 252 49 264 95
rect 195 38 264 49
rect -298 8 -215 24
rect -1158 -39 -862 -34
rect -1158 -40 -815 -39
rect -1158 -85 -862 -40
rect -298 -44 -281 8
rect -229 3 -215 8
rect 195 3 254 38
rect -229 -43 254 3
rect -229 -44 -215 -43
rect -298 -59 -215 -44
rect -1158 -90 -815 -85
rect -1158 -100 -862 -90
rect -1158 -698 -1092 -100
rect 99 -239 145 -132
rect 86 -251 162 -239
rect 86 -303 98 -251
rect 150 -303 162 -251
rect 86 -315 162 -303
rect 99 -352 145 -315
rect 315 -352 361 445
rect 531 255 577 354
rect 531 243 598 255
rect 531 191 534 243
rect 586 191 598 243
rect 531 179 598 191
rect 531 132 577 179
rect 494 15 572 27
rect 494 -14 508 15
rect 453 -37 508 -14
rect 560 -14 572 15
rect 747 -14 793 352
rect 963 256 1011 352
rect 949 244 1025 256
rect 949 192 961 244
rect 1013 192 1025 244
rect 949 180 1025 192
rect 963 132 1011 180
rect 1073 76 1150 91
rect 873 53 934 65
rect 1073 53 1086 76
rect 873 7 884 53
rect 930 24 1086 53
rect 1138 53 1150 76
rect 1138 24 2017 53
rect 930 7 2017 24
rect 873 -5 934 7
rect 560 -37 793 -14
rect 453 -60 793 -37
rect 531 -239 577 -132
rect 511 -251 580 -239
rect 511 -303 523 -251
rect 575 -303 580 -251
rect 511 -315 580 -303
rect 531 -352 577 -315
rect 747 -352 793 -60
rect 1088 -90 1453 -44
rect 963 -239 1015 -132
rect 963 -251 1028 -239
rect 963 -303 964 -251
rect 1016 -303 1028 -251
rect 963 -315 1028 -303
rect 963 -352 1015 -315
rect -35 -460 241 -448
rect -35 -506 183 -460
rect 229 -506 241 -460
rect -35 -518 241 -506
rect 408 -463 485 -450
rect 408 -515 420 -463
rect 472 -515 485 -463
rect -998 -528 -86 -519
rect -998 -580 -938 -528
rect -886 -529 -86 -528
rect -886 -580 -792 -529
rect -998 -581 -792 -580
rect -740 -532 -86 -529
rect -740 -533 -155 -532
rect -740 -581 -461 -533
rect -998 -585 -461 -581
rect -409 -534 -155 -533
rect -409 -585 -315 -534
rect -998 -586 -315 -585
rect -263 -584 -155 -534
rect -103 -584 -86 -532
rect -263 -586 -86 -584
rect -998 -600 -86 -586
rect -35 -698 31 -518
rect 408 -527 485 -515
rect 640 -474 697 -463
rect 1088 -474 1134 -90
rect 640 -520 651 -474
rect 697 -520 1134 -474
rect 640 -531 697 -520
rect 315 -674 361 -579
rect -1158 -764 31 -698
rect 300 -686 376 -674
rect 300 -738 312 -686
rect 364 -738 376 -686
rect 300 -750 376 -738
rect 99 -835 145 -763
rect 315 -799 361 -750
rect -144 -881 145 -835
rect -144 -1112 -98 -881
rect 747 -927 793 -579
rect 950 -657 1026 -645
rect 950 -709 962 -657
rect 1014 -709 1026 -657
rect 950 -721 1026 -709
rect 1119 -816 1196 -803
rect 1119 -868 1131 -816
rect 1183 -868 1196 -816
rect 1119 -880 1196 -868
rect 1446 -927 1571 -521
rect 1677 -927 1802 -520
rect 1925 -927 2050 -520
rect 2137 -927 2262 -520
rect -1 -962 2262 -927
rect -1 -963 398 -962
rect -1 -964 230 -963
rect -1 -1016 34 -964
rect 86 -1015 230 -964
rect 282 -1014 398 -963
rect 450 -1008 526 -962
rect 572 -1008 675 -962
rect 721 -1008 2262 -962
rect 450 -1014 2262 -1008
rect 282 -1015 2262 -1014
rect 86 -1016 2262 -1015
rect -1 -1048 2262 -1016
rect 941 -1112 1018 -1110
rect -144 -1122 1018 -1112
rect -144 -1158 953 -1122
rect 941 -1174 953 -1158
rect 1005 -1174 1018 -1122
rect 941 -1186 1018 -1174
<< via1 >>
rect 90 191 142 243
rect -281 -44 -229 8
rect 98 -303 150 -251
rect 534 191 586 243
rect 508 -37 560 15
rect 961 192 1013 244
rect 1086 24 1138 76
rect 523 -303 575 -251
rect 964 -303 1016 -251
rect 420 -466 472 -463
rect 420 -512 423 -466
rect 423 -512 469 -466
rect 469 -512 472 -466
rect 420 -515 472 -512
rect -938 -580 -886 -528
rect -792 -581 -740 -529
rect -461 -585 -409 -533
rect -315 -586 -263 -534
rect -155 -584 -103 -532
rect 312 -738 364 -686
rect 962 -709 1014 -657
rect 1131 -822 1183 -816
rect 1131 -868 1177 -822
rect 1177 -868 1183 -822
rect 34 -1016 86 -964
rect 230 -1015 282 -963
rect 398 -1014 450 -962
rect 953 -1174 1005 -1122
<< metal2 >>
rect 78 246 145 255
rect 535 246 598 255
rect 949 246 1025 256
rect 78 244 1025 246
rect 78 243 961 244
rect 78 191 90 243
rect 142 191 534 243
rect 586 192 961 243
rect 1013 192 1025 244
rect 586 191 1025 192
rect 78 188 1025 191
rect 78 179 145 188
rect 535 179 598 188
rect 949 180 1025 188
rect 1073 76 1150 91
rect 1073 53 1086 76
rect -298 10 -215 24
rect -298 -46 -286 10
rect -230 8 -215 10
rect -229 -44 -215 8
rect 494 15 572 27
rect 494 -4 508 15
rect -230 -46 -215 -44
rect -298 -59 -215 -46
rect -99 -37 508 -4
rect 560 -4 572 15
rect 1049 24 1086 53
rect 1138 53 1150 76
rect 1138 24 1186 53
rect 1049 -3 1186 24
rect 560 -37 701 -4
rect -99 -60 701 -37
rect -99 -374 -43 -60
rect 86 -247 162 -239
rect 511 -247 580 -239
rect 963 -247 1028 -239
rect 86 -251 1028 -247
rect 86 -303 98 -251
rect 150 -303 523 -251
rect 575 -303 964 -251
rect 1016 -303 1028 -251
rect 86 -307 1028 -303
rect 86 -315 162 -307
rect 511 -315 580 -307
rect 963 -315 1028 -307
rect -99 -430 38 -374
rect -1040 -528 -81 -518
rect -1040 -580 -938 -528
rect -886 -529 -81 -528
rect -886 -580 -792 -529
rect -1040 -581 -792 -580
rect -740 -532 -81 -529
rect -740 -533 -155 -532
rect -740 -581 -461 -533
rect -1040 -585 -461 -581
rect -409 -534 -155 -533
rect -409 -585 -315 -534
rect -1040 -586 -315 -585
rect -263 -584 -155 -534
rect -103 -584 -81 -532
rect -263 -586 -81 -584
rect -1040 -596 -81 -586
rect -986 -943 -908 -596
rect -748 -943 -670 -596
rect -986 -947 -670 -943
rect -531 -947 -453 -596
rect -331 -943 -253 -596
rect -159 -943 -81 -596
rect -18 -684 38 -430
rect 408 -461 485 -450
rect 408 -517 419 -461
rect 475 -517 485 -461
rect 408 -527 485 -517
rect 950 -657 1026 -645
rect 300 -684 376 -674
rect -18 -686 376 -684
rect -18 -738 312 -686
rect 364 -738 376 -686
rect -18 -740 376 -738
rect 300 -750 376 -740
rect 950 -709 962 -657
rect 1014 -709 1026 -657
rect 950 -721 1026 -709
rect -331 -947 -81 -943
rect -986 -962 467 -947
rect -986 -963 398 -962
rect -986 -964 230 -963
rect -986 -1016 34 -964
rect 86 -1015 230 -964
rect 282 -1014 398 -963
rect 450 -1014 467 -962
rect 282 -1015 467 -1014
rect 86 -1016 467 -1015
rect -986 -1021 467 -1016
rect -748 -1025 467 -1021
rect 950 -1110 1018 -721
rect 1130 -759 1186 -3
rect 1129 -803 1186 -759
rect 1119 -816 1196 -803
rect 1119 -868 1131 -816
rect 1183 -868 1196 -816
rect 1119 -880 1196 -868
rect 941 -1122 1018 -1110
rect 941 -1174 953 -1122
rect 1005 -1174 1018 -1122
rect 941 -1186 1018 -1174
<< via2 >>
rect -286 8 -230 10
rect -286 -44 -281 8
rect -281 -44 -230 8
rect -286 -46 -230 -44
rect 419 -463 475 -461
rect 419 -515 420 -463
rect 420 -515 472 -463
rect 472 -515 475 -463
rect 419 -517 475 -515
<< metal3 >>
rect -297 10 -216 24
rect -297 -46 -286 10
rect -230 -46 -216 10
rect -297 -58 -216 -46
rect -288 -447 -229 -58
rect -288 -450 467 -447
rect -288 -461 485 -450
rect -288 -506 419 -461
rect 408 -517 419 -506
rect 475 -517 485 -461
rect 408 -527 485 -517
use inverter_magic  inverter_magic_0
timestamp 1713185578
transform 1 0 1117 0 1 -31
box 0 -569 1108 580
use inverter_magic  inverter_magic_1
timestamp 1713185578
transform 1 0 -1146 0 1 -31
box 0 -569 1108 580
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_0
timestamp 1713185578
transform 1 0 878 0 1 -689
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_1
timestamp 1713185578
transform 1 0 230 0 1 -689
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_2
timestamp 1713185578
transform 1 0 446 0 1 -689
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_3
timestamp 1713185578
transform 1 0 662 0 1 -689
box -168 -180 168 180
use pmos_3p3_VZX6F7  pmos_3p3_VZX6F7_0
timestamp 1713185578
transform 1 0 770 0 1 -242
box -338 -242 338 242
use pmos_3p3_VZX6F7  pmos_3p3_VZX6F7_1
timestamp 1713185578
transform 1 0 338 0 1 242
box -338 -242 338 242
use pmos_3p3_VZX6F7  pmos_3p3_VZX6F7_2
timestamp 1713185578
transform 1 0 770 0 1 242
box -338 -242 338 242
use pmos_3p3_VZX6F7  pmos_3p3_VZX6F7_3
timestamp 1713185578
transform 1 0 338 0 1 -242
box -338 -242 338 242
<< labels >>
flabel psubdiffcont 549 -984 549 -984 0 FreeSans 750 0 0 0 VSS
flabel metal1 s 144 -488 144 -488 0 FreeSans 750 0 0 0 A
port 1 nsew
flabel metal1 s 984 -497 984 -497 0 FreeSans 750 0 0 0 B
port 2 nsew
flabel metal1 s 764 -22 764 -22 0 FreeSans 750 0 0 0 OUT
port 3 nsew
flabel metal1 s -50 483 -50 483 0 FreeSans 1250 0 0 0 VDD
port 4 nsew
<< end >>
