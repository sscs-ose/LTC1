magic
tech gf180mcuC
magscale 1 10
timestamp 1691670472
<< nwell >>
rect 0 310 1172 901
<< pwell >>
rect 222 0 822 236
<< nmos >>
rect 334 68 390 168
rect 494 68 550 168
rect 654 68 710 168
<< pmos >>
rect 174 440 230 640
rect 334 440 390 640
rect 494 440 550 640
rect 654 440 710 640
rect 942 440 998 640
<< ndiff >>
rect 246 155 334 168
rect 246 81 259 155
rect 305 81 334 155
rect 246 68 334 81
rect 390 155 494 168
rect 390 81 419 155
rect 465 81 494 155
rect 390 68 494 81
rect 550 155 654 168
rect 550 81 579 155
rect 625 81 654 155
rect 550 68 654 81
rect 710 155 798 168
rect 710 81 739 155
rect 785 81 798 155
rect 710 68 798 81
<< pdiff >>
rect 86 627 174 640
rect 86 453 99 627
rect 145 453 174 627
rect 86 440 174 453
rect 230 627 334 640
rect 230 453 259 627
rect 305 453 334 627
rect 230 440 334 453
rect 390 627 494 640
rect 390 453 419 627
rect 465 453 494 627
rect 390 440 494 453
rect 550 627 654 640
rect 550 453 579 627
rect 625 453 654 627
rect 550 440 654 453
rect 710 627 798 640
rect 710 453 739 627
rect 785 453 798 627
rect 710 440 798 453
rect 854 627 942 640
rect 854 453 867 627
rect 913 453 942 627
rect 854 440 942 453
rect 998 627 1086 640
rect 998 453 1027 627
rect 1073 453 1086 627
rect 998 440 1086 453
<< ndiffc >>
rect 259 81 305 155
rect 419 81 465 155
rect 579 81 625 155
rect 739 81 785 155
<< pdiffc >>
rect 99 453 145 627
rect 259 453 305 627
rect 419 453 465 627
rect 579 453 625 627
rect 739 453 785 627
rect 867 453 913 627
rect 1027 453 1073 627
<< psubdiff >>
rect 251 -161 793 -148
rect 251 -207 264 -161
rect 310 -207 358 -161
rect 404 -207 452 -161
rect 498 -207 546 -161
rect 592 -207 640 -161
rect 686 -207 734 -161
rect 780 -207 793 -161
rect 251 -220 793 -207
<< nsubdiff >>
rect 24 855 1143 868
rect 24 809 37 855
rect 83 809 131 855
rect 177 809 225 855
rect 271 809 319 855
rect 365 809 413 855
rect 459 809 507 855
rect 553 809 601 855
rect 647 809 708 855
rect 754 809 802 855
rect 848 809 896 855
rect 942 809 990 855
rect 1036 809 1084 855
rect 1130 809 1143 855
rect 24 796 1143 809
<< psubdiffcont >>
rect 264 -207 310 -161
rect 358 -207 404 -161
rect 452 -207 498 -161
rect 546 -207 592 -161
rect 640 -207 686 -161
rect 734 -207 780 -161
<< nsubdiffcont >>
rect 37 809 83 855
rect 131 809 177 855
rect 225 809 271 855
rect 319 809 365 855
rect 413 809 459 855
rect 507 809 553 855
rect 601 809 647 855
rect 708 809 754 855
rect 802 809 848 855
rect 896 809 942 855
rect 990 809 1036 855
rect 1084 809 1130 855
<< polysilicon >>
rect 174 640 230 684
rect 334 640 390 684
rect 494 640 550 684
rect 654 640 710 684
rect 942 640 998 684
rect 174 420 230 440
rect 334 420 390 440
rect 174 364 390 420
rect 178 297 250 305
rect 334 297 390 364
rect 178 292 390 297
rect 178 246 191 292
rect 237 246 390 292
rect 178 241 390 246
rect 178 233 250 241
rect 334 168 390 241
rect 494 420 550 440
rect 654 420 710 440
rect 494 364 710 420
rect 494 168 550 364
rect 622 276 694 284
rect 942 276 998 440
rect 622 271 998 276
rect 622 225 635 271
rect 681 225 998 271
rect 622 220 998 225
rect 622 212 710 220
rect 654 168 710 212
rect 334 24 390 68
rect 132 -24 204 -16
rect 494 -24 550 68
rect 654 24 710 68
rect 132 -29 550 -24
rect 132 -75 145 -29
rect 191 -75 550 -29
rect 132 -80 550 -75
rect 132 -88 204 -80
<< polycontact >>
rect 191 246 237 292
rect 635 225 681 271
rect 145 -75 191 -29
<< metal1 >>
rect 0 855 1172 888
rect 0 809 37 855
rect 83 809 131 855
rect 177 809 225 855
rect 271 809 319 855
rect 365 809 413 855
rect 459 809 507 855
rect 553 809 601 855
rect 647 809 708 855
rect 754 809 802 855
rect 848 809 896 855
rect 942 809 990 855
rect 1036 809 1084 855
rect 1130 809 1172 855
rect 0 776 1172 809
rect 99 627 145 638
rect 99 396 145 453
rect 259 627 305 776
rect 259 442 305 453
rect 419 684 785 730
rect 419 627 465 684
rect 419 396 465 453
rect 99 350 465 396
rect 579 627 625 638
rect 180 297 248 303
rect 97 292 248 297
rect 97 246 191 292
rect 237 246 248 292
rect 579 282 625 453
rect 739 627 785 684
rect 739 442 785 453
rect 867 627 913 638
rect 867 344 913 453
rect 1027 627 1073 776
rect 1027 442 1073 453
rect 867 298 1087 344
rect 579 271 692 282
rect 579 258 635 271
rect 97 241 248 246
rect 180 235 248 241
rect 419 225 635 258
rect 681 225 692 271
rect 867 228 913 298
rect 419 214 692 225
rect 419 212 625 214
rect 259 155 305 166
rect 134 -29 202 -18
rect 100 -75 145 -29
rect 191 -75 202 -29
rect 134 -86 202 -75
rect 259 -128 305 81
rect 419 155 465 212
rect 739 182 913 228
rect 419 70 465 81
rect 579 155 625 166
rect 579 -128 625 81
rect 739 155 785 182
rect 739 70 785 81
rect 222 -161 822 -128
rect 222 -207 264 -161
rect 310 -207 358 -161
rect 404 -207 452 -161
rect 498 -207 546 -161
rect 592 -207 640 -161
rect 686 -207 734 -161
rect 780 -207 822 -161
rect 222 -240 822 -207
<< labels >>
flabel metal1 577 832 577 832 0 FreeSans 320 0 0 0 VDD
port 5 nsew
flabel metal1 530 -184 530 -184 0 FreeSans 320 0 0 0 VSS
port 6 nsew
flabel polycontact 214 269 214 269 0 FreeSans 320 0 0 0 A
port 7 nsew
flabel polycontact 168 -52 168 -52 0 FreeSans 320 0 0 0 B
port 8 nsew
flabel metal1 1064 322 1064 322 0 FreeSans 320 0 0 0 OUT
port 4 nsew
<< end >>
