magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2136 -2042 2136 2042
<< polysilicon >>
rect -136 23 136 42
rect -136 -23 -117 23
rect 117 -23 136 23
rect -136 -42 136 -23
<< polycontact >>
rect -117 -23 117 23
<< metal1 >>
rect -128 23 128 34
rect -128 -23 -117 23
rect 117 -23 128 23
rect -128 -34 128 -23
<< end >>
