magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1262 -1073 1262 1073
<< metal1 >>
rect -262 67 262 73
rect -262 41 -256 67
rect -230 41 -202 67
rect -176 41 -148 67
rect -122 41 -94 67
rect -68 41 -40 67
rect -14 41 14 67
rect 40 41 68 67
rect 94 41 122 67
rect 148 41 176 67
rect 202 41 230 67
rect 256 41 262 67
rect -262 13 262 41
rect -262 -13 -256 13
rect -230 -13 -202 13
rect -176 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 176 13
rect 202 -13 230 13
rect 256 -13 262 13
rect -262 -41 262 -13
rect -262 -67 -256 -41
rect -230 -67 -202 -41
rect -176 -67 -148 -41
rect -122 -67 -94 -41
rect -68 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 68 -41
rect 94 -67 122 -41
rect 148 -67 176 -41
rect 202 -67 230 -41
rect 256 -67 262 -41
rect -262 -73 262 -67
<< via1 >>
rect -256 41 -230 67
rect -202 41 -176 67
rect -148 41 -122 67
rect -94 41 -68 67
rect -40 41 -14 67
rect 14 41 40 67
rect 68 41 94 67
rect 122 41 148 67
rect 176 41 202 67
rect 230 41 256 67
rect -256 -13 -230 13
rect -202 -13 -176 13
rect -148 -13 -122 13
rect -94 -13 -68 13
rect -40 -13 -14 13
rect 14 -13 40 13
rect 68 -13 94 13
rect 122 -13 148 13
rect 176 -13 202 13
rect 230 -13 256 13
rect -256 -67 -230 -41
rect -202 -67 -176 -41
rect -148 -67 -122 -41
rect -94 -67 -68 -41
rect -40 -67 -14 -41
rect 14 -67 40 -41
rect 68 -67 94 -41
rect 122 -67 148 -41
rect 176 -67 202 -41
rect 230 -67 256 -41
<< metal2 >>
rect -262 67 262 73
rect -262 41 -256 67
rect -230 41 -202 67
rect -176 41 -148 67
rect -122 41 -94 67
rect -68 41 -40 67
rect -14 41 14 67
rect 40 41 68 67
rect 94 41 122 67
rect 148 41 176 67
rect 202 41 230 67
rect 256 41 262 67
rect -262 13 262 41
rect -262 -13 -256 13
rect -230 -13 -202 13
rect -176 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 176 13
rect 202 -13 230 13
rect 256 -13 262 13
rect -262 -41 262 -13
rect -262 -67 -256 -41
rect -230 -67 -202 -41
rect -176 -67 -148 -41
rect -122 -67 -94 -41
rect -68 -67 -40 -41
rect -14 -67 14 -41
rect 40 -67 68 -41
rect 94 -67 122 -41
rect 148 -67 176 -41
rect 202 -67 230 -41
rect 256 -67 262 -41
rect -262 -73 262 -67
<< end >>
