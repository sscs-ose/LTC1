magic
tech gf180mcuC
magscale 1 10
timestamp 1698845364
<< nwell >>
rect 71 2748 5251 2749
rect -4931 1088 -2920 2741
rect -2528 1095 -517 2748
rect 71 1096 7118 2748
rect 5511 1095 7118 1096
rect -4931 -4072 -2920 -940
rect -2528 -4065 -517 -933
rect 61 -996 945 -61
rect 1831 -933 5251 -932
rect 61 -3937 945 -2211
rect 1831 -4064 7118 -933
rect 5511 -4065 7118 -4064
rect 1653 -6092 1892 -6091
rect 71 -6093 5251 -6092
rect -4931 -7753 -2920 -6100
rect -2528 -7746 -517 -6093
rect 71 -7744 7118 -6093
rect 71 -7745 3438 -7744
rect 3644 -7745 7118 -7744
rect 5250 -7746 7118 -7745
rect 5250 -7747 5512 -7746
<< pwell >>
rect -4869 232 -4589 904
rect -4465 232 -4185 904
rect -4062 232 -2982 904
rect -2466 239 -2186 911
rect -2062 239 -1782 911
rect -1659 239 -579 911
rect 133 240 413 912
rect 536 240 1616 912
rect 1893 240 2973 912
rect 3096 240 3376 912
rect 3706 240 3986 912
rect 4109 240 5189 912
rect 5573 239 6653 911
rect 6776 239 7056 911
rect -4869 -756 -4589 -84
rect -4465 -756 -4185 -84
rect -4062 -756 -2982 -84
rect -2466 -749 -2186 -77
rect -2062 -749 -1782 -77
rect -1659 -749 -579 -77
rect 1893 -748 2173 -76
rect 2296 -748 3376 -76
rect 3706 -748 4786 -76
rect 4909 -748 5189 -76
rect 5573 -749 5853 -77
rect 5976 -749 7056 -77
rect 123 -1519 883 -1047
rect 123 -2160 883 -1688
rect -4869 -4928 -4589 -4256
rect -4465 -4928 -4185 -4256
rect -4062 -4928 -2982 -4256
rect -2466 -4921 -2186 -4249
rect -2062 -4921 -1782 -4249
rect -1659 -4921 -579 -4249
rect 123 -4460 883 -3988
rect 1893 -4920 2173 -4248
rect 2296 -4920 3376 -4248
rect 3706 -4920 4786 -4248
rect 4909 -4920 5189 -4248
rect 5573 -4921 5853 -4249
rect 5976 -4921 7056 -4249
rect -4869 -5916 -4589 -5244
rect -4465 -5916 -4185 -5244
rect -4062 -5916 -2982 -5244
rect -2466 -5909 -2186 -5237
rect -2062 -5909 -1782 -5237
rect -1659 -5909 -579 -5237
rect 133 -5908 413 -5236
rect 536 -5908 1616 -5236
rect 1893 -5908 2973 -5236
rect 3096 -5908 3376 -5236
rect 3706 -5908 3986 -5236
rect 4109 -5908 5189 -5236
rect 5573 -5909 6653 -5237
rect 6776 -5909 7056 -5237
<< nmos >>
rect -4757 636 -4701 836
rect -4353 636 -4297 836
rect -3950 636 -3894 836
rect -3790 636 -3734 836
rect -3630 636 -3574 836
rect -3470 636 -3414 836
rect -3310 636 -3254 836
rect -3150 636 -3094 836
rect -2354 643 -2298 843
rect -1950 643 -1894 843
rect -1547 643 -1491 843
rect -1387 643 -1331 843
rect -1227 643 -1171 843
rect -1067 643 -1011 843
rect -907 643 -851 843
rect -747 643 -691 843
rect 245 644 301 844
rect 648 644 704 844
rect 808 644 864 844
rect 968 644 1024 844
rect 1128 644 1184 844
rect 1288 644 1344 844
rect 1448 644 1504 844
rect 2005 644 2061 844
rect 2165 644 2221 844
rect 2325 644 2381 844
rect 2485 644 2541 844
rect 2645 644 2701 844
rect 2805 644 2861 844
rect 3208 644 3264 844
rect 3818 644 3874 844
rect 4221 644 4277 844
rect 4381 644 4437 844
rect 4541 644 4597 844
rect 4701 644 4757 844
rect 4861 644 4917 844
rect 5021 644 5077 844
rect 5685 643 5741 843
rect 5845 643 5901 843
rect 6005 643 6061 843
rect 6165 643 6221 843
rect 6325 643 6381 843
rect 6485 643 6541 843
rect 6888 643 6944 843
rect -4757 300 -4701 500
rect -4353 300 -4297 500
rect -3950 300 -3894 500
rect -3790 300 -3734 500
rect -3630 300 -3574 500
rect -3470 300 -3414 500
rect -3310 300 -3254 500
rect -3150 300 -3094 500
rect -2354 307 -2298 507
rect -1950 307 -1894 507
rect -1547 307 -1491 507
rect -1387 307 -1331 507
rect -1227 307 -1171 507
rect -1067 307 -1011 507
rect -907 307 -851 507
rect -747 307 -691 507
rect 245 308 301 508
rect 648 308 704 508
rect 808 308 864 508
rect 968 308 1024 508
rect 1128 308 1184 508
rect 1288 308 1344 508
rect 1448 308 1504 508
rect 2005 308 2061 508
rect 2165 308 2221 508
rect 2325 308 2381 508
rect 2485 308 2541 508
rect 2645 308 2701 508
rect 2805 308 2861 508
rect 3208 308 3264 508
rect 3818 308 3874 508
rect 4221 308 4277 508
rect 4381 308 4437 508
rect 4541 308 4597 508
rect 4701 308 4757 508
rect 4861 308 4917 508
rect 5021 308 5077 508
rect 5685 307 5741 507
rect 5845 307 5901 507
rect 6005 307 6061 507
rect 6165 307 6221 507
rect 6325 307 6381 507
rect 6485 307 6541 507
rect 6888 307 6944 507
rect -4757 -352 -4701 -152
rect -4353 -352 -4297 -152
rect -3950 -352 -3894 -152
rect -3790 -352 -3734 -152
rect -3630 -352 -3574 -152
rect -3470 -352 -3414 -152
rect -3310 -352 -3254 -152
rect -3150 -352 -3094 -152
rect -2354 -345 -2298 -145
rect -1950 -345 -1894 -145
rect -1547 -345 -1491 -145
rect -1387 -345 -1331 -145
rect -1227 -345 -1171 -145
rect -1067 -345 -1011 -145
rect -907 -345 -851 -145
rect -747 -345 -691 -145
rect -4757 -688 -4701 -488
rect -4353 -688 -4297 -488
rect -3950 -688 -3894 -488
rect -3790 -688 -3734 -488
rect -3630 -688 -3574 -488
rect -3470 -688 -3414 -488
rect -3310 -688 -3254 -488
rect -3150 -688 -3094 -488
rect -2354 -681 -2298 -481
rect -1950 -681 -1894 -481
rect -1547 -681 -1491 -481
rect -1387 -681 -1331 -481
rect -1227 -681 -1171 -481
rect -1067 -681 -1011 -481
rect -907 -681 -851 -481
rect -747 -681 -691 -481
rect 2005 -344 2061 -144
rect 2408 -344 2464 -144
rect 2568 -344 2624 -144
rect 2728 -344 2784 -144
rect 2888 -344 2944 -144
rect 3048 -344 3104 -144
rect 3208 -344 3264 -144
rect 3818 -344 3874 -144
rect 3978 -344 4034 -144
rect 4138 -344 4194 -144
rect 4298 -344 4354 -144
rect 4458 -344 4514 -144
rect 4618 -344 4674 -144
rect 5021 -344 5077 -144
rect 5685 -345 5741 -145
rect 6088 -345 6144 -145
rect 6248 -345 6304 -145
rect 6408 -345 6464 -145
rect 6568 -345 6624 -145
rect 6728 -345 6784 -145
rect 6888 -345 6944 -145
rect 2005 -680 2061 -480
rect 2408 -680 2464 -480
rect 2568 -680 2624 -480
rect 2728 -680 2784 -480
rect 2888 -680 2944 -480
rect 3048 -680 3104 -480
rect 3208 -680 3264 -480
rect 3818 -680 3874 -480
rect 3978 -680 4034 -480
rect 4138 -680 4194 -480
rect 4298 -680 4354 -480
rect 4458 -680 4514 -480
rect 4618 -680 4674 -480
rect 5021 -680 5077 -480
rect 5685 -681 5741 -481
rect 6088 -681 6144 -481
rect 6248 -681 6304 -481
rect 6408 -681 6464 -481
rect 6568 -681 6624 -481
rect 6728 -681 6784 -481
rect 6888 -681 6944 -481
rect 235 -1215 291 -1115
rect 395 -1215 451 -1115
rect 555 -1215 611 -1115
rect 715 -1215 771 -1115
rect 235 -1451 291 -1351
rect 395 -1451 451 -1351
rect 555 -1451 611 -1351
rect 715 -1451 771 -1351
rect 235 -1856 291 -1756
rect 395 -1856 451 -1756
rect 555 -1856 611 -1756
rect 715 -1856 771 -1756
rect 235 -2092 291 -1992
rect 395 -2092 451 -1992
rect 555 -2092 611 -1992
rect 715 -2092 771 -1992
rect 235 -4156 291 -4056
rect 395 -4156 451 -4056
rect 555 -4156 611 -4056
rect 715 -4156 771 -4056
rect -4757 -4524 -4701 -4324
rect -4353 -4524 -4297 -4324
rect -3950 -4524 -3894 -4324
rect -3790 -4524 -3734 -4324
rect -3630 -4524 -3574 -4324
rect -3470 -4524 -3414 -4324
rect -3310 -4524 -3254 -4324
rect -3150 -4524 -3094 -4324
rect -2354 -4517 -2298 -4317
rect -1950 -4517 -1894 -4317
rect -1547 -4517 -1491 -4317
rect -1387 -4517 -1331 -4317
rect -1227 -4517 -1171 -4317
rect -1067 -4517 -1011 -4317
rect -907 -4517 -851 -4317
rect -747 -4517 -691 -4317
rect 235 -4392 291 -4292
rect 395 -4392 451 -4292
rect 555 -4392 611 -4292
rect 715 -4392 771 -4292
rect 2005 -4516 2061 -4316
rect 2408 -4516 2464 -4316
rect 2568 -4516 2624 -4316
rect 2728 -4516 2784 -4316
rect 2888 -4516 2944 -4316
rect 3048 -4516 3104 -4316
rect 3208 -4516 3264 -4316
rect 3818 -4516 3874 -4316
rect 3978 -4516 4034 -4316
rect 4138 -4516 4194 -4316
rect 4298 -4516 4354 -4316
rect 4458 -4516 4514 -4316
rect 4618 -4516 4674 -4316
rect 5021 -4516 5077 -4316
rect 5685 -4517 5741 -4317
rect 6088 -4517 6144 -4317
rect 6248 -4517 6304 -4317
rect 6408 -4517 6464 -4317
rect 6568 -4517 6624 -4317
rect 6728 -4517 6784 -4317
rect 6888 -4517 6944 -4317
rect -4757 -4860 -4701 -4660
rect -4353 -4860 -4297 -4660
rect -3950 -4860 -3894 -4660
rect -3790 -4860 -3734 -4660
rect -3630 -4860 -3574 -4660
rect -3470 -4860 -3414 -4660
rect -3310 -4860 -3254 -4660
rect -3150 -4860 -3094 -4660
rect -2354 -4853 -2298 -4653
rect -1950 -4853 -1894 -4653
rect -1547 -4853 -1491 -4653
rect -1387 -4853 -1331 -4653
rect -1227 -4853 -1171 -4653
rect -1067 -4853 -1011 -4653
rect -907 -4853 -851 -4653
rect -747 -4853 -691 -4653
rect 2005 -4852 2061 -4652
rect 2408 -4852 2464 -4652
rect 2568 -4852 2624 -4652
rect 2728 -4852 2784 -4652
rect 2888 -4852 2944 -4652
rect 3048 -4852 3104 -4652
rect 3208 -4852 3264 -4652
rect 3818 -4852 3874 -4652
rect 3978 -4852 4034 -4652
rect 4138 -4852 4194 -4652
rect 4298 -4852 4354 -4652
rect 4458 -4852 4514 -4652
rect 4618 -4852 4674 -4652
rect 5021 -4852 5077 -4652
rect 5685 -4853 5741 -4653
rect 6088 -4853 6144 -4653
rect 6248 -4853 6304 -4653
rect 6408 -4853 6464 -4653
rect 6568 -4853 6624 -4653
rect 6728 -4853 6784 -4653
rect 6888 -4853 6944 -4653
rect -4757 -5512 -4701 -5312
rect -4353 -5512 -4297 -5312
rect -3950 -5512 -3894 -5312
rect -3790 -5512 -3734 -5312
rect -3630 -5512 -3574 -5312
rect -3470 -5512 -3414 -5312
rect -3310 -5512 -3254 -5312
rect -3150 -5512 -3094 -5312
rect -2354 -5505 -2298 -5305
rect -1950 -5505 -1894 -5305
rect -1547 -5505 -1491 -5305
rect -1387 -5505 -1331 -5305
rect -1227 -5505 -1171 -5305
rect -1067 -5505 -1011 -5305
rect -907 -5505 -851 -5305
rect -747 -5505 -691 -5305
rect 245 -5504 301 -5304
rect 648 -5504 704 -5304
rect 808 -5504 864 -5304
rect 968 -5504 1024 -5304
rect 1128 -5504 1184 -5304
rect 1288 -5504 1344 -5304
rect 1448 -5504 1504 -5304
rect 2005 -5504 2061 -5304
rect 2165 -5504 2221 -5304
rect 2325 -5504 2381 -5304
rect 2485 -5504 2541 -5304
rect 2645 -5504 2701 -5304
rect 2805 -5504 2861 -5304
rect 3208 -5504 3264 -5304
rect 3818 -5504 3874 -5304
rect 4221 -5504 4277 -5304
rect 4381 -5504 4437 -5304
rect 4541 -5504 4597 -5304
rect 4701 -5504 4757 -5304
rect 4861 -5504 4917 -5304
rect 5021 -5504 5077 -5304
rect 5685 -5505 5741 -5305
rect 5845 -5505 5901 -5305
rect 6005 -5505 6061 -5305
rect 6165 -5505 6221 -5305
rect 6325 -5505 6381 -5305
rect 6485 -5505 6541 -5305
rect 6888 -5505 6944 -5305
rect -4757 -5848 -4701 -5648
rect -4353 -5848 -4297 -5648
rect -3950 -5848 -3894 -5648
rect -3790 -5848 -3734 -5648
rect -3630 -5848 -3574 -5648
rect -3470 -5848 -3414 -5648
rect -3310 -5848 -3254 -5648
rect -3150 -5848 -3094 -5648
rect -2354 -5841 -2298 -5641
rect -1950 -5841 -1894 -5641
rect -1547 -5841 -1491 -5641
rect -1387 -5841 -1331 -5641
rect -1227 -5841 -1171 -5641
rect -1067 -5841 -1011 -5641
rect -907 -5841 -851 -5641
rect -747 -5841 -691 -5641
rect 245 -5840 301 -5640
rect 648 -5840 704 -5640
rect 808 -5840 864 -5640
rect 968 -5840 1024 -5640
rect 1128 -5840 1184 -5640
rect 1288 -5840 1344 -5640
rect 1448 -5840 1504 -5640
rect 2005 -5840 2061 -5640
rect 2165 -5840 2221 -5640
rect 2325 -5840 2381 -5640
rect 2485 -5840 2541 -5640
rect 2645 -5840 2701 -5640
rect 2805 -5840 2861 -5640
rect 3208 -5840 3264 -5640
rect 3818 -5840 3874 -5640
rect 4221 -5840 4277 -5640
rect 4381 -5840 4437 -5640
rect 4541 -5840 4597 -5640
rect 4701 -5840 4757 -5640
rect 4861 -5840 4917 -5640
rect 5021 -5840 5077 -5640
rect 5685 -5841 5741 -5641
rect 5845 -5841 5901 -5641
rect 6005 -5841 6061 -5641
rect 6165 -5841 6221 -5641
rect 6325 -5841 6381 -5641
rect 6485 -5841 6541 -5641
rect 6888 -5841 6944 -5641
<< pmos >>
rect -4757 2226 -4701 2426
rect -4353 2226 -4297 2426
rect -3950 2226 -3894 2426
rect -3790 2226 -3734 2426
rect -3630 2226 -3574 2426
rect -3470 2226 -3414 2426
rect -3310 2226 -3254 2426
rect -3150 2226 -3094 2426
rect -2354 2233 -2298 2433
rect -1950 2233 -1894 2433
rect -1547 2233 -1491 2433
rect -1387 2233 -1331 2433
rect -1227 2233 -1171 2433
rect -1067 2233 -1011 2433
rect -907 2233 -851 2433
rect -747 2233 -691 2433
rect 245 2234 301 2434
rect 648 2234 704 2434
rect 808 2234 864 2434
rect 968 2234 1024 2434
rect 1128 2234 1184 2434
rect 1288 2234 1344 2434
rect 1448 2234 1504 2434
rect 2005 2234 2061 2434
rect 2165 2234 2221 2434
rect 2325 2234 2381 2434
rect 2485 2234 2541 2434
rect 2645 2234 2701 2434
rect 2805 2234 2861 2434
rect 3208 2234 3264 2434
rect 3818 2234 3874 2434
rect 4221 2234 4277 2434
rect 4381 2234 4437 2434
rect 4541 2234 4597 2434
rect 4701 2234 4757 2434
rect 4861 2234 4917 2434
rect 5021 2234 5077 2434
rect 5685 2233 5741 2433
rect 5845 2233 5901 2433
rect 6005 2233 6061 2433
rect 6165 2233 6221 2433
rect 6325 2233 6381 2433
rect 6485 2233 6541 2433
rect 6888 2233 6944 2433
rect -4757 1890 -4701 2090
rect -4353 1890 -4297 2090
rect -3950 1890 -3894 2090
rect -3790 1890 -3734 2090
rect -3630 1890 -3574 2090
rect -3470 1890 -3414 2090
rect -3310 1890 -3254 2090
rect -3150 1890 -3094 2090
rect -2354 1897 -2298 2097
rect -1950 1897 -1894 2097
rect -1547 1897 -1491 2097
rect -1387 1897 -1331 2097
rect -1227 1897 -1171 2097
rect -1067 1897 -1011 2097
rect -907 1897 -851 2097
rect -747 1897 -691 2097
rect 245 1898 301 2098
rect 648 1898 704 2098
rect 808 1898 864 2098
rect 968 1898 1024 2098
rect 1128 1898 1184 2098
rect 1288 1898 1344 2098
rect 1448 1898 1504 2098
rect 2005 1898 2061 2098
rect 2165 1898 2221 2098
rect 2325 1898 2381 2098
rect 2485 1898 2541 2098
rect 2645 1898 2701 2098
rect 2805 1898 2861 2098
rect 3208 1898 3264 2098
rect 3818 1898 3874 2098
rect 4221 1898 4277 2098
rect 4381 1898 4437 2098
rect 4541 1898 4597 2098
rect 4701 1898 4757 2098
rect 4861 1898 4917 2098
rect 5021 1898 5077 2098
rect 5685 1897 5741 2097
rect 5845 1897 5901 2097
rect 6005 1897 6061 2097
rect 6165 1897 6221 2097
rect 6325 1897 6381 2097
rect 6485 1897 6541 2097
rect 6888 1897 6944 2097
rect -4757 1554 -4701 1754
rect -4353 1554 -4297 1754
rect -3950 1554 -3894 1754
rect -3790 1554 -3734 1754
rect -3630 1554 -3574 1754
rect -3470 1554 -3414 1754
rect -3310 1554 -3254 1754
rect -3150 1554 -3094 1754
rect -2354 1561 -2298 1761
rect -1950 1561 -1894 1761
rect -1547 1561 -1491 1761
rect -1387 1561 -1331 1761
rect -1227 1561 -1171 1761
rect -1067 1561 -1011 1761
rect -907 1561 -851 1761
rect -747 1561 -691 1761
rect 245 1562 301 1762
rect 648 1562 704 1762
rect 808 1562 864 1762
rect 968 1562 1024 1762
rect 1128 1562 1184 1762
rect 1288 1562 1344 1762
rect 1448 1562 1504 1762
rect 2005 1562 2061 1762
rect 2165 1562 2221 1762
rect 2325 1562 2381 1762
rect 2485 1562 2541 1762
rect 2645 1562 2701 1762
rect 2805 1562 2861 1762
rect 3208 1562 3264 1762
rect 3818 1562 3874 1762
rect 4221 1562 4277 1762
rect 4381 1562 4437 1762
rect 4541 1562 4597 1762
rect 4701 1562 4757 1762
rect 4861 1562 4917 1762
rect 5021 1562 5077 1762
rect 5685 1561 5741 1761
rect 5845 1561 5901 1761
rect 6005 1561 6061 1761
rect 6165 1561 6221 1761
rect 6325 1561 6381 1761
rect 6485 1561 6541 1761
rect 6888 1561 6944 1761
rect -4757 1218 -4701 1418
rect -4353 1218 -4297 1418
rect -3950 1218 -3894 1418
rect -3790 1218 -3734 1418
rect -3630 1218 -3574 1418
rect -3470 1218 -3414 1418
rect -3310 1218 -3254 1418
rect -3150 1218 -3094 1418
rect -2354 1225 -2298 1425
rect -1950 1225 -1894 1425
rect -1547 1225 -1491 1425
rect -1387 1225 -1331 1425
rect -1227 1225 -1171 1425
rect -1067 1225 -1011 1425
rect -907 1225 -851 1425
rect -747 1225 -691 1425
rect 245 1226 301 1426
rect 648 1226 704 1426
rect 808 1226 864 1426
rect 968 1226 1024 1426
rect 1128 1226 1184 1426
rect 1288 1226 1344 1426
rect 1448 1226 1504 1426
rect 2005 1226 2061 1426
rect 2165 1226 2221 1426
rect 2325 1226 2381 1426
rect 2485 1226 2541 1426
rect 2645 1226 2701 1426
rect 2805 1226 2861 1426
rect 3208 1226 3264 1426
rect 3818 1226 3874 1426
rect 4221 1226 4277 1426
rect 4381 1226 4437 1426
rect 4541 1226 4597 1426
rect 4701 1226 4757 1426
rect 4861 1226 4917 1426
rect 5021 1226 5077 1426
rect 5685 1225 5741 1425
rect 5845 1225 5901 1425
rect 6005 1225 6061 1425
rect 6165 1225 6221 1425
rect 6325 1225 6381 1425
rect 6485 1225 6541 1425
rect 6888 1225 6944 1425
rect 235 -530 291 -330
rect 395 -530 451 -330
rect 555 -530 611 -330
rect 715 -530 771 -330
rect 235 -866 291 -666
rect 395 -866 451 -666
rect 555 -866 611 -666
rect 715 -866 771 -666
rect -4757 -1270 -4701 -1070
rect -4353 -1270 -4297 -1070
rect -3950 -1270 -3894 -1070
rect -3790 -1270 -3734 -1070
rect -3630 -1270 -3574 -1070
rect -3470 -1270 -3414 -1070
rect -3310 -1270 -3254 -1070
rect -3150 -1270 -3094 -1070
rect -2354 -1263 -2298 -1063
rect -1950 -1263 -1894 -1063
rect -1547 -1263 -1491 -1063
rect -1387 -1263 -1331 -1063
rect -1227 -1263 -1171 -1063
rect -1067 -1263 -1011 -1063
rect -907 -1263 -851 -1063
rect -747 -1263 -691 -1063
rect 2005 -1262 2061 -1062
rect 2408 -1262 2464 -1062
rect 2568 -1262 2624 -1062
rect 2728 -1262 2784 -1062
rect 2888 -1262 2944 -1062
rect 3048 -1262 3104 -1062
rect 3208 -1262 3264 -1062
rect 3818 -1262 3874 -1062
rect 3978 -1262 4034 -1062
rect 4138 -1262 4194 -1062
rect 4298 -1262 4354 -1062
rect 4458 -1262 4514 -1062
rect 4618 -1262 4674 -1062
rect 5021 -1262 5077 -1062
rect -4757 -1606 -4701 -1406
rect -4353 -1606 -4297 -1406
rect -3950 -1606 -3894 -1406
rect -3790 -1606 -3734 -1406
rect -3630 -1606 -3574 -1406
rect -3470 -1606 -3414 -1406
rect -3310 -1606 -3254 -1406
rect -3150 -1606 -3094 -1406
rect -2354 -1599 -2298 -1399
rect -1950 -1599 -1894 -1399
rect -1547 -1599 -1491 -1399
rect -1387 -1599 -1331 -1399
rect -1227 -1599 -1171 -1399
rect -1067 -1599 -1011 -1399
rect -907 -1599 -851 -1399
rect -747 -1599 -691 -1399
rect 5685 -1263 5741 -1063
rect 6088 -1263 6144 -1063
rect 6248 -1263 6304 -1063
rect 6408 -1263 6464 -1063
rect 6568 -1263 6624 -1063
rect 6728 -1263 6784 -1063
rect 6888 -1263 6944 -1063
rect 2005 -1598 2061 -1398
rect 2408 -1598 2464 -1398
rect 2568 -1598 2624 -1398
rect 2728 -1598 2784 -1398
rect 2888 -1598 2944 -1398
rect 3048 -1598 3104 -1398
rect 3208 -1598 3264 -1398
rect 3818 -1598 3874 -1398
rect 3978 -1598 4034 -1398
rect 4138 -1598 4194 -1398
rect 4298 -1598 4354 -1398
rect 4458 -1598 4514 -1398
rect 4618 -1598 4674 -1398
rect 5021 -1598 5077 -1398
rect -4757 -1942 -4701 -1742
rect -4353 -1942 -4297 -1742
rect -3950 -1942 -3894 -1742
rect -3790 -1942 -3734 -1742
rect -3630 -1942 -3574 -1742
rect -3470 -1942 -3414 -1742
rect -3310 -1942 -3254 -1742
rect -3150 -1942 -3094 -1742
rect -2354 -1935 -2298 -1735
rect -1950 -1935 -1894 -1735
rect -1547 -1935 -1491 -1735
rect -1387 -1935 -1331 -1735
rect -1227 -1935 -1171 -1735
rect -1067 -1935 -1011 -1735
rect -907 -1935 -851 -1735
rect -747 -1935 -691 -1735
rect 5685 -1599 5741 -1399
rect 6088 -1599 6144 -1399
rect 6248 -1599 6304 -1399
rect 6408 -1599 6464 -1399
rect 6568 -1599 6624 -1399
rect 6728 -1599 6784 -1399
rect 6888 -1599 6944 -1399
rect 2005 -1934 2061 -1734
rect 2408 -1934 2464 -1734
rect 2568 -1934 2624 -1734
rect 2728 -1934 2784 -1734
rect 2888 -1934 2944 -1734
rect 3048 -1934 3104 -1734
rect 3208 -1934 3264 -1734
rect 3818 -1934 3874 -1734
rect 3978 -1934 4034 -1734
rect 4138 -1934 4194 -1734
rect 4298 -1934 4354 -1734
rect 4458 -1934 4514 -1734
rect 4618 -1934 4674 -1734
rect 5021 -1934 5077 -1734
rect -4757 -2278 -4701 -2078
rect -4353 -2278 -4297 -2078
rect -3950 -2278 -3894 -2078
rect -3790 -2278 -3734 -2078
rect -3630 -2278 -3574 -2078
rect -3470 -2278 -3414 -2078
rect -3310 -2278 -3254 -2078
rect -3150 -2278 -3094 -2078
rect -2354 -2271 -2298 -2071
rect -1950 -2271 -1894 -2071
rect -1547 -2271 -1491 -2071
rect -1387 -2271 -1331 -2071
rect -1227 -2271 -1171 -2071
rect -1067 -2271 -1011 -2071
rect -907 -2271 -851 -2071
rect -747 -2271 -691 -2071
rect 5685 -1935 5741 -1735
rect 6088 -1935 6144 -1735
rect 6248 -1935 6304 -1735
rect 6408 -1935 6464 -1735
rect 6568 -1935 6624 -1735
rect 6728 -1935 6784 -1735
rect 6888 -1935 6944 -1735
rect 2005 -2270 2061 -2070
rect 2408 -2270 2464 -2070
rect 2568 -2270 2624 -2070
rect 2728 -2270 2784 -2070
rect 2888 -2270 2944 -2070
rect 3048 -2270 3104 -2070
rect 3208 -2270 3264 -2070
rect 3818 -2270 3874 -2070
rect 3978 -2270 4034 -2070
rect 4138 -2270 4194 -2070
rect 4298 -2270 4354 -2070
rect 4458 -2270 4514 -2070
rect 4618 -2270 4674 -2070
rect 5021 -2270 5077 -2070
rect 5685 -2271 5741 -2071
rect 6088 -2271 6144 -2071
rect 6248 -2271 6304 -2071
rect 6408 -2271 6464 -2071
rect 6568 -2271 6624 -2071
rect 6728 -2271 6784 -2071
rect 6888 -2271 6944 -2071
rect 235 -2541 291 -2341
rect 395 -2541 451 -2341
rect 555 -2541 611 -2341
rect 715 -2541 771 -2341
rect -4757 -2934 -4701 -2734
rect -4353 -2934 -4297 -2734
rect -3950 -2934 -3894 -2734
rect -3790 -2934 -3734 -2734
rect -3630 -2934 -3574 -2734
rect -3470 -2934 -3414 -2734
rect -3310 -2934 -3254 -2734
rect -3150 -2934 -3094 -2734
rect -2354 -2927 -2298 -2727
rect -1950 -2927 -1894 -2727
rect -1547 -2927 -1491 -2727
rect -1387 -2927 -1331 -2727
rect -1227 -2927 -1171 -2727
rect -1067 -2927 -1011 -2727
rect -907 -2927 -851 -2727
rect -747 -2927 -691 -2727
rect 235 -2877 291 -2677
rect 395 -2877 451 -2677
rect 555 -2877 611 -2677
rect 715 -2877 771 -2677
rect 2005 -2926 2061 -2726
rect 2408 -2926 2464 -2726
rect 2568 -2926 2624 -2726
rect 2728 -2926 2784 -2726
rect 2888 -2926 2944 -2726
rect 3048 -2926 3104 -2726
rect 3208 -2926 3264 -2726
rect 3818 -2926 3874 -2726
rect 3978 -2926 4034 -2726
rect 4138 -2926 4194 -2726
rect 4298 -2926 4354 -2726
rect 4458 -2926 4514 -2726
rect 4618 -2926 4674 -2726
rect 5021 -2926 5077 -2726
rect -4757 -3270 -4701 -3070
rect -4353 -3270 -4297 -3070
rect -3950 -3270 -3894 -3070
rect -3790 -3270 -3734 -3070
rect -3630 -3270 -3574 -3070
rect -3470 -3270 -3414 -3070
rect -3310 -3270 -3254 -3070
rect -3150 -3270 -3094 -3070
rect -2354 -3263 -2298 -3063
rect -1950 -3263 -1894 -3063
rect -1547 -3263 -1491 -3063
rect -1387 -3263 -1331 -3063
rect -1227 -3263 -1171 -3063
rect -1067 -3263 -1011 -3063
rect -907 -3263 -851 -3063
rect -747 -3263 -691 -3063
rect 5685 -2927 5741 -2727
rect 6088 -2927 6144 -2727
rect 6248 -2927 6304 -2727
rect 6408 -2927 6464 -2727
rect 6568 -2927 6624 -2727
rect 6728 -2927 6784 -2727
rect 6888 -2927 6944 -2727
rect 2005 -3262 2061 -3062
rect 2408 -3262 2464 -3062
rect 2568 -3262 2624 -3062
rect 2728 -3262 2784 -3062
rect 2888 -3262 2944 -3062
rect 3048 -3262 3104 -3062
rect 3208 -3262 3264 -3062
rect 3818 -3262 3874 -3062
rect 3978 -3262 4034 -3062
rect 4138 -3262 4194 -3062
rect 4298 -3262 4354 -3062
rect 4458 -3262 4514 -3062
rect 4618 -3262 4674 -3062
rect 5021 -3262 5077 -3062
rect -4757 -3606 -4701 -3406
rect -4353 -3606 -4297 -3406
rect -3950 -3606 -3894 -3406
rect -3790 -3606 -3734 -3406
rect -3630 -3606 -3574 -3406
rect -3470 -3606 -3414 -3406
rect -3310 -3606 -3254 -3406
rect -3150 -3606 -3094 -3406
rect -2354 -3599 -2298 -3399
rect -1950 -3599 -1894 -3399
rect -1547 -3599 -1491 -3399
rect -1387 -3599 -1331 -3399
rect -1227 -3599 -1171 -3399
rect -1067 -3599 -1011 -3399
rect -907 -3599 -851 -3399
rect -747 -3599 -691 -3399
rect 235 -3471 291 -3271
rect 395 -3471 451 -3271
rect 555 -3471 611 -3271
rect 715 -3471 771 -3271
rect 5685 -3263 5741 -3063
rect 6088 -3263 6144 -3063
rect 6248 -3263 6304 -3063
rect 6408 -3263 6464 -3063
rect 6568 -3263 6624 -3063
rect 6728 -3263 6784 -3063
rect 6888 -3263 6944 -3063
rect 2005 -3598 2061 -3398
rect 2408 -3598 2464 -3398
rect 2568 -3598 2624 -3398
rect 2728 -3598 2784 -3398
rect 2888 -3598 2944 -3398
rect 3048 -3598 3104 -3398
rect 3208 -3598 3264 -3398
rect 3818 -3598 3874 -3398
rect 3978 -3598 4034 -3398
rect 4138 -3598 4194 -3398
rect 4298 -3598 4354 -3398
rect 4458 -3598 4514 -3398
rect 4618 -3598 4674 -3398
rect 5021 -3598 5077 -3398
rect -4757 -3942 -4701 -3742
rect -4353 -3942 -4297 -3742
rect -3950 -3942 -3894 -3742
rect -3790 -3942 -3734 -3742
rect -3630 -3942 -3574 -3742
rect -3470 -3942 -3414 -3742
rect -3310 -3942 -3254 -3742
rect -3150 -3942 -3094 -3742
rect -2354 -3935 -2298 -3735
rect -1950 -3935 -1894 -3735
rect -1547 -3935 -1491 -3735
rect -1387 -3935 -1331 -3735
rect -1227 -3935 -1171 -3735
rect -1067 -3935 -1011 -3735
rect -907 -3935 -851 -3735
rect -747 -3935 -691 -3735
rect 235 -3807 291 -3607
rect 395 -3807 451 -3607
rect 555 -3807 611 -3607
rect 715 -3807 771 -3607
rect 5685 -3599 5741 -3399
rect 6088 -3599 6144 -3399
rect 6248 -3599 6304 -3399
rect 6408 -3599 6464 -3399
rect 6568 -3599 6624 -3399
rect 6728 -3599 6784 -3399
rect 6888 -3599 6944 -3399
rect 2005 -3934 2061 -3734
rect 2408 -3934 2464 -3734
rect 2568 -3934 2624 -3734
rect 2728 -3934 2784 -3734
rect 2888 -3934 2944 -3734
rect 3048 -3934 3104 -3734
rect 3208 -3934 3264 -3734
rect 3818 -3934 3874 -3734
rect 3978 -3934 4034 -3734
rect 4138 -3934 4194 -3734
rect 4298 -3934 4354 -3734
rect 4458 -3934 4514 -3734
rect 4618 -3934 4674 -3734
rect 5021 -3934 5077 -3734
rect 5685 -3935 5741 -3735
rect 6088 -3935 6144 -3735
rect 6248 -3935 6304 -3735
rect 6408 -3935 6464 -3735
rect 6568 -3935 6624 -3735
rect 6728 -3935 6784 -3735
rect 6888 -3935 6944 -3735
rect -4757 -6430 -4701 -6230
rect -4353 -6430 -4297 -6230
rect -3950 -6430 -3894 -6230
rect -3790 -6430 -3734 -6230
rect -3630 -6430 -3574 -6230
rect -3470 -6430 -3414 -6230
rect -3310 -6430 -3254 -6230
rect -3150 -6430 -3094 -6230
rect -2354 -6423 -2298 -6223
rect -1950 -6423 -1894 -6223
rect -1547 -6423 -1491 -6223
rect -1387 -6423 -1331 -6223
rect -1227 -6423 -1171 -6223
rect -1067 -6423 -1011 -6223
rect -907 -6423 -851 -6223
rect -747 -6423 -691 -6223
rect 245 -6422 301 -6222
rect 648 -6422 704 -6222
rect 808 -6422 864 -6222
rect 968 -6422 1024 -6222
rect 1128 -6422 1184 -6222
rect 1288 -6422 1344 -6222
rect 1448 -6422 1504 -6222
rect 2005 -6422 2061 -6222
rect 2165 -6422 2221 -6222
rect 2325 -6422 2381 -6222
rect 2485 -6422 2541 -6222
rect 2645 -6422 2701 -6222
rect 2805 -6422 2861 -6222
rect 3208 -6422 3264 -6222
rect 3818 -6422 3874 -6222
rect 4221 -6422 4277 -6222
rect 4381 -6422 4437 -6222
rect 4541 -6422 4597 -6222
rect 4701 -6422 4757 -6222
rect 4861 -6422 4917 -6222
rect 5021 -6422 5077 -6222
rect 5685 -6423 5741 -6223
rect 5845 -6423 5901 -6223
rect 6005 -6423 6061 -6223
rect 6165 -6423 6221 -6223
rect 6325 -6423 6381 -6223
rect 6485 -6423 6541 -6223
rect 6888 -6423 6944 -6223
rect -4757 -6766 -4701 -6566
rect -4353 -6766 -4297 -6566
rect -3950 -6766 -3894 -6566
rect -3790 -6766 -3734 -6566
rect -3630 -6766 -3574 -6566
rect -3470 -6766 -3414 -6566
rect -3310 -6766 -3254 -6566
rect -3150 -6766 -3094 -6566
rect -2354 -6759 -2298 -6559
rect -1950 -6759 -1894 -6559
rect -1547 -6759 -1491 -6559
rect -1387 -6759 -1331 -6559
rect -1227 -6759 -1171 -6559
rect -1067 -6759 -1011 -6559
rect -907 -6759 -851 -6559
rect -747 -6759 -691 -6559
rect 245 -6758 301 -6558
rect 648 -6758 704 -6558
rect 808 -6758 864 -6558
rect 968 -6758 1024 -6558
rect 1128 -6758 1184 -6558
rect 1288 -6758 1344 -6558
rect 1448 -6758 1504 -6558
rect 2005 -6758 2061 -6558
rect 2165 -6758 2221 -6558
rect 2325 -6758 2381 -6558
rect 2485 -6758 2541 -6558
rect 2645 -6758 2701 -6558
rect 2805 -6758 2861 -6558
rect 3208 -6758 3264 -6558
rect 3818 -6758 3874 -6558
rect 4221 -6758 4277 -6558
rect 4381 -6758 4437 -6558
rect 4541 -6758 4597 -6558
rect 4701 -6758 4757 -6558
rect 4861 -6758 4917 -6558
rect 5021 -6758 5077 -6558
rect 5685 -6759 5741 -6559
rect 5845 -6759 5901 -6559
rect 6005 -6759 6061 -6559
rect 6165 -6759 6221 -6559
rect 6325 -6759 6381 -6559
rect 6485 -6759 6541 -6559
rect 6888 -6759 6944 -6559
rect -4757 -7102 -4701 -6902
rect -4353 -7102 -4297 -6902
rect -3950 -7102 -3894 -6902
rect -3790 -7102 -3734 -6902
rect -3630 -7102 -3574 -6902
rect -3470 -7102 -3414 -6902
rect -3310 -7102 -3254 -6902
rect -3150 -7102 -3094 -6902
rect -2354 -7095 -2298 -6895
rect -1950 -7095 -1894 -6895
rect -1547 -7095 -1491 -6895
rect -1387 -7095 -1331 -6895
rect -1227 -7095 -1171 -6895
rect -1067 -7095 -1011 -6895
rect -907 -7095 -851 -6895
rect -747 -7095 -691 -6895
rect 245 -7094 301 -6894
rect 648 -7094 704 -6894
rect 808 -7094 864 -6894
rect 968 -7094 1024 -6894
rect 1128 -7094 1184 -6894
rect 1288 -7094 1344 -6894
rect 1448 -7094 1504 -6894
rect 2005 -7094 2061 -6894
rect 2165 -7094 2221 -6894
rect 2325 -7094 2381 -6894
rect 2485 -7094 2541 -6894
rect 2645 -7094 2701 -6894
rect 2805 -7094 2861 -6894
rect 3208 -7094 3264 -6894
rect 3818 -7094 3874 -6894
rect 4221 -7094 4277 -6894
rect 4381 -7094 4437 -6894
rect 4541 -7094 4597 -6894
rect 4701 -7094 4757 -6894
rect 4861 -7094 4917 -6894
rect 5021 -7094 5077 -6894
rect 5685 -7095 5741 -6895
rect 5845 -7095 5901 -6895
rect 6005 -7095 6061 -6895
rect 6165 -7095 6221 -6895
rect 6325 -7095 6381 -6895
rect 6485 -7095 6541 -6895
rect 6888 -7095 6944 -6895
rect -4757 -7438 -4701 -7238
rect -4353 -7438 -4297 -7238
rect -3950 -7438 -3894 -7238
rect -3790 -7438 -3734 -7238
rect -3630 -7438 -3574 -7238
rect -3470 -7438 -3414 -7238
rect -3310 -7438 -3254 -7238
rect -3150 -7438 -3094 -7238
rect -2354 -7431 -2298 -7231
rect -1950 -7431 -1894 -7231
rect -1547 -7431 -1491 -7231
rect -1387 -7431 -1331 -7231
rect -1227 -7431 -1171 -7231
rect -1067 -7431 -1011 -7231
rect -907 -7431 -851 -7231
rect -747 -7431 -691 -7231
rect 245 -7430 301 -7230
rect 648 -7430 704 -7230
rect 808 -7430 864 -7230
rect 968 -7430 1024 -7230
rect 1128 -7430 1184 -7230
rect 1288 -7430 1344 -7230
rect 1448 -7430 1504 -7230
rect 2005 -7430 2061 -7230
rect 2165 -7430 2221 -7230
rect 2325 -7430 2381 -7230
rect 2485 -7430 2541 -7230
rect 2645 -7430 2701 -7230
rect 2805 -7430 2861 -7230
rect 3208 -7430 3264 -7230
rect 3818 -7430 3874 -7230
rect 4221 -7430 4277 -7230
rect 4381 -7430 4437 -7230
rect 4541 -7430 4597 -7230
rect 4701 -7430 4757 -7230
rect 4861 -7430 4917 -7230
rect 5021 -7430 5077 -7230
rect 5685 -7431 5741 -7231
rect 5845 -7431 5901 -7231
rect 6005 -7431 6061 -7231
rect 6165 -7431 6221 -7231
rect 6325 -7431 6381 -7231
rect 6485 -7431 6541 -7231
rect 6888 -7431 6944 -7231
<< ndiff >>
rect -4845 823 -4757 836
rect -4845 649 -4832 823
rect -4786 649 -4757 823
rect -4845 636 -4757 649
rect -4701 823 -4613 836
rect -4701 649 -4672 823
rect -4626 649 -4613 823
rect -4701 636 -4613 649
rect -4441 823 -4353 836
rect -4441 649 -4428 823
rect -4382 649 -4353 823
rect -4441 636 -4353 649
rect -4297 823 -4209 836
rect -4297 649 -4268 823
rect -4222 649 -4209 823
rect -4297 636 -4209 649
rect -4038 823 -3950 836
rect -4038 649 -4025 823
rect -3979 649 -3950 823
rect -4038 636 -3950 649
rect -3894 823 -3790 836
rect -3894 649 -3865 823
rect -3819 649 -3790 823
rect -3894 636 -3790 649
rect -3734 823 -3630 836
rect -3734 649 -3705 823
rect -3659 649 -3630 823
rect -3734 636 -3630 649
rect -3574 823 -3470 836
rect -3574 649 -3545 823
rect -3499 649 -3470 823
rect -3574 636 -3470 649
rect -3414 823 -3310 836
rect -3414 649 -3385 823
rect -3339 649 -3310 823
rect -3414 636 -3310 649
rect -3254 823 -3150 836
rect -3254 649 -3225 823
rect -3179 649 -3150 823
rect -3254 636 -3150 649
rect -3094 823 -3006 836
rect -3094 649 -3065 823
rect -3019 649 -3006 823
rect -3094 636 -3006 649
rect -2442 830 -2354 843
rect -2442 656 -2429 830
rect -2383 656 -2354 830
rect -2442 643 -2354 656
rect -2298 830 -2210 843
rect -2298 656 -2269 830
rect -2223 656 -2210 830
rect -2298 643 -2210 656
rect -2038 830 -1950 843
rect -2038 656 -2025 830
rect -1979 656 -1950 830
rect -2038 643 -1950 656
rect -1894 830 -1806 843
rect -1894 656 -1865 830
rect -1819 656 -1806 830
rect -1894 643 -1806 656
rect -1635 830 -1547 843
rect -1635 656 -1622 830
rect -1576 656 -1547 830
rect -1635 643 -1547 656
rect -1491 830 -1387 843
rect -1491 656 -1462 830
rect -1416 656 -1387 830
rect -1491 643 -1387 656
rect -1331 830 -1227 843
rect -1331 656 -1302 830
rect -1256 656 -1227 830
rect -1331 643 -1227 656
rect -1171 830 -1067 843
rect -1171 656 -1142 830
rect -1096 656 -1067 830
rect -1171 643 -1067 656
rect -1011 830 -907 843
rect -1011 656 -982 830
rect -936 656 -907 830
rect -1011 643 -907 656
rect -851 830 -747 843
rect -851 656 -822 830
rect -776 656 -747 830
rect -851 643 -747 656
rect -691 830 -603 843
rect -691 656 -662 830
rect -616 656 -603 830
rect -691 643 -603 656
rect 157 831 245 844
rect 157 657 170 831
rect 216 657 245 831
rect 157 644 245 657
rect 301 831 389 844
rect 301 657 330 831
rect 376 657 389 831
rect 301 644 389 657
rect 560 831 648 844
rect 560 657 573 831
rect 619 657 648 831
rect 560 644 648 657
rect 704 831 808 844
rect 704 657 733 831
rect 779 657 808 831
rect 704 644 808 657
rect 864 831 968 844
rect 864 657 893 831
rect 939 657 968 831
rect 864 644 968 657
rect 1024 831 1128 844
rect 1024 657 1053 831
rect 1099 657 1128 831
rect 1024 644 1128 657
rect 1184 831 1288 844
rect 1184 657 1213 831
rect 1259 657 1288 831
rect 1184 644 1288 657
rect 1344 831 1448 844
rect 1344 657 1373 831
rect 1419 657 1448 831
rect 1344 644 1448 657
rect 1504 831 1592 844
rect 1504 657 1533 831
rect 1579 657 1592 831
rect 1504 644 1592 657
rect 1917 831 2005 844
rect 1917 657 1930 831
rect 1976 657 2005 831
rect 1917 644 2005 657
rect 2061 831 2165 844
rect 2061 657 2090 831
rect 2136 657 2165 831
rect 2061 644 2165 657
rect 2221 831 2325 844
rect 2221 657 2250 831
rect 2296 657 2325 831
rect 2221 644 2325 657
rect 2381 831 2485 844
rect 2381 657 2410 831
rect 2456 657 2485 831
rect 2381 644 2485 657
rect 2541 831 2645 844
rect 2541 657 2570 831
rect 2616 657 2645 831
rect 2541 644 2645 657
rect 2701 831 2805 844
rect 2701 657 2730 831
rect 2776 657 2805 831
rect 2701 644 2805 657
rect 2861 831 2949 844
rect 2861 657 2890 831
rect 2936 657 2949 831
rect 2861 644 2949 657
rect 3120 831 3208 844
rect 3120 657 3133 831
rect 3179 657 3208 831
rect 3120 644 3208 657
rect 3264 831 3352 844
rect 3264 657 3293 831
rect 3339 657 3352 831
rect 3264 644 3352 657
rect 3730 831 3818 844
rect 3730 657 3743 831
rect 3789 657 3818 831
rect 3730 644 3818 657
rect 3874 831 3962 844
rect 3874 657 3903 831
rect 3949 657 3962 831
rect 3874 644 3962 657
rect 4133 831 4221 844
rect 4133 657 4146 831
rect 4192 657 4221 831
rect 4133 644 4221 657
rect 4277 831 4381 844
rect 4277 657 4306 831
rect 4352 657 4381 831
rect 4277 644 4381 657
rect 4437 831 4541 844
rect 4437 657 4466 831
rect 4512 657 4541 831
rect 4437 644 4541 657
rect 4597 831 4701 844
rect 4597 657 4626 831
rect 4672 657 4701 831
rect 4597 644 4701 657
rect 4757 831 4861 844
rect 4757 657 4786 831
rect 4832 657 4861 831
rect 4757 644 4861 657
rect 4917 831 5021 844
rect 4917 657 4946 831
rect 4992 657 5021 831
rect 4917 644 5021 657
rect 5077 831 5165 844
rect 5077 657 5106 831
rect 5152 657 5165 831
rect 5077 644 5165 657
rect 5597 830 5685 843
rect 5597 656 5610 830
rect 5656 656 5685 830
rect 5597 643 5685 656
rect 5741 830 5845 843
rect 5741 656 5770 830
rect 5816 656 5845 830
rect 5741 643 5845 656
rect 5901 830 6005 843
rect 5901 656 5930 830
rect 5976 656 6005 830
rect 5901 643 6005 656
rect 6061 830 6165 843
rect 6061 656 6090 830
rect 6136 656 6165 830
rect 6061 643 6165 656
rect 6221 830 6325 843
rect 6221 656 6250 830
rect 6296 656 6325 830
rect 6221 643 6325 656
rect 6381 830 6485 843
rect 6381 656 6410 830
rect 6456 656 6485 830
rect 6381 643 6485 656
rect 6541 830 6629 843
rect 6541 656 6570 830
rect 6616 656 6629 830
rect 6541 643 6629 656
rect 6800 830 6888 843
rect 6800 656 6813 830
rect 6859 656 6888 830
rect 6800 643 6888 656
rect 6944 830 7032 843
rect 6944 656 6973 830
rect 7019 656 7032 830
rect 6944 643 7032 656
rect -4845 487 -4757 500
rect -4845 313 -4832 487
rect -4786 313 -4757 487
rect -4845 300 -4757 313
rect -4701 487 -4613 500
rect -4701 313 -4672 487
rect -4626 313 -4613 487
rect -4701 300 -4613 313
rect -4441 487 -4353 500
rect -4441 313 -4428 487
rect -4382 313 -4353 487
rect -4441 300 -4353 313
rect -4297 487 -4209 500
rect -4297 313 -4268 487
rect -4222 313 -4209 487
rect -4297 300 -4209 313
rect -4038 487 -3950 500
rect -4038 313 -4025 487
rect -3979 313 -3950 487
rect -4038 300 -3950 313
rect -3894 487 -3790 500
rect -3894 313 -3865 487
rect -3819 313 -3790 487
rect -3894 300 -3790 313
rect -3734 487 -3630 500
rect -3734 313 -3705 487
rect -3659 313 -3630 487
rect -3734 300 -3630 313
rect -3574 487 -3470 500
rect -3574 313 -3545 487
rect -3499 313 -3470 487
rect -3574 300 -3470 313
rect -3414 487 -3310 500
rect -3414 313 -3385 487
rect -3339 313 -3310 487
rect -3414 300 -3310 313
rect -3254 487 -3150 500
rect -3254 313 -3225 487
rect -3179 313 -3150 487
rect -3254 300 -3150 313
rect -3094 487 -3006 500
rect -3094 313 -3065 487
rect -3019 313 -3006 487
rect -3094 300 -3006 313
rect -2442 494 -2354 507
rect -2442 320 -2429 494
rect -2383 320 -2354 494
rect -2442 307 -2354 320
rect -2298 494 -2210 507
rect -2298 320 -2269 494
rect -2223 320 -2210 494
rect -2298 307 -2210 320
rect -2038 494 -1950 507
rect -2038 320 -2025 494
rect -1979 320 -1950 494
rect -2038 307 -1950 320
rect -1894 494 -1806 507
rect -1894 320 -1865 494
rect -1819 320 -1806 494
rect -1894 307 -1806 320
rect -1635 494 -1547 507
rect -1635 320 -1622 494
rect -1576 320 -1547 494
rect -1635 307 -1547 320
rect -1491 494 -1387 507
rect -1491 320 -1462 494
rect -1416 320 -1387 494
rect -1491 307 -1387 320
rect -1331 494 -1227 507
rect -1331 320 -1302 494
rect -1256 320 -1227 494
rect -1331 307 -1227 320
rect -1171 494 -1067 507
rect -1171 320 -1142 494
rect -1096 320 -1067 494
rect -1171 307 -1067 320
rect -1011 494 -907 507
rect -1011 320 -982 494
rect -936 320 -907 494
rect -1011 307 -907 320
rect -851 494 -747 507
rect -851 320 -822 494
rect -776 320 -747 494
rect -851 307 -747 320
rect -691 494 -603 507
rect -691 320 -662 494
rect -616 320 -603 494
rect -691 307 -603 320
rect 157 495 245 508
rect 157 321 170 495
rect 216 321 245 495
rect 157 308 245 321
rect 301 495 389 508
rect 301 321 330 495
rect 376 321 389 495
rect 301 308 389 321
rect 560 495 648 508
rect 560 321 573 495
rect 619 321 648 495
rect 560 308 648 321
rect 704 495 808 508
rect 704 321 733 495
rect 779 321 808 495
rect 704 308 808 321
rect 864 495 968 508
rect 864 321 893 495
rect 939 321 968 495
rect 864 308 968 321
rect 1024 495 1128 508
rect 1024 321 1053 495
rect 1099 321 1128 495
rect 1024 308 1128 321
rect 1184 495 1288 508
rect 1184 321 1213 495
rect 1259 321 1288 495
rect 1184 308 1288 321
rect 1344 495 1448 508
rect 1344 321 1373 495
rect 1419 321 1448 495
rect 1344 308 1448 321
rect 1504 495 1592 508
rect 1504 321 1533 495
rect 1579 321 1592 495
rect 1504 308 1592 321
rect 1917 495 2005 508
rect 1917 321 1930 495
rect 1976 321 2005 495
rect 1917 308 2005 321
rect 2061 495 2165 508
rect 2061 321 2090 495
rect 2136 321 2165 495
rect 2061 308 2165 321
rect 2221 495 2325 508
rect 2221 321 2250 495
rect 2296 321 2325 495
rect 2221 308 2325 321
rect 2381 495 2485 508
rect 2381 321 2410 495
rect 2456 321 2485 495
rect 2381 308 2485 321
rect 2541 495 2645 508
rect 2541 321 2570 495
rect 2616 321 2645 495
rect 2541 308 2645 321
rect 2701 495 2805 508
rect 2701 321 2730 495
rect 2776 321 2805 495
rect 2701 308 2805 321
rect 2861 495 2949 508
rect 2861 321 2890 495
rect 2936 321 2949 495
rect 2861 308 2949 321
rect 3120 495 3208 508
rect 3120 321 3133 495
rect 3179 321 3208 495
rect 3120 308 3208 321
rect 3264 495 3352 508
rect 3264 321 3293 495
rect 3339 321 3352 495
rect 3264 308 3352 321
rect 3730 495 3818 508
rect 3730 321 3743 495
rect 3789 321 3818 495
rect 3730 308 3818 321
rect 3874 495 3962 508
rect 3874 321 3903 495
rect 3949 321 3962 495
rect 3874 308 3962 321
rect 4133 495 4221 508
rect 4133 321 4146 495
rect 4192 321 4221 495
rect 4133 308 4221 321
rect 4277 495 4381 508
rect 4277 321 4306 495
rect 4352 321 4381 495
rect 4277 308 4381 321
rect 4437 495 4541 508
rect 4437 321 4466 495
rect 4512 321 4541 495
rect 4437 308 4541 321
rect 4597 495 4701 508
rect 4597 321 4626 495
rect 4672 321 4701 495
rect 4597 308 4701 321
rect 4757 495 4861 508
rect 4757 321 4786 495
rect 4832 321 4861 495
rect 4757 308 4861 321
rect 4917 495 5021 508
rect 4917 321 4946 495
rect 4992 321 5021 495
rect 4917 308 5021 321
rect 5077 495 5165 508
rect 5077 321 5106 495
rect 5152 321 5165 495
rect 5077 308 5165 321
rect 5597 494 5685 507
rect 5597 320 5610 494
rect 5656 320 5685 494
rect 5597 307 5685 320
rect 5741 494 5845 507
rect 5741 320 5770 494
rect 5816 320 5845 494
rect 5741 307 5845 320
rect 5901 494 6005 507
rect 5901 320 5930 494
rect 5976 320 6005 494
rect 5901 307 6005 320
rect 6061 494 6165 507
rect 6061 320 6090 494
rect 6136 320 6165 494
rect 6061 307 6165 320
rect 6221 494 6325 507
rect 6221 320 6250 494
rect 6296 320 6325 494
rect 6221 307 6325 320
rect 6381 494 6485 507
rect 6381 320 6410 494
rect 6456 320 6485 494
rect 6381 307 6485 320
rect 6541 494 6629 507
rect 6541 320 6570 494
rect 6616 320 6629 494
rect 6541 307 6629 320
rect 6800 494 6888 507
rect 6800 320 6813 494
rect 6859 320 6888 494
rect 6800 307 6888 320
rect 6944 494 7032 507
rect 6944 320 6973 494
rect 7019 320 7032 494
rect 6944 307 7032 320
rect -4845 -165 -4757 -152
rect -4845 -339 -4832 -165
rect -4786 -339 -4757 -165
rect -4845 -352 -4757 -339
rect -4701 -165 -4613 -152
rect -4701 -339 -4672 -165
rect -4626 -339 -4613 -165
rect -4701 -352 -4613 -339
rect -4441 -165 -4353 -152
rect -4441 -339 -4428 -165
rect -4382 -339 -4353 -165
rect -4441 -352 -4353 -339
rect -4297 -165 -4209 -152
rect -4297 -339 -4268 -165
rect -4222 -339 -4209 -165
rect -4297 -352 -4209 -339
rect -4038 -165 -3950 -152
rect -4038 -339 -4025 -165
rect -3979 -339 -3950 -165
rect -4038 -352 -3950 -339
rect -3894 -165 -3790 -152
rect -3894 -339 -3865 -165
rect -3819 -339 -3790 -165
rect -3894 -352 -3790 -339
rect -3734 -165 -3630 -152
rect -3734 -339 -3705 -165
rect -3659 -339 -3630 -165
rect -3734 -352 -3630 -339
rect -3574 -165 -3470 -152
rect -3574 -339 -3545 -165
rect -3499 -339 -3470 -165
rect -3574 -352 -3470 -339
rect -3414 -165 -3310 -152
rect -3414 -339 -3385 -165
rect -3339 -339 -3310 -165
rect -3414 -352 -3310 -339
rect -3254 -165 -3150 -152
rect -3254 -339 -3225 -165
rect -3179 -339 -3150 -165
rect -3254 -352 -3150 -339
rect -3094 -165 -3006 -152
rect -3094 -339 -3065 -165
rect -3019 -339 -3006 -165
rect -3094 -352 -3006 -339
rect -2442 -158 -2354 -145
rect -2442 -332 -2429 -158
rect -2383 -332 -2354 -158
rect -2442 -345 -2354 -332
rect -2298 -158 -2210 -145
rect -2298 -332 -2269 -158
rect -2223 -332 -2210 -158
rect -2298 -345 -2210 -332
rect -2038 -158 -1950 -145
rect -2038 -332 -2025 -158
rect -1979 -332 -1950 -158
rect -2038 -345 -1950 -332
rect -1894 -158 -1806 -145
rect -1894 -332 -1865 -158
rect -1819 -332 -1806 -158
rect -1894 -345 -1806 -332
rect -1635 -158 -1547 -145
rect -1635 -332 -1622 -158
rect -1576 -332 -1547 -158
rect -1635 -345 -1547 -332
rect -1491 -158 -1387 -145
rect -1491 -332 -1462 -158
rect -1416 -332 -1387 -158
rect -1491 -345 -1387 -332
rect -1331 -158 -1227 -145
rect -1331 -332 -1302 -158
rect -1256 -332 -1227 -158
rect -1331 -345 -1227 -332
rect -1171 -158 -1067 -145
rect -1171 -332 -1142 -158
rect -1096 -332 -1067 -158
rect -1171 -345 -1067 -332
rect -1011 -158 -907 -145
rect -1011 -332 -982 -158
rect -936 -332 -907 -158
rect -1011 -345 -907 -332
rect -851 -158 -747 -145
rect -851 -332 -822 -158
rect -776 -332 -747 -158
rect -851 -345 -747 -332
rect -691 -158 -603 -145
rect -691 -332 -662 -158
rect -616 -332 -603 -158
rect 1917 -157 2005 -144
rect -691 -345 -603 -332
rect -4845 -501 -4757 -488
rect -4845 -675 -4832 -501
rect -4786 -675 -4757 -501
rect -4845 -688 -4757 -675
rect -4701 -501 -4613 -488
rect -4701 -675 -4672 -501
rect -4626 -675 -4613 -501
rect -4701 -688 -4613 -675
rect -4441 -501 -4353 -488
rect -4441 -675 -4428 -501
rect -4382 -675 -4353 -501
rect -4441 -688 -4353 -675
rect -4297 -501 -4209 -488
rect -4297 -675 -4268 -501
rect -4222 -675 -4209 -501
rect -4297 -688 -4209 -675
rect -4038 -501 -3950 -488
rect -4038 -675 -4025 -501
rect -3979 -675 -3950 -501
rect -4038 -688 -3950 -675
rect -3894 -501 -3790 -488
rect -3894 -675 -3865 -501
rect -3819 -675 -3790 -501
rect -3894 -688 -3790 -675
rect -3734 -501 -3630 -488
rect -3734 -675 -3705 -501
rect -3659 -675 -3630 -501
rect -3734 -688 -3630 -675
rect -3574 -501 -3470 -488
rect -3574 -675 -3545 -501
rect -3499 -675 -3470 -501
rect -3574 -688 -3470 -675
rect -3414 -501 -3310 -488
rect -3414 -675 -3385 -501
rect -3339 -675 -3310 -501
rect -3414 -688 -3310 -675
rect -3254 -501 -3150 -488
rect -3254 -675 -3225 -501
rect -3179 -675 -3150 -501
rect -3254 -688 -3150 -675
rect -3094 -501 -3006 -488
rect -3094 -675 -3065 -501
rect -3019 -675 -3006 -501
rect -3094 -688 -3006 -675
rect -2442 -494 -2354 -481
rect -2442 -668 -2429 -494
rect -2383 -668 -2354 -494
rect -2442 -681 -2354 -668
rect -2298 -494 -2210 -481
rect -2298 -668 -2269 -494
rect -2223 -668 -2210 -494
rect -2298 -681 -2210 -668
rect -2038 -494 -1950 -481
rect -2038 -668 -2025 -494
rect -1979 -668 -1950 -494
rect -2038 -681 -1950 -668
rect -1894 -494 -1806 -481
rect -1894 -668 -1865 -494
rect -1819 -668 -1806 -494
rect -1894 -681 -1806 -668
rect -1635 -494 -1547 -481
rect -1635 -668 -1622 -494
rect -1576 -668 -1547 -494
rect -1635 -681 -1547 -668
rect -1491 -494 -1387 -481
rect -1491 -668 -1462 -494
rect -1416 -668 -1387 -494
rect -1491 -681 -1387 -668
rect -1331 -494 -1227 -481
rect -1331 -668 -1302 -494
rect -1256 -668 -1227 -494
rect -1331 -681 -1227 -668
rect -1171 -494 -1067 -481
rect -1171 -668 -1142 -494
rect -1096 -668 -1067 -494
rect -1171 -681 -1067 -668
rect -1011 -494 -907 -481
rect -1011 -668 -982 -494
rect -936 -668 -907 -494
rect -1011 -681 -907 -668
rect -851 -494 -747 -481
rect -851 -668 -822 -494
rect -776 -668 -747 -494
rect -851 -681 -747 -668
rect -691 -494 -603 -481
rect -691 -668 -662 -494
rect -616 -668 -603 -494
rect 1917 -331 1930 -157
rect 1976 -331 2005 -157
rect 1917 -344 2005 -331
rect 2061 -157 2149 -144
rect 2061 -331 2090 -157
rect 2136 -331 2149 -157
rect 2061 -344 2149 -331
rect 2320 -157 2408 -144
rect 2320 -331 2333 -157
rect 2379 -331 2408 -157
rect 2320 -344 2408 -331
rect 2464 -157 2568 -144
rect 2464 -331 2493 -157
rect 2539 -331 2568 -157
rect 2464 -344 2568 -331
rect 2624 -157 2728 -144
rect 2624 -331 2653 -157
rect 2699 -331 2728 -157
rect 2624 -344 2728 -331
rect 2784 -157 2888 -144
rect 2784 -331 2813 -157
rect 2859 -331 2888 -157
rect 2784 -344 2888 -331
rect 2944 -157 3048 -144
rect 2944 -331 2973 -157
rect 3019 -331 3048 -157
rect 2944 -344 3048 -331
rect 3104 -157 3208 -144
rect 3104 -331 3133 -157
rect 3179 -331 3208 -157
rect 3104 -344 3208 -331
rect 3264 -157 3352 -144
rect 3264 -331 3293 -157
rect 3339 -331 3352 -157
rect 3264 -344 3352 -331
rect 3730 -157 3818 -144
rect 3730 -331 3743 -157
rect 3789 -331 3818 -157
rect 3730 -344 3818 -331
rect 3874 -157 3978 -144
rect 3874 -331 3903 -157
rect 3949 -331 3978 -157
rect 3874 -344 3978 -331
rect 4034 -157 4138 -144
rect 4034 -331 4063 -157
rect 4109 -331 4138 -157
rect 4034 -344 4138 -331
rect 4194 -157 4298 -144
rect 4194 -331 4223 -157
rect 4269 -331 4298 -157
rect 4194 -344 4298 -331
rect 4354 -157 4458 -144
rect 4354 -331 4383 -157
rect 4429 -331 4458 -157
rect 4354 -344 4458 -331
rect 4514 -157 4618 -144
rect 4514 -331 4543 -157
rect 4589 -331 4618 -157
rect 4514 -344 4618 -331
rect 4674 -157 4762 -144
rect 4674 -331 4703 -157
rect 4749 -331 4762 -157
rect 4674 -344 4762 -331
rect 4933 -157 5021 -144
rect 4933 -331 4946 -157
rect 4992 -331 5021 -157
rect 4933 -344 5021 -331
rect 5077 -157 5165 -144
rect 5077 -331 5106 -157
rect 5152 -331 5165 -157
rect 5077 -344 5165 -331
rect 5597 -158 5685 -145
rect 5597 -332 5610 -158
rect 5656 -332 5685 -158
rect 5597 -345 5685 -332
rect 5741 -158 5829 -145
rect 5741 -332 5770 -158
rect 5816 -332 5829 -158
rect 5741 -345 5829 -332
rect 6000 -158 6088 -145
rect 6000 -332 6013 -158
rect 6059 -332 6088 -158
rect 6000 -345 6088 -332
rect 6144 -158 6248 -145
rect 6144 -332 6173 -158
rect 6219 -332 6248 -158
rect 6144 -345 6248 -332
rect 6304 -158 6408 -145
rect 6304 -332 6333 -158
rect 6379 -332 6408 -158
rect 6304 -345 6408 -332
rect 6464 -158 6568 -145
rect 6464 -332 6493 -158
rect 6539 -332 6568 -158
rect 6464 -345 6568 -332
rect 6624 -158 6728 -145
rect 6624 -332 6653 -158
rect 6699 -332 6728 -158
rect 6624 -345 6728 -332
rect 6784 -158 6888 -145
rect 6784 -332 6813 -158
rect 6859 -332 6888 -158
rect 6784 -345 6888 -332
rect 6944 -158 7032 -145
rect 6944 -332 6973 -158
rect 7019 -332 7032 -158
rect 6944 -345 7032 -332
rect 1917 -493 2005 -480
rect -691 -681 -603 -668
rect 1917 -667 1930 -493
rect 1976 -667 2005 -493
rect 1917 -680 2005 -667
rect 2061 -493 2149 -480
rect 2061 -667 2090 -493
rect 2136 -667 2149 -493
rect 2061 -680 2149 -667
rect 2320 -493 2408 -480
rect 2320 -667 2333 -493
rect 2379 -667 2408 -493
rect 2320 -680 2408 -667
rect 2464 -493 2568 -480
rect 2464 -667 2493 -493
rect 2539 -667 2568 -493
rect 2464 -680 2568 -667
rect 2624 -493 2728 -480
rect 2624 -667 2653 -493
rect 2699 -667 2728 -493
rect 2624 -680 2728 -667
rect 2784 -493 2888 -480
rect 2784 -667 2813 -493
rect 2859 -667 2888 -493
rect 2784 -680 2888 -667
rect 2944 -493 3048 -480
rect 2944 -667 2973 -493
rect 3019 -667 3048 -493
rect 2944 -680 3048 -667
rect 3104 -493 3208 -480
rect 3104 -667 3133 -493
rect 3179 -667 3208 -493
rect 3104 -680 3208 -667
rect 3264 -493 3352 -480
rect 3264 -667 3293 -493
rect 3339 -667 3352 -493
rect 3264 -680 3352 -667
rect 3730 -493 3818 -480
rect 3730 -667 3743 -493
rect 3789 -667 3818 -493
rect 3730 -680 3818 -667
rect 3874 -493 3978 -480
rect 3874 -667 3903 -493
rect 3949 -667 3978 -493
rect 3874 -680 3978 -667
rect 4034 -493 4138 -480
rect 4034 -667 4063 -493
rect 4109 -667 4138 -493
rect 4034 -680 4138 -667
rect 4194 -493 4298 -480
rect 4194 -667 4223 -493
rect 4269 -667 4298 -493
rect 4194 -680 4298 -667
rect 4354 -493 4458 -480
rect 4354 -667 4383 -493
rect 4429 -667 4458 -493
rect 4354 -680 4458 -667
rect 4514 -493 4618 -480
rect 4514 -667 4543 -493
rect 4589 -667 4618 -493
rect 4514 -680 4618 -667
rect 4674 -493 4762 -480
rect 4674 -667 4703 -493
rect 4749 -667 4762 -493
rect 4674 -680 4762 -667
rect 4933 -493 5021 -480
rect 4933 -667 4946 -493
rect 4992 -667 5021 -493
rect 4933 -680 5021 -667
rect 5077 -493 5165 -480
rect 5077 -667 5106 -493
rect 5152 -667 5165 -493
rect 5077 -680 5165 -667
rect 5597 -494 5685 -481
rect 5597 -668 5610 -494
rect 5656 -668 5685 -494
rect 5597 -681 5685 -668
rect 5741 -494 5829 -481
rect 5741 -668 5770 -494
rect 5816 -668 5829 -494
rect 5741 -681 5829 -668
rect 6000 -494 6088 -481
rect 6000 -668 6013 -494
rect 6059 -668 6088 -494
rect 6000 -681 6088 -668
rect 6144 -494 6248 -481
rect 6144 -668 6173 -494
rect 6219 -668 6248 -494
rect 6144 -681 6248 -668
rect 6304 -494 6408 -481
rect 6304 -668 6333 -494
rect 6379 -668 6408 -494
rect 6304 -681 6408 -668
rect 6464 -494 6568 -481
rect 6464 -668 6493 -494
rect 6539 -668 6568 -494
rect 6464 -681 6568 -668
rect 6624 -494 6728 -481
rect 6624 -668 6653 -494
rect 6699 -668 6728 -494
rect 6624 -681 6728 -668
rect 6784 -494 6888 -481
rect 6784 -668 6813 -494
rect 6859 -668 6888 -494
rect 6784 -681 6888 -668
rect 6944 -494 7032 -481
rect 6944 -668 6973 -494
rect 7019 -668 7032 -494
rect 6944 -681 7032 -668
rect 147 -1128 235 -1115
rect 147 -1202 160 -1128
rect 206 -1202 235 -1128
rect 147 -1215 235 -1202
rect 291 -1128 395 -1115
rect 291 -1202 320 -1128
rect 366 -1202 395 -1128
rect 291 -1215 395 -1202
rect 451 -1128 555 -1115
rect 451 -1202 480 -1128
rect 526 -1202 555 -1128
rect 451 -1215 555 -1202
rect 611 -1128 715 -1115
rect 611 -1202 640 -1128
rect 686 -1202 715 -1128
rect 611 -1215 715 -1202
rect 771 -1128 859 -1115
rect 771 -1202 800 -1128
rect 846 -1202 859 -1128
rect 771 -1215 859 -1202
rect 147 -1364 235 -1351
rect 147 -1438 160 -1364
rect 206 -1438 235 -1364
rect 147 -1451 235 -1438
rect 291 -1364 395 -1351
rect 291 -1438 320 -1364
rect 366 -1438 395 -1364
rect 291 -1451 395 -1438
rect 451 -1364 555 -1351
rect 451 -1438 480 -1364
rect 526 -1438 555 -1364
rect 451 -1451 555 -1438
rect 611 -1364 715 -1351
rect 611 -1438 640 -1364
rect 686 -1438 715 -1364
rect 611 -1451 715 -1438
rect 771 -1364 859 -1351
rect 771 -1438 800 -1364
rect 846 -1438 859 -1364
rect 771 -1451 859 -1438
rect 147 -1769 235 -1756
rect 147 -1843 160 -1769
rect 206 -1843 235 -1769
rect 147 -1856 235 -1843
rect 291 -1769 395 -1756
rect 291 -1843 320 -1769
rect 366 -1843 395 -1769
rect 291 -1856 395 -1843
rect 451 -1769 555 -1756
rect 451 -1843 480 -1769
rect 526 -1843 555 -1769
rect 451 -1856 555 -1843
rect 611 -1769 715 -1756
rect 611 -1843 640 -1769
rect 686 -1843 715 -1769
rect 611 -1856 715 -1843
rect 771 -1769 859 -1756
rect 771 -1843 800 -1769
rect 846 -1843 859 -1769
rect 771 -1856 859 -1843
rect 147 -2005 235 -1992
rect 147 -2079 160 -2005
rect 206 -2079 235 -2005
rect 147 -2092 235 -2079
rect 291 -2005 395 -1992
rect 291 -2079 320 -2005
rect 366 -2079 395 -2005
rect 291 -2092 395 -2079
rect 451 -2005 555 -1992
rect 451 -2079 480 -2005
rect 526 -2079 555 -2005
rect 451 -2092 555 -2079
rect 611 -2005 715 -1992
rect 611 -2079 640 -2005
rect 686 -2079 715 -2005
rect 611 -2092 715 -2079
rect 771 -2005 859 -1992
rect 771 -2079 800 -2005
rect 846 -2079 859 -2005
rect 771 -2092 859 -2079
rect 147 -4069 235 -4056
rect 147 -4143 160 -4069
rect 206 -4143 235 -4069
rect 147 -4156 235 -4143
rect 291 -4069 395 -4056
rect 291 -4143 320 -4069
rect 366 -4143 395 -4069
rect 291 -4156 395 -4143
rect 451 -4069 555 -4056
rect 451 -4143 480 -4069
rect 526 -4143 555 -4069
rect 451 -4156 555 -4143
rect 611 -4069 715 -4056
rect 611 -4143 640 -4069
rect 686 -4143 715 -4069
rect 611 -4156 715 -4143
rect 771 -4069 859 -4056
rect 771 -4143 800 -4069
rect 846 -4143 859 -4069
rect 771 -4156 859 -4143
rect 147 -4305 235 -4292
rect -4845 -4337 -4757 -4324
rect -4845 -4511 -4832 -4337
rect -4786 -4511 -4757 -4337
rect -4845 -4524 -4757 -4511
rect -4701 -4337 -4613 -4324
rect -4701 -4511 -4672 -4337
rect -4626 -4511 -4613 -4337
rect -4701 -4524 -4613 -4511
rect -4441 -4337 -4353 -4324
rect -4441 -4511 -4428 -4337
rect -4382 -4511 -4353 -4337
rect -4441 -4524 -4353 -4511
rect -4297 -4337 -4209 -4324
rect -4297 -4511 -4268 -4337
rect -4222 -4511 -4209 -4337
rect -4297 -4524 -4209 -4511
rect -4038 -4337 -3950 -4324
rect -4038 -4511 -4025 -4337
rect -3979 -4511 -3950 -4337
rect -4038 -4524 -3950 -4511
rect -3894 -4337 -3790 -4324
rect -3894 -4511 -3865 -4337
rect -3819 -4511 -3790 -4337
rect -3894 -4524 -3790 -4511
rect -3734 -4337 -3630 -4324
rect -3734 -4511 -3705 -4337
rect -3659 -4511 -3630 -4337
rect -3734 -4524 -3630 -4511
rect -3574 -4337 -3470 -4324
rect -3574 -4511 -3545 -4337
rect -3499 -4511 -3470 -4337
rect -3574 -4524 -3470 -4511
rect -3414 -4337 -3310 -4324
rect -3414 -4511 -3385 -4337
rect -3339 -4511 -3310 -4337
rect -3414 -4524 -3310 -4511
rect -3254 -4337 -3150 -4324
rect -3254 -4511 -3225 -4337
rect -3179 -4511 -3150 -4337
rect -3254 -4524 -3150 -4511
rect -3094 -4337 -3006 -4324
rect -3094 -4511 -3065 -4337
rect -3019 -4511 -3006 -4337
rect -3094 -4524 -3006 -4511
rect -2442 -4330 -2354 -4317
rect -2442 -4504 -2429 -4330
rect -2383 -4504 -2354 -4330
rect -2442 -4517 -2354 -4504
rect -2298 -4330 -2210 -4317
rect -2298 -4504 -2269 -4330
rect -2223 -4504 -2210 -4330
rect -2298 -4517 -2210 -4504
rect -2038 -4330 -1950 -4317
rect -2038 -4504 -2025 -4330
rect -1979 -4504 -1950 -4330
rect -2038 -4517 -1950 -4504
rect -1894 -4330 -1806 -4317
rect -1894 -4504 -1865 -4330
rect -1819 -4504 -1806 -4330
rect -1894 -4517 -1806 -4504
rect -1635 -4330 -1547 -4317
rect -1635 -4504 -1622 -4330
rect -1576 -4504 -1547 -4330
rect -1635 -4517 -1547 -4504
rect -1491 -4330 -1387 -4317
rect -1491 -4504 -1462 -4330
rect -1416 -4504 -1387 -4330
rect -1491 -4517 -1387 -4504
rect -1331 -4330 -1227 -4317
rect -1331 -4504 -1302 -4330
rect -1256 -4504 -1227 -4330
rect -1331 -4517 -1227 -4504
rect -1171 -4330 -1067 -4317
rect -1171 -4504 -1142 -4330
rect -1096 -4504 -1067 -4330
rect -1171 -4517 -1067 -4504
rect -1011 -4330 -907 -4317
rect -1011 -4504 -982 -4330
rect -936 -4504 -907 -4330
rect -1011 -4517 -907 -4504
rect -851 -4330 -747 -4317
rect -851 -4504 -822 -4330
rect -776 -4504 -747 -4330
rect -851 -4517 -747 -4504
rect -691 -4330 -603 -4317
rect -691 -4504 -662 -4330
rect -616 -4504 -603 -4330
rect 147 -4379 160 -4305
rect 206 -4379 235 -4305
rect 147 -4392 235 -4379
rect 291 -4305 395 -4292
rect 291 -4379 320 -4305
rect 366 -4379 395 -4305
rect 291 -4392 395 -4379
rect 451 -4305 555 -4292
rect 451 -4379 480 -4305
rect 526 -4379 555 -4305
rect 451 -4392 555 -4379
rect 611 -4305 715 -4292
rect 611 -4379 640 -4305
rect 686 -4379 715 -4305
rect 611 -4392 715 -4379
rect 771 -4305 859 -4292
rect 771 -4379 800 -4305
rect 846 -4379 859 -4305
rect 771 -4392 859 -4379
rect 1917 -4329 2005 -4316
rect -691 -4517 -603 -4504
rect 1917 -4503 1930 -4329
rect 1976 -4503 2005 -4329
rect 1917 -4516 2005 -4503
rect 2061 -4329 2149 -4316
rect 2061 -4503 2090 -4329
rect 2136 -4503 2149 -4329
rect 2061 -4516 2149 -4503
rect 2320 -4329 2408 -4316
rect 2320 -4503 2333 -4329
rect 2379 -4503 2408 -4329
rect 2320 -4516 2408 -4503
rect 2464 -4329 2568 -4316
rect 2464 -4503 2493 -4329
rect 2539 -4503 2568 -4329
rect 2464 -4516 2568 -4503
rect 2624 -4329 2728 -4316
rect 2624 -4503 2653 -4329
rect 2699 -4503 2728 -4329
rect 2624 -4516 2728 -4503
rect 2784 -4329 2888 -4316
rect 2784 -4503 2813 -4329
rect 2859 -4503 2888 -4329
rect 2784 -4516 2888 -4503
rect 2944 -4329 3048 -4316
rect 2944 -4503 2973 -4329
rect 3019 -4503 3048 -4329
rect 2944 -4516 3048 -4503
rect 3104 -4329 3208 -4316
rect 3104 -4503 3133 -4329
rect 3179 -4503 3208 -4329
rect 3104 -4516 3208 -4503
rect 3264 -4329 3352 -4316
rect 3264 -4503 3293 -4329
rect 3339 -4503 3352 -4329
rect 3264 -4516 3352 -4503
rect 3730 -4329 3818 -4316
rect 3730 -4503 3743 -4329
rect 3789 -4503 3818 -4329
rect 3730 -4516 3818 -4503
rect 3874 -4329 3978 -4316
rect 3874 -4503 3903 -4329
rect 3949 -4503 3978 -4329
rect 3874 -4516 3978 -4503
rect 4034 -4329 4138 -4316
rect 4034 -4503 4063 -4329
rect 4109 -4503 4138 -4329
rect 4034 -4516 4138 -4503
rect 4194 -4329 4298 -4316
rect 4194 -4503 4223 -4329
rect 4269 -4503 4298 -4329
rect 4194 -4516 4298 -4503
rect 4354 -4329 4458 -4316
rect 4354 -4503 4383 -4329
rect 4429 -4503 4458 -4329
rect 4354 -4516 4458 -4503
rect 4514 -4329 4618 -4316
rect 4514 -4503 4543 -4329
rect 4589 -4503 4618 -4329
rect 4514 -4516 4618 -4503
rect 4674 -4329 4762 -4316
rect 4674 -4503 4703 -4329
rect 4749 -4503 4762 -4329
rect 4674 -4516 4762 -4503
rect 4933 -4329 5021 -4316
rect 4933 -4503 4946 -4329
rect 4992 -4503 5021 -4329
rect 4933 -4516 5021 -4503
rect 5077 -4329 5165 -4316
rect 5077 -4503 5106 -4329
rect 5152 -4503 5165 -4329
rect 5077 -4516 5165 -4503
rect 5597 -4330 5685 -4317
rect 5597 -4504 5610 -4330
rect 5656 -4504 5685 -4330
rect 5597 -4517 5685 -4504
rect 5741 -4330 5829 -4317
rect 5741 -4504 5770 -4330
rect 5816 -4504 5829 -4330
rect 5741 -4517 5829 -4504
rect 6000 -4330 6088 -4317
rect 6000 -4504 6013 -4330
rect 6059 -4504 6088 -4330
rect 6000 -4517 6088 -4504
rect 6144 -4330 6248 -4317
rect 6144 -4504 6173 -4330
rect 6219 -4504 6248 -4330
rect 6144 -4517 6248 -4504
rect 6304 -4330 6408 -4317
rect 6304 -4504 6333 -4330
rect 6379 -4504 6408 -4330
rect 6304 -4517 6408 -4504
rect 6464 -4330 6568 -4317
rect 6464 -4504 6493 -4330
rect 6539 -4504 6568 -4330
rect 6464 -4517 6568 -4504
rect 6624 -4330 6728 -4317
rect 6624 -4504 6653 -4330
rect 6699 -4504 6728 -4330
rect 6624 -4517 6728 -4504
rect 6784 -4330 6888 -4317
rect 6784 -4504 6813 -4330
rect 6859 -4504 6888 -4330
rect 6784 -4517 6888 -4504
rect 6944 -4330 7032 -4317
rect 6944 -4504 6973 -4330
rect 7019 -4504 7032 -4330
rect 6944 -4517 7032 -4504
rect -4845 -4673 -4757 -4660
rect -4845 -4847 -4832 -4673
rect -4786 -4847 -4757 -4673
rect -4845 -4860 -4757 -4847
rect -4701 -4673 -4613 -4660
rect -4701 -4847 -4672 -4673
rect -4626 -4847 -4613 -4673
rect -4701 -4860 -4613 -4847
rect -4441 -4673 -4353 -4660
rect -4441 -4847 -4428 -4673
rect -4382 -4847 -4353 -4673
rect -4441 -4860 -4353 -4847
rect -4297 -4673 -4209 -4660
rect -4297 -4847 -4268 -4673
rect -4222 -4847 -4209 -4673
rect -4297 -4860 -4209 -4847
rect -4038 -4673 -3950 -4660
rect -4038 -4847 -4025 -4673
rect -3979 -4847 -3950 -4673
rect -4038 -4860 -3950 -4847
rect -3894 -4673 -3790 -4660
rect -3894 -4847 -3865 -4673
rect -3819 -4847 -3790 -4673
rect -3894 -4860 -3790 -4847
rect -3734 -4673 -3630 -4660
rect -3734 -4847 -3705 -4673
rect -3659 -4847 -3630 -4673
rect -3734 -4860 -3630 -4847
rect -3574 -4673 -3470 -4660
rect -3574 -4847 -3545 -4673
rect -3499 -4847 -3470 -4673
rect -3574 -4860 -3470 -4847
rect -3414 -4673 -3310 -4660
rect -3414 -4847 -3385 -4673
rect -3339 -4847 -3310 -4673
rect -3414 -4860 -3310 -4847
rect -3254 -4673 -3150 -4660
rect -3254 -4847 -3225 -4673
rect -3179 -4847 -3150 -4673
rect -3254 -4860 -3150 -4847
rect -3094 -4673 -3006 -4660
rect -3094 -4847 -3065 -4673
rect -3019 -4847 -3006 -4673
rect -3094 -4860 -3006 -4847
rect -2442 -4666 -2354 -4653
rect -2442 -4840 -2429 -4666
rect -2383 -4840 -2354 -4666
rect -2442 -4853 -2354 -4840
rect -2298 -4666 -2210 -4653
rect -2298 -4840 -2269 -4666
rect -2223 -4840 -2210 -4666
rect -2298 -4853 -2210 -4840
rect -2038 -4666 -1950 -4653
rect -2038 -4840 -2025 -4666
rect -1979 -4840 -1950 -4666
rect -2038 -4853 -1950 -4840
rect -1894 -4666 -1806 -4653
rect -1894 -4840 -1865 -4666
rect -1819 -4840 -1806 -4666
rect -1894 -4853 -1806 -4840
rect -1635 -4666 -1547 -4653
rect -1635 -4840 -1622 -4666
rect -1576 -4840 -1547 -4666
rect -1635 -4853 -1547 -4840
rect -1491 -4666 -1387 -4653
rect -1491 -4840 -1462 -4666
rect -1416 -4840 -1387 -4666
rect -1491 -4853 -1387 -4840
rect -1331 -4666 -1227 -4653
rect -1331 -4840 -1302 -4666
rect -1256 -4840 -1227 -4666
rect -1331 -4853 -1227 -4840
rect -1171 -4666 -1067 -4653
rect -1171 -4840 -1142 -4666
rect -1096 -4840 -1067 -4666
rect -1171 -4853 -1067 -4840
rect -1011 -4666 -907 -4653
rect -1011 -4840 -982 -4666
rect -936 -4840 -907 -4666
rect -1011 -4853 -907 -4840
rect -851 -4666 -747 -4653
rect -851 -4840 -822 -4666
rect -776 -4840 -747 -4666
rect -851 -4853 -747 -4840
rect -691 -4666 -603 -4653
rect -691 -4840 -662 -4666
rect -616 -4840 -603 -4666
rect -691 -4853 -603 -4840
rect 1917 -4665 2005 -4652
rect 1917 -4839 1930 -4665
rect 1976 -4839 2005 -4665
rect 1917 -4852 2005 -4839
rect 2061 -4665 2149 -4652
rect 2061 -4839 2090 -4665
rect 2136 -4839 2149 -4665
rect 2061 -4852 2149 -4839
rect 2320 -4665 2408 -4652
rect 2320 -4839 2333 -4665
rect 2379 -4839 2408 -4665
rect 2320 -4852 2408 -4839
rect 2464 -4665 2568 -4652
rect 2464 -4839 2493 -4665
rect 2539 -4839 2568 -4665
rect 2464 -4852 2568 -4839
rect 2624 -4665 2728 -4652
rect 2624 -4839 2653 -4665
rect 2699 -4839 2728 -4665
rect 2624 -4852 2728 -4839
rect 2784 -4665 2888 -4652
rect 2784 -4839 2813 -4665
rect 2859 -4839 2888 -4665
rect 2784 -4852 2888 -4839
rect 2944 -4665 3048 -4652
rect 2944 -4839 2973 -4665
rect 3019 -4839 3048 -4665
rect 2944 -4852 3048 -4839
rect 3104 -4665 3208 -4652
rect 3104 -4839 3133 -4665
rect 3179 -4839 3208 -4665
rect 3104 -4852 3208 -4839
rect 3264 -4665 3352 -4652
rect 3264 -4839 3293 -4665
rect 3339 -4839 3352 -4665
rect 3264 -4852 3352 -4839
rect 3730 -4665 3818 -4652
rect 3730 -4839 3743 -4665
rect 3789 -4839 3818 -4665
rect 3730 -4852 3818 -4839
rect 3874 -4665 3978 -4652
rect 3874 -4839 3903 -4665
rect 3949 -4839 3978 -4665
rect 3874 -4852 3978 -4839
rect 4034 -4665 4138 -4652
rect 4034 -4839 4063 -4665
rect 4109 -4839 4138 -4665
rect 4034 -4852 4138 -4839
rect 4194 -4665 4298 -4652
rect 4194 -4839 4223 -4665
rect 4269 -4839 4298 -4665
rect 4194 -4852 4298 -4839
rect 4354 -4665 4458 -4652
rect 4354 -4839 4383 -4665
rect 4429 -4839 4458 -4665
rect 4354 -4852 4458 -4839
rect 4514 -4665 4618 -4652
rect 4514 -4839 4543 -4665
rect 4589 -4839 4618 -4665
rect 4514 -4852 4618 -4839
rect 4674 -4665 4762 -4652
rect 4674 -4839 4703 -4665
rect 4749 -4839 4762 -4665
rect 4674 -4852 4762 -4839
rect 4933 -4665 5021 -4652
rect 4933 -4839 4946 -4665
rect 4992 -4839 5021 -4665
rect 4933 -4852 5021 -4839
rect 5077 -4665 5165 -4652
rect 5077 -4839 5106 -4665
rect 5152 -4839 5165 -4665
rect 5077 -4852 5165 -4839
rect 5597 -4666 5685 -4653
rect 5597 -4840 5610 -4666
rect 5656 -4840 5685 -4666
rect 5597 -4853 5685 -4840
rect 5741 -4666 5829 -4653
rect 5741 -4840 5770 -4666
rect 5816 -4840 5829 -4666
rect 5741 -4853 5829 -4840
rect 6000 -4666 6088 -4653
rect 6000 -4840 6013 -4666
rect 6059 -4840 6088 -4666
rect 6000 -4853 6088 -4840
rect 6144 -4666 6248 -4653
rect 6144 -4840 6173 -4666
rect 6219 -4840 6248 -4666
rect 6144 -4853 6248 -4840
rect 6304 -4666 6408 -4653
rect 6304 -4840 6333 -4666
rect 6379 -4840 6408 -4666
rect 6304 -4853 6408 -4840
rect 6464 -4666 6568 -4653
rect 6464 -4840 6493 -4666
rect 6539 -4840 6568 -4666
rect 6464 -4853 6568 -4840
rect 6624 -4666 6728 -4653
rect 6624 -4840 6653 -4666
rect 6699 -4840 6728 -4666
rect 6624 -4853 6728 -4840
rect 6784 -4666 6888 -4653
rect 6784 -4840 6813 -4666
rect 6859 -4840 6888 -4666
rect 6784 -4853 6888 -4840
rect 6944 -4666 7032 -4653
rect 6944 -4840 6973 -4666
rect 7019 -4840 7032 -4666
rect 6944 -4853 7032 -4840
rect -4845 -5325 -4757 -5312
rect -4845 -5499 -4832 -5325
rect -4786 -5499 -4757 -5325
rect -4845 -5512 -4757 -5499
rect -4701 -5325 -4613 -5312
rect -4701 -5499 -4672 -5325
rect -4626 -5499 -4613 -5325
rect -4701 -5512 -4613 -5499
rect -4441 -5325 -4353 -5312
rect -4441 -5499 -4428 -5325
rect -4382 -5499 -4353 -5325
rect -4441 -5512 -4353 -5499
rect -4297 -5325 -4209 -5312
rect -4297 -5499 -4268 -5325
rect -4222 -5499 -4209 -5325
rect -4297 -5512 -4209 -5499
rect -4038 -5325 -3950 -5312
rect -4038 -5499 -4025 -5325
rect -3979 -5499 -3950 -5325
rect -4038 -5512 -3950 -5499
rect -3894 -5325 -3790 -5312
rect -3894 -5499 -3865 -5325
rect -3819 -5499 -3790 -5325
rect -3894 -5512 -3790 -5499
rect -3734 -5325 -3630 -5312
rect -3734 -5499 -3705 -5325
rect -3659 -5499 -3630 -5325
rect -3734 -5512 -3630 -5499
rect -3574 -5325 -3470 -5312
rect -3574 -5499 -3545 -5325
rect -3499 -5499 -3470 -5325
rect -3574 -5512 -3470 -5499
rect -3414 -5325 -3310 -5312
rect -3414 -5499 -3385 -5325
rect -3339 -5499 -3310 -5325
rect -3414 -5512 -3310 -5499
rect -3254 -5325 -3150 -5312
rect -3254 -5499 -3225 -5325
rect -3179 -5499 -3150 -5325
rect -3254 -5512 -3150 -5499
rect -3094 -5325 -3006 -5312
rect -3094 -5499 -3065 -5325
rect -3019 -5499 -3006 -5325
rect -3094 -5512 -3006 -5499
rect -2442 -5318 -2354 -5305
rect -2442 -5492 -2429 -5318
rect -2383 -5492 -2354 -5318
rect -2442 -5505 -2354 -5492
rect -2298 -5318 -2210 -5305
rect -2298 -5492 -2269 -5318
rect -2223 -5492 -2210 -5318
rect -2298 -5505 -2210 -5492
rect -2038 -5318 -1950 -5305
rect -2038 -5492 -2025 -5318
rect -1979 -5492 -1950 -5318
rect -2038 -5505 -1950 -5492
rect -1894 -5318 -1806 -5305
rect -1894 -5492 -1865 -5318
rect -1819 -5492 -1806 -5318
rect -1894 -5505 -1806 -5492
rect -1635 -5318 -1547 -5305
rect -1635 -5492 -1622 -5318
rect -1576 -5492 -1547 -5318
rect -1635 -5505 -1547 -5492
rect -1491 -5318 -1387 -5305
rect -1491 -5492 -1462 -5318
rect -1416 -5492 -1387 -5318
rect -1491 -5505 -1387 -5492
rect -1331 -5318 -1227 -5305
rect -1331 -5492 -1302 -5318
rect -1256 -5492 -1227 -5318
rect -1331 -5505 -1227 -5492
rect -1171 -5318 -1067 -5305
rect -1171 -5492 -1142 -5318
rect -1096 -5492 -1067 -5318
rect -1171 -5505 -1067 -5492
rect -1011 -5318 -907 -5305
rect -1011 -5492 -982 -5318
rect -936 -5492 -907 -5318
rect -1011 -5505 -907 -5492
rect -851 -5318 -747 -5305
rect -851 -5492 -822 -5318
rect -776 -5492 -747 -5318
rect -851 -5505 -747 -5492
rect -691 -5318 -603 -5305
rect -691 -5492 -662 -5318
rect -616 -5492 -603 -5318
rect -691 -5505 -603 -5492
rect 157 -5317 245 -5304
rect 157 -5491 170 -5317
rect 216 -5491 245 -5317
rect 157 -5504 245 -5491
rect 301 -5317 389 -5304
rect 301 -5491 330 -5317
rect 376 -5491 389 -5317
rect 301 -5504 389 -5491
rect 560 -5317 648 -5304
rect 560 -5491 573 -5317
rect 619 -5491 648 -5317
rect 560 -5504 648 -5491
rect 704 -5317 808 -5304
rect 704 -5491 733 -5317
rect 779 -5491 808 -5317
rect 704 -5504 808 -5491
rect 864 -5317 968 -5304
rect 864 -5491 893 -5317
rect 939 -5491 968 -5317
rect 864 -5504 968 -5491
rect 1024 -5317 1128 -5304
rect 1024 -5491 1053 -5317
rect 1099 -5491 1128 -5317
rect 1024 -5504 1128 -5491
rect 1184 -5317 1288 -5304
rect 1184 -5491 1213 -5317
rect 1259 -5491 1288 -5317
rect 1184 -5504 1288 -5491
rect 1344 -5317 1448 -5304
rect 1344 -5491 1373 -5317
rect 1419 -5491 1448 -5317
rect 1344 -5504 1448 -5491
rect 1504 -5317 1592 -5304
rect 1504 -5491 1533 -5317
rect 1579 -5491 1592 -5317
rect 1504 -5504 1592 -5491
rect 1917 -5317 2005 -5304
rect 1917 -5491 1930 -5317
rect 1976 -5491 2005 -5317
rect 1917 -5504 2005 -5491
rect 2061 -5317 2165 -5304
rect 2061 -5491 2090 -5317
rect 2136 -5491 2165 -5317
rect 2061 -5504 2165 -5491
rect 2221 -5317 2325 -5304
rect 2221 -5491 2250 -5317
rect 2296 -5491 2325 -5317
rect 2221 -5504 2325 -5491
rect 2381 -5317 2485 -5304
rect 2381 -5491 2410 -5317
rect 2456 -5491 2485 -5317
rect 2381 -5504 2485 -5491
rect 2541 -5317 2645 -5304
rect 2541 -5491 2570 -5317
rect 2616 -5491 2645 -5317
rect 2541 -5504 2645 -5491
rect 2701 -5317 2805 -5304
rect 2701 -5491 2730 -5317
rect 2776 -5491 2805 -5317
rect 2701 -5504 2805 -5491
rect 2861 -5317 2949 -5304
rect 2861 -5491 2890 -5317
rect 2936 -5491 2949 -5317
rect 2861 -5504 2949 -5491
rect 3120 -5317 3208 -5304
rect 3120 -5491 3133 -5317
rect 3179 -5491 3208 -5317
rect 3120 -5504 3208 -5491
rect 3264 -5317 3352 -5304
rect 3264 -5491 3293 -5317
rect 3339 -5491 3352 -5317
rect 3264 -5504 3352 -5491
rect 3730 -5317 3818 -5304
rect 3730 -5491 3743 -5317
rect 3789 -5491 3818 -5317
rect 3730 -5504 3818 -5491
rect 3874 -5317 3962 -5304
rect 3874 -5491 3903 -5317
rect 3949 -5491 3962 -5317
rect 3874 -5504 3962 -5491
rect 4133 -5317 4221 -5304
rect 4133 -5491 4146 -5317
rect 4192 -5491 4221 -5317
rect 4133 -5504 4221 -5491
rect 4277 -5317 4381 -5304
rect 4277 -5491 4306 -5317
rect 4352 -5491 4381 -5317
rect 4277 -5504 4381 -5491
rect 4437 -5317 4541 -5304
rect 4437 -5491 4466 -5317
rect 4512 -5491 4541 -5317
rect 4437 -5504 4541 -5491
rect 4597 -5317 4701 -5304
rect 4597 -5491 4626 -5317
rect 4672 -5491 4701 -5317
rect 4597 -5504 4701 -5491
rect 4757 -5317 4861 -5304
rect 4757 -5491 4786 -5317
rect 4832 -5491 4861 -5317
rect 4757 -5504 4861 -5491
rect 4917 -5317 5021 -5304
rect 4917 -5491 4946 -5317
rect 4992 -5491 5021 -5317
rect 4917 -5504 5021 -5491
rect 5077 -5317 5165 -5304
rect 5077 -5491 5106 -5317
rect 5152 -5491 5165 -5317
rect 5077 -5504 5165 -5491
rect 5597 -5318 5685 -5305
rect 5597 -5492 5610 -5318
rect 5656 -5492 5685 -5318
rect 5597 -5505 5685 -5492
rect 5741 -5318 5845 -5305
rect 5741 -5492 5770 -5318
rect 5816 -5492 5845 -5318
rect 5741 -5505 5845 -5492
rect 5901 -5318 6005 -5305
rect 5901 -5492 5930 -5318
rect 5976 -5492 6005 -5318
rect 5901 -5505 6005 -5492
rect 6061 -5318 6165 -5305
rect 6061 -5492 6090 -5318
rect 6136 -5492 6165 -5318
rect 6061 -5505 6165 -5492
rect 6221 -5318 6325 -5305
rect 6221 -5492 6250 -5318
rect 6296 -5492 6325 -5318
rect 6221 -5505 6325 -5492
rect 6381 -5318 6485 -5305
rect 6381 -5492 6410 -5318
rect 6456 -5492 6485 -5318
rect 6381 -5505 6485 -5492
rect 6541 -5318 6629 -5305
rect 6541 -5492 6570 -5318
rect 6616 -5492 6629 -5318
rect 6541 -5505 6629 -5492
rect 6800 -5318 6888 -5305
rect 6800 -5492 6813 -5318
rect 6859 -5492 6888 -5318
rect 6800 -5505 6888 -5492
rect 6944 -5318 7032 -5305
rect 6944 -5492 6973 -5318
rect 7019 -5492 7032 -5318
rect 6944 -5505 7032 -5492
rect -4845 -5661 -4757 -5648
rect -4845 -5835 -4832 -5661
rect -4786 -5835 -4757 -5661
rect -4845 -5848 -4757 -5835
rect -4701 -5661 -4613 -5648
rect -4701 -5835 -4672 -5661
rect -4626 -5835 -4613 -5661
rect -4701 -5848 -4613 -5835
rect -4441 -5661 -4353 -5648
rect -4441 -5835 -4428 -5661
rect -4382 -5835 -4353 -5661
rect -4441 -5848 -4353 -5835
rect -4297 -5661 -4209 -5648
rect -4297 -5835 -4268 -5661
rect -4222 -5835 -4209 -5661
rect -4297 -5848 -4209 -5835
rect -4038 -5661 -3950 -5648
rect -4038 -5835 -4025 -5661
rect -3979 -5835 -3950 -5661
rect -4038 -5848 -3950 -5835
rect -3894 -5661 -3790 -5648
rect -3894 -5835 -3865 -5661
rect -3819 -5835 -3790 -5661
rect -3894 -5848 -3790 -5835
rect -3734 -5661 -3630 -5648
rect -3734 -5835 -3705 -5661
rect -3659 -5835 -3630 -5661
rect -3734 -5848 -3630 -5835
rect -3574 -5661 -3470 -5648
rect -3574 -5835 -3545 -5661
rect -3499 -5835 -3470 -5661
rect -3574 -5848 -3470 -5835
rect -3414 -5661 -3310 -5648
rect -3414 -5835 -3385 -5661
rect -3339 -5835 -3310 -5661
rect -3414 -5848 -3310 -5835
rect -3254 -5661 -3150 -5648
rect -3254 -5835 -3225 -5661
rect -3179 -5835 -3150 -5661
rect -3254 -5848 -3150 -5835
rect -3094 -5661 -3006 -5648
rect -3094 -5835 -3065 -5661
rect -3019 -5835 -3006 -5661
rect -3094 -5848 -3006 -5835
rect -2442 -5654 -2354 -5641
rect -2442 -5828 -2429 -5654
rect -2383 -5828 -2354 -5654
rect -2442 -5841 -2354 -5828
rect -2298 -5654 -2210 -5641
rect -2298 -5828 -2269 -5654
rect -2223 -5828 -2210 -5654
rect -2298 -5841 -2210 -5828
rect -2038 -5654 -1950 -5641
rect -2038 -5828 -2025 -5654
rect -1979 -5828 -1950 -5654
rect -2038 -5841 -1950 -5828
rect -1894 -5654 -1806 -5641
rect -1894 -5828 -1865 -5654
rect -1819 -5828 -1806 -5654
rect -1894 -5841 -1806 -5828
rect -1635 -5654 -1547 -5641
rect -1635 -5828 -1622 -5654
rect -1576 -5828 -1547 -5654
rect -1635 -5841 -1547 -5828
rect -1491 -5654 -1387 -5641
rect -1491 -5828 -1462 -5654
rect -1416 -5828 -1387 -5654
rect -1491 -5841 -1387 -5828
rect -1331 -5654 -1227 -5641
rect -1331 -5828 -1302 -5654
rect -1256 -5828 -1227 -5654
rect -1331 -5841 -1227 -5828
rect -1171 -5654 -1067 -5641
rect -1171 -5828 -1142 -5654
rect -1096 -5828 -1067 -5654
rect -1171 -5841 -1067 -5828
rect -1011 -5654 -907 -5641
rect -1011 -5828 -982 -5654
rect -936 -5828 -907 -5654
rect -1011 -5841 -907 -5828
rect -851 -5654 -747 -5641
rect -851 -5828 -822 -5654
rect -776 -5828 -747 -5654
rect -851 -5841 -747 -5828
rect -691 -5654 -603 -5641
rect -691 -5828 -662 -5654
rect -616 -5828 -603 -5654
rect -691 -5841 -603 -5828
rect 157 -5653 245 -5640
rect 157 -5827 170 -5653
rect 216 -5827 245 -5653
rect 157 -5840 245 -5827
rect 301 -5653 389 -5640
rect 301 -5827 330 -5653
rect 376 -5827 389 -5653
rect 301 -5840 389 -5827
rect 560 -5653 648 -5640
rect 560 -5827 573 -5653
rect 619 -5827 648 -5653
rect 560 -5840 648 -5827
rect 704 -5653 808 -5640
rect 704 -5827 733 -5653
rect 779 -5827 808 -5653
rect 704 -5840 808 -5827
rect 864 -5653 968 -5640
rect 864 -5827 893 -5653
rect 939 -5827 968 -5653
rect 864 -5840 968 -5827
rect 1024 -5653 1128 -5640
rect 1024 -5827 1053 -5653
rect 1099 -5827 1128 -5653
rect 1024 -5840 1128 -5827
rect 1184 -5653 1288 -5640
rect 1184 -5827 1213 -5653
rect 1259 -5827 1288 -5653
rect 1184 -5840 1288 -5827
rect 1344 -5653 1448 -5640
rect 1344 -5827 1373 -5653
rect 1419 -5827 1448 -5653
rect 1344 -5840 1448 -5827
rect 1504 -5653 1592 -5640
rect 1504 -5827 1533 -5653
rect 1579 -5827 1592 -5653
rect 1504 -5840 1592 -5827
rect 1917 -5653 2005 -5640
rect 1917 -5827 1930 -5653
rect 1976 -5827 2005 -5653
rect 1917 -5840 2005 -5827
rect 2061 -5653 2165 -5640
rect 2061 -5827 2090 -5653
rect 2136 -5827 2165 -5653
rect 2061 -5840 2165 -5827
rect 2221 -5653 2325 -5640
rect 2221 -5827 2250 -5653
rect 2296 -5827 2325 -5653
rect 2221 -5840 2325 -5827
rect 2381 -5653 2485 -5640
rect 2381 -5827 2410 -5653
rect 2456 -5827 2485 -5653
rect 2381 -5840 2485 -5827
rect 2541 -5653 2645 -5640
rect 2541 -5827 2570 -5653
rect 2616 -5827 2645 -5653
rect 2541 -5840 2645 -5827
rect 2701 -5653 2805 -5640
rect 2701 -5827 2730 -5653
rect 2776 -5827 2805 -5653
rect 2701 -5840 2805 -5827
rect 2861 -5653 2949 -5640
rect 2861 -5827 2890 -5653
rect 2936 -5827 2949 -5653
rect 2861 -5840 2949 -5827
rect 3120 -5653 3208 -5640
rect 3120 -5827 3133 -5653
rect 3179 -5827 3208 -5653
rect 3120 -5840 3208 -5827
rect 3264 -5653 3352 -5640
rect 3264 -5827 3293 -5653
rect 3339 -5827 3352 -5653
rect 3264 -5840 3352 -5827
rect 3730 -5653 3818 -5640
rect 3730 -5827 3743 -5653
rect 3789 -5827 3818 -5653
rect 3730 -5840 3818 -5827
rect 3874 -5653 3962 -5640
rect 3874 -5827 3903 -5653
rect 3949 -5827 3962 -5653
rect 3874 -5840 3962 -5827
rect 4133 -5653 4221 -5640
rect 4133 -5827 4146 -5653
rect 4192 -5827 4221 -5653
rect 4133 -5840 4221 -5827
rect 4277 -5653 4381 -5640
rect 4277 -5827 4306 -5653
rect 4352 -5827 4381 -5653
rect 4277 -5840 4381 -5827
rect 4437 -5653 4541 -5640
rect 4437 -5827 4466 -5653
rect 4512 -5827 4541 -5653
rect 4437 -5840 4541 -5827
rect 4597 -5653 4701 -5640
rect 4597 -5827 4626 -5653
rect 4672 -5827 4701 -5653
rect 4597 -5840 4701 -5827
rect 4757 -5653 4861 -5640
rect 4757 -5827 4786 -5653
rect 4832 -5827 4861 -5653
rect 4757 -5840 4861 -5827
rect 4917 -5653 5021 -5640
rect 4917 -5827 4946 -5653
rect 4992 -5827 5021 -5653
rect 4917 -5840 5021 -5827
rect 5077 -5653 5165 -5640
rect 5077 -5827 5106 -5653
rect 5152 -5827 5165 -5653
rect 5077 -5840 5165 -5827
rect 5597 -5654 5685 -5641
rect 5597 -5828 5610 -5654
rect 5656 -5828 5685 -5654
rect 5597 -5841 5685 -5828
rect 5741 -5654 5845 -5641
rect 5741 -5828 5770 -5654
rect 5816 -5828 5845 -5654
rect 5741 -5841 5845 -5828
rect 5901 -5654 6005 -5641
rect 5901 -5828 5930 -5654
rect 5976 -5828 6005 -5654
rect 5901 -5841 6005 -5828
rect 6061 -5654 6165 -5641
rect 6061 -5828 6090 -5654
rect 6136 -5828 6165 -5654
rect 6061 -5841 6165 -5828
rect 6221 -5654 6325 -5641
rect 6221 -5828 6250 -5654
rect 6296 -5828 6325 -5654
rect 6221 -5841 6325 -5828
rect 6381 -5654 6485 -5641
rect 6381 -5828 6410 -5654
rect 6456 -5828 6485 -5654
rect 6381 -5841 6485 -5828
rect 6541 -5654 6629 -5641
rect 6541 -5828 6570 -5654
rect 6616 -5828 6629 -5654
rect 6541 -5841 6629 -5828
rect 6800 -5654 6888 -5641
rect 6800 -5828 6813 -5654
rect 6859 -5828 6888 -5654
rect 6800 -5841 6888 -5828
rect 6944 -5654 7032 -5641
rect 6944 -5828 6973 -5654
rect 7019 -5828 7032 -5654
rect 6944 -5841 7032 -5828
<< pdiff >>
rect -4845 2413 -4757 2426
rect -4845 2239 -4832 2413
rect -4786 2239 -4757 2413
rect -4845 2226 -4757 2239
rect -4701 2413 -4613 2426
rect -4701 2239 -4672 2413
rect -4626 2239 -4613 2413
rect -4701 2226 -4613 2239
rect -4441 2413 -4353 2426
rect -4441 2239 -4428 2413
rect -4382 2239 -4353 2413
rect -4441 2226 -4353 2239
rect -4297 2413 -4209 2426
rect -4297 2239 -4268 2413
rect -4222 2239 -4209 2413
rect -4297 2226 -4209 2239
rect -4038 2413 -3950 2426
rect -4038 2239 -4025 2413
rect -3979 2239 -3950 2413
rect -4038 2226 -3950 2239
rect -3894 2413 -3790 2426
rect -3894 2239 -3865 2413
rect -3819 2239 -3790 2413
rect -3894 2226 -3790 2239
rect -3734 2413 -3630 2426
rect -3734 2239 -3705 2413
rect -3659 2239 -3630 2413
rect -3734 2226 -3630 2239
rect -3574 2413 -3470 2426
rect -3574 2239 -3545 2413
rect -3499 2239 -3470 2413
rect -3574 2226 -3470 2239
rect -3414 2413 -3310 2426
rect -3414 2239 -3385 2413
rect -3339 2239 -3310 2413
rect -3414 2226 -3310 2239
rect -3254 2413 -3150 2426
rect -3254 2239 -3225 2413
rect -3179 2239 -3150 2413
rect -3254 2226 -3150 2239
rect -3094 2413 -3006 2426
rect -3094 2239 -3065 2413
rect -3019 2239 -3006 2413
rect -3094 2226 -3006 2239
rect -2442 2420 -2354 2433
rect -2442 2246 -2429 2420
rect -2383 2246 -2354 2420
rect -2442 2233 -2354 2246
rect -2298 2420 -2210 2433
rect -2298 2246 -2269 2420
rect -2223 2246 -2210 2420
rect -2298 2233 -2210 2246
rect -2038 2420 -1950 2433
rect -2038 2246 -2025 2420
rect -1979 2246 -1950 2420
rect -2038 2233 -1950 2246
rect -1894 2420 -1806 2433
rect -1894 2246 -1865 2420
rect -1819 2246 -1806 2420
rect -1894 2233 -1806 2246
rect -1635 2420 -1547 2433
rect -1635 2246 -1622 2420
rect -1576 2246 -1547 2420
rect -1635 2233 -1547 2246
rect -1491 2420 -1387 2433
rect -1491 2246 -1462 2420
rect -1416 2246 -1387 2420
rect -1491 2233 -1387 2246
rect -1331 2420 -1227 2433
rect -1331 2246 -1302 2420
rect -1256 2246 -1227 2420
rect -1331 2233 -1227 2246
rect -1171 2420 -1067 2433
rect -1171 2246 -1142 2420
rect -1096 2246 -1067 2420
rect -1171 2233 -1067 2246
rect -1011 2420 -907 2433
rect -1011 2246 -982 2420
rect -936 2246 -907 2420
rect -1011 2233 -907 2246
rect -851 2420 -747 2433
rect -851 2246 -822 2420
rect -776 2246 -747 2420
rect -851 2233 -747 2246
rect -691 2420 -603 2433
rect -691 2246 -662 2420
rect -616 2246 -603 2420
rect -691 2233 -603 2246
rect 157 2421 245 2434
rect 157 2247 170 2421
rect 216 2247 245 2421
rect 157 2234 245 2247
rect 301 2421 389 2434
rect 301 2247 330 2421
rect 376 2247 389 2421
rect 301 2234 389 2247
rect 560 2421 648 2434
rect 560 2247 573 2421
rect 619 2247 648 2421
rect 560 2234 648 2247
rect 704 2421 808 2434
rect 704 2247 733 2421
rect 779 2247 808 2421
rect 704 2234 808 2247
rect 864 2421 968 2434
rect 864 2247 893 2421
rect 939 2247 968 2421
rect 864 2234 968 2247
rect 1024 2421 1128 2434
rect 1024 2247 1053 2421
rect 1099 2247 1128 2421
rect 1024 2234 1128 2247
rect 1184 2421 1288 2434
rect 1184 2247 1213 2421
rect 1259 2247 1288 2421
rect 1184 2234 1288 2247
rect 1344 2421 1448 2434
rect 1344 2247 1373 2421
rect 1419 2247 1448 2421
rect 1344 2234 1448 2247
rect 1504 2421 1592 2434
rect 1504 2247 1533 2421
rect 1579 2247 1592 2421
rect 1504 2234 1592 2247
rect 1917 2421 2005 2434
rect 1917 2247 1930 2421
rect 1976 2247 2005 2421
rect 1917 2234 2005 2247
rect 2061 2421 2165 2434
rect 2061 2247 2090 2421
rect 2136 2247 2165 2421
rect 2061 2234 2165 2247
rect 2221 2421 2325 2434
rect 2221 2247 2250 2421
rect 2296 2247 2325 2421
rect 2221 2234 2325 2247
rect 2381 2421 2485 2434
rect 2381 2247 2410 2421
rect 2456 2247 2485 2421
rect 2381 2234 2485 2247
rect 2541 2421 2645 2434
rect 2541 2247 2570 2421
rect 2616 2247 2645 2421
rect 2541 2234 2645 2247
rect 2701 2421 2805 2434
rect 2701 2247 2730 2421
rect 2776 2247 2805 2421
rect 2701 2234 2805 2247
rect 2861 2421 2949 2434
rect 2861 2247 2890 2421
rect 2936 2247 2949 2421
rect 2861 2234 2949 2247
rect 3120 2421 3208 2434
rect 3120 2247 3133 2421
rect 3179 2247 3208 2421
rect 3120 2234 3208 2247
rect 3264 2421 3352 2434
rect 3264 2247 3293 2421
rect 3339 2247 3352 2421
rect 3264 2234 3352 2247
rect 3730 2421 3818 2434
rect 3730 2247 3743 2421
rect 3789 2247 3818 2421
rect 3730 2234 3818 2247
rect 3874 2421 3962 2434
rect 3874 2247 3903 2421
rect 3949 2247 3962 2421
rect 3874 2234 3962 2247
rect 4133 2421 4221 2434
rect 4133 2247 4146 2421
rect 4192 2247 4221 2421
rect 4133 2234 4221 2247
rect 4277 2421 4381 2434
rect 4277 2247 4306 2421
rect 4352 2247 4381 2421
rect 4277 2234 4381 2247
rect 4437 2421 4541 2434
rect 4437 2247 4466 2421
rect 4512 2247 4541 2421
rect 4437 2234 4541 2247
rect 4597 2421 4701 2434
rect 4597 2247 4626 2421
rect 4672 2247 4701 2421
rect 4597 2234 4701 2247
rect 4757 2421 4861 2434
rect 4757 2247 4786 2421
rect 4832 2247 4861 2421
rect 4757 2234 4861 2247
rect 4917 2421 5021 2434
rect 4917 2247 4946 2421
rect 4992 2247 5021 2421
rect 4917 2234 5021 2247
rect 5077 2421 5165 2434
rect 5077 2247 5106 2421
rect 5152 2247 5165 2421
rect 5077 2234 5165 2247
rect 5597 2420 5685 2433
rect 5597 2246 5610 2420
rect 5656 2246 5685 2420
rect 5597 2233 5685 2246
rect 5741 2420 5845 2433
rect 5741 2246 5770 2420
rect 5816 2246 5845 2420
rect 5741 2233 5845 2246
rect 5901 2420 6005 2433
rect 5901 2246 5930 2420
rect 5976 2246 6005 2420
rect 5901 2233 6005 2246
rect 6061 2420 6165 2433
rect 6061 2246 6090 2420
rect 6136 2246 6165 2420
rect 6061 2233 6165 2246
rect 6221 2420 6325 2433
rect 6221 2246 6250 2420
rect 6296 2246 6325 2420
rect 6221 2233 6325 2246
rect 6381 2420 6485 2433
rect 6381 2246 6410 2420
rect 6456 2246 6485 2420
rect 6381 2233 6485 2246
rect 6541 2420 6629 2433
rect 6541 2246 6570 2420
rect 6616 2246 6629 2420
rect 6541 2233 6629 2246
rect 6800 2420 6888 2433
rect 6800 2246 6813 2420
rect 6859 2246 6888 2420
rect 6800 2233 6888 2246
rect 6944 2420 7032 2433
rect 6944 2246 6973 2420
rect 7019 2246 7032 2420
rect 6944 2233 7032 2246
rect -4845 2077 -4757 2090
rect -4845 1903 -4832 2077
rect -4786 1903 -4757 2077
rect -4845 1890 -4757 1903
rect -4701 2077 -4613 2090
rect -4701 1903 -4672 2077
rect -4626 1903 -4613 2077
rect -4701 1890 -4613 1903
rect -4441 2077 -4353 2090
rect -4441 1903 -4428 2077
rect -4382 1903 -4353 2077
rect -4441 1890 -4353 1903
rect -4297 2077 -4209 2090
rect -4297 1903 -4268 2077
rect -4222 1903 -4209 2077
rect -4297 1890 -4209 1903
rect -4038 2077 -3950 2090
rect -4038 1903 -4025 2077
rect -3979 1903 -3950 2077
rect -4038 1890 -3950 1903
rect -3894 2077 -3790 2090
rect -3894 1903 -3865 2077
rect -3819 1903 -3790 2077
rect -3894 1890 -3790 1903
rect -3734 2077 -3630 2090
rect -3734 1903 -3705 2077
rect -3659 1903 -3630 2077
rect -3734 1890 -3630 1903
rect -3574 2077 -3470 2090
rect -3574 1903 -3545 2077
rect -3499 1903 -3470 2077
rect -3574 1890 -3470 1903
rect -3414 2077 -3310 2090
rect -3414 1903 -3385 2077
rect -3339 1903 -3310 2077
rect -3414 1890 -3310 1903
rect -3254 2077 -3150 2090
rect -3254 1903 -3225 2077
rect -3179 1903 -3150 2077
rect -3254 1890 -3150 1903
rect -3094 2077 -3006 2090
rect -3094 1903 -3065 2077
rect -3019 1903 -3006 2077
rect -3094 1890 -3006 1903
rect -2442 2084 -2354 2097
rect -2442 1910 -2429 2084
rect -2383 1910 -2354 2084
rect -2442 1897 -2354 1910
rect -2298 2084 -2210 2097
rect -2298 1910 -2269 2084
rect -2223 1910 -2210 2084
rect -2298 1897 -2210 1910
rect -2038 2084 -1950 2097
rect -2038 1910 -2025 2084
rect -1979 1910 -1950 2084
rect -2038 1897 -1950 1910
rect -1894 2084 -1806 2097
rect -1894 1910 -1865 2084
rect -1819 1910 -1806 2084
rect -1894 1897 -1806 1910
rect -1635 2084 -1547 2097
rect -1635 1910 -1622 2084
rect -1576 1910 -1547 2084
rect -1635 1897 -1547 1910
rect -1491 2084 -1387 2097
rect -1491 1910 -1462 2084
rect -1416 1910 -1387 2084
rect -1491 1897 -1387 1910
rect -1331 2084 -1227 2097
rect -1331 1910 -1302 2084
rect -1256 1910 -1227 2084
rect -1331 1897 -1227 1910
rect -1171 2084 -1067 2097
rect -1171 1910 -1142 2084
rect -1096 1910 -1067 2084
rect -1171 1897 -1067 1910
rect -1011 2084 -907 2097
rect -1011 1910 -982 2084
rect -936 1910 -907 2084
rect -1011 1897 -907 1910
rect -851 2084 -747 2097
rect -851 1910 -822 2084
rect -776 1910 -747 2084
rect -851 1897 -747 1910
rect -691 2084 -603 2097
rect -691 1910 -662 2084
rect -616 1910 -603 2084
rect -691 1897 -603 1910
rect 157 2085 245 2098
rect 157 1911 170 2085
rect 216 1911 245 2085
rect 157 1898 245 1911
rect 301 2085 389 2098
rect 301 1911 330 2085
rect 376 1911 389 2085
rect 301 1898 389 1911
rect 560 2085 648 2098
rect 560 1911 573 2085
rect 619 1911 648 2085
rect 560 1898 648 1911
rect 704 2085 808 2098
rect 704 1911 733 2085
rect 779 1911 808 2085
rect 704 1898 808 1911
rect 864 2085 968 2098
rect 864 1911 893 2085
rect 939 1911 968 2085
rect 864 1898 968 1911
rect 1024 2085 1128 2098
rect 1024 1911 1053 2085
rect 1099 1911 1128 2085
rect 1024 1898 1128 1911
rect 1184 2085 1288 2098
rect 1184 1911 1213 2085
rect 1259 1911 1288 2085
rect 1184 1898 1288 1911
rect 1344 2085 1448 2098
rect 1344 1911 1373 2085
rect 1419 1911 1448 2085
rect 1344 1898 1448 1911
rect 1504 2085 1592 2098
rect 1504 1911 1533 2085
rect 1579 1911 1592 2085
rect 1504 1898 1592 1911
rect 1917 2085 2005 2098
rect 1917 1911 1930 2085
rect 1976 1911 2005 2085
rect 1917 1898 2005 1911
rect 2061 2085 2165 2098
rect 2061 1911 2090 2085
rect 2136 1911 2165 2085
rect 2061 1898 2165 1911
rect 2221 2085 2325 2098
rect 2221 1911 2250 2085
rect 2296 1911 2325 2085
rect 2221 1898 2325 1911
rect 2381 2085 2485 2098
rect 2381 1911 2410 2085
rect 2456 1911 2485 2085
rect 2381 1898 2485 1911
rect 2541 2085 2645 2098
rect 2541 1911 2570 2085
rect 2616 1911 2645 2085
rect 2541 1898 2645 1911
rect 2701 2085 2805 2098
rect 2701 1911 2730 2085
rect 2776 1911 2805 2085
rect 2701 1898 2805 1911
rect 2861 2085 2949 2098
rect 2861 1911 2890 2085
rect 2936 1911 2949 2085
rect 2861 1898 2949 1911
rect 3120 2085 3208 2098
rect 3120 1911 3133 2085
rect 3179 1911 3208 2085
rect 3120 1898 3208 1911
rect 3264 2085 3352 2098
rect 3264 1911 3293 2085
rect 3339 1911 3352 2085
rect 3264 1898 3352 1911
rect 3730 2085 3818 2098
rect 3730 1911 3743 2085
rect 3789 1911 3818 2085
rect 3730 1898 3818 1911
rect 3874 2085 3962 2098
rect 3874 1911 3903 2085
rect 3949 1911 3962 2085
rect 3874 1898 3962 1911
rect 4133 2085 4221 2098
rect 4133 1911 4146 2085
rect 4192 1911 4221 2085
rect 4133 1898 4221 1911
rect 4277 2085 4381 2098
rect 4277 1911 4306 2085
rect 4352 1911 4381 2085
rect 4277 1898 4381 1911
rect 4437 2085 4541 2098
rect 4437 1911 4466 2085
rect 4512 1911 4541 2085
rect 4437 1898 4541 1911
rect 4597 2085 4701 2098
rect 4597 1911 4626 2085
rect 4672 1911 4701 2085
rect 4597 1898 4701 1911
rect 4757 2085 4861 2098
rect 4757 1911 4786 2085
rect 4832 1911 4861 2085
rect 4757 1898 4861 1911
rect 4917 2085 5021 2098
rect 4917 1911 4946 2085
rect 4992 1911 5021 2085
rect 4917 1898 5021 1911
rect 5077 2085 5165 2098
rect 5077 1911 5106 2085
rect 5152 1911 5165 2085
rect 5077 1898 5165 1911
rect 5597 2084 5685 2097
rect 5597 1910 5610 2084
rect 5656 1910 5685 2084
rect 5597 1897 5685 1910
rect 5741 2084 5845 2097
rect 5741 1910 5770 2084
rect 5816 1910 5845 2084
rect 5741 1897 5845 1910
rect 5901 2084 6005 2097
rect 5901 1910 5930 2084
rect 5976 1910 6005 2084
rect 5901 1897 6005 1910
rect 6061 2084 6165 2097
rect 6061 1910 6090 2084
rect 6136 1910 6165 2084
rect 6061 1897 6165 1910
rect 6221 2084 6325 2097
rect 6221 1910 6250 2084
rect 6296 1910 6325 2084
rect 6221 1897 6325 1910
rect 6381 2084 6485 2097
rect 6381 1910 6410 2084
rect 6456 1910 6485 2084
rect 6381 1897 6485 1910
rect 6541 2084 6629 2097
rect 6541 1910 6570 2084
rect 6616 1910 6629 2084
rect 6541 1897 6629 1910
rect 6800 2084 6888 2097
rect 6800 1910 6813 2084
rect 6859 1910 6888 2084
rect 6800 1897 6888 1910
rect 6944 2084 7032 2097
rect 6944 1910 6973 2084
rect 7019 1910 7032 2084
rect 6944 1897 7032 1910
rect -4845 1741 -4757 1754
rect -4845 1567 -4832 1741
rect -4786 1567 -4757 1741
rect -4845 1554 -4757 1567
rect -4701 1741 -4613 1754
rect -4701 1567 -4672 1741
rect -4626 1567 -4613 1741
rect -4701 1554 -4613 1567
rect -4441 1741 -4353 1754
rect -4441 1567 -4428 1741
rect -4382 1567 -4353 1741
rect -4441 1554 -4353 1567
rect -4297 1741 -4209 1754
rect -4297 1567 -4268 1741
rect -4222 1567 -4209 1741
rect -4297 1554 -4209 1567
rect -4038 1741 -3950 1754
rect -4038 1567 -4025 1741
rect -3979 1567 -3950 1741
rect -4038 1554 -3950 1567
rect -3894 1741 -3790 1754
rect -3894 1567 -3865 1741
rect -3819 1567 -3790 1741
rect -3894 1554 -3790 1567
rect -3734 1741 -3630 1754
rect -3734 1567 -3705 1741
rect -3659 1567 -3630 1741
rect -3734 1554 -3630 1567
rect -3574 1741 -3470 1754
rect -3574 1567 -3545 1741
rect -3499 1567 -3470 1741
rect -3574 1554 -3470 1567
rect -3414 1741 -3310 1754
rect -3414 1567 -3385 1741
rect -3339 1567 -3310 1741
rect -3414 1554 -3310 1567
rect -3254 1741 -3150 1754
rect -3254 1567 -3225 1741
rect -3179 1567 -3150 1741
rect -3254 1554 -3150 1567
rect -3094 1741 -3006 1754
rect -3094 1567 -3065 1741
rect -3019 1567 -3006 1741
rect -3094 1554 -3006 1567
rect -2442 1748 -2354 1761
rect -2442 1574 -2429 1748
rect -2383 1574 -2354 1748
rect -2442 1561 -2354 1574
rect -2298 1748 -2210 1761
rect -2298 1574 -2269 1748
rect -2223 1574 -2210 1748
rect -2298 1561 -2210 1574
rect -2038 1748 -1950 1761
rect -2038 1574 -2025 1748
rect -1979 1574 -1950 1748
rect -2038 1561 -1950 1574
rect -1894 1748 -1806 1761
rect -1894 1574 -1865 1748
rect -1819 1574 -1806 1748
rect -1894 1561 -1806 1574
rect -1635 1748 -1547 1761
rect -1635 1574 -1622 1748
rect -1576 1574 -1547 1748
rect -1635 1561 -1547 1574
rect -1491 1748 -1387 1761
rect -1491 1574 -1462 1748
rect -1416 1574 -1387 1748
rect -1491 1561 -1387 1574
rect -1331 1748 -1227 1761
rect -1331 1574 -1302 1748
rect -1256 1574 -1227 1748
rect -1331 1561 -1227 1574
rect -1171 1748 -1067 1761
rect -1171 1574 -1142 1748
rect -1096 1574 -1067 1748
rect -1171 1561 -1067 1574
rect -1011 1748 -907 1761
rect -1011 1574 -982 1748
rect -936 1574 -907 1748
rect -1011 1561 -907 1574
rect -851 1748 -747 1761
rect -851 1574 -822 1748
rect -776 1574 -747 1748
rect -851 1561 -747 1574
rect -691 1748 -603 1761
rect -691 1574 -662 1748
rect -616 1574 -603 1748
rect -691 1561 -603 1574
rect 157 1749 245 1762
rect 157 1575 170 1749
rect 216 1575 245 1749
rect 157 1562 245 1575
rect 301 1749 389 1762
rect 301 1575 330 1749
rect 376 1575 389 1749
rect 301 1562 389 1575
rect 560 1749 648 1762
rect 560 1575 573 1749
rect 619 1575 648 1749
rect 560 1562 648 1575
rect 704 1749 808 1762
rect 704 1575 733 1749
rect 779 1575 808 1749
rect 704 1562 808 1575
rect 864 1749 968 1762
rect 864 1575 893 1749
rect 939 1575 968 1749
rect 864 1562 968 1575
rect 1024 1749 1128 1762
rect 1024 1575 1053 1749
rect 1099 1575 1128 1749
rect 1024 1562 1128 1575
rect 1184 1749 1288 1762
rect 1184 1575 1213 1749
rect 1259 1575 1288 1749
rect 1184 1562 1288 1575
rect 1344 1749 1448 1762
rect 1344 1575 1373 1749
rect 1419 1575 1448 1749
rect 1344 1562 1448 1575
rect 1504 1749 1592 1762
rect 1504 1575 1533 1749
rect 1579 1575 1592 1749
rect 1504 1562 1592 1575
rect 1917 1749 2005 1762
rect 1917 1575 1930 1749
rect 1976 1575 2005 1749
rect 1917 1562 2005 1575
rect 2061 1749 2165 1762
rect 2061 1575 2090 1749
rect 2136 1575 2165 1749
rect 2061 1562 2165 1575
rect 2221 1749 2325 1762
rect 2221 1575 2250 1749
rect 2296 1575 2325 1749
rect 2221 1562 2325 1575
rect 2381 1749 2485 1762
rect 2381 1575 2410 1749
rect 2456 1575 2485 1749
rect 2381 1562 2485 1575
rect 2541 1749 2645 1762
rect 2541 1575 2570 1749
rect 2616 1575 2645 1749
rect 2541 1562 2645 1575
rect 2701 1749 2805 1762
rect 2701 1575 2730 1749
rect 2776 1575 2805 1749
rect 2701 1562 2805 1575
rect 2861 1749 2949 1762
rect 2861 1575 2890 1749
rect 2936 1575 2949 1749
rect 2861 1562 2949 1575
rect 3120 1749 3208 1762
rect 3120 1575 3133 1749
rect 3179 1575 3208 1749
rect 3120 1562 3208 1575
rect 3264 1749 3352 1762
rect 3264 1575 3293 1749
rect 3339 1575 3352 1749
rect 3264 1562 3352 1575
rect 3730 1749 3818 1762
rect 3730 1575 3743 1749
rect 3789 1575 3818 1749
rect 3730 1562 3818 1575
rect 3874 1749 3962 1762
rect 3874 1575 3903 1749
rect 3949 1575 3962 1749
rect 3874 1562 3962 1575
rect 4133 1749 4221 1762
rect 4133 1575 4146 1749
rect 4192 1575 4221 1749
rect 4133 1562 4221 1575
rect 4277 1749 4381 1762
rect 4277 1575 4306 1749
rect 4352 1575 4381 1749
rect 4277 1562 4381 1575
rect 4437 1749 4541 1762
rect 4437 1575 4466 1749
rect 4512 1575 4541 1749
rect 4437 1562 4541 1575
rect 4597 1749 4701 1762
rect 4597 1575 4626 1749
rect 4672 1575 4701 1749
rect 4597 1562 4701 1575
rect 4757 1749 4861 1762
rect 4757 1575 4786 1749
rect 4832 1575 4861 1749
rect 4757 1562 4861 1575
rect 4917 1749 5021 1762
rect 4917 1575 4946 1749
rect 4992 1575 5021 1749
rect 4917 1562 5021 1575
rect 5077 1749 5165 1762
rect 5077 1575 5106 1749
rect 5152 1575 5165 1749
rect 5077 1562 5165 1575
rect 5597 1748 5685 1761
rect 5597 1574 5610 1748
rect 5656 1574 5685 1748
rect 5597 1561 5685 1574
rect 5741 1748 5845 1761
rect 5741 1574 5770 1748
rect 5816 1574 5845 1748
rect 5741 1561 5845 1574
rect 5901 1748 6005 1761
rect 5901 1574 5930 1748
rect 5976 1574 6005 1748
rect 5901 1561 6005 1574
rect 6061 1748 6165 1761
rect 6061 1574 6090 1748
rect 6136 1574 6165 1748
rect 6061 1561 6165 1574
rect 6221 1748 6325 1761
rect 6221 1574 6250 1748
rect 6296 1574 6325 1748
rect 6221 1561 6325 1574
rect 6381 1748 6485 1761
rect 6381 1574 6410 1748
rect 6456 1574 6485 1748
rect 6381 1561 6485 1574
rect 6541 1748 6629 1761
rect 6541 1574 6570 1748
rect 6616 1574 6629 1748
rect 6541 1561 6629 1574
rect 6800 1748 6888 1761
rect 6800 1574 6813 1748
rect 6859 1574 6888 1748
rect 6800 1561 6888 1574
rect 6944 1748 7032 1761
rect 6944 1574 6973 1748
rect 7019 1574 7032 1748
rect 6944 1561 7032 1574
rect -4845 1405 -4757 1418
rect -4845 1231 -4832 1405
rect -4786 1231 -4757 1405
rect -4845 1218 -4757 1231
rect -4701 1405 -4613 1418
rect -4701 1231 -4672 1405
rect -4626 1231 -4613 1405
rect -4701 1218 -4613 1231
rect -4441 1405 -4353 1418
rect -4441 1231 -4428 1405
rect -4382 1231 -4353 1405
rect -4441 1218 -4353 1231
rect -4297 1405 -4209 1418
rect -4297 1231 -4268 1405
rect -4222 1231 -4209 1405
rect -4297 1218 -4209 1231
rect -4038 1405 -3950 1418
rect -4038 1231 -4025 1405
rect -3979 1231 -3950 1405
rect -4038 1218 -3950 1231
rect -3894 1405 -3790 1418
rect -3894 1231 -3865 1405
rect -3819 1231 -3790 1405
rect -3894 1218 -3790 1231
rect -3734 1405 -3630 1418
rect -3734 1231 -3705 1405
rect -3659 1231 -3630 1405
rect -3734 1218 -3630 1231
rect -3574 1405 -3470 1418
rect -3574 1231 -3545 1405
rect -3499 1231 -3470 1405
rect -3574 1218 -3470 1231
rect -3414 1405 -3310 1418
rect -3414 1231 -3385 1405
rect -3339 1231 -3310 1405
rect -3414 1218 -3310 1231
rect -3254 1405 -3150 1418
rect -3254 1231 -3225 1405
rect -3179 1231 -3150 1405
rect -3254 1218 -3150 1231
rect -3094 1405 -3006 1418
rect -3094 1231 -3065 1405
rect -3019 1231 -3006 1405
rect -3094 1218 -3006 1231
rect -2442 1412 -2354 1425
rect -2442 1238 -2429 1412
rect -2383 1238 -2354 1412
rect -2442 1225 -2354 1238
rect -2298 1412 -2210 1425
rect -2298 1238 -2269 1412
rect -2223 1238 -2210 1412
rect -2298 1225 -2210 1238
rect -2038 1412 -1950 1425
rect -2038 1238 -2025 1412
rect -1979 1238 -1950 1412
rect -2038 1225 -1950 1238
rect -1894 1412 -1806 1425
rect -1894 1238 -1865 1412
rect -1819 1238 -1806 1412
rect -1894 1225 -1806 1238
rect -1635 1412 -1547 1425
rect -1635 1238 -1622 1412
rect -1576 1238 -1547 1412
rect -1635 1225 -1547 1238
rect -1491 1412 -1387 1425
rect -1491 1238 -1462 1412
rect -1416 1238 -1387 1412
rect -1491 1225 -1387 1238
rect -1331 1412 -1227 1425
rect -1331 1238 -1302 1412
rect -1256 1238 -1227 1412
rect -1331 1225 -1227 1238
rect -1171 1412 -1067 1425
rect -1171 1238 -1142 1412
rect -1096 1238 -1067 1412
rect -1171 1225 -1067 1238
rect -1011 1412 -907 1425
rect -1011 1238 -982 1412
rect -936 1238 -907 1412
rect -1011 1225 -907 1238
rect -851 1412 -747 1425
rect -851 1238 -822 1412
rect -776 1238 -747 1412
rect -851 1225 -747 1238
rect -691 1412 -603 1425
rect -691 1238 -662 1412
rect -616 1238 -603 1412
rect -691 1225 -603 1238
rect 157 1413 245 1426
rect 157 1239 170 1413
rect 216 1239 245 1413
rect 157 1226 245 1239
rect 301 1413 389 1426
rect 301 1239 330 1413
rect 376 1239 389 1413
rect 301 1226 389 1239
rect 560 1413 648 1426
rect 560 1239 573 1413
rect 619 1239 648 1413
rect 560 1226 648 1239
rect 704 1413 808 1426
rect 704 1239 733 1413
rect 779 1239 808 1413
rect 704 1226 808 1239
rect 864 1413 968 1426
rect 864 1239 893 1413
rect 939 1239 968 1413
rect 864 1226 968 1239
rect 1024 1413 1128 1426
rect 1024 1239 1053 1413
rect 1099 1239 1128 1413
rect 1024 1226 1128 1239
rect 1184 1413 1288 1426
rect 1184 1239 1213 1413
rect 1259 1239 1288 1413
rect 1184 1226 1288 1239
rect 1344 1413 1448 1426
rect 1344 1239 1373 1413
rect 1419 1239 1448 1413
rect 1344 1226 1448 1239
rect 1504 1413 1592 1426
rect 1504 1239 1533 1413
rect 1579 1239 1592 1413
rect 1504 1226 1592 1239
rect 1917 1413 2005 1426
rect 1917 1239 1930 1413
rect 1976 1239 2005 1413
rect 1917 1226 2005 1239
rect 2061 1413 2165 1426
rect 2061 1239 2090 1413
rect 2136 1239 2165 1413
rect 2061 1226 2165 1239
rect 2221 1413 2325 1426
rect 2221 1239 2250 1413
rect 2296 1239 2325 1413
rect 2221 1226 2325 1239
rect 2381 1413 2485 1426
rect 2381 1239 2410 1413
rect 2456 1239 2485 1413
rect 2381 1226 2485 1239
rect 2541 1413 2645 1426
rect 2541 1239 2570 1413
rect 2616 1239 2645 1413
rect 2541 1226 2645 1239
rect 2701 1413 2805 1426
rect 2701 1239 2730 1413
rect 2776 1239 2805 1413
rect 2701 1226 2805 1239
rect 2861 1413 2949 1426
rect 2861 1239 2890 1413
rect 2936 1239 2949 1413
rect 2861 1226 2949 1239
rect 3120 1413 3208 1426
rect 3120 1239 3133 1413
rect 3179 1239 3208 1413
rect 3120 1226 3208 1239
rect 3264 1413 3352 1426
rect 3264 1239 3293 1413
rect 3339 1239 3352 1413
rect 3264 1226 3352 1239
rect 3730 1413 3818 1426
rect 3730 1239 3743 1413
rect 3789 1239 3818 1413
rect 3730 1226 3818 1239
rect 3874 1413 3962 1426
rect 3874 1239 3903 1413
rect 3949 1239 3962 1413
rect 3874 1226 3962 1239
rect 4133 1413 4221 1426
rect 4133 1239 4146 1413
rect 4192 1239 4221 1413
rect 4133 1226 4221 1239
rect 4277 1413 4381 1426
rect 4277 1239 4306 1413
rect 4352 1239 4381 1413
rect 4277 1226 4381 1239
rect 4437 1413 4541 1426
rect 4437 1239 4466 1413
rect 4512 1239 4541 1413
rect 4437 1226 4541 1239
rect 4597 1413 4701 1426
rect 4597 1239 4626 1413
rect 4672 1239 4701 1413
rect 4597 1226 4701 1239
rect 4757 1413 4861 1426
rect 4757 1239 4786 1413
rect 4832 1239 4861 1413
rect 4757 1226 4861 1239
rect 4917 1413 5021 1426
rect 4917 1239 4946 1413
rect 4992 1239 5021 1413
rect 4917 1226 5021 1239
rect 5077 1413 5165 1426
rect 5077 1239 5106 1413
rect 5152 1239 5165 1413
rect 5077 1226 5165 1239
rect 5597 1412 5685 1425
rect 5597 1238 5610 1412
rect 5656 1238 5685 1412
rect 5597 1225 5685 1238
rect 5741 1412 5845 1425
rect 5741 1238 5770 1412
rect 5816 1238 5845 1412
rect 5741 1225 5845 1238
rect 5901 1412 6005 1425
rect 5901 1238 5930 1412
rect 5976 1238 6005 1412
rect 5901 1225 6005 1238
rect 6061 1412 6165 1425
rect 6061 1238 6090 1412
rect 6136 1238 6165 1412
rect 6061 1225 6165 1238
rect 6221 1412 6325 1425
rect 6221 1238 6250 1412
rect 6296 1238 6325 1412
rect 6221 1225 6325 1238
rect 6381 1412 6485 1425
rect 6381 1238 6410 1412
rect 6456 1238 6485 1412
rect 6381 1225 6485 1238
rect 6541 1412 6629 1425
rect 6541 1238 6570 1412
rect 6616 1238 6629 1412
rect 6541 1225 6629 1238
rect 6800 1412 6888 1425
rect 6800 1238 6813 1412
rect 6859 1238 6888 1412
rect 6800 1225 6888 1238
rect 6944 1412 7032 1425
rect 6944 1238 6973 1412
rect 7019 1238 7032 1412
rect 6944 1225 7032 1238
rect 147 -343 235 -330
rect 147 -517 160 -343
rect 206 -517 235 -343
rect 147 -530 235 -517
rect 291 -343 395 -330
rect 291 -517 320 -343
rect 366 -517 395 -343
rect 291 -530 395 -517
rect 451 -343 555 -330
rect 451 -517 480 -343
rect 526 -517 555 -343
rect 451 -530 555 -517
rect 611 -343 715 -330
rect 611 -517 640 -343
rect 686 -517 715 -343
rect 611 -530 715 -517
rect 771 -343 859 -330
rect 771 -517 800 -343
rect 846 -517 859 -343
rect 771 -530 859 -517
rect 147 -679 235 -666
rect 147 -853 160 -679
rect 206 -853 235 -679
rect 147 -866 235 -853
rect 291 -679 395 -666
rect 291 -853 320 -679
rect 366 -853 395 -679
rect 291 -866 395 -853
rect 451 -679 555 -666
rect 451 -853 480 -679
rect 526 -853 555 -679
rect 451 -866 555 -853
rect 611 -679 715 -666
rect 611 -853 640 -679
rect 686 -853 715 -679
rect 611 -866 715 -853
rect 771 -679 859 -666
rect 771 -853 800 -679
rect 846 -853 859 -679
rect 771 -866 859 -853
rect -4845 -1083 -4757 -1070
rect -4845 -1257 -4832 -1083
rect -4786 -1257 -4757 -1083
rect -4845 -1270 -4757 -1257
rect -4701 -1083 -4613 -1070
rect -4701 -1257 -4672 -1083
rect -4626 -1257 -4613 -1083
rect -4701 -1270 -4613 -1257
rect -4441 -1083 -4353 -1070
rect -4441 -1257 -4428 -1083
rect -4382 -1257 -4353 -1083
rect -4441 -1270 -4353 -1257
rect -4297 -1083 -4209 -1070
rect -4297 -1257 -4268 -1083
rect -4222 -1257 -4209 -1083
rect -4297 -1270 -4209 -1257
rect -4038 -1083 -3950 -1070
rect -4038 -1257 -4025 -1083
rect -3979 -1257 -3950 -1083
rect -4038 -1270 -3950 -1257
rect -3894 -1083 -3790 -1070
rect -3894 -1257 -3865 -1083
rect -3819 -1257 -3790 -1083
rect -3894 -1270 -3790 -1257
rect -3734 -1083 -3630 -1070
rect -3734 -1257 -3705 -1083
rect -3659 -1257 -3630 -1083
rect -3734 -1270 -3630 -1257
rect -3574 -1083 -3470 -1070
rect -3574 -1257 -3545 -1083
rect -3499 -1257 -3470 -1083
rect -3574 -1270 -3470 -1257
rect -3414 -1083 -3310 -1070
rect -3414 -1257 -3385 -1083
rect -3339 -1257 -3310 -1083
rect -3414 -1270 -3310 -1257
rect -3254 -1083 -3150 -1070
rect -3254 -1257 -3225 -1083
rect -3179 -1257 -3150 -1083
rect -3254 -1270 -3150 -1257
rect -3094 -1083 -3006 -1070
rect -3094 -1257 -3065 -1083
rect -3019 -1257 -3006 -1083
rect -3094 -1270 -3006 -1257
rect -2442 -1076 -2354 -1063
rect -2442 -1250 -2429 -1076
rect -2383 -1250 -2354 -1076
rect -2442 -1263 -2354 -1250
rect -2298 -1076 -2210 -1063
rect -2298 -1250 -2269 -1076
rect -2223 -1250 -2210 -1076
rect -2298 -1263 -2210 -1250
rect -2038 -1076 -1950 -1063
rect -2038 -1250 -2025 -1076
rect -1979 -1250 -1950 -1076
rect -2038 -1263 -1950 -1250
rect -1894 -1076 -1806 -1063
rect -1894 -1250 -1865 -1076
rect -1819 -1250 -1806 -1076
rect -1894 -1263 -1806 -1250
rect -1635 -1076 -1547 -1063
rect -1635 -1250 -1622 -1076
rect -1576 -1250 -1547 -1076
rect -1635 -1263 -1547 -1250
rect -1491 -1076 -1387 -1063
rect -1491 -1250 -1462 -1076
rect -1416 -1250 -1387 -1076
rect -1491 -1263 -1387 -1250
rect -1331 -1076 -1227 -1063
rect -1331 -1250 -1302 -1076
rect -1256 -1250 -1227 -1076
rect -1331 -1263 -1227 -1250
rect -1171 -1076 -1067 -1063
rect -1171 -1250 -1142 -1076
rect -1096 -1250 -1067 -1076
rect -1171 -1263 -1067 -1250
rect -1011 -1076 -907 -1063
rect -1011 -1250 -982 -1076
rect -936 -1250 -907 -1076
rect -1011 -1263 -907 -1250
rect -851 -1076 -747 -1063
rect -851 -1250 -822 -1076
rect -776 -1250 -747 -1076
rect -851 -1263 -747 -1250
rect -691 -1076 -603 -1063
rect -691 -1250 -662 -1076
rect -616 -1250 -603 -1076
rect 1917 -1075 2005 -1062
rect -691 -1263 -603 -1250
rect 1917 -1249 1930 -1075
rect 1976 -1249 2005 -1075
rect 1917 -1262 2005 -1249
rect 2061 -1075 2149 -1062
rect 2061 -1249 2090 -1075
rect 2136 -1249 2149 -1075
rect 2061 -1262 2149 -1249
rect 2320 -1075 2408 -1062
rect 2320 -1249 2333 -1075
rect 2379 -1249 2408 -1075
rect 2320 -1262 2408 -1249
rect 2464 -1075 2568 -1062
rect 2464 -1249 2493 -1075
rect 2539 -1249 2568 -1075
rect 2464 -1262 2568 -1249
rect 2624 -1075 2728 -1062
rect 2624 -1249 2653 -1075
rect 2699 -1249 2728 -1075
rect 2624 -1262 2728 -1249
rect 2784 -1075 2888 -1062
rect 2784 -1249 2813 -1075
rect 2859 -1249 2888 -1075
rect 2784 -1262 2888 -1249
rect 2944 -1075 3048 -1062
rect 2944 -1249 2973 -1075
rect 3019 -1249 3048 -1075
rect 2944 -1262 3048 -1249
rect 3104 -1075 3208 -1062
rect 3104 -1249 3133 -1075
rect 3179 -1249 3208 -1075
rect 3104 -1262 3208 -1249
rect 3264 -1075 3352 -1062
rect 3264 -1249 3293 -1075
rect 3339 -1249 3352 -1075
rect 3264 -1262 3352 -1249
rect 3730 -1075 3818 -1062
rect 3730 -1249 3743 -1075
rect 3789 -1249 3818 -1075
rect 3730 -1262 3818 -1249
rect 3874 -1075 3978 -1062
rect 3874 -1249 3903 -1075
rect 3949 -1249 3978 -1075
rect 3874 -1262 3978 -1249
rect 4034 -1075 4138 -1062
rect 4034 -1249 4063 -1075
rect 4109 -1249 4138 -1075
rect 4034 -1262 4138 -1249
rect 4194 -1075 4298 -1062
rect 4194 -1249 4223 -1075
rect 4269 -1249 4298 -1075
rect 4194 -1262 4298 -1249
rect 4354 -1075 4458 -1062
rect 4354 -1249 4383 -1075
rect 4429 -1249 4458 -1075
rect 4354 -1262 4458 -1249
rect 4514 -1075 4618 -1062
rect 4514 -1249 4543 -1075
rect 4589 -1249 4618 -1075
rect 4514 -1262 4618 -1249
rect 4674 -1075 4762 -1062
rect 4674 -1249 4703 -1075
rect 4749 -1249 4762 -1075
rect 4674 -1262 4762 -1249
rect 4933 -1075 5021 -1062
rect 4933 -1249 4946 -1075
rect 4992 -1249 5021 -1075
rect 4933 -1262 5021 -1249
rect 5077 -1075 5165 -1062
rect 5077 -1249 5106 -1075
rect 5152 -1249 5165 -1075
rect 5077 -1262 5165 -1249
rect 5597 -1076 5685 -1063
rect 5597 -1250 5610 -1076
rect 5656 -1250 5685 -1076
rect -4845 -1419 -4757 -1406
rect -4845 -1593 -4832 -1419
rect -4786 -1593 -4757 -1419
rect -4845 -1606 -4757 -1593
rect -4701 -1419 -4613 -1406
rect -4701 -1593 -4672 -1419
rect -4626 -1593 -4613 -1419
rect -4701 -1606 -4613 -1593
rect -4441 -1419 -4353 -1406
rect -4441 -1593 -4428 -1419
rect -4382 -1593 -4353 -1419
rect -4441 -1606 -4353 -1593
rect -4297 -1419 -4209 -1406
rect -4297 -1593 -4268 -1419
rect -4222 -1593 -4209 -1419
rect -4297 -1606 -4209 -1593
rect -4038 -1419 -3950 -1406
rect -4038 -1593 -4025 -1419
rect -3979 -1593 -3950 -1419
rect -4038 -1606 -3950 -1593
rect -3894 -1419 -3790 -1406
rect -3894 -1593 -3865 -1419
rect -3819 -1593 -3790 -1419
rect -3894 -1606 -3790 -1593
rect -3734 -1419 -3630 -1406
rect -3734 -1593 -3705 -1419
rect -3659 -1593 -3630 -1419
rect -3734 -1606 -3630 -1593
rect -3574 -1419 -3470 -1406
rect -3574 -1593 -3545 -1419
rect -3499 -1593 -3470 -1419
rect -3574 -1606 -3470 -1593
rect -3414 -1419 -3310 -1406
rect -3414 -1593 -3385 -1419
rect -3339 -1593 -3310 -1419
rect -3414 -1606 -3310 -1593
rect -3254 -1419 -3150 -1406
rect -3254 -1593 -3225 -1419
rect -3179 -1593 -3150 -1419
rect -3254 -1606 -3150 -1593
rect -3094 -1419 -3006 -1406
rect -3094 -1593 -3065 -1419
rect -3019 -1593 -3006 -1419
rect -3094 -1606 -3006 -1593
rect -2442 -1412 -2354 -1399
rect -2442 -1586 -2429 -1412
rect -2383 -1586 -2354 -1412
rect -2442 -1599 -2354 -1586
rect -2298 -1412 -2210 -1399
rect -2298 -1586 -2269 -1412
rect -2223 -1586 -2210 -1412
rect -2298 -1599 -2210 -1586
rect -2038 -1412 -1950 -1399
rect -2038 -1586 -2025 -1412
rect -1979 -1586 -1950 -1412
rect -2038 -1599 -1950 -1586
rect -1894 -1412 -1806 -1399
rect -1894 -1586 -1865 -1412
rect -1819 -1586 -1806 -1412
rect -1894 -1599 -1806 -1586
rect -1635 -1412 -1547 -1399
rect -1635 -1586 -1622 -1412
rect -1576 -1586 -1547 -1412
rect -1635 -1599 -1547 -1586
rect -1491 -1412 -1387 -1399
rect -1491 -1586 -1462 -1412
rect -1416 -1586 -1387 -1412
rect -1491 -1599 -1387 -1586
rect -1331 -1412 -1227 -1399
rect -1331 -1586 -1302 -1412
rect -1256 -1586 -1227 -1412
rect -1331 -1599 -1227 -1586
rect -1171 -1412 -1067 -1399
rect -1171 -1586 -1142 -1412
rect -1096 -1586 -1067 -1412
rect -1171 -1599 -1067 -1586
rect -1011 -1412 -907 -1399
rect -1011 -1586 -982 -1412
rect -936 -1586 -907 -1412
rect -1011 -1599 -907 -1586
rect -851 -1412 -747 -1399
rect -851 -1586 -822 -1412
rect -776 -1586 -747 -1412
rect -851 -1599 -747 -1586
rect -691 -1412 -603 -1399
rect -691 -1586 -662 -1412
rect -616 -1586 -603 -1412
rect 5597 -1263 5685 -1250
rect 5741 -1076 5829 -1063
rect 5741 -1250 5770 -1076
rect 5816 -1250 5829 -1076
rect 5741 -1263 5829 -1250
rect 6000 -1076 6088 -1063
rect 6000 -1250 6013 -1076
rect 6059 -1250 6088 -1076
rect 6000 -1263 6088 -1250
rect 6144 -1076 6248 -1063
rect 6144 -1250 6173 -1076
rect 6219 -1250 6248 -1076
rect 6144 -1263 6248 -1250
rect 6304 -1076 6408 -1063
rect 6304 -1250 6333 -1076
rect 6379 -1250 6408 -1076
rect 6304 -1263 6408 -1250
rect 6464 -1076 6568 -1063
rect 6464 -1250 6493 -1076
rect 6539 -1250 6568 -1076
rect 6464 -1263 6568 -1250
rect 6624 -1076 6728 -1063
rect 6624 -1250 6653 -1076
rect 6699 -1250 6728 -1076
rect 6624 -1263 6728 -1250
rect 6784 -1076 6888 -1063
rect 6784 -1250 6813 -1076
rect 6859 -1250 6888 -1076
rect 6784 -1263 6888 -1250
rect 6944 -1076 7032 -1063
rect 6944 -1250 6973 -1076
rect 7019 -1250 7032 -1076
rect 6944 -1263 7032 -1250
rect 1917 -1411 2005 -1398
rect -691 -1599 -603 -1586
rect 1917 -1585 1930 -1411
rect 1976 -1585 2005 -1411
rect 1917 -1598 2005 -1585
rect 2061 -1411 2149 -1398
rect 2061 -1585 2090 -1411
rect 2136 -1585 2149 -1411
rect 2061 -1598 2149 -1585
rect 2320 -1411 2408 -1398
rect 2320 -1585 2333 -1411
rect 2379 -1585 2408 -1411
rect 2320 -1598 2408 -1585
rect 2464 -1411 2568 -1398
rect 2464 -1585 2493 -1411
rect 2539 -1585 2568 -1411
rect 2464 -1598 2568 -1585
rect 2624 -1411 2728 -1398
rect 2624 -1585 2653 -1411
rect 2699 -1585 2728 -1411
rect 2624 -1598 2728 -1585
rect 2784 -1411 2888 -1398
rect 2784 -1585 2813 -1411
rect 2859 -1585 2888 -1411
rect 2784 -1598 2888 -1585
rect 2944 -1411 3048 -1398
rect 2944 -1585 2973 -1411
rect 3019 -1585 3048 -1411
rect 2944 -1598 3048 -1585
rect 3104 -1411 3208 -1398
rect 3104 -1585 3133 -1411
rect 3179 -1585 3208 -1411
rect 3104 -1598 3208 -1585
rect 3264 -1411 3352 -1398
rect 3264 -1585 3293 -1411
rect 3339 -1585 3352 -1411
rect 3264 -1598 3352 -1585
rect 3730 -1411 3818 -1398
rect 3730 -1585 3743 -1411
rect 3789 -1585 3818 -1411
rect 3730 -1598 3818 -1585
rect 3874 -1411 3978 -1398
rect 3874 -1585 3903 -1411
rect 3949 -1585 3978 -1411
rect 3874 -1598 3978 -1585
rect 4034 -1411 4138 -1398
rect 4034 -1585 4063 -1411
rect 4109 -1585 4138 -1411
rect 4034 -1598 4138 -1585
rect 4194 -1411 4298 -1398
rect 4194 -1585 4223 -1411
rect 4269 -1585 4298 -1411
rect 4194 -1598 4298 -1585
rect 4354 -1411 4458 -1398
rect 4354 -1585 4383 -1411
rect 4429 -1585 4458 -1411
rect 4354 -1598 4458 -1585
rect 4514 -1411 4618 -1398
rect 4514 -1585 4543 -1411
rect 4589 -1585 4618 -1411
rect 4514 -1598 4618 -1585
rect 4674 -1411 4762 -1398
rect 4674 -1585 4703 -1411
rect 4749 -1585 4762 -1411
rect 4674 -1598 4762 -1585
rect 4933 -1411 5021 -1398
rect 4933 -1585 4946 -1411
rect 4992 -1585 5021 -1411
rect 4933 -1598 5021 -1585
rect 5077 -1411 5165 -1398
rect 5077 -1585 5106 -1411
rect 5152 -1585 5165 -1411
rect 5077 -1598 5165 -1585
rect 5597 -1412 5685 -1399
rect 5597 -1586 5610 -1412
rect 5656 -1586 5685 -1412
rect -4845 -1755 -4757 -1742
rect -4845 -1929 -4832 -1755
rect -4786 -1929 -4757 -1755
rect -4845 -1942 -4757 -1929
rect -4701 -1755 -4613 -1742
rect -4701 -1929 -4672 -1755
rect -4626 -1929 -4613 -1755
rect -4701 -1942 -4613 -1929
rect -4441 -1755 -4353 -1742
rect -4441 -1929 -4428 -1755
rect -4382 -1929 -4353 -1755
rect -4441 -1942 -4353 -1929
rect -4297 -1755 -4209 -1742
rect -4297 -1929 -4268 -1755
rect -4222 -1929 -4209 -1755
rect -4297 -1942 -4209 -1929
rect -4038 -1755 -3950 -1742
rect -4038 -1929 -4025 -1755
rect -3979 -1929 -3950 -1755
rect -4038 -1942 -3950 -1929
rect -3894 -1755 -3790 -1742
rect -3894 -1929 -3865 -1755
rect -3819 -1929 -3790 -1755
rect -3894 -1942 -3790 -1929
rect -3734 -1755 -3630 -1742
rect -3734 -1929 -3705 -1755
rect -3659 -1929 -3630 -1755
rect -3734 -1942 -3630 -1929
rect -3574 -1755 -3470 -1742
rect -3574 -1929 -3545 -1755
rect -3499 -1929 -3470 -1755
rect -3574 -1942 -3470 -1929
rect -3414 -1755 -3310 -1742
rect -3414 -1929 -3385 -1755
rect -3339 -1929 -3310 -1755
rect -3414 -1942 -3310 -1929
rect -3254 -1755 -3150 -1742
rect -3254 -1929 -3225 -1755
rect -3179 -1929 -3150 -1755
rect -3254 -1942 -3150 -1929
rect -3094 -1755 -3006 -1742
rect -3094 -1929 -3065 -1755
rect -3019 -1929 -3006 -1755
rect -3094 -1942 -3006 -1929
rect -2442 -1748 -2354 -1735
rect -2442 -1922 -2429 -1748
rect -2383 -1922 -2354 -1748
rect -2442 -1935 -2354 -1922
rect -2298 -1748 -2210 -1735
rect -2298 -1922 -2269 -1748
rect -2223 -1922 -2210 -1748
rect -2298 -1935 -2210 -1922
rect -2038 -1748 -1950 -1735
rect -2038 -1922 -2025 -1748
rect -1979 -1922 -1950 -1748
rect -2038 -1935 -1950 -1922
rect -1894 -1748 -1806 -1735
rect -1894 -1922 -1865 -1748
rect -1819 -1922 -1806 -1748
rect -1894 -1935 -1806 -1922
rect -1635 -1748 -1547 -1735
rect -1635 -1922 -1622 -1748
rect -1576 -1922 -1547 -1748
rect -1635 -1935 -1547 -1922
rect -1491 -1748 -1387 -1735
rect -1491 -1922 -1462 -1748
rect -1416 -1922 -1387 -1748
rect -1491 -1935 -1387 -1922
rect -1331 -1748 -1227 -1735
rect -1331 -1922 -1302 -1748
rect -1256 -1922 -1227 -1748
rect -1331 -1935 -1227 -1922
rect -1171 -1748 -1067 -1735
rect -1171 -1922 -1142 -1748
rect -1096 -1922 -1067 -1748
rect -1171 -1935 -1067 -1922
rect -1011 -1748 -907 -1735
rect -1011 -1922 -982 -1748
rect -936 -1922 -907 -1748
rect -1011 -1935 -907 -1922
rect -851 -1748 -747 -1735
rect -851 -1922 -822 -1748
rect -776 -1922 -747 -1748
rect -851 -1935 -747 -1922
rect -691 -1748 -603 -1735
rect -691 -1922 -662 -1748
rect -616 -1922 -603 -1748
rect 5597 -1599 5685 -1586
rect 5741 -1412 5829 -1399
rect 5741 -1586 5770 -1412
rect 5816 -1586 5829 -1412
rect 5741 -1599 5829 -1586
rect 6000 -1412 6088 -1399
rect 6000 -1586 6013 -1412
rect 6059 -1586 6088 -1412
rect 6000 -1599 6088 -1586
rect 6144 -1412 6248 -1399
rect 6144 -1586 6173 -1412
rect 6219 -1586 6248 -1412
rect 6144 -1599 6248 -1586
rect 6304 -1412 6408 -1399
rect 6304 -1586 6333 -1412
rect 6379 -1586 6408 -1412
rect 6304 -1599 6408 -1586
rect 6464 -1412 6568 -1399
rect 6464 -1586 6493 -1412
rect 6539 -1586 6568 -1412
rect 6464 -1599 6568 -1586
rect 6624 -1412 6728 -1399
rect 6624 -1586 6653 -1412
rect 6699 -1586 6728 -1412
rect 6624 -1599 6728 -1586
rect 6784 -1412 6888 -1399
rect 6784 -1586 6813 -1412
rect 6859 -1586 6888 -1412
rect 6784 -1599 6888 -1586
rect 6944 -1412 7032 -1399
rect 6944 -1586 6973 -1412
rect 7019 -1586 7032 -1412
rect 6944 -1599 7032 -1586
rect 1917 -1747 2005 -1734
rect -691 -1935 -603 -1922
rect 1917 -1921 1930 -1747
rect 1976 -1921 2005 -1747
rect 1917 -1934 2005 -1921
rect 2061 -1747 2149 -1734
rect 2061 -1921 2090 -1747
rect 2136 -1921 2149 -1747
rect 2061 -1934 2149 -1921
rect 2320 -1747 2408 -1734
rect 2320 -1921 2333 -1747
rect 2379 -1921 2408 -1747
rect 2320 -1934 2408 -1921
rect 2464 -1747 2568 -1734
rect 2464 -1921 2493 -1747
rect 2539 -1921 2568 -1747
rect 2464 -1934 2568 -1921
rect 2624 -1747 2728 -1734
rect 2624 -1921 2653 -1747
rect 2699 -1921 2728 -1747
rect 2624 -1934 2728 -1921
rect 2784 -1747 2888 -1734
rect 2784 -1921 2813 -1747
rect 2859 -1921 2888 -1747
rect 2784 -1934 2888 -1921
rect 2944 -1747 3048 -1734
rect 2944 -1921 2973 -1747
rect 3019 -1921 3048 -1747
rect 2944 -1934 3048 -1921
rect 3104 -1747 3208 -1734
rect 3104 -1921 3133 -1747
rect 3179 -1921 3208 -1747
rect 3104 -1934 3208 -1921
rect 3264 -1747 3352 -1734
rect 3264 -1921 3293 -1747
rect 3339 -1921 3352 -1747
rect 3264 -1934 3352 -1921
rect 3730 -1747 3818 -1734
rect 3730 -1921 3743 -1747
rect 3789 -1921 3818 -1747
rect 3730 -1934 3818 -1921
rect 3874 -1747 3978 -1734
rect 3874 -1921 3903 -1747
rect 3949 -1921 3978 -1747
rect 3874 -1934 3978 -1921
rect 4034 -1747 4138 -1734
rect 4034 -1921 4063 -1747
rect 4109 -1921 4138 -1747
rect 4034 -1934 4138 -1921
rect 4194 -1747 4298 -1734
rect 4194 -1921 4223 -1747
rect 4269 -1921 4298 -1747
rect 4194 -1934 4298 -1921
rect 4354 -1747 4458 -1734
rect 4354 -1921 4383 -1747
rect 4429 -1921 4458 -1747
rect 4354 -1934 4458 -1921
rect 4514 -1747 4618 -1734
rect 4514 -1921 4543 -1747
rect 4589 -1921 4618 -1747
rect 4514 -1934 4618 -1921
rect 4674 -1747 4762 -1734
rect 4674 -1921 4703 -1747
rect 4749 -1921 4762 -1747
rect 4674 -1934 4762 -1921
rect 4933 -1747 5021 -1734
rect 4933 -1921 4946 -1747
rect 4992 -1921 5021 -1747
rect 4933 -1934 5021 -1921
rect 5077 -1747 5165 -1734
rect 5077 -1921 5106 -1747
rect 5152 -1921 5165 -1747
rect 5077 -1934 5165 -1921
rect 5597 -1748 5685 -1735
rect 5597 -1922 5610 -1748
rect 5656 -1922 5685 -1748
rect -4845 -2091 -4757 -2078
rect -4845 -2265 -4832 -2091
rect -4786 -2265 -4757 -2091
rect -4845 -2278 -4757 -2265
rect -4701 -2091 -4613 -2078
rect -4701 -2265 -4672 -2091
rect -4626 -2265 -4613 -2091
rect -4701 -2278 -4613 -2265
rect -4441 -2091 -4353 -2078
rect -4441 -2265 -4428 -2091
rect -4382 -2265 -4353 -2091
rect -4441 -2278 -4353 -2265
rect -4297 -2091 -4209 -2078
rect -4297 -2265 -4268 -2091
rect -4222 -2265 -4209 -2091
rect -4297 -2278 -4209 -2265
rect -4038 -2091 -3950 -2078
rect -4038 -2265 -4025 -2091
rect -3979 -2265 -3950 -2091
rect -4038 -2278 -3950 -2265
rect -3894 -2091 -3790 -2078
rect -3894 -2265 -3865 -2091
rect -3819 -2265 -3790 -2091
rect -3894 -2278 -3790 -2265
rect -3734 -2091 -3630 -2078
rect -3734 -2265 -3705 -2091
rect -3659 -2265 -3630 -2091
rect -3734 -2278 -3630 -2265
rect -3574 -2091 -3470 -2078
rect -3574 -2265 -3545 -2091
rect -3499 -2265 -3470 -2091
rect -3574 -2278 -3470 -2265
rect -3414 -2091 -3310 -2078
rect -3414 -2265 -3385 -2091
rect -3339 -2265 -3310 -2091
rect -3414 -2278 -3310 -2265
rect -3254 -2091 -3150 -2078
rect -3254 -2265 -3225 -2091
rect -3179 -2265 -3150 -2091
rect -3254 -2278 -3150 -2265
rect -3094 -2091 -3006 -2078
rect -3094 -2265 -3065 -2091
rect -3019 -2265 -3006 -2091
rect -3094 -2278 -3006 -2265
rect -2442 -2084 -2354 -2071
rect -2442 -2258 -2429 -2084
rect -2383 -2258 -2354 -2084
rect -2442 -2271 -2354 -2258
rect -2298 -2084 -2210 -2071
rect -2298 -2258 -2269 -2084
rect -2223 -2258 -2210 -2084
rect -2298 -2271 -2210 -2258
rect -2038 -2084 -1950 -2071
rect -2038 -2258 -2025 -2084
rect -1979 -2258 -1950 -2084
rect -2038 -2271 -1950 -2258
rect -1894 -2084 -1806 -2071
rect -1894 -2258 -1865 -2084
rect -1819 -2258 -1806 -2084
rect -1894 -2271 -1806 -2258
rect -1635 -2084 -1547 -2071
rect -1635 -2258 -1622 -2084
rect -1576 -2258 -1547 -2084
rect -1635 -2271 -1547 -2258
rect -1491 -2084 -1387 -2071
rect -1491 -2258 -1462 -2084
rect -1416 -2258 -1387 -2084
rect -1491 -2271 -1387 -2258
rect -1331 -2084 -1227 -2071
rect -1331 -2258 -1302 -2084
rect -1256 -2258 -1227 -2084
rect -1331 -2271 -1227 -2258
rect -1171 -2084 -1067 -2071
rect -1171 -2258 -1142 -2084
rect -1096 -2258 -1067 -2084
rect -1171 -2271 -1067 -2258
rect -1011 -2084 -907 -2071
rect -1011 -2258 -982 -2084
rect -936 -2258 -907 -2084
rect -1011 -2271 -907 -2258
rect -851 -2084 -747 -2071
rect -851 -2258 -822 -2084
rect -776 -2258 -747 -2084
rect -851 -2271 -747 -2258
rect -691 -2084 -603 -2071
rect -691 -2258 -662 -2084
rect -616 -2258 -603 -2084
rect 5597 -1935 5685 -1922
rect 5741 -1748 5829 -1735
rect 5741 -1922 5770 -1748
rect 5816 -1922 5829 -1748
rect 5741 -1935 5829 -1922
rect 6000 -1748 6088 -1735
rect 6000 -1922 6013 -1748
rect 6059 -1922 6088 -1748
rect 6000 -1935 6088 -1922
rect 6144 -1748 6248 -1735
rect 6144 -1922 6173 -1748
rect 6219 -1922 6248 -1748
rect 6144 -1935 6248 -1922
rect 6304 -1748 6408 -1735
rect 6304 -1922 6333 -1748
rect 6379 -1922 6408 -1748
rect 6304 -1935 6408 -1922
rect 6464 -1748 6568 -1735
rect 6464 -1922 6493 -1748
rect 6539 -1922 6568 -1748
rect 6464 -1935 6568 -1922
rect 6624 -1748 6728 -1735
rect 6624 -1922 6653 -1748
rect 6699 -1922 6728 -1748
rect 6624 -1935 6728 -1922
rect 6784 -1748 6888 -1735
rect 6784 -1922 6813 -1748
rect 6859 -1922 6888 -1748
rect 6784 -1935 6888 -1922
rect 6944 -1748 7032 -1735
rect 6944 -1922 6973 -1748
rect 7019 -1922 7032 -1748
rect 6944 -1935 7032 -1922
rect 1917 -2083 2005 -2070
rect -691 -2271 -603 -2258
rect 1917 -2257 1930 -2083
rect 1976 -2257 2005 -2083
rect 1917 -2270 2005 -2257
rect 2061 -2083 2149 -2070
rect 2061 -2257 2090 -2083
rect 2136 -2257 2149 -2083
rect 2061 -2270 2149 -2257
rect 2320 -2083 2408 -2070
rect 2320 -2257 2333 -2083
rect 2379 -2257 2408 -2083
rect 2320 -2270 2408 -2257
rect 2464 -2083 2568 -2070
rect 2464 -2257 2493 -2083
rect 2539 -2257 2568 -2083
rect 2464 -2270 2568 -2257
rect 2624 -2083 2728 -2070
rect 2624 -2257 2653 -2083
rect 2699 -2257 2728 -2083
rect 2624 -2270 2728 -2257
rect 2784 -2083 2888 -2070
rect 2784 -2257 2813 -2083
rect 2859 -2257 2888 -2083
rect 2784 -2270 2888 -2257
rect 2944 -2083 3048 -2070
rect 2944 -2257 2973 -2083
rect 3019 -2257 3048 -2083
rect 2944 -2270 3048 -2257
rect 3104 -2083 3208 -2070
rect 3104 -2257 3133 -2083
rect 3179 -2257 3208 -2083
rect 3104 -2270 3208 -2257
rect 3264 -2083 3352 -2070
rect 3264 -2257 3293 -2083
rect 3339 -2257 3352 -2083
rect 3264 -2270 3352 -2257
rect 3730 -2083 3818 -2070
rect 3730 -2257 3743 -2083
rect 3789 -2257 3818 -2083
rect 3730 -2270 3818 -2257
rect 3874 -2083 3978 -2070
rect 3874 -2257 3903 -2083
rect 3949 -2257 3978 -2083
rect 3874 -2270 3978 -2257
rect 4034 -2083 4138 -2070
rect 4034 -2257 4063 -2083
rect 4109 -2257 4138 -2083
rect 4034 -2270 4138 -2257
rect 4194 -2083 4298 -2070
rect 4194 -2257 4223 -2083
rect 4269 -2257 4298 -2083
rect 4194 -2270 4298 -2257
rect 4354 -2083 4458 -2070
rect 4354 -2257 4383 -2083
rect 4429 -2257 4458 -2083
rect 4354 -2270 4458 -2257
rect 4514 -2083 4618 -2070
rect 4514 -2257 4543 -2083
rect 4589 -2257 4618 -2083
rect 4514 -2270 4618 -2257
rect 4674 -2083 4762 -2070
rect 4674 -2257 4703 -2083
rect 4749 -2257 4762 -2083
rect 4674 -2270 4762 -2257
rect 4933 -2083 5021 -2070
rect 4933 -2257 4946 -2083
rect 4992 -2257 5021 -2083
rect 4933 -2270 5021 -2257
rect 5077 -2083 5165 -2070
rect 5077 -2257 5106 -2083
rect 5152 -2257 5165 -2083
rect 5077 -2270 5165 -2257
rect 5597 -2084 5685 -2071
rect 5597 -2258 5610 -2084
rect 5656 -2258 5685 -2084
rect 5597 -2271 5685 -2258
rect 5741 -2084 5829 -2071
rect 5741 -2258 5770 -2084
rect 5816 -2258 5829 -2084
rect 5741 -2271 5829 -2258
rect 6000 -2084 6088 -2071
rect 6000 -2258 6013 -2084
rect 6059 -2258 6088 -2084
rect 6000 -2271 6088 -2258
rect 6144 -2084 6248 -2071
rect 6144 -2258 6173 -2084
rect 6219 -2258 6248 -2084
rect 6144 -2271 6248 -2258
rect 6304 -2084 6408 -2071
rect 6304 -2258 6333 -2084
rect 6379 -2258 6408 -2084
rect 6304 -2271 6408 -2258
rect 6464 -2084 6568 -2071
rect 6464 -2258 6493 -2084
rect 6539 -2258 6568 -2084
rect 6464 -2271 6568 -2258
rect 6624 -2084 6728 -2071
rect 6624 -2258 6653 -2084
rect 6699 -2258 6728 -2084
rect 6624 -2271 6728 -2258
rect 6784 -2084 6888 -2071
rect 6784 -2258 6813 -2084
rect 6859 -2258 6888 -2084
rect 6784 -2271 6888 -2258
rect 6944 -2084 7032 -2071
rect 6944 -2258 6973 -2084
rect 7019 -2258 7032 -2084
rect 6944 -2271 7032 -2258
rect 147 -2354 235 -2341
rect 147 -2528 160 -2354
rect 206 -2528 235 -2354
rect 147 -2541 235 -2528
rect 291 -2354 395 -2341
rect 291 -2528 320 -2354
rect 366 -2528 395 -2354
rect 291 -2541 395 -2528
rect 451 -2354 555 -2341
rect 451 -2528 480 -2354
rect 526 -2528 555 -2354
rect 451 -2541 555 -2528
rect 611 -2354 715 -2341
rect 611 -2528 640 -2354
rect 686 -2528 715 -2354
rect 611 -2541 715 -2528
rect 771 -2354 859 -2341
rect 771 -2528 800 -2354
rect 846 -2528 859 -2354
rect 771 -2541 859 -2528
rect 147 -2690 235 -2677
rect -4845 -2747 -4757 -2734
rect -4845 -2921 -4832 -2747
rect -4786 -2921 -4757 -2747
rect -4845 -2934 -4757 -2921
rect -4701 -2747 -4613 -2734
rect -4701 -2921 -4672 -2747
rect -4626 -2921 -4613 -2747
rect -4701 -2934 -4613 -2921
rect -4441 -2747 -4353 -2734
rect -4441 -2921 -4428 -2747
rect -4382 -2921 -4353 -2747
rect -4441 -2934 -4353 -2921
rect -4297 -2747 -4209 -2734
rect -4297 -2921 -4268 -2747
rect -4222 -2921 -4209 -2747
rect -4297 -2934 -4209 -2921
rect -4038 -2747 -3950 -2734
rect -4038 -2921 -4025 -2747
rect -3979 -2921 -3950 -2747
rect -4038 -2934 -3950 -2921
rect -3894 -2747 -3790 -2734
rect -3894 -2921 -3865 -2747
rect -3819 -2921 -3790 -2747
rect -3894 -2934 -3790 -2921
rect -3734 -2747 -3630 -2734
rect -3734 -2921 -3705 -2747
rect -3659 -2921 -3630 -2747
rect -3734 -2934 -3630 -2921
rect -3574 -2747 -3470 -2734
rect -3574 -2921 -3545 -2747
rect -3499 -2921 -3470 -2747
rect -3574 -2934 -3470 -2921
rect -3414 -2747 -3310 -2734
rect -3414 -2921 -3385 -2747
rect -3339 -2921 -3310 -2747
rect -3414 -2934 -3310 -2921
rect -3254 -2747 -3150 -2734
rect -3254 -2921 -3225 -2747
rect -3179 -2921 -3150 -2747
rect -3254 -2934 -3150 -2921
rect -3094 -2747 -3006 -2734
rect -3094 -2921 -3065 -2747
rect -3019 -2921 -3006 -2747
rect -3094 -2934 -3006 -2921
rect -2442 -2740 -2354 -2727
rect -2442 -2914 -2429 -2740
rect -2383 -2914 -2354 -2740
rect -2442 -2927 -2354 -2914
rect -2298 -2740 -2210 -2727
rect -2298 -2914 -2269 -2740
rect -2223 -2914 -2210 -2740
rect -2298 -2927 -2210 -2914
rect -2038 -2740 -1950 -2727
rect -2038 -2914 -2025 -2740
rect -1979 -2914 -1950 -2740
rect -2038 -2927 -1950 -2914
rect -1894 -2740 -1806 -2727
rect -1894 -2914 -1865 -2740
rect -1819 -2914 -1806 -2740
rect -1894 -2927 -1806 -2914
rect -1635 -2740 -1547 -2727
rect -1635 -2914 -1622 -2740
rect -1576 -2914 -1547 -2740
rect -1635 -2927 -1547 -2914
rect -1491 -2740 -1387 -2727
rect -1491 -2914 -1462 -2740
rect -1416 -2914 -1387 -2740
rect -1491 -2927 -1387 -2914
rect -1331 -2740 -1227 -2727
rect -1331 -2914 -1302 -2740
rect -1256 -2914 -1227 -2740
rect -1331 -2927 -1227 -2914
rect -1171 -2740 -1067 -2727
rect -1171 -2914 -1142 -2740
rect -1096 -2914 -1067 -2740
rect -1171 -2927 -1067 -2914
rect -1011 -2740 -907 -2727
rect -1011 -2914 -982 -2740
rect -936 -2914 -907 -2740
rect -1011 -2927 -907 -2914
rect -851 -2740 -747 -2727
rect -851 -2914 -822 -2740
rect -776 -2914 -747 -2740
rect -851 -2927 -747 -2914
rect -691 -2740 -603 -2727
rect -691 -2914 -662 -2740
rect -616 -2914 -603 -2740
rect 147 -2864 160 -2690
rect 206 -2864 235 -2690
rect 147 -2877 235 -2864
rect 291 -2690 395 -2677
rect 291 -2864 320 -2690
rect 366 -2864 395 -2690
rect 291 -2877 395 -2864
rect 451 -2690 555 -2677
rect 451 -2864 480 -2690
rect 526 -2864 555 -2690
rect 451 -2877 555 -2864
rect 611 -2690 715 -2677
rect 611 -2864 640 -2690
rect 686 -2864 715 -2690
rect 611 -2877 715 -2864
rect 771 -2690 859 -2677
rect 771 -2864 800 -2690
rect 846 -2864 859 -2690
rect 771 -2877 859 -2864
rect 1917 -2739 2005 -2726
rect -691 -2927 -603 -2914
rect 1917 -2913 1930 -2739
rect 1976 -2913 2005 -2739
rect 1917 -2926 2005 -2913
rect 2061 -2739 2149 -2726
rect 2061 -2913 2090 -2739
rect 2136 -2913 2149 -2739
rect 2061 -2926 2149 -2913
rect 2320 -2739 2408 -2726
rect 2320 -2913 2333 -2739
rect 2379 -2913 2408 -2739
rect 2320 -2926 2408 -2913
rect 2464 -2739 2568 -2726
rect 2464 -2913 2493 -2739
rect 2539 -2913 2568 -2739
rect 2464 -2926 2568 -2913
rect 2624 -2739 2728 -2726
rect 2624 -2913 2653 -2739
rect 2699 -2913 2728 -2739
rect 2624 -2926 2728 -2913
rect 2784 -2739 2888 -2726
rect 2784 -2913 2813 -2739
rect 2859 -2913 2888 -2739
rect 2784 -2926 2888 -2913
rect 2944 -2739 3048 -2726
rect 2944 -2913 2973 -2739
rect 3019 -2913 3048 -2739
rect 2944 -2926 3048 -2913
rect 3104 -2739 3208 -2726
rect 3104 -2913 3133 -2739
rect 3179 -2913 3208 -2739
rect 3104 -2926 3208 -2913
rect 3264 -2739 3352 -2726
rect 3264 -2913 3293 -2739
rect 3339 -2913 3352 -2739
rect 3264 -2926 3352 -2913
rect 3730 -2739 3818 -2726
rect 3730 -2913 3743 -2739
rect 3789 -2913 3818 -2739
rect 3730 -2926 3818 -2913
rect 3874 -2739 3978 -2726
rect 3874 -2913 3903 -2739
rect 3949 -2913 3978 -2739
rect 3874 -2926 3978 -2913
rect 4034 -2739 4138 -2726
rect 4034 -2913 4063 -2739
rect 4109 -2913 4138 -2739
rect 4034 -2926 4138 -2913
rect 4194 -2739 4298 -2726
rect 4194 -2913 4223 -2739
rect 4269 -2913 4298 -2739
rect 4194 -2926 4298 -2913
rect 4354 -2739 4458 -2726
rect 4354 -2913 4383 -2739
rect 4429 -2913 4458 -2739
rect 4354 -2926 4458 -2913
rect 4514 -2739 4618 -2726
rect 4514 -2913 4543 -2739
rect 4589 -2913 4618 -2739
rect 4514 -2926 4618 -2913
rect 4674 -2739 4762 -2726
rect 4674 -2913 4703 -2739
rect 4749 -2913 4762 -2739
rect 4674 -2926 4762 -2913
rect 4933 -2739 5021 -2726
rect 4933 -2913 4946 -2739
rect 4992 -2913 5021 -2739
rect 4933 -2926 5021 -2913
rect 5077 -2739 5165 -2726
rect 5077 -2913 5106 -2739
rect 5152 -2913 5165 -2739
rect 5077 -2926 5165 -2913
rect 5597 -2740 5685 -2727
rect 5597 -2914 5610 -2740
rect 5656 -2914 5685 -2740
rect -4845 -3083 -4757 -3070
rect -4845 -3257 -4832 -3083
rect -4786 -3257 -4757 -3083
rect -4845 -3270 -4757 -3257
rect -4701 -3083 -4613 -3070
rect -4701 -3257 -4672 -3083
rect -4626 -3257 -4613 -3083
rect -4701 -3270 -4613 -3257
rect -4441 -3083 -4353 -3070
rect -4441 -3257 -4428 -3083
rect -4382 -3257 -4353 -3083
rect -4441 -3270 -4353 -3257
rect -4297 -3083 -4209 -3070
rect -4297 -3257 -4268 -3083
rect -4222 -3257 -4209 -3083
rect -4297 -3270 -4209 -3257
rect -4038 -3083 -3950 -3070
rect -4038 -3257 -4025 -3083
rect -3979 -3257 -3950 -3083
rect -4038 -3270 -3950 -3257
rect -3894 -3083 -3790 -3070
rect -3894 -3257 -3865 -3083
rect -3819 -3257 -3790 -3083
rect -3894 -3270 -3790 -3257
rect -3734 -3083 -3630 -3070
rect -3734 -3257 -3705 -3083
rect -3659 -3257 -3630 -3083
rect -3734 -3270 -3630 -3257
rect -3574 -3083 -3470 -3070
rect -3574 -3257 -3545 -3083
rect -3499 -3257 -3470 -3083
rect -3574 -3270 -3470 -3257
rect -3414 -3083 -3310 -3070
rect -3414 -3257 -3385 -3083
rect -3339 -3257 -3310 -3083
rect -3414 -3270 -3310 -3257
rect -3254 -3083 -3150 -3070
rect -3254 -3257 -3225 -3083
rect -3179 -3257 -3150 -3083
rect -3254 -3270 -3150 -3257
rect -3094 -3083 -3006 -3070
rect -3094 -3257 -3065 -3083
rect -3019 -3257 -3006 -3083
rect -3094 -3270 -3006 -3257
rect -2442 -3076 -2354 -3063
rect -2442 -3250 -2429 -3076
rect -2383 -3250 -2354 -3076
rect -2442 -3263 -2354 -3250
rect -2298 -3076 -2210 -3063
rect -2298 -3250 -2269 -3076
rect -2223 -3250 -2210 -3076
rect -2298 -3263 -2210 -3250
rect -2038 -3076 -1950 -3063
rect -2038 -3250 -2025 -3076
rect -1979 -3250 -1950 -3076
rect -2038 -3263 -1950 -3250
rect -1894 -3076 -1806 -3063
rect -1894 -3250 -1865 -3076
rect -1819 -3250 -1806 -3076
rect -1894 -3263 -1806 -3250
rect -1635 -3076 -1547 -3063
rect -1635 -3250 -1622 -3076
rect -1576 -3250 -1547 -3076
rect -1635 -3263 -1547 -3250
rect -1491 -3076 -1387 -3063
rect -1491 -3250 -1462 -3076
rect -1416 -3250 -1387 -3076
rect -1491 -3263 -1387 -3250
rect -1331 -3076 -1227 -3063
rect -1331 -3250 -1302 -3076
rect -1256 -3250 -1227 -3076
rect -1331 -3263 -1227 -3250
rect -1171 -3076 -1067 -3063
rect -1171 -3250 -1142 -3076
rect -1096 -3250 -1067 -3076
rect -1171 -3263 -1067 -3250
rect -1011 -3076 -907 -3063
rect -1011 -3250 -982 -3076
rect -936 -3250 -907 -3076
rect -1011 -3263 -907 -3250
rect -851 -3076 -747 -3063
rect -851 -3250 -822 -3076
rect -776 -3250 -747 -3076
rect -851 -3263 -747 -3250
rect -691 -3076 -603 -3063
rect -691 -3250 -662 -3076
rect -616 -3250 -603 -3076
rect 5597 -2927 5685 -2914
rect 5741 -2740 5829 -2727
rect 5741 -2914 5770 -2740
rect 5816 -2914 5829 -2740
rect 5741 -2927 5829 -2914
rect 6000 -2740 6088 -2727
rect 6000 -2914 6013 -2740
rect 6059 -2914 6088 -2740
rect 6000 -2927 6088 -2914
rect 6144 -2740 6248 -2727
rect 6144 -2914 6173 -2740
rect 6219 -2914 6248 -2740
rect 6144 -2927 6248 -2914
rect 6304 -2740 6408 -2727
rect 6304 -2914 6333 -2740
rect 6379 -2914 6408 -2740
rect 6304 -2927 6408 -2914
rect 6464 -2740 6568 -2727
rect 6464 -2914 6493 -2740
rect 6539 -2914 6568 -2740
rect 6464 -2927 6568 -2914
rect 6624 -2740 6728 -2727
rect 6624 -2914 6653 -2740
rect 6699 -2914 6728 -2740
rect 6624 -2927 6728 -2914
rect 6784 -2740 6888 -2727
rect 6784 -2914 6813 -2740
rect 6859 -2914 6888 -2740
rect 6784 -2927 6888 -2914
rect 6944 -2740 7032 -2727
rect 6944 -2914 6973 -2740
rect 7019 -2914 7032 -2740
rect 6944 -2927 7032 -2914
rect 1917 -3075 2005 -3062
rect -691 -3263 -603 -3250
rect 1917 -3249 1930 -3075
rect 1976 -3249 2005 -3075
rect 1917 -3262 2005 -3249
rect 2061 -3075 2149 -3062
rect 2061 -3249 2090 -3075
rect 2136 -3249 2149 -3075
rect 2061 -3262 2149 -3249
rect 2320 -3075 2408 -3062
rect 2320 -3249 2333 -3075
rect 2379 -3249 2408 -3075
rect 2320 -3262 2408 -3249
rect 2464 -3075 2568 -3062
rect 2464 -3249 2493 -3075
rect 2539 -3249 2568 -3075
rect 2464 -3262 2568 -3249
rect 2624 -3075 2728 -3062
rect 2624 -3249 2653 -3075
rect 2699 -3249 2728 -3075
rect 2624 -3262 2728 -3249
rect 2784 -3075 2888 -3062
rect 2784 -3249 2813 -3075
rect 2859 -3249 2888 -3075
rect 2784 -3262 2888 -3249
rect 2944 -3075 3048 -3062
rect 2944 -3249 2973 -3075
rect 3019 -3249 3048 -3075
rect 2944 -3262 3048 -3249
rect 3104 -3075 3208 -3062
rect 3104 -3249 3133 -3075
rect 3179 -3249 3208 -3075
rect 3104 -3262 3208 -3249
rect 3264 -3075 3352 -3062
rect 3264 -3249 3293 -3075
rect 3339 -3249 3352 -3075
rect 3264 -3262 3352 -3249
rect 3730 -3075 3818 -3062
rect 3730 -3249 3743 -3075
rect 3789 -3249 3818 -3075
rect 3730 -3262 3818 -3249
rect 3874 -3075 3978 -3062
rect 3874 -3249 3903 -3075
rect 3949 -3249 3978 -3075
rect 3874 -3262 3978 -3249
rect 4034 -3075 4138 -3062
rect 4034 -3249 4063 -3075
rect 4109 -3249 4138 -3075
rect 4034 -3262 4138 -3249
rect 4194 -3075 4298 -3062
rect 4194 -3249 4223 -3075
rect 4269 -3249 4298 -3075
rect 4194 -3262 4298 -3249
rect 4354 -3075 4458 -3062
rect 4354 -3249 4383 -3075
rect 4429 -3249 4458 -3075
rect 4354 -3262 4458 -3249
rect 4514 -3075 4618 -3062
rect 4514 -3249 4543 -3075
rect 4589 -3249 4618 -3075
rect 4514 -3262 4618 -3249
rect 4674 -3075 4762 -3062
rect 4674 -3249 4703 -3075
rect 4749 -3249 4762 -3075
rect 4674 -3262 4762 -3249
rect 4933 -3075 5021 -3062
rect 4933 -3249 4946 -3075
rect 4992 -3249 5021 -3075
rect 4933 -3262 5021 -3249
rect 5077 -3075 5165 -3062
rect 5077 -3249 5106 -3075
rect 5152 -3249 5165 -3075
rect 5077 -3262 5165 -3249
rect 5597 -3076 5685 -3063
rect 5597 -3250 5610 -3076
rect 5656 -3250 5685 -3076
rect 147 -3284 235 -3271
rect -4845 -3419 -4757 -3406
rect -4845 -3593 -4832 -3419
rect -4786 -3593 -4757 -3419
rect -4845 -3606 -4757 -3593
rect -4701 -3419 -4613 -3406
rect -4701 -3593 -4672 -3419
rect -4626 -3593 -4613 -3419
rect -4701 -3606 -4613 -3593
rect -4441 -3419 -4353 -3406
rect -4441 -3593 -4428 -3419
rect -4382 -3593 -4353 -3419
rect -4441 -3606 -4353 -3593
rect -4297 -3419 -4209 -3406
rect -4297 -3593 -4268 -3419
rect -4222 -3593 -4209 -3419
rect -4297 -3606 -4209 -3593
rect -4038 -3419 -3950 -3406
rect -4038 -3593 -4025 -3419
rect -3979 -3593 -3950 -3419
rect -4038 -3606 -3950 -3593
rect -3894 -3419 -3790 -3406
rect -3894 -3593 -3865 -3419
rect -3819 -3593 -3790 -3419
rect -3894 -3606 -3790 -3593
rect -3734 -3419 -3630 -3406
rect -3734 -3593 -3705 -3419
rect -3659 -3593 -3630 -3419
rect -3734 -3606 -3630 -3593
rect -3574 -3419 -3470 -3406
rect -3574 -3593 -3545 -3419
rect -3499 -3593 -3470 -3419
rect -3574 -3606 -3470 -3593
rect -3414 -3419 -3310 -3406
rect -3414 -3593 -3385 -3419
rect -3339 -3593 -3310 -3419
rect -3414 -3606 -3310 -3593
rect -3254 -3419 -3150 -3406
rect -3254 -3593 -3225 -3419
rect -3179 -3593 -3150 -3419
rect -3254 -3606 -3150 -3593
rect -3094 -3419 -3006 -3406
rect -3094 -3593 -3065 -3419
rect -3019 -3593 -3006 -3419
rect -3094 -3606 -3006 -3593
rect -2442 -3412 -2354 -3399
rect -2442 -3586 -2429 -3412
rect -2383 -3586 -2354 -3412
rect -2442 -3599 -2354 -3586
rect -2298 -3412 -2210 -3399
rect -2298 -3586 -2269 -3412
rect -2223 -3586 -2210 -3412
rect -2298 -3599 -2210 -3586
rect -2038 -3412 -1950 -3399
rect -2038 -3586 -2025 -3412
rect -1979 -3586 -1950 -3412
rect -2038 -3599 -1950 -3586
rect -1894 -3412 -1806 -3399
rect -1894 -3586 -1865 -3412
rect -1819 -3586 -1806 -3412
rect -1894 -3599 -1806 -3586
rect -1635 -3412 -1547 -3399
rect -1635 -3586 -1622 -3412
rect -1576 -3586 -1547 -3412
rect -1635 -3599 -1547 -3586
rect -1491 -3412 -1387 -3399
rect -1491 -3586 -1462 -3412
rect -1416 -3586 -1387 -3412
rect -1491 -3599 -1387 -3586
rect -1331 -3412 -1227 -3399
rect -1331 -3586 -1302 -3412
rect -1256 -3586 -1227 -3412
rect -1331 -3599 -1227 -3586
rect -1171 -3412 -1067 -3399
rect -1171 -3586 -1142 -3412
rect -1096 -3586 -1067 -3412
rect -1171 -3599 -1067 -3586
rect -1011 -3412 -907 -3399
rect -1011 -3586 -982 -3412
rect -936 -3586 -907 -3412
rect -1011 -3599 -907 -3586
rect -851 -3412 -747 -3399
rect -851 -3586 -822 -3412
rect -776 -3586 -747 -3412
rect -851 -3599 -747 -3586
rect -691 -3412 -603 -3399
rect -691 -3586 -662 -3412
rect -616 -3586 -603 -3412
rect 147 -3458 160 -3284
rect 206 -3458 235 -3284
rect 147 -3471 235 -3458
rect 291 -3284 395 -3271
rect 291 -3458 320 -3284
rect 366 -3458 395 -3284
rect 291 -3471 395 -3458
rect 451 -3284 555 -3271
rect 451 -3458 480 -3284
rect 526 -3458 555 -3284
rect 451 -3471 555 -3458
rect 611 -3284 715 -3271
rect 611 -3458 640 -3284
rect 686 -3458 715 -3284
rect 611 -3471 715 -3458
rect 771 -3284 859 -3271
rect 771 -3458 800 -3284
rect 846 -3458 859 -3284
rect 5597 -3263 5685 -3250
rect 5741 -3076 5829 -3063
rect 5741 -3250 5770 -3076
rect 5816 -3250 5829 -3076
rect 5741 -3263 5829 -3250
rect 6000 -3076 6088 -3063
rect 6000 -3250 6013 -3076
rect 6059 -3250 6088 -3076
rect 6000 -3263 6088 -3250
rect 6144 -3076 6248 -3063
rect 6144 -3250 6173 -3076
rect 6219 -3250 6248 -3076
rect 6144 -3263 6248 -3250
rect 6304 -3076 6408 -3063
rect 6304 -3250 6333 -3076
rect 6379 -3250 6408 -3076
rect 6304 -3263 6408 -3250
rect 6464 -3076 6568 -3063
rect 6464 -3250 6493 -3076
rect 6539 -3250 6568 -3076
rect 6464 -3263 6568 -3250
rect 6624 -3076 6728 -3063
rect 6624 -3250 6653 -3076
rect 6699 -3250 6728 -3076
rect 6624 -3263 6728 -3250
rect 6784 -3076 6888 -3063
rect 6784 -3250 6813 -3076
rect 6859 -3250 6888 -3076
rect 6784 -3263 6888 -3250
rect 6944 -3076 7032 -3063
rect 6944 -3250 6973 -3076
rect 7019 -3250 7032 -3076
rect 6944 -3263 7032 -3250
rect 771 -3471 859 -3458
rect 1917 -3411 2005 -3398
rect -691 -3599 -603 -3586
rect 1917 -3585 1930 -3411
rect 1976 -3585 2005 -3411
rect 1917 -3598 2005 -3585
rect 2061 -3411 2149 -3398
rect 2061 -3585 2090 -3411
rect 2136 -3585 2149 -3411
rect 2061 -3598 2149 -3585
rect 2320 -3411 2408 -3398
rect 2320 -3585 2333 -3411
rect 2379 -3585 2408 -3411
rect 2320 -3598 2408 -3585
rect 2464 -3411 2568 -3398
rect 2464 -3585 2493 -3411
rect 2539 -3585 2568 -3411
rect 2464 -3598 2568 -3585
rect 2624 -3411 2728 -3398
rect 2624 -3585 2653 -3411
rect 2699 -3585 2728 -3411
rect 2624 -3598 2728 -3585
rect 2784 -3411 2888 -3398
rect 2784 -3585 2813 -3411
rect 2859 -3585 2888 -3411
rect 2784 -3598 2888 -3585
rect 2944 -3411 3048 -3398
rect 2944 -3585 2973 -3411
rect 3019 -3585 3048 -3411
rect 2944 -3598 3048 -3585
rect 3104 -3411 3208 -3398
rect 3104 -3585 3133 -3411
rect 3179 -3585 3208 -3411
rect 3104 -3598 3208 -3585
rect 3264 -3411 3352 -3398
rect 3264 -3585 3293 -3411
rect 3339 -3585 3352 -3411
rect 3264 -3598 3352 -3585
rect 3730 -3411 3818 -3398
rect 3730 -3585 3743 -3411
rect 3789 -3585 3818 -3411
rect 3730 -3598 3818 -3585
rect 3874 -3411 3978 -3398
rect 3874 -3585 3903 -3411
rect 3949 -3585 3978 -3411
rect 3874 -3598 3978 -3585
rect 4034 -3411 4138 -3398
rect 4034 -3585 4063 -3411
rect 4109 -3585 4138 -3411
rect 4034 -3598 4138 -3585
rect 4194 -3411 4298 -3398
rect 4194 -3585 4223 -3411
rect 4269 -3585 4298 -3411
rect 4194 -3598 4298 -3585
rect 4354 -3411 4458 -3398
rect 4354 -3585 4383 -3411
rect 4429 -3585 4458 -3411
rect 4354 -3598 4458 -3585
rect 4514 -3411 4618 -3398
rect 4514 -3585 4543 -3411
rect 4589 -3585 4618 -3411
rect 4514 -3598 4618 -3585
rect 4674 -3411 4762 -3398
rect 4674 -3585 4703 -3411
rect 4749 -3585 4762 -3411
rect 4674 -3598 4762 -3585
rect 4933 -3411 5021 -3398
rect 4933 -3585 4946 -3411
rect 4992 -3585 5021 -3411
rect 4933 -3598 5021 -3585
rect 5077 -3411 5165 -3398
rect 5077 -3585 5106 -3411
rect 5152 -3585 5165 -3411
rect 5077 -3598 5165 -3585
rect 5597 -3412 5685 -3399
rect 5597 -3586 5610 -3412
rect 5656 -3586 5685 -3412
rect 147 -3620 235 -3607
rect -4845 -3755 -4757 -3742
rect -4845 -3929 -4832 -3755
rect -4786 -3929 -4757 -3755
rect -4845 -3942 -4757 -3929
rect -4701 -3755 -4613 -3742
rect -4701 -3929 -4672 -3755
rect -4626 -3929 -4613 -3755
rect -4701 -3942 -4613 -3929
rect -4441 -3755 -4353 -3742
rect -4441 -3929 -4428 -3755
rect -4382 -3929 -4353 -3755
rect -4441 -3942 -4353 -3929
rect -4297 -3755 -4209 -3742
rect -4297 -3929 -4268 -3755
rect -4222 -3929 -4209 -3755
rect -4297 -3942 -4209 -3929
rect -4038 -3755 -3950 -3742
rect -4038 -3929 -4025 -3755
rect -3979 -3929 -3950 -3755
rect -4038 -3942 -3950 -3929
rect -3894 -3755 -3790 -3742
rect -3894 -3929 -3865 -3755
rect -3819 -3929 -3790 -3755
rect -3894 -3942 -3790 -3929
rect -3734 -3755 -3630 -3742
rect -3734 -3929 -3705 -3755
rect -3659 -3929 -3630 -3755
rect -3734 -3942 -3630 -3929
rect -3574 -3755 -3470 -3742
rect -3574 -3929 -3545 -3755
rect -3499 -3929 -3470 -3755
rect -3574 -3942 -3470 -3929
rect -3414 -3755 -3310 -3742
rect -3414 -3929 -3385 -3755
rect -3339 -3929 -3310 -3755
rect -3414 -3942 -3310 -3929
rect -3254 -3755 -3150 -3742
rect -3254 -3929 -3225 -3755
rect -3179 -3929 -3150 -3755
rect -3254 -3942 -3150 -3929
rect -3094 -3755 -3006 -3742
rect -3094 -3929 -3065 -3755
rect -3019 -3929 -3006 -3755
rect -3094 -3942 -3006 -3929
rect -2442 -3748 -2354 -3735
rect -2442 -3922 -2429 -3748
rect -2383 -3922 -2354 -3748
rect -2442 -3935 -2354 -3922
rect -2298 -3748 -2210 -3735
rect -2298 -3922 -2269 -3748
rect -2223 -3922 -2210 -3748
rect -2298 -3935 -2210 -3922
rect -2038 -3748 -1950 -3735
rect -2038 -3922 -2025 -3748
rect -1979 -3922 -1950 -3748
rect -2038 -3935 -1950 -3922
rect -1894 -3748 -1806 -3735
rect -1894 -3922 -1865 -3748
rect -1819 -3922 -1806 -3748
rect -1894 -3935 -1806 -3922
rect -1635 -3748 -1547 -3735
rect -1635 -3922 -1622 -3748
rect -1576 -3922 -1547 -3748
rect -1635 -3935 -1547 -3922
rect -1491 -3748 -1387 -3735
rect -1491 -3922 -1462 -3748
rect -1416 -3922 -1387 -3748
rect -1491 -3935 -1387 -3922
rect -1331 -3748 -1227 -3735
rect -1331 -3922 -1302 -3748
rect -1256 -3922 -1227 -3748
rect -1331 -3935 -1227 -3922
rect -1171 -3748 -1067 -3735
rect -1171 -3922 -1142 -3748
rect -1096 -3922 -1067 -3748
rect -1171 -3935 -1067 -3922
rect -1011 -3748 -907 -3735
rect -1011 -3922 -982 -3748
rect -936 -3922 -907 -3748
rect -1011 -3935 -907 -3922
rect -851 -3748 -747 -3735
rect -851 -3922 -822 -3748
rect -776 -3922 -747 -3748
rect -851 -3935 -747 -3922
rect -691 -3748 -603 -3735
rect -691 -3922 -662 -3748
rect -616 -3922 -603 -3748
rect 147 -3794 160 -3620
rect 206 -3794 235 -3620
rect 147 -3807 235 -3794
rect 291 -3620 395 -3607
rect 291 -3794 320 -3620
rect 366 -3794 395 -3620
rect 291 -3807 395 -3794
rect 451 -3620 555 -3607
rect 451 -3794 480 -3620
rect 526 -3794 555 -3620
rect 451 -3807 555 -3794
rect 611 -3620 715 -3607
rect 611 -3794 640 -3620
rect 686 -3794 715 -3620
rect 611 -3807 715 -3794
rect 771 -3620 859 -3607
rect 771 -3794 800 -3620
rect 846 -3794 859 -3620
rect 5597 -3599 5685 -3586
rect 5741 -3412 5829 -3399
rect 5741 -3586 5770 -3412
rect 5816 -3586 5829 -3412
rect 5741 -3599 5829 -3586
rect 6000 -3412 6088 -3399
rect 6000 -3586 6013 -3412
rect 6059 -3586 6088 -3412
rect 6000 -3599 6088 -3586
rect 6144 -3412 6248 -3399
rect 6144 -3586 6173 -3412
rect 6219 -3586 6248 -3412
rect 6144 -3599 6248 -3586
rect 6304 -3412 6408 -3399
rect 6304 -3586 6333 -3412
rect 6379 -3586 6408 -3412
rect 6304 -3599 6408 -3586
rect 6464 -3412 6568 -3399
rect 6464 -3586 6493 -3412
rect 6539 -3586 6568 -3412
rect 6464 -3599 6568 -3586
rect 6624 -3412 6728 -3399
rect 6624 -3586 6653 -3412
rect 6699 -3586 6728 -3412
rect 6624 -3599 6728 -3586
rect 6784 -3412 6888 -3399
rect 6784 -3586 6813 -3412
rect 6859 -3586 6888 -3412
rect 6784 -3599 6888 -3586
rect 6944 -3412 7032 -3399
rect 6944 -3586 6973 -3412
rect 7019 -3586 7032 -3412
rect 6944 -3599 7032 -3586
rect 771 -3807 859 -3794
rect 1917 -3747 2005 -3734
rect -691 -3935 -603 -3922
rect 1917 -3921 1930 -3747
rect 1976 -3921 2005 -3747
rect 1917 -3934 2005 -3921
rect 2061 -3747 2149 -3734
rect 2061 -3921 2090 -3747
rect 2136 -3921 2149 -3747
rect 2061 -3934 2149 -3921
rect 2320 -3747 2408 -3734
rect 2320 -3921 2333 -3747
rect 2379 -3921 2408 -3747
rect 2320 -3934 2408 -3921
rect 2464 -3747 2568 -3734
rect 2464 -3921 2493 -3747
rect 2539 -3921 2568 -3747
rect 2464 -3934 2568 -3921
rect 2624 -3747 2728 -3734
rect 2624 -3921 2653 -3747
rect 2699 -3921 2728 -3747
rect 2624 -3934 2728 -3921
rect 2784 -3747 2888 -3734
rect 2784 -3921 2813 -3747
rect 2859 -3921 2888 -3747
rect 2784 -3934 2888 -3921
rect 2944 -3747 3048 -3734
rect 2944 -3921 2973 -3747
rect 3019 -3921 3048 -3747
rect 2944 -3934 3048 -3921
rect 3104 -3747 3208 -3734
rect 3104 -3921 3133 -3747
rect 3179 -3921 3208 -3747
rect 3104 -3934 3208 -3921
rect 3264 -3747 3352 -3734
rect 3264 -3921 3293 -3747
rect 3339 -3921 3352 -3747
rect 3264 -3934 3352 -3921
rect 3730 -3747 3818 -3734
rect 3730 -3921 3743 -3747
rect 3789 -3921 3818 -3747
rect 3730 -3934 3818 -3921
rect 3874 -3747 3978 -3734
rect 3874 -3921 3903 -3747
rect 3949 -3921 3978 -3747
rect 3874 -3934 3978 -3921
rect 4034 -3747 4138 -3734
rect 4034 -3921 4063 -3747
rect 4109 -3921 4138 -3747
rect 4034 -3934 4138 -3921
rect 4194 -3747 4298 -3734
rect 4194 -3921 4223 -3747
rect 4269 -3921 4298 -3747
rect 4194 -3934 4298 -3921
rect 4354 -3747 4458 -3734
rect 4354 -3921 4383 -3747
rect 4429 -3921 4458 -3747
rect 4354 -3934 4458 -3921
rect 4514 -3747 4618 -3734
rect 4514 -3921 4543 -3747
rect 4589 -3921 4618 -3747
rect 4514 -3934 4618 -3921
rect 4674 -3747 4762 -3734
rect 4674 -3921 4703 -3747
rect 4749 -3921 4762 -3747
rect 4674 -3934 4762 -3921
rect 4933 -3747 5021 -3734
rect 4933 -3921 4946 -3747
rect 4992 -3921 5021 -3747
rect 4933 -3934 5021 -3921
rect 5077 -3747 5165 -3734
rect 5077 -3921 5106 -3747
rect 5152 -3921 5165 -3747
rect 5077 -3934 5165 -3921
rect 5597 -3748 5685 -3735
rect 5597 -3922 5610 -3748
rect 5656 -3922 5685 -3748
rect 5597 -3935 5685 -3922
rect 5741 -3748 5829 -3735
rect 5741 -3922 5770 -3748
rect 5816 -3922 5829 -3748
rect 5741 -3935 5829 -3922
rect 6000 -3748 6088 -3735
rect 6000 -3922 6013 -3748
rect 6059 -3922 6088 -3748
rect 6000 -3935 6088 -3922
rect 6144 -3748 6248 -3735
rect 6144 -3922 6173 -3748
rect 6219 -3922 6248 -3748
rect 6144 -3935 6248 -3922
rect 6304 -3748 6408 -3735
rect 6304 -3922 6333 -3748
rect 6379 -3922 6408 -3748
rect 6304 -3935 6408 -3922
rect 6464 -3748 6568 -3735
rect 6464 -3922 6493 -3748
rect 6539 -3922 6568 -3748
rect 6464 -3935 6568 -3922
rect 6624 -3748 6728 -3735
rect 6624 -3922 6653 -3748
rect 6699 -3922 6728 -3748
rect 6624 -3935 6728 -3922
rect 6784 -3748 6888 -3735
rect 6784 -3922 6813 -3748
rect 6859 -3922 6888 -3748
rect 6784 -3935 6888 -3922
rect 6944 -3748 7032 -3735
rect 6944 -3922 6973 -3748
rect 7019 -3922 7032 -3748
rect 6944 -3935 7032 -3922
rect -4845 -6243 -4757 -6230
rect -4845 -6417 -4832 -6243
rect -4786 -6417 -4757 -6243
rect -4845 -6430 -4757 -6417
rect -4701 -6243 -4613 -6230
rect -4701 -6417 -4672 -6243
rect -4626 -6417 -4613 -6243
rect -4701 -6430 -4613 -6417
rect -4441 -6243 -4353 -6230
rect -4441 -6417 -4428 -6243
rect -4382 -6417 -4353 -6243
rect -4441 -6430 -4353 -6417
rect -4297 -6243 -4209 -6230
rect -4297 -6417 -4268 -6243
rect -4222 -6417 -4209 -6243
rect -4297 -6430 -4209 -6417
rect -4038 -6243 -3950 -6230
rect -4038 -6417 -4025 -6243
rect -3979 -6417 -3950 -6243
rect -4038 -6430 -3950 -6417
rect -3894 -6243 -3790 -6230
rect -3894 -6417 -3865 -6243
rect -3819 -6417 -3790 -6243
rect -3894 -6430 -3790 -6417
rect -3734 -6243 -3630 -6230
rect -3734 -6417 -3705 -6243
rect -3659 -6417 -3630 -6243
rect -3734 -6430 -3630 -6417
rect -3574 -6243 -3470 -6230
rect -3574 -6417 -3545 -6243
rect -3499 -6417 -3470 -6243
rect -3574 -6430 -3470 -6417
rect -3414 -6243 -3310 -6230
rect -3414 -6417 -3385 -6243
rect -3339 -6417 -3310 -6243
rect -3414 -6430 -3310 -6417
rect -3254 -6243 -3150 -6230
rect -3254 -6417 -3225 -6243
rect -3179 -6417 -3150 -6243
rect -3254 -6430 -3150 -6417
rect -3094 -6243 -3006 -6230
rect -3094 -6417 -3065 -6243
rect -3019 -6417 -3006 -6243
rect -3094 -6430 -3006 -6417
rect -2442 -6236 -2354 -6223
rect -2442 -6410 -2429 -6236
rect -2383 -6410 -2354 -6236
rect -2442 -6423 -2354 -6410
rect -2298 -6236 -2210 -6223
rect -2298 -6410 -2269 -6236
rect -2223 -6410 -2210 -6236
rect -2298 -6423 -2210 -6410
rect -2038 -6236 -1950 -6223
rect -2038 -6410 -2025 -6236
rect -1979 -6410 -1950 -6236
rect -2038 -6423 -1950 -6410
rect -1894 -6236 -1806 -6223
rect -1894 -6410 -1865 -6236
rect -1819 -6410 -1806 -6236
rect -1894 -6423 -1806 -6410
rect -1635 -6236 -1547 -6223
rect -1635 -6410 -1622 -6236
rect -1576 -6410 -1547 -6236
rect -1635 -6423 -1547 -6410
rect -1491 -6236 -1387 -6223
rect -1491 -6410 -1462 -6236
rect -1416 -6410 -1387 -6236
rect -1491 -6423 -1387 -6410
rect -1331 -6236 -1227 -6223
rect -1331 -6410 -1302 -6236
rect -1256 -6410 -1227 -6236
rect -1331 -6423 -1227 -6410
rect -1171 -6236 -1067 -6223
rect -1171 -6410 -1142 -6236
rect -1096 -6410 -1067 -6236
rect -1171 -6423 -1067 -6410
rect -1011 -6236 -907 -6223
rect -1011 -6410 -982 -6236
rect -936 -6410 -907 -6236
rect -1011 -6423 -907 -6410
rect -851 -6236 -747 -6223
rect -851 -6410 -822 -6236
rect -776 -6410 -747 -6236
rect -851 -6423 -747 -6410
rect -691 -6236 -603 -6223
rect -691 -6410 -662 -6236
rect -616 -6410 -603 -6236
rect -691 -6423 -603 -6410
rect 157 -6235 245 -6222
rect 157 -6409 170 -6235
rect 216 -6409 245 -6235
rect 157 -6422 245 -6409
rect 301 -6235 389 -6222
rect 301 -6409 330 -6235
rect 376 -6409 389 -6235
rect 301 -6422 389 -6409
rect 560 -6235 648 -6222
rect 560 -6409 573 -6235
rect 619 -6409 648 -6235
rect 560 -6422 648 -6409
rect 704 -6235 808 -6222
rect 704 -6409 733 -6235
rect 779 -6409 808 -6235
rect 704 -6422 808 -6409
rect 864 -6235 968 -6222
rect 864 -6409 893 -6235
rect 939 -6409 968 -6235
rect 864 -6422 968 -6409
rect 1024 -6235 1128 -6222
rect 1024 -6409 1053 -6235
rect 1099 -6409 1128 -6235
rect 1024 -6422 1128 -6409
rect 1184 -6235 1288 -6222
rect 1184 -6409 1213 -6235
rect 1259 -6409 1288 -6235
rect 1184 -6422 1288 -6409
rect 1344 -6235 1448 -6222
rect 1344 -6409 1373 -6235
rect 1419 -6409 1448 -6235
rect 1344 -6422 1448 -6409
rect 1504 -6235 1592 -6222
rect 1504 -6409 1533 -6235
rect 1579 -6409 1592 -6235
rect 1504 -6422 1592 -6409
rect 1917 -6235 2005 -6222
rect 1917 -6409 1930 -6235
rect 1976 -6409 2005 -6235
rect 1917 -6422 2005 -6409
rect 2061 -6235 2165 -6222
rect 2061 -6409 2090 -6235
rect 2136 -6409 2165 -6235
rect 2061 -6422 2165 -6409
rect 2221 -6235 2325 -6222
rect 2221 -6409 2250 -6235
rect 2296 -6409 2325 -6235
rect 2221 -6422 2325 -6409
rect 2381 -6235 2485 -6222
rect 2381 -6409 2410 -6235
rect 2456 -6409 2485 -6235
rect 2381 -6422 2485 -6409
rect 2541 -6235 2645 -6222
rect 2541 -6409 2570 -6235
rect 2616 -6409 2645 -6235
rect 2541 -6422 2645 -6409
rect 2701 -6235 2805 -6222
rect 2701 -6409 2730 -6235
rect 2776 -6409 2805 -6235
rect 2701 -6422 2805 -6409
rect 2861 -6235 2949 -6222
rect 2861 -6409 2890 -6235
rect 2936 -6409 2949 -6235
rect 2861 -6422 2949 -6409
rect 3120 -6235 3208 -6222
rect 3120 -6409 3133 -6235
rect 3179 -6409 3208 -6235
rect 3120 -6422 3208 -6409
rect 3264 -6235 3352 -6222
rect 3264 -6409 3293 -6235
rect 3339 -6409 3352 -6235
rect 3264 -6422 3352 -6409
rect 3730 -6235 3818 -6222
rect 3730 -6409 3743 -6235
rect 3789 -6409 3818 -6235
rect 3730 -6422 3818 -6409
rect 3874 -6235 3962 -6222
rect 3874 -6409 3903 -6235
rect 3949 -6409 3962 -6235
rect 3874 -6422 3962 -6409
rect 4133 -6235 4221 -6222
rect 4133 -6409 4146 -6235
rect 4192 -6409 4221 -6235
rect 4133 -6422 4221 -6409
rect 4277 -6235 4381 -6222
rect 4277 -6409 4306 -6235
rect 4352 -6409 4381 -6235
rect 4277 -6422 4381 -6409
rect 4437 -6235 4541 -6222
rect 4437 -6409 4466 -6235
rect 4512 -6409 4541 -6235
rect 4437 -6422 4541 -6409
rect 4597 -6235 4701 -6222
rect 4597 -6409 4626 -6235
rect 4672 -6409 4701 -6235
rect 4597 -6422 4701 -6409
rect 4757 -6235 4861 -6222
rect 4757 -6409 4786 -6235
rect 4832 -6409 4861 -6235
rect 4757 -6422 4861 -6409
rect 4917 -6235 5021 -6222
rect 4917 -6409 4946 -6235
rect 4992 -6409 5021 -6235
rect 4917 -6422 5021 -6409
rect 5077 -6235 5165 -6222
rect 5077 -6409 5106 -6235
rect 5152 -6409 5165 -6235
rect 5077 -6422 5165 -6409
rect 5597 -6236 5685 -6223
rect 5597 -6410 5610 -6236
rect 5656 -6410 5685 -6236
rect 5597 -6423 5685 -6410
rect 5741 -6236 5845 -6223
rect 5741 -6410 5770 -6236
rect 5816 -6410 5845 -6236
rect 5741 -6423 5845 -6410
rect 5901 -6236 6005 -6223
rect 5901 -6410 5930 -6236
rect 5976 -6410 6005 -6236
rect 5901 -6423 6005 -6410
rect 6061 -6236 6165 -6223
rect 6061 -6410 6090 -6236
rect 6136 -6410 6165 -6236
rect 6061 -6423 6165 -6410
rect 6221 -6236 6325 -6223
rect 6221 -6410 6250 -6236
rect 6296 -6410 6325 -6236
rect 6221 -6423 6325 -6410
rect 6381 -6236 6485 -6223
rect 6381 -6410 6410 -6236
rect 6456 -6410 6485 -6236
rect 6381 -6423 6485 -6410
rect 6541 -6236 6629 -6223
rect 6541 -6410 6570 -6236
rect 6616 -6410 6629 -6236
rect 6541 -6423 6629 -6410
rect 6800 -6236 6888 -6223
rect 6800 -6410 6813 -6236
rect 6859 -6410 6888 -6236
rect 6800 -6423 6888 -6410
rect 6944 -6236 7032 -6223
rect 6944 -6410 6973 -6236
rect 7019 -6410 7032 -6236
rect 6944 -6423 7032 -6410
rect -4845 -6579 -4757 -6566
rect -4845 -6753 -4832 -6579
rect -4786 -6753 -4757 -6579
rect -4845 -6766 -4757 -6753
rect -4701 -6579 -4613 -6566
rect -4701 -6753 -4672 -6579
rect -4626 -6753 -4613 -6579
rect -4701 -6766 -4613 -6753
rect -4441 -6579 -4353 -6566
rect -4441 -6753 -4428 -6579
rect -4382 -6753 -4353 -6579
rect -4441 -6766 -4353 -6753
rect -4297 -6579 -4209 -6566
rect -4297 -6753 -4268 -6579
rect -4222 -6753 -4209 -6579
rect -4297 -6766 -4209 -6753
rect -4038 -6579 -3950 -6566
rect -4038 -6753 -4025 -6579
rect -3979 -6753 -3950 -6579
rect -4038 -6766 -3950 -6753
rect -3894 -6579 -3790 -6566
rect -3894 -6753 -3865 -6579
rect -3819 -6753 -3790 -6579
rect -3894 -6766 -3790 -6753
rect -3734 -6579 -3630 -6566
rect -3734 -6753 -3705 -6579
rect -3659 -6753 -3630 -6579
rect -3734 -6766 -3630 -6753
rect -3574 -6579 -3470 -6566
rect -3574 -6753 -3545 -6579
rect -3499 -6753 -3470 -6579
rect -3574 -6766 -3470 -6753
rect -3414 -6579 -3310 -6566
rect -3414 -6753 -3385 -6579
rect -3339 -6753 -3310 -6579
rect -3414 -6766 -3310 -6753
rect -3254 -6579 -3150 -6566
rect -3254 -6753 -3225 -6579
rect -3179 -6753 -3150 -6579
rect -3254 -6766 -3150 -6753
rect -3094 -6579 -3006 -6566
rect -3094 -6753 -3065 -6579
rect -3019 -6753 -3006 -6579
rect -3094 -6766 -3006 -6753
rect -2442 -6572 -2354 -6559
rect -2442 -6746 -2429 -6572
rect -2383 -6746 -2354 -6572
rect -2442 -6759 -2354 -6746
rect -2298 -6572 -2210 -6559
rect -2298 -6746 -2269 -6572
rect -2223 -6746 -2210 -6572
rect -2298 -6759 -2210 -6746
rect -2038 -6572 -1950 -6559
rect -2038 -6746 -2025 -6572
rect -1979 -6746 -1950 -6572
rect -2038 -6759 -1950 -6746
rect -1894 -6572 -1806 -6559
rect -1894 -6746 -1865 -6572
rect -1819 -6746 -1806 -6572
rect -1894 -6759 -1806 -6746
rect -1635 -6572 -1547 -6559
rect -1635 -6746 -1622 -6572
rect -1576 -6746 -1547 -6572
rect -1635 -6759 -1547 -6746
rect -1491 -6572 -1387 -6559
rect -1491 -6746 -1462 -6572
rect -1416 -6746 -1387 -6572
rect -1491 -6759 -1387 -6746
rect -1331 -6572 -1227 -6559
rect -1331 -6746 -1302 -6572
rect -1256 -6746 -1227 -6572
rect -1331 -6759 -1227 -6746
rect -1171 -6572 -1067 -6559
rect -1171 -6746 -1142 -6572
rect -1096 -6746 -1067 -6572
rect -1171 -6759 -1067 -6746
rect -1011 -6572 -907 -6559
rect -1011 -6746 -982 -6572
rect -936 -6746 -907 -6572
rect -1011 -6759 -907 -6746
rect -851 -6572 -747 -6559
rect -851 -6746 -822 -6572
rect -776 -6746 -747 -6572
rect -851 -6759 -747 -6746
rect -691 -6572 -603 -6559
rect -691 -6746 -662 -6572
rect -616 -6746 -603 -6572
rect -691 -6759 -603 -6746
rect 157 -6571 245 -6558
rect 157 -6745 170 -6571
rect 216 -6745 245 -6571
rect 157 -6758 245 -6745
rect 301 -6571 389 -6558
rect 301 -6745 330 -6571
rect 376 -6745 389 -6571
rect 301 -6758 389 -6745
rect 560 -6571 648 -6558
rect 560 -6745 573 -6571
rect 619 -6745 648 -6571
rect 560 -6758 648 -6745
rect 704 -6571 808 -6558
rect 704 -6745 733 -6571
rect 779 -6745 808 -6571
rect 704 -6758 808 -6745
rect 864 -6571 968 -6558
rect 864 -6745 893 -6571
rect 939 -6745 968 -6571
rect 864 -6758 968 -6745
rect 1024 -6571 1128 -6558
rect 1024 -6745 1053 -6571
rect 1099 -6745 1128 -6571
rect 1024 -6758 1128 -6745
rect 1184 -6571 1288 -6558
rect 1184 -6745 1213 -6571
rect 1259 -6745 1288 -6571
rect 1184 -6758 1288 -6745
rect 1344 -6571 1448 -6558
rect 1344 -6745 1373 -6571
rect 1419 -6745 1448 -6571
rect 1344 -6758 1448 -6745
rect 1504 -6571 1592 -6558
rect 1504 -6745 1533 -6571
rect 1579 -6745 1592 -6571
rect 1504 -6758 1592 -6745
rect 1917 -6571 2005 -6558
rect 1917 -6745 1930 -6571
rect 1976 -6745 2005 -6571
rect 1917 -6758 2005 -6745
rect 2061 -6571 2165 -6558
rect 2061 -6745 2090 -6571
rect 2136 -6745 2165 -6571
rect 2061 -6758 2165 -6745
rect 2221 -6571 2325 -6558
rect 2221 -6745 2250 -6571
rect 2296 -6745 2325 -6571
rect 2221 -6758 2325 -6745
rect 2381 -6571 2485 -6558
rect 2381 -6745 2410 -6571
rect 2456 -6745 2485 -6571
rect 2381 -6758 2485 -6745
rect 2541 -6571 2645 -6558
rect 2541 -6745 2570 -6571
rect 2616 -6745 2645 -6571
rect 2541 -6758 2645 -6745
rect 2701 -6571 2805 -6558
rect 2701 -6745 2730 -6571
rect 2776 -6745 2805 -6571
rect 2701 -6758 2805 -6745
rect 2861 -6571 2949 -6558
rect 2861 -6745 2890 -6571
rect 2936 -6745 2949 -6571
rect 2861 -6758 2949 -6745
rect 3120 -6571 3208 -6558
rect 3120 -6745 3133 -6571
rect 3179 -6745 3208 -6571
rect 3120 -6758 3208 -6745
rect 3264 -6571 3352 -6558
rect 3264 -6745 3293 -6571
rect 3339 -6745 3352 -6571
rect 3264 -6758 3352 -6745
rect 3730 -6571 3818 -6558
rect 3730 -6745 3743 -6571
rect 3789 -6745 3818 -6571
rect 3730 -6758 3818 -6745
rect 3874 -6571 3962 -6558
rect 3874 -6745 3903 -6571
rect 3949 -6745 3962 -6571
rect 3874 -6758 3962 -6745
rect 4133 -6571 4221 -6558
rect 4133 -6745 4146 -6571
rect 4192 -6745 4221 -6571
rect 4133 -6758 4221 -6745
rect 4277 -6571 4381 -6558
rect 4277 -6745 4306 -6571
rect 4352 -6745 4381 -6571
rect 4277 -6758 4381 -6745
rect 4437 -6571 4541 -6558
rect 4437 -6745 4466 -6571
rect 4512 -6745 4541 -6571
rect 4437 -6758 4541 -6745
rect 4597 -6571 4701 -6558
rect 4597 -6745 4626 -6571
rect 4672 -6745 4701 -6571
rect 4597 -6758 4701 -6745
rect 4757 -6571 4861 -6558
rect 4757 -6745 4786 -6571
rect 4832 -6745 4861 -6571
rect 4757 -6758 4861 -6745
rect 4917 -6571 5021 -6558
rect 4917 -6745 4946 -6571
rect 4992 -6745 5021 -6571
rect 4917 -6758 5021 -6745
rect 5077 -6571 5165 -6558
rect 5077 -6745 5106 -6571
rect 5152 -6745 5165 -6571
rect 5077 -6758 5165 -6745
rect 5597 -6572 5685 -6559
rect 5597 -6746 5610 -6572
rect 5656 -6746 5685 -6572
rect 5597 -6759 5685 -6746
rect 5741 -6572 5845 -6559
rect 5741 -6746 5770 -6572
rect 5816 -6746 5845 -6572
rect 5741 -6759 5845 -6746
rect 5901 -6572 6005 -6559
rect 5901 -6746 5930 -6572
rect 5976 -6746 6005 -6572
rect 5901 -6759 6005 -6746
rect 6061 -6572 6165 -6559
rect 6061 -6746 6090 -6572
rect 6136 -6746 6165 -6572
rect 6061 -6759 6165 -6746
rect 6221 -6572 6325 -6559
rect 6221 -6746 6250 -6572
rect 6296 -6746 6325 -6572
rect 6221 -6759 6325 -6746
rect 6381 -6572 6485 -6559
rect 6381 -6746 6410 -6572
rect 6456 -6746 6485 -6572
rect 6381 -6759 6485 -6746
rect 6541 -6572 6629 -6559
rect 6541 -6746 6570 -6572
rect 6616 -6746 6629 -6572
rect 6541 -6759 6629 -6746
rect 6800 -6572 6888 -6559
rect 6800 -6746 6813 -6572
rect 6859 -6746 6888 -6572
rect 6800 -6759 6888 -6746
rect 6944 -6572 7032 -6559
rect 6944 -6746 6973 -6572
rect 7019 -6746 7032 -6572
rect 6944 -6759 7032 -6746
rect -4845 -6915 -4757 -6902
rect -4845 -7089 -4832 -6915
rect -4786 -7089 -4757 -6915
rect -4845 -7102 -4757 -7089
rect -4701 -6915 -4613 -6902
rect -4701 -7089 -4672 -6915
rect -4626 -7089 -4613 -6915
rect -4701 -7102 -4613 -7089
rect -4441 -6915 -4353 -6902
rect -4441 -7089 -4428 -6915
rect -4382 -7089 -4353 -6915
rect -4441 -7102 -4353 -7089
rect -4297 -6915 -4209 -6902
rect -4297 -7089 -4268 -6915
rect -4222 -7089 -4209 -6915
rect -4297 -7102 -4209 -7089
rect -4038 -6915 -3950 -6902
rect -4038 -7089 -4025 -6915
rect -3979 -7089 -3950 -6915
rect -4038 -7102 -3950 -7089
rect -3894 -6915 -3790 -6902
rect -3894 -7089 -3865 -6915
rect -3819 -7089 -3790 -6915
rect -3894 -7102 -3790 -7089
rect -3734 -6915 -3630 -6902
rect -3734 -7089 -3705 -6915
rect -3659 -7089 -3630 -6915
rect -3734 -7102 -3630 -7089
rect -3574 -6915 -3470 -6902
rect -3574 -7089 -3545 -6915
rect -3499 -7089 -3470 -6915
rect -3574 -7102 -3470 -7089
rect -3414 -6915 -3310 -6902
rect -3414 -7089 -3385 -6915
rect -3339 -7089 -3310 -6915
rect -3414 -7102 -3310 -7089
rect -3254 -6915 -3150 -6902
rect -3254 -7089 -3225 -6915
rect -3179 -7089 -3150 -6915
rect -3254 -7102 -3150 -7089
rect -3094 -6915 -3006 -6902
rect -3094 -7089 -3065 -6915
rect -3019 -7089 -3006 -6915
rect -3094 -7102 -3006 -7089
rect -2442 -6908 -2354 -6895
rect -2442 -7082 -2429 -6908
rect -2383 -7082 -2354 -6908
rect -2442 -7095 -2354 -7082
rect -2298 -6908 -2210 -6895
rect -2298 -7082 -2269 -6908
rect -2223 -7082 -2210 -6908
rect -2298 -7095 -2210 -7082
rect -2038 -6908 -1950 -6895
rect -2038 -7082 -2025 -6908
rect -1979 -7082 -1950 -6908
rect -2038 -7095 -1950 -7082
rect -1894 -6908 -1806 -6895
rect -1894 -7082 -1865 -6908
rect -1819 -7082 -1806 -6908
rect -1894 -7095 -1806 -7082
rect -1635 -6908 -1547 -6895
rect -1635 -7082 -1622 -6908
rect -1576 -7082 -1547 -6908
rect -1635 -7095 -1547 -7082
rect -1491 -6908 -1387 -6895
rect -1491 -7082 -1462 -6908
rect -1416 -7082 -1387 -6908
rect -1491 -7095 -1387 -7082
rect -1331 -6908 -1227 -6895
rect -1331 -7082 -1302 -6908
rect -1256 -7082 -1227 -6908
rect -1331 -7095 -1227 -7082
rect -1171 -6908 -1067 -6895
rect -1171 -7082 -1142 -6908
rect -1096 -7082 -1067 -6908
rect -1171 -7095 -1067 -7082
rect -1011 -6908 -907 -6895
rect -1011 -7082 -982 -6908
rect -936 -7082 -907 -6908
rect -1011 -7095 -907 -7082
rect -851 -6908 -747 -6895
rect -851 -7082 -822 -6908
rect -776 -7082 -747 -6908
rect -851 -7095 -747 -7082
rect -691 -6908 -603 -6895
rect -691 -7082 -662 -6908
rect -616 -7082 -603 -6908
rect -691 -7095 -603 -7082
rect 157 -6907 245 -6894
rect 157 -7081 170 -6907
rect 216 -7081 245 -6907
rect 157 -7094 245 -7081
rect 301 -6907 389 -6894
rect 301 -7081 330 -6907
rect 376 -7081 389 -6907
rect 301 -7094 389 -7081
rect 560 -6907 648 -6894
rect 560 -7081 573 -6907
rect 619 -7081 648 -6907
rect 560 -7094 648 -7081
rect 704 -6907 808 -6894
rect 704 -7081 733 -6907
rect 779 -7081 808 -6907
rect 704 -7094 808 -7081
rect 864 -6907 968 -6894
rect 864 -7081 893 -6907
rect 939 -7081 968 -6907
rect 864 -7094 968 -7081
rect 1024 -6907 1128 -6894
rect 1024 -7081 1053 -6907
rect 1099 -7081 1128 -6907
rect 1024 -7094 1128 -7081
rect 1184 -6907 1288 -6894
rect 1184 -7081 1213 -6907
rect 1259 -7081 1288 -6907
rect 1184 -7094 1288 -7081
rect 1344 -6907 1448 -6894
rect 1344 -7081 1373 -6907
rect 1419 -7081 1448 -6907
rect 1344 -7094 1448 -7081
rect 1504 -6907 1592 -6894
rect 1504 -7081 1533 -6907
rect 1579 -7081 1592 -6907
rect 1504 -7094 1592 -7081
rect 1917 -6907 2005 -6894
rect 1917 -7081 1930 -6907
rect 1976 -7081 2005 -6907
rect 1917 -7094 2005 -7081
rect 2061 -6907 2165 -6894
rect 2061 -7081 2090 -6907
rect 2136 -7081 2165 -6907
rect 2061 -7094 2165 -7081
rect 2221 -6907 2325 -6894
rect 2221 -7081 2250 -6907
rect 2296 -7081 2325 -6907
rect 2221 -7094 2325 -7081
rect 2381 -6907 2485 -6894
rect 2381 -7081 2410 -6907
rect 2456 -7081 2485 -6907
rect 2381 -7094 2485 -7081
rect 2541 -6907 2645 -6894
rect 2541 -7081 2570 -6907
rect 2616 -7081 2645 -6907
rect 2541 -7094 2645 -7081
rect 2701 -6907 2805 -6894
rect 2701 -7081 2730 -6907
rect 2776 -7081 2805 -6907
rect 2701 -7094 2805 -7081
rect 2861 -6907 2949 -6894
rect 2861 -7081 2890 -6907
rect 2936 -7081 2949 -6907
rect 2861 -7094 2949 -7081
rect 3120 -6907 3208 -6894
rect 3120 -7081 3133 -6907
rect 3179 -7081 3208 -6907
rect 3120 -7094 3208 -7081
rect 3264 -6907 3352 -6894
rect 3264 -7081 3293 -6907
rect 3339 -7081 3352 -6907
rect 3264 -7094 3352 -7081
rect 3730 -6907 3818 -6894
rect 3730 -7081 3743 -6907
rect 3789 -7081 3818 -6907
rect 3730 -7094 3818 -7081
rect 3874 -6907 3962 -6894
rect 3874 -7081 3903 -6907
rect 3949 -7081 3962 -6907
rect 3874 -7094 3962 -7081
rect 4133 -6907 4221 -6894
rect 4133 -7081 4146 -6907
rect 4192 -7081 4221 -6907
rect 4133 -7094 4221 -7081
rect 4277 -6907 4381 -6894
rect 4277 -7081 4306 -6907
rect 4352 -7081 4381 -6907
rect 4277 -7094 4381 -7081
rect 4437 -6907 4541 -6894
rect 4437 -7081 4466 -6907
rect 4512 -7081 4541 -6907
rect 4437 -7094 4541 -7081
rect 4597 -6907 4701 -6894
rect 4597 -7081 4626 -6907
rect 4672 -7081 4701 -6907
rect 4597 -7094 4701 -7081
rect 4757 -6907 4861 -6894
rect 4757 -7081 4786 -6907
rect 4832 -7081 4861 -6907
rect 4757 -7094 4861 -7081
rect 4917 -6907 5021 -6894
rect 4917 -7081 4946 -6907
rect 4992 -7081 5021 -6907
rect 4917 -7094 5021 -7081
rect 5077 -6907 5165 -6894
rect 5077 -7081 5106 -6907
rect 5152 -7081 5165 -6907
rect 5077 -7094 5165 -7081
rect 5597 -6908 5685 -6895
rect 5597 -7082 5610 -6908
rect 5656 -7082 5685 -6908
rect 5597 -7095 5685 -7082
rect 5741 -6908 5845 -6895
rect 5741 -7082 5770 -6908
rect 5816 -7082 5845 -6908
rect 5741 -7095 5845 -7082
rect 5901 -6908 6005 -6895
rect 5901 -7082 5930 -6908
rect 5976 -7082 6005 -6908
rect 5901 -7095 6005 -7082
rect 6061 -6908 6165 -6895
rect 6061 -7082 6090 -6908
rect 6136 -7082 6165 -6908
rect 6061 -7095 6165 -7082
rect 6221 -6908 6325 -6895
rect 6221 -7082 6250 -6908
rect 6296 -7082 6325 -6908
rect 6221 -7095 6325 -7082
rect 6381 -6908 6485 -6895
rect 6381 -7082 6410 -6908
rect 6456 -7082 6485 -6908
rect 6381 -7095 6485 -7082
rect 6541 -6908 6629 -6895
rect 6541 -7082 6570 -6908
rect 6616 -7082 6629 -6908
rect 6541 -7095 6629 -7082
rect 6800 -6908 6888 -6895
rect 6800 -7082 6813 -6908
rect 6859 -7082 6888 -6908
rect 6800 -7095 6888 -7082
rect 6944 -6908 7032 -6895
rect 6944 -7082 6973 -6908
rect 7019 -7082 7032 -6908
rect 6944 -7095 7032 -7082
rect -4845 -7251 -4757 -7238
rect -4845 -7425 -4832 -7251
rect -4786 -7425 -4757 -7251
rect -4845 -7438 -4757 -7425
rect -4701 -7251 -4613 -7238
rect -4701 -7425 -4672 -7251
rect -4626 -7425 -4613 -7251
rect -4701 -7438 -4613 -7425
rect -4441 -7251 -4353 -7238
rect -4441 -7425 -4428 -7251
rect -4382 -7425 -4353 -7251
rect -4441 -7438 -4353 -7425
rect -4297 -7251 -4209 -7238
rect -4297 -7425 -4268 -7251
rect -4222 -7425 -4209 -7251
rect -4297 -7438 -4209 -7425
rect -4038 -7251 -3950 -7238
rect -4038 -7425 -4025 -7251
rect -3979 -7425 -3950 -7251
rect -4038 -7438 -3950 -7425
rect -3894 -7251 -3790 -7238
rect -3894 -7425 -3865 -7251
rect -3819 -7425 -3790 -7251
rect -3894 -7438 -3790 -7425
rect -3734 -7251 -3630 -7238
rect -3734 -7425 -3705 -7251
rect -3659 -7425 -3630 -7251
rect -3734 -7438 -3630 -7425
rect -3574 -7251 -3470 -7238
rect -3574 -7425 -3545 -7251
rect -3499 -7425 -3470 -7251
rect -3574 -7438 -3470 -7425
rect -3414 -7251 -3310 -7238
rect -3414 -7425 -3385 -7251
rect -3339 -7425 -3310 -7251
rect -3414 -7438 -3310 -7425
rect -3254 -7251 -3150 -7238
rect -3254 -7425 -3225 -7251
rect -3179 -7425 -3150 -7251
rect -3254 -7438 -3150 -7425
rect -3094 -7251 -3006 -7238
rect -3094 -7425 -3065 -7251
rect -3019 -7425 -3006 -7251
rect -3094 -7438 -3006 -7425
rect -2442 -7244 -2354 -7231
rect -2442 -7418 -2429 -7244
rect -2383 -7418 -2354 -7244
rect -2442 -7431 -2354 -7418
rect -2298 -7244 -2210 -7231
rect -2298 -7418 -2269 -7244
rect -2223 -7418 -2210 -7244
rect -2298 -7431 -2210 -7418
rect -2038 -7244 -1950 -7231
rect -2038 -7418 -2025 -7244
rect -1979 -7418 -1950 -7244
rect -2038 -7431 -1950 -7418
rect -1894 -7244 -1806 -7231
rect -1894 -7418 -1865 -7244
rect -1819 -7418 -1806 -7244
rect -1894 -7431 -1806 -7418
rect -1635 -7244 -1547 -7231
rect -1635 -7418 -1622 -7244
rect -1576 -7418 -1547 -7244
rect -1635 -7431 -1547 -7418
rect -1491 -7244 -1387 -7231
rect -1491 -7418 -1462 -7244
rect -1416 -7418 -1387 -7244
rect -1491 -7431 -1387 -7418
rect -1331 -7244 -1227 -7231
rect -1331 -7418 -1302 -7244
rect -1256 -7418 -1227 -7244
rect -1331 -7431 -1227 -7418
rect -1171 -7244 -1067 -7231
rect -1171 -7418 -1142 -7244
rect -1096 -7418 -1067 -7244
rect -1171 -7431 -1067 -7418
rect -1011 -7244 -907 -7231
rect -1011 -7418 -982 -7244
rect -936 -7418 -907 -7244
rect -1011 -7431 -907 -7418
rect -851 -7244 -747 -7231
rect -851 -7418 -822 -7244
rect -776 -7418 -747 -7244
rect -851 -7431 -747 -7418
rect -691 -7244 -603 -7231
rect -691 -7418 -662 -7244
rect -616 -7418 -603 -7244
rect -691 -7431 -603 -7418
rect 157 -7243 245 -7230
rect 157 -7417 170 -7243
rect 216 -7417 245 -7243
rect 157 -7430 245 -7417
rect 301 -7243 389 -7230
rect 301 -7417 330 -7243
rect 376 -7417 389 -7243
rect 301 -7430 389 -7417
rect 560 -7243 648 -7230
rect 560 -7417 573 -7243
rect 619 -7417 648 -7243
rect 560 -7430 648 -7417
rect 704 -7243 808 -7230
rect 704 -7417 733 -7243
rect 779 -7417 808 -7243
rect 704 -7430 808 -7417
rect 864 -7243 968 -7230
rect 864 -7417 893 -7243
rect 939 -7417 968 -7243
rect 864 -7430 968 -7417
rect 1024 -7243 1128 -7230
rect 1024 -7417 1053 -7243
rect 1099 -7417 1128 -7243
rect 1024 -7430 1128 -7417
rect 1184 -7243 1288 -7230
rect 1184 -7417 1213 -7243
rect 1259 -7417 1288 -7243
rect 1184 -7430 1288 -7417
rect 1344 -7243 1448 -7230
rect 1344 -7417 1373 -7243
rect 1419 -7417 1448 -7243
rect 1344 -7430 1448 -7417
rect 1504 -7243 1592 -7230
rect 1504 -7417 1533 -7243
rect 1579 -7417 1592 -7243
rect 1504 -7430 1592 -7417
rect 1917 -7243 2005 -7230
rect 1917 -7417 1930 -7243
rect 1976 -7417 2005 -7243
rect 1917 -7430 2005 -7417
rect 2061 -7243 2165 -7230
rect 2061 -7417 2090 -7243
rect 2136 -7417 2165 -7243
rect 2061 -7430 2165 -7417
rect 2221 -7243 2325 -7230
rect 2221 -7417 2250 -7243
rect 2296 -7417 2325 -7243
rect 2221 -7430 2325 -7417
rect 2381 -7243 2485 -7230
rect 2381 -7417 2410 -7243
rect 2456 -7417 2485 -7243
rect 2381 -7430 2485 -7417
rect 2541 -7243 2645 -7230
rect 2541 -7417 2570 -7243
rect 2616 -7417 2645 -7243
rect 2541 -7430 2645 -7417
rect 2701 -7243 2805 -7230
rect 2701 -7417 2730 -7243
rect 2776 -7417 2805 -7243
rect 2701 -7430 2805 -7417
rect 2861 -7243 2949 -7230
rect 2861 -7417 2890 -7243
rect 2936 -7417 2949 -7243
rect 2861 -7430 2949 -7417
rect 3120 -7243 3208 -7230
rect 3120 -7417 3133 -7243
rect 3179 -7417 3208 -7243
rect 3120 -7430 3208 -7417
rect 3264 -7243 3352 -7230
rect 3264 -7417 3293 -7243
rect 3339 -7417 3352 -7243
rect 3264 -7430 3352 -7417
rect 3730 -7243 3818 -7230
rect 3730 -7417 3743 -7243
rect 3789 -7417 3818 -7243
rect 3730 -7430 3818 -7417
rect 3874 -7243 3962 -7230
rect 3874 -7417 3903 -7243
rect 3949 -7417 3962 -7243
rect 3874 -7430 3962 -7417
rect 4133 -7243 4221 -7230
rect 4133 -7417 4146 -7243
rect 4192 -7417 4221 -7243
rect 4133 -7430 4221 -7417
rect 4277 -7243 4381 -7230
rect 4277 -7417 4306 -7243
rect 4352 -7417 4381 -7243
rect 4277 -7430 4381 -7417
rect 4437 -7243 4541 -7230
rect 4437 -7417 4466 -7243
rect 4512 -7417 4541 -7243
rect 4437 -7430 4541 -7417
rect 4597 -7243 4701 -7230
rect 4597 -7417 4626 -7243
rect 4672 -7417 4701 -7243
rect 4597 -7430 4701 -7417
rect 4757 -7243 4861 -7230
rect 4757 -7417 4786 -7243
rect 4832 -7417 4861 -7243
rect 4757 -7430 4861 -7417
rect 4917 -7243 5021 -7230
rect 4917 -7417 4946 -7243
rect 4992 -7417 5021 -7243
rect 4917 -7430 5021 -7417
rect 5077 -7243 5165 -7230
rect 5077 -7417 5106 -7243
rect 5152 -7417 5165 -7243
rect 5077 -7430 5165 -7417
rect 5597 -7244 5685 -7231
rect 5597 -7418 5610 -7244
rect 5656 -7418 5685 -7244
rect 5597 -7431 5685 -7418
rect 5741 -7244 5845 -7231
rect 5741 -7418 5770 -7244
rect 5816 -7418 5845 -7244
rect 5741 -7431 5845 -7418
rect 5901 -7244 6005 -7231
rect 5901 -7418 5930 -7244
rect 5976 -7418 6005 -7244
rect 5901 -7431 6005 -7418
rect 6061 -7244 6165 -7231
rect 6061 -7418 6090 -7244
rect 6136 -7418 6165 -7244
rect 6061 -7431 6165 -7418
rect 6221 -7244 6325 -7231
rect 6221 -7418 6250 -7244
rect 6296 -7418 6325 -7244
rect 6221 -7431 6325 -7418
rect 6381 -7244 6485 -7231
rect 6381 -7418 6410 -7244
rect 6456 -7418 6485 -7244
rect 6381 -7431 6485 -7418
rect 6541 -7244 6629 -7231
rect 6541 -7418 6570 -7244
rect 6616 -7418 6629 -7244
rect 6541 -7431 6629 -7418
rect 6800 -7244 6888 -7231
rect 6800 -7418 6813 -7244
rect 6859 -7418 6888 -7244
rect 6800 -7431 6888 -7418
rect 6944 -7244 7032 -7231
rect 6944 -7418 6973 -7244
rect 7019 -7418 7032 -7244
rect 6944 -7431 7032 -7418
<< ndiffc >>
rect -4832 649 -4786 823
rect -4672 649 -4626 823
rect -4428 649 -4382 823
rect -4268 649 -4222 823
rect -4025 649 -3979 823
rect -3865 649 -3819 823
rect -3705 649 -3659 823
rect -3545 649 -3499 823
rect -3385 649 -3339 823
rect -3225 649 -3179 823
rect -3065 649 -3019 823
rect -2429 656 -2383 830
rect -2269 656 -2223 830
rect -2025 656 -1979 830
rect -1865 656 -1819 830
rect -1622 656 -1576 830
rect -1462 656 -1416 830
rect -1302 656 -1256 830
rect -1142 656 -1096 830
rect -982 656 -936 830
rect -822 656 -776 830
rect -662 656 -616 830
rect 170 657 216 831
rect 330 657 376 831
rect 573 657 619 831
rect 733 657 779 831
rect 893 657 939 831
rect 1053 657 1099 831
rect 1213 657 1259 831
rect 1373 657 1419 831
rect 1533 657 1579 831
rect 1930 657 1976 831
rect 2090 657 2136 831
rect 2250 657 2296 831
rect 2410 657 2456 831
rect 2570 657 2616 831
rect 2730 657 2776 831
rect 2890 657 2936 831
rect 3133 657 3179 831
rect 3293 657 3339 831
rect 3743 657 3789 831
rect 3903 657 3949 831
rect 4146 657 4192 831
rect 4306 657 4352 831
rect 4466 657 4512 831
rect 4626 657 4672 831
rect 4786 657 4832 831
rect 4946 657 4992 831
rect 5106 657 5152 831
rect 5610 656 5656 830
rect 5770 656 5816 830
rect 5930 656 5976 830
rect 6090 656 6136 830
rect 6250 656 6296 830
rect 6410 656 6456 830
rect 6570 656 6616 830
rect 6813 656 6859 830
rect 6973 656 7019 830
rect -4832 313 -4786 487
rect -4672 313 -4626 487
rect -4428 313 -4382 487
rect -4268 313 -4222 487
rect -4025 313 -3979 487
rect -3865 313 -3819 487
rect -3705 313 -3659 487
rect -3545 313 -3499 487
rect -3385 313 -3339 487
rect -3225 313 -3179 487
rect -3065 313 -3019 487
rect -2429 320 -2383 494
rect -2269 320 -2223 494
rect -2025 320 -1979 494
rect -1865 320 -1819 494
rect -1622 320 -1576 494
rect -1462 320 -1416 494
rect -1302 320 -1256 494
rect -1142 320 -1096 494
rect -982 320 -936 494
rect -822 320 -776 494
rect -662 320 -616 494
rect 170 321 216 495
rect 330 321 376 495
rect 573 321 619 495
rect 733 321 779 495
rect 893 321 939 495
rect 1053 321 1099 495
rect 1213 321 1259 495
rect 1373 321 1419 495
rect 1533 321 1579 495
rect 1930 321 1976 495
rect 2090 321 2136 495
rect 2250 321 2296 495
rect 2410 321 2456 495
rect 2570 321 2616 495
rect 2730 321 2776 495
rect 2890 321 2936 495
rect 3133 321 3179 495
rect 3293 321 3339 495
rect 3743 321 3789 495
rect 3903 321 3949 495
rect 4146 321 4192 495
rect 4306 321 4352 495
rect 4466 321 4512 495
rect 4626 321 4672 495
rect 4786 321 4832 495
rect 4946 321 4992 495
rect 5106 321 5152 495
rect 5610 320 5656 494
rect 5770 320 5816 494
rect 5930 320 5976 494
rect 6090 320 6136 494
rect 6250 320 6296 494
rect 6410 320 6456 494
rect 6570 320 6616 494
rect 6813 320 6859 494
rect 6973 320 7019 494
rect -4832 -339 -4786 -165
rect -4672 -339 -4626 -165
rect -4428 -339 -4382 -165
rect -4268 -339 -4222 -165
rect -4025 -339 -3979 -165
rect -3865 -339 -3819 -165
rect -3705 -339 -3659 -165
rect -3545 -339 -3499 -165
rect -3385 -339 -3339 -165
rect -3225 -339 -3179 -165
rect -3065 -339 -3019 -165
rect -2429 -332 -2383 -158
rect -2269 -332 -2223 -158
rect -2025 -332 -1979 -158
rect -1865 -332 -1819 -158
rect -1622 -332 -1576 -158
rect -1462 -332 -1416 -158
rect -1302 -332 -1256 -158
rect -1142 -332 -1096 -158
rect -982 -332 -936 -158
rect -822 -332 -776 -158
rect -662 -332 -616 -158
rect -4832 -675 -4786 -501
rect -4672 -675 -4626 -501
rect -4428 -675 -4382 -501
rect -4268 -675 -4222 -501
rect -4025 -675 -3979 -501
rect -3865 -675 -3819 -501
rect -3705 -675 -3659 -501
rect -3545 -675 -3499 -501
rect -3385 -675 -3339 -501
rect -3225 -675 -3179 -501
rect -3065 -675 -3019 -501
rect -2429 -668 -2383 -494
rect -2269 -668 -2223 -494
rect -2025 -668 -1979 -494
rect -1865 -668 -1819 -494
rect -1622 -668 -1576 -494
rect -1462 -668 -1416 -494
rect -1302 -668 -1256 -494
rect -1142 -668 -1096 -494
rect -982 -668 -936 -494
rect -822 -668 -776 -494
rect -662 -668 -616 -494
rect 1930 -331 1976 -157
rect 2090 -331 2136 -157
rect 2333 -331 2379 -157
rect 2493 -331 2539 -157
rect 2653 -331 2699 -157
rect 2813 -331 2859 -157
rect 2973 -331 3019 -157
rect 3133 -331 3179 -157
rect 3293 -331 3339 -157
rect 3743 -331 3789 -157
rect 3903 -331 3949 -157
rect 4063 -331 4109 -157
rect 4223 -331 4269 -157
rect 4383 -331 4429 -157
rect 4543 -331 4589 -157
rect 4703 -331 4749 -157
rect 4946 -331 4992 -157
rect 5106 -331 5152 -157
rect 5610 -332 5656 -158
rect 5770 -332 5816 -158
rect 6013 -332 6059 -158
rect 6173 -332 6219 -158
rect 6333 -332 6379 -158
rect 6493 -332 6539 -158
rect 6653 -332 6699 -158
rect 6813 -332 6859 -158
rect 6973 -332 7019 -158
rect 1930 -667 1976 -493
rect 2090 -667 2136 -493
rect 2333 -667 2379 -493
rect 2493 -667 2539 -493
rect 2653 -667 2699 -493
rect 2813 -667 2859 -493
rect 2973 -667 3019 -493
rect 3133 -667 3179 -493
rect 3293 -667 3339 -493
rect 3743 -667 3789 -493
rect 3903 -667 3949 -493
rect 4063 -667 4109 -493
rect 4223 -667 4269 -493
rect 4383 -667 4429 -493
rect 4543 -667 4589 -493
rect 4703 -667 4749 -493
rect 4946 -667 4992 -493
rect 5106 -667 5152 -493
rect 5610 -668 5656 -494
rect 5770 -668 5816 -494
rect 6013 -668 6059 -494
rect 6173 -668 6219 -494
rect 6333 -668 6379 -494
rect 6493 -668 6539 -494
rect 6653 -668 6699 -494
rect 6813 -668 6859 -494
rect 6973 -668 7019 -494
rect 160 -1202 206 -1128
rect 320 -1202 366 -1128
rect 480 -1202 526 -1128
rect 640 -1202 686 -1128
rect 800 -1202 846 -1128
rect 160 -1438 206 -1364
rect 320 -1438 366 -1364
rect 480 -1438 526 -1364
rect 640 -1438 686 -1364
rect 800 -1438 846 -1364
rect 160 -1843 206 -1769
rect 320 -1843 366 -1769
rect 480 -1843 526 -1769
rect 640 -1843 686 -1769
rect 800 -1843 846 -1769
rect 160 -2079 206 -2005
rect 320 -2079 366 -2005
rect 480 -2079 526 -2005
rect 640 -2079 686 -2005
rect 800 -2079 846 -2005
rect 160 -4143 206 -4069
rect 320 -4143 366 -4069
rect 480 -4143 526 -4069
rect 640 -4143 686 -4069
rect 800 -4143 846 -4069
rect -4832 -4511 -4786 -4337
rect -4672 -4511 -4626 -4337
rect -4428 -4511 -4382 -4337
rect -4268 -4511 -4222 -4337
rect -4025 -4511 -3979 -4337
rect -3865 -4511 -3819 -4337
rect -3705 -4511 -3659 -4337
rect -3545 -4511 -3499 -4337
rect -3385 -4511 -3339 -4337
rect -3225 -4511 -3179 -4337
rect -3065 -4511 -3019 -4337
rect -2429 -4504 -2383 -4330
rect -2269 -4504 -2223 -4330
rect -2025 -4504 -1979 -4330
rect -1865 -4504 -1819 -4330
rect -1622 -4504 -1576 -4330
rect -1462 -4504 -1416 -4330
rect -1302 -4504 -1256 -4330
rect -1142 -4504 -1096 -4330
rect -982 -4504 -936 -4330
rect -822 -4504 -776 -4330
rect -662 -4504 -616 -4330
rect 160 -4379 206 -4305
rect 320 -4379 366 -4305
rect 480 -4379 526 -4305
rect 640 -4379 686 -4305
rect 800 -4379 846 -4305
rect 1930 -4503 1976 -4329
rect 2090 -4503 2136 -4329
rect 2333 -4503 2379 -4329
rect 2493 -4503 2539 -4329
rect 2653 -4503 2699 -4329
rect 2813 -4503 2859 -4329
rect 2973 -4503 3019 -4329
rect 3133 -4503 3179 -4329
rect 3293 -4503 3339 -4329
rect 3743 -4503 3789 -4329
rect 3903 -4503 3949 -4329
rect 4063 -4503 4109 -4329
rect 4223 -4503 4269 -4329
rect 4383 -4503 4429 -4329
rect 4543 -4503 4589 -4329
rect 4703 -4503 4749 -4329
rect 4946 -4503 4992 -4329
rect 5106 -4503 5152 -4329
rect 5610 -4504 5656 -4330
rect 5770 -4504 5816 -4330
rect 6013 -4504 6059 -4330
rect 6173 -4504 6219 -4330
rect 6333 -4504 6379 -4330
rect 6493 -4504 6539 -4330
rect 6653 -4504 6699 -4330
rect 6813 -4504 6859 -4330
rect 6973 -4504 7019 -4330
rect -4832 -4847 -4786 -4673
rect -4672 -4847 -4626 -4673
rect -4428 -4847 -4382 -4673
rect -4268 -4847 -4222 -4673
rect -4025 -4847 -3979 -4673
rect -3865 -4847 -3819 -4673
rect -3705 -4847 -3659 -4673
rect -3545 -4847 -3499 -4673
rect -3385 -4847 -3339 -4673
rect -3225 -4847 -3179 -4673
rect -3065 -4847 -3019 -4673
rect -2429 -4840 -2383 -4666
rect -2269 -4840 -2223 -4666
rect -2025 -4840 -1979 -4666
rect -1865 -4840 -1819 -4666
rect -1622 -4840 -1576 -4666
rect -1462 -4840 -1416 -4666
rect -1302 -4840 -1256 -4666
rect -1142 -4840 -1096 -4666
rect -982 -4840 -936 -4666
rect -822 -4840 -776 -4666
rect -662 -4840 -616 -4666
rect 1930 -4839 1976 -4665
rect 2090 -4839 2136 -4665
rect 2333 -4839 2379 -4665
rect 2493 -4839 2539 -4665
rect 2653 -4839 2699 -4665
rect 2813 -4839 2859 -4665
rect 2973 -4839 3019 -4665
rect 3133 -4839 3179 -4665
rect 3293 -4839 3339 -4665
rect 3743 -4839 3789 -4665
rect 3903 -4839 3949 -4665
rect 4063 -4839 4109 -4665
rect 4223 -4839 4269 -4665
rect 4383 -4839 4429 -4665
rect 4543 -4839 4589 -4665
rect 4703 -4839 4749 -4665
rect 4946 -4839 4992 -4665
rect 5106 -4839 5152 -4665
rect 5610 -4840 5656 -4666
rect 5770 -4840 5816 -4666
rect 6013 -4840 6059 -4666
rect 6173 -4840 6219 -4666
rect 6333 -4840 6379 -4666
rect 6493 -4840 6539 -4666
rect 6653 -4840 6699 -4666
rect 6813 -4840 6859 -4666
rect 6973 -4840 7019 -4666
rect -4832 -5499 -4786 -5325
rect -4672 -5499 -4626 -5325
rect -4428 -5499 -4382 -5325
rect -4268 -5499 -4222 -5325
rect -4025 -5499 -3979 -5325
rect -3865 -5499 -3819 -5325
rect -3705 -5499 -3659 -5325
rect -3545 -5499 -3499 -5325
rect -3385 -5499 -3339 -5325
rect -3225 -5499 -3179 -5325
rect -3065 -5499 -3019 -5325
rect -2429 -5492 -2383 -5318
rect -2269 -5492 -2223 -5318
rect -2025 -5492 -1979 -5318
rect -1865 -5492 -1819 -5318
rect -1622 -5492 -1576 -5318
rect -1462 -5492 -1416 -5318
rect -1302 -5492 -1256 -5318
rect -1142 -5492 -1096 -5318
rect -982 -5492 -936 -5318
rect -822 -5492 -776 -5318
rect -662 -5492 -616 -5318
rect 170 -5491 216 -5317
rect 330 -5491 376 -5317
rect 573 -5491 619 -5317
rect 733 -5491 779 -5317
rect 893 -5491 939 -5317
rect 1053 -5491 1099 -5317
rect 1213 -5491 1259 -5317
rect 1373 -5491 1419 -5317
rect 1533 -5491 1579 -5317
rect 1930 -5491 1976 -5317
rect 2090 -5491 2136 -5317
rect 2250 -5491 2296 -5317
rect 2410 -5491 2456 -5317
rect 2570 -5491 2616 -5317
rect 2730 -5491 2776 -5317
rect 2890 -5491 2936 -5317
rect 3133 -5491 3179 -5317
rect 3293 -5491 3339 -5317
rect 3743 -5491 3789 -5317
rect 3903 -5491 3949 -5317
rect 4146 -5491 4192 -5317
rect 4306 -5491 4352 -5317
rect 4466 -5491 4512 -5317
rect 4626 -5491 4672 -5317
rect 4786 -5491 4832 -5317
rect 4946 -5491 4992 -5317
rect 5106 -5491 5152 -5317
rect 5610 -5492 5656 -5318
rect 5770 -5492 5816 -5318
rect 5930 -5492 5976 -5318
rect 6090 -5492 6136 -5318
rect 6250 -5492 6296 -5318
rect 6410 -5492 6456 -5318
rect 6570 -5492 6616 -5318
rect 6813 -5492 6859 -5318
rect 6973 -5492 7019 -5318
rect -4832 -5835 -4786 -5661
rect -4672 -5835 -4626 -5661
rect -4428 -5835 -4382 -5661
rect -4268 -5835 -4222 -5661
rect -4025 -5835 -3979 -5661
rect -3865 -5835 -3819 -5661
rect -3705 -5835 -3659 -5661
rect -3545 -5835 -3499 -5661
rect -3385 -5835 -3339 -5661
rect -3225 -5835 -3179 -5661
rect -3065 -5835 -3019 -5661
rect -2429 -5828 -2383 -5654
rect -2269 -5828 -2223 -5654
rect -2025 -5828 -1979 -5654
rect -1865 -5828 -1819 -5654
rect -1622 -5828 -1576 -5654
rect -1462 -5828 -1416 -5654
rect -1302 -5828 -1256 -5654
rect -1142 -5828 -1096 -5654
rect -982 -5828 -936 -5654
rect -822 -5828 -776 -5654
rect -662 -5828 -616 -5654
rect 170 -5827 216 -5653
rect 330 -5827 376 -5653
rect 573 -5827 619 -5653
rect 733 -5827 779 -5653
rect 893 -5827 939 -5653
rect 1053 -5827 1099 -5653
rect 1213 -5827 1259 -5653
rect 1373 -5827 1419 -5653
rect 1533 -5827 1579 -5653
rect 1930 -5827 1976 -5653
rect 2090 -5827 2136 -5653
rect 2250 -5827 2296 -5653
rect 2410 -5827 2456 -5653
rect 2570 -5827 2616 -5653
rect 2730 -5827 2776 -5653
rect 2890 -5827 2936 -5653
rect 3133 -5827 3179 -5653
rect 3293 -5827 3339 -5653
rect 3743 -5827 3789 -5653
rect 3903 -5827 3949 -5653
rect 4146 -5827 4192 -5653
rect 4306 -5827 4352 -5653
rect 4466 -5827 4512 -5653
rect 4626 -5827 4672 -5653
rect 4786 -5827 4832 -5653
rect 4946 -5827 4992 -5653
rect 5106 -5827 5152 -5653
rect 5610 -5828 5656 -5654
rect 5770 -5828 5816 -5654
rect 5930 -5828 5976 -5654
rect 6090 -5828 6136 -5654
rect 6250 -5828 6296 -5654
rect 6410 -5828 6456 -5654
rect 6570 -5828 6616 -5654
rect 6813 -5828 6859 -5654
rect 6973 -5828 7019 -5654
<< pdiffc >>
rect -4832 2239 -4786 2413
rect -4672 2239 -4626 2413
rect -4428 2239 -4382 2413
rect -4268 2239 -4222 2413
rect -4025 2239 -3979 2413
rect -3865 2239 -3819 2413
rect -3705 2239 -3659 2413
rect -3545 2239 -3499 2413
rect -3385 2239 -3339 2413
rect -3225 2239 -3179 2413
rect -3065 2239 -3019 2413
rect -2429 2246 -2383 2420
rect -2269 2246 -2223 2420
rect -2025 2246 -1979 2420
rect -1865 2246 -1819 2420
rect -1622 2246 -1576 2420
rect -1462 2246 -1416 2420
rect -1302 2246 -1256 2420
rect -1142 2246 -1096 2420
rect -982 2246 -936 2420
rect -822 2246 -776 2420
rect -662 2246 -616 2420
rect 170 2247 216 2421
rect 330 2247 376 2421
rect 573 2247 619 2421
rect 733 2247 779 2421
rect 893 2247 939 2421
rect 1053 2247 1099 2421
rect 1213 2247 1259 2421
rect 1373 2247 1419 2421
rect 1533 2247 1579 2421
rect 1930 2247 1976 2421
rect 2090 2247 2136 2421
rect 2250 2247 2296 2421
rect 2410 2247 2456 2421
rect 2570 2247 2616 2421
rect 2730 2247 2776 2421
rect 2890 2247 2936 2421
rect 3133 2247 3179 2421
rect 3293 2247 3339 2421
rect 3743 2247 3789 2421
rect 3903 2247 3949 2421
rect 4146 2247 4192 2421
rect 4306 2247 4352 2421
rect 4466 2247 4512 2421
rect 4626 2247 4672 2421
rect 4786 2247 4832 2421
rect 4946 2247 4992 2421
rect 5106 2247 5152 2421
rect 5610 2246 5656 2420
rect 5770 2246 5816 2420
rect 5930 2246 5976 2420
rect 6090 2246 6136 2420
rect 6250 2246 6296 2420
rect 6410 2246 6456 2420
rect 6570 2246 6616 2420
rect 6813 2246 6859 2420
rect 6973 2246 7019 2420
rect -4832 1903 -4786 2077
rect -4672 1903 -4626 2077
rect -4428 1903 -4382 2077
rect -4268 1903 -4222 2077
rect -4025 1903 -3979 2077
rect -3865 1903 -3819 2077
rect -3705 1903 -3659 2077
rect -3545 1903 -3499 2077
rect -3385 1903 -3339 2077
rect -3225 1903 -3179 2077
rect -3065 1903 -3019 2077
rect -2429 1910 -2383 2084
rect -2269 1910 -2223 2084
rect -2025 1910 -1979 2084
rect -1865 1910 -1819 2084
rect -1622 1910 -1576 2084
rect -1462 1910 -1416 2084
rect -1302 1910 -1256 2084
rect -1142 1910 -1096 2084
rect -982 1910 -936 2084
rect -822 1910 -776 2084
rect -662 1910 -616 2084
rect 170 1911 216 2085
rect 330 1911 376 2085
rect 573 1911 619 2085
rect 733 1911 779 2085
rect 893 1911 939 2085
rect 1053 1911 1099 2085
rect 1213 1911 1259 2085
rect 1373 1911 1419 2085
rect 1533 1911 1579 2085
rect 1930 1911 1976 2085
rect 2090 1911 2136 2085
rect 2250 1911 2296 2085
rect 2410 1911 2456 2085
rect 2570 1911 2616 2085
rect 2730 1911 2776 2085
rect 2890 1911 2936 2085
rect 3133 1911 3179 2085
rect 3293 1911 3339 2085
rect 3743 1911 3789 2085
rect 3903 1911 3949 2085
rect 4146 1911 4192 2085
rect 4306 1911 4352 2085
rect 4466 1911 4512 2085
rect 4626 1911 4672 2085
rect 4786 1911 4832 2085
rect 4946 1911 4992 2085
rect 5106 1911 5152 2085
rect 5610 1910 5656 2084
rect 5770 1910 5816 2084
rect 5930 1910 5976 2084
rect 6090 1910 6136 2084
rect 6250 1910 6296 2084
rect 6410 1910 6456 2084
rect 6570 1910 6616 2084
rect 6813 1910 6859 2084
rect 6973 1910 7019 2084
rect -4832 1567 -4786 1741
rect -4672 1567 -4626 1741
rect -4428 1567 -4382 1741
rect -4268 1567 -4222 1741
rect -4025 1567 -3979 1741
rect -3865 1567 -3819 1741
rect -3705 1567 -3659 1741
rect -3545 1567 -3499 1741
rect -3385 1567 -3339 1741
rect -3225 1567 -3179 1741
rect -3065 1567 -3019 1741
rect -2429 1574 -2383 1748
rect -2269 1574 -2223 1748
rect -2025 1574 -1979 1748
rect -1865 1574 -1819 1748
rect -1622 1574 -1576 1748
rect -1462 1574 -1416 1748
rect -1302 1574 -1256 1748
rect -1142 1574 -1096 1748
rect -982 1574 -936 1748
rect -822 1574 -776 1748
rect -662 1574 -616 1748
rect 170 1575 216 1749
rect 330 1575 376 1749
rect 573 1575 619 1749
rect 733 1575 779 1749
rect 893 1575 939 1749
rect 1053 1575 1099 1749
rect 1213 1575 1259 1749
rect 1373 1575 1419 1749
rect 1533 1575 1579 1749
rect 1930 1575 1976 1749
rect 2090 1575 2136 1749
rect 2250 1575 2296 1749
rect 2410 1575 2456 1749
rect 2570 1575 2616 1749
rect 2730 1575 2776 1749
rect 2890 1575 2936 1749
rect 3133 1575 3179 1749
rect 3293 1575 3339 1749
rect 3743 1575 3789 1749
rect 3903 1575 3949 1749
rect 4146 1575 4192 1749
rect 4306 1575 4352 1749
rect 4466 1575 4512 1749
rect 4626 1575 4672 1749
rect 4786 1575 4832 1749
rect 4946 1575 4992 1749
rect 5106 1575 5152 1749
rect 5610 1574 5656 1748
rect 5770 1574 5816 1748
rect 5930 1574 5976 1748
rect 6090 1574 6136 1748
rect 6250 1574 6296 1748
rect 6410 1574 6456 1748
rect 6570 1574 6616 1748
rect 6813 1574 6859 1748
rect 6973 1574 7019 1748
rect -4832 1231 -4786 1405
rect -4672 1231 -4626 1405
rect -4428 1231 -4382 1405
rect -4268 1231 -4222 1405
rect -4025 1231 -3979 1405
rect -3865 1231 -3819 1405
rect -3705 1231 -3659 1405
rect -3545 1231 -3499 1405
rect -3385 1231 -3339 1405
rect -3225 1231 -3179 1405
rect -3065 1231 -3019 1405
rect -2429 1238 -2383 1412
rect -2269 1238 -2223 1412
rect -2025 1238 -1979 1412
rect -1865 1238 -1819 1412
rect -1622 1238 -1576 1412
rect -1462 1238 -1416 1412
rect -1302 1238 -1256 1412
rect -1142 1238 -1096 1412
rect -982 1238 -936 1412
rect -822 1238 -776 1412
rect -662 1238 -616 1412
rect 170 1239 216 1413
rect 330 1239 376 1413
rect 573 1239 619 1413
rect 733 1239 779 1413
rect 893 1239 939 1413
rect 1053 1239 1099 1413
rect 1213 1239 1259 1413
rect 1373 1239 1419 1413
rect 1533 1239 1579 1413
rect 1930 1239 1976 1413
rect 2090 1239 2136 1413
rect 2250 1239 2296 1413
rect 2410 1239 2456 1413
rect 2570 1239 2616 1413
rect 2730 1239 2776 1413
rect 2890 1239 2936 1413
rect 3133 1239 3179 1413
rect 3293 1239 3339 1413
rect 3743 1239 3789 1413
rect 3903 1239 3949 1413
rect 4146 1239 4192 1413
rect 4306 1239 4352 1413
rect 4466 1239 4512 1413
rect 4626 1239 4672 1413
rect 4786 1239 4832 1413
rect 4946 1239 4992 1413
rect 5106 1239 5152 1413
rect 5610 1238 5656 1412
rect 5770 1238 5816 1412
rect 5930 1238 5976 1412
rect 6090 1238 6136 1412
rect 6250 1238 6296 1412
rect 6410 1238 6456 1412
rect 6570 1238 6616 1412
rect 6813 1238 6859 1412
rect 6973 1238 7019 1412
rect 160 -517 206 -343
rect 320 -517 366 -343
rect 480 -517 526 -343
rect 640 -517 686 -343
rect 800 -517 846 -343
rect 160 -853 206 -679
rect 320 -853 366 -679
rect 480 -853 526 -679
rect 640 -853 686 -679
rect 800 -853 846 -679
rect -4832 -1257 -4786 -1083
rect -4672 -1257 -4626 -1083
rect -4428 -1257 -4382 -1083
rect -4268 -1257 -4222 -1083
rect -4025 -1257 -3979 -1083
rect -3865 -1257 -3819 -1083
rect -3705 -1257 -3659 -1083
rect -3545 -1257 -3499 -1083
rect -3385 -1257 -3339 -1083
rect -3225 -1257 -3179 -1083
rect -3065 -1257 -3019 -1083
rect -2429 -1250 -2383 -1076
rect -2269 -1250 -2223 -1076
rect -2025 -1250 -1979 -1076
rect -1865 -1250 -1819 -1076
rect -1622 -1250 -1576 -1076
rect -1462 -1250 -1416 -1076
rect -1302 -1250 -1256 -1076
rect -1142 -1250 -1096 -1076
rect -982 -1250 -936 -1076
rect -822 -1250 -776 -1076
rect -662 -1250 -616 -1076
rect 1930 -1249 1976 -1075
rect 2090 -1249 2136 -1075
rect 2333 -1249 2379 -1075
rect 2493 -1249 2539 -1075
rect 2653 -1249 2699 -1075
rect 2813 -1249 2859 -1075
rect 2973 -1249 3019 -1075
rect 3133 -1249 3179 -1075
rect 3293 -1249 3339 -1075
rect 3743 -1249 3789 -1075
rect 3903 -1249 3949 -1075
rect 4063 -1249 4109 -1075
rect 4223 -1249 4269 -1075
rect 4383 -1249 4429 -1075
rect 4543 -1249 4589 -1075
rect 4703 -1249 4749 -1075
rect 4946 -1249 4992 -1075
rect 5106 -1249 5152 -1075
rect 5610 -1250 5656 -1076
rect -4832 -1593 -4786 -1419
rect -4672 -1593 -4626 -1419
rect -4428 -1593 -4382 -1419
rect -4268 -1593 -4222 -1419
rect -4025 -1593 -3979 -1419
rect -3865 -1593 -3819 -1419
rect -3705 -1593 -3659 -1419
rect -3545 -1593 -3499 -1419
rect -3385 -1593 -3339 -1419
rect -3225 -1593 -3179 -1419
rect -3065 -1593 -3019 -1419
rect -2429 -1586 -2383 -1412
rect -2269 -1586 -2223 -1412
rect -2025 -1586 -1979 -1412
rect -1865 -1586 -1819 -1412
rect -1622 -1586 -1576 -1412
rect -1462 -1586 -1416 -1412
rect -1302 -1586 -1256 -1412
rect -1142 -1586 -1096 -1412
rect -982 -1586 -936 -1412
rect -822 -1586 -776 -1412
rect -662 -1586 -616 -1412
rect 5770 -1250 5816 -1076
rect 6013 -1250 6059 -1076
rect 6173 -1250 6219 -1076
rect 6333 -1250 6379 -1076
rect 6493 -1250 6539 -1076
rect 6653 -1250 6699 -1076
rect 6813 -1250 6859 -1076
rect 6973 -1250 7019 -1076
rect 1930 -1585 1976 -1411
rect 2090 -1585 2136 -1411
rect 2333 -1585 2379 -1411
rect 2493 -1585 2539 -1411
rect 2653 -1585 2699 -1411
rect 2813 -1585 2859 -1411
rect 2973 -1585 3019 -1411
rect 3133 -1585 3179 -1411
rect 3293 -1585 3339 -1411
rect 3743 -1585 3789 -1411
rect 3903 -1585 3949 -1411
rect 4063 -1585 4109 -1411
rect 4223 -1585 4269 -1411
rect 4383 -1585 4429 -1411
rect 4543 -1585 4589 -1411
rect 4703 -1585 4749 -1411
rect 4946 -1585 4992 -1411
rect 5106 -1585 5152 -1411
rect 5610 -1586 5656 -1412
rect -4832 -1929 -4786 -1755
rect -4672 -1929 -4626 -1755
rect -4428 -1929 -4382 -1755
rect -4268 -1929 -4222 -1755
rect -4025 -1929 -3979 -1755
rect -3865 -1929 -3819 -1755
rect -3705 -1929 -3659 -1755
rect -3545 -1929 -3499 -1755
rect -3385 -1929 -3339 -1755
rect -3225 -1929 -3179 -1755
rect -3065 -1929 -3019 -1755
rect -2429 -1922 -2383 -1748
rect -2269 -1922 -2223 -1748
rect -2025 -1922 -1979 -1748
rect -1865 -1922 -1819 -1748
rect -1622 -1922 -1576 -1748
rect -1462 -1922 -1416 -1748
rect -1302 -1922 -1256 -1748
rect -1142 -1922 -1096 -1748
rect -982 -1922 -936 -1748
rect -822 -1922 -776 -1748
rect -662 -1922 -616 -1748
rect 5770 -1586 5816 -1412
rect 6013 -1586 6059 -1412
rect 6173 -1586 6219 -1412
rect 6333 -1586 6379 -1412
rect 6493 -1586 6539 -1412
rect 6653 -1586 6699 -1412
rect 6813 -1586 6859 -1412
rect 6973 -1586 7019 -1412
rect 1930 -1921 1976 -1747
rect 2090 -1921 2136 -1747
rect 2333 -1921 2379 -1747
rect 2493 -1921 2539 -1747
rect 2653 -1921 2699 -1747
rect 2813 -1921 2859 -1747
rect 2973 -1921 3019 -1747
rect 3133 -1921 3179 -1747
rect 3293 -1921 3339 -1747
rect 3743 -1921 3789 -1747
rect 3903 -1921 3949 -1747
rect 4063 -1921 4109 -1747
rect 4223 -1921 4269 -1747
rect 4383 -1921 4429 -1747
rect 4543 -1921 4589 -1747
rect 4703 -1921 4749 -1747
rect 4946 -1921 4992 -1747
rect 5106 -1921 5152 -1747
rect 5610 -1922 5656 -1748
rect -4832 -2265 -4786 -2091
rect -4672 -2265 -4626 -2091
rect -4428 -2265 -4382 -2091
rect -4268 -2265 -4222 -2091
rect -4025 -2265 -3979 -2091
rect -3865 -2265 -3819 -2091
rect -3705 -2265 -3659 -2091
rect -3545 -2265 -3499 -2091
rect -3385 -2265 -3339 -2091
rect -3225 -2265 -3179 -2091
rect -3065 -2265 -3019 -2091
rect -2429 -2258 -2383 -2084
rect -2269 -2258 -2223 -2084
rect -2025 -2258 -1979 -2084
rect -1865 -2258 -1819 -2084
rect -1622 -2258 -1576 -2084
rect -1462 -2258 -1416 -2084
rect -1302 -2258 -1256 -2084
rect -1142 -2258 -1096 -2084
rect -982 -2258 -936 -2084
rect -822 -2258 -776 -2084
rect -662 -2258 -616 -2084
rect 5770 -1922 5816 -1748
rect 6013 -1922 6059 -1748
rect 6173 -1922 6219 -1748
rect 6333 -1922 6379 -1748
rect 6493 -1922 6539 -1748
rect 6653 -1922 6699 -1748
rect 6813 -1922 6859 -1748
rect 6973 -1922 7019 -1748
rect 1930 -2257 1976 -2083
rect 2090 -2257 2136 -2083
rect 2333 -2257 2379 -2083
rect 2493 -2257 2539 -2083
rect 2653 -2257 2699 -2083
rect 2813 -2257 2859 -2083
rect 2973 -2257 3019 -2083
rect 3133 -2257 3179 -2083
rect 3293 -2257 3339 -2083
rect 3743 -2257 3789 -2083
rect 3903 -2257 3949 -2083
rect 4063 -2257 4109 -2083
rect 4223 -2257 4269 -2083
rect 4383 -2257 4429 -2083
rect 4543 -2257 4589 -2083
rect 4703 -2257 4749 -2083
rect 4946 -2257 4992 -2083
rect 5106 -2257 5152 -2083
rect 5610 -2258 5656 -2084
rect 5770 -2258 5816 -2084
rect 6013 -2258 6059 -2084
rect 6173 -2258 6219 -2084
rect 6333 -2258 6379 -2084
rect 6493 -2258 6539 -2084
rect 6653 -2258 6699 -2084
rect 6813 -2258 6859 -2084
rect 6973 -2258 7019 -2084
rect 160 -2528 206 -2354
rect 320 -2528 366 -2354
rect 480 -2528 526 -2354
rect 640 -2528 686 -2354
rect 800 -2528 846 -2354
rect -4832 -2921 -4786 -2747
rect -4672 -2921 -4626 -2747
rect -4428 -2921 -4382 -2747
rect -4268 -2921 -4222 -2747
rect -4025 -2921 -3979 -2747
rect -3865 -2921 -3819 -2747
rect -3705 -2921 -3659 -2747
rect -3545 -2921 -3499 -2747
rect -3385 -2921 -3339 -2747
rect -3225 -2921 -3179 -2747
rect -3065 -2921 -3019 -2747
rect -2429 -2914 -2383 -2740
rect -2269 -2914 -2223 -2740
rect -2025 -2914 -1979 -2740
rect -1865 -2914 -1819 -2740
rect -1622 -2914 -1576 -2740
rect -1462 -2914 -1416 -2740
rect -1302 -2914 -1256 -2740
rect -1142 -2914 -1096 -2740
rect -982 -2914 -936 -2740
rect -822 -2914 -776 -2740
rect -662 -2914 -616 -2740
rect 160 -2864 206 -2690
rect 320 -2864 366 -2690
rect 480 -2864 526 -2690
rect 640 -2864 686 -2690
rect 800 -2864 846 -2690
rect 1930 -2913 1976 -2739
rect 2090 -2913 2136 -2739
rect 2333 -2913 2379 -2739
rect 2493 -2913 2539 -2739
rect 2653 -2913 2699 -2739
rect 2813 -2913 2859 -2739
rect 2973 -2913 3019 -2739
rect 3133 -2913 3179 -2739
rect 3293 -2913 3339 -2739
rect 3743 -2913 3789 -2739
rect 3903 -2913 3949 -2739
rect 4063 -2913 4109 -2739
rect 4223 -2913 4269 -2739
rect 4383 -2913 4429 -2739
rect 4543 -2913 4589 -2739
rect 4703 -2913 4749 -2739
rect 4946 -2913 4992 -2739
rect 5106 -2913 5152 -2739
rect 5610 -2914 5656 -2740
rect -4832 -3257 -4786 -3083
rect -4672 -3257 -4626 -3083
rect -4428 -3257 -4382 -3083
rect -4268 -3257 -4222 -3083
rect -4025 -3257 -3979 -3083
rect -3865 -3257 -3819 -3083
rect -3705 -3257 -3659 -3083
rect -3545 -3257 -3499 -3083
rect -3385 -3257 -3339 -3083
rect -3225 -3257 -3179 -3083
rect -3065 -3257 -3019 -3083
rect -2429 -3250 -2383 -3076
rect -2269 -3250 -2223 -3076
rect -2025 -3250 -1979 -3076
rect -1865 -3250 -1819 -3076
rect -1622 -3250 -1576 -3076
rect -1462 -3250 -1416 -3076
rect -1302 -3250 -1256 -3076
rect -1142 -3250 -1096 -3076
rect -982 -3250 -936 -3076
rect -822 -3250 -776 -3076
rect -662 -3250 -616 -3076
rect 5770 -2914 5816 -2740
rect 6013 -2914 6059 -2740
rect 6173 -2914 6219 -2740
rect 6333 -2914 6379 -2740
rect 6493 -2914 6539 -2740
rect 6653 -2914 6699 -2740
rect 6813 -2914 6859 -2740
rect 6973 -2914 7019 -2740
rect 1930 -3249 1976 -3075
rect 2090 -3249 2136 -3075
rect 2333 -3249 2379 -3075
rect 2493 -3249 2539 -3075
rect 2653 -3249 2699 -3075
rect 2813 -3249 2859 -3075
rect 2973 -3249 3019 -3075
rect 3133 -3249 3179 -3075
rect 3293 -3249 3339 -3075
rect 3743 -3249 3789 -3075
rect 3903 -3249 3949 -3075
rect 4063 -3249 4109 -3075
rect 4223 -3249 4269 -3075
rect 4383 -3249 4429 -3075
rect 4543 -3249 4589 -3075
rect 4703 -3249 4749 -3075
rect 4946 -3249 4992 -3075
rect 5106 -3249 5152 -3075
rect 5610 -3250 5656 -3076
rect -4832 -3593 -4786 -3419
rect -4672 -3593 -4626 -3419
rect -4428 -3593 -4382 -3419
rect -4268 -3593 -4222 -3419
rect -4025 -3593 -3979 -3419
rect -3865 -3593 -3819 -3419
rect -3705 -3593 -3659 -3419
rect -3545 -3593 -3499 -3419
rect -3385 -3593 -3339 -3419
rect -3225 -3593 -3179 -3419
rect -3065 -3593 -3019 -3419
rect -2429 -3586 -2383 -3412
rect -2269 -3586 -2223 -3412
rect -2025 -3586 -1979 -3412
rect -1865 -3586 -1819 -3412
rect -1622 -3586 -1576 -3412
rect -1462 -3586 -1416 -3412
rect -1302 -3586 -1256 -3412
rect -1142 -3586 -1096 -3412
rect -982 -3586 -936 -3412
rect -822 -3586 -776 -3412
rect -662 -3586 -616 -3412
rect 160 -3458 206 -3284
rect 320 -3458 366 -3284
rect 480 -3458 526 -3284
rect 640 -3458 686 -3284
rect 800 -3458 846 -3284
rect 5770 -3250 5816 -3076
rect 6013 -3250 6059 -3076
rect 6173 -3250 6219 -3076
rect 6333 -3250 6379 -3076
rect 6493 -3250 6539 -3076
rect 6653 -3250 6699 -3076
rect 6813 -3250 6859 -3076
rect 6973 -3250 7019 -3076
rect 1930 -3585 1976 -3411
rect 2090 -3585 2136 -3411
rect 2333 -3585 2379 -3411
rect 2493 -3585 2539 -3411
rect 2653 -3585 2699 -3411
rect 2813 -3585 2859 -3411
rect 2973 -3585 3019 -3411
rect 3133 -3585 3179 -3411
rect 3293 -3585 3339 -3411
rect 3743 -3585 3789 -3411
rect 3903 -3585 3949 -3411
rect 4063 -3585 4109 -3411
rect 4223 -3585 4269 -3411
rect 4383 -3585 4429 -3411
rect 4543 -3585 4589 -3411
rect 4703 -3585 4749 -3411
rect 4946 -3585 4992 -3411
rect 5106 -3585 5152 -3411
rect 5610 -3586 5656 -3412
rect -4832 -3929 -4786 -3755
rect -4672 -3929 -4626 -3755
rect -4428 -3929 -4382 -3755
rect -4268 -3929 -4222 -3755
rect -4025 -3929 -3979 -3755
rect -3865 -3929 -3819 -3755
rect -3705 -3929 -3659 -3755
rect -3545 -3929 -3499 -3755
rect -3385 -3929 -3339 -3755
rect -3225 -3929 -3179 -3755
rect -3065 -3929 -3019 -3755
rect -2429 -3922 -2383 -3748
rect -2269 -3922 -2223 -3748
rect -2025 -3922 -1979 -3748
rect -1865 -3922 -1819 -3748
rect -1622 -3922 -1576 -3748
rect -1462 -3922 -1416 -3748
rect -1302 -3922 -1256 -3748
rect -1142 -3922 -1096 -3748
rect -982 -3922 -936 -3748
rect -822 -3922 -776 -3748
rect -662 -3922 -616 -3748
rect 160 -3794 206 -3620
rect 320 -3794 366 -3620
rect 480 -3794 526 -3620
rect 640 -3794 686 -3620
rect 800 -3794 846 -3620
rect 5770 -3586 5816 -3412
rect 6013 -3586 6059 -3412
rect 6173 -3586 6219 -3412
rect 6333 -3586 6379 -3412
rect 6493 -3586 6539 -3412
rect 6653 -3586 6699 -3412
rect 6813 -3586 6859 -3412
rect 6973 -3586 7019 -3412
rect 1930 -3921 1976 -3747
rect 2090 -3921 2136 -3747
rect 2333 -3921 2379 -3747
rect 2493 -3921 2539 -3747
rect 2653 -3921 2699 -3747
rect 2813 -3921 2859 -3747
rect 2973 -3921 3019 -3747
rect 3133 -3921 3179 -3747
rect 3293 -3921 3339 -3747
rect 3743 -3921 3789 -3747
rect 3903 -3921 3949 -3747
rect 4063 -3921 4109 -3747
rect 4223 -3921 4269 -3747
rect 4383 -3921 4429 -3747
rect 4543 -3921 4589 -3747
rect 4703 -3921 4749 -3747
rect 4946 -3921 4992 -3747
rect 5106 -3921 5152 -3747
rect 5610 -3922 5656 -3748
rect 5770 -3922 5816 -3748
rect 6013 -3922 6059 -3748
rect 6173 -3922 6219 -3748
rect 6333 -3922 6379 -3748
rect 6493 -3922 6539 -3748
rect 6653 -3922 6699 -3748
rect 6813 -3922 6859 -3748
rect 6973 -3922 7019 -3748
rect -4832 -6417 -4786 -6243
rect -4672 -6417 -4626 -6243
rect -4428 -6417 -4382 -6243
rect -4268 -6417 -4222 -6243
rect -4025 -6417 -3979 -6243
rect -3865 -6417 -3819 -6243
rect -3705 -6417 -3659 -6243
rect -3545 -6417 -3499 -6243
rect -3385 -6417 -3339 -6243
rect -3225 -6417 -3179 -6243
rect -3065 -6417 -3019 -6243
rect -2429 -6410 -2383 -6236
rect -2269 -6410 -2223 -6236
rect -2025 -6410 -1979 -6236
rect -1865 -6410 -1819 -6236
rect -1622 -6410 -1576 -6236
rect -1462 -6410 -1416 -6236
rect -1302 -6410 -1256 -6236
rect -1142 -6410 -1096 -6236
rect -982 -6410 -936 -6236
rect -822 -6410 -776 -6236
rect -662 -6410 -616 -6236
rect 170 -6409 216 -6235
rect 330 -6409 376 -6235
rect 573 -6409 619 -6235
rect 733 -6409 779 -6235
rect 893 -6409 939 -6235
rect 1053 -6409 1099 -6235
rect 1213 -6409 1259 -6235
rect 1373 -6409 1419 -6235
rect 1533 -6409 1579 -6235
rect 1930 -6409 1976 -6235
rect 2090 -6409 2136 -6235
rect 2250 -6409 2296 -6235
rect 2410 -6409 2456 -6235
rect 2570 -6409 2616 -6235
rect 2730 -6409 2776 -6235
rect 2890 -6409 2936 -6235
rect 3133 -6409 3179 -6235
rect 3293 -6409 3339 -6235
rect 3743 -6409 3789 -6235
rect 3903 -6409 3949 -6235
rect 4146 -6409 4192 -6235
rect 4306 -6409 4352 -6235
rect 4466 -6409 4512 -6235
rect 4626 -6409 4672 -6235
rect 4786 -6409 4832 -6235
rect 4946 -6409 4992 -6235
rect 5106 -6409 5152 -6235
rect 5610 -6410 5656 -6236
rect 5770 -6410 5816 -6236
rect 5930 -6410 5976 -6236
rect 6090 -6410 6136 -6236
rect 6250 -6410 6296 -6236
rect 6410 -6410 6456 -6236
rect 6570 -6410 6616 -6236
rect 6813 -6410 6859 -6236
rect 6973 -6410 7019 -6236
rect -4832 -6753 -4786 -6579
rect -4672 -6753 -4626 -6579
rect -4428 -6753 -4382 -6579
rect -4268 -6753 -4222 -6579
rect -4025 -6753 -3979 -6579
rect -3865 -6753 -3819 -6579
rect -3705 -6753 -3659 -6579
rect -3545 -6753 -3499 -6579
rect -3385 -6753 -3339 -6579
rect -3225 -6753 -3179 -6579
rect -3065 -6753 -3019 -6579
rect -2429 -6746 -2383 -6572
rect -2269 -6746 -2223 -6572
rect -2025 -6746 -1979 -6572
rect -1865 -6746 -1819 -6572
rect -1622 -6746 -1576 -6572
rect -1462 -6746 -1416 -6572
rect -1302 -6746 -1256 -6572
rect -1142 -6746 -1096 -6572
rect -982 -6746 -936 -6572
rect -822 -6746 -776 -6572
rect -662 -6746 -616 -6572
rect 170 -6745 216 -6571
rect 330 -6745 376 -6571
rect 573 -6745 619 -6571
rect 733 -6745 779 -6571
rect 893 -6745 939 -6571
rect 1053 -6745 1099 -6571
rect 1213 -6745 1259 -6571
rect 1373 -6745 1419 -6571
rect 1533 -6745 1579 -6571
rect 1930 -6745 1976 -6571
rect 2090 -6745 2136 -6571
rect 2250 -6745 2296 -6571
rect 2410 -6745 2456 -6571
rect 2570 -6745 2616 -6571
rect 2730 -6745 2776 -6571
rect 2890 -6745 2936 -6571
rect 3133 -6745 3179 -6571
rect 3293 -6745 3339 -6571
rect 3743 -6745 3789 -6571
rect 3903 -6745 3949 -6571
rect 4146 -6745 4192 -6571
rect 4306 -6745 4352 -6571
rect 4466 -6745 4512 -6571
rect 4626 -6745 4672 -6571
rect 4786 -6745 4832 -6571
rect 4946 -6745 4992 -6571
rect 5106 -6745 5152 -6571
rect 5610 -6746 5656 -6572
rect 5770 -6746 5816 -6572
rect 5930 -6746 5976 -6572
rect 6090 -6746 6136 -6572
rect 6250 -6746 6296 -6572
rect 6410 -6746 6456 -6572
rect 6570 -6746 6616 -6572
rect 6813 -6746 6859 -6572
rect 6973 -6746 7019 -6572
rect -4832 -7089 -4786 -6915
rect -4672 -7089 -4626 -6915
rect -4428 -7089 -4382 -6915
rect -4268 -7089 -4222 -6915
rect -4025 -7089 -3979 -6915
rect -3865 -7089 -3819 -6915
rect -3705 -7089 -3659 -6915
rect -3545 -7089 -3499 -6915
rect -3385 -7089 -3339 -6915
rect -3225 -7089 -3179 -6915
rect -3065 -7089 -3019 -6915
rect -2429 -7082 -2383 -6908
rect -2269 -7082 -2223 -6908
rect -2025 -7082 -1979 -6908
rect -1865 -7082 -1819 -6908
rect -1622 -7082 -1576 -6908
rect -1462 -7082 -1416 -6908
rect -1302 -7082 -1256 -6908
rect -1142 -7082 -1096 -6908
rect -982 -7082 -936 -6908
rect -822 -7082 -776 -6908
rect -662 -7082 -616 -6908
rect 170 -7081 216 -6907
rect 330 -7081 376 -6907
rect 573 -7081 619 -6907
rect 733 -7081 779 -6907
rect 893 -7081 939 -6907
rect 1053 -7081 1099 -6907
rect 1213 -7081 1259 -6907
rect 1373 -7081 1419 -6907
rect 1533 -7081 1579 -6907
rect 1930 -7081 1976 -6907
rect 2090 -7081 2136 -6907
rect 2250 -7081 2296 -6907
rect 2410 -7081 2456 -6907
rect 2570 -7081 2616 -6907
rect 2730 -7081 2776 -6907
rect 2890 -7081 2936 -6907
rect 3133 -7081 3179 -6907
rect 3293 -7081 3339 -6907
rect 3743 -7081 3789 -6907
rect 3903 -7081 3949 -6907
rect 4146 -7081 4192 -6907
rect 4306 -7081 4352 -6907
rect 4466 -7081 4512 -6907
rect 4626 -7081 4672 -6907
rect 4786 -7081 4832 -6907
rect 4946 -7081 4992 -6907
rect 5106 -7081 5152 -6907
rect 5610 -7082 5656 -6908
rect 5770 -7082 5816 -6908
rect 5930 -7082 5976 -6908
rect 6090 -7082 6136 -6908
rect 6250 -7082 6296 -6908
rect 6410 -7082 6456 -6908
rect 6570 -7082 6616 -6908
rect 6813 -7082 6859 -6908
rect 6973 -7082 7019 -6908
rect -4832 -7425 -4786 -7251
rect -4672 -7425 -4626 -7251
rect -4428 -7425 -4382 -7251
rect -4268 -7425 -4222 -7251
rect -4025 -7425 -3979 -7251
rect -3865 -7425 -3819 -7251
rect -3705 -7425 -3659 -7251
rect -3545 -7425 -3499 -7251
rect -3385 -7425 -3339 -7251
rect -3225 -7425 -3179 -7251
rect -3065 -7425 -3019 -7251
rect -2429 -7418 -2383 -7244
rect -2269 -7418 -2223 -7244
rect -2025 -7418 -1979 -7244
rect -1865 -7418 -1819 -7244
rect -1622 -7418 -1576 -7244
rect -1462 -7418 -1416 -7244
rect -1302 -7418 -1256 -7244
rect -1142 -7418 -1096 -7244
rect -982 -7418 -936 -7244
rect -822 -7418 -776 -7244
rect -662 -7418 -616 -7244
rect 170 -7417 216 -7243
rect 330 -7417 376 -7243
rect 573 -7417 619 -7243
rect 733 -7417 779 -7243
rect 893 -7417 939 -7243
rect 1053 -7417 1099 -7243
rect 1213 -7417 1259 -7243
rect 1373 -7417 1419 -7243
rect 1533 -7417 1579 -7243
rect 1930 -7417 1976 -7243
rect 2090 -7417 2136 -7243
rect 2250 -7417 2296 -7243
rect 2410 -7417 2456 -7243
rect 2570 -7417 2616 -7243
rect 2730 -7417 2776 -7243
rect 2890 -7417 2936 -7243
rect 3133 -7417 3179 -7243
rect 3293 -7417 3339 -7243
rect 3743 -7417 3789 -7243
rect 3903 -7417 3949 -7243
rect 4146 -7417 4192 -7243
rect 4306 -7417 4352 -7243
rect 4466 -7417 4512 -7243
rect 4626 -7417 4672 -7243
rect 4786 -7417 4832 -7243
rect 4946 -7417 4992 -7243
rect 5106 -7417 5152 -7243
rect 5610 -7418 5656 -7244
rect 5770 -7418 5816 -7244
rect 5930 -7418 5976 -7244
rect 6090 -7418 6136 -7244
rect 6250 -7418 6296 -7244
rect 6410 -7418 6456 -7244
rect 6570 -7418 6616 -7244
rect 6813 -7418 6859 -7244
rect 6973 -7418 7019 -7244
<< psubdiff >>
rect -4901 101 -2950 131
rect -4901 47 -4688 101
rect -4527 47 -4467 101
rect -4306 47 -4246 101
rect -4085 47 -4025 101
rect -3864 47 -3804 101
rect -3643 47 -3583 101
rect -3422 47 -3362 101
rect -3201 47 -3141 101
rect -2980 47 -2950 101
rect -4901 17 -2950 47
rect -2498 108 -547 138
rect -2498 54 -2285 108
rect -2124 54 -2064 108
rect -1903 54 -1843 108
rect -1682 54 -1622 108
rect -1461 54 -1401 108
rect -1240 54 -1180 108
rect -1019 54 -959 108
rect -798 54 -738 108
rect -577 54 -547 108
rect -2498 24 -547 54
rect 101 109 1648 139
rect 101 55 131 109
rect 292 55 352 109
rect 513 55 573 109
rect 734 55 794 109
rect 955 55 1015 109
rect 1176 55 1236 109
rect 1397 55 1457 109
rect 1618 55 1648 109
rect 101 25 1648 55
rect 1861 109 3408 139
rect 1861 55 1891 109
rect 2052 55 2112 109
rect 2273 55 2333 109
rect 2494 55 2554 109
rect 2715 55 2775 109
rect 2936 55 2996 109
rect 3157 55 3217 109
rect 3378 55 3408 109
rect 1861 25 3408 55
rect 3674 109 5221 139
rect 3674 55 3704 109
rect 3865 55 3925 109
rect 4086 55 4146 109
rect 4307 55 4367 109
rect 4528 55 4588 109
rect 4749 55 4809 109
rect 4970 55 5030 109
rect 5191 55 5221 109
rect 3674 25 5221 55
rect 5541 108 7088 138
rect 5541 54 5571 108
rect 5732 54 5792 108
rect 5953 54 6013 108
rect 6174 54 6234 108
rect 6395 54 6455 108
rect 6616 54 6676 108
rect 6837 54 6897 108
rect 7058 54 7088 108
rect 5541 24 7088 54
rect 93 -1576 908 -1558
rect 93 -1631 115 -1576
rect 879 -1631 908 -1576
rect 93 -1649 908 -1631
rect 93 -4517 908 -4499
rect 93 -4572 115 -4517
rect 879 -4572 908 -4517
rect 93 -4590 908 -4572
rect -4901 -5059 -2950 -5029
rect -4901 -5113 -4688 -5059
rect -4527 -5113 -4467 -5059
rect -4306 -5113 -4246 -5059
rect -4085 -5113 -4025 -5059
rect -3864 -5113 -3804 -5059
rect -3643 -5113 -3583 -5059
rect -3422 -5113 -3362 -5059
rect -3201 -5113 -3141 -5059
rect -2980 -5113 -2950 -5059
rect -4901 -5143 -2950 -5113
rect -2498 -5052 -547 -5022
rect -2498 -5106 -2285 -5052
rect -2124 -5106 -2064 -5052
rect -1903 -5106 -1843 -5052
rect -1682 -5106 -1622 -5052
rect -1461 -5106 -1401 -5052
rect -1240 -5106 -1180 -5052
rect -1019 -5106 -959 -5052
rect -798 -5106 -738 -5052
rect -577 -5106 -547 -5052
rect -2498 -5136 -547 -5106
rect 101 -5051 1648 -5021
rect 101 -5105 131 -5051
rect 292 -5105 352 -5051
rect 513 -5105 573 -5051
rect 734 -5105 794 -5051
rect 955 -5105 1015 -5051
rect 1176 -5105 1236 -5051
rect 1397 -5105 1457 -5051
rect 1618 -5105 1648 -5051
rect 101 -5135 1648 -5105
rect 1861 -5051 3408 -5021
rect 1861 -5105 1891 -5051
rect 2052 -5105 2112 -5051
rect 2273 -5105 2333 -5051
rect 2494 -5105 2554 -5051
rect 2715 -5105 2775 -5051
rect 2936 -5105 2996 -5051
rect 3157 -5105 3217 -5051
rect 3378 -5105 3408 -5051
rect 1861 -5135 3408 -5105
rect 3674 -5051 5221 -5021
rect 3674 -5105 3704 -5051
rect 3865 -5105 3925 -5051
rect 4086 -5105 4146 -5051
rect 4307 -5105 4367 -5051
rect 4528 -5105 4588 -5051
rect 4749 -5105 4809 -5051
rect 4970 -5105 5030 -5051
rect 5191 -5105 5221 -5051
rect 3674 -5135 5221 -5105
rect 5541 -5052 7088 -5022
rect 5541 -5106 5571 -5052
rect 5732 -5106 5792 -5052
rect 5953 -5106 6013 -5052
rect 6174 -5106 6234 -5052
rect 6395 -5106 6455 -5052
rect 6616 -5106 6676 -5052
rect 6837 -5106 6897 -5052
rect 7058 -5106 7088 -5052
rect 5541 -5136 7088 -5106
<< nsubdiff >>
rect -4907 2681 -2950 2711
rect -4907 2627 -4688 2681
rect -4527 2627 -4467 2681
rect -4306 2627 -4246 2681
rect -4085 2627 -4025 2681
rect -3864 2627 -3804 2681
rect -3643 2627 -3583 2681
rect -3422 2627 -3362 2681
rect -3201 2627 -3141 2681
rect -2980 2627 -2950 2681
rect -4907 2597 -2950 2627
rect -2504 2688 -547 2718
rect -2504 2634 -2285 2688
rect -2124 2634 -2064 2688
rect -1903 2634 -1843 2688
rect -1682 2634 -1622 2688
rect -1461 2634 -1401 2688
rect -1240 2634 -1180 2688
rect -1019 2634 -959 2688
rect -798 2634 -738 2688
rect -577 2634 -547 2688
rect -2504 2604 -547 2634
rect 101 2689 1648 2719
rect 101 2635 131 2689
rect 292 2635 352 2689
rect 513 2635 573 2689
rect 734 2635 794 2689
rect 955 2635 1015 2689
rect 1176 2635 1236 2689
rect 1397 2635 1457 2689
rect 1618 2635 1648 2689
rect 101 2605 1648 2635
rect 1861 2689 3408 2719
rect 1861 2635 1891 2689
rect 2052 2635 2112 2689
rect 2273 2635 2333 2689
rect 2494 2635 2554 2689
rect 2715 2635 2775 2689
rect 2936 2635 2996 2689
rect 3157 2635 3217 2689
rect 3378 2635 3408 2689
rect 1861 2605 3408 2635
rect 3674 2689 5221 2719
rect 3674 2635 3704 2689
rect 3865 2635 3925 2689
rect 4086 2635 4146 2689
rect 4307 2635 4367 2689
rect 4528 2635 4588 2689
rect 4749 2635 4809 2689
rect 4970 2635 5030 2689
rect 5191 2635 5221 2689
rect 3674 2605 5221 2635
rect 5541 2688 7088 2718
rect 5541 2634 5571 2688
rect 5732 2634 5792 2688
rect 5953 2634 6013 2688
rect 6174 2634 6234 2688
rect 6395 2634 6455 2688
rect 6616 2634 6676 2688
rect 6837 2634 6897 2688
rect 7058 2634 7088 2688
rect 5541 2604 7088 2634
rect 95 -103 910 -86
rect 95 -163 124 -103
rect 871 -163 910 -103
rect 95 -176 910 -163
rect -4907 -2479 -2950 -2449
rect -4907 -2533 -4688 -2479
rect -4527 -2533 -4467 -2479
rect -4306 -2533 -4246 -2479
rect -4085 -2533 -4025 -2479
rect -3864 -2533 -3804 -2479
rect -3643 -2533 -3583 -2479
rect -3422 -2533 -3362 -2479
rect -3201 -2533 -3141 -2479
rect -2980 -2533 -2950 -2479
rect -4907 -2563 -2950 -2533
rect -2504 -2472 -547 -2442
rect -2504 -2526 -2285 -2472
rect -2124 -2526 -2064 -2472
rect -1903 -2526 -1843 -2472
rect -1682 -2526 -1622 -2472
rect -1461 -2526 -1401 -2472
rect -1240 -2526 -1180 -2472
rect -1019 -2526 -959 -2472
rect -798 -2526 -738 -2472
rect -577 -2526 -547 -2472
rect -2504 -2556 -547 -2526
rect 1861 -2471 3408 -2441
rect 1861 -2525 1891 -2471
rect 2052 -2525 2112 -2471
rect 2273 -2525 2333 -2471
rect 2494 -2525 2554 -2471
rect 2715 -2525 2775 -2471
rect 2936 -2525 2996 -2471
rect 3157 -2525 3217 -2471
rect 3378 -2525 3408 -2471
rect 1861 -2555 3408 -2525
rect 3674 -2471 5221 -2441
rect 3674 -2525 3704 -2471
rect 3865 -2525 3925 -2471
rect 4086 -2525 4146 -2471
rect 4307 -2525 4367 -2471
rect 4528 -2525 4588 -2471
rect 4749 -2525 4809 -2471
rect 4970 -2525 5030 -2471
rect 5191 -2525 5221 -2471
rect 3674 -2555 5221 -2525
rect 5541 -2472 7088 -2442
rect 5541 -2526 5571 -2472
rect 5732 -2526 5792 -2472
rect 5953 -2526 6013 -2472
rect 6174 -2526 6234 -2472
rect 6395 -2526 6455 -2472
rect 6616 -2526 6676 -2472
rect 6837 -2526 6897 -2472
rect 7058 -2526 7088 -2472
rect 5541 -2556 7088 -2526
rect 95 -3044 910 -3027
rect 95 -3104 124 -3044
rect 871 -3104 910 -3044
rect 95 -3121 910 -3104
rect -4907 -7639 -2950 -7609
rect -4907 -7693 -4688 -7639
rect -4527 -7693 -4467 -7639
rect -4306 -7693 -4246 -7639
rect -4085 -7693 -4025 -7639
rect -3864 -7693 -3804 -7639
rect -3643 -7693 -3583 -7639
rect -3422 -7693 -3362 -7639
rect -3201 -7693 -3141 -7639
rect -2980 -7693 -2950 -7639
rect -4907 -7723 -2950 -7693
rect -2504 -7632 -547 -7602
rect -2504 -7686 -2285 -7632
rect -2124 -7686 -2064 -7632
rect -1903 -7686 -1843 -7632
rect -1682 -7686 -1622 -7632
rect -1461 -7686 -1401 -7632
rect -1240 -7686 -1180 -7632
rect -1019 -7686 -959 -7632
rect -798 -7686 -738 -7632
rect -577 -7686 -547 -7632
rect -2504 -7716 -547 -7686
rect 101 -7631 1648 -7601
rect 101 -7685 131 -7631
rect 292 -7685 352 -7631
rect 513 -7685 573 -7631
rect 734 -7685 794 -7631
rect 955 -7685 1015 -7631
rect 1176 -7685 1236 -7631
rect 1397 -7685 1457 -7631
rect 1618 -7685 1648 -7631
rect 101 -7715 1648 -7685
rect 1861 -7631 3408 -7601
rect 1861 -7685 1891 -7631
rect 2052 -7685 2112 -7631
rect 2273 -7685 2333 -7631
rect 2494 -7685 2554 -7631
rect 2715 -7685 2775 -7631
rect 2936 -7685 2996 -7631
rect 3157 -7685 3217 -7631
rect 3378 -7685 3408 -7631
rect 1861 -7715 3408 -7685
rect 3674 -7631 5221 -7601
rect 3674 -7685 3704 -7631
rect 3865 -7685 3925 -7631
rect 4086 -7685 4146 -7631
rect 4307 -7685 4367 -7631
rect 4528 -7685 4588 -7631
rect 4749 -7685 4809 -7631
rect 4970 -7685 5030 -7631
rect 5191 -7685 5221 -7631
rect 3674 -7715 5221 -7685
rect 5541 -7632 7088 -7602
rect 5541 -7686 5571 -7632
rect 5732 -7686 5792 -7632
rect 5953 -7686 6013 -7632
rect 6174 -7686 6234 -7632
rect 6395 -7686 6455 -7632
rect 6616 -7686 6676 -7632
rect 6837 -7686 6897 -7632
rect 7058 -7686 7088 -7632
rect 5541 -7716 7088 -7686
<< psubdiffcont >>
rect -4688 47 -4527 101
rect -4467 47 -4306 101
rect -4246 47 -4085 101
rect -4025 47 -3864 101
rect -3804 47 -3643 101
rect -3583 47 -3422 101
rect -3362 47 -3201 101
rect -3141 47 -2980 101
rect -2285 54 -2124 108
rect -2064 54 -1903 108
rect -1843 54 -1682 108
rect -1622 54 -1461 108
rect -1401 54 -1240 108
rect -1180 54 -1019 108
rect -959 54 -798 108
rect -738 54 -577 108
rect 131 55 292 109
rect 352 55 513 109
rect 573 55 734 109
rect 794 55 955 109
rect 1015 55 1176 109
rect 1236 55 1397 109
rect 1457 55 1618 109
rect 1891 55 2052 109
rect 2112 55 2273 109
rect 2333 55 2494 109
rect 2554 55 2715 109
rect 2775 55 2936 109
rect 2996 55 3157 109
rect 3217 55 3378 109
rect 3704 55 3865 109
rect 3925 55 4086 109
rect 4146 55 4307 109
rect 4367 55 4528 109
rect 4588 55 4749 109
rect 4809 55 4970 109
rect 5030 55 5191 109
rect 5571 54 5732 108
rect 5792 54 5953 108
rect 6013 54 6174 108
rect 6234 54 6395 108
rect 6455 54 6616 108
rect 6676 54 6837 108
rect 6897 54 7058 108
rect 115 -1631 879 -1576
rect 115 -4572 879 -4517
rect -4688 -5113 -4527 -5059
rect -4467 -5113 -4306 -5059
rect -4246 -5113 -4085 -5059
rect -4025 -5113 -3864 -5059
rect -3804 -5113 -3643 -5059
rect -3583 -5113 -3422 -5059
rect -3362 -5113 -3201 -5059
rect -3141 -5113 -2980 -5059
rect -2285 -5106 -2124 -5052
rect -2064 -5106 -1903 -5052
rect -1843 -5106 -1682 -5052
rect -1622 -5106 -1461 -5052
rect -1401 -5106 -1240 -5052
rect -1180 -5106 -1019 -5052
rect -959 -5106 -798 -5052
rect -738 -5106 -577 -5052
rect 131 -5105 292 -5051
rect 352 -5105 513 -5051
rect 573 -5105 734 -5051
rect 794 -5105 955 -5051
rect 1015 -5105 1176 -5051
rect 1236 -5105 1397 -5051
rect 1457 -5105 1618 -5051
rect 1891 -5105 2052 -5051
rect 2112 -5105 2273 -5051
rect 2333 -5105 2494 -5051
rect 2554 -5105 2715 -5051
rect 2775 -5105 2936 -5051
rect 2996 -5105 3157 -5051
rect 3217 -5105 3378 -5051
rect 3704 -5105 3865 -5051
rect 3925 -5105 4086 -5051
rect 4146 -5105 4307 -5051
rect 4367 -5105 4528 -5051
rect 4588 -5105 4749 -5051
rect 4809 -5105 4970 -5051
rect 5030 -5105 5191 -5051
rect 5571 -5106 5732 -5052
rect 5792 -5106 5953 -5052
rect 6013 -5106 6174 -5052
rect 6234 -5106 6395 -5052
rect 6455 -5106 6616 -5052
rect 6676 -5106 6837 -5052
rect 6897 -5106 7058 -5052
<< nsubdiffcont >>
rect -4688 2627 -4527 2681
rect -4467 2627 -4306 2681
rect -4246 2627 -4085 2681
rect -4025 2627 -3864 2681
rect -3804 2627 -3643 2681
rect -3583 2627 -3422 2681
rect -3362 2627 -3201 2681
rect -3141 2627 -2980 2681
rect -2285 2634 -2124 2688
rect -2064 2634 -1903 2688
rect -1843 2634 -1682 2688
rect -1622 2634 -1461 2688
rect -1401 2634 -1240 2688
rect -1180 2634 -1019 2688
rect -959 2634 -798 2688
rect -738 2634 -577 2688
rect 131 2635 292 2689
rect 352 2635 513 2689
rect 573 2635 734 2689
rect 794 2635 955 2689
rect 1015 2635 1176 2689
rect 1236 2635 1397 2689
rect 1457 2635 1618 2689
rect 1891 2635 2052 2689
rect 2112 2635 2273 2689
rect 2333 2635 2494 2689
rect 2554 2635 2715 2689
rect 2775 2635 2936 2689
rect 2996 2635 3157 2689
rect 3217 2635 3378 2689
rect 3704 2635 3865 2689
rect 3925 2635 4086 2689
rect 4146 2635 4307 2689
rect 4367 2635 4528 2689
rect 4588 2635 4749 2689
rect 4809 2635 4970 2689
rect 5030 2635 5191 2689
rect 5571 2634 5732 2688
rect 5792 2634 5953 2688
rect 6013 2634 6174 2688
rect 6234 2634 6395 2688
rect 6455 2634 6616 2688
rect 6676 2634 6837 2688
rect 6897 2634 7058 2688
rect 124 -163 871 -103
rect -4688 -2533 -4527 -2479
rect -4467 -2533 -4306 -2479
rect -4246 -2533 -4085 -2479
rect -4025 -2533 -3864 -2479
rect -3804 -2533 -3643 -2479
rect -3583 -2533 -3422 -2479
rect -3362 -2533 -3201 -2479
rect -3141 -2533 -2980 -2479
rect -2285 -2526 -2124 -2472
rect -2064 -2526 -1903 -2472
rect -1843 -2526 -1682 -2472
rect -1622 -2526 -1461 -2472
rect -1401 -2526 -1240 -2472
rect -1180 -2526 -1019 -2472
rect -959 -2526 -798 -2472
rect -738 -2526 -577 -2472
rect 1891 -2525 2052 -2471
rect 2112 -2525 2273 -2471
rect 2333 -2525 2494 -2471
rect 2554 -2525 2715 -2471
rect 2775 -2525 2936 -2471
rect 2996 -2525 3157 -2471
rect 3217 -2525 3378 -2471
rect 3704 -2525 3865 -2471
rect 3925 -2525 4086 -2471
rect 4146 -2525 4307 -2471
rect 4367 -2525 4528 -2471
rect 4588 -2525 4749 -2471
rect 4809 -2525 4970 -2471
rect 5030 -2525 5191 -2471
rect 5571 -2526 5732 -2472
rect 5792 -2526 5953 -2472
rect 6013 -2526 6174 -2472
rect 6234 -2526 6395 -2472
rect 6455 -2526 6616 -2472
rect 6676 -2526 6837 -2472
rect 6897 -2526 7058 -2472
rect 124 -3104 871 -3044
rect -4688 -7693 -4527 -7639
rect -4467 -7693 -4306 -7639
rect -4246 -7693 -4085 -7639
rect -4025 -7693 -3864 -7639
rect -3804 -7693 -3643 -7639
rect -3583 -7693 -3422 -7639
rect -3362 -7693 -3201 -7639
rect -3141 -7693 -2980 -7639
rect -2285 -7686 -2124 -7632
rect -2064 -7686 -1903 -7632
rect -1843 -7686 -1682 -7632
rect -1622 -7686 -1461 -7632
rect -1401 -7686 -1240 -7632
rect -1180 -7686 -1019 -7632
rect -959 -7686 -798 -7632
rect -738 -7686 -577 -7632
rect 131 -7685 292 -7631
rect 352 -7685 513 -7631
rect 573 -7685 734 -7631
rect 794 -7685 955 -7631
rect 1015 -7685 1176 -7631
rect 1236 -7685 1397 -7631
rect 1457 -7685 1618 -7631
rect 1891 -7685 2052 -7631
rect 2112 -7685 2273 -7631
rect 2333 -7685 2494 -7631
rect 2554 -7685 2715 -7631
rect 2775 -7685 2936 -7631
rect 2996 -7685 3157 -7631
rect 3217 -7685 3378 -7631
rect 3704 -7685 3865 -7631
rect 3925 -7685 4086 -7631
rect 4146 -7685 4307 -7631
rect 4367 -7685 4528 -7631
rect 4588 -7685 4749 -7631
rect 4809 -7685 4970 -7631
rect 5030 -7685 5191 -7631
rect 5571 -7686 5732 -7632
rect 5792 -7686 5953 -7632
rect 6013 -7686 6174 -7632
rect 6234 -7686 6395 -7632
rect 6455 -7686 6616 -7632
rect 6676 -7686 6837 -7632
rect 6897 -7686 7058 -7632
<< polysilicon >>
rect -4757 2426 -4701 2470
rect -4353 2426 -4297 2470
rect -3950 2426 -3894 2470
rect -3790 2426 -3734 2470
rect -3630 2426 -3574 2470
rect -3470 2426 -3414 2470
rect -3310 2426 -3254 2470
rect -3150 2426 -3094 2470
rect -2354 2433 -2298 2477
rect -1950 2433 -1894 2477
rect -1547 2433 -1491 2477
rect -1387 2433 -1331 2477
rect -1227 2433 -1171 2477
rect -1067 2433 -1011 2477
rect -907 2433 -851 2477
rect -747 2433 -691 2477
rect 245 2434 301 2478
rect 648 2434 704 2478
rect 808 2434 864 2478
rect 968 2434 1024 2478
rect 1128 2434 1184 2478
rect 1288 2434 1344 2478
rect 1448 2434 1504 2478
rect 2005 2434 2061 2478
rect 2165 2434 2221 2478
rect 2325 2434 2381 2478
rect 2485 2434 2541 2478
rect 2645 2434 2701 2478
rect 2805 2434 2861 2478
rect 3208 2434 3264 2478
rect 3818 2434 3874 2478
rect 4221 2434 4277 2478
rect 4381 2434 4437 2478
rect 4541 2434 4597 2478
rect 4701 2434 4757 2478
rect 4861 2434 4917 2478
rect 5021 2434 5077 2478
rect 5685 2433 5741 2477
rect 5845 2433 5901 2477
rect 6005 2433 6061 2477
rect 6165 2433 6221 2477
rect 6325 2433 6381 2477
rect 6485 2433 6541 2477
rect 6888 2433 6944 2477
rect -4757 2090 -4701 2226
rect -4353 2090 -4297 2226
rect -4158 2182 -4083 2194
rect -3950 2182 -3894 2226
rect -3790 2182 -3734 2226
rect -3630 2182 -3574 2226
rect -3470 2182 -3414 2226
rect -3310 2182 -3254 2226
rect -3150 2182 -3094 2226
rect -4158 2181 -3094 2182
rect -4158 2135 -4143 2181
rect -4097 2135 -3094 2181
rect -4158 2134 -3094 2135
rect -4158 2120 -4083 2134
rect -3950 2090 -3894 2134
rect -3790 2090 -3734 2134
rect -3630 2090 -3574 2134
rect -3470 2090 -3414 2134
rect -3310 2090 -3254 2134
rect -3150 2090 -3094 2134
rect -2354 2097 -2298 2233
rect -1950 2097 -1894 2233
rect -1755 2189 -1680 2201
rect -1547 2189 -1491 2233
rect -1387 2189 -1331 2233
rect -1227 2189 -1171 2233
rect -1067 2189 -1011 2233
rect -907 2189 -851 2233
rect -747 2189 -691 2233
rect -1755 2188 -691 2189
rect -1755 2142 -1740 2188
rect -1694 2142 -691 2188
rect -1755 2141 -691 2142
rect -1755 2127 -1680 2141
rect -1547 2097 -1491 2141
rect -1387 2097 -1331 2141
rect -1227 2097 -1171 2141
rect -1067 2097 -1011 2141
rect -907 2097 -851 2141
rect -747 2097 -691 2141
rect 245 2098 301 2234
rect 440 2190 515 2202
rect 648 2190 704 2234
rect 808 2190 864 2234
rect 968 2190 1024 2234
rect 1128 2190 1184 2234
rect 1288 2190 1344 2234
rect 1448 2190 1504 2234
rect 440 2189 1504 2190
rect 440 2143 455 2189
rect 501 2143 1504 2189
rect 440 2142 1504 2143
rect 440 2128 515 2142
rect 648 2098 704 2142
rect 808 2098 864 2142
rect 968 2098 1024 2142
rect 1128 2098 1184 2142
rect 1288 2098 1344 2142
rect 1448 2098 1504 2142
rect 2005 2190 2061 2234
rect 2165 2190 2221 2234
rect 2325 2190 2381 2234
rect 2485 2190 2541 2234
rect 2645 2190 2701 2234
rect 2805 2190 2861 2234
rect 2994 2190 3069 2202
rect 2005 2189 3069 2190
rect 2005 2143 3008 2189
rect 3054 2143 3069 2189
rect 2005 2142 3069 2143
rect 2005 2098 2061 2142
rect 2165 2098 2221 2142
rect 2325 2098 2381 2142
rect 2485 2098 2541 2142
rect 2645 2098 2701 2142
rect 2805 2098 2861 2142
rect 2994 2128 3069 2142
rect 3208 2098 3264 2234
rect 3818 2098 3874 2234
rect 4013 2190 4088 2202
rect 4221 2190 4277 2234
rect 4381 2190 4437 2234
rect 4541 2190 4597 2234
rect 4701 2190 4757 2234
rect 4861 2190 4917 2234
rect 5021 2190 5077 2234
rect 4013 2189 5077 2190
rect 4013 2143 4028 2189
rect 4074 2143 5077 2189
rect 4013 2142 5077 2143
rect 4013 2128 4088 2142
rect 4221 2098 4277 2142
rect 4381 2098 4437 2142
rect 4541 2098 4597 2142
rect 4701 2098 4757 2142
rect 4861 2098 4917 2142
rect 5021 2098 5077 2142
rect 5685 2189 5741 2233
rect 5845 2189 5901 2233
rect 6005 2189 6061 2233
rect 6165 2189 6221 2233
rect 6325 2189 6381 2233
rect 6485 2189 6541 2233
rect 6674 2189 6749 2201
rect 5685 2188 6749 2189
rect 5685 2142 6688 2188
rect 6734 2142 6749 2188
rect 5685 2141 6749 2142
rect 5685 2097 5741 2141
rect 5845 2097 5901 2141
rect 6005 2097 6061 2141
rect 6165 2097 6221 2141
rect 6325 2097 6381 2141
rect 6485 2097 6541 2141
rect 6674 2127 6749 2141
rect 6888 2097 6944 2233
rect -4757 1754 -4701 1890
rect -4353 1754 -4297 1890
rect -4158 1846 -4083 1858
rect -3950 1846 -3894 1890
rect -3790 1846 -3734 1890
rect -3630 1846 -3574 1890
rect -3470 1846 -3414 1890
rect -3310 1846 -3254 1890
rect -3150 1846 -3094 1890
rect -4158 1845 -3094 1846
rect -4158 1799 -4143 1845
rect -4097 1799 -3094 1845
rect -4158 1798 -3094 1799
rect -4158 1784 -4083 1798
rect -3950 1754 -3894 1798
rect -3790 1754 -3734 1798
rect -3630 1754 -3574 1798
rect -3470 1754 -3414 1798
rect -3310 1754 -3254 1798
rect -3150 1754 -3094 1798
rect -2354 1761 -2298 1897
rect -1950 1761 -1894 1897
rect -1755 1853 -1680 1865
rect -1547 1853 -1491 1897
rect -1387 1853 -1331 1897
rect -1227 1853 -1171 1897
rect -1067 1853 -1011 1897
rect -907 1853 -851 1897
rect -747 1853 -691 1897
rect -1755 1852 -691 1853
rect -1755 1806 -1740 1852
rect -1694 1806 -691 1852
rect -1755 1805 -691 1806
rect -1755 1791 -1680 1805
rect -1547 1761 -1491 1805
rect -1387 1761 -1331 1805
rect -1227 1761 -1171 1805
rect -1067 1761 -1011 1805
rect -907 1761 -851 1805
rect -747 1761 -691 1805
rect 245 1762 301 1898
rect 440 1854 515 1866
rect 648 1854 704 1898
rect 808 1854 864 1898
rect 968 1854 1024 1898
rect 1128 1854 1184 1898
rect 1288 1854 1344 1898
rect 1448 1854 1504 1898
rect 440 1853 1504 1854
rect 440 1807 455 1853
rect 501 1807 1504 1853
rect 440 1806 1504 1807
rect 440 1792 515 1806
rect 648 1762 704 1806
rect 808 1762 864 1806
rect 968 1762 1024 1806
rect 1128 1762 1184 1806
rect 1288 1762 1344 1806
rect 1448 1762 1504 1806
rect 2005 1854 2061 1898
rect 2165 1854 2221 1898
rect 2325 1854 2381 1898
rect 2485 1854 2541 1898
rect 2645 1854 2701 1898
rect 2805 1854 2861 1898
rect 2994 1854 3069 1866
rect 2005 1853 3069 1854
rect 2005 1807 3008 1853
rect 3054 1807 3069 1853
rect 2005 1806 3069 1807
rect 2005 1762 2061 1806
rect 2165 1762 2221 1806
rect 2325 1762 2381 1806
rect 2485 1762 2541 1806
rect 2645 1762 2701 1806
rect 2805 1762 2861 1806
rect 2994 1792 3069 1806
rect 3208 1762 3264 1898
rect 3818 1762 3874 1898
rect 4013 1854 4088 1866
rect 4221 1854 4277 1898
rect 4381 1854 4437 1898
rect 4541 1854 4597 1898
rect 4701 1854 4757 1898
rect 4861 1854 4917 1898
rect 5021 1854 5077 1898
rect 4013 1853 5077 1854
rect 4013 1807 4028 1853
rect 4074 1807 5077 1853
rect 4013 1806 5077 1807
rect 4013 1792 4088 1806
rect 4221 1762 4277 1806
rect 4381 1762 4437 1806
rect 4541 1762 4597 1806
rect 4701 1762 4757 1806
rect 4861 1762 4917 1806
rect 5021 1762 5077 1806
rect 5685 1853 5741 1897
rect 5845 1853 5901 1897
rect 6005 1853 6061 1897
rect 6165 1853 6221 1897
rect 6325 1853 6381 1897
rect 6485 1853 6541 1897
rect 6674 1853 6749 1865
rect 5685 1852 6749 1853
rect 5685 1806 6688 1852
rect 6734 1806 6749 1852
rect 5685 1805 6749 1806
rect 5685 1761 5741 1805
rect 5845 1761 5901 1805
rect 6005 1761 6061 1805
rect 6165 1761 6221 1805
rect 6325 1761 6381 1805
rect 6485 1761 6541 1805
rect 6674 1791 6749 1805
rect 6888 1761 6944 1897
rect -4757 1418 -4701 1554
rect -4353 1418 -4297 1554
rect -4158 1510 -4083 1522
rect -3950 1510 -3894 1554
rect -3790 1510 -3734 1554
rect -3630 1510 -3574 1554
rect -3470 1510 -3414 1554
rect -3310 1510 -3254 1554
rect -3150 1510 -3094 1554
rect -4158 1509 -3094 1510
rect -4158 1463 -4143 1509
rect -4097 1463 -3094 1509
rect -4158 1462 -3094 1463
rect -4158 1448 -4083 1462
rect -3950 1418 -3894 1462
rect -3790 1418 -3734 1462
rect -3630 1418 -3574 1462
rect -3470 1418 -3414 1462
rect -3310 1418 -3254 1462
rect -3150 1418 -3094 1462
rect -2354 1425 -2298 1561
rect -1950 1425 -1894 1561
rect -1755 1517 -1680 1529
rect -1547 1517 -1491 1561
rect -1387 1517 -1331 1561
rect -1227 1517 -1171 1561
rect -1067 1517 -1011 1561
rect -907 1517 -851 1561
rect -747 1517 -691 1561
rect -1755 1516 -691 1517
rect -1755 1470 -1740 1516
rect -1694 1470 -691 1516
rect -1755 1469 -691 1470
rect -1755 1455 -1680 1469
rect -1547 1425 -1491 1469
rect -1387 1425 -1331 1469
rect -1227 1425 -1171 1469
rect -1067 1425 -1011 1469
rect -907 1425 -851 1469
rect -747 1425 -691 1469
rect 245 1426 301 1562
rect 440 1518 515 1530
rect 648 1518 704 1562
rect 808 1518 864 1562
rect 968 1518 1024 1562
rect 1128 1518 1184 1562
rect 1288 1518 1344 1562
rect 1448 1518 1504 1562
rect 440 1517 1504 1518
rect 440 1471 455 1517
rect 501 1471 1504 1517
rect 440 1470 1504 1471
rect 440 1456 515 1470
rect 648 1426 704 1470
rect 808 1426 864 1470
rect 968 1426 1024 1470
rect 1128 1426 1184 1470
rect 1288 1426 1344 1470
rect 1448 1426 1504 1470
rect 2005 1518 2061 1562
rect 2165 1518 2221 1562
rect 2325 1518 2381 1562
rect 2485 1518 2541 1562
rect 2645 1518 2701 1562
rect 2805 1518 2861 1562
rect 2994 1518 3069 1530
rect 2005 1517 3069 1518
rect 2005 1471 3008 1517
rect 3054 1471 3069 1517
rect 2005 1470 3069 1471
rect 2005 1426 2061 1470
rect 2165 1426 2221 1470
rect 2325 1426 2381 1470
rect 2485 1426 2541 1470
rect 2645 1426 2701 1470
rect 2805 1426 2861 1470
rect 2994 1456 3069 1470
rect 3208 1426 3264 1562
rect 3818 1426 3874 1562
rect 4013 1518 4088 1530
rect 4221 1518 4277 1562
rect 4381 1518 4437 1562
rect 4541 1518 4597 1562
rect 4701 1518 4757 1562
rect 4861 1518 4917 1562
rect 5021 1518 5077 1562
rect 4013 1517 5077 1518
rect 4013 1471 4028 1517
rect 4074 1471 5077 1517
rect 4013 1470 5077 1471
rect 4013 1456 4088 1470
rect 4221 1426 4277 1470
rect 4381 1426 4437 1470
rect 4541 1426 4597 1470
rect 4701 1426 4757 1470
rect 4861 1426 4917 1470
rect 5021 1426 5077 1470
rect 5685 1517 5741 1561
rect 5845 1517 5901 1561
rect 6005 1517 6061 1561
rect 6165 1517 6221 1561
rect 6325 1517 6381 1561
rect 6485 1517 6541 1561
rect 6674 1517 6749 1529
rect 5685 1516 6749 1517
rect 5685 1470 6688 1516
rect 6734 1470 6749 1516
rect 5685 1469 6749 1470
rect 5685 1425 5741 1469
rect 5845 1425 5901 1469
rect 6005 1425 6061 1469
rect 6165 1425 6221 1469
rect 6325 1425 6381 1469
rect 6485 1425 6541 1469
rect 6674 1455 6749 1469
rect 6888 1425 6944 1561
rect -4757 975 -4701 1218
rect -5001 958 -4701 975
rect -5001 912 -4980 958
rect -4934 912 -4882 958
rect -4836 912 -4784 958
rect -4738 912 -4701 958
rect -4353 957 -4297 1218
rect -3950 1147 -3894 1218
rect -3790 1147 -3734 1218
rect -3630 1147 -3574 1218
rect -3470 1147 -3414 1218
rect -3310 1147 -3254 1218
rect -3150 1147 -3094 1218
rect -3950 1097 -3093 1147
rect -2354 982 -2298 1225
rect -5001 895 -4701 912
rect -4757 836 -4701 895
rect -4522 944 -4297 957
rect -4522 936 -4401 944
rect -4522 890 -4508 936
rect -4460 898 -4401 936
rect -4355 898 -4297 944
rect -2598 965 -2298 982
rect -2598 919 -2577 965
rect -2531 919 -2479 965
rect -2433 919 -2381 965
rect -2335 919 -2298 965
rect -1950 964 -1894 1225
rect -1547 1154 -1491 1225
rect -1387 1154 -1331 1225
rect -1227 1154 -1171 1225
rect -1067 1154 -1011 1225
rect -907 1154 -851 1225
rect -747 1154 -691 1225
rect -1547 1104 -690 1154
rect 245 965 301 1226
rect 648 1155 704 1226
rect 808 1155 864 1226
rect 968 1155 1024 1226
rect 1128 1155 1184 1226
rect 1288 1155 1344 1226
rect 1448 1155 1504 1226
rect 2005 1155 2061 1226
rect 2165 1155 2221 1226
rect 2325 1155 2381 1226
rect 2485 1155 2541 1226
rect 2645 1155 2701 1226
rect 2805 1155 2861 1226
rect 648 1105 1505 1155
rect 2004 1105 2861 1155
rect -2598 902 -2298 919
rect -4460 890 -4297 898
rect -4522 885 -4297 890
rect -4522 877 -4446 885
rect -4353 836 -4297 885
rect -3950 836 -3894 880
rect -3790 836 -3734 880
rect -3630 836 -3574 880
rect -3470 836 -3414 880
rect -3310 836 -3254 880
rect -3150 836 -3094 880
rect -2354 843 -2298 902
rect -2119 951 -1894 964
rect -2119 943 -1998 951
rect -2119 897 -2105 943
rect -2057 905 -1998 943
rect -1952 905 -1894 951
rect -2057 897 -1894 905
rect -2119 892 -1894 897
rect -2119 884 -2043 892
rect -1950 843 -1894 892
rect 76 952 301 965
rect 76 944 197 952
rect 76 898 90 944
rect 138 906 197 944
rect 243 906 301 952
rect 138 898 301 906
rect 76 893 301 898
rect -1547 843 -1491 887
rect -1387 843 -1331 887
rect -1227 843 -1171 887
rect -1067 843 -1011 887
rect -907 843 -851 887
rect -747 843 -691 887
rect 76 885 152 893
rect 245 844 301 893
rect 3208 965 3264 1226
rect 3818 965 3874 1226
rect 4221 1155 4277 1226
rect 4381 1155 4437 1226
rect 4541 1155 4597 1226
rect 4701 1155 4757 1226
rect 4861 1155 4917 1226
rect 5021 1155 5077 1226
rect 4221 1105 5078 1155
rect 5685 1154 5741 1225
rect 5845 1154 5901 1225
rect 6005 1154 6061 1225
rect 6165 1154 6221 1225
rect 6325 1154 6381 1225
rect 6485 1154 6541 1225
rect 5684 1104 6541 1154
rect 3208 952 3433 965
rect 3208 906 3266 952
rect 3312 944 3433 952
rect 3312 906 3371 944
rect 3208 898 3371 906
rect 3419 898 3433 944
rect 3208 893 3433 898
rect 648 844 704 888
rect 808 844 864 888
rect 968 844 1024 888
rect 1128 844 1184 888
rect 1288 844 1344 888
rect 1448 844 1504 888
rect 2005 844 2061 888
rect 2165 844 2221 888
rect 2325 844 2381 888
rect 2485 844 2541 888
rect 2645 844 2701 888
rect 2805 844 2861 888
rect 3208 844 3264 893
rect 3357 885 3433 893
rect 3649 952 3874 965
rect 3649 944 3770 952
rect 3649 898 3663 944
rect 3711 906 3770 944
rect 3816 906 3874 952
rect 3711 898 3874 906
rect 3649 893 3874 898
rect 3649 885 3725 893
rect 3818 844 3874 893
rect 6888 964 6944 1225
rect 6888 951 7113 964
rect 6888 905 6946 951
rect 6992 943 7113 951
rect 6992 905 7051 943
rect 6888 897 7051 905
rect 7099 897 7113 943
rect 6888 892 7113 897
rect 4221 844 4277 888
rect 4381 844 4437 888
rect 4541 844 4597 888
rect 4701 844 4757 888
rect 4861 844 4917 888
rect 5021 844 5077 888
rect 5685 843 5741 887
rect 5845 843 5901 887
rect 6005 843 6061 887
rect 6165 843 6221 887
rect 6325 843 6381 887
rect 6485 843 6541 887
rect 6888 843 6944 892
rect 7037 884 7113 892
rect -4757 500 -4701 636
rect -4353 596 -4297 636
rect -3950 596 -3894 636
rect -4353 592 -3894 596
rect -3790 592 -3734 636
rect -3630 592 -3574 636
rect -3470 592 -3414 636
rect -3310 592 -3254 636
rect -3150 592 -3094 636
rect -4353 544 -3094 592
rect -4353 540 -3894 544
rect -4353 500 -4297 540
rect -3950 500 -3894 540
rect -3790 500 -3734 544
rect -3630 500 -3574 544
rect -3470 500 -3414 544
rect -3310 500 -3254 544
rect -3150 500 -3094 544
rect -2354 507 -2298 643
rect -1950 603 -1894 643
rect -1547 603 -1491 643
rect -1950 599 -1491 603
rect -1387 599 -1331 643
rect -1227 599 -1171 643
rect -1067 599 -1011 643
rect -907 599 -851 643
rect -747 599 -691 643
rect -1950 551 -691 599
rect -1950 547 -1491 551
rect -1950 507 -1894 547
rect -1547 507 -1491 547
rect -1387 507 -1331 551
rect -1227 507 -1171 551
rect -1067 507 -1011 551
rect -907 507 -851 551
rect -747 507 -691 551
rect 245 604 301 644
rect 648 604 704 644
rect 245 600 704 604
rect 808 600 864 644
rect 968 600 1024 644
rect 1128 600 1184 644
rect 1288 600 1344 644
rect 1448 600 1504 644
rect 245 552 1504 600
rect 245 548 704 552
rect 245 508 301 548
rect 648 508 704 548
rect 808 508 864 552
rect 968 508 1024 552
rect 1128 508 1184 552
rect 1288 508 1344 552
rect 1448 508 1504 552
rect 2005 600 2061 644
rect 2165 600 2221 644
rect 2325 600 2381 644
rect 2485 600 2541 644
rect 2645 600 2701 644
rect 2805 604 2861 644
rect 3208 604 3264 644
rect 2805 600 3264 604
rect 2005 552 3264 600
rect 2005 508 2061 552
rect 2165 508 2221 552
rect 2325 508 2381 552
rect 2485 508 2541 552
rect 2645 508 2701 552
rect 2805 548 3264 552
rect 2805 508 2861 548
rect 3208 508 3264 548
rect 3818 604 3874 644
rect 4221 604 4277 644
rect 3818 600 4277 604
rect 4381 600 4437 644
rect 4541 600 4597 644
rect 4701 600 4757 644
rect 4861 600 4917 644
rect 5021 600 5077 644
rect 3818 552 5077 600
rect 3818 548 4277 552
rect 3818 508 3874 548
rect 4221 508 4277 548
rect 4381 508 4437 552
rect 4541 508 4597 552
rect 4701 508 4757 552
rect 4861 508 4917 552
rect 5021 508 5077 552
rect 5685 599 5741 643
rect 5845 599 5901 643
rect 6005 599 6061 643
rect 6165 599 6221 643
rect 6325 599 6381 643
rect 6485 603 6541 643
rect 6888 603 6944 643
rect 6485 599 6944 603
rect 5685 551 6944 599
rect 5685 507 5741 551
rect 5845 507 5901 551
rect 6005 507 6061 551
rect 6165 507 6221 551
rect 6325 507 6381 551
rect 6485 547 6944 551
rect 6485 507 6541 547
rect 6888 507 6944 547
rect -4757 256 -4701 300
rect -4353 280 -4297 300
rect -3950 280 -3894 300
rect -3790 280 -3734 300
rect -3630 280 -3574 300
rect -3470 280 -3414 300
rect -3310 280 -3254 300
rect -3150 280 -3094 300
rect -4353 256 -3094 280
rect -2354 263 -2298 307
rect -1950 287 -1894 307
rect -1547 287 -1491 307
rect -1387 287 -1331 307
rect -1227 287 -1171 307
rect -1067 287 -1011 307
rect -907 287 -851 307
rect -747 287 -691 307
rect -1950 263 -691 287
rect 245 288 301 308
rect 648 288 704 308
rect 808 288 864 308
rect 968 288 1024 308
rect 1128 288 1184 308
rect 1288 288 1344 308
rect 1448 288 1504 308
rect 245 264 1504 288
rect 2005 288 2061 308
rect 2165 288 2221 308
rect 2325 288 2381 308
rect 2485 288 2541 308
rect 2645 288 2701 308
rect 2805 288 2861 308
rect 3208 288 3264 308
rect 2005 264 3264 288
rect -4353 224 -3095 256
rect -1950 231 -692 263
rect 245 232 1503 264
rect 2006 232 3264 264
rect 3818 288 3874 308
rect 4221 288 4277 308
rect 4381 288 4437 308
rect 4541 288 4597 308
rect 4701 288 4757 308
rect 4861 288 4917 308
rect 5021 288 5077 308
rect 3818 264 5077 288
rect 5685 287 5741 307
rect 5845 287 5901 307
rect 6005 287 6061 307
rect 6165 287 6221 307
rect 6325 287 6381 307
rect 6485 287 6541 307
rect 6888 287 6944 307
rect 3818 232 5076 264
rect 5685 263 6944 287
rect 5686 231 6944 263
rect -4353 -108 -3095 -76
rect -1950 -101 -692 -69
rect -4757 -152 -4701 -108
rect -4353 -132 -3094 -108
rect -4353 -152 -4297 -132
rect -3950 -152 -3894 -132
rect -3790 -152 -3734 -132
rect -3630 -152 -3574 -132
rect -3470 -152 -3414 -132
rect -3310 -152 -3254 -132
rect -3150 -152 -3094 -132
rect -2354 -145 -2298 -101
rect -1950 -125 -691 -101
rect -1950 -145 -1894 -125
rect -1547 -145 -1491 -125
rect -1387 -145 -1331 -125
rect -1227 -145 -1171 -125
rect -1067 -145 -1011 -125
rect -907 -145 -851 -125
rect -747 -145 -691 -125
rect 2005 -100 3263 -68
rect 3819 -100 5077 -68
rect 2005 -124 3264 -100
rect 2005 -144 2061 -124
rect 2408 -144 2464 -124
rect 2568 -144 2624 -124
rect 2728 -144 2784 -124
rect 2888 -144 2944 -124
rect 3048 -144 3104 -124
rect 3208 -144 3264 -124
rect 3818 -124 5077 -100
rect 3818 -144 3874 -124
rect 3978 -144 4034 -124
rect 4138 -144 4194 -124
rect 4298 -144 4354 -124
rect 4458 -144 4514 -124
rect 4618 -144 4674 -124
rect 5021 -144 5077 -124
rect 5685 -101 6943 -69
rect 5685 -125 6944 -101
rect 235 -330 291 -286
rect 395 -330 451 -286
rect 555 -330 611 -286
rect 715 -330 771 -286
rect -4757 -488 -4701 -352
rect -4353 -392 -4297 -352
rect -3950 -392 -3894 -352
rect -4353 -396 -3894 -392
rect -3790 -396 -3734 -352
rect -3630 -396 -3574 -352
rect -3470 -396 -3414 -352
rect -3310 -396 -3254 -352
rect -3150 -396 -3094 -352
rect -4353 -444 -3094 -396
rect -4353 -448 -3894 -444
rect -4353 -488 -4297 -448
rect -3950 -488 -3894 -448
rect -3790 -488 -3734 -444
rect -3630 -488 -3574 -444
rect -3470 -488 -3414 -444
rect -3310 -488 -3254 -444
rect -3150 -488 -3094 -444
rect -2354 -481 -2298 -345
rect -1950 -385 -1894 -345
rect -1547 -385 -1491 -345
rect -1950 -389 -1491 -385
rect -1387 -389 -1331 -345
rect -1227 -389 -1171 -345
rect -1067 -389 -1011 -345
rect -907 -389 -851 -345
rect -747 -389 -691 -345
rect -1950 -437 -691 -389
rect -1950 -441 -1491 -437
rect -1950 -481 -1894 -441
rect -1547 -481 -1491 -441
rect -1387 -481 -1331 -437
rect -1227 -481 -1171 -437
rect -1067 -481 -1011 -437
rect -907 -481 -851 -437
rect -747 -481 -691 -437
rect 5685 -145 5741 -125
rect 6088 -145 6144 -125
rect 6248 -145 6304 -125
rect 6408 -145 6464 -125
rect 6568 -145 6624 -125
rect 6728 -145 6784 -125
rect 6888 -145 6944 -125
rect 2005 -384 2061 -344
rect 2408 -384 2464 -344
rect 2005 -388 2464 -384
rect 2568 -388 2624 -344
rect 2728 -388 2784 -344
rect 2888 -388 2944 -344
rect 3048 -388 3104 -344
rect 3208 -388 3264 -344
rect 2005 -436 3264 -388
rect 2005 -440 2464 -436
rect 2005 -480 2061 -440
rect 2408 -480 2464 -440
rect 2568 -480 2624 -436
rect 2728 -480 2784 -436
rect 2888 -480 2944 -436
rect 3048 -480 3104 -436
rect 3208 -480 3264 -436
rect 3818 -388 3874 -344
rect 3978 -388 4034 -344
rect 4138 -388 4194 -344
rect 4298 -388 4354 -344
rect 4458 -388 4514 -344
rect 4618 -384 4674 -344
rect 5021 -384 5077 -344
rect 4618 -388 5077 -384
rect 3818 -436 5077 -388
rect 3818 -480 3874 -436
rect 3978 -480 4034 -436
rect 4138 -480 4194 -436
rect 4298 -480 4354 -436
rect 4458 -480 4514 -436
rect 4618 -440 5077 -436
rect 4618 -480 4674 -440
rect 5021 -480 5077 -440
rect 5685 -385 5741 -345
rect 6088 -385 6144 -345
rect 5685 -389 6144 -385
rect 6248 -389 6304 -345
rect 6408 -389 6464 -345
rect 6568 -389 6624 -345
rect 6728 -389 6784 -345
rect 6888 -389 6944 -345
rect 5685 -437 6944 -389
rect 5685 -441 6144 -437
rect 235 -666 291 -530
rect 395 -666 451 -530
rect 555 -666 611 -530
rect 715 -666 771 -530
rect -4757 -747 -4701 -688
rect -5001 -764 -4701 -747
rect -5001 -810 -4980 -764
rect -4934 -810 -4882 -764
rect -4836 -810 -4784 -764
rect -4738 -810 -4701 -764
rect -4522 -737 -4446 -729
rect -4353 -737 -4297 -688
rect -3950 -732 -3894 -688
rect -3790 -732 -3734 -688
rect -3630 -732 -3574 -688
rect -3470 -732 -3414 -688
rect -3310 -732 -3254 -688
rect -3150 -732 -3094 -688
rect -4522 -742 -4297 -737
rect -2354 -740 -2298 -681
rect -4522 -788 -4508 -742
rect -4460 -750 -4297 -742
rect -4460 -788 -4401 -750
rect -4522 -796 -4401 -788
rect -4355 -796 -4297 -750
rect -4522 -809 -4297 -796
rect -5001 -827 -4701 -810
rect -4757 -1070 -4701 -827
rect -4353 -1070 -4297 -809
rect -2598 -757 -2298 -740
rect -2598 -803 -2577 -757
rect -2531 -803 -2479 -757
rect -2433 -803 -2381 -757
rect -2335 -803 -2298 -757
rect -2119 -730 -2043 -722
rect -1950 -730 -1894 -681
rect -1547 -725 -1491 -681
rect -1387 -725 -1331 -681
rect -1227 -725 -1171 -681
rect -1067 -725 -1011 -681
rect -907 -725 -851 -681
rect -747 -725 -691 -681
rect -2119 -735 -1894 -730
rect -2119 -781 -2105 -735
rect -2057 -743 -1894 -735
rect -2057 -781 -1998 -743
rect -2119 -789 -1998 -781
rect -1952 -789 -1894 -743
rect -2119 -802 -1894 -789
rect -2598 -820 -2298 -803
rect -3950 -999 -3093 -949
rect -3950 -1070 -3894 -999
rect -3790 -1070 -3734 -999
rect -3630 -1070 -3574 -999
rect -3470 -1070 -3414 -999
rect -3310 -1070 -3254 -999
rect -3150 -1070 -3094 -999
rect -2354 -1063 -2298 -820
rect -1950 -1063 -1894 -802
rect 5685 -481 5741 -441
rect 6088 -481 6144 -441
rect 6248 -481 6304 -437
rect 6408 -481 6464 -437
rect 6568 -481 6624 -437
rect 6728 -481 6784 -437
rect 6888 -481 6944 -437
rect 1836 -729 1912 -721
rect 2005 -729 2061 -680
rect 2408 -724 2464 -680
rect 2568 -724 2624 -680
rect 2728 -724 2784 -680
rect 2888 -724 2944 -680
rect 3048 -724 3104 -680
rect 3208 -724 3264 -680
rect 3818 -724 3874 -680
rect 3978 -724 4034 -680
rect 4138 -724 4194 -680
rect 4298 -724 4354 -680
rect 4458 -724 4514 -680
rect 4618 -724 4674 -680
rect 1836 -734 2061 -729
rect 1836 -780 1850 -734
rect 1898 -742 2061 -734
rect 1898 -780 1957 -742
rect 1836 -788 1957 -780
rect 2003 -788 2061 -742
rect 1836 -801 2061 -788
rect 235 -910 291 -866
rect 395 -910 451 -866
rect 555 -910 611 -866
rect 715 -910 771 -866
rect -1547 -992 -690 -942
rect 235 -954 771 -910
rect 235 -973 291 -954
rect 189 -986 291 -973
rect -1547 -1063 -1491 -992
rect -1387 -1063 -1331 -992
rect -1227 -1063 -1171 -992
rect -1067 -1063 -1011 -992
rect -907 -1063 -851 -992
rect -747 -1063 -691 -992
rect 189 -1035 205 -986
rect 252 -1035 291 -986
rect 189 -1050 291 -1035
rect 235 -1115 291 -1050
rect 395 -1115 451 -954
rect 555 -1115 611 -954
rect 715 -1115 771 -954
rect 2005 -1062 2061 -801
rect 5021 -729 5077 -680
rect 5170 -729 5246 -721
rect 5021 -734 5246 -729
rect 5021 -742 5184 -734
rect 5021 -788 5079 -742
rect 5125 -780 5184 -742
rect 5232 -780 5246 -734
rect 5125 -788 5246 -780
rect 5021 -801 5246 -788
rect 5516 -730 5592 -722
rect 5685 -730 5741 -681
rect 6088 -725 6144 -681
rect 6248 -725 6304 -681
rect 6408 -725 6464 -681
rect 6568 -725 6624 -681
rect 6728 -725 6784 -681
rect 6888 -725 6944 -681
rect 5516 -735 5741 -730
rect 5516 -781 5530 -735
rect 5578 -743 5741 -735
rect 5578 -781 5637 -743
rect 5516 -789 5637 -781
rect 5683 -789 5741 -743
rect 2408 -991 3265 -941
rect 3817 -991 4674 -941
rect 2408 -1062 2464 -991
rect 2568 -1062 2624 -991
rect 2728 -1062 2784 -991
rect 2888 -1062 2944 -991
rect 3048 -1062 3104 -991
rect 3208 -1062 3264 -991
rect 3818 -1062 3874 -991
rect 3978 -1062 4034 -991
rect 4138 -1062 4194 -991
rect 4298 -1062 4354 -991
rect 4458 -1062 4514 -991
rect 4618 -1062 4674 -991
rect 5021 -1062 5077 -801
rect 5516 -802 5741 -789
rect -4757 -1406 -4701 -1270
rect -4353 -1406 -4297 -1270
rect -4158 -1314 -4083 -1300
rect -3950 -1314 -3894 -1270
rect -3790 -1314 -3734 -1270
rect -3630 -1314 -3574 -1270
rect -3470 -1314 -3414 -1270
rect -3310 -1314 -3254 -1270
rect -3150 -1314 -3094 -1270
rect -4158 -1315 -3094 -1314
rect -4158 -1361 -4143 -1315
rect -4097 -1361 -3094 -1315
rect -4158 -1362 -3094 -1361
rect -4158 -1374 -4083 -1362
rect -3950 -1406 -3894 -1362
rect -3790 -1406 -3734 -1362
rect -3630 -1406 -3574 -1362
rect -3470 -1406 -3414 -1362
rect -3310 -1406 -3254 -1362
rect -3150 -1406 -3094 -1362
rect -2354 -1399 -2298 -1263
rect -1950 -1399 -1894 -1263
rect -1755 -1307 -1680 -1293
rect -1547 -1307 -1491 -1263
rect -1387 -1307 -1331 -1263
rect -1227 -1307 -1171 -1263
rect -1067 -1307 -1011 -1263
rect -907 -1307 -851 -1263
rect -747 -1307 -691 -1263
rect -1755 -1308 -691 -1307
rect -1755 -1354 -1740 -1308
rect -1694 -1354 -691 -1308
rect 235 -1351 291 -1215
rect 395 -1351 451 -1215
rect 555 -1351 611 -1215
rect 715 -1351 771 -1215
rect 5685 -1063 5741 -802
rect 6088 -992 6945 -942
rect 6088 -1063 6144 -992
rect 6248 -1063 6304 -992
rect 6408 -1063 6464 -992
rect 6568 -1063 6624 -992
rect 6728 -1063 6784 -992
rect 6888 -1063 6944 -992
rect -1755 -1355 -691 -1354
rect -1755 -1367 -1680 -1355
rect -1547 -1399 -1491 -1355
rect -1387 -1399 -1331 -1355
rect -1227 -1399 -1171 -1355
rect -1067 -1399 -1011 -1355
rect -907 -1399 -851 -1355
rect -747 -1399 -691 -1355
rect 2005 -1398 2061 -1262
rect 2200 -1306 2275 -1292
rect 2408 -1306 2464 -1262
rect 2568 -1306 2624 -1262
rect 2728 -1306 2784 -1262
rect 2888 -1306 2944 -1262
rect 3048 -1306 3104 -1262
rect 3208 -1306 3264 -1262
rect 2200 -1307 3264 -1306
rect 2200 -1353 2215 -1307
rect 2261 -1353 3264 -1307
rect 2200 -1354 3264 -1353
rect 2200 -1366 2275 -1354
rect 2408 -1398 2464 -1354
rect 2568 -1398 2624 -1354
rect 2728 -1398 2784 -1354
rect 2888 -1398 2944 -1354
rect 3048 -1398 3104 -1354
rect 3208 -1398 3264 -1354
rect 3818 -1306 3874 -1262
rect 3978 -1306 4034 -1262
rect 4138 -1306 4194 -1262
rect 4298 -1306 4354 -1262
rect 4458 -1306 4514 -1262
rect 4618 -1306 4674 -1262
rect 4807 -1306 4882 -1292
rect 3818 -1307 4882 -1306
rect 3818 -1353 4821 -1307
rect 4867 -1353 4882 -1307
rect 3818 -1354 4882 -1353
rect 3818 -1398 3874 -1354
rect 3978 -1398 4034 -1354
rect 4138 -1398 4194 -1354
rect 4298 -1398 4354 -1354
rect 4458 -1398 4514 -1354
rect 4618 -1398 4674 -1354
rect 4807 -1366 4882 -1354
rect 5021 -1398 5077 -1262
rect 235 -1495 291 -1451
rect 395 -1495 451 -1451
rect 555 -1495 611 -1451
rect 715 -1495 771 -1451
rect -4757 -1742 -4701 -1606
rect -4353 -1742 -4297 -1606
rect -4158 -1650 -4083 -1636
rect -3950 -1650 -3894 -1606
rect -3790 -1650 -3734 -1606
rect -3630 -1650 -3574 -1606
rect -3470 -1650 -3414 -1606
rect -3310 -1650 -3254 -1606
rect -3150 -1650 -3094 -1606
rect -4158 -1651 -3094 -1650
rect -4158 -1697 -4143 -1651
rect -4097 -1697 -3094 -1651
rect -4158 -1698 -3094 -1697
rect -4158 -1710 -4083 -1698
rect -3950 -1742 -3894 -1698
rect -3790 -1742 -3734 -1698
rect -3630 -1742 -3574 -1698
rect -3470 -1742 -3414 -1698
rect -3310 -1742 -3254 -1698
rect -3150 -1742 -3094 -1698
rect -2354 -1735 -2298 -1599
rect -1950 -1735 -1894 -1599
rect -1755 -1643 -1680 -1629
rect -1547 -1643 -1491 -1599
rect -1387 -1643 -1331 -1599
rect -1227 -1643 -1171 -1599
rect -1067 -1643 -1011 -1599
rect -907 -1643 -851 -1599
rect -747 -1643 -691 -1599
rect -1755 -1644 -691 -1643
rect -1755 -1690 -1740 -1644
rect -1694 -1690 -691 -1644
rect 5685 -1399 5741 -1263
rect 5880 -1307 5955 -1293
rect 6088 -1307 6144 -1263
rect 6248 -1307 6304 -1263
rect 6408 -1307 6464 -1263
rect 6568 -1307 6624 -1263
rect 6728 -1307 6784 -1263
rect 6888 -1307 6944 -1263
rect 5880 -1308 6944 -1307
rect 5880 -1354 5895 -1308
rect 5941 -1354 6944 -1308
rect 5880 -1355 6944 -1354
rect 5880 -1367 5955 -1355
rect 6088 -1399 6144 -1355
rect 6248 -1399 6304 -1355
rect 6408 -1399 6464 -1355
rect 6568 -1399 6624 -1355
rect 6728 -1399 6784 -1355
rect 6888 -1399 6944 -1355
rect -1755 -1691 -691 -1690
rect -1755 -1703 -1680 -1691
rect -1547 -1735 -1491 -1691
rect -1387 -1735 -1331 -1691
rect -1227 -1735 -1171 -1691
rect -1067 -1735 -1011 -1691
rect -907 -1735 -851 -1691
rect -747 -1735 -691 -1691
rect 235 -1756 291 -1712
rect 395 -1756 451 -1712
rect 555 -1756 611 -1712
rect 715 -1756 771 -1712
rect 2005 -1734 2061 -1598
rect 2200 -1642 2275 -1628
rect 2408 -1642 2464 -1598
rect 2568 -1642 2624 -1598
rect 2728 -1642 2784 -1598
rect 2888 -1642 2944 -1598
rect 3048 -1642 3104 -1598
rect 3208 -1642 3264 -1598
rect 2200 -1643 3264 -1642
rect 2200 -1689 2215 -1643
rect 2261 -1689 3264 -1643
rect 2200 -1690 3264 -1689
rect 2200 -1702 2275 -1690
rect 2408 -1734 2464 -1690
rect 2568 -1734 2624 -1690
rect 2728 -1734 2784 -1690
rect 2888 -1734 2944 -1690
rect 3048 -1734 3104 -1690
rect 3208 -1734 3264 -1690
rect 3818 -1642 3874 -1598
rect 3978 -1642 4034 -1598
rect 4138 -1642 4194 -1598
rect 4298 -1642 4354 -1598
rect 4458 -1642 4514 -1598
rect 4618 -1642 4674 -1598
rect 4807 -1642 4882 -1628
rect 3818 -1643 4882 -1642
rect 3818 -1689 4821 -1643
rect 4867 -1689 4882 -1643
rect 3818 -1690 4882 -1689
rect 3818 -1734 3874 -1690
rect 3978 -1734 4034 -1690
rect 4138 -1734 4194 -1690
rect 4298 -1734 4354 -1690
rect 4458 -1734 4514 -1690
rect 4618 -1734 4674 -1690
rect 4807 -1702 4882 -1690
rect 5021 -1734 5077 -1598
rect -4757 -2078 -4701 -1942
rect -4353 -2078 -4297 -1942
rect -4158 -1986 -4083 -1972
rect -3950 -1986 -3894 -1942
rect -3790 -1986 -3734 -1942
rect -3630 -1986 -3574 -1942
rect -3470 -1986 -3414 -1942
rect -3310 -1986 -3254 -1942
rect -3150 -1986 -3094 -1942
rect -4158 -1987 -3094 -1986
rect -4158 -2033 -4143 -1987
rect -4097 -2033 -3094 -1987
rect -4158 -2034 -3094 -2033
rect -4158 -2046 -4083 -2034
rect -3950 -2078 -3894 -2034
rect -3790 -2078 -3734 -2034
rect -3630 -2078 -3574 -2034
rect -3470 -2078 -3414 -2034
rect -3310 -2078 -3254 -2034
rect -3150 -2078 -3094 -2034
rect -2354 -2071 -2298 -1935
rect -1950 -2071 -1894 -1935
rect -1755 -1979 -1680 -1965
rect -1547 -1979 -1491 -1935
rect -1387 -1979 -1331 -1935
rect -1227 -1979 -1171 -1935
rect -1067 -1979 -1011 -1935
rect -907 -1979 -851 -1935
rect -747 -1979 -691 -1935
rect -1755 -1980 -691 -1979
rect -1755 -2026 -1740 -1980
rect -1694 -2026 -691 -1980
rect 235 -1992 291 -1856
rect 395 -1992 451 -1856
rect 555 -1992 611 -1856
rect 715 -1992 771 -1856
rect 5685 -1735 5741 -1599
rect 5880 -1643 5955 -1629
rect 6088 -1643 6144 -1599
rect 6248 -1643 6304 -1599
rect 6408 -1643 6464 -1599
rect 6568 -1643 6624 -1599
rect 6728 -1643 6784 -1599
rect 6888 -1643 6944 -1599
rect 5880 -1644 6944 -1643
rect 5880 -1690 5895 -1644
rect 5941 -1690 6944 -1644
rect 5880 -1691 6944 -1690
rect 5880 -1703 5955 -1691
rect 6088 -1735 6144 -1691
rect 6248 -1735 6304 -1691
rect 6408 -1735 6464 -1691
rect 6568 -1735 6624 -1691
rect 6728 -1735 6784 -1691
rect 6888 -1735 6944 -1691
rect -1755 -2027 -691 -2026
rect -1755 -2039 -1680 -2027
rect -1547 -2071 -1491 -2027
rect -1387 -2071 -1331 -2027
rect -1227 -2071 -1171 -2027
rect -1067 -2071 -1011 -2027
rect -907 -2071 -851 -2027
rect -747 -2071 -691 -2027
rect 2005 -2070 2061 -1934
rect 2200 -1978 2275 -1964
rect 2408 -1978 2464 -1934
rect 2568 -1978 2624 -1934
rect 2728 -1978 2784 -1934
rect 2888 -1978 2944 -1934
rect 3048 -1978 3104 -1934
rect 3208 -1978 3264 -1934
rect 2200 -1979 3264 -1978
rect 2200 -2025 2215 -1979
rect 2261 -2025 3264 -1979
rect 2200 -2026 3264 -2025
rect 2200 -2038 2275 -2026
rect 2408 -2070 2464 -2026
rect 2568 -2070 2624 -2026
rect 2728 -2070 2784 -2026
rect 2888 -2070 2944 -2026
rect 3048 -2070 3104 -2026
rect 3208 -2070 3264 -2026
rect 3818 -1978 3874 -1934
rect 3978 -1978 4034 -1934
rect 4138 -1978 4194 -1934
rect 4298 -1978 4354 -1934
rect 4458 -1978 4514 -1934
rect 4618 -1978 4674 -1934
rect 4807 -1978 4882 -1964
rect 3818 -1979 4882 -1978
rect 3818 -2025 4821 -1979
rect 4867 -2025 4882 -1979
rect 3818 -2026 4882 -2025
rect 3818 -2070 3874 -2026
rect 3978 -2070 4034 -2026
rect 4138 -2070 4194 -2026
rect 4298 -2070 4354 -2026
rect 4458 -2070 4514 -2026
rect 4618 -2070 4674 -2026
rect 4807 -2038 4882 -2026
rect 5021 -2070 5077 -1934
rect 235 -2157 291 -2092
rect 189 -2172 291 -2157
rect 189 -2221 205 -2172
rect 252 -2221 291 -2172
rect 189 -2234 291 -2221
rect 235 -2253 291 -2234
rect 395 -2253 451 -2092
rect 555 -2253 611 -2092
rect 715 -2253 771 -2092
rect -4757 -2322 -4701 -2278
rect -4353 -2322 -4297 -2278
rect -3950 -2322 -3894 -2278
rect -3790 -2322 -3734 -2278
rect -3630 -2322 -3574 -2278
rect -3470 -2322 -3414 -2278
rect -3310 -2322 -3254 -2278
rect -3150 -2322 -3094 -2278
rect -2354 -2315 -2298 -2271
rect -1950 -2315 -1894 -2271
rect -1547 -2315 -1491 -2271
rect -1387 -2315 -1331 -2271
rect -1227 -2315 -1171 -2271
rect -1067 -2315 -1011 -2271
rect -907 -2315 -851 -2271
rect -747 -2315 -691 -2271
rect 235 -2297 771 -2253
rect 5685 -2071 5741 -1935
rect 5880 -1979 5955 -1965
rect 6088 -1979 6144 -1935
rect 6248 -1979 6304 -1935
rect 6408 -1979 6464 -1935
rect 6568 -1979 6624 -1935
rect 6728 -1979 6784 -1935
rect 6888 -1979 6944 -1935
rect 5880 -1980 6944 -1979
rect 5880 -2026 5895 -1980
rect 5941 -2026 6944 -1980
rect 5880 -2027 6944 -2026
rect 5880 -2039 5955 -2027
rect 6088 -2071 6144 -2027
rect 6248 -2071 6304 -2027
rect 6408 -2071 6464 -2027
rect 6568 -2071 6624 -2027
rect 6728 -2071 6784 -2027
rect 6888 -2071 6944 -2027
rect 235 -2341 291 -2297
rect 395 -2341 451 -2297
rect 555 -2341 611 -2297
rect 715 -2341 771 -2297
rect 2005 -2314 2061 -2270
rect 2408 -2314 2464 -2270
rect 2568 -2314 2624 -2270
rect 2728 -2314 2784 -2270
rect 2888 -2314 2944 -2270
rect 3048 -2314 3104 -2270
rect 3208 -2314 3264 -2270
rect 3818 -2314 3874 -2270
rect 3978 -2314 4034 -2270
rect 4138 -2314 4194 -2270
rect 4298 -2314 4354 -2270
rect 4458 -2314 4514 -2270
rect 4618 -2314 4674 -2270
rect 5021 -2314 5077 -2270
rect 5685 -2315 5741 -2271
rect 6088 -2315 6144 -2271
rect 6248 -2315 6304 -2271
rect 6408 -2315 6464 -2271
rect 6568 -2315 6624 -2271
rect 6728 -2315 6784 -2271
rect 6888 -2315 6944 -2271
rect 235 -2677 291 -2541
rect 395 -2677 451 -2541
rect 555 -2677 611 -2541
rect 715 -2677 771 -2541
rect -4757 -2734 -4701 -2690
rect -4353 -2734 -4297 -2690
rect -3950 -2734 -3894 -2690
rect -3790 -2734 -3734 -2690
rect -3630 -2734 -3574 -2690
rect -3470 -2734 -3414 -2690
rect -3310 -2734 -3254 -2690
rect -3150 -2734 -3094 -2690
rect -2354 -2727 -2298 -2683
rect -1950 -2727 -1894 -2683
rect -1547 -2727 -1491 -2683
rect -1387 -2727 -1331 -2683
rect -1227 -2727 -1171 -2683
rect -1067 -2727 -1011 -2683
rect -907 -2727 -851 -2683
rect -747 -2727 -691 -2683
rect 2005 -2726 2061 -2682
rect 2408 -2726 2464 -2682
rect 2568 -2726 2624 -2682
rect 2728 -2726 2784 -2682
rect 2888 -2726 2944 -2682
rect 3048 -2726 3104 -2682
rect 3208 -2726 3264 -2682
rect 3818 -2726 3874 -2682
rect 3978 -2726 4034 -2682
rect 4138 -2726 4194 -2682
rect 4298 -2726 4354 -2682
rect 4458 -2726 4514 -2682
rect 4618 -2726 4674 -2682
rect 5021 -2726 5077 -2682
rect 235 -2921 291 -2877
rect 395 -2921 451 -2877
rect 555 -2921 611 -2877
rect 715 -2921 771 -2877
rect 5685 -2727 5741 -2683
rect 6088 -2727 6144 -2683
rect 6248 -2727 6304 -2683
rect 6408 -2727 6464 -2683
rect 6568 -2727 6624 -2683
rect 6728 -2727 6784 -2683
rect 6888 -2727 6944 -2683
rect -4757 -3070 -4701 -2934
rect -4353 -3070 -4297 -2934
rect -4158 -2978 -4083 -2966
rect -3950 -2978 -3894 -2934
rect -3790 -2978 -3734 -2934
rect -3630 -2978 -3574 -2934
rect -3470 -2978 -3414 -2934
rect -3310 -2978 -3254 -2934
rect -3150 -2978 -3094 -2934
rect -4158 -2979 -3094 -2978
rect -4158 -3025 -4143 -2979
rect -4097 -3025 -3094 -2979
rect -4158 -3026 -3094 -3025
rect -4158 -3040 -4083 -3026
rect -3950 -3070 -3894 -3026
rect -3790 -3070 -3734 -3026
rect -3630 -3070 -3574 -3026
rect -3470 -3070 -3414 -3026
rect -3310 -3070 -3254 -3026
rect -3150 -3070 -3094 -3026
rect -2354 -3063 -2298 -2927
rect -1950 -3063 -1894 -2927
rect -1755 -2971 -1680 -2959
rect -1547 -2971 -1491 -2927
rect -1387 -2971 -1331 -2927
rect -1227 -2971 -1171 -2927
rect -1067 -2971 -1011 -2927
rect -907 -2971 -851 -2927
rect -747 -2971 -691 -2927
rect -1755 -2972 -691 -2971
rect -1755 -3018 -1740 -2972
rect -1694 -3018 -691 -2972
rect -1755 -3019 -691 -3018
rect -1755 -3033 -1680 -3019
rect -1547 -3063 -1491 -3019
rect -1387 -3063 -1331 -3019
rect -1227 -3063 -1171 -3019
rect -1067 -3063 -1011 -3019
rect -907 -3063 -851 -3019
rect -747 -3063 -691 -3019
rect 2005 -3062 2061 -2926
rect 2200 -2970 2275 -2958
rect 2408 -2970 2464 -2926
rect 2568 -2970 2624 -2926
rect 2728 -2970 2784 -2926
rect 2888 -2970 2944 -2926
rect 3048 -2970 3104 -2926
rect 3208 -2970 3264 -2926
rect 2200 -2971 3264 -2970
rect 2200 -3017 2215 -2971
rect 2261 -3017 3264 -2971
rect 2200 -3018 3264 -3017
rect 2200 -3032 2275 -3018
rect 2408 -3062 2464 -3018
rect 2568 -3062 2624 -3018
rect 2728 -3062 2784 -3018
rect 2888 -3062 2944 -3018
rect 3048 -3062 3104 -3018
rect 3208 -3062 3264 -3018
rect 3818 -2970 3874 -2926
rect 3978 -2970 4034 -2926
rect 4138 -2970 4194 -2926
rect 4298 -2970 4354 -2926
rect 4458 -2970 4514 -2926
rect 4618 -2970 4674 -2926
rect 4807 -2970 4882 -2958
rect 3818 -2971 4882 -2970
rect 3818 -3017 4821 -2971
rect 4867 -3017 4882 -2971
rect 3818 -3018 4882 -3017
rect 3818 -3062 3874 -3018
rect 3978 -3062 4034 -3018
rect 4138 -3062 4194 -3018
rect 4298 -3062 4354 -3018
rect 4458 -3062 4514 -3018
rect 4618 -3062 4674 -3018
rect 4807 -3032 4882 -3018
rect 5021 -3062 5077 -2926
rect -4757 -3406 -4701 -3270
rect -4353 -3406 -4297 -3270
rect -4158 -3314 -4083 -3302
rect -3950 -3314 -3894 -3270
rect -3790 -3314 -3734 -3270
rect -3630 -3314 -3574 -3270
rect -3470 -3314 -3414 -3270
rect -3310 -3314 -3254 -3270
rect -3150 -3314 -3094 -3270
rect -4158 -3315 -3094 -3314
rect -4158 -3361 -4143 -3315
rect -4097 -3361 -3094 -3315
rect -4158 -3362 -3094 -3361
rect -4158 -3376 -4083 -3362
rect -3950 -3406 -3894 -3362
rect -3790 -3406 -3734 -3362
rect -3630 -3406 -3574 -3362
rect -3470 -3406 -3414 -3362
rect -3310 -3406 -3254 -3362
rect -3150 -3406 -3094 -3362
rect -2354 -3399 -2298 -3263
rect -1950 -3399 -1894 -3263
rect -1755 -3307 -1680 -3295
rect -1547 -3307 -1491 -3263
rect -1387 -3307 -1331 -3263
rect -1227 -3307 -1171 -3263
rect -1067 -3307 -1011 -3263
rect -907 -3307 -851 -3263
rect -747 -3307 -691 -3263
rect 235 -3271 291 -3227
rect 395 -3271 451 -3227
rect 555 -3271 611 -3227
rect 715 -3271 771 -3227
rect 5685 -3063 5741 -2927
rect 5880 -2971 5955 -2959
rect 6088 -2971 6144 -2927
rect 6248 -2971 6304 -2927
rect 6408 -2971 6464 -2927
rect 6568 -2971 6624 -2927
rect 6728 -2971 6784 -2927
rect 6888 -2971 6944 -2927
rect 5880 -2972 6944 -2971
rect 5880 -3018 5895 -2972
rect 5941 -3018 6944 -2972
rect 5880 -3019 6944 -3018
rect 5880 -3033 5955 -3019
rect 6088 -3063 6144 -3019
rect 6248 -3063 6304 -3019
rect 6408 -3063 6464 -3019
rect 6568 -3063 6624 -3019
rect 6728 -3063 6784 -3019
rect 6888 -3063 6944 -3019
rect -1755 -3308 -691 -3307
rect -1755 -3354 -1740 -3308
rect -1694 -3354 -691 -3308
rect -1755 -3355 -691 -3354
rect -1755 -3369 -1680 -3355
rect -1547 -3399 -1491 -3355
rect -1387 -3399 -1331 -3355
rect -1227 -3399 -1171 -3355
rect -1067 -3399 -1011 -3355
rect -907 -3399 -851 -3355
rect -747 -3399 -691 -3355
rect 2005 -3398 2061 -3262
rect 2200 -3306 2275 -3294
rect 2408 -3306 2464 -3262
rect 2568 -3306 2624 -3262
rect 2728 -3306 2784 -3262
rect 2888 -3306 2944 -3262
rect 3048 -3306 3104 -3262
rect 3208 -3306 3264 -3262
rect 2200 -3307 3264 -3306
rect 2200 -3353 2215 -3307
rect 2261 -3353 3264 -3307
rect 2200 -3354 3264 -3353
rect 2200 -3368 2275 -3354
rect 2408 -3398 2464 -3354
rect 2568 -3398 2624 -3354
rect 2728 -3398 2784 -3354
rect 2888 -3398 2944 -3354
rect 3048 -3398 3104 -3354
rect 3208 -3398 3264 -3354
rect 3818 -3306 3874 -3262
rect 3978 -3306 4034 -3262
rect 4138 -3306 4194 -3262
rect 4298 -3306 4354 -3262
rect 4458 -3306 4514 -3262
rect 4618 -3306 4674 -3262
rect 4807 -3306 4882 -3294
rect 3818 -3307 4882 -3306
rect 3818 -3353 4821 -3307
rect 4867 -3353 4882 -3307
rect 3818 -3354 4882 -3353
rect 3818 -3398 3874 -3354
rect 3978 -3398 4034 -3354
rect 4138 -3398 4194 -3354
rect 4298 -3398 4354 -3354
rect 4458 -3398 4514 -3354
rect 4618 -3398 4674 -3354
rect 4807 -3368 4882 -3354
rect 5021 -3398 5077 -3262
rect -4757 -3742 -4701 -3606
rect -4353 -3742 -4297 -3606
rect -4158 -3650 -4083 -3638
rect -3950 -3650 -3894 -3606
rect -3790 -3650 -3734 -3606
rect -3630 -3650 -3574 -3606
rect -3470 -3650 -3414 -3606
rect -3310 -3650 -3254 -3606
rect -3150 -3650 -3094 -3606
rect -4158 -3651 -3094 -3650
rect -4158 -3697 -4143 -3651
rect -4097 -3697 -3094 -3651
rect -4158 -3698 -3094 -3697
rect -4158 -3712 -4083 -3698
rect -3950 -3742 -3894 -3698
rect -3790 -3742 -3734 -3698
rect -3630 -3742 -3574 -3698
rect -3470 -3742 -3414 -3698
rect -3310 -3742 -3254 -3698
rect -3150 -3742 -3094 -3698
rect -2354 -3735 -2298 -3599
rect -1950 -3735 -1894 -3599
rect -1755 -3643 -1680 -3631
rect -1547 -3643 -1491 -3599
rect -1387 -3643 -1331 -3599
rect -1227 -3643 -1171 -3599
rect -1067 -3643 -1011 -3599
rect -907 -3643 -851 -3599
rect -747 -3643 -691 -3599
rect 235 -3607 291 -3471
rect 395 -3607 451 -3471
rect 555 -3607 611 -3471
rect 715 -3607 771 -3471
rect 5685 -3399 5741 -3263
rect 5880 -3307 5955 -3295
rect 6088 -3307 6144 -3263
rect 6248 -3307 6304 -3263
rect 6408 -3307 6464 -3263
rect 6568 -3307 6624 -3263
rect 6728 -3307 6784 -3263
rect 6888 -3307 6944 -3263
rect 5880 -3308 6944 -3307
rect 5880 -3354 5895 -3308
rect 5941 -3354 6944 -3308
rect 5880 -3355 6944 -3354
rect 5880 -3369 5955 -3355
rect 6088 -3399 6144 -3355
rect 6248 -3399 6304 -3355
rect 6408 -3399 6464 -3355
rect 6568 -3399 6624 -3355
rect 6728 -3399 6784 -3355
rect 6888 -3399 6944 -3355
rect -1755 -3644 -691 -3643
rect -1755 -3690 -1740 -3644
rect -1694 -3690 -691 -3644
rect -1755 -3691 -691 -3690
rect -1755 -3705 -1680 -3691
rect -1547 -3735 -1491 -3691
rect -1387 -3735 -1331 -3691
rect -1227 -3735 -1171 -3691
rect -1067 -3735 -1011 -3691
rect -907 -3735 -851 -3691
rect -747 -3735 -691 -3691
rect 2005 -3734 2061 -3598
rect 2200 -3642 2275 -3630
rect 2408 -3642 2464 -3598
rect 2568 -3642 2624 -3598
rect 2728 -3642 2784 -3598
rect 2888 -3642 2944 -3598
rect 3048 -3642 3104 -3598
rect 3208 -3642 3264 -3598
rect 2200 -3643 3264 -3642
rect 2200 -3689 2215 -3643
rect 2261 -3689 3264 -3643
rect 2200 -3690 3264 -3689
rect 2200 -3704 2275 -3690
rect 2408 -3734 2464 -3690
rect 2568 -3734 2624 -3690
rect 2728 -3734 2784 -3690
rect 2888 -3734 2944 -3690
rect 3048 -3734 3104 -3690
rect 3208 -3734 3264 -3690
rect 3818 -3642 3874 -3598
rect 3978 -3642 4034 -3598
rect 4138 -3642 4194 -3598
rect 4298 -3642 4354 -3598
rect 4458 -3642 4514 -3598
rect 4618 -3642 4674 -3598
rect 4807 -3642 4882 -3630
rect 3818 -3643 4882 -3642
rect 3818 -3689 4821 -3643
rect 4867 -3689 4882 -3643
rect 3818 -3690 4882 -3689
rect 3818 -3734 3874 -3690
rect 3978 -3734 4034 -3690
rect 4138 -3734 4194 -3690
rect 4298 -3734 4354 -3690
rect 4458 -3734 4514 -3690
rect 4618 -3734 4674 -3690
rect 4807 -3704 4882 -3690
rect 5021 -3734 5077 -3598
rect 235 -3851 291 -3807
rect 395 -3851 451 -3807
rect 555 -3851 611 -3807
rect 715 -3851 771 -3807
rect 235 -3895 771 -3851
rect 235 -3914 291 -3895
rect 189 -3927 291 -3914
rect -4757 -4185 -4701 -3942
rect -5001 -4202 -4701 -4185
rect -5001 -4248 -4980 -4202
rect -4934 -4248 -4882 -4202
rect -4836 -4248 -4784 -4202
rect -4738 -4248 -4701 -4202
rect -4353 -4203 -4297 -3942
rect -3950 -4013 -3894 -3942
rect -3790 -4013 -3734 -3942
rect -3630 -4013 -3574 -3942
rect -3470 -4013 -3414 -3942
rect -3310 -4013 -3254 -3942
rect -3150 -4013 -3094 -3942
rect -3950 -4063 -3093 -4013
rect -2354 -4178 -2298 -3935
rect -5001 -4265 -4701 -4248
rect -4757 -4324 -4701 -4265
rect -4522 -4216 -4297 -4203
rect -4522 -4224 -4401 -4216
rect -4522 -4270 -4508 -4224
rect -4460 -4262 -4401 -4224
rect -4355 -4262 -4297 -4216
rect -2598 -4195 -2298 -4178
rect -2598 -4241 -2577 -4195
rect -2531 -4241 -2479 -4195
rect -2433 -4241 -2381 -4195
rect -2335 -4241 -2298 -4195
rect -1950 -4196 -1894 -3935
rect -1547 -4006 -1491 -3935
rect -1387 -4006 -1331 -3935
rect -1227 -4006 -1171 -3935
rect -1067 -4006 -1011 -3935
rect -907 -4006 -851 -3935
rect -747 -4006 -691 -3935
rect 189 -3976 205 -3927
rect 252 -3976 291 -3927
rect 189 -3991 291 -3976
rect -1547 -4056 -690 -4006
rect 235 -4056 291 -3991
rect 395 -4056 451 -3895
rect 555 -4056 611 -3895
rect 715 -4056 771 -3895
rect 5685 -3735 5741 -3599
rect 5880 -3643 5955 -3631
rect 6088 -3643 6144 -3599
rect 6248 -3643 6304 -3599
rect 6408 -3643 6464 -3599
rect 6568 -3643 6624 -3599
rect 6728 -3643 6784 -3599
rect 6888 -3643 6944 -3599
rect 5880 -3644 6944 -3643
rect 5880 -3690 5895 -3644
rect 5941 -3690 6944 -3644
rect 5880 -3691 6944 -3690
rect 5880 -3705 5955 -3691
rect 6088 -3735 6144 -3691
rect 6248 -3735 6304 -3691
rect 6408 -3735 6464 -3691
rect 6568 -3735 6624 -3691
rect 6728 -3735 6784 -3691
rect 6888 -3735 6944 -3691
rect -2598 -4258 -2298 -4241
rect -4460 -4270 -4297 -4262
rect -4522 -4275 -4297 -4270
rect -4522 -4283 -4446 -4275
rect -4353 -4324 -4297 -4275
rect -3950 -4324 -3894 -4280
rect -3790 -4324 -3734 -4280
rect -3630 -4324 -3574 -4280
rect -3470 -4324 -3414 -4280
rect -3310 -4324 -3254 -4280
rect -3150 -4324 -3094 -4280
rect -2354 -4317 -2298 -4258
rect -2119 -4209 -1894 -4196
rect -2119 -4217 -1998 -4209
rect -2119 -4263 -2105 -4217
rect -2057 -4255 -1998 -4217
rect -1952 -4255 -1894 -4209
rect -2057 -4263 -1894 -4255
rect -2119 -4268 -1894 -4263
rect -2119 -4276 -2043 -4268
rect -1950 -4317 -1894 -4268
rect -1547 -4317 -1491 -4273
rect -1387 -4317 -1331 -4273
rect -1227 -4317 -1171 -4273
rect -1067 -4317 -1011 -4273
rect -907 -4317 -851 -4273
rect -747 -4317 -691 -4273
rect 235 -4292 291 -4156
rect 395 -4292 451 -4156
rect 555 -4292 611 -4156
rect 715 -4292 771 -4156
rect 2005 -4195 2061 -3934
rect 2408 -4005 2464 -3934
rect 2568 -4005 2624 -3934
rect 2728 -4005 2784 -3934
rect 2888 -4005 2944 -3934
rect 3048 -4005 3104 -3934
rect 3208 -4005 3264 -3934
rect 3818 -4005 3874 -3934
rect 3978 -4005 4034 -3934
rect 4138 -4005 4194 -3934
rect 4298 -4005 4354 -3934
rect 4458 -4005 4514 -3934
rect 4618 -4005 4674 -3934
rect 2408 -4055 3265 -4005
rect 3817 -4055 4674 -4005
rect 1836 -4208 2061 -4195
rect 1836 -4216 1957 -4208
rect 1836 -4262 1850 -4216
rect 1898 -4254 1957 -4216
rect 2003 -4254 2061 -4208
rect 1898 -4262 2061 -4254
rect 1836 -4267 2061 -4262
rect 1836 -4275 1912 -4267
rect 2005 -4316 2061 -4267
rect 5021 -4195 5077 -3934
rect 5021 -4208 5246 -4195
rect 5685 -4196 5741 -3935
rect 6088 -4006 6144 -3935
rect 6248 -4006 6304 -3935
rect 6408 -4006 6464 -3935
rect 6568 -4006 6624 -3935
rect 6728 -4006 6784 -3935
rect 6888 -4006 6944 -3935
rect 6088 -4056 6945 -4006
rect 5021 -4254 5079 -4208
rect 5125 -4216 5246 -4208
rect 5125 -4254 5184 -4216
rect 5021 -4262 5184 -4254
rect 5232 -4262 5246 -4216
rect 5021 -4267 5246 -4262
rect 2408 -4316 2464 -4272
rect 2568 -4316 2624 -4272
rect 2728 -4316 2784 -4272
rect 2888 -4316 2944 -4272
rect 3048 -4316 3104 -4272
rect 3208 -4316 3264 -4272
rect 3818 -4316 3874 -4272
rect 3978 -4316 4034 -4272
rect 4138 -4316 4194 -4272
rect 4298 -4316 4354 -4272
rect 4458 -4316 4514 -4272
rect 4618 -4316 4674 -4272
rect 5021 -4316 5077 -4267
rect 5170 -4275 5246 -4267
rect 5516 -4209 5741 -4196
rect 5516 -4217 5637 -4209
rect 5516 -4263 5530 -4217
rect 5578 -4255 5637 -4217
rect 5683 -4255 5741 -4209
rect 5578 -4263 5741 -4255
rect 5516 -4268 5741 -4263
rect 5516 -4276 5592 -4268
rect 235 -4436 291 -4392
rect 395 -4436 451 -4392
rect 555 -4436 611 -4392
rect 715 -4436 771 -4392
rect 5685 -4317 5741 -4268
rect 6088 -4317 6144 -4273
rect 6248 -4317 6304 -4273
rect 6408 -4317 6464 -4273
rect 6568 -4317 6624 -4273
rect 6728 -4317 6784 -4273
rect 6888 -4317 6944 -4273
rect -4757 -4660 -4701 -4524
rect -4353 -4564 -4297 -4524
rect -3950 -4564 -3894 -4524
rect -4353 -4568 -3894 -4564
rect -3790 -4568 -3734 -4524
rect -3630 -4568 -3574 -4524
rect -3470 -4568 -3414 -4524
rect -3310 -4568 -3254 -4524
rect -3150 -4568 -3094 -4524
rect -4353 -4616 -3094 -4568
rect -4353 -4620 -3894 -4616
rect -4353 -4660 -4297 -4620
rect -3950 -4660 -3894 -4620
rect -3790 -4660 -3734 -4616
rect -3630 -4660 -3574 -4616
rect -3470 -4660 -3414 -4616
rect -3310 -4660 -3254 -4616
rect -3150 -4660 -3094 -4616
rect -2354 -4653 -2298 -4517
rect -1950 -4557 -1894 -4517
rect -1547 -4557 -1491 -4517
rect -1950 -4561 -1491 -4557
rect -1387 -4561 -1331 -4517
rect -1227 -4561 -1171 -4517
rect -1067 -4561 -1011 -4517
rect -907 -4561 -851 -4517
rect -747 -4561 -691 -4517
rect -1950 -4609 -691 -4561
rect 2005 -4556 2061 -4516
rect 2408 -4556 2464 -4516
rect 2005 -4560 2464 -4556
rect 2568 -4560 2624 -4516
rect 2728 -4560 2784 -4516
rect 2888 -4560 2944 -4516
rect 3048 -4560 3104 -4516
rect 3208 -4560 3264 -4516
rect -1950 -4613 -1491 -4609
rect -1950 -4653 -1894 -4613
rect -1547 -4653 -1491 -4613
rect -1387 -4653 -1331 -4609
rect -1227 -4653 -1171 -4609
rect -1067 -4653 -1011 -4609
rect -907 -4653 -851 -4609
rect -747 -4653 -691 -4609
rect 2005 -4608 3264 -4560
rect 2005 -4612 2464 -4608
rect 2005 -4652 2061 -4612
rect 2408 -4652 2464 -4612
rect 2568 -4652 2624 -4608
rect 2728 -4652 2784 -4608
rect 2888 -4652 2944 -4608
rect 3048 -4652 3104 -4608
rect 3208 -4652 3264 -4608
rect 3818 -4560 3874 -4516
rect 3978 -4560 4034 -4516
rect 4138 -4560 4194 -4516
rect 4298 -4560 4354 -4516
rect 4458 -4560 4514 -4516
rect 4618 -4556 4674 -4516
rect 5021 -4556 5077 -4516
rect 4618 -4560 5077 -4556
rect 3818 -4608 5077 -4560
rect 3818 -4652 3874 -4608
rect 3978 -4652 4034 -4608
rect 4138 -4652 4194 -4608
rect 4298 -4652 4354 -4608
rect 4458 -4652 4514 -4608
rect 4618 -4612 5077 -4608
rect 4618 -4652 4674 -4612
rect 5021 -4652 5077 -4612
rect 5685 -4557 5741 -4517
rect 6088 -4557 6144 -4517
rect 5685 -4561 6144 -4557
rect 6248 -4561 6304 -4517
rect 6408 -4561 6464 -4517
rect 6568 -4561 6624 -4517
rect 6728 -4561 6784 -4517
rect 6888 -4561 6944 -4517
rect 5685 -4609 6944 -4561
rect 5685 -4613 6144 -4609
rect 5685 -4653 5741 -4613
rect 6088 -4653 6144 -4613
rect 6248 -4653 6304 -4609
rect 6408 -4653 6464 -4609
rect 6568 -4653 6624 -4609
rect 6728 -4653 6784 -4609
rect 6888 -4653 6944 -4609
rect -4757 -4904 -4701 -4860
rect -4353 -4880 -4297 -4860
rect -3950 -4880 -3894 -4860
rect -3790 -4880 -3734 -4860
rect -3630 -4880 -3574 -4860
rect -3470 -4880 -3414 -4860
rect -3310 -4880 -3254 -4860
rect -3150 -4880 -3094 -4860
rect -4353 -4904 -3094 -4880
rect -2354 -4897 -2298 -4853
rect -1950 -4873 -1894 -4853
rect -1547 -4873 -1491 -4853
rect -1387 -4873 -1331 -4853
rect -1227 -4873 -1171 -4853
rect -1067 -4873 -1011 -4853
rect -907 -4873 -851 -4853
rect -747 -4873 -691 -4853
rect -1950 -4897 -691 -4873
rect 2005 -4872 2061 -4852
rect 2408 -4872 2464 -4852
rect 2568 -4872 2624 -4852
rect 2728 -4872 2784 -4852
rect 2888 -4872 2944 -4852
rect 3048 -4872 3104 -4852
rect 3208 -4872 3264 -4852
rect 2005 -4896 3264 -4872
rect 3818 -4872 3874 -4852
rect 3978 -4872 4034 -4852
rect 4138 -4872 4194 -4852
rect 4298 -4872 4354 -4852
rect 4458 -4872 4514 -4852
rect 4618 -4872 4674 -4852
rect 5021 -4872 5077 -4852
rect 3818 -4896 5077 -4872
rect -4353 -4936 -3095 -4904
rect -1950 -4929 -692 -4897
rect 2005 -4928 3263 -4896
rect 3819 -4928 5077 -4896
rect 5685 -4873 5741 -4853
rect 6088 -4873 6144 -4853
rect 6248 -4873 6304 -4853
rect 6408 -4873 6464 -4853
rect 6568 -4873 6624 -4853
rect 6728 -4873 6784 -4853
rect 6888 -4873 6944 -4853
rect 5685 -4897 6944 -4873
rect 5685 -4929 6943 -4897
rect -4353 -5268 -3095 -5236
rect -1950 -5261 -692 -5229
rect 245 -5260 1503 -5228
rect 2006 -5260 3264 -5228
rect -4757 -5312 -4701 -5268
rect -4353 -5292 -3094 -5268
rect -4353 -5312 -4297 -5292
rect -3950 -5312 -3894 -5292
rect -3790 -5312 -3734 -5292
rect -3630 -5312 -3574 -5292
rect -3470 -5312 -3414 -5292
rect -3310 -5312 -3254 -5292
rect -3150 -5312 -3094 -5292
rect -2354 -5305 -2298 -5261
rect -1950 -5285 -691 -5261
rect -1950 -5305 -1894 -5285
rect -1547 -5305 -1491 -5285
rect -1387 -5305 -1331 -5285
rect -1227 -5305 -1171 -5285
rect -1067 -5305 -1011 -5285
rect -907 -5305 -851 -5285
rect -747 -5305 -691 -5285
rect 245 -5284 1504 -5260
rect 245 -5304 301 -5284
rect 648 -5304 704 -5284
rect 808 -5304 864 -5284
rect 968 -5304 1024 -5284
rect 1128 -5304 1184 -5284
rect 1288 -5304 1344 -5284
rect 1448 -5304 1504 -5284
rect 2005 -5284 3264 -5260
rect 2005 -5304 2061 -5284
rect 2165 -5304 2221 -5284
rect 2325 -5304 2381 -5284
rect 2485 -5304 2541 -5284
rect 2645 -5304 2701 -5284
rect 2805 -5304 2861 -5284
rect 3208 -5304 3264 -5284
rect 3818 -5260 5076 -5228
rect 3818 -5284 5077 -5260
rect 5686 -5261 6944 -5229
rect 3818 -5304 3874 -5284
rect 4221 -5304 4277 -5284
rect 4381 -5304 4437 -5284
rect 4541 -5304 4597 -5284
rect 4701 -5304 4757 -5284
rect 4861 -5304 4917 -5284
rect 5021 -5304 5077 -5284
rect 5685 -5285 6944 -5261
rect 5685 -5305 5741 -5285
rect 5845 -5305 5901 -5285
rect 6005 -5305 6061 -5285
rect 6165 -5305 6221 -5285
rect 6325 -5305 6381 -5285
rect 6485 -5305 6541 -5285
rect 6888 -5305 6944 -5285
rect -4757 -5648 -4701 -5512
rect -4353 -5552 -4297 -5512
rect -3950 -5552 -3894 -5512
rect -4353 -5556 -3894 -5552
rect -3790 -5556 -3734 -5512
rect -3630 -5556 -3574 -5512
rect -3470 -5556 -3414 -5512
rect -3310 -5556 -3254 -5512
rect -3150 -5556 -3094 -5512
rect -4353 -5604 -3094 -5556
rect -4353 -5608 -3894 -5604
rect -4353 -5648 -4297 -5608
rect -3950 -5648 -3894 -5608
rect -3790 -5648 -3734 -5604
rect -3630 -5648 -3574 -5604
rect -3470 -5648 -3414 -5604
rect -3310 -5648 -3254 -5604
rect -3150 -5648 -3094 -5604
rect -2354 -5641 -2298 -5505
rect -1950 -5545 -1894 -5505
rect -1547 -5545 -1491 -5505
rect -1950 -5549 -1491 -5545
rect -1387 -5549 -1331 -5505
rect -1227 -5549 -1171 -5505
rect -1067 -5549 -1011 -5505
rect -907 -5549 -851 -5505
rect -747 -5549 -691 -5505
rect -1950 -5597 -691 -5549
rect -1950 -5601 -1491 -5597
rect -1950 -5641 -1894 -5601
rect -1547 -5641 -1491 -5601
rect -1387 -5641 -1331 -5597
rect -1227 -5641 -1171 -5597
rect -1067 -5641 -1011 -5597
rect -907 -5641 -851 -5597
rect -747 -5641 -691 -5597
rect 245 -5544 301 -5504
rect 648 -5544 704 -5504
rect 245 -5548 704 -5544
rect 808 -5548 864 -5504
rect 968 -5548 1024 -5504
rect 1128 -5548 1184 -5504
rect 1288 -5548 1344 -5504
rect 1448 -5548 1504 -5504
rect 245 -5596 1504 -5548
rect 245 -5600 704 -5596
rect 245 -5640 301 -5600
rect 648 -5640 704 -5600
rect 808 -5640 864 -5596
rect 968 -5640 1024 -5596
rect 1128 -5640 1184 -5596
rect 1288 -5640 1344 -5596
rect 1448 -5640 1504 -5596
rect 2005 -5548 2061 -5504
rect 2165 -5548 2221 -5504
rect 2325 -5548 2381 -5504
rect 2485 -5548 2541 -5504
rect 2645 -5548 2701 -5504
rect 2805 -5544 2861 -5504
rect 3208 -5544 3264 -5504
rect 2805 -5548 3264 -5544
rect 2005 -5596 3264 -5548
rect 2005 -5640 2061 -5596
rect 2165 -5640 2221 -5596
rect 2325 -5640 2381 -5596
rect 2485 -5640 2541 -5596
rect 2645 -5640 2701 -5596
rect 2805 -5600 3264 -5596
rect 2805 -5640 2861 -5600
rect 3208 -5640 3264 -5600
rect 3818 -5544 3874 -5504
rect 4221 -5544 4277 -5504
rect 3818 -5548 4277 -5544
rect 4381 -5548 4437 -5504
rect 4541 -5548 4597 -5504
rect 4701 -5548 4757 -5504
rect 4861 -5548 4917 -5504
rect 5021 -5548 5077 -5504
rect 3818 -5596 5077 -5548
rect 3818 -5600 4277 -5596
rect 3818 -5640 3874 -5600
rect 4221 -5640 4277 -5600
rect 4381 -5640 4437 -5596
rect 4541 -5640 4597 -5596
rect 4701 -5640 4757 -5596
rect 4861 -5640 4917 -5596
rect 5021 -5640 5077 -5596
rect 5685 -5549 5741 -5505
rect 5845 -5549 5901 -5505
rect 6005 -5549 6061 -5505
rect 6165 -5549 6221 -5505
rect 6325 -5549 6381 -5505
rect 6485 -5545 6541 -5505
rect 6888 -5545 6944 -5505
rect 6485 -5549 6944 -5545
rect 5685 -5597 6944 -5549
rect 5685 -5641 5741 -5597
rect 5845 -5641 5901 -5597
rect 6005 -5641 6061 -5597
rect 6165 -5641 6221 -5597
rect 6325 -5641 6381 -5597
rect 6485 -5601 6944 -5597
rect 6485 -5641 6541 -5601
rect 6888 -5641 6944 -5601
rect -4757 -5907 -4701 -5848
rect -5001 -5924 -4701 -5907
rect -5001 -5970 -4980 -5924
rect -4934 -5970 -4882 -5924
rect -4836 -5970 -4784 -5924
rect -4738 -5970 -4701 -5924
rect -4522 -5897 -4446 -5889
rect -4353 -5897 -4297 -5848
rect -3950 -5892 -3894 -5848
rect -3790 -5892 -3734 -5848
rect -3630 -5892 -3574 -5848
rect -3470 -5892 -3414 -5848
rect -3310 -5892 -3254 -5848
rect -3150 -5892 -3094 -5848
rect -4522 -5902 -4297 -5897
rect -2354 -5900 -2298 -5841
rect -4522 -5948 -4508 -5902
rect -4460 -5910 -4297 -5902
rect -4460 -5948 -4401 -5910
rect -4522 -5956 -4401 -5948
rect -4355 -5956 -4297 -5910
rect -4522 -5969 -4297 -5956
rect -5001 -5987 -4701 -5970
rect -4757 -6230 -4701 -5987
rect -4353 -6230 -4297 -5969
rect -2598 -5917 -2298 -5900
rect -2598 -5963 -2577 -5917
rect -2531 -5963 -2479 -5917
rect -2433 -5963 -2381 -5917
rect -2335 -5963 -2298 -5917
rect -2119 -5890 -2043 -5882
rect -1950 -5890 -1894 -5841
rect -1547 -5885 -1491 -5841
rect -1387 -5885 -1331 -5841
rect -1227 -5885 -1171 -5841
rect -1067 -5885 -1011 -5841
rect -907 -5885 -851 -5841
rect -747 -5885 -691 -5841
rect -2119 -5895 -1894 -5890
rect -2119 -5941 -2105 -5895
rect -2057 -5903 -1894 -5895
rect -2057 -5941 -1998 -5903
rect -2119 -5949 -1998 -5941
rect -1952 -5949 -1894 -5903
rect -2119 -5962 -1894 -5949
rect 76 -5889 152 -5881
rect 245 -5889 301 -5840
rect 648 -5884 704 -5840
rect 808 -5884 864 -5840
rect 968 -5884 1024 -5840
rect 1128 -5884 1184 -5840
rect 1288 -5884 1344 -5840
rect 1448 -5884 1504 -5840
rect 2005 -5884 2061 -5840
rect 2165 -5884 2221 -5840
rect 2325 -5884 2381 -5840
rect 2485 -5884 2541 -5840
rect 2645 -5884 2701 -5840
rect 2805 -5884 2861 -5840
rect 76 -5894 301 -5889
rect 76 -5940 90 -5894
rect 138 -5902 301 -5894
rect 138 -5940 197 -5902
rect 76 -5948 197 -5940
rect 243 -5948 301 -5902
rect 76 -5961 301 -5948
rect -2598 -5980 -2298 -5963
rect -3950 -6159 -3093 -6109
rect -3950 -6230 -3894 -6159
rect -3790 -6230 -3734 -6159
rect -3630 -6230 -3574 -6159
rect -3470 -6230 -3414 -6159
rect -3310 -6230 -3254 -6159
rect -3150 -6230 -3094 -6159
rect -2354 -6223 -2298 -5980
rect -1950 -6223 -1894 -5962
rect -1547 -6152 -690 -6102
rect -1547 -6223 -1491 -6152
rect -1387 -6223 -1331 -6152
rect -1227 -6223 -1171 -6152
rect -1067 -6223 -1011 -6152
rect -907 -6223 -851 -6152
rect -747 -6223 -691 -6152
rect 245 -6222 301 -5961
rect 3208 -5889 3264 -5840
rect 3357 -5889 3433 -5881
rect 3208 -5894 3433 -5889
rect 3208 -5902 3371 -5894
rect 3208 -5948 3266 -5902
rect 3312 -5940 3371 -5902
rect 3419 -5940 3433 -5894
rect 3312 -5948 3433 -5940
rect 3208 -5961 3433 -5948
rect 3649 -5889 3725 -5881
rect 3818 -5889 3874 -5840
rect 4221 -5884 4277 -5840
rect 4381 -5884 4437 -5840
rect 4541 -5884 4597 -5840
rect 4701 -5884 4757 -5840
rect 4861 -5884 4917 -5840
rect 5021 -5884 5077 -5840
rect 5685 -5885 5741 -5841
rect 5845 -5885 5901 -5841
rect 6005 -5885 6061 -5841
rect 6165 -5885 6221 -5841
rect 6325 -5885 6381 -5841
rect 6485 -5885 6541 -5841
rect 3649 -5894 3874 -5889
rect 3649 -5940 3663 -5894
rect 3711 -5902 3874 -5894
rect 3711 -5940 3770 -5902
rect 3649 -5948 3770 -5940
rect 3816 -5948 3874 -5902
rect 3649 -5961 3874 -5948
rect 648 -6151 1505 -6101
rect 2004 -6151 2861 -6101
rect 648 -6222 704 -6151
rect 808 -6222 864 -6151
rect 968 -6222 1024 -6151
rect 1128 -6222 1184 -6151
rect 1288 -6222 1344 -6151
rect 1448 -6222 1504 -6151
rect 2005 -6222 2061 -6151
rect 2165 -6222 2221 -6151
rect 2325 -6222 2381 -6151
rect 2485 -6222 2541 -6151
rect 2645 -6222 2701 -6151
rect 2805 -6222 2861 -6151
rect 3208 -6222 3264 -5961
rect 3818 -6222 3874 -5961
rect 6888 -5890 6944 -5841
rect 7037 -5890 7113 -5882
rect 6888 -5895 7113 -5890
rect 6888 -5903 7051 -5895
rect 6888 -5949 6946 -5903
rect 6992 -5941 7051 -5903
rect 7099 -5941 7113 -5895
rect 6992 -5949 7113 -5941
rect 6888 -5962 7113 -5949
rect 4221 -6151 5078 -6101
rect 4221 -6222 4277 -6151
rect 4381 -6222 4437 -6151
rect 4541 -6222 4597 -6151
rect 4701 -6222 4757 -6151
rect 4861 -6222 4917 -6151
rect 5021 -6222 5077 -6151
rect 5684 -6152 6541 -6102
rect 5685 -6223 5741 -6152
rect 5845 -6223 5901 -6152
rect 6005 -6223 6061 -6152
rect 6165 -6223 6221 -6152
rect 6325 -6223 6381 -6152
rect 6485 -6223 6541 -6152
rect 6888 -6223 6944 -5962
rect -4757 -6566 -4701 -6430
rect -4353 -6566 -4297 -6430
rect -4158 -6474 -4083 -6460
rect -3950 -6474 -3894 -6430
rect -3790 -6474 -3734 -6430
rect -3630 -6474 -3574 -6430
rect -3470 -6474 -3414 -6430
rect -3310 -6474 -3254 -6430
rect -3150 -6474 -3094 -6430
rect -4158 -6475 -3094 -6474
rect -4158 -6521 -4143 -6475
rect -4097 -6521 -3094 -6475
rect -4158 -6522 -3094 -6521
rect -4158 -6534 -4083 -6522
rect -3950 -6566 -3894 -6522
rect -3790 -6566 -3734 -6522
rect -3630 -6566 -3574 -6522
rect -3470 -6566 -3414 -6522
rect -3310 -6566 -3254 -6522
rect -3150 -6566 -3094 -6522
rect -2354 -6559 -2298 -6423
rect -1950 -6559 -1894 -6423
rect -1755 -6467 -1680 -6453
rect -1547 -6467 -1491 -6423
rect -1387 -6467 -1331 -6423
rect -1227 -6467 -1171 -6423
rect -1067 -6467 -1011 -6423
rect -907 -6467 -851 -6423
rect -747 -6467 -691 -6423
rect -1755 -6468 -691 -6467
rect -1755 -6514 -1740 -6468
rect -1694 -6514 -691 -6468
rect -1755 -6515 -691 -6514
rect -1755 -6527 -1680 -6515
rect -1547 -6559 -1491 -6515
rect -1387 -6559 -1331 -6515
rect -1227 -6559 -1171 -6515
rect -1067 -6559 -1011 -6515
rect -907 -6559 -851 -6515
rect -747 -6559 -691 -6515
rect 245 -6558 301 -6422
rect 440 -6466 515 -6452
rect 648 -6466 704 -6422
rect 808 -6466 864 -6422
rect 968 -6466 1024 -6422
rect 1128 -6466 1184 -6422
rect 1288 -6466 1344 -6422
rect 1448 -6466 1504 -6422
rect 440 -6467 1504 -6466
rect 440 -6513 455 -6467
rect 501 -6513 1504 -6467
rect 440 -6514 1504 -6513
rect 440 -6526 515 -6514
rect 648 -6558 704 -6514
rect 808 -6558 864 -6514
rect 968 -6558 1024 -6514
rect 1128 -6558 1184 -6514
rect 1288 -6558 1344 -6514
rect 1448 -6558 1504 -6514
rect 2005 -6466 2061 -6422
rect 2165 -6466 2221 -6422
rect 2325 -6466 2381 -6422
rect 2485 -6466 2541 -6422
rect 2645 -6466 2701 -6422
rect 2805 -6466 2861 -6422
rect 2994 -6466 3069 -6452
rect 2005 -6467 3069 -6466
rect 2005 -6513 3008 -6467
rect 3054 -6513 3069 -6467
rect 2005 -6514 3069 -6513
rect 2005 -6558 2061 -6514
rect 2165 -6558 2221 -6514
rect 2325 -6558 2381 -6514
rect 2485 -6558 2541 -6514
rect 2645 -6558 2701 -6514
rect 2805 -6558 2861 -6514
rect 2994 -6526 3069 -6514
rect 3208 -6558 3264 -6422
rect 3818 -6558 3874 -6422
rect 4013 -6466 4088 -6452
rect 4221 -6466 4277 -6422
rect 4381 -6466 4437 -6422
rect 4541 -6466 4597 -6422
rect 4701 -6466 4757 -6422
rect 4861 -6466 4917 -6422
rect 5021 -6466 5077 -6422
rect 4013 -6467 5077 -6466
rect 4013 -6513 4028 -6467
rect 4074 -6513 5077 -6467
rect 4013 -6514 5077 -6513
rect 4013 -6526 4088 -6514
rect 4221 -6558 4277 -6514
rect 4381 -6558 4437 -6514
rect 4541 -6558 4597 -6514
rect 4701 -6558 4757 -6514
rect 4861 -6558 4917 -6514
rect 5021 -6558 5077 -6514
rect 5685 -6467 5741 -6423
rect 5845 -6467 5901 -6423
rect 6005 -6467 6061 -6423
rect 6165 -6467 6221 -6423
rect 6325 -6467 6381 -6423
rect 6485 -6467 6541 -6423
rect 6674 -6467 6749 -6453
rect 5685 -6468 6749 -6467
rect 5685 -6514 6688 -6468
rect 6734 -6514 6749 -6468
rect 5685 -6515 6749 -6514
rect 5685 -6559 5741 -6515
rect 5845 -6559 5901 -6515
rect 6005 -6559 6061 -6515
rect 6165 -6559 6221 -6515
rect 6325 -6559 6381 -6515
rect 6485 -6559 6541 -6515
rect 6674 -6527 6749 -6515
rect 6888 -6559 6944 -6423
rect -4757 -6902 -4701 -6766
rect -4353 -6902 -4297 -6766
rect -4158 -6810 -4083 -6796
rect -3950 -6810 -3894 -6766
rect -3790 -6810 -3734 -6766
rect -3630 -6810 -3574 -6766
rect -3470 -6810 -3414 -6766
rect -3310 -6810 -3254 -6766
rect -3150 -6810 -3094 -6766
rect -4158 -6811 -3094 -6810
rect -4158 -6857 -4143 -6811
rect -4097 -6857 -3094 -6811
rect -4158 -6858 -3094 -6857
rect -4158 -6870 -4083 -6858
rect -3950 -6902 -3894 -6858
rect -3790 -6902 -3734 -6858
rect -3630 -6902 -3574 -6858
rect -3470 -6902 -3414 -6858
rect -3310 -6902 -3254 -6858
rect -3150 -6902 -3094 -6858
rect -2354 -6895 -2298 -6759
rect -1950 -6895 -1894 -6759
rect -1755 -6803 -1680 -6789
rect -1547 -6803 -1491 -6759
rect -1387 -6803 -1331 -6759
rect -1227 -6803 -1171 -6759
rect -1067 -6803 -1011 -6759
rect -907 -6803 -851 -6759
rect -747 -6803 -691 -6759
rect -1755 -6804 -691 -6803
rect -1755 -6850 -1740 -6804
rect -1694 -6850 -691 -6804
rect -1755 -6851 -691 -6850
rect -1755 -6863 -1680 -6851
rect -1547 -6895 -1491 -6851
rect -1387 -6895 -1331 -6851
rect -1227 -6895 -1171 -6851
rect -1067 -6895 -1011 -6851
rect -907 -6895 -851 -6851
rect -747 -6895 -691 -6851
rect 245 -6894 301 -6758
rect 440 -6802 515 -6788
rect 648 -6802 704 -6758
rect 808 -6802 864 -6758
rect 968 -6802 1024 -6758
rect 1128 -6802 1184 -6758
rect 1288 -6802 1344 -6758
rect 1448 -6802 1504 -6758
rect 440 -6803 1504 -6802
rect 440 -6849 455 -6803
rect 501 -6849 1504 -6803
rect 440 -6850 1504 -6849
rect 440 -6862 515 -6850
rect 648 -6894 704 -6850
rect 808 -6894 864 -6850
rect 968 -6894 1024 -6850
rect 1128 -6894 1184 -6850
rect 1288 -6894 1344 -6850
rect 1448 -6894 1504 -6850
rect 2005 -6802 2061 -6758
rect 2165 -6802 2221 -6758
rect 2325 -6802 2381 -6758
rect 2485 -6802 2541 -6758
rect 2645 -6802 2701 -6758
rect 2805 -6802 2861 -6758
rect 2994 -6802 3069 -6788
rect 2005 -6803 3069 -6802
rect 2005 -6849 3008 -6803
rect 3054 -6849 3069 -6803
rect 2005 -6850 3069 -6849
rect 2005 -6894 2061 -6850
rect 2165 -6894 2221 -6850
rect 2325 -6894 2381 -6850
rect 2485 -6894 2541 -6850
rect 2645 -6894 2701 -6850
rect 2805 -6894 2861 -6850
rect 2994 -6862 3069 -6850
rect 3208 -6894 3264 -6758
rect 3818 -6894 3874 -6758
rect 4013 -6802 4088 -6788
rect 4221 -6802 4277 -6758
rect 4381 -6802 4437 -6758
rect 4541 -6802 4597 -6758
rect 4701 -6802 4757 -6758
rect 4861 -6802 4917 -6758
rect 5021 -6802 5077 -6758
rect 4013 -6803 5077 -6802
rect 4013 -6849 4028 -6803
rect 4074 -6849 5077 -6803
rect 4013 -6850 5077 -6849
rect 4013 -6862 4088 -6850
rect 4221 -6894 4277 -6850
rect 4381 -6894 4437 -6850
rect 4541 -6894 4597 -6850
rect 4701 -6894 4757 -6850
rect 4861 -6894 4917 -6850
rect 5021 -6894 5077 -6850
rect 5685 -6803 5741 -6759
rect 5845 -6803 5901 -6759
rect 6005 -6803 6061 -6759
rect 6165 -6803 6221 -6759
rect 6325 -6803 6381 -6759
rect 6485 -6803 6541 -6759
rect 6674 -6803 6749 -6789
rect 5685 -6804 6749 -6803
rect 5685 -6850 6688 -6804
rect 6734 -6850 6749 -6804
rect 5685 -6851 6749 -6850
rect 5685 -6895 5741 -6851
rect 5845 -6895 5901 -6851
rect 6005 -6895 6061 -6851
rect 6165 -6895 6221 -6851
rect 6325 -6895 6381 -6851
rect 6485 -6895 6541 -6851
rect 6674 -6863 6749 -6851
rect 6888 -6895 6944 -6759
rect -4757 -7238 -4701 -7102
rect -4353 -7238 -4297 -7102
rect -4158 -7146 -4083 -7132
rect -3950 -7146 -3894 -7102
rect -3790 -7146 -3734 -7102
rect -3630 -7146 -3574 -7102
rect -3470 -7146 -3414 -7102
rect -3310 -7146 -3254 -7102
rect -3150 -7146 -3094 -7102
rect -4158 -7147 -3094 -7146
rect -4158 -7193 -4143 -7147
rect -4097 -7193 -3094 -7147
rect -4158 -7194 -3094 -7193
rect -4158 -7206 -4083 -7194
rect -3950 -7238 -3894 -7194
rect -3790 -7238 -3734 -7194
rect -3630 -7238 -3574 -7194
rect -3470 -7238 -3414 -7194
rect -3310 -7238 -3254 -7194
rect -3150 -7238 -3094 -7194
rect -2354 -7231 -2298 -7095
rect -1950 -7231 -1894 -7095
rect -1755 -7139 -1680 -7125
rect -1547 -7139 -1491 -7095
rect -1387 -7139 -1331 -7095
rect -1227 -7139 -1171 -7095
rect -1067 -7139 -1011 -7095
rect -907 -7139 -851 -7095
rect -747 -7139 -691 -7095
rect -1755 -7140 -691 -7139
rect -1755 -7186 -1740 -7140
rect -1694 -7186 -691 -7140
rect -1755 -7187 -691 -7186
rect -1755 -7199 -1680 -7187
rect -1547 -7231 -1491 -7187
rect -1387 -7231 -1331 -7187
rect -1227 -7231 -1171 -7187
rect -1067 -7231 -1011 -7187
rect -907 -7231 -851 -7187
rect -747 -7231 -691 -7187
rect 245 -7230 301 -7094
rect 440 -7138 515 -7124
rect 648 -7138 704 -7094
rect 808 -7138 864 -7094
rect 968 -7138 1024 -7094
rect 1128 -7138 1184 -7094
rect 1288 -7138 1344 -7094
rect 1448 -7138 1504 -7094
rect 440 -7139 1504 -7138
rect 440 -7185 455 -7139
rect 501 -7185 1504 -7139
rect 440 -7186 1504 -7185
rect 440 -7198 515 -7186
rect 648 -7230 704 -7186
rect 808 -7230 864 -7186
rect 968 -7230 1024 -7186
rect 1128 -7230 1184 -7186
rect 1288 -7230 1344 -7186
rect 1448 -7230 1504 -7186
rect 2005 -7138 2061 -7094
rect 2165 -7138 2221 -7094
rect 2325 -7138 2381 -7094
rect 2485 -7138 2541 -7094
rect 2645 -7138 2701 -7094
rect 2805 -7138 2861 -7094
rect 2994 -7138 3069 -7124
rect 2005 -7139 3069 -7138
rect 2005 -7185 3008 -7139
rect 3054 -7185 3069 -7139
rect 2005 -7186 3069 -7185
rect 2005 -7230 2061 -7186
rect 2165 -7230 2221 -7186
rect 2325 -7230 2381 -7186
rect 2485 -7230 2541 -7186
rect 2645 -7230 2701 -7186
rect 2805 -7230 2861 -7186
rect 2994 -7198 3069 -7186
rect 3208 -7230 3264 -7094
rect 3818 -7230 3874 -7094
rect 4013 -7138 4088 -7124
rect 4221 -7138 4277 -7094
rect 4381 -7138 4437 -7094
rect 4541 -7138 4597 -7094
rect 4701 -7138 4757 -7094
rect 4861 -7138 4917 -7094
rect 5021 -7138 5077 -7094
rect 4013 -7139 5077 -7138
rect 4013 -7185 4028 -7139
rect 4074 -7185 5077 -7139
rect 4013 -7186 5077 -7185
rect 4013 -7198 4088 -7186
rect 4221 -7230 4277 -7186
rect 4381 -7230 4437 -7186
rect 4541 -7230 4597 -7186
rect 4701 -7230 4757 -7186
rect 4861 -7230 4917 -7186
rect 5021 -7230 5077 -7186
rect 5685 -7139 5741 -7095
rect 5845 -7139 5901 -7095
rect 6005 -7139 6061 -7095
rect 6165 -7139 6221 -7095
rect 6325 -7139 6381 -7095
rect 6485 -7139 6541 -7095
rect 6674 -7139 6749 -7125
rect 5685 -7140 6749 -7139
rect 5685 -7186 6688 -7140
rect 6734 -7186 6749 -7140
rect 5685 -7187 6749 -7186
rect 5685 -7231 5741 -7187
rect 5845 -7231 5901 -7187
rect 6005 -7231 6061 -7187
rect 6165 -7231 6221 -7187
rect 6325 -7231 6381 -7187
rect 6485 -7231 6541 -7187
rect 6674 -7199 6749 -7187
rect 6888 -7231 6944 -7095
rect -4757 -7482 -4701 -7438
rect -4353 -7482 -4297 -7438
rect -3950 -7482 -3894 -7438
rect -3790 -7482 -3734 -7438
rect -3630 -7482 -3574 -7438
rect -3470 -7482 -3414 -7438
rect -3310 -7482 -3254 -7438
rect -3150 -7482 -3094 -7438
rect -2354 -7475 -2298 -7431
rect -1950 -7475 -1894 -7431
rect -1547 -7475 -1491 -7431
rect -1387 -7475 -1331 -7431
rect -1227 -7475 -1171 -7431
rect -1067 -7475 -1011 -7431
rect -907 -7475 -851 -7431
rect -747 -7475 -691 -7431
rect 245 -7474 301 -7430
rect 648 -7474 704 -7430
rect 808 -7474 864 -7430
rect 968 -7474 1024 -7430
rect 1128 -7474 1184 -7430
rect 1288 -7474 1344 -7430
rect 1448 -7474 1504 -7430
rect 2005 -7474 2061 -7430
rect 2165 -7474 2221 -7430
rect 2325 -7474 2381 -7430
rect 2485 -7474 2541 -7430
rect 2645 -7474 2701 -7430
rect 2805 -7474 2861 -7430
rect 3208 -7474 3264 -7430
rect 3818 -7474 3874 -7430
rect 4221 -7474 4277 -7430
rect 4381 -7474 4437 -7430
rect 4541 -7474 4597 -7430
rect 4701 -7474 4757 -7430
rect 4861 -7474 4917 -7430
rect 5021 -7474 5077 -7430
rect 5685 -7475 5741 -7431
rect 5845 -7475 5901 -7431
rect 6005 -7475 6061 -7431
rect 6165 -7475 6221 -7431
rect 6325 -7475 6381 -7431
rect 6485 -7475 6541 -7431
rect 6888 -7475 6944 -7431
<< polycontact >>
rect -4143 2135 -4097 2181
rect -1740 2142 -1694 2188
rect 455 2143 501 2189
rect 3008 2143 3054 2189
rect 4028 2143 4074 2189
rect 6688 2142 6734 2188
rect -4143 1799 -4097 1845
rect -1740 1806 -1694 1852
rect 455 1807 501 1853
rect 3008 1807 3054 1853
rect 4028 1807 4074 1853
rect 6688 1806 6734 1852
rect -4143 1463 -4097 1509
rect -1740 1470 -1694 1516
rect 455 1471 501 1517
rect 3008 1471 3054 1517
rect 4028 1471 4074 1517
rect 6688 1470 6734 1516
rect -4980 912 -4934 958
rect -4882 912 -4836 958
rect -4784 912 -4738 958
rect -4508 890 -4460 936
rect -4401 898 -4355 944
rect -2577 919 -2531 965
rect -2479 919 -2433 965
rect -2381 919 -2335 965
rect -2105 897 -2057 943
rect -1998 905 -1952 951
rect 90 898 138 944
rect 197 906 243 952
rect 3266 906 3312 952
rect 3371 898 3419 944
rect 3663 898 3711 944
rect 3770 906 3816 952
rect 6946 905 6992 951
rect 7051 897 7099 943
rect -4980 -810 -4934 -764
rect -4882 -810 -4836 -764
rect -4784 -810 -4738 -764
rect -4508 -788 -4460 -742
rect -4401 -796 -4355 -750
rect -2577 -803 -2531 -757
rect -2479 -803 -2433 -757
rect -2381 -803 -2335 -757
rect -2105 -781 -2057 -735
rect -1998 -789 -1952 -743
rect 1850 -780 1898 -734
rect 1957 -788 2003 -742
rect 205 -1035 252 -986
rect 5079 -788 5125 -742
rect 5184 -780 5232 -734
rect 5530 -781 5578 -735
rect 5637 -789 5683 -743
rect -4143 -1361 -4097 -1315
rect -1740 -1354 -1694 -1308
rect 2215 -1353 2261 -1307
rect 4821 -1353 4867 -1307
rect -4143 -1697 -4097 -1651
rect -1740 -1690 -1694 -1644
rect 5895 -1354 5941 -1308
rect 2215 -1689 2261 -1643
rect 4821 -1689 4867 -1643
rect -4143 -2033 -4097 -1987
rect -1740 -2026 -1694 -1980
rect 5895 -1690 5941 -1644
rect 2215 -2025 2261 -1979
rect 4821 -2025 4867 -1979
rect 205 -2221 252 -2172
rect 5895 -2026 5941 -1980
rect -4143 -3025 -4097 -2979
rect -1740 -3018 -1694 -2972
rect 2215 -3017 2261 -2971
rect 4821 -3017 4867 -2971
rect -4143 -3361 -4097 -3315
rect 5895 -3018 5941 -2972
rect -1740 -3354 -1694 -3308
rect 2215 -3353 2261 -3307
rect 4821 -3353 4867 -3307
rect -4143 -3697 -4097 -3651
rect 5895 -3354 5941 -3308
rect -1740 -3690 -1694 -3644
rect 2215 -3689 2261 -3643
rect 4821 -3689 4867 -3643
rect -4980 -4248 -4934 -4202
rect -4882 -4248 -4836 -4202
rect -4784 -4248 -4738 -4202
rect -4508 -4270 -4460 -4224
rect -4401 -4262 -4355 -4216
rect -2577 -4241 -2531 -4195
rect -2479 -4241 -2433 -4195
rect -2381 -4241 -2335 -4195
rect 205 -3976 252 -3927
rect 5895 -3690 5941 -3644
rect -2105 -4263 -2057 -4217
rect -1998 -4255 -1952 -4209
rect 1850 -4262 1898 -4216
rect 1957 -4254 2003 -4208
rect 5079 -4254 5125 -4208
rect 5184 -4262 5232 -4216
rect 5530 -4263 5578 -4217
rect 5637 -4255 5683 -4209
rect -4980 -5970 -4934 -5924
rect -4882 -5970 -4836 -5924
rect -4784 -5970 -4738 -5924
rect -4508 -5948 -4460 -5902
rect -4401 -5956 -4355 -5910
rect -2577 -5963 -2531 -5917
rect -2479 -5963 -2433 -5917
rect -2381 -5963 -2335 -5917
rect -2105 -5941 -2057 -5895
rect -1998 -5949 -1952 -5903
rect 90 -5940 138 -5894
rect 197 -5948 243 -5902
rect 3266 -5948 3312 -5902
rect 3371 -5940 3419 -5894
rect 3663 -5940 3711 -5894
rect 3770 -5948 3816 -5902
rect 6946 -5949 6992 -5903
rect 7051 -5941 7099 -5895
rect -4143 -6521 -4097 -6475
rect -1740 -6514 -1694 -6468
rect 455 -6513 501 -6467
rect 3008 -6513 3054 -6467
rect 4028 -6513 4074 -6467
rect 6688 -6514 6734 -6468
rect -4143 -6857 -4097 -6811
rect -1740 -6850 -1694 -6804
rect 455 -6849 501 -6803
rect 3008 -6849 3054 -6803
rect 4028 -6849 4074 -6803
rect 6688 -6850 6734 -6804
rect -4143 -7193 -4097 -7147
rect -1740 -7186 -1694 -7140
rect 455 -7185 501 -7139
rect 3008 -7185 3054 -7139
rect 4028 -7185 4074 -7139
rect 6688 -7186 6734 -7140
<< metal1 >>
rect 71 2748 5251 2749
rect -2528 2745 -517 2748
rect 71 2745 7118 2748
rect -4931 2740 -2920 2741
rect -2528 2740 7118 2745
rect -4931 2689 7118 2740
rect -4931 2688 131 2689
rect -4931 2681 -2285 2688
rect -4931 2627 -4688 2681
rect -4527 2627 -4467 2681
rect -4306 2627 -4246 2681
rect -4085 2627 -4025 2681
rect -3864 2627 -3804 2681
rect -3643 2627 -3583 2681
rect -3422 2627 -3362 2681
rect -3201 2627 -3141 2681
rect -2980 2634 -2285 2681
rect -2124 2634 -2064 2688
rect -1903 2634 -1843 2688
rect -1682 2634 -1622 2688
rect -1461 2634 -1401 2688
rect -1240 2634 -1180 2688
rect -1019 2634 -959 2688
rect -798 2634 -738 2688
rect -577 2635 131 2688
rect 292 2635 352 2689
rect 513 2635 573 2689
rect 734 2635 794 2689
rect 955 2635 1015 2689
rect 1176 2635 1236 2689
rect 1397 2635 1457 2689
rect 1618 2635 1891 2689
rect 2052 2635 2112 2689
rect 2273 2635 2333 2689
rect 2494 2635 2554 2689
rect 2715 2635 2775 2689
rect 2936 2635 2996 2689
rect 3157 2635 3217 2689
rect 3378 2635 3704 2689
rect 3865 2635 3925 2689
rect 4086 2635 4146 2689
rect 4307 2635 4367 2689
rect 4528 2635 4588 2689
rect 4749 2635 4809 2689
rect 4970 2635 5030 2689
rect 5191 2688 7118 2689
rect 5191 2635 5571 2688
rect -577 2634 5571 2635
rect 5732 2634 5792 2688
rect 5953 2634 6013 2688
rect 6174 2634 6234 2688
rect 6395 2634 6455 2688
rect 6616 2687 6676 2688
rect 6837 2687 6897 2688
rect 6616 2635 6627 2687
rect 6837 2635 6867 2687
rect 6616 2634 6676 2635
rect 6837 2634 6897 2635
rect 7058 2634 7118 2688
rect -2980 2627 7118 2634
rect -4931 2575 7118 2627
rect -4931 2574 216 2575
rect -4931 2568 -2171 2574
rect -4931 2567 -2920 2568
rect -4832 2413 -4786 2567
rect -4832 2077 -4786 2239
rect -4832 1741 -4786 1903
rect -4832 1405 -4786 1567
rect -4832 1220 -4786 1231
rect -4672 2413 -4626 2424
rect -4672 2077 -4626 2239
rect -4672 1741 -4626 1903
rect -4672 1405 -4626 1567
rect -5214 1204 -5093 1208
rect -5214 1174 -5197 1204
rect -5352 1147 -5197 1174
rect -5140 1147 -5093 1204
rect -5352 1117 -5093 1147
rect -5214 1094 -5093 1117
rect -5214 1037 -5197 1094
rect -5140 1037 -5093 1094
rect -5214 1026 -5093 1037
rect -5040 975 -4978 977
rect -5040 969 -4727 975
rect -5111 958 -4727 969
rect -5111 941 -4980 958
rect -5114 885 -5104 941
rect -5048 885 -4994 941
rect -4934 912 -4882 958
rect -4836 912 -4784 958
rect -4738 912 -4727 958
rect -4938 895 -4727 912
rect -4672 954 -4626 1231
rect -4428 2413 -4382 2567
rect -4025 2470 -3019 2518
rect -4428 2077 -4382 2239
rect -4428 1741 -4382 1903
rect -4428 1405 -4382 1567
rect -4428 1220 -4382 1231
rect -4268 2413 -4222 2424
rect -4268 2180 -4222 2239
rect -4025 2413 -3979 2470
rect -4158 2181 -4083 2194
rect -4158 2180 -4143 2181
rect -4268 2135 -4143 2180
rect -4097 2135 -4083 2181
rect -4268 2134 -4083 2135
rect -4268 2077 -4222 2134
rect -4158 2120 -4083 2134
rect -4268 1844 -4222 1903
rect -4025 2077 -3979 2239
rect -4158 1845 -4083 1858
rect -4158 1844 -4143 1845
rect -4268 1799 -4143 1844
rect -4097 1799 -4083 1845
rect -4268 1798 -4083 1799
rect -4268 1741 -4222 1798
rect -4158 1784 -4083 1798
rect -4268 1508 -4222 1567
rect -4025 1741 -3979 1903
rect -4158 1509 -4083 1522
rect -4158 1508 -4143 1509
rect -4268 1463 -4143 1508
rect -4097 1463 -4083 1509
rect -4268 1462 -4083 1463
rect -4268 1405 -4222 1462
rect -4158 1448 -4083 1462
rect -4522 954 -4328 957
rect -4672 944 -4328 954
rect -4672 936 -4401 944
rect -4938 885 -4887 895
rect -5111 853 -4887 885
rect -4672 891 -4508 936
rect -5197 711 -5101 714
rect -5197 661 -5170 711
rect -5368 654 -5170 661
rect -5113 654 -5101 711
rect -5368 604 -5101 654
rect -5197 601 -5101 604
rect -5197 544 -5170 601
rect -5113 544 -5101 601
rect -5197 540 -5101 544
rect -5040 -615 -4978 853
rect -4832 823 -4786 834
rect -4832 487 -4786 649
rect -4832 161 -4786 313
rect -4672 823 -4626 891
rect -4522 890 -4508 891
rect -4460 898 -4401 936
rect -4355 898 -4328 944
rect -4460 890 -4328 898
rect -4522 885 -4328 890
rect -4522 877 -4446 885
rect -4672 487 -4626 649
rect -4672 302 -4626 313
rect -4428 823 -4382 834
rect -4428 487 -4382 649
rect -4428 161 -4382 313
rect -4268 823 -4222 1231
rect -4025 1405 -3979 1567
rect -3865 2413 -3819 2424
rect -3865 2077 -3819 2239
rect -3865 1741 -3819 1903
rect -3865 1433 -3819 1567
rect -3866 1405 -3819 1433
rect -3866 1387 -3865 1405
rect -4159 1201 -4082 1213
rect -4159 1147 -4145 1201
rect -4091 1197 -4082 1201
rect -4025 1197 -3979 1231
rect -4091 1147 -3979 1197
rect -4159 1089 -3979 1147
rect -3865 1174 -3819 1231
rect -3705 2413 -3659 2470
rect -3705 2077 -3659 2239
rect -3705 1741 -3659 1903
rect -3705 1405 -3659 1567
rect -3545 2413 -3499 2424
rect -3545 2077 -3499 2239
rect -3545 1741 -3499 1903
rect -3545 1405 -3499 1567
rect -3705 1220 -3659 1231
rect -3546 1174 -3499 1231
rect -3385 2413 -3339 2470
rect -3385 2077 -3339 2239
rect -3385 1741 -3339 1903
rect -3385 1405 -3339 1567
rect -3225 2413 -3179 2424
rect -3225 2077 -3179 2239
rect -3225 1741 -3179 1903
rect -3225 1405 -3179 1567
rect -3385 1220 -3339 1231
rect -3226 1174 -3179 1231
rect -3065 2413 -3019 2470
rect -3065 2077 -3019 2239
rect -3065 1741 -3019 1903
rect -3065 1405 -3019 1567
rect -3065 1220 -3019 1231
rect -2429 2420 -2383 2568
rect -2429 2084 -2383 2246
rect -2429 1748 -2383 1910
rect -2429 1412 -2383 1574
rect -2429 1227 -2383 1238
rect -2269 2420 -2223 2431
rect -2269 2084 -2223 2246
rect -2269 1748 -2223 1910
rect -2269 1412 -2223 1574
rect -3865 1172 -3179 1174
rect -3865 1161 -2840 1172
rect -3865 1105 -3020 1161
rect -2964 1105 -2909 1161
rect -2853 1105 -2840 1161
rect -3865 1097 -2840 1105
rect -3865 1095 -3179 1097
rect -4159 1030 -4149 1089
rect -4090 1030 -3979 1089
rect -4159 1017 -3979 1030
rect -4268 487 -4222 649
rect -4268 302 -4222 313
rect -4025 823 -3979 1017
rect -3275 990 -3179 1095
rect -4025 487 -3979 649
rect -4025 255 -3979 313
rect -3865 881 -3179 990
rect -2600 974 -2324 982
rect -2689 965 -2324 974
rect -2689 930 -2577 965
rect -2531 930 -2479 965
rect -3865 823 -3819 881
rect -3865 487 -3819 649
rect -3865 302 -3819 313
rect -3705 823 -3659 834
rect -3705 487 -3659 649
rect -3705 255 -3659 313
rect -3545 823 -3499 881
rect -3545 487 -3499 649
rect -3545 302 -3499 313
rect -3385 823 -3339 834
rect -3385 487 -3339 649
rect -3385 255 -3339 313
rect -3225 823 -3179 881
rect -2691 874 -2681 930
rect -2625 919 -2577 930
rect -2515 919 -2479 930
rect -2433 919 -2381 965
rect -2335 919 -2324 965
rect -2625 874 -2571 919
rect -2515 902 -2324 919
rect -2269 961 -2223 1238
rect -2025 2420 -1979 2574
rect -611 2573 216 2574
rect -1622 2477 -616 2525
rect -2025 2084 -1979 2246
rect -2025 1748 -1979 1910
rect -2025 1412 -1979 1574
rect -2025 1227 -1979 1238
rect -1865 2420 -1819 2431
rect -1865 2187 -1819 2246
rect -1622 2420 -1576 2477
rect -1755 2188 -1680 2201
rect -1755 2187 -1740 2188
rect -1865 2142 -1740 2187
rect -1694 2142 -1680 2188
rect -1865 2141 -1680 2142
rect -1865 2084 -1819 2141
rect -1755 2127 -1680 2141
rect -1865 1851 -1819 1910
rect -1622 2084 -1576 2246
rect -1755 1852 -1680 1865
rect -1755 1851 -1740 1852
rect -1865 1806 -1740 1851
rect -1694 1806 -1680 1852
rect -1865 1805 -1680 1806
rect -1865 1748 -1819 1805
rect -1755 1791 -1680 1805
rect -1865 1515 -1819 1574
rect -1622 1748 -1576 1910
rect -1755 1516 -1680 1529
rect -1755 1515 -1740 1516
rect -1865 1470 -1740 1515
rect -1694 1470 -1680 1516
rect -1865 1469 -1680 1470
rect -1865 1412 -1819 1469
rect -1755 1455 -1680 1469
rect -2119 961 -1925 964
rect -2269 951 -1925 961
rect -2269 943 -1998 951
rect -2515 874 -2481 902
rect -3225 487 -3179 649
rect -3225 302 -3179 313
rect -3065 823 -3019 834
rect -2689 830 -2481 874
rect -2269 898 -2105 943
rect -2429 830 -2383 841
rect -3065 487 -3019 649
rect -3065 255 -3019 313
rect -4025 207 -3019 255
rect -2429 494 -2383 656
rect -2429 168 -2383 320
rect -2269 830 -2223 898
rect -2119 897 -2105 898
rect -2057 905 -1998 943
rect -1952 905 -1925 951
rect -2057 897 -1925 905
rect -2119 892 -1925 897
rect -2119 884 -2043 892
rect -2269 494 -2223 656
rect -2269 309 -2223 320
rect -2025 830 -1979 841
rect -2025 494 -1979 656
rect -2025 168 -1979 320
rect -1865 830 -1819 1238
rect -1622 1412 -1576 1574
rect -1462 2420 -1416 2431
rect -1462 2084 -1416 2246
rect -1462 1748 -1416 1910
rect -1462 1440 -1416 1574
rect -1463 1412 -1416 1440
rect -1463 1394 -1462 1412
rect -1756 1208 -1679 1220
rect -1756 1154 -1742 1208
rect -1688 1204 -1679 1208
rect -1622 1204 -1576 1238
rect -1688 1154 -1576 1204
rect -1756 1096 -1576 1154
rect -1462 1181 -1416 1238
rect -1302 2420 -1256 2477
rect -1302 2084 -1256 2246
rect -1302 1748 -1256 1910
rect -1302 1412 -1256 1574
rect -1142 2420 -1096 2431
rect -1142 2084 -1096 2246
rect -1142 1748 -1096 1910
rect -1142 1412 -1096 1574
rect -1302 1227 -1256 1238
rect -1143 1181 -1096 1238
rect -982 2420 -936 2477
rect -982 2084 -936 2246
rect -982 1748 -936 1910
rect -982 1412 -936 1574
rect -822 2420 -776 2431
rect -822 2084 -776 2246
rect -822 1748 -776 1910
rect -822 1412 -776 1574
rect -982 1227 -936 1238
rect -823 1181 -776 1238
rect -662 2420 -616 2477
rect -662 2084 -616 2246
rect -662 1748 -616 1910
rect -662 1412 -616 1574
rect -662 1227 -616 1238
rect 170 2421 216 2573
rect 573 2478 1579 2526
rect 170 2085 216 2247
rect 170 1749 216 1911
rect 170 1413 216 1575
rect 170 1228 216 1239
rect 330 2421 376 2432
rect 330 2188 376 2247
rect 573 2421 619 2478
rect 440 2189 515 2202
rect 440 2188 455 2189
rect 330 2143 455 2188
rect 501 2143 515 2189
rect 330 2142 515 2143
rect 330 2085 376 2142
rect 440 2128 515 2142
rect 330 1852 376 1911
rect 573 2085 619 2247
rect 440 1853 515 1866
rect 440 1852 455 1853
rect 330 1807 455 1852
rect 501 1807 515 1853
rect 330 1806 515 1807
rect 330 1749 376 1806
rect 440 1792 515 1806
rect 330 1516 376 1575
rect 573 1749 619 1911
rect 440 1517 515 1530
rect 440 1516 455 1517
rect 330 1471 455 1516
rect 501 1471 515 1517
rect 330 1470 515 1471
rect 330 1413 376 1470
rect 440 1456 515 1470
rect 47 1214 124 1223
rect 46 1210 125 1214
rect 46 1188 58 1210
rect -1462 1179 -776 1181
rect -1462 1170 -437 1179
rect -1462 1169 -505 1170
rect -1462 1113 -625 1169
rect -569 1114 -505 1169
rect -449 1114 -437 1170
rect -9 1154 58 1188
rect 114 1154 125 1210
rect -9 1134 125 1154
rect -569 1113 -437 1114
rect -1462 1104 -437 1113
rect -1462 1102 -776 1104
rect -1756 1037 -1746 1096
rect -1687 1037 -1576 1096
rect -1756 1024 -1576 1037
rect -1865 494 -1819 656
rect -1865 309 -1819 320
rect -1622 830 -1576 1024
rect -872 997 -776 1102
rect 46 1100 125 1134
rect 46 1044 58 1100
rect 114 1044 125 1100
rect 46 1028 125 1044
rect -1622 494 -1576 656
rect -1622 262 -1576 320
rect -1462 888 -776 997
rect 76 952 270 965
rect 76 945 197 952
rect -1462 830 -1416 888
rect -1462 494 -1416 656
rect -1462 309 -1416 320
rect -1302 830 -1256 841
rect -1302 494 -1256 656
rect -1302 262 -1256 320
rect -1142 830 -1096 888
rect -1142 494 -1096 656
rect -1142 309 -1096 320
rect -982 830 -936 841
rect -982 494 -936 656
rect -982 262 -936 320
rect -822 830 -776 888
rect -86 944 197 945
rect -86 898 90 944
rect 138 906 197 944
rect 243 906 270 952
rect 138 898 270 906
rect -86 896 270 898
rect -822 494 -776 656
rect -822 309 -776 320
rect -662 830 -616 841
rect -86 821 -40 896
rect 76 893 270 896
rect 76 885 152 893
rect 170 831 216 842
rect -102 805 -13 821
rect -102 748 -84 805
rect -27 748 -13 805
rect -102 732 -13 748
rect -662 494 -616 656
rect -662 262 -616 320
rect -1622 214 -616 262
rect -2528 162 -517 168
rect -2973 161 -517 162
rect -4931 109 -517 161
rect -4931 108 -1009 109
rect -953 108 -899 109
rect -843 108 -789 109
rect -733 108 -679 109
rect -623 108 -517 109
rect -4931 101 -2285 108
rect -4931 47 -4688 101
rect -4527 47 -4467 101
rect -4306 47 -4246 101
rect -4085 47 -4025 101
rect -3864 47 -3804 101
rect -3643 47 -3583 101
rect -3422 47 -3362 101
rect -3201 47 -3141 101
rect -2980 54 -2285 101
rect -2124 54 -2064 108
rect -1903 54 -1843 108
rect -1682 54 -1622 108
rect -1461 54 -1401 108
rect -1240 54 -1180 108
rect -1019 54 -1009 108
rect -798 54 -789 108
rect -577 54 -517 108
rect -2980 53 -1009 54
rect -953 53 -899 54
rect -843 53 -789 54
rect -733 53 -679 54
rect -623 53 -517 54
rect -2980 47 -517 53
rect -4931 -6 -517 47
rect -4931 -10 -2265 -6
rect -4931 -13 -2920 -10
rect -4832 -165 -4786 -13
rect -4832 -501 -4786 -339
rect -5041 -623 -4935 -615
rect -5041 -679 -5016 -623
rect -4960 -679 -4935 -623
rect -5041 -733 -4935 -679
rect -4832 -686 -4786 -675
rect -4672 -165 -4626 -154
rect -4672 -501 -4626 -339
rect -5041 -789 -5016 -733
rect -4960 -747 -4935 -733
rect -4672 -743 -4626 -675
rect -4428 -165 -4382 -13
rect -4025 -107 -3019 -59
rect -4428 -501 -4382 -339
rect -4428 -686 -4382 -675
rect -4268 -165 -4222 -154
rect -4268 -501 -4222 -339
rect -4522 -737 -4446 -729
rect -4522 -742 -4328 -737
rect -4522 -743 -4508 -742
rect -4960 -764 -4727 -747
rect -5041 -804 -4980 -789
rect -5040 -810 -4980 -804
rect -4934 -810 -4882 -764
rect -4836 -810 -4784 -764
rect -4738 -810 -4727 -764
rect -5040 -827 -4727 -810
rect -4672 -788 -4508 -743
rect -4460 -750 -4328 -742
rect -4460 -788 -4401 -750
rect -4672 -796 -4401 -788
rect -4355 -796 -4328 -750
rect -4672 -806 -4328 -796
rect -5194 -914 -5099 -878
rect -5194 -965 -5181 -914
rect -5324 -972 -5181 -965
rect -5123 -972 -5099 -914
rect -5324 -1024 -5099 -972
rect -5324 -1025 -5181 -1024
rect -5194 -1082 -5181 -1025
rect -5123 -1082 -5099 -1024
rect -5194 -1094 -5099 -1082
rect -5189 -1391 -5094 -1381
rect -5189 -1439 -5164 -1391
rect -5254 -1447 -5164 -1439
rect -5108 -1447 -5094 -1391
rect -5254 -1493 -5094 -1447
rect -5189 -1501 -5094 -1493
rect -5189 -1557 -5164 -1501
rect -5108 -1557 -5094 -1501
rect -5189 -1567 -5094 -1557
rect -5209 -3275 -5121 -3268
rect -5209 -3323 -5193 -3275
rect -5288 -3331 -5193 -3323
rect -5137 -3331 -5121 -3275
rect -5288 -3377 -5121 -3331
rect -5209 -3385 -5121 -3377
rect -5209 -3441 -5193 -3385
rect -5137 -3441 -5121 -3385
rect -5209 -3458 -5121 -3441
rect -5189 -3959 -5107 -3947
rect -5336 -3960 -5107 -3959
rect -5336 -4014 -5177 -3960
rect -5189 -4018 -5177 -4014
rect -5119 -4018 -5107 -3960
rect -5189 -4070 -5107 -4018
rect -5189 -4128 -5177 -4070
rect -5119 -4128 -5107 -4070
rect -5189 -4135 -5107 -4128
rect -5040 -4185 -4978 -827
rect -4832 -1083 -4786 -1072
rect -4832 -1419 -4786 -1257
rect -4832 -1755 -4786 -1593
rect -4832 -2091 -4786 -1929
rect -4832 -2419 -4786 -2265
rect -4672 -1083 -4626 -806
rect -4522 -809 -4328 -806
rect -4672 -1419 -4626 -1257
rect -4672 -1755 -4626 -1593
rect -4672 -2091 -4626 -1929
rect -4672 -2276 -4626 -2265
rect -4428 -1083 -4382 -1072
rect -4428 -1419 -4382 -1257
rect -4428 -1755 -4382 -1593
rect -4428 -2091 -4382 -1929
rect -4428 -2419 -4382 -2265
rect -4268 -1083 -4222 -675
rect -4025 -165 -3979 -107
rect -4025 -501 -3979 -339
rect -4025 -869 -3979 -675
rect -3865 -165 -3819 -154
rect -3865 -501 -3819 -339
rect -3865 -733 -3819 -675
rect -3705 -165 -3659 -107
rect -3705 -501 -3659 -339
rect -3705 -686 -3659 -675
rect -3545 -165 -3499 -154
rect -3545 -501 -3499 -339
rect -3545 -733 -3499 -675
rect -3385 -165 -3339 -107
rect -3385 -501 -3339 -339
rect -3385 -686 -3339 -675
rect -3225 -165 -3179 -154
rect -3225 -501 -3179 -339
rect -3225 -733 -3179 -675
rect -3065 -165 -3019 -107
rect -3065 -501 -3019 -339
rect -2429 -158 -2383 -10
rect -2429 -494 -2383 -332
rect -3065 -686 -3019 -675
rect -2601 -624 -2501 -611
rect -2601 -680 -2582 -624
rect -2526 -680 -2501 -624
rect -2429 -679 -2383 -668
rect -2269 -158 -2223 -147
rect -2269 -494 -2223 -332
rect -3865 -842 -3179 -733
rect -2601 -734 -2501 -680
rect -2601 -790 -2582 -734
rect -2526 -740 -2501 -734
rect -2269 -736 -2223 -668
rect -2025 -158 -1979 -6
rect -1622 -100 -616 -52
rect -2025 -494 -1979 -332
rect -2025 -679 -1979 -668
rect -1865 -158 -1819 -147
rect -1865 -494 -1819 -332
rect -2119 -730 -2043 -722
rect -2119 -735 -1925 -730
rect -2119 -736 -2105 -735
rect -2526 -757 -2324 -740
rect -2526 -790 -2479 -757
rect -2601 -803 -2577 -790
rect -2531 -803 -2479 -790
rect -2433 -803 -2381 -757
rect -2335 -803 -2324 -757
rect -2601 -806 -2324 -803
rect -2600 -820 -2324 -806
rect -2269 -781 -2105 -736
rect -2057 -743 -1925 -735
rect -2057 -781 -1998 -743
rect -2269 -789 -1998 -781
rect -1952 -789 -1925 -743
rect -2269 -799 -1925 -789
rect -4159 -882 -3979 -869
rect -4159 -941 -4149 -882
rect -4090 -941 -3979 -882
rect -4159 -999 -3979 -941
rect -3275 -947 -3179 -842
rect -4159 -1053 -4145 -999
rect -4091 -1049 -3979 -999
rect -4091 -1053 -4082 -1049
rect -4159 -1065 -4082 -1053
rect -4268 -1314 -4222 -1257
rect -4025 -1083 -3979 -1049
rect -3865 -949 -3179 -947
rect -3049 -949 -2839 -948
rect -3865 -958 -2839 -949
rect -3865 -1014 -3039 -958
rect -2983 -959 -2839 -958
rect -2983 -1014 -2921 -959
rect -3865 -1015 -2921 -1014
rect -2865 -1015 -2839 -959
rect -3865 -1024 -2839 -1015
rect -3865 -1026 -3179 -1024
rect -3049 -1025 -2839 -1024
rect -3865 -1083 -3819 -1026
rect -4158 -1314 -4083 -1300
rect -4268 -1315 -4083 -1314
rect -4268 -1360 -4143 -1315
rect -4268 -1419 -4222 -1360
rect -4158 -1361 -4143 -1360
rect -4097 -1361 -4083 -1315
rect -4158 -1374 -4083 -1361
rect -4268 -1650 -4222 -1593
rect -4025 -1419 -3979 -1257
rect -3866 -1257 -3865 -1239
rect -3866 -1285 -3819 -1257
rect -4158 -1650 -4083 -1636
rect -4268 -1651 -4083 -1650
rect -4268 -1696 -4143 -1651
rect -4268 -1755 -4222 -1696
rect -4158 -1697 -4143 -1696
rect -4097 -1697 -4083 -1651
rect -4158 -1710 -4083 -1697
rect -4268 -1986 -4222 -1929
rect -4025 -1755 -3979 -1593
rect -4158 -1986 -4083 -1972
rect -4268 -1987 -4083 -1986
rect -4268 -2032 -4143 -1987
rect -4268 -2091 -4222 -2032
rect -4158 -2033 -4143 -2032
rect -4097 -2033 -4083 -1987
rect -4158 -2046 -4083 -2033
rect -4268 -2276 -4222 -2265
rect -4025 -2091 -3979 -1929
rect -4025 -2322 -3979 -2265
rect -3865 -1419 -3819 -1285
rect -3865 -1755 -3819 -1593
rect -3865 -2091 -3819 -1929
rect -3865 -2276 -3819 -2265
rect -3705 -1083 -3659 -1072
rect -3546 -1083 -3499 -1026
rect -3705 -1419 -3659 -1257
rect -3705 -1755 -3659 -1593
rect -3705 -2091 -3659 -1929
rect -3705 -2322 -3659 -2265
rect -3545 -1419 -3499 -1257
rect -3545 -1755 -3499 -1593
rect -3545 -2091 -3499 -1929
rect -3545 -2276 -3499 -2265
rect -3385 -1083 -3339 -1072
rect -3226 -1083 -3179 -1026
rect -3385 -1419 -3339 -1257
rect -3385 -1755 -3339 -1593
rect -3385 -2091 -3339 -1929
rect -3385 -2322 -3339 -2265
rect -3225 -1419 -3179 -1257
rect -3225 -1755 -3179 -1593
rect -3225 -2091 -3179 -1929
rect -3225 -2276 -3179 -2265
rect -3065 -1083 -3019 -1072
rect -3065 -1419 -3019 -1257
rect -3065 -1755 -3019 -1593
rect -3065 -2091 -3019 -1929
rect -3065 -2322 -3019 -2265
rect -4025 -2370 -3019 -2322
rect -2429 -1076 -2383 -1065
rect -2429 -1412 -2383 -1250
rect -2429 -1748 -2383 -1586
rect -2429 -2084 -2383 -1922
rect -2429 -2412 -2383 -2258
rect -2269 -1076 -2223 -799
rect -2119 -802 -1925 -799
rect -2269 -1412 -2223 -1250
rect -2269 -1748 -2223 -1586
rect -2269 -2084 -2223 -1922
rect -2269 -2269 -2223 -2258
rect -2025 -1076 -1979 -1065
rect -2025 -1412 -1979 -1250
rect -2025 -1748 -1979 -1586
rect -2025 -2084 -1979 -1922
rect -2025 -2412 -1979 -2258
rect -1865 -1076 -1819 -668
rect -1622 -158 -1576 -100
rect -1622 -494 -1576 -332
rect -1622 -862 -1576 -668
rect -1462 -158 -1416 -147
rect -1462 -494 -1416 -332
rect -1462 -726 -1416 -668
rect -1302 -158 -1256 -100
rect -1302 -494 -1256 -332
rect -1302 -679 -1256 -668
rect -1142 -158 -1096 -147
rect -1142 -494 -1096 -332
rect -1142 -726 -1096 -668
rect -982 -158 -936 -100
rect -982 -494 -936 -332
rect -982 -679 -936 -668
rect -822 -158 -776 -147
rect -822 -494 -776 -332
rect -822 -726 -776 -668
rect -662 -158 -616 -100
rect -662 -494 -616 -332
rect -662 -679 -616 -668
rect -1462 -835 -776 -726
rect -1756 -875 -1576 -862
rect -1756 -934 -1746 -875
rect -1687 -934 -1576 -875
rect -1756 -992 -1576 -934
rect -872 -940 -776 -835
rect -1756 -1046 -1742 -992
rect -1688 -1042 -1576 -992
rect -1688 -1046 -1679 -1042
rect -1756 -1058 -1679 -1046
rect -1865 -1307 -1819 -1250
rect -1622 -1076 -1576 -1042
rect -1462 -942 -776 -940
rect -1462 -950 -436 -942
rect -1462 -1006 -621 -950
rect -565 -1006 -502 -950
rect -446 -1006 -436 -950
rect -1462 -1017 -436 -1006
rect -98 -983 -40 732
rect 170 495 216 657
rect 170 169 216 321
rect 330 831 376 1239
rect 573 1413 619 1575
rect 733 2421 779 2432
rect 733 2085 779 2247
rect 733 1749 779 1911
rect 733 1441 779 1575
rect 732 1413 779 1441
rect 732 1395 733 1413
rect 438 1209 517 1221
rect 438 1155 453 1209
rect 507 1205 517 1209
rect 573 1205 619 1239
rect 507 1158 619 1205
rect 507 1155 517 1158
rect 438 1099 517 1155
rect 438 1045 453 1099
rect 507 1045 517 1099
rect 438 1033 517 1045
rect 330 495 376 657
rect 330 310 376 321
rect 573 831 619 1158
rect 733 1182 779 1239
rect 893 2421 939 2478
rect 893 2085 939 2247
rect 893 1749 939 1911
rect 893 1413 939 1575
rect 1053 2421 1099 2432
rect 1053 2085 1099 2247
rect 1053 1749 1099 1911
rect 1053 1413 1099 1575
rect 893 1228 939 1239
rect 1052 1182 1099 1239
rect 1213 2421 1259 2478
rect 1213 2085 1259 2247
rect 1213 1749 1259 1911
rect 1213 1413 1259 1575
rect 1373 2421 1419 2432
rect 1373 2085 1419 2247
rect 1373 1749 1419 1911
rect 1373 1413 1419 1575
rect 1213 1228 1259 1239
rect 1372 1182 1419 1239
rect 1533 2421 1579 2478
rect 1533 2085 1579 2247
rect 1533 1749 1579 1911
rect 1533 1413 1579 1575
rect 1533 1228 1579 1239
rect 1930 2478 2936 2526
rect 1930 2421 1976 2478
rect 1930 2085 1976 2247
rect 1930 1749 1976 1911
rect 1930 1413 1976 1575
rect 1930 1228 1976 1239
rect 2090 2421 2136 2432
rect 2090 2085 2136 2247
rect 2090 1749 2136 1911
rect 2090 1413 2136 1575
rect 2250 2421 2296 2478
rect 2250 2085 2296 2247
rect 2250 1749 2296 1911
rect 2250 1413 2296 1575
rect 733 1180 1419 1182
rect 2090 1182 2137 1239
rect 2250 1228 2296 1239
rect 2410 2421 2456 2432
rect 2410 2085 2456 2247
rect 2410 1749 2456 1911
rect 2410 1413 2456 1575
rect 2570 2421 2616 2478
rect 2570 2085 2616 2247
rect 2570 1749 2616 1911
rect 2570 1413 2616 1575
rect 2410 1182 2457 1239
rect 2570 1228 2616 1239
rect 2730 2421 2776 2432
rect 2730 2085 2776 2247
rect 2730 1749 2776 1911
rect 2730 1441 2776 1575
rect 2890 2421 2936 2478
rect 2890 2085 2936 2247
rect 3133 2421 3179 2432
rect 2994 2189 3069 2202
rect 2994 2143 3008 2189
rect 3054 2188 3069 2189
rect 3133 2188 3179 2247
rect 3054 2143 3179 2188
rect 2994 2142 3179 2143
rect 2994 2128 3069 2142
rect 2890 1749 2936 1911
rect 3133 2085 3179 2142
rect 2994 1853 3069 1866
rect 2994 1807 3008 1853
rect 3054 1852 3069 1853
rect 3133 1852 3179 1911
rect 3054 1807 3179 1852
rect 2994 1806 3179 1807
rect 2994 1792 3069 1806
rect 2730 1413 2777 1441
rect 2776 1395 2777 1413
rect 2890 1413 2936 1575
rect 3133 1749 3179 1806
rect 2994 1517 3069 1530
rect 2994 1471 3008 1517
rect 3054 1516 3069 1517
rect 3133 1516 3179 1575
rect 3054 1471 3179 1516
rect 2994 1470 3179 1471
rect 2994 1456 3069 1470
rect 2730 1182 2776 1239
rect 2090 1180 2776 1182
rect 733 1105 2776 1180
rect 733 1103 1419 1105
rect 1323 998 1419 1103
rect 573 495 619 657
rect 573 263 619 321
rect 733 889 1419 998
rect 733 831 779 889
rect 733 495 779 657
rect 733 310 779 321
rect 893 831 939 842
rect 893 495 939 657
rect 893 263 939 321
rect 1053 831 1099 889
rect 1053 495 1099 657
rect 1053 310 1099 321
rect 1213 831 1259 842
rect 1213 495 1259 657
rect 1213 263 1259 321
rect 1373 831 1419 889
rect 1373 495 1419 657
rect 1373 310 1419 321
rect 1533 831 1579 842
rect 1533 495 1579 657
rect 1533 263 1579 321
rect 573 215 1579 263
rect 1708 415 1788 1105
rect 2090 1103 2776 1105
rect 3133 1413 3179 1470
rect 2890 1205 2936 1239
rect 2995 1319 3070 1331
rect 2995 1265 3002 1319
rect 3056 1265 3070 1319
rect 2995 1221 3070 1265
rect 2993 1209 3070 1221
rect 2993 1205 3002 1209
rect 2890 1158 3002 1205
rect 2090 998 2186 1103
rect 2090 889 2776 998
rect 1708 360 1721 415
rect 1776 360 1788 415
rect 1708 305 1788 360
rect 1708 250 1721 305
rect 1776 250 1788 305
rect 1708 238 1788 250
rect 1930 831 1976 842
rect 1930 495 1976 657
rect 1930 263 1976 321
rect 2090 831 2136 889
rect 2090 495 2136 657
rect 2090 310 2136 321
rect 2250 831 2296 842
rect 2250 495 2296 657
rect 2250 263 2296 321
rect 2410 831 2456 889
rect 2410 495 2456 657
rect 2410 310 2456 321
rect 2570 831 2616 842
rect 2570 495 2616 657
rect 2570 263 2616 321
rect 2730 831 2776 889
rect 2730 495 2776 657
rect 2730 310 2776 321
rect 2890 831 2936 1158
rect 2993 1155 3002 1158
rect 3056 1155 3070 1209
rect 2993 1143 3070 1155
rect 2995 1142 3070 1143
rect 2890 495 2936 657
rect 2890 263 2936 321
rect 3133 831 3179 1239
rect 3293 2421 3339 2575
rect 3293 2085 3339 2247
rect 3293 1749 3339 1911
rect 3293 1413 3339 1575
rect 3743 2421 3789 2575
rect 5511 2574 7118 2575
rect 7503 2731 7676 2748
rect 7503 2675 7507 2731
rect 7563 2675 7617 2731
rect 7673 2675 7676 2731
rect 7503 2621 7676 2675
rect 4146 2478 5152 2526
rect 3743 2085 3789 2247
rect 3743 1749 3789 1911
rect 3743 1413 3789 1575
rect 3293 1228 3339 1239
rect 3385 1320 3462 1332
rect 3385 1264 3395 1320
rect 3451 1264 3462 1320
rect 3385 1210 3462 1264
rect 3385 1154 3395 1210
rect 3451 1188 3462 1210
rect 3620 1320 3696 1332
rect 3620 1264 3631 1320
rect 3687 1264 3696 1320
rect 3620 1223 3696 1264
rect 3743 1228 3789 1239
rect 3903 2421 3949 2432
rect 3903 2188 3949 2247
rect 4146 2421 4192 2478
rect 4013 2189 4088 2202
rect 4013 2188 4028 2189
rect 3903 2143 4028 2188
rect 4074 2143 4088 2189
rect 3903 2142 4088 2143
rect 3903 2085 3949 2142
rect 4013 2128 4088 2142
rect 3903 1852 3949 1911
rect 4146 2085 4192 2247
rect 4013 1853 4088 1866
rect 4013 1852 4028 1853
rect 3903 1807 4028 1852
rect 4074 1807 4088 1853
rect 3903 1806 4088 1807
rect 3903 1749 3949 1806
rect 4013 1792 4088 1806
rect 3903 1516 3949 1575
rect 4146 1749 4192 1911
rect 4013 1517 4088 1530
rect 4013 1516 4028 1517
rect 3903 1471 4028 1516
rect 4074 1471 4088 1517
rect 3903 1470 4088 1471
rect 3903 1413 3949 1470
rect 4013 1456 4088 1470
rect 3620 1210 3697 1223
rect 3620 1188 3631 1210
rect 3451 1154 3518 1188
rect 3385 1135 3518 1154
rect 3462 1134 3518 1135
rect 3564 1154 3631 1188
rect 3687 1154 3697 1210
rect 3564 1135 3697 1154
rect 3564 1134 3696 1135
rect 3239 952 3433 965
rect 3239 906 3266 952
rect 3312 945 3433 952
rect 3649 952 3843 965
rect 3649 945 3770 952
rect 3312 944 3770 945
rect 3312 906 3371 944
rect 3239 898 3371 906
rect 3419 898 3663 944
rect 3711 906 3770 944
rect 3816 906 3843 952
rect 3711 898 3843 906
rect 3239 896 3843 898
rect 3239 893 3433 896
rect 3357 885 3433 893
rect 3484 895 3575 896
rect 3133 495 3179 657
rect 3133 310 3179 321
rect 3293 831 3339 842
rect 3293 495 3339 657
rect 3484 466 3530 895
rect 3649 893 3843 896
rect 3649 885 3725 893
rect 3743 831 3789 842
rect 3743 495 3789 657
rect 1930 215 2936 263
rect 3293 169 3339 321
rect 3470 454 3543 466
rect 3470 400 3480 454
rect 3534 400 3543 454
rect 3470 344 3543 400
rect 3470 290 3480 344
rect 3534 290 3543 344
rect 3470 277 3543 290
rect 3743 169 3789 321
rect 3903 831 3949 1239
rect 4146 1413 4192 1575
rect 4306 2421 4352 2432
rect 4306 2085 4352 2247
rect 4306 1749 4352 1911
rect 4306 1441 4352 1575
rect 4305 1413 4352 1441
rect 4305 1395 4306 1413
rect 4012 1209 4089 1221
rect 4012 1155 4026 1209
rect 4080 1205 4089 1209
rect 4146 1205 4192 1239
rect 4080 1158 4192 1205
rect 4080 1155 4089 1158
rect 4012 1143 4089 1155
rect 3903 495 3949 657
rect 3903 310 3949 321
rect 4146 831 4192 1158
rect 4306 1182 4352 1239
rect 4466 2421 4512 2478
rect 4466 2085 4512 2247
rect 4466 1749 4512 1911
rect 4466 1413 4512 1575
rect 4626 2421 4672 2432
rect 4626 2085 4672 2247
rect 4626 1749 4672 1911
rect 4626 1413 4672 1575
rect 4466 1228 4512 1239
rect 4625 1182 4672 1239
rect 4786 2421 4832 2478
rect 4786 2085 4832 2247
rect 4786 1749 4832 1911
rect 4786 1413 4832 1575
rect 4946 2421 4992 2432
rect 4946 2085 4992 2247
rect 4946 1749 4992 1911
rect 4946 1413 4992 1575
rect 4786 1228 4832 1239
rect 4945 1182 4992 1239
rect 5106 2421 5152 2478
rect 5106 2085 5152 2247
rect 5106 1749 5152 1911
rect 5106 1413 5152 1575
rect 5106 1228 5152 1239
rect 5610 2477 6616 2525
rect 5610 2420 5656 2477
rect 5610 2084 5656 2246
rect 5610 1748 5656 1910
rect 5610 1412 5656 1574
rect 5610 1227 5656 1238
rect 5770 2420 5816 2431
rect 5770 2084 5816 2246
rect 5770 1748 5816 1910
rect 5770 1412 5816 1574
rect 5930 2420 5976 2477
rect 5930 2084 5976 2246
rect 5930 1748 5976 1910
rect 5930 1412 5976 1574
rect 4306 1180 4992 1182
rect 5770 1181 5817 1238
rect 5930 1227 5976 1238
rect 6090 2420 6136 2431
rect 6090 2084 6136 2246
rect 6090 1748 6136 1910
rect 6090 1412 6136 1574
rect 6250 2420 6296 2477
rect 6250 2084 6296 2246
rect 6250 1748 6296 1910
rect 6250 1412 6296 1574
rect 6090 1181 6137 1238
rect 6250 1227 6296 1238
rect 6410 2420 6456 2431
rect 6410 2084 6456 2246
rect 6410 1748 6456 1910
rect 6410 1440 6456 1574
rect 6570 2420 6616 2477
rect 6570 2084 6616 2246
rect 6813 2420 6859 2431
rect 6674 2188 6749 2201
rect 6674 2142 6688 2188
rect 6734 2187 6749 2188
rect 6813 2187 6859 2246
rect 6734 2142 6859 2187
rect 6674 2141 6859 2142
rect 6674 2127 6749 2141
rect 6570 1748 6616 1910
rect 6813 2084 6859 2141
rect 6674 1852 6749 1865
rect 6674 1806 6688 1852
rect 6734 1851 6749 1852
rect 6813 1851 6859 1910
rect 6734 1806 6859 1851
rect 6674 1805 6859 1806
rect 6674 1791 6749 1805
rect 6410 1412 6457 1440
rect 6456 1394 6457 1412
rect 6570 1412 6616 1574
rect 6813 1748 6859 1805
rect 6674 1516 6749 1529
rect 6674 1470 6688 1516
rect 6734 1515 6749 1516
rect 6813 1515 6859 1574
rect 6734 1470 6859 1515
rect 6674 1469 6859 1470
rect 6674 1455 6749 1469
rect 6410 1181 6456 1238
rect 4306 1179 5331 1180
rect 5770 1179 6456 1181
rect 4306 1105 6456 1179
rect 4306 1103 4992 1105
rect 4896 998 4992 1103
rect 4146 495 4192 657
rect 4146 263 4192 321
rect 4306 889 4992 998
rect 4306 831 4352 889
rect 4306 495 4352 657
rect 4306 310 4352 321
rect 4466 831 4512 842
rect 4466 495 4512 657
rect 4466 263 4512 321
rect 4626 831 4672 889
rect 4626 495 4672 657
rect 4626 310 4672 321
rect 4786 831 4832 842
rect 4786 495 4832 657
rect 4786 263 4832 321
rect 4946 831 4992 889
rect 5284 1104 6456 1105
rect 4946 495 4992 657
rect 4946 310 4992 321
rect 5106 831 5152 842
rect 5106 495 5152 657
rect 5284 415 5364 1104
rect 5770 1102 6456 1104
rect 6813 1412 6859 1469
rect 6570 1204 6616 1238
rect 6673 1328 6750 1339
rect 6673 1274 6685 1328
rect 6739 1274 6750 1328
rect 6673 1208 6750 1274
rect 6673 1204 6682 1208
rect 6570 1157 6682 1204
rect 5770 997 5866 1102
rect 5770 888 6456 997
rect 5610 830 5656 841
rect 5610 494 5656 656
rect 5106 263 5152 321
rect 4146 215 5152 263
rect 5285 402 5365 415
rect 5285 346 5297 402
rect 5353 346 5365 402
rect 5285 292 5365 346
rect 5285 236 5297 292
rect 5353 236 5365 292
rect 5285 224 5365 236
rect 5610 262 5656 320
rect 5770 830 5816 888
rect 5770 494 5816 656
rect 5770 309 5816 320
rect 5930 830 5976 841
rect 5930 494 5976 656
rect 5930 262 5976 320
rect 6090 830 6136 888
rect 6090 494 6136 656
rect 6090 309 6136 320
rect 6250 830 6296 841
rect 6250 494 6296 656
rect 6250 262 6296 320
rect 6410 830 6456 888
rect 6410 494 6456 656
rect 6410 309 6456 320
rect 6570 830 6616 1157
rect 6673 1154 6682 1157
rect 6736 1154 6750 1208
rect 6673 1142 6750 1154
rect 6570 494 6616 656
rect 6570 262 6616 320
rect 6813 830 6859 1238
rect 6973 2420 7019 2574
rect 7503 2565 7507 2621
rect 7563 2565 7617 2621
rect 7673 2565 7676 2621
rect 7503 2511 7676 2565
rect 7503 2455 7507 2511
rect 7563 2455 7617 2511
rect 7673 2455 7676 2511
rect 7503 2443 7676 2455
rect 6973 2084 7019 2246
rect 6973 1748 7019 1910
rect 6973 1412 7019 1574
rect 6973 1227 7019 1238
rect 7065 1319 7142 1357
rect 7065 1263 7075 1319
rect 7131 1263 7142 1319
rect 7065 1209 7142 1263
rect 7065 1153 7075 1209
rect 7131 1187 7142 1209
rect 7131 1153 7198 1187
rect 7065 1134 7198 1153
rect 7142 1133 7198 1134
rect 6919 951 7113 964
rect 6919 905 6946 951
rect 6992 944 7113 951
rect 6992 943 7234 944
rect 6992 905 7051 943
rect 6919 897 7051 905
rect 7099 915 7234 943
rect 7099 897 7161 915
rect 6919 892 7161 897
rect 7037 884 7161 892
rect 7144 858 7161 884
rect 7218 858 7234 915
rect 6813 494 6859 656
rect 6813 309 6859 320
rect 6973 830 7019 841
rect 7144 805 7234 858
rect 7144 748 7161 805
rect 7218 748 7234 805
rect 7144 739 7234 748
rect 7505 791 7676 2443
rect 7505 774 7678 791
rect 6973 494 7019 656
rect 5610 214 6616 262
rect 71 168 5251 169
rect 6973 168 7019 320
rect 7505 718 7509 774
rect 7565 718 7619 774
rect 7675 718 7678 774
rect 7505 664 7678 718
rect 7505 608 7509 664
rect 7565 608 7619 664
rect 7675 608 7678 664
rect 7505 554 7678 608
rect 7505 498 7509 554
rect 7565 498 7619 554
rect 7675 498 7678 554
rect 7505 486 7678 498
rect 71 114 7412 168
rect 70 58 80 114
rect 136 109 190 114
rect 246 109 300 114
rect 356 109 410 114
rect 466 109 520 114
rect 576 109 7412 114
rect 292 58 300 109
rect 513 58 520 109
rect 71 55 131 58
rect 292 55 352 58
rect 513 55 573 58
rect 734 55 794 109
rect 955 55 1015 109
rect 1176 55 1236 109
rect 1397 55 1457 109
rect 1618 55 1891 109
rect 2052 55 2112 109
rect 2273 55 2333 109
rect 2494 55 2554 109
rect 2715 55 2775 109
rect 2936 55 2996 109
rect 3157 55 3217 109
rect 3378 55 3704 109
rect 3865 55 3925 109
rect 4086 55 4146 109
rect 4307 55 4367 109
rect 4528 55 4588 109
rect 4749 55 4809 109
rect 4970 55 5030 109
rect 5191 108 7412 109
rect 5191 55 5571 108
rect 71 54 5571 55
rect 5732 54 5792 108
rect 5953 54 6013 108
rect 6174 54 6234 108
rect 6395 54 6455 108
rect 6616 54 6676 108
rect 6837 54 6897 108
rect 7058 54 7412 108
rect 71 -5 7412 54
rect 61 -102 945 -61
rect 61 -103 849 -102
rect 61 -163 124 -103
rect 905 -158 945 -102
rect 871 -163 945 -158
rect 61 -200 945 -163
rect 160 -343 206 -200
rect 160 -679 206 -517
rect 160 -864 206 -853
rect 320 -343 366 -332
rect 320 -679 366 -517
rect 189 -983 266 -973
rect -98 -986 266 -983
rect -1462 -1019 -776 -1017
rect -1462 -1076 -1416 -1019
rect -1755 -1307 -1680 -1293
rect -1865 -1308 -1680 -1307
rect -1865 -1353 -1740 -1308
rect -1865 -1412 -1819 -1353
rect -1755 -1354 -1740 -1353
rect -1694 -1354 -1680 -1308
rect -1755 -1367 -1680 -1354
rect -1865 -1643 -1819 -1586
rect -1622 -1412 -1576 -1250
rect -1463 -1250 -1462 -1232
rect -1463 -1278 -1416 -1250
rect -1755 -1643 -1680 -1629
rect -1865 -1644 -1680 -1643
rect -1865 -1689 -1740 -1644
rect -1865 -1748 -1819 -1689
rect -1755 -1690 -1740 -1689
rect -1694 -1690 -1680 -1644
rect -1755 -1703 -1680 -1690
rect -1865 -1979 -1819 -1922
rect -1622 -1748 -1576 -1586
rect -1755 -1979 -1680 -1965
rect -1865 -1980 -1680 -1979
rect -1865 -2025 -1740 -1980
rect -1865 -2084 -1819 -2025
rect -1755 -2026 -1740 -2025
rect -1694 -2026 -1680 -1980
rect -1755 -2039 -1680 -2026
rect -1865 -2269 -1819 -2258
rect -1622 -2084 -1576 -1922
rect -1622 -2315 -1576 -2258
rect -1462 -1412 -1416 -1278
rect -1462 -1748 -1416 -1586
rect -1462 -2084 -1416 -1922
rect -1462 -2269 -1416 -2258
rect -1302 -1076 -1256 -1065
rect -1143 -1076 -1096 -1019
rect -1302 -1412 -1256 -1250
rect -1302 -1748 -1256 -1586
rect -1302 -2084 -1256 -1922
rect -1302 -2315 -1256 -2258
rect -1142 -1412 -1096 -1250
rect -1142 -1748 -1096 -1586
rect -1142 -2084 -1096 -1922
rect -1142 -2269 -1096 -2258
rect -982 -1076 -936 -1065
rect -823 -1076 -776 -1019
rect -98 -1029 205 -986
rect -98 -1030 51 -1029
rect -982 -1412 -936 -1250
rect -982 -1748 -936 -1586
rect -982 -2084 -936 -1922
rect -982 -2315 -936 -2258
rect -822 -1412 -776 -1250
rect -822 -1748 -776 -1586
rect -822 -2084 -776 -1922
rect -822 -2269 -776 -2258
rect -662 -1076 -616 -1065
rect -662 -1412 -616 -1250
rect -98 -1509 -40 -1030
rect 189 -1035 205 -1029
rect 252 -1035 266 -986
rect 189 -1050 266 -1035
rect 320 -984 366 -853
rect 480 -343 526 -200
rect 480 -679 526 -517
rect 480 -864 526 -853
rect 640 -343 686 -332
rect 640 -679 686 -517
rect 640 -984 686 -853
rect 800 -343 846 -200
rect 991 -354 1178 -341
rect 991 -408 1004 -354
rect 1058 -408 1114 -354
rect 1168 -408 1178 -354
rect 991 -420 1178 -408
rect 800 -679 846 -517
rect 800 -864 846 -853
rect 1008 -984 1054 -420
rect 1326 -491 1407 -481
rect 1326 -548 1338 -491
rect 1395 -548 1407 -491
rect 1326 -601 1407 -548
rect 1106 -618 1178 -607
rect 1106 -672 1115 -618
rect 1169 -672 1178 -618
rect 1326 -658 1338 -601
rect 1395 -658 1407 -601
rect 1326 -670 1407 -658
rect 1106 -728 1178 -672
rect 1106 -782 1115 -728
rect 1169 -782 1178 -728
rect 1106 -795 1178 -782
rect 320 -1030 1054 -984
rect 160 -1128 206 -1117
rect 160 -1364 206 -1202
rect -662 -1748 -616 -1586
rect -126 -1519 -31 -1509
rect -126 -1575 -101 -1519
rect -45 -1575 -31 -1519
rect 160 -1531 206 -1438
rect 320 -1128 366 -1030
rect 320 -1364 366 -1202
rect 320 -1449 366 -1438
rect 480 -1128 526 -1117
rect 480 -1364 526 -1202
rect 480 -1531 526 -1438
rect 640 -1128 686 -1030
rect 640 -1364 686 -1202
rect 640 -1449 686 -1438
rect 800 -1128 846 -1117
rect 800 -1364 846 -1202
rect 800 -1531 846 -1438
rect -126 -1629 -31 -1575
rect -126 -1685 -101 -1629
rect -45 -1685 -31 -1629
rect 61 -1576 945 -1531
rect 61 -1631 115 -1576
rect 879 -1577 945 -1576
rect 61 -1634 452 -1631
rect 508 -1633 587 -1631
rect 643 -1632 717 -1631
rect 773 -1632 860 -1631
rect 643 -1633 860 -1632
rect 916 -1633 945 -1577
rect 508 -1634 945 -1633
rect 61 -1676 945 -1634
rect -126 -1695 -31 -1685
rect -662 -2084 -616 -1922
rect -340 -2019 -150 -2011
rect -340 -2075 -328 -2019
rect -272 -2075 -218 -2019
rect -162 -2075 -150 -2019
rect -340 -2082 -150 -2075
rect -662 -2315 -616 -2258
rect -1622 -2363 -616 -2315
rect -2528 -2419 -517 -2412
rect -4931 -2471 -517 -2419
rect -4931 -2472 -1080 -2471
rect -1024 -2472 -970 -2471
rect -914 -2472 -860 -2471
rect -804 -2472 -750 -2471
rect -694 -2472 -640 -2471
rect -584 -2472 -517 -2471
rect -4931 -2479 -2285 -2472
rect -4931 -2533 -4688 -2479
rect -4527 -2533 -4467 -2479
rect -4306 -2533 -4246 -2479
rect -4085 -2533 -4025 -2479
rect -3864 -2533 -3804 -2479
rect -3643 -2533 -3583 -2479
rect -3422 -2533 -3362 -2479
rect -3201 -2533 -3141 -2479
rect -2980 -2526 -2285 -2479
rect -2124 -2526 -2064 -2472
rect -1903 -2526 -1843 -2472
rect -1682 -2526 -1622 -2472
rect -1461 -2526 -1401 -2472
rect -1240 -2526 -1180 -2472
rect -1019 -2526 -970 -2472
rect -798 -2526 -750 -2472
rect -577 -2526 -517 -2472
rect -2980 -2527 -1080 -2526
rect -1024 -2527 -970 -2526
rect -914 -2527 -860 -2526
rect -804 -2527 -750 -2526
rect -694 -2527 -640 -2526
rect -584 -2527 -517 -2526
rect -2980 -2533 -517 -2527
rect -4931 -2586 -517 -2533
rect -4931 -2593 -2920 -2586
rect -4832 -2747 -4786 -2593
rect -4832 -3083 -4786 -2921
rect -4832 -3419 -4786 -3257
rect -4832 -3755 -4786 -3593
rect -4832 -3940 -4786 -3929
rect -4672 -2747 -4626 -2736
rect -4672 -3083 -4626 -2921
rect -4672 -3419 -4626 -3257
rect -4672 -3755 -4626 -3593
rect -5040 -4199 -4727 -4185
rect -5055 -4202 -4727 -4199
rect -5055 -4209 -4980 -4202
rect -5055 -4265 -5030 -4209
rect -4934 -4248 -4882 -4202
rect -4836 -4248 -4784 -4202
rect -4738 -4248 -4727 -4202
rect -4974 -4265 -4727 -4248
rect -4672 -4206 -4626 -3929
rect -4428 -2747 -4382 -2593
rect -4025 -2690 -3019 -2642
rect -4428 -3083 -4382 -2921
rect -4428 -3419 -4382 -3257
rect -4428 -3755 -4382 -3593
rect -4428 -3940 -4382 -3929
rect -4268 -2747 -4222 -2736
rect -4268 -2980 -4222 -2921
rect -4025 -2747 -3979 -2690
rect -4158 -2979 -4083 -2966
rect -4158 -2980 -4143 -2979
rect -4268 -3025 -4143 -2980
rect -4097 -3025 -4083 -2979
rect -4268 -3026 -4083 -3025
rect -4268 -3083 -4222 -3026
rect -4158 -3040 -4083 -3026
rect -4268 -3316 -4222 -3257
rect -4025 -3083 -3979 -2921
rect -4158 -3315 -4083 -3302
rect -4158 -3316 -4143 -3315
rect -4268 -3361 -4143 -3316
rect -4097 -3361 -4083 -3315
rect -4268 -3362 -4083 -3361
rect -4268 -3419 -4222 -3362
rect -4158 -3376 -4083 -3362
rect -4268 -3652 -4222 -3593
rect -4025 -3419 -3979 -3257
rect -4158 -3651 -4083 -3638
rect -4158 -3652 -4143 -3651
rect -4268 -3697 -4143 -3652
rect -4097 -3697 -4083 -3651
rect -4268 -3698 -4083 -3697
rect -4268 -3755 -4222 -3698
rect -4158 -3712 -4083 -3698
rect -4522 -4206 -4328 -4203
rect -4672 -4216 -4328 -4206
rect -4672 -4224 -4401 -4216
rect -5055 -4319 -4960 -4265
rect -5055 -4375 -5030 -4319
rect -4974 -4375 -4960 -4319
rect -4672 -4269 -4508 -4224
rect -5055 -4385 -4960 -4375
rect -4832 -4337 -4786 -4326
rect -5235 -5518 -5162 -5506
rect -5376 -5575 -5225 -5518
rect -5168 -5575 -5162 -5518
rect -5235 -5628 -5162 -5575
rect -5235 -5685 -5225 -5628
rect -5168 -5685 -5162 -5628
rect -5235 -5697 -5162 -5685
rect -5040 -5768 -4978 -4385
rect -4832 -4673 -4786 -4511
rect -4832 -4999 -4786 -4847
rect -4672 -4337 -4626 -4269
rect -4522 -4270 -4508 -4269
rect -4460 -4262 -4401 -4224
rect -4355 -4262 -4328 -4216
rect -4460 -4270 -4328 -4262
rect -4522 -4275 -4328 -4270
rect -4522 -4283 -4446 -4275
rect -4672 -4673 -4626 -4511
rect -4672 -4858 -4626 -4847
rect -4428 -4337 -4382 -4326
rect -4428 -4673 -4382 -4511
rect -4428 -4999 -4382 -4847
rect -4268 -4337 -4222 -3929
rect -4025 -3755 -3979 -3593
rect -3865 -2747 -3819 -2736
rect -3865 -3083 -3819 -2921
rect -3865 -3419 -3819 -3257
rect -3865 -3727 -3819 -3593
rect -3866 -3755 -3819 -3727
rect -3866 -3773 -3865 -3755
rect -4159 -3959 -4082 -3947
rect -4159 -4013 -4145 -3959
rect -4091 -3963 -4082 -3959
rect -4025 -3963 -3979 -3929
rect -4091 -4013 -3979 -3963
rect -4159 -4071 -3979 -4013
rect -3865 -3986 -3819 -3929
rect -3705 -2747 -3659 -2690
rect -3705 -3083 -3659 -2921
rect -3705 -3419 -3659 -3257
rect -3705 -3755 -3659 -3593
rect -3545 -2747 -3499 -2736
rect -3545 -3083 -3499 -2921
rect -3545 -3419 -3499 -3257
rect -3545 -3755 -3499 -3593
rect -3705 -3940 -3659 -3929
rect -3546 -3986 -3499 -3929
rect -3385 -2747 -3339 -2690
rect -3385 -3083 -3339 -2921
rect -3385 -3419 -3339 -3257
rect -3385 -3755 -3339 -3593
rect -3225 -2747 -3179 -2736
rect -3225 -3083 -3179 -2921
rect -3225 -3419 -3179 -3257
rect -3225 -3755 -3179 -3593
rect -3385 -3940 -3339 -3929
rect -3226 -3986 -3179 -3929
rect -3065 -2747 -3019 -2690
rect -3065 -3083 -3019 -2921
rect -3065 -3419 -3019 -3257
rect -3065 -3755 -3019 -3593
rect -3065 -3940 -3019 -3929
rect -2429 -2740 -2383 -2586
rect -2429 -3076 -2383 -2914
rect -2429 -3412 -2383 -3250
rect -2429 -3748 -2383 -3586
rect -2429 -3933 -2383 -3922
rect -2269 -2740 -2223 -2729
rect -2269 -3076 -2223 -2914
rect -2269 -3412 -2223 -3250
rect -2269 -3748 -2223 -3586
rect -3865 -3988 -3179 -3986
rect -3865 -3997 -2840 -3988
rect -3865 -4053 -3040 -3997
rect -2984 -4053 -2919 -3997
rect -2863 -4053 -2840 -3997
rect -3865 -4063 -2840 -4053
rect -3865 -4065 -3179 -4063
rect -4159 -4130 -4149 -4071
rect -4090 -4130 -3979 -4071
rect -4159 -4143 -3979 -4130
rect -4268 -4673 -4222 -4511
rect -4268 -4858 -4222 -4847
rect -4025 -4337 -3979 -4143
rect -3275 -4170 -3179 -4065
rect -4025 -4673 -3979 -4511
rect -4025 -4905 -3979 -4847
rect -3865 -4279 -3179 -4170
rect -2600 -4190 -2324 -4178
rect -3865 -4337 -3819 -4279
rect -3865 -4673 -3819 -4511
rect -3865 -4858 -3819 -4847
rect -3705 -4337 -3659 -4326
rect -3705 -4673 -3659 -4511
rect -3705 -4905 -3659 -4847
rect -3545 -4337 -3499 -4279
rect -3545 -4673 -3499 -4511
rect -3545 -4858 -3499 -4847
rect -3385 -4337 -3339 -4326
rect -3385 -4673 -3339 -4511
rect -3385 -4905 -3339 -4847
rect -3225 -4337 -3179 -4279
rect -2620 -4195 -2324 -4190
rect -2620 -4200 -2577 -4195
rect -2620 -4256 -2595 -4200
rect -2531 -4241 -2479 -4195
rect -2433 -4241 -2381 -4195
rect -2335 -4241 -2324 -4195
rect -2539 -4256 -2324 -4241
rect -2620 -4258 -2324 -4256
rect -2269 -4199 -2223 -3922
rect -2025 -2740 -1979 -2586
rect -1622 -2683 -616 -2635
rect -2025 -3076 -1979 -2914
rect -2025 -3412 -1979 -3250
rect -2025 -3748 -1979 -3586
rect -2025 -3933 -1979 -3922
rect -1865 -2740 -1819 -2729
rect -1865 -2973 -1819 -2914
rect -1622 -2740 -1576 -2683
rect -1755 -2972 -1680 -2959
rect -1755 -2973 -1740 -2972
rect -1865 -3018 -1740 -2973
rect -1694 -3018 -1680 -2972
rect -1865 -3019 -1680 -3018
rect -1865 -3076 -1819 -3019
rect -1755 -3033 -1680 -3019
rect -1865 -3309 -1819 -3250
rect -1622 -3076 -1576 -2914
rect -1755 -3308 -1680 -3295
rect -1755 -3309 -1740 -3308
rect -1865 -3354 -1740 -3309
rect -1694 -3354 -1680 -3308
rect -1865 -3355 -1680 -3354
rect -1865 -3412 -1819 -3355
rect -1755 -3369 -1680 -3355
rect -1865 -3645 -1819 -3586
rect -1622 -3412 -1576 -3250
rect -1755 -3644 -1680 -3631
rect -1755 -3645 -1740 -3644
rect -1865 -3690 -1740 -3645
rect -1694 -3690 -1680 -3644
rect -1865 -3691 -1680 -3690
rect -1865 -3748 -1819 -3691
rect -1755 -3705 -1680 -3691
rect -2119 -4199 -1925 -4196
rect -2269 -4209 -1925 -4199
rect -2269 -4217 -1998 -4209
rect -2620 -4310 -2525 -4258
rect -3225 -4673 -3179 -4511
rect -3225 -4858 -3179 -4847
rect -3065 -4337 -3019 -4326
rect -2620 -4366 -2595 -4310
rect -2539 -4366 -2525 -4310
rect -2269 -4262 -2105 -4217
rect -2620 -4376 -2525 -4366
rect -2429 -4330 -2383 -4319
rect -3065 -4673 -3019 -4511
rect -3065 -4905 -3019 -4847
rect -4025 -4953 -3019 -4905
rect -2429 -4666 -2383 -4504
rect -2429 -4992 -2383 -4840
rect -2269 -4330 -2223 -4262
rect -2119 -4263 -2105 -4262
rect -2057 -4255 -1998 -4217
rect -1952 -4255 -1925 -4209
rect -2057 -4263 -1925 -4255
rect -2119 -4268 -1925 -4263
rect -2119 -4276 -2043 -4268
rect -2269 -4666 -2223 -4504
rect -2269 -4851 -2223 -4840
rect -2025 -4330 -1979 -4319
rect -2025 -4666 -1979 -4504
rect -2025 -4992 -1979 -4840
rect -1865 -4330 -1819 -3922
rect -1622 -3748 -1576 -3586
rect -1462 -2740 -1416 -2729
rect -1462 -3076 -1416 -2914
rect -1462 -3412 -1416 -3250
rect -1462 -3720 -1416 -3586
rect -1463 -3748 -1416 -3720
rect -1463 -3766 -1462 -3748
rect -1756 -3952 -1679 -3940
rect -1756 -4006 -1742 -3952
rect -1688 -3956 -1679 -3952
rect -1622 -3956 -1576 -3922
rect -1688 -4006 -1576 -3956
rect -1756 -4064 -1576 -4006
rect -1462 -3979 -1416 -3922
rect -1302 -2740 -1256 -2683
rect -1302 -3076 -1256 -2914
rect -1302 -3412 -1256 -3250
rect -1302 -3748 -1256 -3586
rect -1142 -2740 -1096 -2729
rect -1142 -3076 -1096 -2914
rect -1142 -3412 -1096 -3250
rect -1142 -3748 -1096 -3586
rect -1302 -3933 -1256 -3922
rect -1143 -3979 -1096 -3922
rect -982 -2740 -936 -2683
rect -982 -3076 -936 -2914
rect -982 -3412 -936 -3250
rect -982 -3748 -936 -3586
rect -822 -2740 -776 -2729
rect -822 -3076 -776 -2914
rect -822 -3412 -776 -3250
rect -822 -3748 -776 -3586
rect -982 -3933 -936 -3922
rect -823 -3979 -776 -3922
rect -662 -2740 -616 -2683
rect -662 -3076 -616 -2914
rect -662 -3412 -616 -3250
rect -662 -3748 -616 -3586
rect -662 -3933 -616 -3922
rect -1462 -3981 -776 -3979
rect -1462 -3989 -437 -3981
rect -1462 -3990 -520 -3989
rect -1462 -4046 -658 -3990
rect -602 -4045 -520 -3990
rect -464 -4045 -437 -3989
rect -602 -4046 -437 -4045
rect -1462 -4056 -437 -4046
rect -1462 -4058 -776 -4056
rect -673 -4057 -437 -4056
rect -1756 -4123 -1746 -4064
rect -1687 -4123 -1576 -4064
rect -1756 -4136 -1576 -4123
rect -1865 -4666 -1819 -4504
rect -1865 -4851 -1819 -4840
rect -1622 -4330 -1576 -4136
rect -872 -4163 -776 -4058
rect -1622 -4666 -1576 -4504
rect -1622 -4898 -1576 -4840
rect -1462 -4272 -776 -4163
rect -1462 -4330 -1416 -4272
rect -1462 -4666 -1416 -4504
rect -1462 -4851 -1416 -4840
rect -1302 -4330 -1256 -4319
rect -1302 -4666 -1256 -4504
rect -1302 -4898 -1256 -4840
rect -1142 -4330 -1096 -4272
rect -1142 -4666 -1096 -4504
rect -1142 -4851 -1096 -4840
rect -982 -4330 -936 -4319
rect -982 -4666 -936 -4504
rect -982 -4898 -936 -4840
rect -822 -4330 -776 -4272
rect -822 -4666 -776 -4504
rect -822 -4851 -776 -4840
rect -662 -4330 -616 -4319
rect -340 -4336 -151 -4324
rect -340 -4396 -331 -4336
rect -271 -4396 -218 -4336
rect -158 -4396 -151 -4336
rect -340 -4408 -151 -4396
rect -662 -4666 -616 -4504
rect -662 -4898 -616 -4840
rect -1622 -4946 -616 -4898
rect -4931 -5000 -2920 -4999
rect -2528 -5000 -517 -4992
rect -4931 -5050 -517 -5000
rect -4931 -5052 -1189 -5050
rect -1133 -5052 -1079 -5050
rect -1023 -5052 -969 -5050
rect -913 -5052 -859 -5050
rect -803 -5052 -749 -5050
rect -693 -5052 -639 -5050
rect -583 -5052 -517 -5050
rect -4931 -5059 -2285 -5052
rect -4931 -5113 -4688 -5059
rect -4527 -5113 -4467 -5059
rect -4306 -5113 -4246 -5059
rect -4085 -5113 -4025 -5059
rect -3864 -5113 -3804 -5059
rect -3643 -5113 -3583 -5059
rect -3422 -5113 -3362 -5059
rect -3201 -5113 -3141 -5059
rect -2980 -5106 -2285 -5059
rect -2124 -5106 -2064 -5052
rect -1903 -5106 -1843 -5052
rect -1682 -5106 -1622 -5052
rect -1461 -5106 -1401 -5052
rect -1240 -5106 -1189 -5052
rect -1019 -5106 -969 -5052
rect -798 -5106 -749 -5052
rect -577 -5106 -517 -5052
rect -2980 -5113 -517 -5106
rect -4931 -5166 -517 -5113
rect -4931 -5173 -2378 -5166
rect -4832 -5325 -4786 -5173
rect -4832 -5661 -4786 -5499
rect -5044 -5778 -4949 -5768
rect -5044 -5834 -5019 -5778
rect -4963 -5834 -4949 -5778
rect -5044 -5888 -4949 -5834
rect -4832 -5846 -4786 -5835
rect -4672 -5325 -4626 -5314
rect -4672 -5661 -4626 -5499
rect -5044 -5944 -5019 -5888
rect -4963 -5907 -4949 -5888
rect -4672 -5903 -4626 -5835
rect -4428 -5325 -4382 -5173
rect -4025 -5267 -3019 -5219
rect -4428 -5661 -4382 -5499
rect -4428 -5846 -4382 -5835
rect -4268 -5325 -4222 -5314
rect -4268 -5661 -4222 -5499
rect -4522 -5897 -4446 -5889
rect -4522 -5902 -4328 -5897
rect -4522 -5903 -4508 -5902
rect -4963 -5924 -4727 -5907
rect -5044 -5954 -4980 -5944
rect -5040 -5970 -4980 -5954
rect -4934 -5970 -4882 -5924
rect -4836 -5970 -4784 -5924
rect -4738 -5970 -4727 -5924
rect -5040 -5986 -4727 -5970
rect -5003 -5987 -4727 -5986
rect -4672 -5948 -4508 -5903
rect -4460 -5910 -4328 -5902
rect -4460 -5948 -4401 -5910
rect -4672 -5956 -4401 -5948
rect -4355 -5956 -4328 -5910
rect -4672 -5966 -4328 -5956
rect -5128 -6049 -5051 -6041
rect -5128 -6106 -5119 -6049
rect -5062 -6106 -5051 -6049
rect -5128 -6157 -5051 -6106
rect -5382 -6159 -5051 -6157
rect -5382 -6216 -5119 -6159
rect -5062 -6216 -5051 -6159
rect -5128 -6228 -5051 -6216
rect -4832 -6243 -4786 -6232
rect -4832 -6579 -4786 -6417
rect -4832 -6915 -4786 -6753
rect -4832 -7251 -4786 -7089
rect -4832 -7579 -4786 -7425
rect -4672 -6243 -4626 -5966
rect -4522 -5969 -4328 -5966
rect -4672 -6579 -4626 -6417
rect -4672 -6915 -4626 -6753
rect -4672 -7251 -4626 -7089
rect -4672 -7436 -4626 -7425
rect -4428 -6243 -4382 -6232
rect -4428 -6579 -4382 -6417
rect -4428 -6915 -4382 -6753
rect -4428 -7251 -4382 -7089
rect -4428 -7579 -4382 -7425
rect -4268 -6243 -4222 -5835
rect -4025 -5325 -3979 -5267
rect -4025 -5661 -3979 -5499
rect -4025 -6029 -3979 -5835
rect -3865 -5325 -3819 -5314
rect -3865 -5661 -3819 -5499
rect -3865 -5893 -3819 -5835
rect -3705 -5325 -3659 -5267
rect -3705 -5661 -3659 -5499
rect -3705 -5846 -3659 -5835
rect -3545 -5325 -3499 -5314
rect -3545 -5661 -3499 -5499
rect -3545 -5893 -3499 -5835
rect -3385 -5325 -3339 -5267
rect -3385 -5661 -3339 -5499
rect -3385 -5846 -3339 -5835
rect -3225 -5325 -3179 -5314
rect -3225 -5661 -3179 -5499
rect -3225 -5893 -3179 -5835
rect -3065 -5325 -3019 -5267
rect -3065 -5661 -3019 -5499
rect -2429 -5318 -2383 -5173
rect -2429 -5654 -2383 -5492
rect -3065 -5846 -3019 -5835
rect -2626 -5782 -2531 -5772
rect -2626 -5838 -2601 -5782
rect -2545 -5838 -2531 -5782
rect -3865 -6002 -3179 -5893
rect -2626 -5892 -2531 -5838
rect -2429 -5839 -2383 -5828
rect -2269 -5318 -2223 -5307
rect -2269 -5654 -2223 -5492
rect -2626 -5948 -2601 -5892
rect -2545 -5900 -2531 -5892
rect -2269 -5896 -2223 -5828
rect -2025 -5318 -1979 -5166
rect -1622 -5260 -616 -5212
rect -2025 -5654 -1979 -5492
rect -2025 -5839 -1979 -5828
rect -1865 -5318 -1819 -5307
rect -1865 -5654 -1819 -5492
rect -2119 -5890 -2043 -5882
rect -2119 -5895 -1925 -5890
rect -2119 -5896 -2105 -5895
rect -2545 -5917 -2324 -5900
rect -2626 -5958 -2577 -5948
rect -2600 -5963 -2577 -5958
rect -2531 -5963 -2479 -5917
rect -2433 -5963 -2381 -5917
rect -2335 -5963 -2324 -5917
rect -2600 -5980 -2324 -5963
rect -2269 -5941 -2105 -5896
rect -2057 -5903 -1925 -5895
rect -2057 -5941 -1998 -5903
rect -2269 -5949 -1998 -5941
rect -1952 -5949 -1925 -5903
rect -2269 -5959 -1925 -5949
rect -4159 -6042 -3979 -6029
rect -4159 -6101 -4149 -6042
rect -4090 -6101 -3979 -6042
rect -4159 -6159 -3979 -6101
rect -3275 -6107 -3179 -6002
rect -4159 -6213 -4145 -6159
rect -4091 -6209 -3979 -6159
rect -4091 -6213 -4082 -6209
rect -4159 -6225 -4082 -6213
rect -4268 -6474 -4222 -6417
rect -4025 -6243 -3979 -6209
rect -3865 -6109 -3179 -6107
rect -3865 -6117 -2840 -6109
rect -3865 -6173 -3038 -6117
rect -2982 -6173 -2908 -6117
rect -2852 -6173 -2840 -6117
rect -3865 -6184 -2840 -6173
rect -3865 -6186 -3179 -6184
rect -3865 -6243 -3819 -6186
rect -4158 -6474 -4083 -6460
rect -4268 -6475 -4083 -6474
rect -4268 -6520 -4143 -6475
rect -4268 -6579 -4222 -6520
rect -4158 -6521 -4143 -6520
rect -4097 -6521 -4083 -6475
rect -4158 -6534 -4083 -6521
rect -4268 -6810 -4222 -6753
rect -4025 -6579 -3979 -6417
rect -3866 -6417 -3865 -6399
rect -3866 -6445 -3819 -6417
rect -4158 -6810 -4083 -6796
rect -4268 -6811 -4083 -6810
rect -4268 -6856 -4143 -6811
rect -4268 -6915 -4222 -6856
rect -4158 -6857 -4143 -6856
rect -4097 -6857 -4083 -6811
rect -4158 -6870 -4083 -6857
rect -4268 -7146 -4222 -7089
rect -4025 -6915 -3979 -6753
rect -4158 -7146 -4083 -7132
rect -4268 -7147 -4083 -7146
rect -4268 -7192 -4143 -7147
rect -4268 -7251 -4222 -7192
rect -4158 -7193 -4143 -7192
rect -4097 -7193 -4083 -7147
rect -4158 -7206 -4083 -7193
rect -4268 -7436 -4222 -7425
rect -4025 -7251 -3979 -7089
rect -4025 -7482 -3979 -7425
rect -3865 -6579 -3819 -6445
rect -3865 -6915 -3819 -6753
rect -3865 -7251 -3819 -7089
rect -3865 -7436 -3819 -7425
rect -3705 -6243 -3659 -6232
rect -3546 -6243 -3499 -6186
rect -3705 -6579 -3659 -6417
rect -3705 -6915 -3659 -6753
rect -3705 -7251 -3659 -7089
rect -3705 -7482 -3659 -7425
rect -3545 -6579 -3499 -6417
rect -3545 -6915 -3499 -6753
rect -3545 -7251 -3499 -7089
rect -3545 -7436 -3499 -7425
rect -3385 -6243 -3339 -6232
rect -3226 -6243 -3179 -6186
rect -3385 -6579 -3339 -6417
rect -3385 -6915 -3339 -6753
rect -3385 -7251 -3339 -7089
rect -3385 -7482 -3339 -7425
rect -3225 -6579 -3179 -6417
rect -3225 -6915 -3179 -6753
rect -3225 -7251 -3179 -7089
rect -3225 -7436 -3179 -7425
rect -3065 -6243 -3019 -6232
rect -3065 -6579 -3019 -6417
rect -3065 -6915 -3019 -6753
rect -3065 -7251 -3019 -7089
rect -3065 -7482 -3019 -7425
rect -4025 -7530 -3019 -7482
rect -2429 -6236 -2383 -6225
rect -2429 -6572 -2383 -6410
rect -2429 -6908 -2383 -6746
rect -2429 -7244 -2383 -7082
rect -2429 -7572 -2383 -7418
rect -2269 -6236 -2223 -5959
rect -2119 -5962 -1925 -5959
rect -2269 -6572 -2223 -6410
rect -2269 -6908 -2223 -6746
rect -2269 -7244 -2223 -7082
rect -2269 -7429 -2223 -7418
rect -2025 -6236 -1979 -6225
rect -2025 -6572 -1979 -6410
rect -2025 -6908 -1979 -6746
rect -2025 -7244 -1979 -7082
rect -2025 -7572 -1979 -7418
rect -1865 -6236 -1819 -5828
rect -1622 -5318 -1576 -5260
rect -1622 -5654 -1576 -5492
rect -1622 -6022 -1576 -5828
rect -1462 -5318 -1416 -5307
rect -1462 -5654 -1416 -5492
rect -1462 -5886 -1416 -5828
rect -1302 -5318 -1256 -5260
rect -1302 -5654 -1256 -5492
rect -1302 -5839 -1256 -5828
rect -1142 -5318 -1096 -5307
rect -1142 -5654 -1096 -5492
rect -1142 -5886 -1096 -5828
rect -982 -5318 -936 -5260
rect -982 -5654 -936 -5492
rect -982 -5839 -936 -5828
rect -822 -5318 -776 -5307
rect -822 -5654 -776 -5492
rect -822 -5886 -776 -5828
rect -662 -5318 -616 -5260
rect -662 -5654 -616 -5492
rect -98 -5642 -40 -1695
rect 160 -1769 206 -1676
rect 160 -2005 206 -1843
rect 7 -2019 92 -2007
rect 7 -2075 24 -2019
rect 80 -2075 92 -2019
rect 7 -2129 92 -2075
rect 160 -2090 206 -2079
rect 320 -1769 366 -1758
rect 320 -2005 366 -1843
rect 7 -2185 24 -2129
rect 80 -2178 92 -2129
rect 189 -2172 266 -2157
rect 189 -2178 205 -2172
rect 80 -2185 205 -2178
rect 7 -2195 205 -2185
rect 17 -2221 205 -2195
rect 252 -2221 266 -2172
rect 17 -2223 266 -2221
rect 60 -2224 266 -2223
rect 189 -2234 266 -2224
rect 320 -2177 366 -2079
rect 480 -1769 526 -1676
rect 480 -2005 526 -1843
rect 480 -2090 526 -2079
rect 640 -1769 686 -1758
rect 640 -2005 686 -1843
rect 640 -2177 686 -2079
rect 800 -1769 846 -1676
rect 800 -2005 846 -1843
rect 800 -2090 846 -2079
rect 746 -2170 935 -2155
rect 746 -2177 756 -2170
rect 320 -2223 756 -2177
rect 160 -2354 206 -2343
rect 160 -2690 206 -2528
rect 160 -3002 206 -2864
rect 320 -2354 366 -2223
rect 320 -2690 366 -2528
rect 320 -2875 366 -2864
rect 480 -2354 526 -2343
rect 480 -2690 526 -2528
rect 480 -3002 526 -2864
rect 640 -2354 686 -2223
rect 746 -2224 756 -2223
rect 810 -2224 866 -2170
rect 920 -2177 935 -2170
rect 920 -2223 946 -2177
rect 920 -2224 935 -2223
rect 746 -2238 935 -2224
rect 640 -2690 686 -2528
rect 640 -2875 686 -2864
rect 800 -2354 846 -2343
rect 800 -2690 846 -2528
rect 800 -3002 846 -2864
rect 61 -3044 945 -3002
rect 61 -3104 124 -3044
rect 871 -3046 945 -3044
rect 922 -3102 945 -3046
rect 871 -3104 945 -3102
rect 61 -3146 945 -3104
rect 160 -3284 206 -3146
rect 160 -3620 206 -3458
rect 160 -3805 206 -3794
rect 320 -3284 366 -3273
rect 320 -3620 366 -3458
rect 189 -3924 266 -3914
rect 23 -3927 266 -3924
rect 23 -3970 205 -3927
rect 23 -4207 69 -3970
rect 189 -3976 205 -3970
rect 252 -3976 266 -3927
rect 189 -3991 266 -3976
rect 320 -3925 366 -3794
rect 480 -3284 526 -3146
rect 480 -3620 526 -3458
rect 480 -3805 526 -3794
rect 640 -3284 686 -3273
rect 640 -3620 686 -3458
rect 640 -3925 686 -3794
rect 800 -3284 846 -3146
rect 800 -3620 846 -3458
rect 800 -3805 846 -3794
rect 749 -3921 941 -3906
rect 749 -3925 765 -3921
rect 320 -3971 765 -3925
rect 160 -4069 206 -4058
rect 7 -4223 86 -4207
rect 7 -4277 19 -4223
rect 73 -4277 86 -4223
rect 7 -4333 86 -4277
rect 7 -4387 19 -4333
rect 73 -4387 86 -4333
rect 7 -4399 86 -4387
rect 160 -4305 206 -4143
rect 160 -4472 206 -4379
rect 320 -4069 366 -3971
rect 320 -4305 366 -4143
rect 320 -4390 366 -4379
rect 480 -4069 526 -4058
rect 480 -4305 526 -4143
rect 480 -4472 526 -4379
rect 640 -4069 686 -3971
rect 749 -3975 765 -3971
rect 819 -3975 875 -3921
rect 929 -3925 941 -3921
rect 929 -3971 946 -3925
rect 929 -3975 941 -3971
rect 749 -3987 941 -3975
rect 640 -4305 686 -4143
rect 640 -4390 686 -4379
rect 800 -4069 846 -4058
rect 800 -4305 846 -4143
rect 800 -4472 846 -4379
rect 61 -4517 945 -4472
rect 1008 -4500 1054 -1030
rect 1118 -2153 1165 -795
rect 1213 -860 1293 -848
rect 1213 -916 1225 -860
rect 1281 -916 1293 -860
rect 1213 -970 1293 -916
rect 1213 -1026 1225 -970
rect 1281 -1026 1293 -970
rect 1213 -1033 1293 -1026
rect 1225 -1898 1272 -1033
rect 1216 -1910 1287 -1898
rect 1216 -1964 1226 -1910
rect 1280 -1964 1287 -1910
rect 1216 -2020 1287 -1964
rect 1216 -2074 1226 -2020
rect 1280 -2074 1287 -2020
rect 1216 -2087 1287 -2074
rect 1104 -2165 1180 -2153
rect 1104 -2219 1115 -2165
rect 1169 -2219 1180 -2165
rect 1104 -2275 1180 -2219
rect 1104 -2329 1115 -2275
rect 1169 -2329 1180 -2275
rect 1104 -2340 1180 -2329
rect 1118 -4072 1165 -2340
rect 1103 -4085 1180 -4072
rect 1103 -4139 1115 -4085
rect 1169 -4139 1180 -4085
rect 1103 -4195 1180 -4139
rect 1103 -4249 1115 -4195
rect 1169 -4249 1180 -4195
rect 1103 -4263 1180 -4249
rect 1226 -4215 1272 -2087
rect 1344 -3796 1391 -670
rect 1469 -1389 1569 -5
rect 1930 -157 1976 -5
rect 3433 -6 3660 -5
rect 2333 -71 3339 -51
rect 2320 -83 3339 -71
rect 3743 -80 4749 -51
rect 2320 -86 3357 -83
rect 2320 -140 2330 -86
rect 2384 -88 3357 -86
rect 2384 -89 3288 -88
rect 2384 -99 2646 -89
rect 2384 -140 2396 -99
rect 1930 -493 1976 -331
rect 1930 -678 1976 -667
rect 2090 -157 2136 -146
rect 2320 -154 2396 -140
rect 2632 -145 2646 -99
rect 2702 -99 2966 -89
rect 2702 -145 2714 -99
rect 2090 -493 2136 -331
rect 1623 -721 1856 -718
rect 1623 -729 1912 -721
rect 1623 -783 1635 -729
rect 1689 -783 1745 -729
rect 1799 -734 2030 -729
rect 1799 -780 1850 -734
rect 1898 -742 2030 -734
rect 1898 -780 1957 -742
rect 1799 -783 1957 -780
rect 1623 -788 1957 -783
rect 2003 -788 2030 -742
rect 1623 -795 2030 -788
rect 1836 -801 2030 -795
rect 1751 -971 1807 -970
rect 1751 -990 1884 -971
rect 1751 -1024 1818 -990
rect 1807 -1046 1818 -1024
rect 1874 -1046 1884 -990
rect 1807 -1059 1884 -1046
rect 1930 -1075 1976 -1064
rect 1458 -1391 1584 -1389
rect 1458 -1447 1492 -1391
rect 1548 -1447 1584 -1391
rect 1458 -1501 1584 -1447
rect 1458 -1557 1492 -1501
rect 1548 -1557 1584 -1501
rect 1458 -1611 1584 -1557
rect 1458 -1667 1492 -1611
rect 1548 -1667 1584 -1611
rect 1458 -1674 1584 -1667
rect 1930 -1411 1976 -1249
rect 1930 -1747 1976 -1585
rect 1930 -2083 1976 -1921
rect 1930 -2411 1976 -2257
rect 2090 -1075 2136 -667
rect 2333 -157 2379 -154
rect 2333 -493 2379 -331
rect 2199 -991 2276 -979
rect 2199 -1045 2213 -991
rect 2267 -994 2276 -991
rect 2333 -994 2379 -667
rect 2493 -157 2539 -146
rect 2632 -147 2714 -145
rect 2953 -145 2966 -99
rect 3022 -99 3288 -89
rect 3022 -145 3035 -99
rect 3275 -144 3288 -99
rect 3344 -144 3357 -88
rect 3275 -145 3357 -144
rect 3718 -86 4749 -80
rect 3718 -88 4768 -86
rect 3718 -90 4378 -88
rect 2493 -493 2539 -331
rect 2493 -725 2539 -667
rect 2653 -157 2699 -147
rect 2653 -493 2699 -331
rect 2653 -678 2699 -667
rect 2813 -157 2859 -146
rect 2953 -147 3035 -145
rect 2813 -493 2859 -331
rect 2813 -725 2859 -667
rect 2973 -157 3019 -147
rect 2973 -493 3019 -331
rect 2973 -678 3019 -667
rect 3133 -157 3179 -146
rect 3133 -493 3179 -331
rect 3133 -725 3179 -667
rect 3293 -157 3339 -145
rect 3718 -146 3735 -90
rect 3791 -91 4378 -90
rect 3791 -99 4057 -91
rect 3791 -146 3804 -99
rect 3718 -151 3804 -146
rect 3293 -493 3339 -331
rect 3293 -678 3339 -667
rect 3743 -157 3789 -151
rect 3743 -493 3789 -331
rect 3743 -678 3789 -667
rect 3903 -157 3949 -146
rect 4041 -147 4057 -99
rect 4113 -99 4378 -91
rect 4113 -147 4127 -99
rect 4361 -144 4378 -99
rect 4434 -99 4768 -88
rect 4434 -144 4447 -99
rect 4361 -146 4447 -144
rect 4041 -151 4127 -147
rect 3903 -493 3949 -331
rect 2493 -834 3179 -725
rect 3083 -939 3179 -834
rect 2267 -1041 2379 -994
rect 2267 -1045 2276 -1041
rect 2199 -1057 2276 -1045
rect 2090 -1306 2136 -1249
rect 2333 -1075 2379 -1041
rect 2493 -941 3179 -939
rect 3903 -725 3949 -667
rect 4063 -157 4109 -151
rect 4063 -493 4109 -331
rect 4063 -678 4109 -667
rect 4223 -157 4269 -146
rect 4223 -493 4269 -331
rect 4223 -725 4269 -667
rect 4383 -157 4429 -146
rect 4383 -493 4429 -331
rect 4383 -678 4429 -667
rect 4543 -157 4589 -146
rect 4686 -153 4699 -99
rect 4753 -153 4768 -99
rect 4686 -157 4768 -153
rect 4686 -164 4703 -157
rect 4543 -493 4589 -331
rect 4543 -725 4589 -667
rect 3903 -834 4589 -725
rect 4749 -164 4768 -157
rect 4946 -157 4992 -146
rect 4703 -493 4749 -331
rect 3903 -939 3999 -834
rect 3903 -941 4589 -939
rect 2493 -1016 4589 -941
rect 2493 -1018 3179 -1016
rect 2493 -1075 2539 -1018
rect 2200 -1306 2275 -1292
rect 2090 -1307 2275 -1306
rect 2090 -1352 2215 -1307
rect 2090 -1411 2136 -1352
rect 2200 -1353 2215 -1352
rect 2261 -1353 2275 -1307
rect 2200 -1366 2275 -1353
rect 2090 -1642 2136 -1585
rect 2333 -1411 2379 -1249
rect 2492 -1249 2493 -1231
rect 2492 -1277 2539 -1249
rect 2200 -1642 2275 -1628
rect 2090 -1643 2275 -1642
rect 2090 -1688 2215 -1643
rect 2090 -1747 2136 -1688
rect 2200 -1689 2215 -1688
rect 2261 -1689 2275 -1643
rect 2200 -1702 2275 -1689
rect 2090 -1978 2136 -1921
rect 2333 -1747 2379 -1585
rect 2200 -1978 2275 -1964
rect 2090 -1979 2275 -1978
rect 2090 -2024 2215 -1979
rect 2090 -2083 2136 -2024
rect 2200 -2025 2215 -2024
rect 2261 -2025 2275 -1979
rect 2200 -2038 2275 -2025
rect 2090 -2268 2136 -2257
rect 2333 -2083 2379 -1921
rect 2333 -2314 2379 -2257
rect 2493 -1411 2539 -1277
rect 2493 -1747 2539 -1585
rect 2493 -2083 2539 -1921
rect 2493 -2268 2539 -2257
rect 2653 -1075 2699 -1064
rect 2812 -1075 2859 -1018
rect 2653 -1411 2699 -1249
rect 2653 -1747 2699 -1585
rect 2653 -2083 2699 -1921
rect 2653 -2314 2699 -2257
rect 2813 -1411 2859 -1249
rect 2813 -1747 2859 -1585
rect 2813 -2083 2859 -1921
rect 2813 -2268 2859 -2257
rect 2973 -1075 3019 -1064
rect 3132 -1075 3179 -1018
rect 2973 -1411 3019 -1249
rect 2973 -1747 3019 -1585
rect 2973 -2083 3019 -1921
rect 2973 -2314 3019 -2257
rect 3133 -1411 3179 -1249
rect 3133 -1747 3179 -1585
rect 3133 -2083 3179 -1921
rect 3133 -2268 3179 -2257
rect 3293 -1075 3339 -1064
rect 3293 -1411 3339 -1249
rect 3492 -1065 3604 -1016
rect 3903 -1018 4589 -1016
rect 3492 -1119 3512 -1065
rect 3566 -1119 3604 -1065
rect 3492 -1175 3604 -1119
rect 3492 -1229 3512 -1175
rect 3566 -1229 3604 -1175
rect 3492 -1254 3604 -1229
rect 3743 -1075 3789 -1064
rect 3293 -1747 3339 -1585
rect 3293 -2083 3339 -1921
rect 3293 -2314 3339 -2257
rect 2333 -2362 3339 -2314
rect 3743 -1411 3789 -1249
rect 3743 -1747 3789 -1585
rect 3743 -2083 3789 -1921
rect 3743 -2314 3789 -2257
rect 3903 -1075 3950 -1018
rect 4063 -1075 4109 -1064
rect 3903 -1411 3949 -1249
rect 3903 -1747 3949 -1585
rect 3903 -2083 3949 -1921
rect 3903 -2268 3949 -2257
rect 4063 -1411 4109 -1249
rect 4063 -1747 4109 -1585
rect 4063 -2083 4109 -1921
rect 4063 -2314 4109 -2257
rect 4223 -1075 4270 -1018
rect 4383 -1075 4429 -1064
rect 4223 -1411 4269 -1249
rect 4223 -1747 4269 -1585
rect 4223 -2083 4269 -1921
rect 4223 -2268 4269 -2257
rect 4383 -1411 4429 -1249
rect 4383 -1747 4429 -1585
rect 4383 -2083 4429 -1921
rect 4383 -2314 4429 -2257
rect 4543 -1075 4589 -1018
rect 4703 -994 4749 -667
rect 4946 -493 4992 -331
rect 4806 -991 4883 -979
rect 4806 -994 4815 -991
rect 4703 -1041 4815 -994
rect 4703 -1075 4749 -1041
rect 4806 -1045 4815 -1041
rect 4869 -1045 4883 -991
rect 4806 -1057 4883 -1045
rect 4589 -1249 4590 -1231
rect 4543 -1277 4590 -1249
rect 4543 -1411 4589 -1277
rect 4543 -1747 4589 -1585
rect 4543 -2083 4589 -1921
rect 4543 -2268 4589 -2257
rect 4703 -1411 4749 -1249
rect 4946 -1075 4992 -667
rect 5106 -157 5152 -5
rect 5511 -6 7412 -5
rect 5106 -493 5152 -331
rect 5610 -158 5656 -6
rect 6013 -100 7019 -52
rect 5106 -678 5152 -667
rect 5384 -460 5457 -444
rect 5384 -514 5394 -460
rect 5448 -514 5457 -460
rect 5384 -570 5457 -514
rect 5384 -624 5394 -570
rect 5448 -624 5457 -570
rect 5227 -721 5337 -720
rect 5170 -729 5337 -721
rect 5052 -733 5337 -729
rect 5052 -734 5269 -733
rect 5052 -742 5184 -734
rect 5052 -788 5079 -742
rect 5125 -780 5184 -742
rect 5232 -780 5269 -734
rect 5125 -788 5269 -780
rect 5052 -789 5269 -788
rect 5325 -789 5337 -733
rect 5384 -733 5457 -624
rect 5610 -494 5656 -332
rect 5610 -679 5656 -668
rect 5770 -158 5816 -147
rect 5770 -494 5816 -332
rect 5516 -730 5592 -722
rect 5516 -733 5710 -730
rect 5384 -735 5710 -733
rect 5384 -781 5530 -735
rect 5578 -743 5710 -735
rect 5578 -781 5637 -743
rect 5384 -782 5637 -781
rect 5052 -801 5337 -789
rect 5255 -843 5337 -801
rect 5516 -789 5637 -782
rect 5683 -789 5710 -743
rect 5516 -802 5710 -789
rect 5255 -899 5269 -843
rect 5325 -899 5337 -843
rect 5255 -914 5337 -899
rect 5275 -971 5331 -970
rect 5461 -971 5564 -970
rect 5198 -990 5331 -971
rect 5198 -1046 5208 -990
rect 5264 -1024 5331 -990
rect 5431 -991 5564 -971
rect 5264 -1046 5275 -1024
rect 5431 -1025 5498 -991
rect 5198 -1059 5275 -1046
rect 5461 -1047 5498 -1025
rect 5554 -1047 5564 -991
rect 4807 -1306 4882 -1292
rect 4946 -1306 4992 -1249
rect 4807 -1307 4992 -1306
rect 4807 -1353 4821 -1307
rect 4867 -1352 4992 -1307
rect 4867 -1353 4882 -1352
rect 4807 -1366 4882 -1353
rect 4703 -1747 4749 -1585
rect 4946 -1411 4992 -1352
rect 4807 -1642 4882 -1628
rect 4946 -1642 4992 -1585
rect 4807 -1643 4992 -1642
rect 4807 -1689 4821 -1643
rect 4867 -1688 4992 -1643
rect 4867 -1689 4882 -1688
rect 4807 -1702 4882 -1689
rect 4703 -2083 4749 -1921
rect 4946 -1747 4992 -1688
rect 4807 -1978 4882 -1964
rect 4946 -1978 4992 -1921
rect 4807 -1979 4992 -1978
rect 4807 -2025 4821 -1979
rect 4867 -2024 4992 -1979
rect 4867 -2025 4882 -2024
rect 4807 -2038 4882 -2025
rect 4703 -2314 4749 -2257
rect 4946 -2083 4992 -2024
rect 4946 -2268 4992 -2257
rect 5106 -1075 5152 -1064
rect 5106 -1411 5152 -1249
rect 5461 -1101 5564 -1047
rect 5461 -1157 5498 -1101
rect 5554 -1157 5564 -1101
rect 5461 -1254 5564 -1157
rect 5610 -1076 5656 -1065
rect 5106 -1747 5152 -1585
rect 5106 -2083 5152 -1921
rect 3743 -2362 4749 -2314
rect 5106 -2411 5152 -2257
rect 5610 -1412 5656 -1250
rect 5610 -1748 5656 -1586
rect 5610 -2084 5656 -1922
rect 1831 -2412 5251 -2411
rect 5610 -2412 5656 -2258
rect 5770 -1076 5816 -668
rect 6013 -158 6059 -100
rect 6013 -494 6059 -332
rect 5878 -992 5956 -980
rect 5878 -1046 5893 -992
rect 5947 -995 5956 -992
rect 6013 -995 6059 -668
rect 6173 -158 6219 -147
rect 6173 -494 6219 -332
rect 6173 -726 6219 -668
rect 6333 -158 6379 -100
rect 6333 -494 6379 -332
rect 6333 -679 6379 -668
rect 6493 -158 6539 -147
rect 6493 -494 6539 -332
rect 6493 -726 6539 -668
rect 6653 -158 6699 -100
rect 6653 -494 6699 -332
rect 6653 -679 6699 -668
rect 6813 -158 6859 -147
rect 6813 -494 6859 -332
rect 6813 -726 6859 -668
rect 6973 -158 7019 -100
rect 6973 -494 7019 -332
rect 6973 -679 7019 -668
rect 6173 -754 6859 -726
rect 7066 -747 7145 -731
rect 7066 -754 7078 -747
rect 6173 -801 7078 -754
rect 7132 -801 7145 -747
rect 6173 -835 7145 -801
rect 6661 -857 7145 -835
rect 6661 -911 7078 -857
rect 7132 -911 7145 -857
rect 6661 -940 7145 -911
rect 5947 -1042 6059 -995
rect 5947 -1046 5956 -1042
rect 5878 -1102 5956 -1046
rect 5878 -1156 5893 -1102
rect 5947 -1156 5956 -1102
rect 5878 -1175 5956 -1156
rect 6013 -1076 6059 -1042
rect 5770 -1307 5816 -1250
rect 6173 -942 7145 -940
rect 6173 -967 7198 -942
rect 6173 -1017 7078 -967
rect 6173 -1019 6859 -1017
rect 6173 -1076 6219 -1019
rect 5880 -1307 5955 -1293
rect 5770 -1308 5955 -1307
rect 5770 -1353 5895 -1308
rect 5770 -1412 5816 -1353
rect 5880 -1354 5895 -1353
rect 5941 -1354 5955 -1308
rect 5880 -1367 5955 -1354
rect 5770 -1643 5816 -1586
rect 6013 -1412 6059 -1250
rect 6172 -1250 6173 -1232
rect 6172 -1278 6219 -1250
rect 5880 -1643 5955 -1629
rect 5770 -1644 5955 -1643
rect 5770 -1689 5895 -1644
rect 5770 -1748 5816 -1689
rect 5880 -1690 5895 -1689
rect 5941 -1690 5955 -1644
rect 5880 -1703 5955 -1690
rect 5770 -1979 5816 -1922
rect 6013 -1748 6059 -1586
rect 5880 -1979 5955 -1965
rect 5770 -1980 5955 -1979
rect 5770 -2025 5895 -1980
rect 5770 -2084 5816 -2025
rect 5880 -2026 5895 -2025
rect 5941 -2026 5955 -1980
rect 5880 -2039 5955 -2026
rect 5770 -2269 5816 -2258
rect 6013 -2084 6059 -1922
rect 6013 -2315 6059 -2258
rect 6173 -1412 6219 -1278
rect 6173 -1748 6219 -1586
rect 6173 -2084 6219 -1922
rect 6173 -2269 6219 -2258
rect 6333 -1076 6379 -1065
rect 6492 -1076 6539 -1019
rect 6333 -1412 6379 -1250
rect 6333 -1748 6379 -1586
rect 6333 -2084 6379 -1922
rect 6333 -2315 6379 -2258
rect 6493 -1412 6539 -1250
rect 6493 -1748 6539 -1586
rect 6493 -2084 6539 -1922
rect 6493 -2269 6539 -2258
rect 6653 -1076 6699 -1065
rect 6812 -1076 6859 -1019
rect 7066 -1021 7078 -1017
rect 7132 -1017 7198 -967
rect 7132 -1021 7146 -1017
rect 7066 -1034 7146 -1021
rect 6653 -1412 6699 -1250
rect 6653 -1748 6699 -1586
rect 6653 -2084 6699 -1922
rect 6653 -2315 6699 -2258
rect 6813 -1412 6859 -1250
rect 6813 -1748 6859 -1586
rect 6813 -2084 6859 -1922
rect 6813 -2269 6859 -2258
rect 6973 -1076 7019 -1065
rect 6973 -1412 7019 -1250
rect 6973 -1748 7019 -1586
rect 6973 -2084 7019 -1922
rect 6973 -2315 7019 -2258
rect 6013 -2363 7019 -2315
rect 1831 -2450 7118 -2412
rect 1682 -2471 7118 -2450
rect 1682 -2525 1891 -2471
rect 2052 -2525 2112 -2471
rect 2273 -2525 2333 -2471
rect 2494 -2525 2554 -2471
rect 2715 -2525 2775 -2471
rect 2936 -2525 2996 -2471
rect 3157 -2525 3217 -2471
rect 3378 -2525 3704 -2471
rect 3865 -2525 3925 -2471
rect 4086 -2525 4146 -2471
rect 4307 -2525 4367 -2471
rect 4528 -2525 4588 -2471
rect 4749 -2525 4809 -2471
rect 4970 -2525 5030 -2471
rect 5191 -2472 7118 -2471
rect 5191 -2525 5571 -2472
rect 1682 -2526 5571 -2525
rect 5732 -2526 5792 -2472
rect 5953 -2526 6013 -2472
rect 6174 -2526 6234 -2472
rect 6395 -2526 6455 -2472
rect 6616 -2473 6676 -2472
rect 6837 -2473 6897 -2472
rect 6616 -2525 6627 -2473
rect 6837 -2525 6867 -2473
rect 6616 -2526 6676 -2525
rect 6837 -2526 6897 -2525
rect 7058 -2526 7118 -2472
rect 1682 -2550 7118 -2526
rect 1682 -2850 1782 -2550
rect 1831 -2585 7118 -2550
rect 1930 -2739 1976 -2585
rect 3416 -2586 3682 -2585
rect 2333 -2682 3339 -2634
rect 1666 -2861 1794 -2850
rect 1666 -2917 1702 -2861
rect 1758 -2917 1794 -2861
rect 1666 -2971 1794 -2917
rect 1666 -3027 1702 -2971
rect 1758 -3027 1794 -2971
rect 1666 -3081 1794 -3027
rect 1666 -3137 1702 -3081
rect 1758 -3137 1794 -3081
rect 1666 -3143 1794 -3137
rect 1930 -3075 1976 -2913
rect 1930 -3411 1976 -3249
rect 1930 -3747 1976 -3585
rect 1323 -3808 1405 -3796
rect 1323 -3865 1333 -3808
rect 1390 -3865 1405 -3808
rect 1323 -3918 1405 -3865
rect 1323 -3975 1333 -3918
rect 1390 -3975 1405 -3918
rect 1930 -3932 1976 -3921
rect 2090 -2739 2136 -2728
rect 2090 -2972 2136 -2913
rect 2333 -2739 2379 -2682
rect 2200 -2971 2275 -2958
rect 2200 -2972 2215 -2971
rect 2090 -3017 2215 -2972
rect 2261 -3017 2275 -2971
rect 2090 -3018 2275 -3017
rect 2090 -3075 2136 -3018
rect 2200 -3032 2275 -3018
rect 2090 -3308 2136 -3249
rect 2333 -3075 2379 -2913
rect 2200 -3307 2275 -3294
rect 2200 -3308 2215 -3307
rect 2090 -3353 2215 -3308
rect 2261 -3353 2275 -3307
rect 2090 -3354 2275 -3353
rect 2090 -3411 2136 -3354
rect 2200 -3368 2275 -3354
rect 2090 -3644 2136 -3585
rect 2333 -3411 2379 -3249
rect 2200 -3643 2275 -3630
rect 2200 -3644 2215 -3643
rect 2090 -3689 2215 -3644
rect 2261 -3689 2275 -3643
rect 2090 -3690 2275 -3689
rect 2090 -3747 2136 -3690
rect 2200 -3704 2275 -3690
rect 1807 -3950 1884 -3937
rect 1807 -3972 1818 -3950
rect 1323 -3989 1405 -3975
rect 1751 -4006 1818 -3972
rect 1874 -4006 1884 -3950
rect 1751 -4025 1884 -4006
rect 1751 -4026 1807 -4025
rect 1836 -4208 2030 -4195
rect 1836 -4215 1957 -4208
rect 1226 -4216 1957 -4215
rect 1226 -4262 1850 -4216
rect 1898 -4254 1957 -4216
rect 2003 -4254 2030 -4208
rect 1898 -4262 2030 -4254
rect 1226 -4264 2030 -4262
rect 1836 -4267 2030 -4264
rect 1836 -4275 1912 -4267
rect 1930 -4329 1976 -4318
rect 61 -4572 115 -4517
rect 879 -4572 945 -4517
rect 61 -4611 945 -4572
rect 991 -4512 1180 -4500
rect 991 -4566 1004 -4512
rect 1058 -4566 1114 -4512
rect 1168 -4566 1180 -4512
rect 991 -4579 1180 -4566
rect 311 -4991 405 -4611
rect 1930 -4665 1976 -4503
rect 1674 -4991 1837 -4990
rect 1930 -4991 1976 -4839
rect 2090 -4329 2136 -3921
rect 2333 -3747 2379 -3585
rect 2493 -2739 2539 -2728
rect 2493 -3075 2539 -2913
rect 2493 -3411 2539 -3249
rect 2493 -3719 2539 -3585
rect 2492 -3747 2539 -3719
rect 2492 -3765 2493 -3747
rect 2199 -3951 2276 -3939
rect 2199 -4005 2213 -3951
rect 2267 -3955 2276 -3951
rect 2333 -3955 2379 -3921
rect 2267 -4002 2379 -3955
rect 2267 -4005 2276 -4002
rect 2199 -4017 2276 -4005
rect 2090 -4665 2136 -4503
rect 2333 -4329 2379 -4002
rect 2493 -3978 2539 -3921
rect 2653 -2739 2699 -2682
rect 2653 -3075 2699 -2913
rect 2653 -3411 2699 -3249
rect 2653 -3747 2699 -3585
rect 2813 -2739 2859 -2728
rect 2813 -3075 2859 -2913
rect 2813 -3411 2859 -3249
rect 2813 -3747 2859 -3585
rect 2653 -3932 2699 -3921
rect 2812 -3978 2859 -3921
rect 2973 -2739 3019 -2682
rect 2973 -3075 3019 -2913
rect 2973 -3411 3019 -3249
rect 2973 -3747 3019 -3585
rect 3133 -2739 3179 -2728
rect 3133 -3075 3179 -2913
rect 3133 -3411 3179 -3249
rect 3133 -3747 3179 -3585
rect 2973 -3932 3019 -3921
rect 3132 -3978 3179 -3921
rect 3293 -2739 3339 -2682
rect 3293 -3075 3339 -2913
rect 3293 -3411 3339 -3249
rect 3293 -3747 3339 -3585
rect 3743 -2682 4749 -2634
rect 3743 -2739 3789 -2682
rect 3743 -3075 3789 -2913
rect 3743 -3411 3789 -3249
rect 3743 -3747 3789 -3585
rect 3293 -3932 3339 -3921
rect 3520 -3823 3602 -3810
rect 3520 -3881 3533 -3823
rect 3591 -3881 3602 -3823
rect 2493 -3980 3179 -3978
rect 3520 -3933 3602 -3881
rect 3743 -3932 3789 -3921
rect 3903 -2739 3949 -2728
rect 3903 -3075 3949 -2913
rect 3903 -3411 3949 -3249
rect 3903 -3747 3949 -3585
rect 4063 -2739 4109 -2682
rect 4063 -3075 4109 -2913
rect 4063 -3411 4109 -3249
rect 4063 -3747 4109 -3585
rect 3520 -3980 3533 -3933
rect 2493 -3991 3533 -3980
rect 3591 -3980 3602 -3933
rect 3903 -3978 3950 -3921
rect 4063 -3932 4109 -3921
rect 4223 -2739 4269 -2728
rect 4223 -3075 4269 -2913
rect 4223 -3411 4269 -3249
rect 4223 -3747 4269 -3585
rect 4383 -2739 4429 -2682
rect 4383 -3075 4429 -2913
rect 4383 -3411 4429 -3249
rect 4383 -3747 4429 -3585
rect 4223 -3978 4270 -3921
rect 4383 -3932 4429 -3921
rect 4543 -2739 4589 -2728
rect 4543 -3075 4589 -2913
rect 4543 -3411 4589 -3249
rect 4543 -3719 4589 -3585
rect 4703 -2739 4749 -2682
rect 4703 -3075 4749 -2913
rect 4946 -2739 4992 -2728
rect 4807 -2971 4882 -2958
rect 4807 -3017 4821 -2971
rect 4867 -2972 4882 -2971
rect 4946 -2972 4992 -2913
rect 4867 -3017 4992 -2972
rect 4807 -3018 4992 -3017
rect 4807 -3032 4882 -3018
rect 4703 -3411 4749 -3249
rect 4946 -3075 4992 -3018
rect 4807 -3307 4882 -3294
rect 4807 -3353 4821 -3307
rect 4867 -3308 4882 -3307
rect 4946 -3308 4992 -3249
rect 4867 -3353 4992 -3308
rect 4807 -3354 4992 -3353
rect 4807 -3368 4882 -3354
rect 4543 -3747 4590 -3719
rect 4589 -3765 4590 -3747
rect 4703 -3747 4749 -3585
rect 4946 -3411 4992 -3354
rect 4807 -3643 4882 -3630
rect 4807 -3689 4821 -3643
rect 4867 -3644 4882 -3643
rect 4946 -3644 4992 -3585
rect 4867 -3689 4992 -3644
rect 4807 -3690 4992 -3689
rect 4807 -3704 4882 -3690
rect 4543 -3978 4589 -3921
rect 3903 -3980 4589 -3978
rect 3591 -3991 4589 -3980
rect 2493 -4055 4589 -3991
rect 2493 -4057 3179 -4055
rect 3083 -4162 3179 -4057
rect 2333 -4665 2379 -4503
rect 2090 -4850 2136 -4839
rect 2327 -4839 2333 -4833
rect 2493 -4271 3179 -4162
rect 2493 -4329 2539 -4271
rect 2493 -4665 2539 -4503
rect 2379 -4837 2403 -4833
rect 2327 -4891 2337 -4839
rect 2391 -4891 2403 -4837
rect 2653 -4329 2699 -4318
rect 2653 -4665 2699 -4503
rect 2493 -4850 2539 -4839
rect 2625 -4832 2653 -4822
rect 2813 -4329 2859 -4271
rect 2813 -4665 2859 -4503
rect 2699 -4832 2717 -4822
rect 2327 -4897 2403 -4891
rect 2625 -4888 2645 -4832
rect 2701 -4888 2717 -4832
rect 2973 -4329 3019 -4318
rect 2973 -4665 3019 -4503
rect 2813 -4850 2859 -4839
rect 2952 -4839 2973 -4835
rect 3133 -4329 3179 -4271
rect 3903 -4057 4589 -4055
rect 4703 -3955 4749 -3921
rect 4946 -3747 4992 -3690
rect 4806 -3951 4883 -3939
rect 4806 -3955 4815 -3951
rect 4703 -4002 4815 -3955
rect 3903 -4162 3999 -4057
rect 3903 -4271 4589 -4162
rect 3133 -4665 3179 -4503
rect 3019 -4839 3037 -4835
rect 2952 -4845 3037 -4839
rect 2625 -4897 2717 -4888
rect 2952 -4897 2966 -4845
rect 2327 -4901 2966 -4897
rect 3022 -4897 3037 -4845
rect 3293 -4329 3339 -4318
rect 3293 -4665 3339 -4503
rect 3133 -4850 3179 -4839
rect 3271 -4839 3293 -4837
rect 3743 -4329 3789 -4318
rect 3743 -4665 3789 -4503
rect 3339 -4839 3349 -4837
rect 3271 -4848 3349 -4839
rect 3271 -4897 3283 -4848
rect 3022 -4901 3283 -4897
rect 2327 -4904 3283 -4901
rect 3339 -4904 3349 -4848
rect 2327 -4906 3349 -4904
rect 2333 -4916 3349 -4906
rect 3732 -4839 3743 -4834
rect 3903 -4329 3949 -4271
rect 3903 -4665 3949 -4503
rect 3789 -4839 3813 -4834
rect 3732 -4848 3813 -4839
rect 3732 -4904 3745 -4848
rect 3801 -4897 3813 -4848
rect 4063 -4329 4109 -4318
rect 4063 -4665 4109 -4503
rect 3903 -4850 3949 -4839
rect 4044 -4839 4063 -4828
rect 4223 -4329 4269 -4271
rect 4223 -4665 4269 -4503
rect 4109 -4839 4125 -4828
rect 4044 -4846 4125 -4839
rect 4044 -4897 4057 -4846
rect 3801 -4902 4057 -4897
rect 4113 -4897 4125 -4846
rect 4383 -4329 4429 -4318
rect 4383 -4665 4429 -4503
rect 4223 -4850 4269 -4839
rect 4364 -4839 4383 -4830
rect 4543 -4329 4589 -4271
rect 4543 -4665 4589 -4503
rect 4429 -4839 4445 -4830
rect 4364 -4843 4445 -4839
rect 4364 -4897 4377 -4843
rect 4113 -4899 4377 -4897
rect 4433 -4897 4445 -4843
rect 4703 -4329 4749 -4002
rect 4806 -4005 4815 -4002
rect 4869 -4005 4883 -3951
rect 4806 -4017 4883 -4005
rect 4703 -4665 4749 -4503
rect 4543 -4850 4589 -4839
rect 4683 -4839 4703 -4828
rect 4946 -4329 4992 -3921
rect 5106 -2739 5152 -2585
rect 5511 -2586 7118 -2585
rect 5106 -3075 5152 -2913
rect 5106 -3411 5152 -3249
rect 5106 -3747 5152 -3585
rect 5610 -2740 5656 -2586
rect 6013 -2683 7019 -2635
rect 5610 -3076 5656 -2914
rect 5610 -3412 5656 -3250
rect 5610 -3748 5656 -3586
rect 5106 -3932 5152 -3921
rect 5487 -3841 5564 -3822
rect 5487 -3897 5498 -3841
rect 5554 -3897 5564 -3841
rect 5198 -3950 5275 -3937
rect 5198 -4006 5208 -3950
rect 5264 -3972 5275 -3950
rect 5487 -3951 5564 -3897
rect 5610 -3933 5656 -3922
rect 5770 -2740 5816 -2729
rect 5770 -2973 5816 -2914
rect 6013 -2740 6059 -2683
rect 5880 -2972 5955 -2959
rect 5880 -2973 5895 -2972
rect 5770 -3018 5895 -2973
rect 5941 -3018 5955 -2972
rect 5770 -3019 5955 -3018
rect 5770 -3076 5816 -3019
rect 5880 -3033 5955 -3019
rect 5770 -3309 5816 -3250
rect 6013 -3076 6059 -2914
rect 5880 -3308 5955 -3295
rect 5880 -3309 5895 -3308
rect 5770 -3354 5895 -3309
rect 5941 -3354 5955 -3308
rect 5770 -3355 5955 -3354
rect 5770 -3412 5816 -3355
rect 5880 -3369 5955 -3355
rect 5770 -3645 5816 -3586
rect 6013 -3412 6059 -3250
rect 5880 -3644 5955 -3631
rect 5880 -3645 5895 -3644
rect 5770 -3690 5895 -3645
rect 5941 -3690 5955 -3644
rect 5770 -3691 5955 -3690
rect 5770 -3748 5816 -3691
rect 5880 -3705 5955 -3691
rect 6013 -3748 6059 -3586
rect 6173 -2740 6219 -2729
rect 6173 -3076 6219 -2914
rect 6173 -3412 6219 -3250
rect 6173 -3720 6219 -3586
rect 5264 -4006 5331 -3972
rect 5487 -3973 5498 -3951
rect 5198 -4025 5331 -4006
rect 5275 -4026 5331 -4025
rect 5431 -4007 5498 -3973
rect 5554 -4007 5564 -3951
rect 5431 -4027 5564 -4007
rect 5244 -4099 5322 -4083
rect 5244 -4155 5253 -4099
rect 5309 -4155 5322 -4099
rect 5244 -4195 5322 -4155
rect 5052 -4202 5322 -4195
rect 5052 -4208 5324 -4202
rect 5052 -4254 5079 -4208
rect 5125 -4209 5324 -4208
rect 5125 -4216 5253 -4209
rect 5125 -4254 5184 -4216
rect 5052 -4262 5184 -4254
rect 5232 -4262 5253 -4216
rect 5052 -4265 5253 -4262
rect 5309 -4215 5324 -4209
rect 5516 -4209 5710 -4196
rect 5309 -4264 5331 -4215
rect 5421 -4216 5470 -4215
rect 5516 -4216 5637 -4209
rect 5421 -4217 5637 -4216
rect 5421 -4263 5530 -4217
rect 5578 -4255 5637 -4217
rect 5683 -4255 5710 -4209
rect 5578 -4263 5710 -4255
rect 5309 -4265 5324 -4264
rect 5052 -4267 5324 -4265
rect 5170 -4275 5324 -4267
rect 5243 -4276 5324 -4275
rect 5421 -4265 5710 -4263
rect 4946 -4665 4992 -4503
rect 4749 -4839 4771 -4828
rect 4683 -4843 4771 -4839
rect 4683 -4897 4699 -4843
rect 4753 -4897 4771 -4843
rect 4946 -4850 4992 -4839
rect 5106 -4329 5152 -4318
rect 5421 -4329 5470 -4265
rect 5516 -4268 5710 -4265
rect 5516 -4276 5592 -4268
rect 5106 -4665 5152 -4503
rect 5412 -4343 5484 -4329
rect 5412 -4397 5419 -4343
rect 5473 -4397 5484 -4343
rect 5412 -4453 5484 -4397
rect 5412 -4507 5419 -4453
rect 5473 -4507 5484 -4453
rect 5412 -4522 5484 -4507
rect 5610 -4330 5656 -4319
rect 4433 -4899 4771 -4897
rect 4113 -4902 4771 -4899
rect 3801 -4904 4771 -4902
rect 3732 -4909 4771 -4904
rect 2333 -4945 3339 -4916
rect 3732 -4920 4749 -4909
rect 3743 -4945 4749 -4920
rect 5106 -4991 5152 -4839
rect 5610 -4666 5656 -4504
rect 71 -4992 5251 -4991
rect 5610 -4992 5656 -4840
rect 5770 -4330 5816 -3922
rect 5876 -3842 5956 -3836
rect 5876 -3896 5889 -3842
rect 5943 -3896 5956 -3842
rect 5876 -3952 5956 -3896
rect 5876 -4006 5893 -3952
rect 5947 -3956 5956 -3952
rect 6172 -3748 6219 -3720
rect 6172 -3766 6173 -3748
rect 6013 -3956 6059 -3922
rect 5947 -4003 6059 -3956
rect 5947 -4006 5956 -4003
rect 5876 -4018 5956 -4006
rect 5770 -4666 5816 -4504
rect 5770 -4851 5816 -4840
rect 6013 -4330 6059 -4003
rect 6173 -3979 6219 -3922
rect 6333 -2740 6379 -2683
rect 6333 -3076 6379 -2914
rect 6333 -3412 6379 -3250
rect 6333 -3748 6379 -3586
rect 6493 -2740 6539 -2729
rect 6493 -3076 6539 -2914
rect 6493 -3412 6539 -3250
rect 6493 -3748 6539 -3586
rect 6333 -3933 6379 -3922
rect 6492 -3979 6539 -3922
rect 6653 -2740 6699 -2683
rect 6653 -3076 6699 -2914
rect 6653 -3412 6699 -3250
rect 6653 -3748 6699 -3586
rect 6813 -2740 6859 -2729
rect 6813 -3076 6859 -2914
rect 6813 -3412 6859 -3250
rect 6813 -3748 6859 -3586
rect 6653 -3933 6699 -3922
rect 6812 -3979 6859 -3922
rect 6973 -2740 7019 -2683
rect 6973 -3076 7019 -2914
rect 6973 -3412 7019 -3250
rect 6973 -3748 7019 -3586
rect 6973 -3933 7019 -3922
rect 6173 -3981 6859 -3979
rect 7084 -3977 7162 -3964
rect 7084 -3981 7096 -3977
rect 6173 -4031 7096 -3981
rect 7150 -3981 7162 -3977
rect 7150 -4031 7198 -3981
rect 6173 -4056 7198 -4031
rect 6173 -4058 7162 -4056
rect 6675 -4087 7162 -4058
rect 6675 -4141 7096 -4087
rect 7150 -4141 7162 -4087
rect 6675 -4163 7162 -4141
rect 6013 -4666 6059 -4504
rect 6013 -4898 6059 -4840
rect 6173 -4197 7162 -4163
rect 6173 -4231 7096 -4197
rect 6173 -4272 6859 -4231
rect 7084 -4251 7096 -4231
rect 7150 -4251 7162 -4197
rect 7084 -4268 7162 -4251
rect 6173 -4330 6219 -4272
rect 6173 -4666 6219 -4504
rect 6173 -4851 6219 -4840
rect 6333 -4330 6379 -4319
rect 6333 -4666 6379 -4504
rect 6333 -4898 6379 -4840
rect 6493 -4330 6539 -4272
rect 6493 -4666 6539 -4504
rect 6493 -4851 6539 -4840
rect 6653 -4330 6699 -4319
rect 6653 -4666 6699 -4504
rect 6653 -4898 6699 -4840
rect 6813 -4330 6859 -4272
rect 6813 -4666 6859 -4504
rect 6813 -4851 6859 -4840
rect 6973 -4330 7019 -4319
rect 6973 -4666 7019 -4504
rect 6973 -4898 7019 -4840
rect 6013 -4946 7019 -4898
rect 7245 -4992 7412 -6
rect 71 -5050 7412 -4992
rect 71 -5106 86 -5050
rect 142 -5051 196 -5050
rect 252 -5051 306 -5050
rect 362 -5051 416 -5050
rect 472 -5051 526 -5050
rect 582 -5051 636 -5050
rect 692 -5051 746 -5050
rect 802 -5051 7412 -5050
rect 292 -5105 306 -5051
rect 513 -5105 526 -5051
rect 734 -5105 746 -5051
rect 955 -5105 1015 -5051
rect 1176 -5105 1236 -5051
rect 1397 -5105 1457 -5051
rect 1618 -5105 1891 -5051
rect 2052 -5105 2112 -5051
rect 2273 -5105 2333 -5051
rect 2494 -5105 2554 -5051
rect 2715 -5105 2775 -5051
rect 2936 -5105 2996 -5051
rect 3157 -5105 3217 -5051
rect 3378 -5105 3704 -5051
rect 3865 -5105 3925 -5051
rect 4086 -5105 4146 -5051
rect 4307 -5105 4367 -5051
rect 4528 -5105 4588 -5051
rect 4749 -5105 4809 -5051
rect 4970 -5105 5030 -5051
rect 5191 -5052 7412 -5051
rect 5191 -5105 5571 -5052
rect 142 -5106 196 -5105
rect 252 -5106 306 -5105
rect 362 -5106 416 -5105
rect 472 -5106 526 -5105
rect 582 -5106 636 -5105
rect 692 -5106 746 -5105
rect 802 -5106 5571 -5105
rect 5732 -5106 5792 -5052
rect 5953 -5106 6013 -5052
rect 6174 -5106 6234 -5052
rect 6395 -5106 6455 -5052
rect 6616 -5106 6676 -5052
rect 6837 -5106 6897 -5052
rect 7058 -5106 7412 -5052
rect 71 -5164 7412 -5106
rect 71 -5165 3438 -5164
rect 3644 -5165 7412 -5164
rect 170 -5317 216 -5165
rect 573 -5259 1579 -5211
rect -97 -5646 -16 -5642
rect -97 -5703 -85 -5646
rect -28 -5703 -16 -5646
rect -97 -5756 -16 -5703
rect -97 -5813 -85 -5756
rect -28 -5813 -16 -5756
rect -97 -5823 -16 -5813
rect 170 -5653 216 -5491
rect -662 -5839 -616 -5828
rect -1462 -5995 -776 -5886
rect -86 -5892 -40 -5823
rect 170 -5838 216 -5827
rect 330 -5317 376 -5306
rect 330 -5653 376 -5491
rect 76 -5889 152 -5881
rect 76 -5892 270 -5889
rect -86 -5894 270 -5892
rect -86 -5940 90 -5894
rect 138 -5902 270 -5894
rect 138 -5940 197 -5902
rect -86 -5941 197 -5940
rect 76 -5948 197 -5941
rect 243 -5948 270 -5902
rect 76 -5961 270 -5948
rect -1756 -6035 -1576 -6022
rect -1756 -6094 -1746 -6035
rect -1687 -6094 -1576 -6035
rect -1756 -6152 -1576 -6094
rect -872 -6100 -776 -5995
rect -1756 -6206 -1742 -6152
rect -1688 -6202 -1576 -6152
rect -1688 -6206 -1679 -6202
rect -1756 -6218 -1679 -6206
rect -1865 -6467 -1819 -6410
rect -1622 -6236 -1576 -6202
rect -1462 -6102 -776 -6100
rect 47 -6041 124 -6027
rect 47 -6097 57 -6041
rect 113 -6097 124 -6041
rect -1462 -6110 -437 -6102
rect -1462 -6166 -633 -6110
rect -577 -6166 -508 -6110
rect -452 -6166 -437 -6110
rect 47 -6130 124 -6097
rect -1462 -6177 -437 -6166
rect -9 -6150 124 -6130
rect -1462 -6179 -776 -6177
rect -1462 -6236 -1416 -6179
rect -1755 -6467 -1680 -6453
rect -1865 -6468 -1680 -6467
rect -1865 -6513 -1740 -6468
rect -1865 -6572 -1819 -6513
rect -1755 -6514 -1740 -6513
rect -1694 -6514 -1680 -6468
rect -1755 -6527 -1680 -6514
rect -1865 -6803 -1819 -6746
rect -1622 -6572 -1576 -6410
rect -1463 -6410 -1462 -6392
rect -1463 -6438 -1416 -6410
rect -1755 -6803 -1680 -6789
rect -1865 -6804 -1680 -6803
rect -1865 -6849 -1740 -6804
rect -1865 -6908 -1819 -6849
rect -1755 -6850 -1740 -6849
rect -1694 -6850 -1680 -6804
rect -1755 -6863 -1680 -6850
rect -1865 -7139 -1819 -7082
rect -1622 -6908 -1576 -6746
rect -1755 -7139 -1680 -7125
rect -1865 -7140 -1680 -7139
rect -1865 -7185 -1740 -7140
rect -1865 -7244 -1819 -7185
rect -1755 -7186 -1740 -7185
rect -1694 -7186 -1680 -7140
rect -1755 -7199 -1680 -7186
rect -1865 -7429 -1819 -7418
rect -1622 -7244 -1576 -7082
rect -1622 -7475 -1576 -7418
rect -1462 -6572 -1416 -6438
rect -1462 -6908 -1416 -6746
rect -1462 -7244 -1416 -7082
rect -1462 -7429 -1416 -7418
rect -1302 -6236 -1256 -6225
rect -1143 -6236 -1096 -6179
rect -1302 -6572 -1256 -6410
rect -1302 -6908 -1256 -6746
rect -1302 -7244 -1256 -7082
rect -1302 -7475 -1256 -7418
rect -1142 -6572 -1096 -6410
rect -1142 -6908 -1096 -6746
rect -1142 -7244 -1096 -7082
rect -1142 -7429 -1096 -7418
rect -982 -6236 -936 -6225
rect -823 -6236 -776 -6179
rect -9 -6184 58 -6150
rect 47 -6206 58 -6184
rect 114 -6206 124 -6150
rect 47 -6220 124 -6206
rect -982 -6572 -936 -6410
rect -982 -6908 -936 -6746
rect -982 -7244 -936 -7082
rect -982 -7475 -936 -7418
rect -822 -6572 -776 -6410
rect -822 -6908 -776 -6746
rect -822 -7244 -776 -7082
rect -822 -7429 -776 -7418
rect -662 -6236 -616 -6225
rect -662 -6572 -616 -6410
rect -662 -6908 -616 -6746
rect -662 -7244 -616 -7082
rect -662 -7475 -616 -7418
rect -1622 -7523 -616 -7475
rect 170 -6235 216 -6224
rect 170 -6571 216 -6409
rect 170 -6907 216 -6745
rect 170 -7243 216 -7081
rect 170 -7571 216 -7417
rect 330 -6235 376 -5827
rect 573 -5317 619 -5259
rect 573 -5653 619 -5491
rect 439 -6040 516 -6028
rect 439 -6096 448 -6040
rect 504 -6096 516 -6040
rect 439 -6151 516 -6096
rect 439 -6205 453 -6151
rect 507 -6154 516 -6151
rect 573 -6154 619 -5827
rect 733 -5317 779 -5306
rect 733 -5653 779 -5491
rect 733 -5885 779 -5827
rect 893 -5317 939 -5259
rect 893 -5653 939 -5491
rect 893 -5838 939 -5827
rect 1053 -5317 1099 -5306
rect 1053 -5653 1099 -5491
rect 1053 -5885 1099 -5827
rect 1213 -5317 1259 -5259
rect 1213 -5653 1259 -5491
rect 1213 -5838 1259 -5827
rect 1373 -5317 1419 -5306
rect 1373 -5653 1419 -5491
rect 1373 -5885 1419 -5827
rect 1533 -5317 1579 -5259
rect 1930 -5259 2936 -5211
rect 1930 -5317 1976 -5259
rect 1533 -5653 1579 -5491
rect 1533 -5838 1579 -5827
rect 1715 -5337 1795 -5324
rect 1715 -5392 1728 -5337
rect 1783 -5392 1795 -5337
rect 1715 -5447 1795 -5392
rect 1715 -5502 1728 -5447
rect 1783 -5502 1795 -5447
rect 733 -5994 1419 -5885
rect 1323 -6099 1419 -5994
rect 507 -6201 619 -6154
rect 507 -6205 516 -6201
rect 439 -6217 516 -6205
rect 330 -6466 376 -6409
rect 573 -6235 619 -6201
rect 733 -6101 1419 -6099
rect 1715 -6101 1795 -5502
rect 1930 -5653 1976 -5491
rect 1930 -5838 1976 -5827
rect 2090 -5317 2136 -5306
rect 2090 -5653 2136 -5491
rect 2090 -5885 2136 -5827
rect 2250 -5317 2296 -5259
rect 2250 -5653 2296 -5491
rect 2250 -5838 2296 -5827
rect 2410 -5317 2456 -5306
rect 2410 -5653 2456 -5491
rect 2410 -5885 2456 -5827
rect 2570 -5317 2616 -5259
rect 2570 -5653 2616 -5491
rect 2570 -5838 2616 -5827
rect 2730 -5317 2776 -5306
rect 2730 -5653 2776 -5491
rect 2730 -5885 2776 -5827
rect 2090 -5994 2776 -5885
rect 2890 -5317 2936 -5259
rect 2890 -5653 2936 -5491
rect 2090 -6099 2186 -5994
rect 2090 -6101 2776 -6099
rect 733 -6176 2776 -6101
rect 733 -6178 1419 -6176
rect 1715 -6177 1795 -6176
rect 733 -6235 779 -6178
rect 440 -6466 515 -6452
rect 330 -6467 515 -6466
rect 330 -6512 455 -6467
rect 330 -6571 376 -6512
rect 440 -6513 455 -6512
rect 501 -6513 515 -6467
rect 440 -6526 515 -6513
rect 330 -6802 376 -6745
rect 573 -6571 619 -6409
rect 732 -6409 733 -6391
rect 732 -6437 779 -6409
rect 440 -6802 515 -6788
rect 330 -6803 515 -6802
rect 330 -6848 455 -6803
rect 330 -6907 376 -6848
rect 440 -6849 455 -6848
rect 501 -6849 515 -6803
rect 440 -6862 515 -6849
rect 330 -7138 376 -7081
rect 573 -6907 619 -6745
rect 440 -7138 515 -7124
rect 330 -7139 515 -7138
rect 330 -7184 455 -7139
rect 330 -7243 376 -7184
rect 440 -7185 455 -7184
rect 501 -7185 515 -7139
rect 440 -7198 515 -7185
rect 330 -7428 376 -7417
rect 573 -7243 619 -7081
rect 573 -7474 619 -7417
rect 733 -6571 779 -6437
rect 733 -6907 779 -6745
rect 733 -7243 779 -7081
rect 733 -7428 779 -7417
rect 893 -6235 939 -6224
rect 1052 -6235 1099 -6178
rect 893 -6571 939 -6409
rect 893 -6907 939 -6745
rect 893 -7243 939 -7081
rect 893 -7474 939 -7417
rect 1053 -6571 1099 -6409
rect 1053 -6907 1099 -6745
rect 1053 -7243 1099 -7081
rect 1053 -7428 1099 -7417
rect 1213 -6235 1259 -6224
rect 1372 -6235 1419 -6178
rect 2090 -6178 2776 -6176
rect 1213 -6571 1259 -6409
rect 1213 -6907 1259 -6745
rect 1213 -7243 1259 -7081
rect 1213 -7474 1259 -7417
rect 1373 -6571 1419 -6409
rect 1373 -6907 1419 -6745
rect 1373 -7243 1419 -7081
rect 1373 -7428 1419 -7417
rect 1533 -6235 1579 -6224
rect 1533 -6571 1579 -6409
rect 1533 -6907 1579 -6745
rect 1533 -7243 1579 -7081
rect 1533 -7474 1579 -7417
rect 573 -7522 1579 -7474
rect 1930 -6235 1976 -6224
rect 1930 -6571 1976 -6409
rect 1930 -6907 1976 -6745
rect 1930 -7243 1976 -7081
rect 1930 -7474 1976 -7417
rect 2090 -6235 2137 -6178
rect 2250 -6235 2296 -6224
rect 2090 -6571 2136 -6409
rect 2090 -6907 2136 -6745
rect 2090 -7243 2136 -7081
rect 2090 -7428 2136 -7417
rect 2250 -6571 2296 -6409
rect 2250 -6907 2296 -6745
rect 2250 -7243 2296 -7081
rect 2250 -7474 2296 -7417
rect 2410 -6235 2457 -6178
rect 2570 -6235 2616 -6224
rect 2410 -6571 2456 -6409
rect 2410 -6907 2456 -6745
rect 2410 -7243 2456 -7081
rect 2410 -7428 2456 -7417
rect 2570 -6571 2616 -6409
rect 2570 -6907 2616 -6745
rect 2570 -7243 2616 -7081
rect 2570 -7474 2616 -7417
rect 2730 -6235 2776 -6178
rect 2890 -6154 2936 -5827
rect 3133 -5317 3179 -5306
rect 3133 -5653 3179 -5491
rect 2990 -6041 3070 -6034
rect 2990 -6095 3002 -6041
rect 3056 -6095 3070 -6041
rect 2990 -6151 3070 -6095
rect 2990 -6154 3002 -6151
rect 2890 -6201 3002 -6154
rect 2890 -6235 2936 -6201
rect 2990 -6205 3002 -6201
rect 3056 -6205 3070 -6151
rect 2990 -6217 3070 -6205
rect 2776 -6409 2777 -6391
rect 2730 -6437 2777 -6409
rect 2730 -6571 2776 -6437
rect 2730 -6907 2776 -6745
rect 2730 -7243 2776 -7081
rect 2730 -7428 2776 -7417
rect 2890 -6571 2936 -6409
rect 3133 -6235 3179 -5827
rect 3293 -5317 3339 -5165
rect 3293 -5653 3339 -5491
rect 3470 -5310 3543 -5297
rect 3470 -5364 3480 -5310
rect 3534 -5364 3543 -5310
rect 3470 -5420 3543 -5364
rect 3470 -5474 3480 -5420
rect 3534 -5474 3543 -5420
rect 3470 -5493 3543 -5474
rect 3743 -5317 3789 -5165
rect 5247 -5166 7412 -5165
rect 7505 -2281 7676 486
rect 7747 -746 7936 -730
rect 7747 -802 7758 -746
rect 7814 -802 7868 -746
rect 7924 -802 7936 -746
rect 7747 -856 7936 -802
rect 7747 -912 7758 -856
rect 7814 -912 7868 -856
rect 7924 -912 7936 -856
rect 7747 -966 7936 -912
rect 7747 -1022 7758 -966
rect 7814 -1022 7868 -966
rect 7924 -1022 7936 -966
rect 7747 -1034 7936 -1022
rect 7505 -2298 7678 -2281
rect 7505 -2354 7509 -2298
rect 7565 -2354 7619 -2298
rect 7675 -2354 7678 -2298
rect 7505 -2408 7678 -2354
rect 7505 -2464 7509 -2408
rect 7565 -2464 7619 -2408
rect 7675 -2464 7678 -2408
rect 7505 -2518 7678 -2464
rect 7505 -2574 7509 -2518
rect 7565 -2574 7619 -2518
rect 7675 -2574 7678 -2518
rect 7505 -2586 7678 -2574
rect 4146 -5259 5152 -5211
rect 3293 -5838 3339 -5827
rect 3357 -5889 3433 -5881
rect 3239 -5892 3433 -5889
rect 3484 -5892 3530 -5493
rect 3743 -5653 3789 -5491
rect 3743 -5838 3789 -5827
rect 3903 -5317 3949 -5306
rect 3903 -5653 3949 -5491
rect 3649 -5889 3725 -5881
rect 3649 -5892 3843 -5889
rect 3239 -5894 3843 -5892
rect 3239 -5902 3371 -5894
rect 3239 -5948 3266 -5902
rect 3312 -5940 3371 -5902
rect 3419 -5940 3663 -5894
rect 3711 -5902 3843 -5894
rect 3711 -5940 3770 -5902
rect 3312 -5941 3770 -5940
rect 3312 -5948 3433 -5941
rect 3239 -5961 3433 -5948
rect 3649 -5948 3770 -5941
rect 3816 -5948 3843 -5902
rect 3649 -5961 3843 -5948
rect 3620 -6040 3697 -6028
rect 3620 -6096 3631 -6040
rect 3687 -6096 3697 -6040
rect 3620 -6130 3697 -6096
rect 3462 -6131 3518 -6130
rect 3385 -6150 3518 -6131
rect 3385 -6206 3395 -6150
rect 3451 -6184 3518 -6150
rect 3564 -6150 3697 -6130
rect 3564 -6184 3631 -6150
rect 3451 -6206 3462 -6184
rect 3385 -6219 3462 -6206
rect 3620 -6206 3631 -6184
rect 3687 -6206 3697 -6150
rect 3620 -6219 3697 -6206
rect 2994 -6466 3069 -6452
rect 3133 -6466 3179 -6409
rect 2994 -6467 3179 -6466
rect 2994 -6513 3008 -6467
rect 3054 -6512 3179 -6467
rect 3054 -6513 3069 -6512
rect 2994 -6526 3069 -6513
rect 2890 -6907 2936 -6745
rect 3133 -6571 3179 -6512
rect 2994 -6802 3069 -6788
rect 3133 -6802 3179 -6745
rect 2994 -6803 3179 -6802
rect 2994 -6849 3008 -6803
rect 3054 -6848 3179 -6803
rect 3054 -6849 3069 -6848
rect 2994 -6862 3069 -6849
rect 2890 -7243 2936 -7081
rect 3133 -6907 3179 -6848
rect 2994 -7138 3069 -7124
rect 3133 -7138 3179 -7081
rect 2994 -7139 3179 -7138
rect 2994 -7185 3008 -7139
rect 3054 -7184 3179 -7139
rect 3054 -7185 3069 -7184
rect 2994 -7198 3069 -7185
rect 2890 -7474 2936 -7417
rect 3133 -7243 3179 -7184
rect 3133 -7428 3179 -7417
rect 3293 -6235 3339 -6224
rect 3293 -6571 3339 -6409
rect 3293 -6907 3339 -6745
rect 3293 -7243 3339 -7081
rect 1930 -7522 2936 -7474
rect 1675 -7571 1838 -7570
rect 3293 -7571 3339 -7417
rect 3743 -6235 3789 -6224
rect 3743 -6571 3789 -6409
rect 3743 -6907 3789 -6745
rect 3743 -7243 3789 -7081
rect 3743 -7571 3789 -7417
rect 3903 -6235 3949 -5827
rect 4146 -5317 4192 -5259
rect 4146 -5653 4192 -5491
rect 4012 -6041 4089 -6033
rect 4011 -6097 4021 -6041
rect 4077 -6097 4089 -6041
rect 4012 -6151 4089 -6097
rect 4012 -6205 4026 -6151
rect 4080 -6154 4089 -6151
rect 4146 -6154 4192 -5827
rect 4306 -5317 4352 -5306
rect 4306 -5653 4352 -5491
rect 4306 -5885 4352 -5827
rect 4466 -5317 4512 -5259
rect 4466 -5653 4512 -5491
rect 4466 -5838 4512 -5827
rect 4626 -5317 4672 -5306
rect 4626 -5653 4672 -5491
rect 4626 -5885 4672 -5827
rect 4786 -5317 4832 -5259
rect 4786 -5653 4832 -5491
rect 4786 -5838 4832 -5827
rect 4946 -5317 4992 -5306
rect 4946 -5653 4992 -5491
rect 4946 -5885 4992 -5827
rect 5106 -5317 5152 -5259
rect 5610 -5260 6616 -5212
rect 5610 -5318 5656 -5260
rect 5106 -5653 5152 -5491
rect 5106 -5838 5152 -5827
rect 5321 -5342 5408 -5327
rect 5321 -5398 5335 -5342
rect 5391 -5398 5408 -5342
rect 5321 -5452 5408 -5398
rect 5321 -5508 5335 -5452
rect 5391 -5508 5408 -5452
rect 4306 -5994 4992 -5885
rect 4896 -6099 4992 -5994
rect 4080 -6201 4192 -6154
rect 4080 -6205 4089 -6201
rect 4012 -6217 4089 -6205
rect 3903 -6466 3949 -6409
rect 4146 -6235 4192 -6201
rect 4306 -6101 4992 -6099
rect 5321 -6101 5408 -5508
rect 5610 -5654 5656 -5492
rect 5610 -5839 5656 -5828
rect 5770 -5318 5816 -5307
rect 5770 -5654 5816 -5492
rect 5770 -5886 5816 -5828
rect 5930 -5318 5976 -5260
rect 5930 -5654 5976 -5492
rect 5930 -5839 5976 -5828
rect 6090 -5318 6136 -5307
rect 6090 -5654 6136 -5492
rect 6090 -5886 6136 -5828
rect 6250 -5318 6296 -5260
rect 6250 -5654 6296 -5492
rect 6250 -5839 6296 -5828
rect 6410 -5318 6456 -5307
rect 6410 -5654 6456 -5492
rect 6410 -5886 6456 -5828
rect 5770 -5995 6456 -5886
rect 6570 -5318 6616 -5260
rect 6570 -5654 6616 -5492
rect 5770 -6100 5866 -5995
rect 4306 -6102 5539 -6101
rect 5770 -6102 6456 -6100
rect 4306 -6176 6456 -6102
rect 4306 -6178 4992 -6176
rect 5285 -6177 6456 -6176
rect 4306 -6235 4352 -6178
rect 4013 -6466 4088 -6452
rect 3903 -6467 4088 -6466
rect 3903 -6512 4028 -6467
rect 3903 -6571 3949 -6512
rect 4013 -6513 4028 -6512
rect 4074 -6513 4088 -6467
rect 4013 -6526 4088 -6513
rect 3903 -6802 3949 -6745
rect 4146 -6571 4192 -6409
rect 4305 -6409 4306 -6391
rect 4305 -6437 4352 -6409
rect 4013 -6802 4088 -6788
rect 3903 -6803 4088 -6802
rect 3903 -6848 4028 -6803
rect 3903 -6907 3949 -6848
rect 4013 -6849 4028 -6848
rect 4074 -6849 4088 -6803
rect 4013 -6862 4088 -6849
rect 3903 -7138 3949 -7081
rect 4146 -6907 4192 -6745
rect 4013 -7138 4088 -7124
rect 3903 -7139 4088 -7138
rect 3903 -7184 4028 -7139
rect 3903 -7243 3949 -7184
rect 4013 -7185 4028 -7184
rect 4074 -7185 4088 -7139
rect 4013 -7198 4088 -7185
rect 3903 -7428 3949 -7417
rect 4146 -7243 4192 -7081
rect 4146 -7474 4192 -7417
rect 4306 -6571 4352 -6437
rect 4306 -6907 4352 -6745
rect 4306 -7243 4352 -7081
rect 4306 -7428 4352 -7417
rect 4466 -6235 4512 -6224
rect 4625 -6235 4672 -6178
rect 4466 -6571 4512 -6409
rect 4466 -6907 4512 -6745
rect 4466 -7243 4512 -7081
rect 4466 -7474 4512 -7417
rect 4626 -6571 4672 -6409
rect 4626 -6907 4672 -6745
rect 4626 -7243 4672 -7081
rect 4626 -7428 4672 -7417
rect 4786 -6235 4832 -6224
rect 4945 -6235 4992 -6178
rect 5770 -6179 6456 -6177
rect 4786 -6571 4832 -6409
rect 4786 -6907 4832 -6745
rect 4786 -7243 4832 -7081
rect 4786 -7474 4832 -7417
rect 4946 -6571 4992 -6409
rect 4946 -6907 4992 -6745
rect 4946 -7243 4992 -7081
rect 4946 -7428 4992 -7417
rect 5106 -6235 5152 -6224
rect 5106 -6571 5152 -6409
rect 5106 -6907 5152 -6745
rect 5106 -7243 5152 -7081
rect 5106 -7474 5152 -7417
rect 4146 -7522 5152 -7474
rect 5610 -6236 5656 -6225
rect 5610 -6572 5656 -6410
rect 5610 -6908 5656 -6746
rect 5610 -7244 5656 -7082
rect 5610 -7475 5656 -7418
rect 5770 -6236 5817 -6179
rect 5930 -6236 5976 -6225
rect 5770 -6572 5816 -6410
rect 5770 -6908 5816 -6746
rect 5770 -7244 5816 -7082
rect 5770 -7429 5816 -7418
rect 5930 -6572 5976 -6410
rect 5930 -6908 5976 -6746
rect 5930 -7244 5976 -7082
rect 5930 -7475 5976 -7418
rect 6090 -6236 6137 -6179
rect 6250 -6236 6296 -6225
rect 6090 -6572 6136 -6410
rect 6090 -6908 6136 -6746
rect 6090 -7244 6136 -7082
rect 6090 -7429 6136 -7418
rect 6250 -6572 6296 -6410
rect 6250 -6908 6296 -6746
rect 6250 -7244 6296 -7082
rect 6250 -7475 6296 -7418
rect 6410 -6236 6456 -6179
rect 6570 -6155 6616 -5828
rect 6813 -5318 6859 -5307
rect 6813 -5654 6859 -5492
rect 6673 -6042 6750 -6030
rect 6673 -6096 6682 -6042
rect 6736 -6096 6750 -6042
rect 6673 -6152 6750 -6096
rect 6673 -6155 6682 -6152
rect 6570 -6202 6682 -6155
rect 6570 -6236 6616 -6202
rect 6673 -6206 6682 -6202
rect 6736 -6206 6750 -6152
rect 6673 -6218 6750 -6206
rect 6456 -6410 6457 -6392
rect 6410 -6438 6457 -6410
rect 6410 -6572 6456 -6438
rect 6410 -6908 6456 -6746
rect 6410 -7244 6456 -7082
rect 6410 -7429 6456 -7418
rect 6570 -6572 6616 -6410
rect 6813 -6236 6859 -5828
rect 6973 -5318 7019 -5166
rect 6973 -5654 7019 -5492
rect 6973 -5839 7019 -5828
rect 7085 -5756 7176 -5742
rect 7085 -5810 7108 -5756
rect 7162 -5810 7176 -5756
rect 7085 -5866 7176 -5810
rect 7085 -5882 7108 -5866
rect 7037 -5890 7108 -5882
rect 6919 -5895 7108 -5890
rect 6919 -5903 7051 -5895
rect 6919 -5949 6946 -5903
rect 6992 -5941 7051 -5903
rect 7099 -5920 7108 -5895
rect 7162 -5893 7176 -5866
rect 7162 -5920 7198 -5893
rect 7099 -5941 7198 -5920
rect 6992 -5942 7198 -5941
rect 6992 -5944 7176 -5942
rect 6992 -5949 7113 -5944
rect 6919 -5962 7113 -5949
rect 7066 -6131 7143 -6130
rect 7066 -6132 7198 -6131
rect 7065 -6151 7198 -6132
rect 7065 -6207 7075 -6151
rect 7131 -6185 7198 -6151
rect 7131 -6207 7143 -6185
rect 7065 -6220 7143 -6207
rect 6674 -6467 6749 -6453
rect 6813 -6467 6859 -6410
rect 6674 -6468 6859 -6467
rect 6674 -6514 6688 -6468
rect 6734 -6513 6859 -6468
rect 6734 -6514 6749 -6513
rect 6674 -6527 6749 -6514
rect 6570 -6908 6616 -6746
rect 6813 -6572 6859 -6513
rect 6674 -6803 6749 -6789
rect 6813 -6803 6859 -6746
rect 6674 -6804 6859 -6803
rect 6674 -6850 6688 -6804
rect 6734 -6849 6859 -6804
rect 6734 -6850 6749 -6849
rect 6674 -6863 6749 -6850
rect 6570 -7244 6616 -7082
rect 6813 -6908 6859 -6849
rect 6674 -7139 6749 -7125
rect 6813 -7139 6859 -7082
rect 6674 -7140 6859 -7139
rect 6674 -7186 6688 -7140
rect 6734 -7185 6859 -7140
rect 6734 -7186 6749 -7185
rect 6674 -7199 6749 -7186
rect 6570 -7475 6616 -7418
rect 6813 -7244 6859 -7185
rect 6813 -7429 6859 -7418
rect 6973 -6236 7019 -6225
rect 7066 -6261 7143 -6220
rect 7066 -6317 7075 -6261
rect 7131 -6317 7143 -6261
rect 7066 -6334 7143 -6317
rect 6973 -6572 7019 -6410
rect 6973 -6908 7019 -6746
rect 6973 -7244 7019 -7082
rect 5610 -7523 6616 -7475
rect 71 -7572 5251 -7571
rect 6973 -7572 7019 -7418
rect 7505 -7441 7676 -2586
rect 7753 -3963 7936 -1034
rect 7744 -3976 7936 -3963
rect 7744 -4032 7753 -3976
rect 7809 -4032 7863 -3976
rect 7919 -4032 7936 -3976
rect 7744 -4086 7936 -4032
rect 7744 -4142 7753 -4086
rect 7809 -4142 7863 -4086
rect 7919 -4142 7936 -4086
rect 7744 -4196 7936 -4142
rect 7744 -4252 7753 -4196
rect 7809 -4252 7863 -4196
rect 7919 -4252 7936 -4196
rect 7744 -4267 7936 -4252
rect 7505 -7458 7678 -7441
rect 7505 -7514 7509 -7458
rect 7565 -7514 7619 -7458
rect 7675 -7514 7678 -7458
rect 7505 -7568 7678 -7514
rect -2528 -7579 7118 -7572
rect -4931 -7631 7118 -7579
rect -4931 -7632 131 -7631
rect -4931 -7639 -2285 -7632
rect -4931 -7693 -4688 -7639
rect -4527 -7693 -4467 -7639
rect -4306 -7693 -4246 -7639
rect -4085 -7693 -4025 -7639
rect -3864 -7693 -3804 -7639
rect -3643 -7693 -3583 -7639
rect -3422 -7693 -3362 -7639
rect -3201 -7693 -3141 -7639
rect -2980 -7686 -2285 -7639
rect -2124 -7686 -2064 -7632
rect -1903 -7686 -1843 -7632
rect -1682 -7686 -1622 -7632
rect -1461 -7686 -1401 -7632
rect -1240 -7686 -1180 -7632
rect -1019 -7686 -959 -7632
rect -798 -7686 -738 -7632
rect -577 -7685 131 -7632
rect 292 -7685 352 -7631
rect 513 -7685 573 -7631
rect 734 -7685 794 -7631
rect 955 -7685 1015 -7631
rect 1176 -7685 1236 -7631
rect 1397 -7685 1457 -7631
rect 1618 -7685 1891 -7631
rect 2052 -7685 2112 -7631
rect 2273 -7685 2333 -7631
rect 2494 -7685 2554 -7631
rect 2715 -7685 2775 -7631
rect 2936 -7685 2996 -7631
rect 3157 -7685 3217 -7631
rect 3378 -7685 3704 -7631
rect 3865 -7685 3925 -7631
rect 4086 -7685 4146 -7631
rect 4307 -7685 4367 -7631
rect 4528 -7685 4588 -7631
rect 4749 -7685 4809 -7631
rect 4970 -7685 5030 -7631
rect 5191 -7632 7118 -7631
rect 5191 -7685 5571 -7632
rect -577 -7686 5571 -7685
rect 5732 -7686 5792 -7632
rect 5953 -7686 6013 -7632
rect 6174 -7686 6234 -7632
rect 6395 -7686 6455 -7632
rect 6616 -7633 6676 -7632
rect 6837 -7633 6897 -7632
rect 6616 -7685 6627 -7633
rect 6837 -7685 6867 -7633
rect 6616 -7686 6676 -7685
rect 6837 -7686 6897 -7685
rect 7058 -7686 7118 -7632
rect -2980 -7693 7118 -7686
rect -4931 -7742 7118 -7693
rect -4931 -7746 -517 -7742
rect 71 -7745 7118 -7742
rect -4931 -7752 -2426 -7746
rect 3434 -7747 3656 -7745
rect 5511 -7746 7118 -7745
rect 7505 -7624 7509 -7568
rect 7565 -7624 7619 -7568
rect 7675 -7624 7678 -7568
rect 7505 -7678 7678 -7624
rect 7505 -7734 7509 -7678
rect 7565 -7734 7619 -7678
rect 7675 -7734 7678 -7678
rect 7505 -7746 7678 -7734
rect -4931 -7753 -2920 -7752
<< via1 >>
rect 6507 2635 6561 2687
rect 6627 2635 6676 2687
rect 6676 2635 6681 2687
rect 6747 2635 6801 2687
rect 6867 2635 6897 2687
rect 6897 2635 6921 2687
rect 6987 2635 7041 2687
rect -5197 1147 -5140 1204
rect -5197 1037 -5140 1094
rect -5104 885 -5048 941
rect -4994 912 -4980 941
rect -4980 912 -4938 941
rect -4994 885 -4938 912
rect -5170 654 -5113 711
rect -5170 544 -5113 601
rect -4145 1147 -4091 1201
rect -3020 1105 -2964 1161
rect -2909 1105 -2853 1161
rect -4149 1030 -4090 1089
rect -2681 874 -2625 930
rect -2571 919 -2531 930
rect -2531 919 -2515 930
rect -2571 874 -2515 919
rect -1742 1154 -1688 1208
rect -625 1113 -569 1169
rect -505 1114 -449 1170
rect 58 1154 114 1210
rect -1746 1037 -1687 1096
rect 58 1044 114 1100
rect -84 748 -27 805
rect -1009 108 -953 109
rect -899 108 -843 109
rect -789 108 -733 109
rect -679 108 -623 109
rect -1009 54 -959 108
rect -959 54 -953 108
rect -899 54 -843 108
rect -789 54 -738 108
rect -738 54 -733 108
rect -679 54 -623 108
rect -1009 53 -953 54
rect -899 53 -843 54
rect -789 53 -733 54
rect -679 53 -623 54
rect -5016 -679 -4960 -623
rect -5016 -764 -4960 -733
rect -5016 -789 -4980 -764
rect -4980 -789 -4960 -764
rect -5181 -972 -5123 -914
rect -5181 -1082 -5123 -1024
rect -5164 -1447 -5108 -1391
rect -5164 -1557 -5108 -1501
rect -5193 -3331 -5137 -3275
rect -5193 -3441 -5137 -3385
rect -5177 -4018 -5119 -3960
rect -5177 -4128 -5119 -4070
rect -2582 -680 -2526 -624
rect -2582 -757 -2526 -734
rect -2582 -790 -2577 -757
rect -2577 -790 -2531 -757
rect -2531 -790 -2526 -757
rect -4149 -941 -4090 -882
rect -4145 -1053 -4091 -999
rect -3039 -1014 -2983 -958
rect -2921 -1015 -2865 -959
rect -1746 -934 -1687 -875
rect -1742 -1046 -1688 -992
rect -621 -1006 -565 -950
rect -502 -1006 -446 -950
rect 453 1155 507 1209
rect 453 1045 507 1099
rect 3002 1265 3056 1319
rect 1721 360 1776 415
rect 1721 250 1776 305
rect 3002 1155 3056 1209
rect 7507 2675 7563 2731
rect 7617 2675 7673 2731
rect 3395 1264 3451 1320
rect 3395 1154 3451 1210
rect 3631 1264 3687 1320
rect 3631 1154 3687 1210
rect 3480 400 3534 454
rect 3480 290 3534 344
rect 4026 1155 4080 1209
rect 6685 1274 6739 1328
rect 5297 346 5353 402
rect 5297 236 5353 292
rect 6682 1154 6736 1208
rect 7507 2565 7563 2621
rect 7617 2565 7673 2621
rect 7507 2455 7563 2511
rect 7617 2455 7673 2511
rect 7075 1263 7131 1319
rect 7075 1153 7131 1209
rect 7161 858 7218 915
rect 7161 748 7218 805
rect 7509 718 7565 774
rect 7619 718 7675 774
rect 7509 608 7565 664
rect 7619 608 7675 664
rect 7509 498 7565 554
rect 7619 498 7675 554
rect 80 109 136 114
rect 190 109 246 114
rect 300 109 356 114
rect 410 109 466 114
rect 520 109 576 114
rect 80 58 131 109
rect 131 58 136 109
rect 190 58 246 109
rect 300 58 352 109
rect 352 58 356 109
rect 410 58 466 109
rect 520 58 573 109
rect 573 58 576 109
rect 849 -103 905 -102
rect 352 -159 408 -103
rect 477 -161 533 -105
rect 592 -161 648 -105
rect 719 -160 775 -104
rect 849 -158 871 -103
rect 871 -158 905 -103
rect 1004 -408 1058 -354
rect 1114 -408 1168 -354
rect 1338 -548 1395 -491
rect 1115 -672 1169 -618
rect 1338 -658 1395 -601
rect 1115 -782 1169 -728
rect -101 -1575 -45 -1519
rect -101 -1685 -45 -1629
rect 452 -1631 508 -1578
rect 587 -1631 643 -1577
rect 717 -1631 773 -1576
rect 860 -1631 879 -1577
rect 879 -1631 916 -1577
rect 452 -1634 508 -1631
rect 587 -1633 643 -1631
rect 717 -1632 773 -1631
rect 860 -1633 916 -1631
rect -328 -2075 -272 -2019
rect -218 -2075 -162 -2019
rect -1080 -2472 -1024 -2471
rect -970 -2472 -914 -2471
rect -860 -2472 -804 -2471
rect -750 -2472 -694 -2471
rect -640 -2472 -584 -2471
rect -1080 -2526 -1024 -2472
rect -970 -2526 -959 -2472
rect -959 -2526 -914 -2472
rect -860 -2526 -804 -2472
rect -750 -2526 -738 -2472
rect -738 -2526 -694 -2472
rect -640 -2526 -584 -2472
rect -1080 -2527 -1024 -2526
rect -970 -2527 -914 -2526
rect -860 -2527 -804 -2526
rect -750 -2527 -694 -2526
rect -640 -2527 -584 -2526
rect -5030 -4248 -4980 -4209
rect -4980 -4248 -4974 -4209
rect -5030 -4265 -4974 -4248
rect -5030 -4375 -4974 -4319
rect -5225 -5575 -5168 -5518
rect -5225 -5685 -5168 -5628
rect -4145 -4013 -4091 -3959
rect -3040 -4053 -2984 -3997
rect -2919 -4053 -2863 -3997
rect -4149 -4130 -4090 -4071
rect -2595 -4241 -2577 -4200
rect -2577 -4241 -2539 -4200
rect -2595 -4256 -2539 -4241
rect -2595 -4366 -2539 -4310
rect -1742 -4006 -1688 -3952
rect -658 -4046 -602 -3990
rect -520 -4045 -464 -3989
rect -1746 -4123 -1687 -4064
rect -331 -4396 -271 -4336
rect -218 -4396 -158 -4336
rect -1189 -5052 -1133 -5050
rect -1079 -5052 -1023 -5050
rect -969 -5052 -913 -5050
rect -859 -5052 -803 -5050
rect -749 -5052 -693 -5050
rect -639 -5052 -583 -5050
rect -1189 -5106 -1180 -5052
rect -1180 -5106 -1133 -5052
rect -1079 -5106 -1023 -5052
rect -969 -5106 -959 -5052
rect -959 -5106 -913 -5052
rect -859 -5106 -803 -5052
rect -749 -5106 -738 -5052
rect -738 -5106 -693 -5052
rect -639 -5106 -583 -5052
rect -5019 -5834 -4963 -5778
rect -5019 -5924 -4963 -5888
rect -5019 -5944 -4980 -5924
rect -4980 -5944 -4963 -5924
rect -5119 -6106 -5062 -6049
rect -5119 -6216 -5062 -6159
rect -2601 -5838 -2545 -5782
rect -2601 -5917 -2545 -5892
rect -2601 -5948 -2577 -5917
rect -2577 -5948 -2545 -5917
rect -4149 -6101 -4090 -6042
rect -4145 -6213 -4091 -6159
rect -3038 -6173 -2982 -6117
rect -2908 -6173 -2852 -6117
rect 24 -2075 80 -2019
rect 24 -2185 80 -2129
rect 756 -2224 810 -2170
rect 866 -2224 920 -2170
rect 395 -3103 451 -3047
rect 513 -3101 569 -3045
rect 637 -3100 693 -3044
rect 746 -3100 802 -3044
rect 866 -3102 871 -3046
rect 871 -3102 922 -3046
rect 19 -4277 73 -4223
rect 19 -4387 73 -4333
rect 765 -3975 819 -3921
rect 875 -3975 929 -3921
rect 1225 -916 1281 -860
rect 1225 -1026 1281 -970
rect 1226 -1964 1280 -1910
rect 1226 -2074 1280 -2020
rect 1115 -2219 1169 -2165
rect 1115 -2329 1169 -2275
rect 1115 -4139 1169 -4085
rect 1115 -4249 1169 -4195
rect 2330 -140 2384 -86
rect 2646 -145 2702 -89
rect 1635 -783 1689 -729
rect 1745 -783 1799 -729
rect 1818 -1046 1874 -990
rect 1492 -1447 1548 -1391
rect 1492 -1557 1548 -1501
rect 1492 -1667 1548 -1611
rect 2213 -1045 2267 -991
rect 2966 -145 3022 -89
rect 3288 -144 3344 -88
rect 3735 -146 3791 -90
rect 4057 -147 4113 -91
rect 4378 -144 4434 -88
rect 4699 -153 4753 -99
rect 3512 -1119 3566 -1065
rect 3512 -1229 3566 -1175
rect 4815 -1045 4869 -991
rect 5394 -514 5448 -460
rect 5394 -624 5448 -570
rect 5269 -789 5325 -733
rect 5269 -899 5325 -843
rect 5208 -1046 5264 -990
rect 5498 -1047 5554 -991
rect 5498 -1157 5554 -1101
rect 5893 -1046 5947 -992
rect 7078 -801 7132 -747
rect 7078 -911 7132 -857
rect 5893 -1156 5947 -1102
rect 7078 -1021 7132 -967
rect 6507 -2525 6561 -2473
rect 6627 -2525 6676 -2473
rect 6676 -2525 6681 -2473
rect 6747 -2525 6801 -2473
rect 6867 -2525 6897 -2473
rect 6897 -2525 6921 -2473
rect 6987 -2525 7041 -2473
rect 1702 -2917 1758 -2861
rect 1702 -3027 1758 -2971
rect 1702 -3137 1758 -3081
rect 1333 -3865 1390 -3808
rect 1333 -3975 1390 -3918
rect 1818 -4006 1874 -3950
rect 1004 -4566 1058 -4512
rect 1114 -4566 1168 -4512
rect 2213 -4005 2267 -3951
rect 3533 -3881 3591 -3823
rect 3533 -3991 3591 -3933
rect 2337 -4839 2379 -4837
rect 2379 -4839 2391 -4837
rect 2337 -4891 2391 -4839
rect 2645 -4839 2653 -4832
rect 2653 -4839 2699 -4832
rect 2699 -4839 2701 -4832
rect 2645 -4888 2701 -4839
rect 2966 -4901 3022 -4845
rect 3283 -4904 3339 -4848
rect 3745 -4904 3801 -4848
rect 4057 -4902 4113 -4846
rect 4377 -4899 4433 -4843
rect 4815 -4005 4869 -3951
rect 5498 -3897 5554 -3841
rect 5208 -4006 5264 -3950
rect 5498 -4007 5554 -3951
rect 5253 -4155 5309 -4099
rect 5253 -4265 5309 -4209
rect 4699 -4897 4753 -4843
rect 5419 -4397 5473 -4343
rect 5419 -4507 5473 -4453
rect 5889 -3896 5943 -3842
rect 5893 -4006 5947 -3952
rect 7096 -4031 7150 -3977
rect 7096 -4141 7150 -4087
rect 7096 -4251 7150 -4197
rect 86 -5051 142 -5050
rect 196 -5051 252 -5050
rect 306 -5051 362 -5050
rect 416 -5051 472 -5050
rect 526 -5051 582 -5050
rect 636 -5051 692 -5050
rect 746 -5051 802 -5050
rect 86 -5105 131 -5051
rect 131 -5105 142 -5051
rect 196 -5105 252 -5051
rect 306 -5105 352 -5051
rect 352 -5105 362 -5051
rect 416 -5105 472 -5051
rect 526 -5105 573 -5051
rect 573 -5105 582 -5051
rect 636 -5105 692 -5051
rect 746 -5105 794 -5051
rect 794 -5105 802 -5051
rect 86 -5106 142 -5105
rect 196 -5106 252 -5105
rect 306 -5106 362 -5105
rect 416 -5106 472 -5105
rect 526 -5106 582 -5105
rect 636 -5106 692 -5105
rect 746 -5106 802 -5105
rect -85 -5703 -28 -5646
rect -85 -5813 -28 -5756
rect -1746 -6094 -1687 -6035
rect -1742 -6206 -1688 -6152
rect 57 -6097 113 -6041
rect -633 -6166 -577 -6110
rect -508 -6166 -452 -6110
rect 58 -6206 114 -6150
rect 448 -6096 504 -6040
rect 453 -6205 507 -6151
rect 1728 -5392 1783 -5337
rect 1728 -5502 1783 -5447
rect 3002 -6095 3056 -6041
rect 3002 -6205 3056 -6151
rect 3480 -5364 3534 -5310
rect 3480 -5474 3534 -5420
rect 7758 -802 7814 -746
rect 7868 -802 7924 -746
rect 7758 -912 7814 -856
rect 7868 -912 7924 -856
rect 7758 -1022 7814 -966
rect 7868 -1022 7924 -966
rect 7509 -2354 7565 -2298
rect 7619 -2354 7675 -2298
rect 7509 -2464 7565 -2408
rect 7619 -2464 7675 -2408
rect 7509 -2574 7565 -2518
rect 7619 -2574 7675 -2518
rect 3631 -6096 3687 -6040
rect 3395 -6206 3451 -6150
rect 3631 -6206 3687 -6150
rect 4021 -6097 4077 -6041
rect 4026 -6205 4080 -6151
rect 5335 -5398 5391 -5342
rect 5335 -5508 5391 -5452
rect 6682 -6096 6736 -6042
rect 6682 -6206 6736 -6152
rect 7108 -5810 7162 -5756
rect 7108 -5920 7162 -5866
rect 7075 -6207 7131 -6151
rect 7075 -6317 7131 -6261
rect 7753 -4032 7809 -3976
rect 7863 -4032 7919 -3976
rect 7753 -4142 7809 -4086
rect 7863 -4142 7919 -4086
rect 7753 -4252 7809 -4196
rect 7863 -4252 7919 -4196
rect 7509 -7514 7565 -7458
rect 7619 -7514 7675 -7458
rect 6507 -7685 6561 -7633
rect 6627 -7685 6676 -7633
rect 6676 -7685 6681 -7633
rect 6747 -7685 6801 -7633
rect 6867 -7685 6897 -7633
rect 6897 -7685 6921 -7633
rect 6987 -7685 7041 -7633
rect 7509 -7624 7565 -7568
rect 7619 -7624 7675 -7568
rect 7509 -7734 7565 -7678
rect 7619 -7734 7675 -7678
<< metal2 >>
rect 6445 2731 7676 2748
rect 6445 2687 7507 2731
rect 6445 2635 6507 2687
rect 6561 2635 6627 2687
rect 6681 2635 6747 2687
rect 6801 2635 6867 2687
rect 6921 2635 6987 2687
rect 7041 2675 7507 2687
rect 7563 2675 7617 2731
rect 7673 2675 7676 2731
rect 7041 2635 7676 2675
rect 6445 2621 7676 2635
rect 6445 2574 7507 2621
rect 7503 2565 7507 2574
rect 7563 2565 7617 2621
rect 7673 2565 7676 2621
rect 7503 2511 7676 2565
rect -3019 2367 7142 2480
rect 7503 2455 7507 2511
rect 7563 2455 7617 2511
rect 7673 2455 7676 2511
rect 7503 2443 7676 2455
rect -5214 1204 -5093 1208
rect -5214 1147 -5197 1204
rect -5140 1202 -5093 1204
rect -4159 1202 -4082 1213
rect -5140 1201 -4082 1202
rect -5140 1147 -4145 1201
rect -4091 1147 -4082 1201
rect -3019 1172 -2906 2367
rect -591 1933 3696 2047
rect -1756 1209 -1679 1220
rect -2593 1208 -1679 1209
rect -5214 1094 -4082 1147
rect -3028 1161 -2840 1172
rect -3028 1105 -3020 1161
rect -2964 1105 -2909 1161
rect -2853 1105 -2840 1161
rect -3028 1097 -2840 1105
rect -2593 1154 -1742 1208
rect -1688 1154 -1679 1208
rect -591 1180 -477 1933
rect -174 1655 3070 1684
rect -174 1599 -159 1655
rect -103 1653 3070 1655
rect -103 1599 -40 1653
rect -174 1597 -40 1599
rect 16 1597 67 1653
rect 123 1597 3070 1653
rect -174 1568 3070 1597
rect 2943 1319 3070 1568
rect 3385 1320 3462 1332
rect 3385 1319 3395 1320
rect 2943 1265 3002 1319
rect 3056 1265 3395 1319
rect 2943 1264 3395 1265
rect 3451 1264 3462 1320
rect -59 1221 129 1223
rect -59 1210 517 1221
rect -59 1206 57 1210
rect -591 1179 -449 1180
rect -3020 1095 -2964 1097
rect -2593 1096 -1679 1154
rect -637 1170 -437 1179
rect -637 1169 -505 1170
rect -637 1113 -625 1169
rect -569 1114 -505 1169
rect -449 1114 -437 1170
rect -569 1113 -437 1114
rect -637 1104 -437 1113
rect -59 1150 -47 1206
rect 9 1154 57 1206
rect 114 1209 517 1210
rect 114 1155 453 1209
rect 507 1155 517 1209
rect 114 1154 517 1155
rect 9 1150 517 1154
rect -625 1103 -569 1104
rect -5214 1037 -5197 1094
rect -5140 1089 -4082 1094
rect -5140 1037 -4149 1089
rect -5214 1030 -4149 1037
rect -4090 1030 -4082 1089
rect -2593 1037 -1746 1096
rect -1687 1037 -1679 1096
rect -2593 1033 -1679 1037
rect -5214 1026 -4082 1030
rect -4159 1017 -4082 1026
rect -5111 958 -4887 969
rect -2689 958 -2481 974
rect -5111 941 -2481 958
rect -5111 885 -5104 941
rect -5048 885 -4994 941
rect -4938 930 -2481 941
rect -4938 885 -2681 930
rect -5111 874 -2681 885
rect -2625 874 -2571 930
rect -2515 874 -2481 930
rect -5111 868 -2481 874
rect -5111 853 -4887 868
rect -2689 830 -2481 868
rect -5197 711 -5101 714
rect -5197 654 -5170 711
rect -5113 699 -5101 711
rect -2219 699 -2062 1033
rect -1756 1024 -1679 1033
rect -59 1101 517 1150
rect 2943 1210 3462 1264
rect 2943 1209 3395 1210
rect 2943 1155 3002 1209
rect 3056 1155 3395 1209
rect 2943 1154 3395 1155
rect 3451 1154 3462 1210
rect 2943 1142 3070 1154
rect 3385 1135 3462 1154
rect 3573 1320 3696 1933
rect 3573 1264 3631 1320
rect 3687 1264 3696 1320
rect 3573 1223 3696 1264
rect 6673 1328 6750 1339
rect 6673 1274 6685 1328
rect 6739 1306 6750 1328
rect 7018 1319 7142 2367
rect 7018 1306 7075 1319
rect 6739 1274 7075 1306
rect 6673 1263 7075 1274
rect 7131 1263 7142 1319
rect 3573 1210 3697 1223
rect 4012 1210 4089 1221
rect 3573 1154 3631 1210
rect 3687 1209 4089 1210
rect 3687 1155 4026 1209
rect 4080 1155 4089 1209
rect 3687 1154 4089 1155
rect 3573 1135 3697 1154
rect 4012 1143 4089 1154
rect 6673 1209 7142 1263
rect 6673 1208 7075 1209
rect 6673 1154 6682 1208
rect 6736 1154 7075 1208
rect 6673 1153 7075 1154
rect 7131 1153 7142 1209
rect 6673 1142 6750 1153
rect 3573 1134 3696 1135
rect 7018 1126 7142 1153
rect -59 1045 -47 1101
rect 9 1100 517 1101
rect 9 1045 58 1100
rect -59 1044 58 1045
rect 114 1099 517 1100
rect 114 1053 453 1099
rect 114 1044 129 1053
rect -59 1028 129 1044
rect 438 1045 453 1053
rect 507 1045 517 1099
rect 438 1033 517 1045
rect 7144 915 7234 944
rect 7144 858 7161 915
rect 7218 858 7234 915
rect -102 805 -13 821
rect 7144 805 7234 858
rect -102 748 -84 805
rect -27 748 7161 805
rect 7218 748 7234 805
rect -102 732 -13 748
rect 7144 739 7234 748
rect 7505 774 7678 791
rect -5113 654 -2062 699
rect 7505 718 7509 774
rect 7565 718 7619 774
rect 7675 718 7678 774
rect 7505 682 7678 718
rect -5197 601 -2062 654
rect -5197 544 -5170 601
rect -5113 544 -2062 601
rect -5197 542 -2062 544
rect 824 664 7678 682
rect 824 608 7509 664
rect 7565 608 7619 664
rect 7675 608 7678 664
rect 824 554 7678 608
rect -5197 540 -5101 542
rect 824 540 7509 554
rect -1023 114 645 170
rect -1023 109 80 114
rect -1023 53 -1009 109
rect -953 53 -899 109
rect -843 53 -789 109
rect -733 53 -679 109
rect -623 58 80 109
rect 136 58 190 114
rect 246 58 300 114
rect 356 58 410 114
rect 466 58 520 114
rect 576 58 645 114
rect -623 53 645 58
rect -1023 -6 645 53
rect 824 -74 966 540
rect 7505 498 7509 540
rect 7565 498 7619 554
rect 7675 498 7678 554
rect 7505 486 7678 498
rect 3470 454 3543 466
rect 342 -102 966 -74
rect 342 -103 849 -102
rect 342 -159 352 -103
rect 408 -104 849 -103
rect 408 -105 719 -104
rect 408 -159 477 -105
rect 342 -161 477 -159
rect 533 -161 592 -105
rect 648 -160 719 -105
rect 775 -158 849 -104
rect 905 -158 966 -102
rect 1708 415 1788 430
rect 1708 360 1721 415
rect 1776 360 1788 415
rect 1708 305 1788 360
rect 1708 250 1721 305
rect 1776 250 1788 305
rect 3470 400 3480 454
rect 3534 400 3543 454
rect 3470 344 3543 400
rect 3470 290 3480 344
rect 3534 290 3543 344
rect 3470 277 3543 290
rect 5285 402 5365 415
rect 5285 346 5297 402
rect 5353 346 5365 402
rect 5285 292 5365 346
rect 1708 -71 1788 250
rect 1708 -86 3363 -71
rect 1708 -140 2330 -86
rect 2384 -88 3363 -86
rect 2384 -89 3288 -88
rect 2384 -140 2646 -89
rect 1708 -145 2646 -140
rect 2702 -145 2966 -89
rect 3022 -144 3288 -89
rect 3344 -144 3363 -88
rect 3022 -145 3363 -144
rect 1708 -154 3363 -145
rect 2646 -155 2702 -154
rect 2966 -155 3022 -154
rect 775 -160 966 -158
rect 648 -161 966 -160
rect 342 -174 966 -161
rect 991 -350 1178 -341
rect 3482 -350 3538 277
rect 5285 236 5297 292
rect 5353 236 5365 292
rect 3718 -86 3804 -80
rect 4041 -86 4127 -80
rect 4361 -86 4447 -75
rect 5285 -86 5365 236
rect 3718 -88 5365 -86
rect 3718 -90 4378 -88
rect 3718 -146 3735 -90
rect 3791 -91 4378 -90
rect 3791 -146 4057 -91
rect 3718 -147 4057 -146
rect 4113 -144 4378 -91
rect 4434 -99 5365 -88
rect 4434 -144 4699 -99
rect 4113 -147 4699 -144
rect 3718 -153 4699 -147
rect 4753 -153 5365 -99
rect 3718 -164 5365 -153
rect 991 -354 3538 -350
rect 991 -408 1004 -354
rect 1058 -408 1114 -354
rect 1168 -406 3538 -354
rect 1168 -408 1178 -406
rect 991 -420 1178 -408
rect 5384 -460 5457 -444
rect 1326 -491 1407 -481
rect 1326 -548 1338 -491
rect 1395 -548 1407 -491
rect 1326 -568 1407 -548
rect 5384 -514 5394 -460
rect 5448 -514 5457 -460
rect 5384 -568 5457 -514
rect 1326 -570 5457 -568
rect 1326 -601 5394 -570
rect -5041 -623 -4935 -615
rect -5041 -679 -5016 -623
rect -4960 -659 -4935 -623
rect -2601 -624 -2501 -611
rect -2601 -659 -2582 -624
rect -4960 -679 -2582 -659
rect -5041 -680 -2582 -679
rect -2526 -680 -2501 -624
rect -5041 -733 -2501 -680
rect -5041 -789 -5016 -733
rect -4960 -734 -2501 -733
rect -4960 -770 -2582 -734
rect -4960 -789 -4935 -770
rect -5041 -804 -4935 -789
rect -2601 -790 -2582 -770
rect -2526 -790 -2501 -734
rect -2601 -806 -2501 -790
rect 1106 -618 1178 -607
rect 1106 -672 1115 -618
rect 1169 -672 1178 -618
rect 1326 -658 1338 -601
rect 1395 -624 5394 -601
rect 5448 -624 5457 -570
rect 1395 -625 5457 -624
rect 1395 -658 1407 -625
rect 5384 -635 5457 -625
rect 1326 -670 1407 -658
rect 1106 -726 1178 -672
rect 1623 -726 1856 -718
rect 1106 -728 1856 -726
rect 1106 -782 1115 -728
rect 1169 -729 1856 -728
rect 1169 -782 1635 -729
rect 1106 -795 1178 -782
rect 1623 -783 1635 -782
rect 1689 -783 1745 -729
rect 1799 -783 1856 -729
rect 1623 -795 1856 -783
rect 5255 -733 5337 -720
rect 5255 -789 5269 -733
rect 5325 -789 5337 -733
rect 5255 -843 5337 -789
rect 1213 -858 1293 -848
rect 5255 -858 5269 -843
rect 1213 -860 5269 -858
rect -4159 -878 -4082 -869
rect -1756 -871 -1679 -862
rect -5194 -882 -4082 -878
rect -5194 -914 -4149 -882
rect -5194 -972 -5181 -914
rect -5123 -941 -4149 -914
rect -4090 -941 -4082 -882
rect -5123 -972 -4082 -941
rect -2593 -875 -1679 -871
rect -2593 -934 -1746 -875
rect -1687 -934 -1679 -875
rect -5194 -999 -4082 -972
rect -5194 -1024 -4145 -999
rect -5194 -1082 -5181 -1024
rect -5123 -1053 -4145 -1024
rect -4091 -1053 -4082 -999
rect -3049 -958 -2839 -948
rect -3049 -1014 -3039 -958
rect -2983 -959 -2839 -958
rect -2983 -1014 -2921 -959
rect -3049 -1015 -2921 -1014
rect -2865 -1015 -2839 -959
rect -3049 -1025 -2839 -1015
rect -2593 -992 -1679 -934
rect 1213 -916 1225 -860
rect 1281 -899 5269 -860
rect 5325 -899 5337 -843
rect 1281 -914 5337 -899
rect 7066 -747 7145 -731
rect 7066 -801 7078 -747
rect 7132 -801 7145 -747
rect 7066 -808 7145 -801
rect 7747 -746 7936 -730
rect 7747 -802 7758 -746
rect 7814 -802 7868 -746
rect 7924 -802 7936 -746
rect 7747 -808 7936 -802
rect 7066 -856 7936 -808
rect 7066 -857 7758 -856
rect 7066 -911 7078 -857
rect 7132 -911 7758 -857
rect 7066 -912 7758 -911
rect 7814 -912 7868 -856
rect 7924 -912 7936 -856
rect 1281 -916 1293 -914
rect -621 -942 -565 -940
rect -502 -942 -446 -940
rect -2593 -1046 -1742 -992
rect -1688 -1046 -1679 -992
rect -630 -950 -436 -942
rect -630 -1006 -621 -950
rect -565 -1006 -502 -950
rect -446 -1006 -436 -950
rect -630 -1017 -436 -1006
rect 1213 -970 1293 -916
rect 7066 -966 7936 -912
rect 7066 -967 7758 -966
rect 1213 -1026 1225 -970
rect 1281 -1026 1293 -970
rect 1213 -1033 1293 -1026
rect 1807 -990 1884 -971
rect 2199 -990 2276 -979
rect -2593 -1047 -1679 -1046
rect -5123 -1054 -4082 -1053
rect -5123 -1082 -5099 -1054
rect -4159 -1065 -4082 -1054
rect -5194 -1094 -5099 -1082
rect -5189 -1386 -5094 -1381
rect -2279 -1386 -2122 -1047
rect -1756 -1058 -1679 -1047
rect 1807 -1046 1818 -990
rect 1874 -991 2276 -990
rect 1874 -1045 2213 -991
rect 2267 -1045 2276 -991
rect 4806 -990 4883 -979
rect 5198 -990 5275 -971
rect 4806 -991 5208 -990
rect 1874 -1046 2276 -1045
rect 1807 -1059 1884 -1046
rect 2199 -1057 2276 -1046
rect 3492 -1065 3604 -1016
rect 4806 -1045 4815 -991
rect 4869 -1045 5208 -991
rect 4806 -1046 5208 -1045
rect 5264 -1046 5275 -990
rect 4806 -1057 4883 -1046
rect 5198 -1059 5275 -1046
rect 5442 -980 5564 -970
rect 5442 -991 5956 -980
rect 5442 -1047 5498 -991
rect 5554 -992 5956 -991
rect 5554 -1046 5893 -992
rect 5947 -1046 5956 -992
rect 7066 -1021 7078 -967
rect 7132 -1021 7758 -967
rect 7066 -1022 7758 -1021
rect 7814 -1022 7868 -966
rect 7924 -1022 7936 -966
rect 7066 -1034 7146 -1022
rect 7747 -1034 7936 -1022
rect 5554 -1047 5956 -1046
rect 3492 -1119 3512 -1065
rect 3566 -1119 3604 -1065
rect 3492 -1142 3604 -1119
rect 5442 -1101 5956 -1047
rect 5442 -1142 5498 -1101
rect 3492 -1157 5498 -1142
rect 5554 -1102 5956 -1101
rect 5554 -1156 5893 -1102
rect 5947 -1156 5956 -1102
rect 5554 -1157 5956 -1156
rect 3492 -1174 5956 -1157
rect 3492 -1175 5564 -1174
rect 5878 -1175 5956 -1174
rect 3492 -1229 3512 -1175
rect 3566 -1229 5564 -1175
rect 3492 -1254 5564 -1229
rect -5189 -1391 -2122 -1386
rect -5189 -1447 -5164 -1391
rect -5108 -1447 -2122 -1391
rect -5189 -1501 -2122 -1447
rect -5189 -1557 -5164 -1501
rect -5108 -1543 -2122 -1501
rect 1458 -1391 1584 -1389
rect 1458 -1447 1492 -1391
rect 1548 -1447 1584 -1391
rect 1458 -1501 1584 -1447
rect -126 -1519 -31 -1509
rect -5108 -1557 -5094 -1543
rect -5189 -1567 -5094 -1557
rect -126 -1575 -101 -1519
rect -45 -1575 -31 -1519
rect 1458 -1557 1492 -1501
rect 1548 -1557 1584 -1501
rect 1458 -1559 1584 -1557
rect -126 -1629 -31 -1575
rect -126 -1635 -101 -1629
rect -5286 -1685 -101 -1635
rect -45 -1685 -31 -1629
rect 441 -1576 1584 -1559
rect 441 -1577 717 -1576
rect 441 -1578 587 -1577
rect 441 -1634 452 -1578
rect 508 -1633 587 -1578
rect 643 -1632 717 -1577
rect 773 -1577 1584 -1576
rect 773 -1632 860 -1577
rect 643 -1633 860 -1632
rect 916 -1611 1584 -1577
rect 916 -1633 1492 -1611
rect 508 -1634 1492 -1633
rect 441 -1667 1492 -1634
rect 1548 -1667 1584 -1611
rect 441 -1674 1584 -1667
rect -5286 -1691 -31 -1685
rect -126 -1695 -31 -1691
rect 1216 -1910 1287 -1898
rect 1216 -1964 1226 -1910
rect 1280 -1964 1287 -1910
rect -340 -2019 -150 -2011
rect 7 -2019 92 -2007
rect 1216 -2019 1287 -1964
rect -5292 -2075 -328 -2019
rect -272 -2075 -218 -2019
rect -162 -2075 24 -2019
rect 80 -2020 1287 -2019
rect 80 -2074 1226 -2020
rect 1280 -2074 1287 -2020
rect 80 -2075 1287 -2074
rect -340 -2082 -150 -2075
rect 7 -2129 92 -2075
rect 1216 -2087 1287 -2075
rect 7 -2185 24 -2129
rect 80 -2185 92 -2129
rect 7 -2195 92 -2185
rect 746 -2166 935 -2155
rect 1104 -2165 1180 -2153
rect 1104 -2166 1115 -2165
rect 746 -2170 1115 -2166
rect 746 -2224 756 -2170
rect 810 -2224 866 -2170
rect 920 -2219 1115 -2170
rect 1169 -2219 1180 -2165
rect 920 -2222 1180 -2219
rect 920 -2224 935 -2222
rect 746 -2238 935 -2224
rect 1104 -2275 1180 -2222
rect 1104 -2329 1115 -2275
rect 1169 -2329 1180 -2275
rect 1104 -2340 1180 -2329
rect 7505 -2298 7678 -2281
rect 7505 -2354 7509 -2298
rect 7565 -2354 7619 -2298
rect 7675 -2354 7678 -2298
rect 7505 -2408 7678 -2354
rect 7505 -2412 7509 -2408
rect -1090 -2428 -518 -2412
rect -1090 -2471 -258 -2428
rect -1090 -2527 -1080 -2471
rect -1024 -2527 -970 -2471
rect -914 -2527 -860 -2471
rect -804 -2527 -750 -2471
rect -694 -2527 -640 -2471
rect -584 -2527 -258 -2471
rect -1090 -2552 -258 -2527
rect -1090 -2585 -518 -2552
rect -382 -3020 -258 -2552
rect 6445 -2464 7509 -2412
rect 7565 -2464 7619 -2408
rect 7675 -2464 7678 -2408
rect 6445 -2473 7678 -2464
rect 6445 -2525 6507 -2473
rect 6561 -2525 6627 -2473
rect 6681 -2525 6747 -2473
rect 6801 -2525 6867 -2473
rect 6921 -2525 6987 -2473
rect 7041 -2518 7678 -2473
rect 7041 -2525 7509 -2518
rect 6445 -2574 7509 -2525
rect 7565 -2574 7619 -2518
rect 7675 -2574 7678 -2518
rect 6445 -2586 7678 -2574
rect 1666 -2861 1794 -2850
rect 1666 -2917 1702 -2861
rect 1758 -2917 1794 -2861
rect 1666 -2971 1794 -2917
rect 373 -3020 922 -3019
rect 1666 -3020 1702 -2971
rect -382 -3027 1702 -3020
rect 1758 -3027 1794 -2971
rect -382 -3044 1794 -3027
rect -382 -3045 637 -3044
rect -382 -3047 513 -3045
rect -382 -3103 395 -3047
rect 451 -3101 513 -3047
rect 569 -3100 637 -3045
rect 693 -3100 746 -3044
rect 802 -3046 1794 -3044
rect 802 -3100 866 -3046
rect 569 -3101 866 -3100
rect 451 -3102 866 -3101
rect 922 -3081 1794 -3046
rect 922 -3102 1702 -3081
rect 451 -3103 1702 -3102
rect -382 -3137 1702 -3103
rect 1758 -3137 1794 -3081
rect -382 -3143 1794 -3137
rect -382 -3144 1702 -3143
rect -5193 -3268 -5137 -3265
rect -5209 -3275 -5121 -3268
rect -5209 -3331 -5193 -3275
rect -5137 -3293 -5121 -3275
rect -5137 -3331 -2150 -3293
rect -5209 -3385 -2150 -3331
rect -5209 -3441 -5193 -3385
rect -5137 -3407 -2150 -3385
rect -5137 -3441 -5121 -3407
rect -5209 -3458 -5121 -3441
rect -5189 -3958 -5107 -3947
rect -4159 -3958 -4082 -3947
rect -2264 -3951 -2150 -3407
rect 1323 -3808 1405 -3796
rect 1323 -3865 1333 -3808
rect 1390 -3865 1405 -3808
rect 749 -3918 941 -3906
rect 1323 -3918 1405 -3865
rect 749 -3921 1333 -3918
rect -1756 -3951 -1679 -3940
rect -5189 -3959 -4082 -3958
rect -5189 -3960 -4145 -3959
rect -5189 -4018 -5177 -3960
rect -5119 -4013 -4145 -3960
rect -4091 -4013 -4082 -3959
rect -2593 -3952 -1679 -3951
rect -3040 -3988 -2984 -3987
rect -2919 -3988 -2863 -3987
rect -5119 -4018 -4082 -4013
rect -5189 -4070 -4082 -4018
rect -3050 -3997 -2840 -3988
rect -3050 -4053 -3040 -3997
rect -2984 -4053 -2919 -3997
rect -2863 -4053 -2840 -3997
rect -3050 -4063 -2840 -4053
rect -2593 -4006 -1742 -3952
rect -1688 -4006 -1679 -3952
rect 749 -3975 765 -3921
rect 819 -3975 875 -3921
rect 929 -3975 1333 -3921
rect 1390 -3975 1405 -3918
rect 3520 -3823 5564 -3765
rect 3520 -3881 3533 -3823
rect 3591 -3838 5564 -3823
rect 5876 -3838 5956 -3836
rect 3591 -3841 5956 -3838
rect 3591 -3881 5498 -3841
rect 3520 -3933 3602 -3881
rect -658 -3981 -602 -3980
rect -520 -3981 -464 -3979
rect -5189 -4128 -5177 -4070
rect -5119 -4071 -4082 -4070
rect -5119 -4128 -4149 -4071
rect -5189 -4130 -4149 -4128
rect -4090 -4130 -4082 -4071
rect -2593 -4064 -1679 -4006
rect -673 -3989 -437 -3981
rect 749 -3987 941 -3975
rect 1323 -3989 1405 -3975
rect 1807 -3950 1884 -3937
rect 2199 -3950 2276 -3939
rect -673 -3990 -520 -3989
rect -673 -4046 -658 -3990
rect -602 -4045 -520 -3990
rect -464 -4045 -437 -3989
rect 1807 -4006 1818 -3950
rect 1874 -3951 2276 -3950
rect 1874 -4005 2213 -3951
rect 2267 -4005 2276 -3951
rect 1874 -4006 2276 -4005
rect 1807 -4025 1884 -4006
rect 2199 -4017 2276 -4006
rect 3520 -3991 3533 -3933
rect 3591 -3991 3602 -3933
rect 5487 -3897 5498 -3881
rect 5554 -3842 5956 -3841
rect 5554 -3896 5889 -3842
rect 5943 -3896 5956 -3842
rect 5554 -3897 5956 -3896
rect 3520 -4017 3602 -3991
rect 4806 -3950 4883 -3939
rect 5198 -3950 5275 -3937
rect 4806 -3951 5208 -3950
rect 4806 -4005 4815 -3951
rect 4869 -4005 5208 -3951
rect 4806 -4006 5208 -4005
rect 5264 -4006 5275 -3950
rect 4806 -4017 4883 -4006
rect 5198 -4025 5275 -4006
rect 5487 -3951 5956 -3897
rect 5487 -4007 5498 -3951
rect 5554 -3952 5956 -3951
rect 5554 -4006 5893 -3952
rect 5947 -4006 5956 -3952
rect 5554 -4007 5956 -4006
rect 5487 -4027 5564 -4007
rect 5876 -4018 5956 -4007
rect 7084 -3976 7162 -3964
rect 7744 -3976 7933 -3963
rect 7084 -3977 7753 -3976
rect -602 -4046 -437 -4045
rect -673 -4057 -437 -4046
rect 7084 -4031 7096 -3977
rect 7150 -4031 7753 -3977
rect 7084 -4032 7753 -4031
rect 7809 -4032 7863 -3976
rect 7919 -4032 7933 -3976
rect -2593 -4123 -1746 -4064
rect -1687 -4123 -1679 -4064
rect -2593 -4127 -1679 -4123
rect -5189 -4134 -4082 -4130
rect -5189 -4135 -5107 -4134
rect -4159 -4143 -4082 -4134
rect -1756 -4136 -1679 -4127
rect 1103 -4084 1180 -4072
rect 5244 -4084 5322 -4083
rect 1103 -4085 5322 -4084
rect 1103 -4139 1115 -4085
rect 1169 -4099 5322 -4085
rect 1169 -4139 5253 -4099
rect 1103 -4140 5253 -4139
rect -5055 -4209 -4960 -4199
rect -5055 -4265 -5030 -4209
rect -4974 -4224 -4960 -4209
rect -2620 -4200 -2525 -4190
rect -2620 -4224 -2595 -4200
rect -4974 -4256 -2595 -4224
rect -2539 -4256 -2525 -4200
rect 1103 -4195 1180 -4140
rect -4974 -4265 -2525 -4256
rect -5055 -4310 -2525 -4265
rect -5055 -4319 -2595 -4310
rect -5055 -4375 -5030 -4319
rect -4974 -4344 -2595 -4319
rect -4974 -4375 -4960 -4344
rect -5055 -4385 -4960 -4375
rect -2620 -4366 -2595 -4344
rect -2539 -4366 -2525 -4310
rect 7 -4223 86 -4207
rect 7 -4277 19 -4223
rect 73 -4277 86 -4223
rect 1103 -4249 1115 -4195
rect 1169 -4249 1180 -4195
rect 1103 -4263 1180 -4249
rect 5244 -4155 5253 -4140
rect 5309 -4155 5322 -4099
rect 5244 -4202 5322 -4155
rect 7084 -4086 7933 -4032
rect 7084 -4087 7753 -4086
rect 7084 -4141 7096 -4087
rect 7150 -4141 7753 -4087
rect 7084 -4142 7753 -4141
rect 7809 -4142 7863 -4086
rect 7919 -4142 7933 -4086
rect 7084 -4175 7933 -4142
rect 7084 -4197 7162 -4175
rect 5244 -4209 5324 -4202
rect 5244 -4265 5253 -4209
rect 5309 -4265 5324 -4209
rect 5244 -4276 5324 -4265
rect 7084 -4251 7096 -4197
rect 7150 -4251 7162 -4197
rect 7084 -4268 7162 -4251
rect 7744 -4196 7933 -4175
rect 7744 -4252 7753 -4196
rect 7809 -4252 7863 -4196
rect 7919 -4252 7933 -4196
rect 7744 -4267 7933 -4252
rect -2620 -4376 -2525 -4366
rect -340 -4336 -151 -4324
rect 7 -4333 86 -4277
rect 7 -4336 19 -4333
rect -340 -4396 -331 -4336
rect -271 -4396 -218 -4336
rect -158 -4387 19 -4336
rect 73 -4336 86 -4333
rect 5412 -4336 5484 -4329
rect 73 -4343 5484 -4336
rect 73 -4387 5419 -4343
rect -158 -4396 5419 -4387
rect -340 -4408 -79 -4396
rect 7 -4399 86 -4396
rect 5412 -4397 5419 -4396
rect 5473 -4397 5484 -4343
rect -139 -4513 -79 -4408
rect 5412 -4453 5484 -4397
rect -5306 -4573 -79 -4513
rect 991 -4512 1180 -4500
rect 991 -4566 1004 -4512
rect 1058 -4566 1114 -4512
rect 1168 -4514 1180 -4512
rect 5412 -4507 5419 -4453
rect 5473 -4507 5484 -4453
rect 1168 -4566 3535 -4514
rect 5412 -4522 5484 -4507
rect 991 -4570 3535 -4566
rect 991 -4579 1180 -4570
rect 2625 -4832 2717 -4822
rect 1715 -4837 2403 -4833
rect 2625 -4837 2645 -4832
rect 1715 -4891 2337 -4837
rect 2391 -4888 2645 -4837
rect 2701 -4837 2717 -4832
rect 2952 -4837 3037 -4835
rect 2701 -4845 3349 -4837
rect 2701 -4888 2966 -4845
rect 2391 -4891 2966 -4888
rect 1715 -4901 2966 -4891
rect 3022 -4848 3349 -4845
rect 3022 -4901 3283 -4848
rect 1715 -4904 3283 -4901
rect 3339 -4904 3349 -4848
rect 1715 -4906 3349 -4904
rect -1209 -5050 867 -4988
rect -1209 -5106 -1189 -5050
rect -1133 -5106 -1079 -5050
rect -1023 -5106 -969 -5050
rect -913 -5106 -859 -5050
rect -803 -5106 -749 -5050
rect -693 -5106 -639 -5050
rect -583 -5106 86 -5050
rect 142 -5106 196 -5050
rect 252 -5106 306 -5050
rect 362 -5106 416 -5050
rect 472 -5106 526 -5050
rect 582 -5106 636 -5050
rect 692 -5106 746 -5050
rect 802 -5106 867 -5050
rect -1209 -5165 867 -5106
rect 1715 -5337 1795 -4906
rect 2371 -4916 3349 -4906
rect 2371 -4917 3325 -4916
rect 3479 -5297 3535 -4570
rect 4708 -4828 5408 -4827
rect 3732 -4842 3813 -4834
rect 4044 -4842 4125 -4828
rect 4364 -4842 4445 -4830
rect 4683 -4842 5408 -4828
rect 3732 -4843 5408 -4842
rect 3732 -4846 4377 -4843
rect 3732 -4848 4057 -4846
rect 3732 -4904 3745 -4848
rect 3801 -4898 4057 -4848
rect 3801 -4904 3813 -4898
rect 3732 -4920 3813 -4904
rect 4044 -4902 4057 -4898
rect 4113 -4898 4377 -4846
rect 4113 -4902 4125 -4898
rect 4044 -4914 4125 -4902
rect 4364 -4899 4377 -4898
rect 4433 -4897 4699 -4843
rect 4753 -4897 5408 -4843
rect 4433 -4898 5408 -4897
rect 4433 -4899 4445 -4898
rect 4364 -4916 4445 -4899
rect 4683 -4909 5408 -4898
rect 4708 -4929 5408 -4909
rect 1715 -5392 1728 -5337
rect 1783 -5392 1795 -5337
rect 1715 -5447 1795 -5392
rect 1715 -5502 1728 -5447
rect 1783 -5502 1795 -5447
rect 3470 -5310 3543 -5297
rect 3470 -5364 3480 -5310
rect 3534 -5364 3543 -5310
rect 3470 -5420 3543 -5364
rect 3470 -5474 3480 -5420
rect 3534 -5474 3543 -5420
rect 3470 -5493 3543 -5474
rect 5321 -5342 5408 -4929
rect 5321 -5398 5335 -5342
rect 5391 -5398 5408 -5342
rect 5321 -5452 5408 -5398
rect 1715 -5504 1795 -5502
rect -5235 -5518 -5162 -5506
rect 5321 -5508 5335 -5452
rect 5391 -5508 5408 -5452
rect 5321 -5515 5408 -5508
rect -5235 -5575 -5225 -5518
rect -5168 -5575 -2149 -5518
rect -5235 -5628 -2149 -5575
rect -5235 -5685 -5225 -5628
rect -5168 -5632 -2149 -5628
rect -5168 -5685 -5162 -5632
rect -5235 -5697 -5162 -5685
rect -5044 -5778 -4949 -5768
rect -5044 -5834 -5019 -5778
rect -4963 -5824 -4949 -5778
rect -2626 -5782 -2531 -5772
rect -2626 -5824 -2601 -5782
rect -4963 -5834 -2601 -5824
rect -5044 -5838 -2601 -5834
rect -2545 -5838 -2531 -5782
rect -5044 -5888 -2531 -5838
rect -5044 -5944 -5019 -5888
rect -4963 -5892 -2531 -5888
rect -4963 -5944 -2601 -5892
rect -5044 -5954 -4949 -5944
rect -2626 -5948 -2601 -5944
rect -2545 -5948 -2531 -5892
rect -2626 -5958 -2531 -5948
rect -4159 -6038 -4082 -6029
rect -2263 -6031 -2149 -5632
rect -97 -5646 -16 -5642
rect -97 -5703 -85 -5646
rect -28 -5703 -16 -5646
rect -97 -5704 -16 -5703
rect -97 -5756 7176 -5704
rect -97 -5813 -85 -5756
rect -28 -5810 7108 -5756
rect 7162 -5810 7176 -5756
rect -28 -5813 7176 -5810
rect -97 -5823 -16 -5813
rect 7085 -5866 7176 -5813
rect 7085 -5920 7108 -5866
rect 7162 -5920 7176 -5866
rect 7085 -5944 7176 -5920
rect -1756 -6031 -1679 -6022
rect -5128 -6042 -4082 -6038
rect -5128 -6049 -4149 -6042
rect -5128 -6106 -5119 -6049
rect -5062 -6101 -4149 -6049
rect -4090 -6101 -4082 -6042
rect -5062 -6106 -4082 -6101
rect -5128 -6159 -4082 -6106
rect -2593 -6035 -1679 -6031
rect -2593 -6094 -1746 -6035
rect -1687 -6094 -1679 -6035
rect -3038 -6109 -2982 -6107
rect -2908 -6109 -2852 -6107
rect -5128 -6216 -5119 -6159
rect -5062 -6213 -4145 -6159
rect -4091 -6213 -4082 -6159
rect -3046 -6117 -2840 -6109
rect -3046 -6173 -3038 -6117
rect -2982 -6173 -2908 -6117
rect -2852 -6173 -2840 -6117
rect -3046 -6184 -2840 -6173
rect -2593 -6152 -1679 -6094
rect -80 -6041 124 -6026
rect -80 -6047 57 -6041
rect -633 -6102 -577 -6100
rect -508 -6102 -452 -6100
rect -5062 -6214 -4082 -6213
rect -5062 -6216 -5035 -6214
rect -5128 -6228 -5051 -6216
rect -4159 -6225 -4082 -6214
rect -2981 -7364 -2867 -6184
rect -2593 -6206 -1742 -6152
rect -1688 -6206 -1679 -6152
rect -641 -6110 -437 -6102
rect -641 -6166 -633 -6110
rect -577 -6166 -508 -6110
rect -452 -6166 -437 -6110
rect -641 -6177 -437 -6166
rect -80 -6103 -61 -6047
rect -5 -6097 57 -6047
rect 113 -6071 124 -6041
rect 439 -6040 516 -6028
rect 439 -6071 448 -6040
rect 113 -6096 448 -6071
rect 504 -6096 516 -6040
rect 113 -6097 516 -6096
rect -5 -6103 516 -6097
rect -80 -6150 516 -6103
rect -80 -6157 58 -6150
rect -2593 -6207 -1679 -6206
rect -1756 -6218 -1679 -6207
rect -574 -6986 -460 -6177
rect -80 -6213 -61 -6157
rect -5 -6206 58 -6157
rect 114 -6151 516 -6150
rect 114 -6205 453 -6151
rect 507 -6205 516 -6151
rect 114 -6206 516 -6205
rect -5 -6213 124 -6206
rect -80 -6220 124 -6213
rect 439 -6217 516 -6206
rect 2943 -6041 3070 -6034
rect 2943 -6095 3002 -6041
rect 3056 -6095 3070 -6041
rect 2943 -6150 3070 -6095
rect 3573 -6040 3697 -6028
rect 4021 -6033 4077 -6031
rect 3573 -6096 3631 -6040
rect 3687 -6073 3697 -6040
rect 4012 -6041 4089 -6033
rect 4012 -6073 4021 -6041
rect 3687 -6096 4021 -6073
rect 3573 -6097 4021 -6096
rect 4077 -6097 4089 -6041
rect 3385 -6150 3462 -6131
rect 2943 -6151 3395 -6150
rect 2943 -6205 3002 -6151
rect 3056 -6205 3395 -6151
rect 2943 -6206 3395 -6205
rect 3451 -6206 3462 -6150
rect 2943 -6217 3070 -6206
rect 2943 -6564 3059 -6217
rect 3385 -6219 3462 -6206
rect 3573 -6150 4089 -6097
rect 3573 -6206 3631 -6150
rect 3687 -6151 4089 -6150
rect 3687 -6205 4026 -6151
rect 4080 -6205 4089 -6151
rect 3687 -6206 4089 -6205
rect 3573 -6219 3697 -6206
rect 4012 -6217 4089 -6206
rect 6673 -6042 6750 -6030
rect 6673 -6096 6682 -6042
rect 6736 -6096 6750 -6042
rect 6673 -6151 6750 -6096
rect 7066 -6132 7143 -6130
rect 7017 -6151 7143 -6132
rect 6673 -6152 7075 -6151
rect 6673 -6206 6682 -6152
rect 6736 -6206 7075 -6152
rect 6673 -6207 7075 -6206
rect 7131 -6207 7143 -6151
rect 6673 -6218 6750 -6207
rect -315 -6592 3059 -6564
rect -315 -6648 -300 -6592
rect -244 -6593 3059 -6592
rect -244 -6594 -84 -6593
rect -244 -6648 -189 -6594
rect -315 -6650 -189 -6648
rect -133 -6649 -84 -6594
rect -28 -6649 3059 -6593
rect -133 -6650 3059 -6649
rect -315 -6680 3059 -6650
rect 3573 -6986 3687 -6219
rect -574 -7100 3687 -6986
rect 7017 -6261 7143 -6207
rect 7017 -6317 7075 -6261
rect 7131 -6317 7143 -6261
rect 7017 -6334 7143 -6317
rect 7017 -7364 7142 -6334
rect -2981 -7478 7142 -7364
rect 7505 -7458 7678 -7441
rect 7505 -7514 7509 -7458
rect 7565 -7514 7619 -7458
rect 7675 -7514 7678 -7458
rect 7505 -7568 7678 -7514
rect 7505 -7572 7509 -7568
rect 6445 -7624 7509 -7572
rect 7565 -7624 7619 -7568
rect 7675 -7624 7678 -7568
rect 6445 -7633 7678 -7624
rect 6445 -7685 6507 -7633
rect 6561 -7685 6627 -7633
rect 6681 -7685 6747 -7633
rect 6801 -7685 6867 -7633
rect 6921 -7685 6987 -7633
rect 7041 -7678 7678 -7633
rect 7041 -7685 7509 -7678
rect 6445 -7734 7509 -7685
rect 7565 -7734 7619 -7678
rect 7675 -7734 7678 -7678
rect 6445 -7746 7678 -7734
<< via2 >>
rect -159 1599 -103 1655
rect -40 1597 16 1653
rect 67 1597 123 1653
rect -47 1150 9 1206
rect 57 1154 58 1210
rect 58 1154 113 1210
rect -47 1045 9 1101
rect 58 1044 114 1100
rect -3039 -1014 -2983 -958
rect -2921 -1015 -2865 -959
rect -621 -1006 -565 -950
rect -502 -1006 -446 -950
rect -3040 -4053 -2984 -3997
rect -2919 -4053 -2863 -3997
rect -658 -4046 -602 -3990
rect -520 -4045 -464 -3989
rect -61 -6103 -5 -6047
rect 57 -6097 113 -6041
rect -61 -6213 -5 -6157
rect 58 -6206 114 -6150
rect -300 -6648 -244 -6592
rect -189 -6650 -133 -6594
rect -84 -6649 -28 -6593
<< metal3 >>
rect -2973 1655 138 1684
rect -2973 1599 -159 1655
rect -103 1653 138 1655
rect -103 1599 -40 1653
rect -2973 1597 -40 1599
rect 16 1597 67 1653
rect 123 1597 138 1653
rect -2973 1568 138 1597
rect -2973 -948 -2857 1568
rect -59 1210 129 1223
rect -59 1207 57 1210
rect -609 1206 57 1207
rect -609 1150 -47 1206
rect 9 1154 57 1206
rect 113 1154 129 1210
rect 9 1150 129 1154
rect -609 1101 129 1150
rect -609 1063 -47 1101
rect -609 -942 -465 1063
rect -59 1045 -47 1063
rect 9 1100 129 1101
rect 9 1045 58 1100
rect -59 1044 58 1045
rect 114 1044 129 1100
rect -59 1028 129 1044
rect -3049 -958 -2839 -948
rect -630 -950 -436 -942
rect -3049 -1014 -3039 -958
rect -2983 -959 -2839 -958
rect -2983 -1014 -2921 -959
rect -3049 -1015 -2921 -1014
rect -2865 -1015 -2839 -959
rect -631 -1006 -621 -950
rect -565 -1006 -502 -950
rect -446 -1006 -436 -950
rect -3049 -1025 -2839 -1015
rect -630 -1017 -436 -1006
rect -3050 -3997 -2840 -3988
rect -3050 -4053 -3040 -3997
rect -2984 -4053 -2919 -3997
rect -2863 -4053 -2840 -3997
rect -3050 -4063 -2840 -4053
rect -673 -3989 -437 -3981
rect -673 -3990 -520 -3989
rect -673 -4046 -658 -3990
rect -602 -4045 -520 -3990
rect -464 -4045 -437 -3989
rect -602 -4046 -437 -4045
rect -673 -4057 -437 -4046
rect -2998 -6564 -2882 -4063
rect -612 -6038 -454 -4057
rect -80 -6038 124 -6026
rect -612 -6041 124 -6038
rect -612 -6047 57 -6041
rect -612 -6103 -61 -6047
rect -5 -6097 57 -6047
rect 113 -6097 124 -6041
rect -5 -6103 124 -6097
rect -612 -6150 124 -6103
rect -612 -6157 58 -6150
rect -612 -6196 -61 -6157
rect -80 -6213 -61 -6196
rect -5 -6206 58 -6157
rect 114 -6206 124 -6150
rect -5 -6213 124 -6206
rect -80 -6220 124 -6213
rect -2998 -6592 -15 -6564
rect -2998 -6648 -300 -6592
rect -244 -6593 -15 -6592
rect -244 -6594 -84 -6593
rect -244 -6648 -189 -6594
rect -2998 -6650 -189 -6648
rect -133 -6649 -84 -6594
rect -28 -6649 -15 -6593
rect -133 -6650 -15 -6649
rect -2998 -6680 -15 -6650
<< labels >>
flabel metal1 -249 -4375 -249 -4375 0 FreeSans 800 0 0 0 S2
port 33 nsew
flabel via1 -286 -2051 -286 -2051 0 FreeSans 800 0 0 0 S1
port 34 nsew
flabel metal1 -62 -890 -62 -890 0 FreeSans 800 0 0 0 S0
port 3 nsew
flabel metal1 7779 -1906 7779 -1906 0 FreeSans 1120 0 0 0 Vout
port 36 nsew
flabel metal1 5373 2647 5373 2647 0 FreeSans 1600 0 0 0 VDD
port 38 nsew
flabel metal1 7170 -5116 7170 -5116 0 FreeSans 1600 0 0 0 VSS
port 40 nsew
flabel metal1 -5348 -6192 -5348 -6192 0 FreeSans 480 0 0 0 A5
port 29 nsew
flabel metal1 -5362 -5551 -5362 -5551 0 FreeSans 480 0 0 0 A1
port 30 nsew
flabel metal1 -5266 -3998 -5266 -3998 0 FreeSans 480 0 0 0 A3
port 43 nsew
flabel metal1 -5266 1147 -5266 1147 0 FreeSans 480 0 0 0 A6
port 27 nsew
flabel metal1 -5320 626 -5320 626 0 FreeSans 480 0 0 0 A2
port 26 nsew
flabel metal1 -5235 -1468 -5235 -1468 0 FreeSans 480 0 0 0 A4
port 28 nsew
flabel metal1 -5242 -3352 -5242 -3352 0 FreeSans 480 0 0 0 A7
port 45 nsew
flabel metal1 -5245 -994 -5245 -994 0 FreeSans 480 0 0 0 A0
port 6 nsew
flabel metal1 -5011 -24 -5010 -23 0 FreeSans 1600 0 0 0 ENA
port 47 nsew
flabel metal1 -2940 -4010 -2940 -4010 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_1.B
flabel nsubdiffcont -3722 -2511 -3722 -2511 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_1.VDD
flabel psubdiffcont -3731 -5090 -3731 -5090 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_1.VSS
flabel metal2 -4973 -4035 -4973 -4035 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_1.A
flabel metal1 -5002 -4208 -5002 -4208 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_1.CLK
flabel metal1 -2940 -6162 -2940 -6162 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_2.B
flabel nsubdiffcont -3722 -7661 -3722 -7661 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_2.VDD
flabel psubdiffcont -3731 -5082 -3731 -5082 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_2.VSS
flabel metal2 -4973 -6137 -4973 -6137 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_2.A
flabel metal1 -5002 -5964 -5002 -5964 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_2.CLK
flabel metal1 -537 -6155 -537 -6155 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_4.B
flabel nsubdiffcont -1319 -7654 -1319 -7654 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_4.VDD
flabel psubdiffcont -1328 -5075 -1328 -5075 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_4.VSS
flabel metal2 -2570 -6130 -2570 -6130 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_4.A
flabel metal1 -2599 -5957 -2599 -5957 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_4.CLK
flabel metal1 -537 -4003 -537 -4003 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_5.B
flabel nsubdiffcont -1319 -2504 -1319 -2504 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_5.VDD
flabel psubdiffcont -1328 -5083 -1328 -5083 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_5.VSS
flabel metal2 -2570 -4028 -2570 -4028 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_5.A
flabel metal1 -2599 -4201 -2599 -4201 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_5.CLK
flabel metal1 1658 -6154 1658 -6154 0 FreeSans 800 0 0 0 TG_magic_4.B
flabel nsubdiffcont 876 -7653 876 -7653 0 FreeSans 800 0 0 0 TG_magic_4.VDD
flabel psubdiffcont 867 -5074 867 -5074 0 FreeSans 800 0 0 0 TG_magic_4.VSS
flabel metal1 72 -5914 72 -5914 0 FreeSans 800 0 0 0 TG_magic_4.CLK
flabel metal1 44 -6159 44 -6159 0 FreeSans 800 0 0 0 TG_magic_4.A
flabel metal1 1851 -6154 1851 -6154 0 FreeSans 800 0 0 0 TG_magic_1.B
flabel nsubdiffcont 2633 -7653 2633 -7653 0 FreeSans 800 0 0 0 TG_magic_1.VDD
flabel psubdiffcont 2642 -5074 2642 -5074 0 FreeSans 800 0 0 0 TG_magic_1.VSS
flabel metal1 3437 -5914 3437 -5914 0 FreeSans 800 0 0 0 TG_magic_1.CLK
flabel metal1 3465 -6159 3465 -6159 0 FreeSans 800 0 0 0 TG_magic_1.A
flabel metal1 5231 -6154 5231 -6154 0 FreeSans 800 0 0 0 TG_magic_2.B
flabel nsubdiffcont 4449 -7653 4449 -7653 0 FreeSans 800 0 0 0 TG_magic_2.VDD
flabel psubdiffcont 4440 -5074 4440 -5074 0 FreeSans 800 0 0 0 TG_magic_2.VSS
flabel metal1 3645 -5914 3645 -5914 0 FreeSans 800 0 0 0 TG_magic_2.CLK
flabel metal1 3617 -6159 3617 -6159 0 FreeSans 800 0 0 0 TG_magic_2.A
flabel metal1 3664 -4002 3664 -4002 0 FreeSans 800 0 0 0 TG_magic_7.B
flabel nsubdiffcont 4446 -2503 4446 -2503 0 FreeSans 800 0 0 0 TG_magic_7.VDD
flabel psubdiffcont 4455 -5082 4455 -5082 0 FreeSans 800 0 0 0 TG_magic_7.VSS
flabel metal1 5250 -4242 5250 -4242 0 FreeSans 800 0 0 0 TG_magic_7.CLK
flabel metal1 5278 -3997 5278 -3997 0 FreeSans 800 0 0 0 TG_magic_7.A
flabel metal1 3418 -4002 3418 -4002 0 FreeSans 800 0 0 0 TG_magic_9.B
flabel nsubdiffcont 2636 -2503 2636 -2503 0 FreeSans 800 0 0 0 TG_magic_9.VDD
flabel psubdiffcont 2627 -5082 2627 -5082 0 FreeSans 800 0 0 0 TG_magic_9.VSS
flabel metal1 1832 -4242 1832 -4242 0 FreeSans 800 0 0 0 TG_magic_9.CLK
flabel metal1 1804 -3997 1804 -3997 0 FreeSans 800 0 0 0 TG_magic_9.A
flabel metal1 7098 -4003 7098 -4003 0 FreeSans 800 0 0 0 TG_magic_12.B
flabel nsubdiffcont 6316 -2504 6316 -2504 0 FreeSans 800 0 0 0 TG_magic_12.VDD
flabel psubdiffcont 6307 -5083 6307 -5083 0 FreeSans 800 0 0 0 TG_magic_12.VSS
flabel metal1 5512 -4243 5512 -4243 0 FreeSans 800 0 0 0 TG_magic_12.CLK
flabel metal1 5484 -3998 5484 -3998 0 FreeSans 800 0 0 0 TG_magic_12.A
flabel metal1 5531 -6155 5531 -6155 0 FreeSans 800 0 0 0 TG_magic_13.B
flabel nsubdiffcont 6313 -7654 6313 -7654 0 FreeSans 800 0 0 0 TG_magic_13.VDD
flabel psubdiffcont 6322 -5075 6322 -5075 0 FreeSans 800 0 0 0 TG_magic_13.VSS
flabel metal1 7117 -5915 7117 -5915 0 FreeSans 800 0 0 0 TG_magic_13.CLK
flabel metal1 7145 -6160 7145 -6160 0 FreeSans 800 0 0 0 TG_magic_13.A
flabel metal1 -2940 -1002 -2940 -1002 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_0.B
flabel nsubdiffcont -3722 -2501 -3722 -2501 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_0.VDD
flabel psubdiffcont -3731 78 -3731 78 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_0.VSS
flabel metal2 -4973 -977 -4973 -977 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_0.A
flabel metal1 -5002 -804 -5002 -804 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_0.CLK
flabel metal1 -537 -995 -537 -995 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_6.B
flabel nsubdiffcont -1319 -2494 -1319 -2494 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_6.VDD
flabel psubdiffcont -1328 85 -1328 85 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_6.VSS
flabel metal2 -2570 -970 -2570 -970 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_6.A
flabel metal1 -2599 -797 -2599 -797 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_6.CLK
flabel nsubdiffcont 495 -3074 495 -3074 0 FreeSans 800 0 0 0 INVERTER_MUX_1.VDD
flabel psubdiffcont 486 -4555 489 -4552 0 FreeSans 800 0 0 0 INVERTER_MUX_1.VSS
flabel metal1 88 -3954 88 -3954 0 FreeSans 800 0 0 0 INVERTER_MUX_1.IN
flabel metal1 912 -3948 912 -3948 0 FreeSans 800 0 0 0 INVERTER_MUX_1.OUT
flabel nsubdiffcont 495 -3074 495 -3074 0 FreeSans 800 0 0 0 INVERTER_MUX_2.VDD
flabel psubdiffcont 486 -1596 489 -1593 0 FreeSans 800 0 0 0 INVERTER_MUX_2.VSS
flabel metal1 88 -2194 88 -2194 0 FreeSans 800 0 0 0 INVERTER_MUX_2.IN
flabel metal1 912 -2200 912 -2200 0 FreeSans 800 0 0 0 INVERTER_MUX_2.OUT
flabel metal1 3418 -994 3418 -994 0 FreeSans 800 0 0 0 TG_magic_0.B
flabel nsubdiffcont 2636 -2493 2636 -2493 0 FreeSans 800 0 0 0 TG_magic_0.VDD
flabel psubdiffcont 2627 86 2627 86 0 FreeSans 800 0 0 0 TG_magic_0.VSS
flabel metal1 1832 -754 1832 -754 0 FreeSans 800 0 0 0 TG_magic_0.CLK
flabel metal1 1804 -999 1804 -999 0 FreeSans 800 0 0 0 TG_magic_0.A
flabel metal1 3664 -994 3664 -994 0 FreeSans 800 0 0 0 TG_magic_5.B
flabel nsubdiffcont 4446 -2493 4446 -2493 0 FreeSans 800 0 0 0 TG_magic_5.VDD
flabel psubdiffcont 4455 86 4455 86 0 FreeSans 800 0 0 0 TG_magic_5.VSS
flabel metal1 5250 -754 5250 -754 0 FreeSans 800 0 0 0 TG_magic_5.CLK
flabel metal1 5278 -999 5278 -999 0 FreeSans 800 0 0 0 TG_magic_5.A
flabel metal1 7098 -995 7098 -995 0 FreeSans 800 0 0 0 TG_magic_8.B
flabel nsubdiffcont 6316 -2494 6316 -2494 0 FreeSans 800 0 0 0 TG_magic_8.VDD
flabel psubdiffcont 6307 85 6307 85 0 FreeSans 800 0 0 0 TG_magic_8.VSS
flabel metal1 5512 -755 5512 -755 0 FreeSans 800 0 0 0 TG_magic_8.CLK
flabel metal1 5484 -1000 5484 -1000 0 FreeSans 800 0 0 0 TG_magic_8.A
flabel metal1 -2940 1150 -2940 1150 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_3.B
flabel nsubdiffcont -3722 2649 -3722 2649 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_3.VDD
flabel psubdiffcont -3731 70 -3731 70 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_3.VSS
flabel metal2 -4973 1125 -4973 1125 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_3.A
flabel metal1 -5002 952 -5002 952 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_3.CLK
flabel metal1 -537 1157 -537 1157 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_7.B
flabel nsubdiffcont -1319 2656 -1319 2656 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_7.VDD
flabel psubdiffcont -1328 77 -1328 77 0 FreeSans 800 0 0 0 TG_GATE_SWITCH_magic_7.VSS
flabel metal2 -2570 1132 -2570 1132 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_7.A
flabel metal1 -2599 959 -2599 959 0 FreeSans 1600 0 0 0 TG_GATE_SWITCH_magic_7.CLK
flabel nsubdiffcont 495 -133 495 -133 0 FreeSans 800 0 0 0 INVERTER_MUX_0.VDD
flabel psubdiffcont 486 -1614 489 -1611 0 FreeSans 800 0 0 0 INVERTER_MUX_0.VSS
flabel metal1 88 -1013 88 -1013 0 FreeSans 800 0 0 0 INVERTER_MUX_0.IN
flabel metal1 912 -1007 912 -1007 0 FreeSans 800 0 0 0 INVERTER_MUX_0.OUT
flabel metal1 1658 1158 1658 1158 0 FreeSans 800 0 0 0 TG_magic_10.B
flabel nsubdiffcont 876 2657 876 2657 0 FreeSans 800 0 0 0 TG_magic_10.VDD
flabel psubdiffcont 867 78 867 78 0 FreeSans 800 0 0 0 TG_magic_10.VSS
flabel metal1 72 918 72 918 0 FreeSans 800 0 0 0 TG_magic_10.CLK
flabel metal1 44 1163 44 1163 0 FreeSans 800 0 0 0 TG_magic_10.A
flabel metal1 1851 1158 1851 1158 0 FreeSans 800 0 0 0 TG_magic_6.B
flabel nsubdiffcont 2633 2657 2633 2657 0 FreeSans 800 0 0 0 TG_magic_6.VDD
flabel psubdiffcont 2642 78 2642 78 0 FreeSans 800 0 0 0 TG_magic_6.VSS
flabel metal1 3437 918 3437 918 0 FreeSans 800 0 0 0 TG_magic_6.CLK
flabel metal1 3465 1163 3465 1163 0 FreeSans 800 0 0 0 TG_magic_6.A
flabel metal1 5231 1158 5231 1158 0 FreeSans 800 0 0 0 TG_magic_11.B
flabel nsubdiffcont 4449 2657 4449 2657 0 FreeSans 800 0 0 0 TG_magic_11.VDD
flabel psubdiffcont 4440 78 4440 78 0 FreeSans 800 0 0 0 TG_magic_11.VSS
flabel metal1 3645 918 3645 918 0 FreeSans 800 0 0 0 TG_magic_11.CLK
flabel metal1 3617 1163 3617 1163 0 FreeSans 800 0 0 0 TG_magic_11.A
flabel metal1 5531 1157 5531 1157 0 FreeSans 800 0 0 0 TG_magic_3.B
flabel nsubdiffcont 6313 2656 6313 2656 0 FreeSans 800 0 0 0 TG_magic_3.VDD
flabel psubdiffcont 6322 77 6322 77 0 FreeSans 800 0 0 0 TG_magic_3.VSS
flabel metal1 7117 917 7117 917 0 FreeSans 800 0 0 0 TG_magic_3.CLK
flabel metal1 7145 1162 7145 1162 0 FreeSans 800 0 0 0 TG_magic_3.A
<< end >>
