magic
tech gf180mcuC
magscale 1 10
timestamp 1692077799
<< nwell >>
rect 418 310 1302 828
<< pwell >>
rect 0 0 1720 236
<< nmos >>
rect 112 68 168 168
rect 272 68 328 168
rect 432 68 488 168
rect 592 68 648 168
rect 752 68 808 168
rect 912 68 968 168
rect 1072 68 1128 168
rect 1232 68 1288 168
rect 1392 68 1448 168
rect 1552 68 1608 168
<< pmos >>
rect 592 440 648 640
rect 752 440 808 640
rect 912 440 968 640
rect 1072 440 1128 640
<< ndiff >>
rect 24 155 112 168
rect 24 81 37 155
rect 83 81 112 155
rect 24 68 112 81
rect 168 155 272 168
rect 168 81 197 155
rect 243 81 272 155
rect 168 68 272 81
rect 328 155 432 168
rect 328 81 357 155
rect 403 81 432 155
rect 328 68 432 81
rect 488 155 592 168
rect 488 81 517 155
rect 563 81 592 155
rect 488 68 592 81
rect 648 155 752 168
rect 648 81 677 155
rect 723 81 752 155
rect 648 68 752 81
rect 808 155 912 168
rect 808 81 837 155
rect 883 81 912 155
rect 808 68 912 81
rect 968 155 1072 168
rect 968 81 997 155
rect 1043 81 1072 155
rect 968 68 1072 81
rect 1128 155 1232 168
rect 1128 81 1157 155
rect 1203 81 1232 155
rect 1128 68 1232 81
rect 1288 155 1392 168
rect 1288 81 1317 155
rect 1363 81 1392 155
rect 1288 68 1392 81
rect 1448 155 1552 168
rect 1448 81 1477 155
rect 1523 81 1552 155
rect 1448 68 1552 81
rect 1608 155 1696 168
rect 1608 81 1637 155
rect 1683 81 1696 155
rect 1608 68 1696 81
<< pdiff >>
rect 504 627 592 640
rect 504 453 517 627
rect 563 453 592 627
rect 504 440 592 453
rect 648 627 752 640
rect 648 453 677 627
rect 723 453 752 627
rect 648 440 752 453
rect 808 627 912 640
rect 808 453 837 627
rect 883 453 912 627
rect 808 440 912 453
rect 968 627 1072 640
rect 968 453 997 627
rect 1043 453 1072 627
rect 968 440 1072 453
rect 1128 627 1216 640
rect 1128 453 1157 627
rect 1203 453 1216 627
rect 1128 440 1216 453
<< ndiffc >>
rect 37 81 83 155
rect 197 81 243 155
rect 357 81 403 155
rect 517 81 563 155
rect 677 81 723 155
rect 837 81 883 155
rect 997 81 1043 155
rect 1157 81 1203 155
rect 1317 81 1363 155
rect 1477 81 1523 155
rect 1637 81 1683 155
<< pdiffc >>
rect 517 453 563 627
rect 677 453 723 627
rect 837 453 883 627
rect 997 453 1043 627
rect 1157 453 1203 627
<< psubdiff >>
rect 24 -228 1695 -215
rect 24 -274 37 -228
rect 83 -274 131 -228
rect 177 -274 225 -228
rect 271 -274 319 -228
rect 365 -274 413 -228
rect 459 -274 507 -228
rect 553 -274 601 -228
rect 647 -274 695 -228
rect 741 -274 789 -228
rect 835 -274 883 -228
rect 929 -274 977 -228
rect 1023 -274 1071 -228
rect 1117 -274 1165 -228
rect 1211 -274 1259 -228
rect 1305 -274 1353 -228
rect 1399 -274 1447 -228
rect 1493 -274 1541 -228
rect 1587 -274 1635 -228
rect 1681 -274 1695 -228
rect 24 -287 1695 -274
<< nsubdiff >>
rect 448 782 1272 795
rect 448 736 461 782
rect 507 736 555 782
rect 601 736 649 782
rect 695 736 743 782
rect 789 736 837 782
rect 883 736 931 782
rect 977 736 1025 782
rect 1071 736 1119 782
rect 1165 736 1213 782
rect 1259 736 1272 782
rect 448 723 1272 736
<< psubdiffcont >>
rect 37 -274 83 -228
rect 131 -274 177 -228
rect 225 -274 271 -228
rect 319 -274 365 -228
rect 413 -274 459 -228
rect 507 -274 553 -228
rect 601 -274 647 -228
rect 695 -274 741 -228
rect 789 -274 835 -228
rect 883 -274 929 -228
rect 977 -274 1023 -228
rect 1071 -274 1117 -228
rect 1165 -274 1211 -228
rect 1259 -274 1305 -228
rect 1353 -274 1399 -228
rect 1447 -274 1493 -228
rect 1541 -274 1587 -228
rect 1635 -274 1681 -228
<< nsubdiffcont >>
rect 461 736 507 782
rect 555 736 601 782
rect 649 736 695 782
rect 743 736 789 782
rect 837 736 883 782
rect 931 736 977 782
rect 1025 736 1071 782
rect 1119 736 1165 782
rect 1213 736 1259 782
<< polysilicon >>
rect 592 640 648 684
rect 752 640 808 684
rect 912 640 968 684
rect 1072 640 1128 684
rect 279 396 357 405
rect 592 396 648 440
rect 279 392 648 396
rect 279 345 292 392
rect 339 345 648 392
rect 279 340 648 345
rect 279 332 357 340
rect 112 168 168 212
rect 272 168 328 212
rect 432 168 488 340
rect 592 168 648 212
rect 752 168 808 440
rect 912 316 968 440
rect 1072 420 1128 440
rect 1072 385 1608 420
rect 1072 364 1303 385
rect 1290 339 1303 364
rect 1349 364 1608 385
rect 1349 339 1362 364
rect 1290 326 1362 339
rect 912 260 1128 316
rect 912 168 968 212
rect 1072 168 1128 260
rect 1232 168 1288 212
rect 1392 168 1448 212
rect 1552 168 1608 364
rect 112 48 168 68
rect 272 48 328 68
rect 432 48 488 68
rect 112 -8 488 48
rect 592 48 648 68
rect 752 48 808 68
rect 912 48 968 68
rect 592 -8 968 48
rect 1072 48 1128 68
rect 1232 48 1288 68
rect 1392 48 1448 68
rect 1072 -8 1448 48
rect 1552 24 1608 68
rect 573 -82 647 -73
rect 695 -82 751 -8
rect 573 -86 751 -82
rect 573 -138 586 -86
rect 634 -138 751 -86
rect 1392 -55 1448 -8
rect 1599 -55 1672 -46
rect 1392 -59 1672 -55
rect 1392 -106 1612 -59
rect 1659 -106 1672 -59
rect 1392 -111 1672 -106
rect 1599 -119 1672 -111
rect 573 -151 647 -138
<< polycontact >>
rect 292 345 339 392
rect 1303 339 1349 385
rect 586 -138 634 -86
rect 1612 -106 1659 -59
<< metal1 >>
rect 418 782 1302 815
rect 418 736 461 782
rect 507 736 555 782
rect 601 736 649 782
rect 695 736 743 782
rect 789 736 837 782
rect 883 736 931 782
rect 977 736 1025 782
rect 1071 736 1119 782
rect 1165 736 1213 782
rect 1259 736 1302 782
rect 418 703 1302 736
rect 675 638 721 703
rect 517 627 563 638
rect 675 627 723 638
rect 675 609 677 627
rect 279 396 350 403
rect 199 392 350 396
rect 199 345 292 392
rect 339 345 350 392
rect 199 340 350 345
rect 279 334 350 340
rect 517 385 563 453
rect 677 442 723 453
rect 837 627 883 638
rect 837 385 883 453
rect 997 627 1043 703
rect 997 442 1043 453
rect 1157 627 1203 638
rect 1203 453 1783 488
rect 1157 442 1783 453
rect 1292 385 1360 396
rect 517 339 1303 385
rect 1349 339 1360 385
rect 517 258 563 339
rect 1292 328 1360 339
rect 37 212 563 258
rect 677 212 1363 258
rect 37 155 83 212
rect 37 70 83 81
rect 197 155 243 166
rect 197 24 243 81
rect 357 155 403 212
rect 357 70 403 81
rect 517 155 563 166
rect 517 24 563 81
rect 677 155 723 212
rect 677 70 723 81
rect 837 155 883 166
rect 837 24 883 81
rect 997 155 1043 212
rect 997 70 1043 81
rect 1157 155 1203 166
rect 197 -22 883 24
rect 585 -85 645 -75
rect 483 -86 645 -85
rect 483 -138 586 -86
rect 634 -138 645 -86
rect 483 -141 645 -138
rect 585 -149 645 -141
rect 1157 -195 1203 81
rect 1317 155 1363 212
rect 1317 70 1363 81
rect 1477 155 1523 166
rect 1477 -195 1523 81
rect 1637 155 1683 442
rect 1637 70 1683 81
rect 1601 -56 1659 -48
rect 1601 -59 1780 -56
rect 1601 -106 1612 -59
rect 1659 -106 1780 -59
rect 1601 -112 1780 -106
rect 1601 -117 1659 -112
rect 4 -228 1715 -195
rect 4 -274 37 -228
rect 83 -274 131 -228
rect 177 -274 225 -228
rect 271 -274 319 -228
rect 365 -274 413 -228
rect 459 -274 507 -228
rect 553 -274 601 -228
rect 647 -274 695 -228
rect 741 -274 789 -228
rect 835 -274 883 -228
rect 929 -274 977 -228
rect 1023 -274 1071 -228
rect 1117 -274 1165 -228
rect 1211 -274 1259 -228
rect 1305 -274 1353 -228
rect 1399 -274 1447 -228
rect 1493 -274 1541 -228
rect 1587 -274 1635 -228
rect 1681 -274 1715 -228
rect 4 -307 1715 -274
<< labels >>
flabel metal1 493 -115 493 -115 0 FreeSans 320 0 0 0 B
port 2 nsew
flabel metal1 1760 462 1760 462 0 FreeSans 320 0 0 0 OUT
port 5 nsew
flabel nsubdiffcont 860 759 860 759 0 FreeSans 320 0 0 0 VDD
port 6 nsew
flabel psubdiff 858 -251 858 -251 0 FreeSans 320 0 0 0 VSS
port 8 nsew
flabel metal1 1770 -86 1770 -86 0 FreeSans 320 180 0 0 C
port 3 nsew
flabel metal1 213 362 213 362 0 FreeSans 320 0 0 0 A
port 1 nsew
<< end >>
