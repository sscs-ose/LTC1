magic
tech gf180mcuC
magscale 1 10
timestamp 1695119997
<< metal1 >>
rect 2619 2592 2695 2594
rect 508 2584 2696 2592
rect 508 2525 519 2584
rect 571 2545 2629 2584
rect 571 2525 583 2545
rect 508 2512 583 2525
rect 2619 2531 2629 2545
rect 2687 2545 2696 2584
rect 2687 2531 2695 2545
rect 2619 2514 2695 2531
rect 342 2508 414 2509
rect -156 2466 414 2508
rect -156 2358 838 2466
rect 343 2357 838 2358
rect 1183 2357 1969 2466
rect 2437 2462 2534 2464
rect 2902 2462 2983 2588
rect 2437 2452 2983 2462
rect 2437 2386 2454 2452
rect 2516 2386 2983 2452
rect 2437 2381 2983 2386
rect 2437 2378 2534 2381
rect 1813 2314 1969 2357
rect 1813 2299 3723 2314
rect 508 2268 583 2276
rect 508 2209 518 2268
rect 570 2209 583 2268
rect 508 2200 583 2209
rect 386 2078 458 2089
rect 386 2062 396 2078
rect -347 1996 -30 2043
rect 264 2020 396 2062
rect 448 2020 458 2078
rect 264 2007 458 2020
rect 386 2006 458 2007
rect 524 1948 571 2200
rect 1813 2187 3636 2299
rect 3709 2187 3723 2299
rect 1813 2166 3723 2187
rect 1165 2014 1214 2015
rect 317 1901 571 1948
rect 647 1953 864 2000
rect 1165 1967 1918 2014
rect 1165 1966 1214 1967
rect -285 1699 -198 1710
rect -285 1634 -277 1699
rect -211 1634 -198 1699
rect -285 1620 -198 1634
rect 460 1702 530 1710
rect 460 1630 469 1702
rect 522 1684 530 1702
rect 647 1684 694 1953
rect 1326 1917 1412 1919
rect 1181 1904 1412 1917
rect 1181 1860 1337 1904
rect 1326 1845 1337 1860
rect 1397 1845 1412 1904
rect 1326 1831 1412 1845
rect 1863 1814 1918 1967
rect 2379 1824 2673 1871
rect 522 1637 694 1684
rect 1862 1759 2101 1814
rect 522 1630 530 1637
rect 460 1620 530 1630
rect 1862 1567 1917 1759
rect 2477 1747 2545 1748
rect 2474 1730 2545 1747
rect 2626 1734 2673 1824
rect 2474 1669 2484 1730
rect 2539 1669 2545 1730
rect 2474 1653 2545 1669
rect 2618 1733 2673 1734
rect 2748 1774 2959 1823
rect 3459 1811 3540 1821
rect 3283 1810 3828 1811
rect 2618 1720 2697 1733
rect 2618 1668 2628 1720
rect 2685 1668 2697 1720
rect 2618 1652 2697 1668
rect 1855 1555 1918 1567
rect 1855 1503 1862 1555
rect 1914 1503 1918 1555
rect 1855 1490 1918 1503
rect 275 1475 415 1476
rect 14 1370 416 1475
rect 2574 1466 2635 1487
rect 757 1417 897 1418
rect 734 1370 1299 1417
rect 2574 1404 2579 1466
rect 2631 1404 2635 1466
rect 2574 1388 2635 1404
rect -364 1305 2504 1370
rect -364 1254 2447 1305
rect -365 1231 2447 1254
rect -365 1175 2504 1231
rect -365 1140 897 1175
rect -365 1138 -280 1140
rect -2 1139 897 1140
rect 532 1134 897 1139
rect 639 1133 897 1134
rect 2586 904 2632 1388
rect 2748 966 2808 1774
rect 3283 1763 3469 1810
rect 3459 1754 3469 1763
rect 3528 1763 3828 1810
rect 3528 1754 3540 1763
rect 3459 1745 3540 1754
rect 2857 1724 2930 1727
rect 2857 1672 2873 1724
rect 2928 1672 2930 1724
rect 2857 1667 2930 1672
rect 2863 1309 3426 1381
rect 2863 1232 2886 1309
rect 2974 1232 3426 1309
rect 2863 1074 3426 1232
rect 612 882 692 888
rect 612 844 626 882
rect 680 879 692 882
rect 484 814 626 844
rect 682 818 692 879
rect 1322 858 1410 870
rect 1322 837 1339 858
rect 680 814 692 818
rect 484 787 692 814
rect 612 786 692 787
rect 1194 800 1339 837
rect 1397 800 1410 858
rect 2484 845 2632 904
rect 2725 954 2823 966
rect 2725 881 2744 954
rect 2812 881 2823 954
rect 2725 865 2823 881
rect 1194 780 1410 800
rect 1322 778 1410 780
rect 1480 764 1568 779
rect -133 704 136 751
rect 827 740 859 741
rect -133 554 -86 704
rect 430 685 859 740
rect 1480 732 1492 764
rect 827 683 859 685
rect 1147 690 1492 732
rect 1554 732 1568 764
rect 1983 763 2089 810
rect 1983 735 2030 763
rect 2383 743 2631 798
rect 1554 690 1618 732
rect 1147 682 1618 690
rect 1945 682 2030 735
rect 2577 692 2631 743
rect 3336 786 3468 787
rect 3599 786 3809 787
rect 3336 785 3809 786
rect 3336 731 3338 785
rect 3394 731 3809 785
rect 3394 728 3430 731
rect 1147 677 1576 682
rect 2577 645 2995 692
rect 3458 663 3540 674
rect 3458 662 3474 663
rect 2577 560 2630 645
rect 3279 611 3474 662
rect 3526 611 3540 663
rect 3279 606 3540 611
rect 3459 598 3540 606
rect -141 542 -63 554
rect -141 490 -126 542
rect -72 490 -63 542
rect -141 477 -63 490
rect 2562 544 2638 560
rect 2562 490 2577 544
rect 2630 490 2638 544
rect 2562 477 2638 490
rect -264 373 3788 381
rect -265 336 3788 373
rect -265 212 3629 336
rect 3710 212 3788 336
rect -265 154 3788 212
rect -265 146 3787 154
<< via1 >>
rect 519 2525 571 2584
rect 2629 2531 2687 2584
rect 2454 2386 2516 2452
rect 518 2209 570 2268
rect 396 2020 448 2078
rect 3636 2187 3709 2299
rect -277 1634 -211 1699
rect 469 1630 522 1702
rect 1337 1845 1397 1904
rect 2484 1669 2539 1730
rect 2628 1668 2685 1720
rect 1862 1503 1914 1555
rect 2579 1404 2631 1466
rect 2447 1231 2514 1305
rect 3469 1754 3528 1810
rect 2873 1672 2928 1724
rect 2886 1232 2974 1309
rect 626 879 680 882
rect 626 818 682 879
rect 626 814 680 818
rect 1339 800 1397 858
rect 2744 881 2812 954
rect 1492 690 1554 764
rect 3338 728 3394 785
rect 3474 611 3526 663
rect -126 490 -72 542
rect 2577 490 2630 544
rect 3629 212 3710 336
<< metal2 >>
rect 508 2584 583 2592
rect 508 2525 519 2584
rect 571 2525 583 2584
rect 508 2268 583 2525
rect 2618 2584 2697 2592
rect 2618 2531 2629 2584
rect 2687 2531 2697 2584
rect 2437 2459 2534 2464
rect 508 2209 518 2268
rect 570 2209 583 2268
rect 508 2200 583 2209
rect 1329 2452 2534 2459
rect 1329 2386 2454 2452
rect 2516 2386 2534 2452
rect 1329 2379 2534 2386
rect 388 2078 692 2086
rect 388 2020 396 2078
rect 448 2020 692 2078
rect 388 2007 692 2020
rect -285 1702 530 1710
rect -285 1699 469 1702
rect -285 1634 -277 1699
rect -211 1634 469 1699
rect -285 1630 469 1634
rect 522 1630 530 1702
rect -285 1620 530 1630
rect 613 882 692 2007
rect 1329 1918 1409 2379
rect 2437 2378 2534 2379
rect 613 814 626 882
rect 680 879 692 882
rect 682 818 692 879
rect 1328 1904 1411 1918
rect 1328 1845 1337 1904
rect 1397 1845 1411 1904
rect 1328 870 1411 1845
rect 2477 1747 2545 1748
rect 2466 1741 2545 1747
rect 680 814 692 818
rect 613 788 692 814
rect 1322 858 1411 870
rect 1322 800 1339 858
rect 1397 800 1411 858
rect 1322 784 1411 800
rect 1483 1730 2545 1741
rect 1483 1669 2484 1730
rect 2539 1669 2545 1730
rect 1483 1658 2545 1669
rect 1322 778 1410 784
rect 1483 764 1566 1658
rect 2466 1653 2545 1658
rect 2618 1733 2697 2531
rect 3621 2299 3723 2314
rect 3621 2187 3636 2299
rect 3709 2187 3723 2299
rect 3459 1810 3540 1821
rect 3459 1754 3469 1810
rect 3528 1754 3540 1810
rect 3459 1745 3540 1754
rect 2618 1724 2945 1733
rect 2618 1720 2873 1724
rect 2618 1668 2628 1720
rect 2685 1672 2873 1720
rect 2928 1672 2945 1724
rect 2685 1668 2945 1672
rect 2466 1652 2526 1653
rect 2618 1652 2945 1668
rect 1855 1563 1917 1567
rect 1855 1555 2635 1563
rect 1855 1503 1862 1555
rect 1914 1503 2635 1555
rect 1855 1493 2635 1503
rect 1855 1491 1918 1493
rect 2574 1466 2635 1493
rect 2574 1404 2579 1466
rect 2631 1404 2635 1466
rect 2574 1386 2635 1404
rect 2864 1330 3003 1333
rect 2432 1309 3003 1330
rect 2432 1305 2886 1309
rect 2432 1231 2447 1305
rect 2514 1232 2886 1305
rect 2974 1232 3003 1309
rect 2514 1231 3003 1232
rect 2432 1213 3003 1231
rect 1483 690 1492 764
rect 1554 690 1566 764
rect 2711 954 2827 972
rect 2711 881 2744 954
rect 2812 881 2827 954
rect 2711 812 2827 881
rect 2711 785 3402 812
rect 2711 728 3338 785
rect 3394 728 3402 785
rect 2711 698 3402 728
rect 2711 696 3320 698
rect 1483 682 1566 690
rect 3470 674 3534 1745
rect 3458 663 3540 674
rect 3458 611 3474 663
rect 3526 611 3540 663
rect 3458 606 3540 611
rect 3459 598 3540 606
rect -141 542 -63 554
rect -141 490 -126 542
rect -72 541 -63 542
rect 2563 544 2638 560
rect 2563 541 2577 544
rect -72 490 2577 541
rect 2630 490 2638 544
rect -141 481 2638 490
rect -141 477 -63 481
rect 2563 477 2638 481
rect 3621 336 3723 2187
rect 3621 212 3629 336
rect 3710 212 3723 336
rect 3621 146 3723 212
use inv  inv_0
timestamp 1695119997
transform 1 0 1629 0 1 236
box -61 58 345 1028
use inv_my_mag  inv_my_mag_0
timestamp 1695119997
transform 1 0 1629 0 1 236
box -61 58 345 1028
use nand2  nand2_0
timestamp 1694691991
transform 1 0 799 0 -1 2278
box -70 -188 502 863
use nand2  nand2_1
timestamp 1694691991
transform 1 0 2032 0 1 485
box -70 -188 502 863
use nand2  nand2_2
timestamp 1694691991
transform 1 0 79 0 1 426
box -70 -188 502 863
use nand2  nand2_3
timestamp 1694691991
transform 1 0 796 0 1 419
box -70 -188 502 863
use nand2  nand2_4
timestamp 1694691991
transform 1 0 2928 0 1 367
box -70 -188 502 863
use nand2  nand2_5
timestamp 1694691991
transform 1 0 2028 0 -1 2088
box -70 -188 502 863
use nand2  nand2_6
timestamp 1694691991
transform -1 0 3364 0 -1 2088
box -70 -188 502 863
use nand2  nand2_7
timestamp 1694691991
transform 1 0 -87 0 -1 2321
box -70 -188 502 863
<< labels >>
flabel metal1 -330 2030 -330 2030 0 FreeSans 480 0 0 0 D
port 1 nsew
flabel metal1 -300 1210 -300 1210 0 FreeSans 480 0 0 0 VDD
port 3 nsew
flabel metal1 3440 220 3440 220 0 FreeSans 480 0 0 0 VSS
port 4 nsew
flabel metal1 2943 2541 2943 2541 0 FreeSans 480 0 0 0 RST
port 7 nsew
flabel via1 -244 1667 -244 1667 0 FreeSans 480 0 0 0 CLK
port 8 nsew
flabel metal1 3801 1790 3801 1790 0 FreeSans 480 0 0 0 Q
port 9 nsew
flabel metal1 3782 760 3782 760 0 FreeSans 480 0 0 0 QB
port 10 nsew
<< end >>
