magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2079 -4959 2921 2525
<< nwell >>
rect 0 364 892 525
<< psubdiff >>
rect 179 -2894 680 -2873
rect 179 -2895 415 -2894
rect 179 -2941 251 -2895
rect 297 -2940 415 -2895
rect 461 -2895 680 -2894
rect 461 -2940 535 -2895
rect 297 -2941 535 -2940
rect 581 -2941 680 -2895
rect 179 -2959 680 -2941
<< nsubdiff >>
rect 316 483 633 500
rect 316 437 358 483
rect 404 437 465 483
rect 511 437 569 483
rect 615 437 633 483
rect 316 422 633 437
<< psubdiffcont >>
rect 251 -2941 297 -2895
rect 415 -2940 461 -2894
rect 535 -2941 581 -2895
<< nsubdiffcont >>
rect 358 437 404 483
rect 465 437 511 483
rect 569 437 615 483
<< polysilicon >>
rect 174 -86 286 16
rect 390 -86 502 16
rect 606 -86 718 16
rect 174 -570 286 -398
rect 390 -570 502 -398
rect 606 -570 718 -398
rect 174 -1054 286 -882
rect 390 -1054 502 -882
rect 606 -1054 718 -882
rect 174 -1538 286 -1366
rect 390 -1538 502 -1366
rect 606 -1404 718 -1366
rect 578 -1439 718 -1404
rect 578 -1485 611 -1439
rect 657 -1485 718 -1439
rect 578 -1510 718 -1485
rect 606 -1538 718 -1510
rect 174 -2022 286 -1850
rect 390 -1890 502 -1850
rect 361 -1916 502 -1890
rect 361 -1962 400 -1916
rect 446 -1962 502 -1916
rect 361 -1984 502 -1962
rect 390 -2022 502 -1984
rect 606 -2022 718 -1850
rect 174 -2377 286 -2332
rect 172 -2390 286 -2377
rect 172 -2436 187 -2390
rect 233 -2436 286 -2390
rect 172 -2464 286 -2436
rect 390 -2464 502 -2331
rect 606 -2464 718 -2332
rect 174 -2465 286 -2464
<< polycontact >>
rect 611 -1485 657 -1439
rect 400 -1962 446 -1916
rect 187 -2436 233 -2390
<< metal1 >>
rect 71 483 741 500
rect 71 437 358 483
rect 404 437 465 483
rect 511 437 569 483
rect 615 437 741 483
rect 71 422 741 437
rect -40 -1431 41 -1421
rect -79 -1438 41 -1431
rect -79 -1490 -25 -1438
rect 27 -1490 41 -1438
rect -79 -1497 41 -1490
rect -40 -1507 41 -1497
rect -54 -1913 50 -1902
rect -54 -1965 -15 -1913
rect 37 -1965 50 -1913
rect -54 -1973 50 -1965
rect 99 -2288 145 422
rect 315 -1691 361 282
rect 531 -1202 577 282
rect 433 -1203 577 -1202
rect 218 -1741 361 -1691
rect 423 -1252 577 -1203
rect 423 -1681 477 -1252
rect 531 -1320 577 -1252
rect 747 -1167 793 282
rect 747 -1255 921 -1167
rect 588 -1435 679 -1419
rect 588 -1487 607 -1435
rect 659 -1487 679 -1435
rect 588 -1507 679 -1487
rect 531 -1681 577 -1584
rect 423 -1731 577 -1681
rect 218 -2173 267 -1741
rect 315 -1804 361 -1741
rect 379 -1912 465 -1894
rect 379 -1964 396 -1912
rect 448 -1964 465 -1912
rect 379 -1982 465 -1964
rect 315 -2173 361 -2068
rect 218 -2223 361 -2173
rect 315 -2288 361 -2223
rect 531 -2288 577 -1731
rect 174 -2388 246 -2377
rect 128 -2390 246 -2388
rect 128 -2436 187 -2390
rect 233 -2436 246 -2390
rect 747 -2417 793 -1255
rect 128 -2437 246 -2436
rect 174 -2448 246 -2437
rect 315 -2464 793 -2417
rect 99 -2777 145 -2510
rect 315 -2730 361 -2464
rect 531 -2777 577 -2510
rect 747 -2730 793 -2464
rect 99 -2823 577 -2777
rect 99 -2874 145 -2823
rect 332 -2874 680 -2873
rect 76 -2894 821 -2874
rect 76 -2895 415 -2894
rect 76 -2941 251 -2895
rect 297 -2940 415 -2895
rect 461 -2895 821 -2894
rect 461 -2940 535 -2895
rect 297 -2941 535 -2940
rect 581 -2941 821 -2895
rect 76 -2959 821 -2941
<< via1 >>
rect -25 -1490 27 -1438
rect -15 -1965 37 -1913
rect 607 -1439 659 -1435
rect 607 -1485 611 -1439
rect 611 -1485 657 -1439
rect 657 -1485 659 -1439
rect 607 -1487 659 -1485
rect 396 -1916 448 -1912
rect 396 -1962 400 -1916
rect 400 -1962 446 -1916
rect 446 -1962 448 -1916
rect 396 -1964 448 -1962
<< metal2 >>
rect -40 -1427 41 -1421
rect 588 -1427 679 -1419
rect -40 -1435 679 -1427
rect -40 -1438 607 -1435
rect -40 -1490 -25 -1438
rect 27 -1487 607 -1438
rect 659 -1487 679 -1435
rect 27 -1490 679 -1487
rect -40 -1498 679 -1490
rect -40 -1499 367 -1498
rect -40 -1507 41 -1499
rect 588 -1507 679 -1498
rect 379 -1902 465 -1894
rect -28 -1912 465 -1902
rect -28 -1913 396 -1912
rect -28 -1965 -15 -1913
rect 37 -1964 396 -1913
rect 448 -1964 465 -1912
rect 37 -1965 465 -1964
rect -28 -1973 465 -1965
rect 379 -1982 465 -1973
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_0
timestamp 1713185578
transform 1 0 230 0 1 -2620
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_1
timestamp 1713185578
transform 1 0 446 0 1 -2620
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_2
timestamp 1713185578
transform 1 0 662 0 1 -2620
box -168 -180 168 180
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_0
timestamp 1713185578
transform 1 0 662 0 1 -2178
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_1
timestamp 1713185578
transform 1 0 230 0 1 -2178
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_2
timestamp 1713185578
transform 1 0 446 0 1 -2178
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_3
timestamp 1713185578
transform 1 0 662 0 1 -1210
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_4
timestamp 1713185578
transform 1 0 446 0 1 -1210
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_5
timestamp 1713185578
transform 1 0 230 0 1 -1210
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_6
timestamp 1713185578
transform 1 0 230 0 1 -1694
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_7
timestamp 1713185578
transform 1 0 446 0 1 -1694
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_8
timestamp 1713185578
transform 1 0 662 0 1 -1694
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_9
timestamp 1713185578
transform 1 0 230 0 1 -726
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_10
timestamp 1713185578
transform 1 0 446 0 1 -726
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_11
timestamp 1713185578
transform 1 0 662 0 1 -726
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_12
timestamp 1713185578
transform 1 0 230 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_13
timestamp 1713185578
transform 1 0 446 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_14
timestamp 1713185578
transform 1 0 662 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_15
timestamp 1713185578
transform 1 0 662 0 1 172
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_16
timestamp 1713185578
transform 1 0 446 0 1 172
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_17
timestamp 1713185578
transform 1 0 230 0 1 172
box -230 -242 230 242
<< labels >>
flabel nsubdiffcont 382 462 382 462 0 FreeSans 750 0 0 0 VDD
flabel psubdiffcont 438 -2917 438 -2917 0 FreeSans 750 0 0 0 VSS
flabel metal1 s 144 -2414 144 -2414 0 FreeSans 750 0 0 0 A
port 1 nsew
flabel metal1 s -50 -1942 -50 -1942 0 FreeSans 750 0 0 0 B
port 2 nsew
flabel metal1 s -64 -1470 -64 -1470 0 FreeSans 750 0 0 0 C
port 3 nsew
flabel metal1 s 882 -1219 882 -1219 0 FreeSans 750 0 0 0 VOUT
port 4 nsew
<< end >>
