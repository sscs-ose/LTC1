magic
tech gf180mcuC
magscale 1 10
timestamp 1714562775
<< nwell >>
rect -55208 23853 56994 26259
rect 42596 16872 42621 16920
rect 32263 15615 32288 15663
rect 42484 9484 42514 9533
rect 42549 9113 42618 9393
rect 32153 8241 32176 8290
rect 12548 7418 12843 7429
rect 12394 7364 12849 7418
rect 12394 7284 12854 7364
rect 12399 7230 12854 7284
rect 16000 163 18007 966
rect 20198 872 20535 1341
rect 49364 -2053 50681 -1322
rect -5034 -4592 -4812 -4205
rect -3927 -4592 -3705 -4205
rect 30742 -6464 31342 -6437
rect 30367 -6647 31342 -6464
rect 30742 -6768 31342 -6647
rect 49417 -6744 50748 -6013
rect 51686 -16258 52943 -15579
rect 11508 -19432 11706 -19109
rect 12748 -19430 12933 -19109
rect 8294 -21029 8626 -20953
rect 5973 -21454 6890 -21380
rect -2958 -22110 -2779 -22057
rect -2958 -22114 -2788 -22110
rect -2764 -22114 -2751 -22079
rect -2958 -22362 -1818 -22114
rect -2958 -22365 -2450 -22362
rect -1858 -22365 -1818 -22362
rect -2958 -22453 -1818 -22365
<< pwell >>
rect 12625 -11234 12862 -11042
rect 13033 -11425 13601 -11231
rect 3933 -23198 4327 -22962
rect -157 -23989 120 -23772
<< psubdiff >>
rect 9554 -1908 22354 -1669
rect 9486 -15322 44085 -14251
rect -55858 -29624 54839 -29479
rect -55858 -29952 -55497 -29624
rect -55172 -29952 -55002 -29624
rect -54677 -29952 -54507 -29624
rect -54182 -29952 -54012 -29624
rect -53687 -29952 -53517 -29624
rect -53192 -29952 -53022 -29624
rect -52697 -29952 -52527 -29624
rect -52202 -29952 -52032 -29624
rect -51707 -29952 -51537 -29624
rect -51212 -29952 -51042 -29624
rect -50717 -29952 -50547 -29624
rect -50222 -29952 -50052 -29624
rect -49727 -29952 -49557 -29624
rect -49232 -29952 -49062 -29624
rect -48737 -29952 -48567 -29624
rect -48242 -29952 -48072 -29624
rect -47747 -29952 -47577 -29624
rect -47252 -29952 -47082 -29624
rect -46757 -29952 -46587 -29624
rect -46262 -29952 -46092 -29624
rect -45767 -29952 -45597 -29624
rect -45272 -29952 -45102 -29624
rect -44777 -29952 -44607 -29624
rect -44282 -29952 -44112 -29624
rect -43787 -29952 -43617 -29624
rect -43292 -29952 -43122 -29624
rect -42797 -29952 -42627 -29624
rect -42302 -29952 -42132 -29624
rect -41807 -29952 -41637 -29624
rect -41312 -29952 -41142 -29624
rect -40817 -29952 -40647 -29624
rect -40322 -29952 -40152 -29624
rect -39827 -29952 -39657 -29624
rect -39332 -29952 -39162 -29624
rect -38837 -29952 -38667 -29624
rect -38342 -29952 -38172 -29624
rect -37847 -29952 -37677 -29624
rect -37352 -29952 -37182 -29624
rect -36857 -29952 -36687 -29624
rect -36362 -29952 -36192 -29624
rect -35867 -29952 -35697 -29624
rect -35372 -29952 -35202 -29624
rect -34877 -29952 -34707 -29624
rect -34382 -29952 -34212 -29624
rect -33887 -29952 -33717 -29624
rect -33392 -29952 -33222 -29624
rect -32897 -29952 -32727 -29624
rect -32402 -29952 -32232 -29624
rect -31907 -29952 -31737 -29624
rect -31412 -29952 -31242 -29624
rect -30917 -29952 -30747 -29624
rect -30422 -29952 -30252 -29624
rect -29927 -29952 -29757 -29624
rect -29432 -29952 -29262 -29624
rect -28937 -29952 -28767 -29624
rect -28442 -29952 -28272 -29624
rect -27947 -29952 -27777 -29624
rect -27452 -29952 -27282 -29624
rect -26957 -29952 -26787 -29624
rect -26462 -29952 -26292 -29624
rect -25967 -29952 -25797 -29624
rect -25472 -29952 -25302 -29624
rect -24977 -29952 -24807 -29624
rect -24482 -29952 -24312 -29624
rect -23987 -29952 -23817 -29624
rect -23492 -29952 -23322 -29624
rect -22997 -29952 -22827 -29624
rect -22502 -29952 -22332 -29624
rect -22007 -29952 -21837 -29624
rect -21512 -29952 -21342 -29624
rect -21017 -29952 -20847 -29624
rect -20522 -29952 -20352 -29624
rect -20027 -29952 -19857 -29624
rect -19532 -29952 -19362 -29624
rect -19037 -29952 -18867 -29624
rect -18542 -29952 -18372 -29624
rect -18047 -29952 -17877 -29624
rect -17552 -29952 -17382 -29624
rect -17057 -29952 -16887 -29624
rect -16562 -29952 -16392 -29624
rect -16067 -29952 -15897 -29624
rect -15572 -29952 -15402 -29624
rect -15077 -29952 -14907 -29624
rect -14582 -29952 -14412 -29624
rect -14087 -29952 -13917 -29624
rect -13592 -29952 -13422 -29624
rect -13097 -29952 -12927 -29624
rect -12602 -29952 -12432 -29624
rect -12107 -29952 -11937 -29624
rect -11612 -29952 -11442 -29624
rect -11117 -29952 -10947 -29624
rect -10622 -29952 -10452 -29624
rect -10127 -29952 -9957 -29624
rect -9632 -29952 -9462 -29624
rect -9137 -29952 -8967 -29624
rect -8642 -29952 -8472 -29624
rect -8147 -29952 -7977 -29624
rect -7652 -29952 -7482 -29624
rect -7157 -29952 -6987 -29624
rect -6662 -29952 -6492 -29624
rect -6167 -29952 -5997 -29624
rect -5672 -29952 -5502 -29624
rect -5177 -29952 -5007 -29624
rect -4682 -29952 -4512 -29624
rect -4187 -29952 -4017 -29624
rect -3692 -29952 -3522 -29624
rect -3197 -29952 -3027 -29624
rect -2702 -29952 -2532 -29624
rect -2207 -29952 -2037 -29624
rect -1712 -29952 -1542 -29624
rect -1217 -29952 -1047 -29624
rect -722 -29952 -552 -29624
rect -227 -29952 -57 -29624
rect 268 -29952 438 -29624
rect 763 -29952 933 -29624
rect 1258 -29952 1428 -29624
rect 1753 -29952 1923 -29624
rect 2248 -29952 2418 -29624
rect 2743 -29952 2913 -29624
rect 3238 -29952 3408 -29624
rect 3733 -29952 3903 -29624
rect 4228 -29952 4398 -29624
rect 4723 -29952 4893 -29624
rect 5218 -29952 5388 -29624
rect 5713 -29952 5883 -29624
rect 6208 -29952 6378 -29624
rect 6703 -29952 6873 -29624
rect 7198 -29952 7368 -29624
rect 7693 -29952 7863 -29624
rect 8188 -29952 8358 -29624
rect 8683 -29952 8853 -29624
rect 9178 -29952 9348 -29624
rect 9673 -29952 9843 -29624
rect 10168 -29952 10338 -29624
rect 10663 -29952 10833 -29624
rect 11158 -29952 11328 -29624
rect 11653 -29952 11823 -29624
rect 12148 -29952 12318 -29624
rect 12643 -29952 12813 -29624
rect 13138 -29952 13308 -29624
rect 13633 -29952 13803 -29624
rect 14128 -29952 14298 -29624
rect 14623 -29952 14793 -29624
rect 15118 -29952 15288 -29624
rect 15613 -29952 15783 -29624
rect 16108 -29952 16278 -29624
rect 16603 -29952 16773 -29624
rect 17098 -29952 17268 -29624
rect 17593 -29952 17763 -29624
rect 18088 -29952 18258 -29624
rect 18583 -29952 18753 -29624
rect 19078 -29952 19248 -29624
rect 19573 -29952 19743 -29624
rect 20068 -29952 20238 -29624
rect 20563 -29952 20733 -29624
rect 21058 -29952 21228 -29624
rect 21553 -29952 21723 -29624
rect 22048 -29952 22218 -29624
rect 22543 -29952 22713 -29624
rect 23038 -29952 23208 -29624
rect 23533 -29952 23703 -29624
rect 24028 -29952 24198 -29624
rect 24523 -29952 24693 -29624
rect 25018 -29952 25188 -29624
rect 25513 -29952 25683 -29624
rect 26008 -29952 26178 -29624
rect 26503 -29952 26673 -29624
rect 26998 -29952 27168 -29624
rect 27493 -29952 27663 -29624
rect 27988 -29952 28158 -29624
rect 28483 -29952 28653 -29624
rect 28978 -29952 29148 -29624
rect 29473 -29952 29643 -29624
rect 29968 -29952 30138 -29624
rect 30463 -29952 30633 -29624
rect 30958 -29952 31128 -29624
rect 31453 -29952 31623 -29624
rect 31948 -29952 32118 -29624
rect 32443 -29952 32613 -29624
rect 32938 -29952 33108 -29624
rect 33433 -29952 33603 -29624
rect 33928 -29952 34098 -29624
rect 34423 -29952 34593 -29624
rect 34918 -29952 35088 -29624
rect 35413 -29952 35583 -29624
rect 35908 -29952 36078 -29624
rect 36403 -29952 36573 -29624
rect 36898 -29952 37068 -29624
rect 37393 -29952 37563 -29624
rect 37888 -29952 38058 -29624
rect 38383 -29952 38553 -29624
rect 38878 -29952 39048 -29624
rect 39373 -29952 39543 -29624
rect 39868 -29952 40038 -29624
rect 40363 -29952 40533 -29624
rect 40858 -29952 41028 -29624
rect 41353 -29952 41523 -29624
rect 41848 -29952 42018 -29624
rect 42343 -29952 42513 -29624
rect 42838 -29952 43008 -29624
rect 43333 -29952 43503 -29624
rect 43828 -29952 43998 -29624
rect 44323 -29952 44493 -29624
rect 44818 -29952 44988 -29624
rect 45313 -29952 45483 -29624
rect 45808 -29952 45978 -29624
rect 46303 -29952 46473 -29624
rect 46798 -29952 46968 -29624
rect 47293 -29952 47463 -29624
rect 47788 -29952 47958 -29624
rect 48283 -29952 48453 -29624
rect 48778 -29952 48948 -29624
rect 49273 -29952 49443 -29624
rect 49768 -29952 49938 -29624
rect 50263 -29952 50433 -29624
rect 50758 -29952 50928 -29624
rect 51253 -29952 51423 -29624
rect 51748 -29952 51918 -29624
rect 52243 -29952 52413 -29624
rect 52738 -29952 52908 -29624
rect 53233 -29952 53403 -29624
rect 53728 -29952 53898 -29624
rect 54223 -29952 54839 -29624
rect -55858 -30100 54839 -29952
rect -55858 -30428 -55497 -30100
rect -55172 -30428 -55002 -30100
rect -54677 -30428 -54507 -30100
rect -54182 -30428 -54012 -30100
rect -53687 -30428 -53517 -30100
rect -53192 -30428 -53022 -30100
rect -52697 -30428 -52527 -30100
rect -52202 -30428 -52032 -30100
rect -51707 -30428 -51537 -30100
rect -51212 -30428 -51042 -30100
rect -50717 -30428 -50547 -30100
rect -50222 -30428 -50052 -30100
rect -49727 -30428 -49557 -30100
rect -49232 -30428 -49062 -30100
rect -48737 -30428 -48567 -30100
rect -48242 -30428 -48072 -30100
rect -47747 -30428 -47577 -30100
rect -47252 -30428 -47082 -30100
rect -46757 -30428 -46587 -30100
rect -46262 -30428 -46092 -30100
rect -45767 -30428 -45597 -30100
rect -45272 -30428 -45102 -30100
rect -44777 -30428 -44607 -30100
rect -44282 -30428 -44112 -30100
rect -43787 -30428 -43617 -30100
rect -43292 -30428 -43122 -30100
rect -42797 -30428 -42627 -30100
rect -42302 -30428 -42132 -30100
rect -41807 -30428 -41637 -30100
rect -41312 -30428 -41142 -30100
rect -40817 -30428 -40647 -30100
rect -40322 -30428 -40152 -30100
rect -39827 -30428 -39657 -30100
rect -39332 -30428 -39162 -30100
rect -38837 -30428 -38667 -30100
rect -38342 -30428 -38172 -30100
rect -37847 -30428 -37677 -30100
rect -37352 -30428 -37182 -30100
rect -36857 -30428 -36687 -30100
rect -36362 -30428 -36192 -30100
rect -35867 -30428 -35697 -30100
rect -35372 -30428 -35202 -30100
rect -34877 -30428 -34707 -30100
rect -34382 -30428 -34212 -30100
rect -33887 -30428 -33717 -30100
rect -33392 -30428 -33222 -30100
rect -32897 -30428 -32727 -30100
rect -32402 -30428 -32232 -30100
rect -31907 -30428 -31737 -30100
rect -31412 -30428 -31242 -30100
rect -30917 -30428 -30747 -30100
rect -30422 -30428 -30252 -30100
rect -29927 -30428 -29757 -30100
rect -29432 -30428 -29262 -30100
rect -28937 -30428 -28767 -30100
rect -28442 -30428 -28272 -30100
rect -27947 -30428 -27777 -30100
rect -27452 -30428 -27282 -30100
rect -26957 -30428 -26787 -30100
rect -26462 -30428 -26292 -30100
rect -25967 -30428 -25797 -30100
rect -25472 -30428 -25302 -30100
rect -24977 -30428 -24807 -30100
rect -24482 -30428 -24312 -30100
rect -23987 -30428 -23817 -30100
rect -23492 -30428 -23322 -30100
rect -22997 -30428 -22827 -30100
rect -22502 -30428 -22332 -30100
rect -22007 -30428 -21837 -30100
rect -21512 -30428 -21342 -30100
rect -21017 -30428 -20847 -30100
rect -20522 -30428 -20352 -30100
rect -20027 -30428 -19857 -30100
rect -19532 -30428 -19362 -30100
rect -19037 -30428 -18867 -30100
rect -18542 -30428 -18372 -30100
rect -18047 -30428 -17877 -30100
rect -17552 -30428 -17382 -30100
rect -17057 -30428 -16887 -30100
rect -16562 -30428 -16392 -30100
rect -16067 -30428 -15897 -30100
rect -15572 -30428 -15402 -30100
rect -15077 -30428 -14907 -30100
rect -14582 -30428 -14412 -30100
rect -14087 -30428 -13917 -30100
rect -13592 -30428 -13422 -30100
rect -13097 -30428 -12927 -30100
rect -12602 -30428 -12432 -30100
rect -12107 -30428 -11937 -30100
rect -11612 -30428 -11442 -30100
rect -11117 -30428 -10947 -30100
rect -10622 -30428 -10452 -30100
rect -10127 -30428 -9957 -30100
rect -9632 -30428 -9462 -30100
rect -9137 -30428 -8967 -30100
rect -8642 -30428 -8472 -30100
rect -8147 -30428 -7977 -30100
rect -7652 -30428 -7482 -30100
rect -7157 -30428 -6987 -30100
rect -6662 -30428 -6492 -30100
rect -6167 -30428 -5997 -30100
rect -5672 -30428 -5502 -30100
rect -5177 -30428 -5007 -30100
rect -4682 -30428 -4512 -30100
rect -4187 -30428 -4017 -30100
rect -3692 -30428 -3522 -30100
rect -3197 -30428 -3027 -30100
rect -2702 -30428 -2532 -30100
rect -2207 -30428 -2037 -30100
rect -1712 -30428 -1542 -30100
rect -1217 -30428 -1047 -30100
rect -722 -30428 -552 -30100
rect -227 -30428 -57 -30100
rect 268 -30428 438 -30100
rect 763 -30428 933 -30100
rect 1258 -30428 1428 -30100
rect 1753 -30428 1923 -30100
rect 2248 -30428 2418 -30100
rect 2743 -30428 2913 -30100
rect 3238 -30428 3408 -30100
rect 3733 -30428 3903 -30100
rect 4228 -30428 4398 -30100
rect 4723 -30428 4893 -30100
rect 5218 -30428 5388 -30100
rect 5713 -30428 5883 -30100
rect 6208 -30428 6378 -30100
rect 6703 -30428 6873 -30100
rect 7198 -30428 7368 -30100
rect 7693 -30428 7863 -30100
rect 8188 -30428 8358 -30100
rect 8683 -30428 8853 -30100
rect 9178 -30428 9348 -30100
rect 9673 -30428 9843 -30100
rect 10168 -30428 10338 -30100
rect 10663 -30428 10833 -30100
rect 11158 -30428 11328 -30100
rect 11653 -30428 11823 -30100
rect 12148 -30428 12318 -30100
rect 12643 -30428 12813 -30100
rect 13138 -30428 13308 -30100
rect 13633 -30428 13803 -30100
rect 14128 -30428 14298 -30100
rect 14623 -30428 14793 -30100
rect 15118 -30428 15288 -30100
rect 15613 -30428 15783 -30100
rect 16108 -30428 16278 -30100
rect 16603 -30428 16773 -30100
rect 17098 -30428 17268 -30100
rect 17593 -30428 17763 -30100
rect 18088 -30428 18258 -30100
rect 18583 -30428 18753 -30100
rect 19078 -30428 19248 -30100
rect 19573 -30428 19743 -30100
rect 20068 -30428 20238 -30100
rect 20563 -30428 20733 -30100
rect 21058 -30428 21228 -30100
rect 21553 -30428 21723 -30100
rect 22048 -30428 22218 -30100
rect 22543 -30428 22713 -30100
rect 23038 -30428 23208 -30100
rect 23533 -30428 23703 -30100
rect 24028 -30428 24198 -30100
rect 24523 -30428 24693 -30100
rect 25018 -30428 25188 -30100
rect 25513 -30428 25683 -30100
rect 26008 -30428 26178 -30100
rect 26503 -30428 26673 -30100
rect 26998 -30428 27168 -30100
rect 27493 -30428 27663 -30100
rect 27988 -30428 28158 -30100
rect 28483 -30428 28653 -30100
rect 28978 -30428 29148 -30100
rect 29473 -30428 29643 -30100
rect 29968 -30428 30138 -30100
rect 30463 -30428 30633 -30100
rect 30958 -30428 31128 -30100
rect 31453 -30428 31623 -30100
rect 31948 -30428 32118 -30100
rect 32443 -30428 32613 -30100
rect 32938 -30428 33108 -30100
rect 33433 -30428 33603 -30100
rect 33928 -30428 34098 -30100
rect 34423 -30428 34593 -30100
rect 34918 -30428 35088 -30100
rect 35413 -30428 35583 -30100
rect 35908 -30428 36078 -30100
rect 36403 -30428 36573 -30100
rect 36898 -30428 37068 -30100
rect 37393 -30428 37563 -30100
rect 37888 -30428 38058 -30100
rect 38383 -30428 38553 -30100
rect 38878 -30428 39048 -30100
rect 39373 -30428 39543 -30100
rect 39868 -30428 40038 -30100
rect 40363 -30428 40533 -30100
rect 40858 -30428 41028 -30100
rect 41353 -30428 41523 -30100
rect 41848 -30428 42018 -30100
rect 42343 -30428 42513 -30100
rect 42838 -30428 43008 -30100
rect 43333 -30428 43503 -30100
rect 43828 -30428 43998 -30100
rect 44323 -30428 44493 -30100
rect 44818 -30428 44988 -30100
rect 45313 -30428 45483 -30100
rect 45808 -30428 45978 -30100
rect 46303 -30428 46473 -30100
rect 46798 -30428 46968 -30100
rect 47293 -30428 47463 -30100
rect 47788 -30428 47958 -30100
rect 48283 -30428 48453 -30100
rect 48778 -30428 48948 -30100
rect 49273 -30428 49443 -30100
rect 49768 -30428 49938 -30100
rect 50263 -30428 50433 -30100
rect 50758 -30428 50928 -30100
rect 51253 -30428 51423 -30100
rect 51748 -30428 51918 -30100
rect 52243 -30428 52413 -30100
rect 52738 -30428 52908 -30100
rect 53233 -30428 53403 -30100
rect 53728 -30428 53898 -30100
rect 54223 -30428 54839 -30100
rect -55858 -30576 54839 -30428
rect -55858 -30904 -55497 -30576
rect -55172 -30904 -55002 -30576
rect -54677 -30904 -54507 -30576
rect -54182 -30904 -54012 -30576
rect -53687 -30904 -53517 -30576
rect -53192 -30904 -53022 -30576
rect -52697 -30904 -52527 -30576
rect -52202 -30904 -52032 -30576
rect -51707 -30904 -51537 -30576
rect -51212 -30904 -51042 -30576
rect -50717 -30904 -50547 -30576
rect -50222 -30904 -50052 -30576
rect -49727 -30904 -49557 -30576
rect -49232 -30904 -49062 -30576
rect -48737 -30904 -48567 -30576
rect -48242 -30904 -48072 -30576
rect -47747 -30904 -47577 -30576
rect -47252 -30904 -47082 -30576
rect -46757 -30904 -46587 -30576
rect -46262 -30904 -46092 -30576
rect -45767 -30904 -45597 -30576
rect -45272 -30904 -45102 -30576
rect -44777 -30904 -44607 -30576
rect -44282 -30904 -44112 -30576
rect -43787 -30904 -43617 -30576
rect -43292 -30904 -43122 -30576
rect -42797 -30904 -42627 -30576
rect -42302 -30904 -42132 -30576
rect -41807 -30904 -41637 -30576
rect -41312 -30904 -41142 -30576
rect -40817 -30904 -40647 -30576
rect -40322 -30904 -40152 -30576
rect -39827 -30904 -39657 -30576
rect -39332 -30904 -39162 -30576
rect -38837 -30904 -38667 -30576
rect -38342 -30904 -38172 -30576
rect -37847 -30904 -37677 -30576
rect -37352 -30904 -37182 -30576
rect -36857 -30904 -36687 -30576
rect -36362 -30904 -36192 -30576
rect -35867 -30904 -35697 -30576
rect -35372 -30904 -35202 -30576
rect -34877 -30904 -34707 -30576
rect -34382 -30904 -34212 -30576
rect -33887 -30904 -33717 -30576
rect -33392 -30904 -33222 -30576
rect -32897 -30904 -32727 -30576
rect -32402 -30904 -32232 -30576
rect -31907 -30904 -31737 -30576
rect -31412 -30904 -31242 -30576
rect -30917 -30904 -30747 -30576
rect -30422 -30904 -30252 -30576
rect -29927 -30904 -29757 -30576
rect -29432 -30904 -29262 -30576
rect -28937 -30904 -28767 -30576
rect -28442 -30904 -28272 -30576
rect -27947 -30904 -27777 -30576
rect -27452 -30904 -27282 -30576
rect -26957 -30904 -26787 -30576
rect -26462 -30904 -26292 -30576
rect -25967 -30904 -25797 -30576
rect -25472 -30904 -25302 -30576
rect -24977 -30904 -24807 -30576
rect -24482 -30904 -24312 -30576
rect -23987 -30904 -23817 -30576
rect -23492 -30904 -23322 -30576
rect -22997 -30904 -22827 -30576
rect -22502 -30904 -22332 -30576
rect -22007 -30904 -21837 -30576
rect -21512 -30904 -21342 -30576
rect -21017 -30904 -20847 -30576
rect -20522 -30904 -20352 -30576
rect -20027 -30904 -19857 -30576
rect -19532 -30904 -19362 -30576
rect -19037 -30904 -18867 -30576
rect -18542 -30904 -18372 -30576
rect -18047 -30904 -17877 -30576
rect -17552 -30904 -17382 -30576
rect -17057 -30904 -16887 -30576
rect -16562 -30904 -16392 -30576
rect -16067 -30904 -15897 -30576
rect -15572 -30904 -15402 -30576
rect -15077 -30904 -14907 -30576
rect -14582 -30904 -14412 -30576
rect -14087 -30904 -13917 -30576
rect -13592 -30904 -13422 -30576
rect -13097 -30904 -12927 -30576
rect -12602 -30904 -12432 -30576
rect -12107 -30904 -11937 -30576
rect -11612 -30904 -11442 -30576
rect -11117 -30904 -10947 -30576
rect -10622 -30904 -10452 -30576
rect -10127 -30904 -9957 -30576
rect -9632 -30904 -9462 -30576
rect -9137 -30904 -8967 -30576
rect -8642 -30904 -8472 -30576
rect -8147 -30904 -7977 -30576
rect -7652 -30904 -7482 -30576
rect -7157 -30904 -6987 -30576
rect -6662 -30904 -6492 -30576
rect -6167 -30904 -5997 -30576
rect -5672 -30904 -5502 -30576
rect -5177 -30904 -5007 -30576
rect -4682 -30904 -4512 -30576
rect -4187 -30904 -4017 -30576
rect -3692 -30904 -3522 -30576
rect -3197 -30904 -3027 -30576
rect -2702 -30904 -2532 -30576
rect -2207 -30904 -2037 -30576
rect -1712 -30904 -1542 -30576
rect -1217 -30904 -1047 -30576
rect -722 -30904 -552 -30576
rect -227 -30904 -57 -30576
rect 268 -30904 438 -30576
rect 763 -30904 933 -30576
rect 1258 -30904 1428 -30576
rect 1753 -30904 1923 -30576
rect 2248 -30904 2418 -30576
rect 2743 -30904 2913 -30576
rect 3238 -30904 3408 -30576
rect 3733 -30904 3903 -30576
rect 4228 -30904 4398 -30576
rect 4723 -30904 4893 -30576
rect 5218 -30904 5388 -30576
rect 5713 -30904 5883 -30576
rect 6208 -30904 6378 -30576
rect 6703 -30904 6873 -30576
rect 7198 -30904 7368 -30576
rect 7693 -30904 7863 -30576
rect 8188 -30904 8358 -30576
rect 8683 -30904 8853 -30576
rect 9178 -30904 9348 -30576
rect 9673 -30904 9843 -30576
rect 10168 -30904 10338 -30576
rect 10663 -30904 10833 -30576
rect 11158 -30904 11328 -30576
rect 11653 -30904 11823 -30576
rect 12148 -30904 12318 -30576
rect 12643 -30904 12813 -30576
rect 13138 -30904 13308 -30576
rect 13633 -30904 13803 -30576
rect 14128 -30904 14298 -30576
rect 14623 -30904 14793 -30576
rect 15118 -30904 15288 -30576
rect 15613 -30904 15783 -30576
rect 16108 -30904 16278 -30576
rect 16603 -30904 16773 -30576
rect 17098 -30904 17268 -30576
rect 17593 -30904 17763 -30576
rect 18088 -30904 18258 -30576
rect 18583 -30904 18753 -30576
rect 19078 -30904 19248 -30576
rect 19573 -30904 19743 -30576
rect 20068 -30904 20238 -30576
rect 20563 -30904 20733 -30576
rect 21058 -30904 21228 -30576
rect 21553 -30904 21723 -30576
rect 22048 -30904 22218 -30576
rect 22543 -30904 22713 -30576
rect 23038 -30904 23208 -30576
rect 23533 -30904 23703 -30576
rect 24028 -30904 24198 -30576
rect 24523 -30904 24693 -30576
rect 25018 -30904 25188 -30576
rect 25513 -30904 25683 -30576
rect 26008 -30904 26178 -30576
rect 26503 -30904 26673 -30576
rect 26998 -30904 27168 -30576
rect 27493 -30904 27663 -30576
rect 27988 -30904 28158 -30576
rect 28483 -30904 28653 -30576
rect 28978 -30904 29148 -30576
rect 29473 -30904 29643 -30576
rect 29968 -30904 30138 -30576
rect 30463 -30904 30633 -30576
rect 30958 -30904 31128 -30576
rect 31453 -30904 31623 -30576
rect 31948 -30904 32118 -30576
rect 32443 -30904 32613 -30576
rect 32938 -30904 33108 -30576
rect 33433 -30904 33603 -30576
rect 33928 -30904 34098 -30576
rect 34423 -30904 34593 -30576
rect 34918 -30904 35088 -30576
rect 35413 -30904 35583 -30576
rect 35908 -30904 36078 -30576
rect 36403 -30904 36573 -30576
rect 36898 -30904 37068 -30576
rect 37393 -30904 37563 -30576
rect 37888 -30904 38058 -30576
rect 38383 -30904 38553 -30576
rect 38878 -30904 39048 -30576
rect 39373 -30904 39543 -30576
rect 39868 -30904 40038 -30576
rect 40363 -30904 40533 -30576
rect 40858 -30904 41028 -30576
rect 41353 -30904 41523 -30576
rect 41848 -30904 42018 -30576
rect 42343 -30904 42513 -30576
rect 42838 -30904 43008 -30576
rect 43333 -30904 43503 -30576
rect 43828 -30904 43998 -30576
rect 44323 -30904 44493 -30576
rect 44818 -30904 44988 -30576
rect 45313 -30904 45483 -30576
rect 45808 -30904 45978 -30576
rect 46303 -30904 46473 -30576
rect 46798 -30904 46968 -30576
rect 47293 -30904 47463 -30576
rect 47788 -30904 47958 -30576
rect 48283 -30904 48453 -30576
rect 48778 -30904 48948 -30576
rect 49273 -30904 49443 -30576
rect 49768 -30904 49938 -30576
rect 50263 -30904 50433 -30576
rect 50758 -30904 50928 -30576
rect 51253 -30904 51423 -30576
rect 51748 -30904 51918 -30576
rect 52243 -30904 52413 -30576
rect 52738 -30904 52908 -30576
rect 53233 -30904 53403 -30576
rect 53728 -30904 53898 -30576
rect 54223 -30904 54839 -30576
rect -55858 -31052 54839 -30904
rect -55858 -31380 -55497 -31052
rect -55172 -31380 -55002 -31052
rect -54677 -31380 -54507 -31052
rect -54182 -31380 -54012 -31052
rect -53687 -31380 -53517 -31052
rect -53192 -31380 -53022 -31052
rect -52697 -31380 -52527 -31052
rect -52202 -31380 -52032 -31052
rect -51707 -31380 -51537 -31052
rect -51212 -31380 -51042 -31052
rect -50717 -31380 -50547 -31052
rect -50222 -31380 -50052 -31052
rect -49727 -31380 -49557 -31052
rect -49232 -31380 -49062 -31052
rect -48737 -31380 -48567 -31052
rect -48242 -31380 -48072 -31052
rect -47747 -31380 -47577 -31052
rect -47252 -31380 -47082 -31052
rect -46757 -31380 -46587 -31052
rect -46262 -31380 -46092 -31052
rect -45767 -31380 -45597 -31052
rect -45272 -31380 -45102 -31052
rect -44777 -31380 -44607 -31052
rect -44282 -31380 -44112 -31052
rect -43787 -31380 -43617 -31052
rect -43292 -31380 -43122 -31052
rect -42797 -31380 -42627 -31052
rect -42302 -31380 -42132 -31052
rect -41807 -31380 -41637 -31052
rect -41312 -31380 -41142 -31052
rect -40817 -31380 -40647 -31052
rect -40322 -31380 -40152 -31052
rect -39827 -31380 -39657 -31052
rect -39332 -31380 -39162 -31052
rect -38837 -31380 -38667 -31052
rect -38342 -31380 -38172 -31052
rect -37847 -31380 -37677 -31052
rect -37352 -31380 -37182 -31052
rect -36857 -31380 -36687 -31052
rect -36362 -31380 -36192 -31052
rect -35867 -31380 -35697 -31052
rect -35372 -31380 -35202 -31052
rect -34877 -31380 -34707 -31052
rect -34382 -31380 -34212 -31052
rect -33887 -31380 -33717 -31052
rect -33392 -31380 -33222 -31052
rect -32897 -31380 -32727 -31052
rect -32402 -31380 -32232 -31052
rect -31907 -31380 -31737 -31052
rect -31412 -31380 -31242 -31052
rect -30917 -31380 -30747 -31052
rect -30422 -31380 -30252 -31052
rect -29927 -31380 -29757 -31052
rect -29432 -31380 -29262 -31052
rect -28937 -31380 -28767 -31052
rect -28442 -31380 -28272 -31052
rect -27947 -31380 -27777 -31052
rect -27452 -31380 -27282 -31052
rect -26957 -31380 -26787 -31052
rect -26462 -31380 -26292 -31052
rect -25967 -31380 -25797 -31052
rect -25472 -31380 -25302 -31052
rect -24977 -31380 -24807 -31052
rect -24482 -31380 -24312 -31052
rect -23987 -31380 -23817 -31052
rect -23492 -31380 -23322 -31052
rect -22997 -31380 -22827 -31052
rect -22502 -31380 -22332 -31052
rect -22007 -31380 -21837 -31052
rect -21512 -31380 -21342 -31052
rect -21017 -31380 -20847 -31052
rect -20522 -31380 -20352 -31052
rect -20027 -31380 -19857 -31052
rect -19532 -31380 -19362 -31052
rect -19037 -31380 -18867 -31052
rect -18542 -31380 -18372 -31052
rect -18047 -31380 -17877 -31052
rect -17552 -31380 -17382 -31052
rect -17057 -31380 -16887 -31052
rect -16562 -31380 -16392 -31052
rect -16067 -31380 -15897 -31052
rect -15572 -31380 -15402 -31052
rect -15077 -31380 -14907 -31052
rect -14582 -31380 -14412 -31052
rect -14087 -31380 -13917 -31052
rect -13592 -31380 -13422 -31052
rect -13097 -31380 -12927 -31052
rect -12602 -31380 -12432 -31052
rect -12107 -31380 -11937 -31052
rect -11612 -31380 -11442 -31052
rect -11117 -31380 -10947 -31052
rect -10622 -31380 -10452 -31052
rect -10127 -31380 -9957 -31052
rect -9632 -31380 -9462 -31052
rect -9137 -31380 -8967 -31052
rect -8642 -31380 -8472 -31052
rect -8147 -31380 -7977 -31052
rect -7652 -31380 -7482 -31052
rect -7157 -31380 -6987 -31052
rect -6662 -31380 -6492 -31052
rect -6167 -31380 -5997 -31052
rect -5672 -31380 -5502 -31052
rect -5177 -31380 -5007 -31052
rect -4682 -31380 -4512 -31052
rect -4187 -31380 -4017 -31052
rect -3692 -31380 -3522 -31052
rect -3197 -31380 -3027 -31052
rect -2702 -31380 -2532 -31052
rect -2207 -31380 -2037 -31052
rect -1712 -31380 -1542 -31052
rect -1217 -31380 -1047 -31052
rect -722 -31380 -552 -31052
rect -227 -31380 -57 -31052
rect 268 -31380 438 -31052
rect 763 -31380 933 -31052
rect 1258 -31380 1428 -31052
rect 1753 -31380 1923 -31052
rect 2248 -31380 2418 -31052
rect 2743 -31380 2913 -31052
rect 3238 -31380 3408 -31052
rect 3733 -31380 3903 -31052
rect 4228 -31380 4398 -31052
rect 4723 -31380 4893 -31052
rect 5218 -31380 5388 -31052
rect 5713 -31380 5883 -31052
rect 6208 -31380 6378 -31052
rect 6703 -31380 6873 -31052
rect 7198 -31380 7368 -31052
rect 7693 -31380 7863 -31052
rect 8188 -31380 8358 -31052
rect 8683 -31380 8853 -31052
rect 9178 -31380 9348 -31052
rect 9673 -31380 9843 -31052
rect 10168 -31380 10338 -31052
rect 10663 -31380 10833 -31052
rect 11158 -31380 11328 -31052
rect 11653 -31380 11823 -31052
rect 12148 -31380 12318 -31052
rect 12643 -31380 12813 -31052
rect 13138 -31380 13308 -31052
rect 13633 -31380 13803 -31052
rect 14128 -31380 14298 -31052
rect 14623 -31380 14793 -31052
rect 15118 -31380 15288 -31052
rect 15613 -31380 15783 -31052
rect 16108 -31380 16278 -31052
rect 16603 -31380 16773 -31052
rect 17098 -31380 17268 -31052
rect 17593 -31380 17763 -31052
rect 18088 -31380 18258 -31052
rect 18583 -31380 18753 -31052
rect 19078 -31380 19248 -31052
rect 19573 -31380 19743 -31052
rect 20068 -31380 20238 -31052
rect 20563 -31380 20733 -31052
rect 21058 -31380 21228 -31052
rect 21553 -31380 21723 -31052
rect 22048 -31380 22218 -31052
rect 22543 -31380 22713 -31052
rect 23038 -31380 23208 -31052
rect 23533 -31380 23703 -31052
rect 24028 -31380 24198 -31052
rect 24523 -31380 24693 -31052
rect 25018 -31380 25188 -31052
rect 25513 -31380 25683 -31052
rect 26008 -31380 26178 -31052
rect 26503 -31380 26673 -31052
rect 26998 -31380 27168 -31052
rect 27493 -31380 27663 -31052
rect 27988 -31380 28158 -31052
rect 28483 -31380 28653 -31052
rect 28978 -31380 29148 -31052
rect 29473 -31380 29643 -31052
rect 29968 -31380 30138 -31052
rect 30463 -31380 30633 -31052
rect 30958 -31380 31128 -31052
rect 31453 -31380 31623 -31052
rect 31948 -31380 32118 -31052
rect 32443 -31380 32613 -31052
rect 32938 -31380 33108 -31052
rect 33433 -31380 33603 -31052
rect 33928 -31380 34098 -31052
rect 34423 -31380 34593 -31052
rect 34918 -31380 35088 -31052
rect 35413 -31380 35583 -31052
rect 35908 -31380 36078 -31052
rect 36403 -31380 36573 -31052
rect 36898 -31380 37068 -31052
rect 37393 -31380 37563 -31052
rect 37888 -31380 38058 -31052
rect 38383 -31380 38553 -31052
rect 38878 -31380 39048 -31052
rect 39373 -31380 39543 -31052
rect 39868 -31380 40038 -31052
rect 40363 -31380 40533 -31052
rect 40858 -31380 41028 -31052
rect 41353 -31380 41523 -31052
rect 41848 -31380 42018 -31052
rect 42343 -31380 42513 -31052
rect 42838 -31380 43008 -31052
rect 43333 -31380 43503 -31052
rect 43828 -31380 43998 -31052
rect 44323 -31380 44493 -31052
rect 44818 -31380 44988 -31052
rect 45313 -31380 45483 -31052
rect 45808 -31380 45978 -31052
rect 46303 -31380 46473 -31052
rect 46798 -31380 46968 -31052
rect 47293 -31380 47463 -31052
rect 47788 -31380 47958 -31052
rect 48283 -31380 48453 -31052
rect 48778 -31380 48948 -31052
rect 49273 -31380 49443 -31052
rect 49768 -31380 49938 -31052
rect 50263 -31380 50433 -31052
rect 50758 -31380 50928 -31052
rect 51253 -31380 51423 -31052
rect 51748 -31380 51918 -31052
rect 52243 -31380 52413 -31052
rect 52738 -31380 52908 -31052
rect 53233 -31380 53403 -31052
rect 53728 -31380 53898 -31052
rect 54223 -31380 54839 -31052
rect -55858 -31528 54839 -31380
rect -55858 -31856 -55497 -31528
rect -55172 -31856 -55002 -31528
rect -54677 -31856 -54507 -31528
rect -54182 -31856 -54012 -31528
rect -53687 -31856 -53517 -31528
rect -53192 -31856 -53022 -31528
rect -52697 -31856 -52527 -31528
rect -52202 -31856 -52032 -31528
rect -51707 -31856 -51537 -31528
rect -51212 -31856 -51042 -31528
rect -50717 -31856 -50547 -31528
rect -50222 -31856 -50052 -31528
rect -49727 -31856 -49557 -31528
rect -49232 -31856 -49062 -31528
rect -48737 -31856 -48567 -31528
rect -48242 -31856 -48072 -31528
rect -47747 -31856 -47577 -31528
rect -47252 -31856 -47082 -31528
rect -46757 -31856 -46587 -31528
rect -46262 -31856 -46092 -31528
rect -45767 -31856 -45597 -31528
rect -45272 -31856 -45102 -31528
rect -44777 -31856 -44607 -31528
rect -44282 -31856 -44112 -31528
rect -43787 -31856 -43617 -31528
rect -43292 -31856 -43122 -31528
rect -42797 -31856 -42627 -31528
rect -42302 -31856 -42132 -31528
rect -41807 -31856 -41637 -31528
rect -41312 -31856 -41142 -31528
rect -40817 -31856 -40647 -31528
rect -40322 -31856 -40152 -31528
rect -39827 -31856 -39657 -31528
rect -39332 -31856 -39162 -31528
rect -38837 -31856 -38667 -31528
rect -38342 -31856 -38172 -31528
rect -37847 -31856 -37677 -31528
rect -37352 -31856 -37182 -31528
rect -36857 -31856 -36687 -31528
rect -36362 -31856 -36192 -31528
rect -35867 -31856 -35697 -31528
rect -35372 -31856 -35202 -31528
rect -34877 -31856 -34707 -31528
rect -34382 -31856 -34212 -31528
rect -33887 -31856 -33717 -31528
rect -33392 -31856 -33222 -31528
rect -32897 -31856 -32727 -31528
rect -32402 -31856 -32232 -31528
rect -31907 -31856 -31737 -31528
rect -31412 -31856 -31242 -31528
rect -30917 -31856 -30747 -31528
rect -30422 -31856 -30252 -31528
rect -29927 -31856 -29757 -31528
rect -29432 -31856 -29262 -31528
rect -28937 -31856 -28767 -31528
rect -28442 -31856 -28272 -31528
rect -27947 -31856 -27777 -31528
rect -27452 -31856 -27282 -31528
rect -26957 -31856 -26787 -31528
rect -26462 -31856 -26292 -31528
rect -25967 -31856 -25797 -31528
rect -25472 -31856 -25302 -31528
rect -24977 -31856 -24807 -31528
rect -24482 -31856 -24312 -31528
rect -23987 -31856 -23817 -31528
rect -23492 -31856 -23322 -31528
rect -22997 -31856 -22827 -31528
rect -22502 -31856 -22332 -31528
rect -22007 -31856 -21837 -31528
rect -21512 -31856 -21342 -31528
rect -21017 -31856 -20847 -31528
rect -20522 -31856 -20352 -31528
rect -20027 -31856 -19857 -31528
rect -19532 -31856 -19362 -31528
rect -19037 -31856 -18867 -31528
rect -18542 -31856 -18372 -31528
rect -18047 -31856 -17877 -31528
rect -17552 -31856 -17382 -31528
rect -17057 -31856 -16887 -31528
rect -16562 -31856 -16392 -31528
rect -16067 -31856 -15897 -31528
rect -15572 -31856 -15402 -31528
rect -15077 -31856 -14907 -31528
rect -14582 -31856 -14412 -31528
rect -14087 -31856 -13917 -31528
rect -13592 -31856 -13422 -31528
rect -13097 -31856 -12927 -31528
rect -12602 -31856 -12432 -31528
rect -12107 -31856 -11937 -31528
rect -11612 -31856 -11442 -31528
rect -11117 -31856 -10947 -31528
rect -10622 -31856 -10452 -31528
rect -10127 -31856 -9957 -31528
rect -9632 -31856 -9462 -31528
rect -9137 -31856 -8967 -31528
rect -8642 -31856 -8472 -31528
rect -8147 -31856 -7977 -31528
rect -7652 -31856 -7482 -31528
rect -7157 -31856 -6987 -31528
rect -6662 -31856 -6492 -31528
rect -6167 -31856 -5997 -31528
rect -5672 -31856 -5502 -31528
rect -5177 -31856 -5007 -31528
rect -4682 -31856 -4512 -31528
rect -4187 -31856 -4017 -31528
rect -3692 -31856 -3522 -31528
rect -3197 -31856 -3027 -31528
rect -2702 -31856 -2532 -31528
rect -2207 -31856 -2037 -31528
rect -1712 -31856 -1542 -31528
rect -1217 -31856 -1047 -31528
rect -722 -31856 -552 -31528
rect -227 -31856 -57 -31528
rect 268 -31856 438 -31528
rect 763 -31856 933 -31528
rect 1258 -31856 1428 -31528
rect 1753 -31856 1923 -31528
rect 2248 -31856 2418 -31528
rect 2743 -31856 2913 -31528
rect 3238 -31856 3408 -31528
rect 3733 -31856 3903 -31528
rect 4228 -31856 4398 -31528
rect 4723 -31856 4893 -31528
rect 5218 -31856 5388 -31528
rect 5713 -31856 5883 -31528
rect 6208 -31856 6378 -31528
rect 6703 -31856 6873 -31528
rect 7198 -31856 7368 -31528
rect 7693 -31856 7863 -31528
rect 8188 -31856 8358 -31528
rect 8683 -31856 8853 -31528
rect 9178 -31856 9348 -31528
rect 9673 -31856 9843 -31528
rect 10168 -31856 10338 -31528
rect 10663 -31856 10833 -31528
rect 11158 -31856 11328 -31528
rect 11653 -31856 11823 -31528
rect 12148 -31856 12318 -31528
rect 12643 -31856 12813 -31528
rect 13138 -31856 13308 -31528
rect 13633 -31856 13803 -31528
rect 14128 -31856 14298 -31528
rect 14623 -31856 14793 -31528
rect 15118 -31856 15288 -31528
rect 15613 -31856 15783 -31528
rect 16108 -31856 16278 -31528
rect 16603 -31856 16773 -31528
rect 17098 -31856 17268 -31528
rect 17593 -31856 17763 -31528
rect 18088 -31856 18258 -31528
rect 18583 -31856 18753 -31528
rect 19078 -31856 19248 -31528
rect 19573 -31856 19743 -31528
rect 20068 -31856 20238 -31528
rect 20563 -31856 20733 -31528
rect 21058 -31856 21228 -31528
rect 21553 -31856 21723 -31528
rect 22048 -31856 22218 -31528
rect 22543 -31856 22713 -31528
rect 23038 -31856 23208 -31528
rect 23533 -31856 23703 -31528
rect 24028 -31856 24198 -31528
rect 24523 -31856 24693 -31528
rect 25018 -31856 25188 -31528
rect 25513 -31856 25683 -31528
rect 26008 -31856 26178 -31528
rect 26503 -31856 26673 -31528
rect 26998 -31856 27168 -31528
rect 27493 -31856 27663 -31528
rect 27988 -31856 28158 -31528
rect 28483 -31856 28653 -31528
rect 28978 -31856 29148 -31528
rect 29473 -31856 29643 -31528
rect 29968 -31856 30138 -31528
rect 30463 -31856 30633 -31528
rect 30958 -31856 31128 -31528
rect 31453 -31856 31623 -31528
rect 31948 -31856 32118 -31528
rect 32443 -31856 32613 -31528
rect 32938 -31856 33108 -31528
rect 33433 -31856 33603 -31528
rect 33928 -31856 34098 -31528
rect 34423 -31856 34593 -31528
rect 34918 -31856 35088 -31528
rect 35413 -31856 35583 -31528
rect 35908 -31856 36078 -31528
rect 36403 -31856 36573 -31528
rect 36898 -31856 37068 -31528
rect 37393 -31856 37563 -31528
rect 37888 -31856 38058 -31528
rect 38383 -31856 38553 -31528
rect 38878 -31856 39048 -31528
rect 39373 -31856 39543 -31528
rect 39868 -31856 40038 -31528
rect 40363 -31856 40533 -31528
rect 40858 -31856 41028 -31528
rect 41353 -31856 41523 -31528
rect 41848 -31856 42018 -31528
rect 42343 -31856 42513 -31528
rect 42838 -31856 43008 -31528
rect 43333 -31856 43503 -31528
rect 43828 -31856 43998 -31528
rect 44323 -31856 44493 -31528
rect 44818 -31856 44988 -31528
rect 45313 -31856 45483 -31528
rect 45808 -31856 45978 -31528
rect 46303 -31856 46473 -31528
rect 46798 -31856 46968 -31528
rect 47293 -31856 47463 -31528
rect 47788 -31856 47958 -31528
rect 48283 -31856 48453 -31528
rect 48778 -31856 48948 -31528
rect 49273 -31856 49443 -31528
rect 49768 -31856 49938 -31528
rect 50263 -31856 50433 -31528
rect 50758 -31856 50928 -31528
rect 51253 -31856 51423 -31528
rect 51748 -31856 51918 -31528
rect 52243 -31856 52413 -31528
rect 52738 -31856 52908 -31528
rect 53233 -31856 53403 -31528
rect 53728 -31856 53898 -31528
rect 54223 -31856 54839 -31528
rect -55858 -32147 54839 -31856
<< nsubdiff >>
rect -54929 26103 -54529 26166
rect -54929 25814 -54870 26103
rect -54596 25814 -54529 26103
rect -54929 25766 -54529 25814
rect -54352 26103 -53952 26166
rect -54352 25814 -54293 26103
rect -54019 25814 -53952 26103
rect -54352 25766 -53952 25814
rect -53775 26103 -53375 26166
rect -53775 25814 -53716 26103
rect -53442 25814 -53375 26103
rect -53775 25766 -53375 25814
rect -53198 26103 -52798 26166
rect -53198 25814 -53139 26103
rect -52865 25814 -52798 26103
rect -53198 25766 -52798 25814
rect -52621 26103 -52221 26166
rect -52621 25814 -52562 26103
rect -52288 25814 -52221 26103
rect -52621 25766 -52221 25814
rect -52044 26103 -51644 26166
rect -52044 25814 -51985 26103
rect -51711 25814 -51644 26103
rect -52044 25766 -51644 25814
rect -51467 26103 -51067 26166
rect -51467 25814 -51408 26103
rect -51134 25814 -51067 26103
rect -51467 25766 -51067 25814
rect -50890 26103 -50490 26166
rect -50890 25814 -50831 26103
rect -50557 25814 -50490 26103
rect -50890 25766 -50490 25814
rect -50313 26103 -49913 26166
rect -50313 25814 -50254 26103
rect -49980 25814 -49913 26103
rect -50313 25766 -49913 25814
rect -49736 26103 -49336 26166
rect -49736 25814 -49677 26103
rect -49403 25814 -49336 26103
rect -49736 25766 -49336 25814
rect -49159 26103 -48759 26166
rect -49159 25814 -49100 26103
rect -48826 25814 -48759 26103
rect -49159 25766 -48759 25814
rect -48582 26103 -48182 26166
rect -48582 25814 -48523 26103
rect -48249 25814 -48182 26103
rect -48582 25766 -48182 25814
rect -48005 26103 -47605 26166
rect -48005 25814 -47946 26103
rect -47672 25814 -47605 26103
rect -48005 25766 -47605 25814
rect -47428 26103 -47028 26166
rect -47428 25814 -47369 26103
rect -47095 25814 -47028 26103
rect -47428 25766 -47028 25814
rect -46851 26103 -46451 26166
rect -46851 25814 -46792 26103
rect -46518 25814 -46451 26103
rect -46851 25766 -46451 25814
rect -46274 26103 -45874 26166
rect -46274 25814 -46215 26103
rect -45941 25814 -45874 26103
rect -46274 25766 -45874 25814
rect -45697 26103 -45297 26166
rect -45697 25814 -45638 26103
rect -45364 25814 -45297 26103
rect -45697 25766 -45297 25814
rect -45120 26103 -44720 26166
rect -45120 25814 -45061 26103
rect -44787 25814 -44720 26103
rect -45120 25766 -44720 25814
rect -44543 26103 -44143 26166
rect -44543 25814 -44484 26103
rect -44210 25814 -44143 26103
rect -44543 25766 -44143 25814
rect -43966 26103 -43566 26166
rect -43966 25814 -43907 26103
rect -43633 25814 -43566 26103
rect -43966 25766 -43566 25814
rect -43389 26103 -42989 26166
rect -43389 25814 -43330 26103
rect -43056 25814 -42989 26103
rect -43389 25766 -42989 25814
rect -42812 26103 -42412 26166
rect -42812 25814 -42753 26103
rect -42479 25814 -42412 26103
rect -42812 25766 -42412 25814
rect -42235 26103 -41835 26166
rect -42235 25814 -42176 26103
rect -41902 25814 -41835 26103
rect -42235 25766 -41835 25814
rect -41658 26103 -41258 26166
rect -41658 25814 -41599 26103
rect -41325 25814 -41258 26103
rect -41658 25766 -41258 25814
rect -41081 26103 -40681 26166
rect -41081 25814 -41022 26103
rect -40748 25814 -40681 26103
rect -41081 25766 -40681 25814
rect -40504 26103 -40104 26166
rect -40504 25814 -40445 26103
rect -40171 25814 -40104 26103
rect -40504 25766 -40104 25814
rect -39927 26103 -39527 26166
rect -39927 25814 -39868 26103
rect -39594 25814 -39527 26103
rect -39927 25766 -39527 25814
rect -39350 26103 -38950 26166
rect -39350 25814 -39291 26103
rect -39017 25814 -38950 26103
rect -39350 25766 -38950 25814
rect -38773 26103 -38373 26166
rect -38773 25814 -38714 26103
rect -38440 25814 -38373 26103
rect -38773 25766 -38373 25814
rect -38196 26103 -37796 26166
rect -38196 25814 -38137 26103
rect -37863 25814 -37796 26103
rect -38196 25766 -37796 25814
rect -37619 26103 -37219 26166
rect -37619 25814 -37560 26103
rect -37286 25814 -37219 26103
rect -37619 25766 -37219 25814
rect -37042 26103 -36642 26166
rect -37042 25814 -36983 26103
rect -36709 25814 -36642 26103
rect -37042 25766 -36642 25814
rect -36465 26103 -36065 26166
rect -36465 25814 -36406 26103
rect -36132 25814 -36065 26103
rect -36465 25766 -36065 25814
rect -35888 26103 -35488 26166
rect -35888 25814 -35829 26103
rect -35555 25814 -35488 26103
rect -35888 25766 -35488 25814
rect -35311 26103 -34911 26166
rect -35311 25814 -35252 26103
rect -34978 25814 -34911 26103
rect -35311 25766 -34911 25814
rect -34734 26103 -34334 26166
rect -34734 25814 -34675 26103
rect -34401 25814 -34334 26103
rect -34734 25766 -34334 25814
rect -34157 26103 -33757 26166
rect -34157 25814 -34098 26103
rect -33824 25814 -33757 26103
rect -34157 25766 -33757 25814
rect -33580 26103 -33180 26166
rect -33580 25814 -33521 26103
rect -33247 25814 -33180 26103
rect -33580 25766 -33180 25814
rect -33003 26103 -32603 26166
rect -33003 25814 -32944 26103
rect -32670 25814 -32603 26103
rect -33003 25766 -32603 25814
rect -32426 26103 -32026 26166
rect -32426 25814 -32367 26103
rect -32093 25814 -32026 26103
rect -32426 25766 -32026 25814
rect -31849 26103 -31449 26166
rect -31849 25814 -31790 26103
rect -31516 25814 -31449 26103
rect -31849 25766 -31449 25814
rect -31272 26103 -30872 26166
rect -31272 25814 -31213 26103
rect -30939 25814 -30872 26103
rect -31272 25766 -30872 25814
rect -30695 26103 -30295 26166
rect -30695 25814 -30636 26103
rect -30362 25814 -30295 26103
rect -30695 25766 -30295 25814
rect -30118 26103 -29718 26166
rect -30118 25814 -30059 26103
rect -29785 25814 -29718 26103
rect -30118 25766 -29718 25814
rect -29541 26103 -29141 26166
rect -29541 25814 -29482 26103
rect -29208 25814 -29141 26103
rect -29541 25766 -29141 25814
rect -28964 26103 -28564 26166
rect -28964 25814 -28905 26103
rect -28631 25814 -28564 26103
rect -28964 25766 -28564 25814
rect -28387 26103 -27987 26166
rect -28387 25814 -28328 26103
rect -28054 25814 -27987 26103
rect -28387 25766 -27987 25814
rect -27810 26103 -27410 26166
rect -27810 25814 -27751 26103
rect -27477 25814 -27410 26103
rect -27810 25766 -27410 25814
rect -27233 26103 -26833 26166
rect -27233 25814 -27174 26103
rect -26900 25814 -26833 26103
rect -27233 25766 -26833 25814
rect -26656 26103 -26256 26166
rect -26656 25814 -26597 26103
rect -26323 25814 -26256 26103
rect -26656 25766 -26256 25814
rect -26079 26103 -25679 26166
rect -26079 25814 -26020 26103
rect -25746 25814 -25679 26103
rect -26079 25766 -25679 25814
rect -25502 26103 -25102 26166
rect -25502 25814 -25443 26103
rect -25169 25814 -25102 26103
rect -25502 25766 -25102 25814
rect -24925 26103 -24525 26166
rect -24925 25814 -24866 26103
rect -24592 25814 -24525 26103
rect -24925 25766 -24525 25814
rect -24348 26103 -23948 26166
rect -24348 25814 -24289 26103
rect -24015 25814 -23948 26103
rect -24348 25766 -23948 25814
rect -23771 26103 -23371 26166
rect -23771 25814 -23712 26103
rect -23438 25814 -23371 26103
rect -23771 25766 -23371 25814
rect -23194 26103 -22794 26166
rect -23194 25814 -23135 26103
rect -22861 25814 -22794 26103
rect -23194 25766 -22794 25814
rect -22617 26103 -22217 26166
rect -22617 25814 -22558 26103
rect -22284 25814 -22217 26103
rect -22617 25766 -22217 25814
rect -22040 26103 -21640 26166
rect -22040 25814 -21981 26103
rect -21707 25814 -21640 26103
rect -22040 25766 -21640 25814
rect -21463 26103 -21063 26166
rect -21463 25814 -21404 26103
rect -21130 25814 -21063 26103
rect -21463 25766 -21063 25814
rect -20886 26103 -20486 26166
rect -20886 25814 -20827 26103
rect -20553 25814 -20486 26103
rect -20886 25766 -20486 25814
rect -20309 26103 -19909 26166
rect -20309 25814 -20250 26103
rect -19976 25814 -19909 26103
rect -20309 25766 -19909 25814
rect -19732 26103 -19332 26166
rect -19732 25814 -19673 26103
rect -19399 25814 -19332 26103
rect -19732 25766 -19332 25814
rect -19155 26103 -18755 26166
rect -19155 25814 -19096 26103
rect -18822 25814 -18755 26103
rect -19155 25766 -18755 25814
rect -18578 26103 -18178 26166
rect -18578 25814 -18519 26103
rect -18245 25814 -18178 26103
rect -18578 25766 -18178 25814
rect -18001 26103 -17601 26166
rect -18001 25814 -17942 26103
rect -17668 25814 -17601 26103
rect -18001 25766 -17601 25814
rect -17424 26103 -17024 26166
rect -17424 25814 -17365 26103
rect -17091 25814 -17024 26103
rect -17424 25766 -17024 25814
rect -16847 26103 -16447 26166
rect -16847 25814 -16788 26103
rect -16514 25814 -16447 26103
rect -16847 25766 -16447 25814
rect -16270 26103 -15870 26166
rect -16270 25814 -16211 26103
rect -15937 25814 -15870 26103
rect -16270 25766 -15870 25814
rect -15693 26103 -15293 26166
rect -15693 25814 -15634 26103
rect -15360 25814 -15293 26103
rect -15693 25766 -15293 25814
rect -15116 26103 -14716 26166
rect -15116 25814 -15057 26103
rect -14783 25814 -14716 26103
rect -15116 25766 -14716 25814
rect -14539 26103 -14139 26166
rect -14539 25814 -14480 26103
rect -14206 25814 -14139 26103
rect -14539 25766 -14139 25814
rect -13962 26103 -13562 26166
rect -13962 25814 -13903 26103
rect -13629 25814 -13562 26103
rect -13962 25766 -13562 25814
rect -13385 26103 -12985 26166
rect -13385 25814 -13326 26103
rect -13052 25814 -12985 26103
rect -13385 25766 -12985 25814
rect -12808 26103 -12408 26166
rect -12808 25814 -12749 26103
rect -12475 25814 -12408 26103
rect -12808 25766 -12408 25814
rect -12231 26103 -11831 26166
rect -12231 25814 -12172 26103
rect -11898 25814 -11831 26103
rect -12231 25766 -11831 25814
rect -11654 26103 -11254 26166
rect -11654 25814 -11595 26103
rect -11321 25814 -11254 26103
rect -11654 25766 -11254 25814
rect -11077 26103 -10677 26166
rect -11077 25814 -11018 26103
rect -10744 25814 -10677 26103
rect -11077 25766 -10677 25814
rect -10500 26103 -10100 26166
rect -10500 25814 -10441 26103
rect -10167 25814 -10100 26103
rect -10500 25766 -10100 25814
rect -9923 26103 -9523 26166
rect -9923 25814 -9864 26103
rect -9590 25814 -9523 26103
rect -9923 25766 -9523 25814
rect -9346 26103 -8946 26166
rect -9346 25814 -9287 26103
rect -9013 25814 -8946 26103
rect -9346 25766 -8946 25814
rect -8769 26103 -8369 26166
rect -8769 25814 -8710 26103
rect -8436 25814 -8369 26103
rect -8769 25766 -8369 25814
rect -8192 26103 -7792 26166
rect -8192 25814 -8133 26103
rect -7859 25814 -7792 26103
rect -8192 25766 -7792 25814
rect -7615 26103 -7215 26166
rect -7615 25814 -7556 26103
rect -7282 25814 -7215 26103
rect -7615 25766 -7215 25814
rect -7038 26103 -6638 26166
rect -7038 25814 -6979 26103
rect -6705 25814 -6638 26103
rect -7038 25766 -6638 25814
rect -6461 26103 -6061 26166
rect -6461 25814 -6402 26103
rect -6128 25814 -6061 26103
rect -6461 25766 -6061 25814
rect -5884 26103 -5484 26166
rect -5884 25814 -5825 26103
rect -5551 25814 -5484 26103
rect -5884 25766 -5484 25814
rect -5307 26103 -4907 26166
rect -5307 25814 -5248 26103
rect -4974 25814 -4907 26103
rect -5307 25766 -4907 25814
rect -4730 26103 -4330 26166
rect -4730 25814 -4671 26103
rect -4397 25814 -4330 26103
rect -4730 25766 -4330 25814
rect -4153 26103 -3753 26166
rect -4153 25814 -4094 26103
rect -3820 25814 -3753 26103
rect -4153 25766 -3753 25814
rect -3576 26103 -3176 26166
rect -3576 25814 -3517 26103
rect -3243 25814 -3176 26103
rect -3576 25766 -3176 25814
rect -2999 26103 -2599 26166
rect -2999 25814 -2940 26103
rect -2666 25814 -2599 26103
rect -2999 25766 -2599 25814
rect -2422 26103 -2022 26166
rect -2422 25814 -2363 26103
rect -2089 25814 -2022 26103
rect -2422 25766 -2022 25814
rect -1845 26103 -1445 26166
rect -1845 25814 -1786 26103
rect -1512 25814 -1445 26103
rect -1845 25766 -1445 25814
rect -1268 26103 -868 26166
rect -1268 25814 -1209 26103
rect -935 25814 -868 26103
rect -1268 25766 -868 25814
rect -691 26103 -291 26166
rect -691 25814 -632 26103
rect -358 25814 -291 26103
rect -691 25766 -291 25814
rect -114 26103 286 26166
rect -114 25814 -55 26103
rect 219 25814 286 26103
rect -114 25766 286 25814
rect 463 26103 863 26166
rect 463 25814 522 26103
rect 796 25814 863 26103
rect 463 25766 863 25814
rect 1040 26103 1440 26166
rect 1040 25814 1099 26103
rect 1373 25814 1440 26103
rect 1040 25766 1440 25814
rect 1617 26103 2017 26166
rect 1617 25814 1676 26103
rect 1950 25814 2017 26103
rect 1617 25766 2017 25814
rect 2194 26103 2594 26166
rect 2194 25814 2253 26103
rect 2527 25814 2594 26103
rect 2194 25766 2594 25814
rect 2771 26103 3171 26166
rect 2771 25814 2830 26103
rect 3104 25814 3171 26103
rect 2771 25766 3171 25814
rect 3348 26103 3748 26166
rect 3348 25814 3407 26103
rect 3681 25814 3748 26103
rect 3348 25766 3748 25814
rect 3925 26103 4325 26166
rect 3925 25814 3984 26103
rect 4258 25814 4325 26103
rect 3925 25766 4325 25814
rect 4502 26103 4902 26166
rect 4502 25814 4561 26103
rect 4835 25814 4902 26103
rect 4502 25766 4902 25814
rect 5079 26103 5479 26166
rect 5079 25814 5138 26103
rect 5412 25814 5479 26103
rect 5079 25766 5479 25814
rect 5656 26103 6056 26166
rect 5656 25814 5715 26103
rect 5989 25814 6056 26103
rect 5656 25766 6056 25814
rect 6233 26103 6633 26166
rect 6233 25814 6292 26103
rect 6566 25814 6633 26103
rect 6233 25766 6633 25814
rect 6810 26103 7210 26166
rect 6810 25814 6869 26103
rect 7143 25814 7210 26103
rect 6810 25766 7210 25814
rect 7387 26103 7787 26166
rect 7387 25814 7446 26103
rect 7720 25814 7787 26103
rect 7387 25766 7787 25814
rect 7964 26103 8364 26166
rect 7964 25814 8023 26103
rect 8297 25814 8364 26103
rect 7964 25766 8364 25814
rect 8541 26103 8941 26166
rect 8541 25814 8600 26103
rect 8874 25814 8941 26103
rect 8541 25766 8941 25814
rect 9118 26103 9518 26166
rect 9118 25814 9177 26103
rect 9451 25814 9518 26103
rect 9118 25766 9518 25814
rect 9695 26103 10095 26166
rect 9695 25814 9754 26103
rect 10028 25814 10095 26103
rect 9695 25766 10095 25814
rect 10272 26103 10672 26166
rect 10272 25814 10331 26103
rect 10605 25814 10672 26103
rect 10272 25766 10672 25814
rect 10849 26103 11249 26166
rect 10849 25814 10908 26103
rect 11182 25814 11249 26103
rect 10849 25766 11249 25814
rect 11426 26103 11826 26166
rect 11426 25814 11485 26103
rect 11759 25814 11826 26103
rect 11426 25766 11826 25814
rect 12003 26103 12403 26166
rect 12003 25814 12062 26103
rect 12336 25814 12403 26103
rect 12003 25766 12403 25814
rect 12580 26103 12980 26166
rect 12580 25814 12639 26103
rect 12913 25814 12980 26103
rect 12580 25766 12980 25814
rect 13157 26103 13557 26166
rect 13157 25814 13216 26103
rect 13490 25814 13557 26103
rect 13157 25766 13557 25814
rect 13734 26103 14134 26166
rect 13734 25814 13793 26103
rect 14067 25814 14134 26103
rect 13734 25766 14134 25814
rect 14311 26103 14711 26166
rect 14311 25814 14370 26103
rect 14644 25814 14711 26103
rect 14311 25766 14711 25814
rect 14888 26103 15288 26166
rect 14888 25814 14947 26103
rect 15221 25814 15288 26103
rect 14888 25766 15288 25814
rect 15465 26103 15865 26166
rect 15465 25814 15524 26103
rect 15798 25814 15865 26103
rect 15465 25766 15865 25814
rect 16042 26103 16442 26166
rect 16042 25814 16101 26103
rect 16375 25814 16442 26103
rect 16042 25766 16442 25814
rect 16619 26103 17019 26166
rect 16619 25814 16678 26103
rect 16952 25814 17019 26103
rect 16619 25766 17019 25814
rect 17196 26103 17596 26166
rect 17196 25814 17255 26103
rect 17529 25814 17596 26103
rect 17196 25766 17596 25814
rect 17773 26103 18173 26166
rect 17773 25814 17832 26103
rect 18106 25814 18173 26103
rect 17773 25766 18173 25814
rect 18350 26103 18750 26166
rect 18350 25814 18409 26103
rect 18683 25814 18750 26103
rect 18350 25766 18750 25814
rect 18927 26103 19327 26166
rect 18927 25814 18986 26103
rect 19260 25814 19327 26103
rect 18927 25766 19327 25814
rect 19504 26103 19904 26166
rect 19504 25814 19563 26103
rect 19837 25814 19904 26103
rect 19504 25766 19904 25814
rect 20081 26103 20481 26166
rect 20081 25814 20140 26103
rect 20414 25814 20481 26103
rect 20081 25766 20481 25814
rect 20658 26103 21058 26166
rect 20658 25814 20717 26103
rect 20991 25814 21058 26103
rect 20658 25766 21058 25814
rect 21235 26103 21635 26166
rect 21235 25814 21294 26103
rect 21568 25814 21635 26103
rect 21235 25766 21635 25814
rect 21812 26103 22212 26166
rect 21812 25814 21871 26103
rect 22145 25814 22212 26103
rect 21812 25766 22212 25814
rect 22389 26103 22789 26166
rect 22389 25814 22448 26103
rect 22722 25814 22789 26103
rect 22389 25766 22789 25814
rect 22966 26103 23366 26166
rect 22966 25814 23025 26103
rect 23299 25814 23366 26103
rect 22966 25766 23366 25814
rect 23543 26103 23943 26166
rect 23543 25814 23602 26103
rect 23876 25814 23943 26103
rect 23543 25766 23943 25814
rect 24120 26103 24520 26166
rect 24120 25814 24179 26103
rect 24453 25814 24520 26103
rect 24120 25766 24520 25814
rect 24697 26103 25097 26166
rect 24697 25814 24756 26103
rect 25030 25814 25097 26103
rect 24697 25766 25097 25814
rect 25274 26103 25674 26166
rect 25274 25814 25333 26103
rect 25607 25814 25674 26103
rect 25274 25766 25674 25814
rect 25851 26103 26251 26166
rect 25851 25814 25910 26103
rect 26184 25814 26251 26103
rect 25851 25766 26251 25814
rect 26428 26103 26828 26166
rect 26428 25814 26487 26103
rect 26761 25814 26828 26103
rect 26428 25766 26828 25814
rect 27005 26103 27405 26166
rect 27005 25814 27064 26103
rect 27338 25814 27405 26103
rect 27005 25766 27405 25814
rect 27582 26103 27982 26166
rect 27582 25814 27641 26103
rect 27915 25814 27982 26103
rect 27582 25766 27982 25814
rect 28159 26103 28559 26166
rect 28159 25814 28218 26103
rect 28492 25814 28559 26103
rect 28159 25766 28559 25814
rect 28736 26103 29136 26166
rect 28736 25814 28795 26103
rect 29069 25814 29136 26103
rect 28736 25766 29136 25814
rect 29313 26103 29713 26166
rect 29313 25814 29372 26103
rect 29646 25814 29713 26103
rect 29313 25766 29713 25814
rect 29890 26103 30290 26166
rect 29890 25814 29949 26103
rect 30223 25814 30290 26103
rect 29890 25766 30290 25814
rect 30467 26103 30867 26166
rect 30467 25814 30526 26103
rect 30800 25814 30867 26103
rect 30467 25766 30867 25814
rect 31044 26103 31444 26166
rect 31044 25814 31103 26103
rect 31377 25814 31444 26103
rect 31044 25766 31444 25814
rect 31621 26103 32021 26166
rect 31621 25814 31680 26103
rect 31954 25814 32021 26103
rect 31621 25766 32021 25814
rect 32198 26103 32598 26166
rect 32198 25814 32257 26103
rect 32531 25814 32598 26103
rect 32198 25766 32598 25814
rect 32775 26103 33175 26166
rect 32775 25814 32834 26103
rect 33108 25814 33175 26103
rect 32775 25766 33175 25814
rect 33352 26103 33752 26166
rect 33352 25814 33411 26103
rect 33685 25814 33752 26103
rect 33352 25766 33752 25814
rect 33929 26103 34329 26166
rect 33929 25814 33988 26103
rect 34262 25814 34329 26103
rect 33929 25766 34329 25814
rect 34506 26103 34906 26166
rect 34506 25814 34565 26103
rect 34839 25814 34906 26103
rect 34506 25766 34906 25814
rect 35083 26103 35483 26166
rect 35083 25814 35142 26103
rect 35416 25814 35483 26103
rect 35083 25766 35483 25814
rect 35660 26103 36060 26166
rect 35660 25814 35719 26103
rect 35993 25814 36060 26103
rect 35660 25766 36060 25814
rect 36237 26103 36637 26166
rect 36237 25814 36296 26103
rect 36570 25814 36637 26103
rect 36237 25766 36637 25814
rect 36814 26103 37214 26166
rect 36814 25814 36873 26103
rect 37147 25814 37214 26103
rect 36814 25766 37214 25814
rect 37391 26103 37791 26166
rect 37391 25814 37450 26103
rect 37724 25814 37791 26103
rect 37391 25766 37791 25814
rect 37968 26103 38368 26166
rect 37968 25814 38027 26103
rect 38301 25814 38368 26103
rect 37968 25766 38368 25814
rect 38545 26103 38945 26166
rect 38545 25814 38604 26103
rect 38878 25814 38945 26103
rect 38545 25766 38945 25814
rect 39122 26103 39522 26166
rect 39122 25814 39181 26103
rect 39455 25814 39522 26103
rect 39122 25766 39522 25814
rect 39699 26103 40099 26166
rect 39699 25814 39758 26103
rect 40032 25814 40099 26103
rect 39699 25766 40099 25814
rect 40276 26103 40676 26166
rect 40276 25814 40335 26103
rect 40609 25814 40676 26103
rect 40276 25766 40676 25814
rect 40853 26103 41253 26166
rect 40853 25814 40912 26103
rect 41186 25814 41253 26103
rect 40853 25766 41253 25814
rect 41430 26103 41830 26166
rect 41430 25814 41489 26103
rect 41763 25814 41830 26103
rect 41430 25766 41830 25814
rect 42007 26103 42407 26166
rect 42007 25814 42066 26103
rect 42340 25814 42407 26103
rect 42007 25766 42407 25814
rect 42584 26103 42984 26166
rect 42584 25814 42643 26103
rect 42917 25814 42984 26103
rect 42584 25766 42984 25814
rect 43161 26103 43561 26166
rect 43161 25814 43220 26103
rect 43494 25814 43561 26103
rect 43161 25766 43561 25814
rect 43738 26103 44138 26166
rect 43738 25814 43797 26103
rect 44071 25814 44138 26103
rect 43738 25766 44138 25814
rect 44315 26103 44715 26166
rect 44315 25814 44374 26103
rect 44648 25814 44715 26103
rect 44315 25766 44715 25814
rect 44892 26103 45292 26166
rect 44892 25814 44951 26103
rect 45225 25814 45292 26103
rect 44892 25766 45292 25814
rect 45469 26103 45869 26166
rect 45469 25814 45528 26103
rect 45802 25814 45869 26103
rect 45469 25766 45869 25814
rect 46046 26103 46446 26166
rect 46046 25814 46105 26103
rect 46379 25814 46446 26103
rect 46046 25766 46446 25814
rect 46623 26103 47023 26166
rect 46623 25814 46682 26103
rect 46956 25814 47023 26103
rect 46623 25766 47023 25814
rect 47200 26103 47600 26166
rect 47200 25814 47259 26103
rect 47533 25814 47600 26103
rect 47200 25766 47600 25814
rect 47777 26103 48177 26166
rect 47777 25814 47836 26103
rect 48110 25814 48177 26103
rect 47777 25766 48177 25814
rect 48354 26103 48754 26166
rect 48354 25814 48413 26103
rect 48687 25814 48754 26103
rect 48354 25766 48754 25814
rect 48931 26103 49331 26166
rect 48931 25814 48990 26103
rect 49264 25814 49331 26103
rect 48931 25766 49331 25814
rect 49508 26103 49908 26166
rect 49508 25814 49567 26103
rect 49841 25814 49908 26103
rect 49508 25766 49908 25814
rect 50085 26103 50485 26166
rect 50085 25814 50144 26103
rect 50418 25814 50485 26103
rect 50085 25766 50485 25814
rect 50662 26103 51062 26166
rect 50662 25814 50721 26103
rect 50995 25814 51062 26103
rect 50662 25766 51062 25814
rect 51239 26103 51639 26166
rect 51239 25814 51298 26103
rect 51572 25814 51639 26103
rect 51239 25766 51639 25814
rect 51816 26103 52216 26166
rect 51816 25814 51875 26103
rect 52149 25814 52216 26103
rect 51816 25766 52216 25814
rect 52393 26103 52793 26166
rect 52393 25814 52452 26103
rect 52726 25814 52793 26103
rect 52393 25766 52793 25814
rect 52970 26103 53370 26166
rect 52970 25814 53029 26103
rect 53303 25814 53370 26103
rect 52970 25766 53370 25814
rect 53547 26103 53947 26166
rect 53547 25814 53606 26103
rect 53880 25814 53947 26103
rect 53547 25766 53947 25814
rect 54124 26103 54524 26166
rect 54124 25814 54183 26103
rect 54457 25814 54524 26103
rect 54124 25766 54524 25814
rect 54701 26103 55101 26166
rect 54701 25814 54760 26103
rect 55034 25814 55101 26103
rect 54701 25766 55101 25814
rect 55278 26103 55678 26166
rect 55278 25814 55337 26103
rect 55611 25814 55678 26103
rect 55278 25766 55678 25814
rect 55855 26103 56255 26166
rect 55855 25814 55914 26103
rect 56188 25814 56255 26103
rect 55855 25766 56255 25814
rect -54929 25545 -54529 25608
rect -54929 25256 -54870 25545
rect -54596 25256 -54529 25545
rect -54929 25208 -54529 25256
rect -54352 25545 -53952 25608
rect -54352 25256 -54293 25545
rect -54019 25256 -53952 25545
rect -54352 25208 -53952 25256
rect -53775 25545 -53375 25608
rect -53775 25256 -53716 25545
rect -53442 25256 -53375 25545
rect -53775 25208 -53375 25256
rect -53198 25545 -52798 25608
rect -53198 25256 -53139 25545
rect -52865 25256 -52798 25545
rect -53198 25208 -52798 25256
rect -52621 25545 -52221 25608
rect -52621 25256 -52562 25545
rect -52288 25256 -52221 25545
rect -52621 25208 -52221 25256
rect -52044 25545 -51644 25608
rect -52044 25256 -51985 25545
rect -51711 25256 -51644 25545
rect -52044 25208 -51644 25256
rect -51467 25545 -51067 25608
rect -51467 25256 -51408 25545
rect -51134 25256 -51067 25545
rect -51467 25208 -51067 25256
rect -50890 25545 -50490 25608
rect -50890 25256 -50831 25545
rect -50557 25256 -50490 25545
rect -50890 25208 -50490 25256
rect -50313 25545 -49913 25608
rect -50313 25256 -50254 25545
rect -49980 25256 -49913 25545
rect -50313 25208 -49913 25256
rect -49736 25545 -49336 25608
rect -49736 25256 -49677 25545
rect -49403 25256 -49336 25545
rect -49736 25208 -49336 25256
rect -49159 25545 -48759 25608
rect -49159 25256 -49100 25545
rect -48826 25256 -48759 25545
rect -49159 25208 -48759 25256
rect -48582 25545 -48182 25608
rect -48582 25256 -48523 25545
rect -48249 25256 -48182 25545
rect -48582 25208 -48182 25256
rect -48005 25545 -47605 25608
rect -48005 25256 -47946 25545
rect -47672 25256 -47605 25545
rect -48005 25208 -47605 25256
rect -47428 25545 -47028 25608
rect -47428 25256 -47369 25545
rect -47095 25256 -47028 25545
rect -47428 25208 -47028 25256
rect -46851 25545 -46451 25608
rect -46851 25256 -46792 25545
rect -46518 25256 -46451 25545
rect -46851 25208 -46451 25256
rect -46274 25545 -45874 25608
rect -46274 25256 -46215 25545
rect -45941 25256 -45874 25545
rect -46274 25208 -45874 25256
rect -45697 25545 -45297 25608
rect -45697 25256 -45638 25545
rect -45364 25256 -45297 25545
rect -45697 25208 -45297 25256
rect -45120 25545 -44720 25608
rect -45120 25256 -45061 25545
rect -44787 25256 -44720 25545
rect -45120 25208 -44720 25256
rect -44543 25545 -44143 25608
rect -44543 25256 -44484 25545
rect -44210 25256 -44143 25545
rect -44543 25208 -44143 25256
rect -43966 25545 -43566 25608
rect -43966 25256 -43907 25545
rect -43633 25256 -43566 25545
rect -43966 25208 -43566 25256
rect -43389 25545 -42989 25608
rect -43389 25256 -43330 25545
rect -43056 25256 -42989 25545
rect -43389 25208 -42989 25256
rect -42812 25545 -42412 25608
rect -42812 25256 -42753 25545
rect -42479 25256 -42412 25545
rect -42812 25208 -42412 25256
rect -42235 25545 -41835 25608
rect -42235 25256 -42176 25545
rect -41902 25256 -41835 25545
rect -42235 25208 -41835 25256
rect -41658 25545 -41258 25608
rect -41658 25256 -41599 25545
rect -41325 25256 -41258 25545
rect -41658 25208 -41258 25256
rect -41081 25545 -40681 25608
rect -41081 25256 -41022 25545
rect -40748 25256 -40681 25545
rect -41081 25208 -40681 25256
rect -40504 25545 -40104 25608
rect -40504 25256 -40445 25545
rect -40171 25256 -40104 25545
rect -40504 25208 -40104 25256
rect -39927 25545 -39527 25608
rect -39927 25256 -39868 25545
rect -39594 25256 -39527 25545
rect -39927 25208 -39527 25256
rect -39350 25545 -38950 25608
rect -39350 25256 -39291 25545
rect -39017 25256 -38950 25545
rect -39350 25208 -38950 25256
rect -38773 25545 -38373 25608
rect -38773 25256 -38714 25545
rect -38440 25256 -38373 25545
rect -38773 25208 -38373 25256
rect -38196 25545 -37796 25608
rect -38196 25256 -38137 25545
rect -37863 25256 -37796 25545
rect -38196 25208 -37796 25256
rect -37619 25545 -37219 25608
rect -37619 25256 -37560 25545
rect -37286 25256 -37219 25545
rect -37619 25208 -37219 25256
rect -37042 25545 -36642 25608
rect -37042 25256 -36983 25545
rect -36709 25256 -36642 25545
rect -37042 25208 -36642 25256
rect -36465 25545 -36065 25608
rect -36465 25256 -36406 25545
rect -36132 25256 -36065 25545
rect -36465 25208 -36065 25256
rect -35888 25545 -35488 25608
rect -35888 25256 -35829 25545
rect -35555 25256 -35488 25545
rect -35888 25208 -35488 25256
rect -35311 25545 -34911 25608
rect -35311 25256 -35252 25545
rect -34978 25256 -34911 25545
rect -35311 25208 -34911 25256
rect -34734 25545 -34334 25608
rect -34734 25256 -34675 25545
rect -34401 25256 -34334 25545
rect -34734 25208 -34334 25256
rect -34157 25545 -33757 25608
rect -34157 25256 -34098 25545
rect -33824 25256 -33757 25545
rect -34157 25208 -33757 25256
rect -33580 25545 -33180 25608
rect -33580 25256 -33521 25545
rect -33247 25256 -33180 25545
rect -33580 25208 -33180 25256
rect -33003 25545 -32603 25608
rect -33003 25256 -32944 25545
rect -32670 25256 -32603 25545
rect -33003 25208 -32603 25256
rect -32426 25545 -32026 25608
rect -32426 25256 -32367 25545
rect -32093 25256 -32026 25545
rect -32426 25208 -32026 25256
rect -31849 25545 -31449 25608
rect -31849 25256 -31790 25545
rect -31516 25256 -31449 25545
rect -31849 25208 -31449 25256
rect -31272 25545 -30872 25608
rect -31272 25256 -31213 25545
rect -30939 25256 -30872 25545
rect -31272 25208 -30872 25256
rect -30695 25545 -30295 25608
rect -30695 25256 -30636 25545
rect -30362 25256 -30295 25545
rect -30695 25208 -30295 25256
rect -30118 25545 -29718 25608
rect -30118 25256 -30059 25545
rect -29785 25256 -29718 25545
rect -30118 25208 -29718 25256
rect -29541 25545 -29141 25608
rect -29541 25256 -29482 25545
rect -29208 25256 -29141 25545
rect -29541 25208 -29141 25256
rect -28964 25545 -28564 25608
rect -28964 25256 -28905 25545
rect -28631 25256 -28564 25545
rect -28964 25208 -28564 25256
rect -28387 25545 -27987 25608
rect -28387 25256 -28328 25545
rect -28054 25256 -27987 25545
rect -28387 25208 -27987 25256
rect -27810 25545 -27410 25608
rect -27810 25256 -27751 25545
rect -27477 25256 -27410 25545
rect -27810 25208 -27410 25256
rect -27233 25545 -26833 25608
rect -27233 25256 -27174 25545
rect -26900 25256 -26833 25545
rect -27233 25208 -26833 25256
rect -26656 25545 -26256 25608
rect -26656 25256 -26597 25545
rect -26323 25256 -26256 25545
rect -26656 25208 -26256 25256
rect -26079 25545 -25679 25608
rect -26079 25256 -26020 25545
rect -25746 25256 -25679 25545
rect -26079 25208 -25679 25256
rect -25502 25545 -25102 25608
rect -25502 25256 -25443 25545
rect -25169 25256 -25102 25545
rect -25502 25208 -25102 25256
rect -24925 25545 -24525 25608
rect -24925 25256 -24866 25545
rect -24592 25256 -24525 25545
rect -24925 25208 -24525 25256
rect -24348 25545 -23948 25608
rect -24348 25256 -24289 25545
rect -24015 25256 -23948 25545
rect -24348 25208 -23948 25256
rect -23771 25545 -23371 25608
rect -23771 25256 -23712 25545
rect -23438 25256 -23371 25545
rect -23771 25208 -23371 25256
rect -23194 25545 -22794 25608
rect -23194 25256 -23135 25545
rect -22861 25256 -22794 25545
rect -23194 25208 -22794 25256
rect -22617 25545 -22217 25608
rect -22617 25256 -22558 25545
rect -22284 25256 -22217 25545
rect -22617 25208 -22217 25256
rect -22040 25545 -21640 25608
rect -22040 25256 -21981 25545
rect -21707 25256 -21640 25545
rect -22040 25208 -21640 25256
rect -21463 25545 -21063 25608
rect -21463 25256 -21404 25545
rect -21130 25256 -21063 25545
rect -21463 25208 -21063 25256
rect -20886 25545 -20486 25608
rect -20886 25256 -20827 25545
rect -20553 25256 -20486 25545
rect -20886 25208 -20486 25256
rect -20309 25545 -19909 25608
rect -20309 25256 -20250 25545
rect -19976 25256 -19909 25545
rect -20309 25208 -19909 25256
rect -19732 25545 -19332 25608
rect -19732 25256 -19673 25545
rect -19399 25256 -19332 25545
rect -19732 25208 -19332 25256
rect -19155 25545 -18755 25608
rect -19155 25256 -19096 25545
rect -18822 25256 -18755 25545
rect -19155 25208 -18755 25256
rect -18578 25545 -18178 25608
rect -18578 25256 -18519 25545
rect -18245 25256 -18178 25545
rect -18578 25208 -18178 25256
rect -18001 25545 -17601 25608
rect -18001 25256 -17942 25545
rect -17668 25256 -17601 25545
rect -18001 25208 -17601 25256
rect -17424 25545 -17024 25608
rect -17424 25256 -17365 25545
rect -17091 25256 -17024 25545
rect -17424 25208 -17024 25256
rect -16847 25545 -16447 25608
rect -16847 25256 -16788 25545
rect -16514 25256 -16447 25545
rect -16847 25208 -16447 25256
rect -16270 25545 -15870 25608
rect -16270 25256 -16211 25545
rect -15937 25256 -15870 25545
rect -16270 25208 -15870 25256
rect -15693 25545 -15293 25608
rect -15693 25256 -15634 25545
rect -15360 25256 -15293 25545
rect -15693 25208 -15293 25256
rect -15116 25545 -14716 25608
rect -15116 25256 -15057 25545
rect -14783 25256 -14716 25545
rect -15116 25208 -14716 25256
rect -14539 25545 -14139 25608
rect -14539 25256 -14480 25545
rect -14206 25256 -14139 25545
rect -14539 25208 -14139 25256
rect -13962 25545 -13562 25608
rect -13962 25256 -13903 25545
rect -13629 25256 -13562 25545
rect -13962 25208 -13562 25256
rect -13385 25545 -12985 25608
rect -13385 25256 -13326 25545
rect -13052 25256 -12985 25545
rect -13385 25208 -12985 25256
rect -12808 25545 -12408 25608
rect -12808 25256 -12749 25545
rect -12475 25256 -12408 25545
rect -12808 25208 -12408 25256
rect -12231 25545 -11831 25608
rect -12231 25256 -12172 25545
rect -11898 25256 -11831 25545
rect -12231 25208 -11831 25256
rect -11654 25545 -11254 25608
rect -11654 25256 -11595 25545
rect -11321 25256 -11254 25545
rect -11654 25208 -11254 25256
rect -11077 25545 -10677 25608
rect -11077 25256 -11018 25545
rect -10744 25256 -10677 25545
rect -11077 25208 -10677 25256
rect -10500 25545 -10100 25608
rect -10500 25256 -10441 25545
rect -10167 25256 -10100 25545
rect -10500 25208 -10100 25256
rect -9923 25545 -9523 25608
rect -9923 25256 -9864 25545
rect -9590 25256 -9523 25545
rect -9923 25208 -9523 25256
rect -9346 25545 -8946 25608
rect -9346 25256 -9287 25545
rect -9013 25256 -8946 25545
rect -9346 25208 -8946 25256
rect -8769 25545 -8369 25608
rect -8769 25256 -8710 25545
rect -8436 25256 -8369 25545
rect -8769 25208 -8369 25256
rect -8192 25545 -7792 25608
rect -8192 25256 -8133 25545
rect -7859 25256 -7792 25545
rect -8192 25208 -7792 25256
rect -7615 25545 -7215 25608
rect -7615 25256 -7556 25545
rect -7282 25256 -7215 25545
rect -7615 25208 -7215 25256
rect -7038 25545 -6638 25608
rect -7038 25256 -6979 25545
rect -6705 25256 -6638 25545
rect -7038 25208 -6638 25256
rect -6461 25545 -6061 25608
rect -6461 25256 -6402 25545
rect -6128 25256 -6061 25545
rect -6461 25208 -6061 25256
rect -5884 25545 -5484 25608
rect -5884 25256 -5825 25545
rect -5551 25256 -5484 25545
rect -5884 25208 -5484 25256
rect -5307 25545 -4907 25608
rect -5307 25256 -5248 25545
rect -4974 25256 -4907 25545
rect -5307 25208 -4907 25256
rect -4730 25545 -4330 25608
rect -4730 25256 -4671 25545
rect -4397 25256 -4330 25545
rect -4730 25208 -4330 25256
rect -4153 25545 -3753 25608
rect -4153 25256 -4094 25545
rect -3820 25256 -3753 25545
rect -4153 25208 -3753 25256
rect -3576 25545 -3176 25608
rect -3576 25256 -3517 25545
rect -3243 25256 -3176 25545
rect -3576 25208 -3176 25256
rect -2999 25545 -2599 25608
rect -2999 25256 -2940 25545
rect -2666 25256 -2599 25545
rect -2999 25208 -2599 25256
rect -2422 25545 -2022 25608
rect -2422 25256 -2363 25545
rect -2089 25256 -2022 25545
rect -2422 25208 -2022 25256
rect -1845 25545 -1445 25608
rect -1845 25256 -1786 25545
rect -1512 25256 -1445 25545
rect -1845 25208 -1445 25256
rect -1268 25545 -868 25608
rect -1268 25256 -1209 25545
rect -935 25256 -868 25545
rect -1268 25208 -868 25256
rect -691 25545 -291 25608
rect -691 25256 -632 25545
rect -358 25256 -291 25545
rect -691 25208 -291 25256
rect -114 25545 286 25608
rect -114 25256 -55 25545
rect 219 25256 286 25545
rect -114 25208 286 25256
rect 463 25545 863 25608
rect 463 25256 522 25545
rect 796 25256 863 25545
rect 463 25208 863 25256
rect 1040 25545 1440 25608
rect 1040 25256 1099 25545
rect 1373 25256 1440 25545
rect 1040 25208 1440 25256
rect 1617 25545 2017 25608
rect 1617 25256 1676 25545
rect 1950 25256 2017 25545
rect 1617 25208 2017 25256
rect 2194 25545 2594 25608
rect 2194 25256 2253 25545
rect 2527 25256 2594 25545
rect 2194 25208 2594 25256
rect 2771 25545 3171 25608
rect 2771 25256 2830 25545
rect 3104 25256 3171 25545
rect 2771 25208 3171 25256
rect 3348 25545 3748 25608
rect 3348 25256 3407 25545
rect 3681 25256 3748 25545
rect 3348 25208 3748 25256
rect 3925 25545 4325 25608
rect 3925 25256 3984 25545
rect 4258 25256 4325 25545
rect 3925 25208 4325 25256
rect 4502 25545 4902 25608
rect 4502 25256 4561 25545
rect 4835 25256 4902 25545
rect 4502 25208 4902 25256
rect 5079 25545 5479 25608
rect 5079 25256 5138 25545
rect 5412 25256 5479 25545
rect 5079 25208 5479 25256
rect 5656 25545 6056 25608
rect 5656 25256 5715 25545
rect 5989 25256 6056 25545
rect 5656 25208 6056 25256
rect 6233 25545 6633 25608
rect 6233 25256 6292 25545
rect 6566 25256 6633 25545
rect 6233 25208 6633 25256
rect 6810 25545 7210 25608
rect 6810 25256 6869 25545
rect 7143 25256 7210 25545
rect 6810 25208 7210 25256
rect 7387 25545 7787 25608
rect 7387 25256 7446 25545
rect 7720 25256 7787 25545
rect 7387 25208 7787 25256
rect 7964 25545 8364 25608
rect 7964 25256 8023 25545
rect 8297 25256 8364 25545
rect 7964 25208 8364 25256
rect 8541 25545 8941 25608
rect 8541 25256 8600 25545
rect 8874 25256 8941 25545
rect 8541 25208 8941 25256
rect 9118 25545 9518 25608
rect 9118 25256 9177 25545
rect 9451 25256 9518 25545
rect 9118 25208 9518 25256
rect 9695 25545 10095 25608
rect 9695 25256 9754 25545
rect 10028 25256 10095 25545
rect 9695 25208 10095 25256
rect 10272 25545 10672 25608
rect 10272 25256 10331 25545
rect 10605 25256 10672 25545
rect 10272 25208 10672 25256
rect 10849 25545 11249 25608
rect 10849 25256 10908 25545
rect 11182 25256 11249 25545
rect 10849 25208 11249 25256
rect 11426 25545 11826 25608
rect 11426 25256 11485 25545
rect 11759 25256 11826 25545
rect 11426 25208 11826 25256
rect 12003 25545 12403 25608
rect 12003 25256 12062 25545
rect 12336 25256 12403 25545
rect 12003 25208 12403 25256
rect 12580 25545 12980 25608
rect 12580 25256 12639 25545
rect 12913 25256 12980 25545
rect 12580 25208 12980 25256
rect 13157 25545 13557 25608
rect 13157 25256 13216 25545
rect 13490 25256 13557 25545
rect 13157 25208 13557 25256
rect 13734 25545 14134 25608
rect 13734 25256 13793 25545
rect 14067 25256 14134 25545
rect 13734 25208 14134 25256
rect 14311 25545 14711 25608
rect 14311 25256 14370 25545
rect 14644 25256 14711 25545
rect 14311 25208 14711 25256
rect 14888 25545 15288 25608
rect 14888 25256 14947 25545
rect 15221 25256 15288 25545
rect 14888 25208 15288 25256
rect 15465 25545 15865 25608
rect 15465 25256 15524 25545
rect 15798 25256 15865 25545
rect 15465 25208 15865 25256
rect 16042 25545 16442 25608
rect 16042 25256 16101 25545
rect 16375 25256 16442 25545
rect 16042 25208 16442 25256
rect 16619 25545 17019 25608
rect 16619 25256 16678 25545
rect 16952 25256 17019 25545
rect 16619 25208 17019 25256
rect 17196 25545 17596 25608
rect 17196 25256 17255 25545
rect 17529 25256 17596 25545
rect 17196 25208 17596 25256
rect 17773 25545 18173 25608
rect 17773 25256 17832 25545
rect 18106 25256 18173 25545
rect 17773 25208 18173 25256
rect 18350 25545 18750 25608
rect 18350 25256 18409 25545
rect 18683 25256 18750 25545
rect 18350 25208 18750 25256
rect 18927 25545 19327 25608
rect 18927 25256 18986 25545
rect 19260 25256 19327 25545
rect 18927 25208 19327 25256
rect 19504 25545 19904 25608
rect 19504 25256 19563 25545
rect 19837 25256 19904 25545
rect 19504 25208 19904 25256
rect 20081 25545 20481 25608
rect 20081 25256 20140 25545
rect 20414 25256 20481 25545
rect 20081 25208 20481 25256
rect 20658 25545 21058 25608
rect 20658 25256 20717 25545
rect 20991 25256 21058 25545
rect 20658 25208 21058 25256
rect 21235 25545 21635 25608
rect 21235 25256 21294 25545
rect 21568 25256 21635 25545
rect 21235 25208 21635 25256
rect 21812 25545 22212 25608
rect 21812 25256 21871 25545
rect 22145 25256 22212 25545
rect 21812 25208 22212 25256
rect 22389 25545 22789 25608
rect 22389 25256 22448 25545
rect 22722 25256 22789 25545
rect 22389 25208 22789 25256
rect 22966 25545 23366 25608
rect 22966 25256 23025 25545
rect 23299 25256 23366 25545
rect 22966 25208 23366 25256
rect 23543 25545 23943 25608
rect 23543 25256 23602 25545
rect 23876 25256 23943 25545
rect 23543 25208 23943 25256
rect 24120 25545 24520 25608
rect 24120 25256 24179 25545
rect 24453 25256 24520 25545
rect 24120 25208 24520 25256
rect 24697 25545 25097 25608
rect 24697 25256 24756 25545
rect 25030 25256 25097 25545
rect 24697 25208 25097 25256
rect 25274 25545 25674 25608
rect 25274 25256 25333 25545
rect 25607 25256 25674 25545
rect 25274 25208 25674 25256
rect 25851 25545 26251 25608
rect 25851 25256 25910 25545
rect 26184 25256 26251 25545
rect 25851 25208 26251 25256
rect 26428 25545 26828 25608
rect 26428 25256 26487 25545
rect 26761 25256 26828 25545
rect 26428 25208 26828 25256
rect 27005 25545 27405 25608
rect 27005 25256 27064 25545
rect 27338 25256 27405 25545
rect 27005 25208 27405 25256
rect 27582 25545 27982 25608
rect 27582 25256 27641 25545
rect 27915 25256 27982 25545
rect 27582 25208 27982 25256
rect 28159 25545 28559 25608
rect 28159 25256 28218 25545
rect 28492 25256 28559 25545
rect 28159 25208 28559 25256
rect 28736 25545 29136 25608
rect 28736 25256 28795 25545
rect 29069 25256 29136 25545
rect 28736 25208 29136 25256
rect 29313 25545 29713 25608
rect 29313 25256 29372 25545
rect 29646 25256 29713 25545
rect 29313 25208 29713 25256
rect 29890 25545 30290 25608
rect 29890 25256 29949 25545
rect 30223 25256 30290 25545
rect 29890 25208 30290 25256
rect 30467 25545 30867 25608
rect 30467 25256 30526 25545
rect 30800 25256 30867 25545
rect 30467 25208 30867 25256
rect 31044 25545 31444 25608
rect 31044 25256 31103 25545
rect 31377 25256 31444 25545
rect 31044 25208 31444 25256
rect 31621 25545 32021 25608
rect 31621 25256 31680 25545
rect 31954 25256 32021 25545
rect 31621 25208 32021 25256
rect 32198 25545 32598 25608
rect 32198 25256 32257 25545
rect 32531 25256 32598 25545
rect 32198 25208 32598 25256
rect 32775 25545 33175 25608
rect 32775 25256 32834 25545
rect 33108 25256 33175 25545
rect 32775 25208 33175 25256
rect 33352 25545 33752 25608
rect 33352 25256 33411 25545
rect 33685 25256 33752 25545
rect 33352 25208 33752 25256
rect 33929 25545 34329 25608
rect 33929 25256 33988 25545
rect 34262 25256 34329 25545
rect 33929 25208 34329 25256
rect 34506 25545 34906 25608
rect 34506 25256 34565 25545
rect 34839 25256 34906 25545
rect 34506 25208 34906 25256
rect 35083 25545 35483 25608
rect 35083 25256 35142 25545
rect 35416 25256 35483 25545
rect 35083 25208 35483 25256
rect 35660 25545 36060 25608
rect 35660 25256 35719 25545
rect 35993 25256 36060 25545
rect 35660 25208 36060 25256
rect 36237 25545 36637 25608
rect 36237 25256 36296 25545
rect 36570 25256 36637 25545
rect 36237 25208 36637 25256
rect 36814 25545 37214 25608
rect 36814 25256 36873 25545
rect 37147 25256 37214 25545
rect 36814 25208 37214 25256
rect 37391 25545 37791 25608
rect 37391 25256 37450 25545
rect 37724 25256 37791 25545
rect 37391 25208 37791 25256
rect 37968 25545 38368 25608
rect 37968 25256 38027 25545
rect 38301 25256 38368 25545
rect 37968 25208 38368 25256
rect 38545 25545 38945 25608
rect 38545 25256 38604 25545
rect 38878 25256 38945 25545
rect 38545 25208 38945 25256
rect 39122 25545 39522 25608
rect 39122 25256 39181 25545
rect 39455 25256 39522 25545
rect 39122 25208 39522 25256
rect 39699 25545 40099 25608
rect 39699 25256 39758 25545
rect 40032 25256 40099 25545
rect 39699 25208 40099 25256
rect 40276 25545 40676 25608
rect 40276 25256 40335 25545
rect 40609 25256 40676 25545
rect 40276 25208 40676 25256
rect 40853 25545 41253 25608
rect 40853 25256 40912 25545
rect 41186 25256 41253 25545
rect 40853 25208 41253 25256
rect 41430 25545 41830 25608
rect 41430 25256 41489 25545
rect 41763 25256 41830 25545
rect 41430 25208 41830 25256
rect 42007 25545 42407 25608
rect 42007 25256 42066 25545
rect 42340 25256 42407 25545
rect 42007 25208 42407 25256
rect 42584 25545 42984 25608
rect 42584 25256 42643 25545
rect 42917 25256 42984 25545
rect 42584 25208 42984 25256
rect 43161 25545 43561 25608
rect 43161 25256 43220 25545
rect 43494 25256 43561 25545
rect 43161 25208 43561 25256
rect 43738 25545 44138 25608
rect 43738 25256 43797 25545
rect 44071 25256 44138 25545
rect 43738 25208 44138 25256
rect 44315 25545 44715 25608
rect 44315 25256 44374 25545
rect 44648 25256 44715 25545
rect 44315 25208 44715 25256
rect 44892 25545 45292 25608
rect 44892 25256 44951 25545
rect 45225 25256 45292 25545
rect 44892 25208 45292 25256
rect 45469 25545 45869 25608
rect 45469 25256 45528 25545
rect 45802 25256 45869 25545
rect 45469 25208 45869 25256
rect 46046 25545 46446 25608
rect 46046 25256 46105 25545
rect 46379 25256 46446 25545
rect 46046 25208 46446 25256
rect 46623 25545 47023 25608
rect 46623 25256 46682 25545
rect 46956 25256 47023 25545
rect 46623 25208 47023 25256
rect 47200 25545 47600 25608
rect 47200 25256 47259 25545
rect 47533 25256 47600 25545
rect 47200 25208 47600 25256
rect 47777 25545 48177 25608
rect 47777 25256 47836 25545
rect 48110 25256 48177 25545
rect 47777 25208 48177 25256
rect 48354 25545 48754 25608
rect 48354 25256 48413 25545
rect 48687 25256 48754 25545
rect 48354 25208 48754 25256
rect 48931 25545 49331 25608
rect 48931 25256 48990 25545
rect 49264 25256 49331 25545
rect 48931 25208 49331 25256
rect 49508 25545 49908 25608
rect 49508 25256 49567 25545
rect 49841 25256 49908 25545
rect 49508 25208 49908 25256
rect 50085 25545 50485 25608
rect 50085 25256 50144 25545
rect 50418 25256 50485 25545
rect 50085 25208 50485 25256
rect 50662 25545 51062 25608
rect 50662 25256 50721 25545
rect 50995 25256 51062 25545
rect 50662 25208 51062 25256
rect 51239 25545 51639 25608
rect 51239 25256 51298 25545
rect 51572 25256 51639 25545
rect 51239 25208 51639 25256
rect 51816 25545 52216 25608
rect 51816 25256 51875 25545
rect 52149 25256 52216 25545
rect 51816 25208 52216 25256
rect 52393 25545 52793 25608
rect 52393 25256 52452 25545
rect 52726 25256 52793 25545
rect 52393 25208 52793 25256
rect 52970 25545 53370 25608
rect 52970 25256 53029 25545
rect 53303 25256 53370 25545
rect 52970 25208 53370 25256
rect 53547 25545 53947 25608
rect 53547 25256 53606 25545
rect 53880 25256 53947 25545
rect 53547 25208 53947 25256
rect 54124 25545 54524 25608
rect 54124 25256 54183 25545
rect 54457 25256 54524 25545
rect 54124 25208 54524 25256
rect 54701 25545 55101 25608
rect 54701 25256 54760 25545
rect 55034 25256 55101 25545
rect 54701 25208 55101 25256
rect 55278 25545 55678 25608
rect 55278 25256 55337 25545
rect 55611 25256 55678 25545
rect 55278 25208 55678 25256
rect 55855 25545 56255 25608
rect 55855 25256 55914 25545
rect 56188 25256 56255 25545
rect 55855 25208 56255 25256
rect -54929 24987 -54529 25050
rect -54929 24698 -54870 24987
rect -54596 24698 -54529 24987
rect -54929 24650 -54529 24698
rect -54352 24987 -53952 25050
rect -54352 24698 -54293 24987
rect -54019 24698 -53952 24987
rect -54352 24650 -53952 24698
rect -53775 24987 -53375 25050
rect -53775 24698 -53716 24987
rect -53442 24698 -53375 24987
rect -53775 24650 -53375 24698
rect -53198 24987 -52798 25050
rect -53198 24698 -53139 24987
rect -52865 24698 -52798 24987
rect -53198 24650 -52798 24698
rect -52621 24987 -52221 25050
rect -52621 24698 -52562 24987
rect -52288 24698 -52221 24987
rect -52621 24650 -52221 24698
rect -52044 24987 -51644 25050
rect -52044 24698 -51985 24987
rect -51711 24698 -51644 24987
rect -52044 24650 -51644 24698
rect -51467 24987 -51067 25050
rect -51467 24698 -51408 24987
rect -51134 24698 -51067 24987
rect -51467 24650 -51067 24698
rect -50890 24987 -50490 25050
rect -50890 24698 -50831 24987
rect -50557 24698 -50490 24987
rect -50890 24650 -50490 24698
rect -50313 24987 -49913 25050
rect -50313 24698 -50254 24987
rect -49980 24698 -49913 24987
rect -50313 24650 -49913 24698
rect -49736 24987 -49336 25050
rect -49736 24698 -49677 24987
rect -49403 24698 -49336 24987
rect -49736 24650 -49336 24698
rect -49159 24987 -48759 25050
rect -49159 24698 -49100 24987
rect -48826 24698 -48759 24987
rect -49159 24650 -48759 24698
rect -48582 24987 -48182 25050
rect -48582 24698 -48523 24987
rect -48249 24698 -48182 24987
rect -48582 24650 -48182 24698
rect -48005 24987 -47605 25050
rect -48005 24698 -47946 24987
rect -47672 24698 -47605 24987
rect -48005 24650 -47605 24698
rect -47428 24987 -47028 25050
rect -47428 24698 -47369 24987
rect -47095 24698 -47028 24987
rect -47428 24650 -47028 24698
rect -46851 24987 -46451 25050
rect -46851 24698 -46792 24987
rect -46518 24698 -46451 24987
rect -46851 24650 -46451 24698
rect -46274 24987 -45874 25050
rect -46274 24698 -46215 24987
rect -45941 24698 -45874 24987
rect -46274 24650 -45874 24698
rect -45697 24987 -45297 25050
rect -45697 24698 -45638 24987
rect -45364 24698 -45297 24987
rect -45697 24650 -45297 24698
rect -45120 24987 -44720 25050
rect -45120 24698 -45061 24987
rect -44787 24698 -44720 24987
rect -45120 24650 -44720 24698
rect -44543 24987 -44143 25050
rect -44543 24698 -44484 24987
rect -44210 24698 -44143 24987
rect -44543 24650 -44143 24698
rect -43966 24987 -43566 25050
rect -43966 24698 -43907 24987
rect -43633 24698 -43566 24987
rect -43966 24650 -43566 24698
rect -43389 24987 -42989 25050
rect -43389 24698 -43330 24987
rect -43056 24698 -42989 24987
rect -43389 24650 -42989 24698
rect -42812 24987 -42412 25050
rect -42812 24698 -42753 24987
rect -42479 24698 -42412 24987
rect -42812 24650 -42412 24698
rect -42235 24987 -41835 25050
rect -42235 24698 -42176 24987
rect -41902 24698 -41835 24987
rect -42235 24650 -41835 24698
rect -41658 24987 -41258 25050
rect -41658 24698 -41599 24987
rect -41325 24698 -41258 24987
rect -41658 24650 -41258 24698
rect -41081 24987 -40681 25050
rect -41081 24698 -41022 24987
rect -40748 24698 -40681 24987
rect -41081 24650 -40681 24698
rect -40504 24987 -40104 25050
rect -40504 24698 -40445 24987
rect -40171 24698 -40104 24987
rect -40504 24650 -40104 24698
rect -39927 24987 -39527 25050
rect -39927 24698 -39868 24987
rect -39594 24698 -39527 24987
rect -39927 24650 -39527 24698
rect -39350 24987 -38950 25050
rect -39350 24698 -39291 24987
rect -39017 24698 -38950 24987
rect -39350 24650 -38950 24698
rect -38773 24987 -38373 25050
rect -38773 24698 -38714 24987
rect -38440 24698 -38373 24987
rect -38773 24650 -38373 24698
rect -38196 24987 -37796 25050
rect -38196 24698 -38137 24987
rect -37863 24698 -37796 24987
rect -38196 24650 -37796 24698
rect -37619 24987 -37219 25050
rect -37619 24698 -37560 24987
rect -37286 24698 -37219 24987
rect -37619 24650 -37219 24698
rect -37042 24987 -36642 25050
rect -37042 24698 -36983 24987
rect -36709 24698 -36642 24987
rect -37042 24650 -36642 24698
rect -36465 24987 -36065 25050
rect -36465 24698 -36406 24987
rect -36132 24698 -36065 24987
rect -36465 24650 -36065 24698
rect -35888 24987 -35488 25050
rect -35888 24698 -35829 24987
rect -35555 24698 -35488 24987
rect -35888 24650 -35488 24698
rect -35311 24987 -34911 25050
rect -35311 24698 -35252 24987
rect -34978 24698 -34911 24987
rect -35311 24650 -34911 24698
rect -34734 24987 -34334 25050
rect -34734 24698 -34675 24987
rect -34401 24698 -34334 24987
rect -34734 24650 -34334 24698
rect -34157 24987 -33757 25050
rect -34157 24698 -34098 24987
rect -33824 24698 -33757 24987
rect -34157 24650 -33757 24698
rect -33580 24987 -33180 25050
rect -33580 24698 -33521 24987
rect -33247 24698 -33180 24987
rect -33580 24650 -33180 24698
rect -33003 24987 -32603 25050
rect -33003 24698 -32944 24987
rect -32670 24698 -32603 24987
rect -33003 24650 -32603 24698
rect -32426 24987 -32026 25050
rect -32426 24698 -32367 24987
rect -32093 24698 -32026 24987
rect -32426 24650 -32026 24698
rect -31849 24987 -31449 25050
rect -31849 24698 -31790 24987
rect -31516 24698 -31449 24987
rect -31849 24650 -31449 24698
rect -31272 24987 -30872 25050
rect -31272 24698 -31213 24987
rect -30939 24698 -30872 24987
rect -31272 24650 -30872 24698
rect -30695 24987 -30295 25050
rect -30695 24698 -30636 24987
rect -30362 24698 -30295 24987
rect -30695 24650 -30295 24698
rect -30118 24987 -29718 25050
rect -30118 24698 -30059 24987
rect -29785 24698 -29718 24987
rect -30118 24650 -29718 24698
rect -29541 24987 -29141 25050
rect -29541 24698 -29482 24987
rect -29208 24698 -29141 24987
rect -29541 24650 -29141 24698
rect -28964 24987 -28564 25050
rect -28964 24698 -28905 24987
rect -28631 24698 -28564 24987
rect -28964 24650 -28564 24698
rect -28387 24987 -27987 25050
rect -28387 24698 -28328 24987
rect -28054 24698 -27987 24987
rect -28387 24650 -27987 24698
rect -27810 24987 -27410 25050
rect -27810 24698 -27751 24987
rect -27477 24698 -27410 24987
rect -27810 24650 -27410 24698
rect -27233 24987 -26833 25050
rect -27233 24698 -27174 24987
rect -26900 24698 -26833 24987
rect -27233 24650 -26833 24698
rect -26656 24987 -26256 25050
rect -26656 24698 -26597 24987
rect -26323 24698 -26256 24987
rect -26656 24650 -26256 24698
rect -26079 24987 -25679 25050
rect -26079 24698 -26020 24987
rect -25746 24698 -25679 24987
rect -26079 24650 -25679 24698
rect -25502 24987 -25102 25050
rect -25502 24698 -25443 24987
rect -25169 24698 -25102 24987
rect -25502 24650 -25102 24698
rect -24925 24987 -24525 25050
rect -24925 24698 -24866 24987
rect -24592 24698 -24525 24987
rect -24925 24650 -24525 24698
rect -24348 24987 -23948 25050
rect -24348 24698 -24289 24987
rect -24015 24698 -23948 24987
rect -24348 24650 -23948 24698
rect -23771 24987 -23371 25050
rect -23771 24698 -23712 24987
rect -23438 24698 -23371 24987
rect -23771 24650 -23371 24698
rect -23194 24987 -22794 25050
rect -23194 24698 -23135 24987
rect -22861 24698 -22794 24987
rect -23194 24650 -22794 24698
rect -22617 24987 -22217 25050
rect -22617 24698 -22558 24987
rect -22284 24698 -22217 24987
rect -22617 24650 -22217 24698
rect -22040 24987 -21640 25050
rect -22040 24698 -21981 24987
rect -21707 24698 -21640 24987
rect -22040 24650 -21640 24698
rect -21463 24987 -21063 25050
rect -21463 24698 -21404 24987
rect -21130 24698 -21063 24987
rect -21463 24650 -21063 24698
rect -20886 24987 -20486 25050
rect -20886 24698 -20827 24987
rect -20553 24698 -20486 24987
rect -20886 24650 -20486 24698
rect -20309 24987 -19909 25050
rect -20309 24698 -20250 24987
rect -19976 24698 -19909 24987
rect -20309 24650 -19909 24698
rect -19732 24987 -19332 25050
rect -19732 24698 -19673 24987
rect -19399 24698 -19332 24987
rect -19732 24650 -19332 24698
rect -19155 24987 -18755 25050
rect -19155 24698 -19096 24987
rect -18822 24698 -18755 24987
rect -19155 24650 -18755 24698
rect -18578 24987 -18178 25050
rect -18578 24698 -18519 24987
rect -18245 24698 -18178 24987
rect -18578 24650 -18178 24698
rect -18001 24987 -17601 25050
rect -18001 24698 -17942 24987
rect -17668 24698 -17601 24987
rect -18001 24650 -17601 24698
rect -17424 24987 -17024 25050
rect -17424 24698 -17365 24987
rect -17091 24698 -17024 24987
rect -17424 24650 -17024 24698
rect -16847 24987 -16447 25050
rect -16847 24698 -16788 24987
rect -16514 24698 -16447 24987
rect -16847 24650 -16447 24698
rect -16270 24987 -15870 25050
rect -16270 24698 -16211 24987
rect -15937 24698 -15870 24987
rect -16270 24650 -15870 24698
rect -15693 24987 -15293 25050
rect -15693 24698 -15634 24987
rect -15360 24698 -15293 24987
rect -15693 24650 -15293 24698
rect -15116 24987 -14716 25050
rect -15116 24698 -15057 24987
rect -14783 24698 -14716 24987
rect -15116 24650 -14716 24698
rect -14539 24987 -14139 25050
rect -14539 24698 -14480 24987
rect -14206 24698 -14139 24987
rect -14539 24650 -14139 24698
rect -13962 24987 -13562 25050
rect -13962 24698 -13903 24987
rect -13629 24698 -13562 24987
rect -13962 24650 -13562 24698
rect -13385 24987 -12985 25050
rect -13385 24698 -13326 24987
rect -13052 24698 -12985 24987
rect -13385 24650 -12985 24698
rect -12808 24987 -12408 25050
rect -12808 24698 -12749 24987
rect -12475 24698 -12408 24987
rect -12808 24650 -12408 24698
rect -12231 24987 -11831 25050
rect -12231 24698 -12172 24987
rect -11898 24698 -11831 24987
rect -12231 24650 -11831 24698
rect -11654 24987 -11254 25050
rect -11654 24698 -11595 24987
rect -11321 24698 -11254 24987
rect -11654 24650 -11254 24698
rect -11077 24987 -10677 25050
rect -11077 24698 -11018 24987
rect -10744 24698 -10677 24987
rect -11077 24650 -10677 24698
rect -10500 24987 -10100 25050
rect -10500 24698 -10441 24987
rect -10167 24698 -10100 24987
rect -10500 24650 -10100 24698
rect -9923 24987 -9523 25050
rect -9923 24698 -9864 24987
rect -9590 24698 -9523 24987
rect -9923 24650 -9523 24698
rect -9346 24987 -8946 25050
rect -9346 24698 -9287 24987
rect -9013 24698 -8946 24987
rect -9346 24650 -8946 24698
rect -8769 24987 -8369 25050
rect -8769 24698 -8710 24987
rect -8436 24698 -8369 24987
rect -8769 24650 -8369 24698
rect -8192 24987 -7792 25050
rect -8192 24698 -8133 24987
rect -7859 24698 -7792 24987
rect -8192 24650 -7792 24698
rect -7615 24987 -7215 25050
rect -7615 24698 -7556 24987
rect -7282 24698 -7215 24987
rect -7615 24650 -7215 24698
rect -7038 24987 -6638 25050
rect -7038 24698 -6979 24987
rect -6705 24698 -6638 24987
rect -7038 24650 -6638 24698
rect -6461 24987 -6061 25050
rect -6461 24698 -6402 24987
rect -6128 24698 -6061 24987
rect -6461 24650 -6061 24698
rect -5884 24987 -5484 25050
rect -5884 24698 -5825 24987
rect -5551 24698 -5484 24987
rect -5884 24650 -5484 24698
rect -5307 24987 -4907 25050
rect -5307 24698 -5248 24987
rect -4974 24698 -4907 24987
rect -5307 24650 -4907 24698
rect -4730 24987 -4330 25050
rect -4730 24698 -4671 24987
rect -4397 24698 -4330 24987
rect -4730 24650 -4330 24698
rect -4153 24987 -3753 25050
rect -4153 24698 -4094 24987
rect -3820 24698 -3753 24987
rect -4153 24650 -3753 24698
rect -3576 24987 -3176 25050
rect -3576 24698 -3517 24987
rect -3243 24698 -3176 24987
rect -3576 24650 -3176 24698
rect -2999 24987 -2599 25050
rect -2999 24698 -2940 24987
rect -2666 24698 -2599 24987
rect -2999 24650 -2599 24698
rect -2422 24987 -2022 25050
rect -2422 24698 -2363 24987
rect -2089 24698 -2022 24987
rect -2422 24650 -2022 24698
rect -1845 24987 -1445 25050
rect -1845 24698 -1786 24987
rect -1512 24698 -1445 24987
rect -1845 24650 -1445 24698
rect -1268 24987 -868 25050
rect -1268 24698 -1209 24987
rect -935 24698 -868 24987
rect -1268 24650 -868 24698
rect -691 24987 -291 25050
rect -691 24698 -632 24987
rect -358 24698 -291 24987
rect -691 24650 -291 24698
rect -114 24987 286 25050
rect -114 24698 -55 24987
rect 219 24698 286 24987
rect -114 24650 286 24698
rect 463 24987 863 25050
rect 463 24698 522 24987
rect 796 24698 863 24987
rect 463 24650 863 24698
rect 1040 24987 1440 25050
rect 1040 24698 1099 24987
rect 1373 24698 1440 24987
rect 1040 24650 1440 24698
rect 1617 24987 2017 25050
rect 1617 24698 1676 24987
rect 1950 24698 2017 24987
rect 1617 24650 2017 24698
rect 2194 24987 2594 25050
rect 2194 24698 2253 24987
rect 2527 24698 2594 24987
rect 2194 24650 2594 24698
rect 2771 24987 3171 25050
rect 2771 24698 2830 24987
rect 3104 24698 3171 24987
rect 2771 24650 3171 24698
rect 3348 24987 3748 25050
rect 3348 24698 3407 24987
rect 3681 24698 3748 24987
rect 3348 24650 3748 24698
rect 3925 24987 4325 25050
rect 3925 24698 3984 24987
rect 4258 24698 4325 24987
rect 3925 24650 4325 24698
rect 4502 24987 4902 25050
rect 4502 24698 4561 24987
rect 4835 24698 4902 24987
rect 4502 24650 4902 24698
rect 5079 24987 5479 25050
rect 5079 24698 5138 24987
rect 5412 24698 5479 24987
rect 5079 24650 5479 24698
rect 5656 24987 6056 25050
rect 5656 24698 5715 24987
rect 5989 24698 6056 24987
rect 5656 24650 6056 24698
rect 6233 24987 6633 25050
rect 6233 24698 6292 24987
rect 6566 24698 6633 24987
rect 6233 24650 6633 24698
rect 6810 24987 7210 25050
rect 6810 24698 6869 24987
rect 7143 24698 7210 24987
rect 6810 24650 7210 24698
rect 7387 24987 7787 25050
rect 7387 24698 7446 24987
rect 7720 24698 7787 24987
rect 7387 24650 7787 24698
rect 7964 24987 8364 25050
rect 7964 24698 8023 24987
rect 8297 24698 8364 24987
rect 7964 24650 8364 24698
rect 8541 24987 8941 25050
rect 8541 24698 8600 24987
rect 8874 24698 8941 24987
rect 8541 24650 8941 24698
rect 9118 24987 9518 25050
rect 9118 24698 9177 24987
rect 9451 24698 9518 24987
rect 9118 24650 9518 24698
rect 9695 24987 10095 25050
rect 9695 24698 9754 24987
rect 10028 24698 10095 24987
rect 9695 24650 10095 24698
rect 10272 24987 10672 25050
rect 10272 24698 10331 24987
rect 10605 24698 10672 24987
rect 10272 24650 10672 24698
rect 10849 24987 11249 25050
rect 10849 24698 10908 24987
rect 11182 24698 11249 24987
rect 10849 24650 11249 24698
rect 11426 24987 11826 25050
rect 11426 24698 11485 24987
rect 11759 24698 11826 24987
rect 11426 24650 11826 24698
rect 12003 24987 12403 25050
rect 12003 24698 12062 24987
rect 12336 24698 12403 24987
rect 12003 24650 12403 24698
rect 12580 24987 12980 25050
rect 12580 24698 12639 24987
rect 12913 24698 12980 24987
rect 12580 24650 12980 24698
rect 13157 24987 13557 25050
rect 13157 24698 13216 24987
rect 13490 24698 13557 24987
rect 13157 24650 13557 24698
rect 13734 24987 14134 25050
rect 13734 24698 13793 24987
rect 14067 24698 14134 24987
rect 13734 24650 14134 24698
rect 14311 24987 14711 25050
rect 14311 24698 14370 24987
rect 14644 24698 14711 24987
rect 14311 24650 14711 24698
rect 14888 24987 15288 25050
rect 14888 24698 14947 24987
rect 15221 24698 15288 24987
rect 14888 24650 15288 24698
rect 15465 24987 15865 25050
rect 15465 24698 15524 24987
rect 15798 24698 15865 24987
rect 15465 24650 15865 24698
rect 16042 24987 16442 25050
rect 16042 24698 16101 24987
rect 16375 24698 16442 24987
rect 16042 24650 16442 24698
rect 16619 24987 17019 25050
rect 16619 24698 16678 24987
rect 16952 24698 17019 24987
rect 16619 24650 17019 24698
rect 17196 24987 17596 25050
rect 17196 24698 17255 24987
rect 17529 24698 17596 24987
rect 17196 24650 17596 24698
rect 17773 24987 18173 25050
rect 17773 24698 17832 24987
rect 18106 24698 18173 24987
rect 17773 24650 18173 24698
rect 18350 24987 18750 25050
rect 18350 24698 18409 24987
rect 18683 24698 18750 24987
rect 18350 24650 18750 24698
rect 18927 24987 19327 25050
rect 18927 24698 18986 24987
rect 19260 24698 19327 24987
rect 18927 24650 19327 24698
rect 19504 24987 19904 25050
rect 19504 24698 19563 24987
rect 19837 24698 19904 24987
rect 19504 24650 19904 24698
rect 20081 24987 20481 25050
rect 20081 24698 20140 24987
rect 20414 24698 20481 24987
rect 20081 24650 20481 24698
rect 20658 24987 21058 25050
rect 20658 24698 20717 24987
rect 20991 24698 21058 24987
rect 20658 24650 21058 24698
rect 21235 24987 21635 25050
rect 21235 24698 21294 24987
rect 21568 24698 21635 24987
rect 21235 24650 21635 24698
rect 21812 24987 22212 25050
rect 21812 24698 21871 24987
rect 22145 24698 22212 24987
rect 21812 24650 22212 24698
rect 22389 24987 22789 25050
rect 22389 24698 22448 24987
rect 22722 24698 22789 24987
rect 22389 24650 22789 24698
rect 22966 24987 23366 25050
rect 22966 24698 23025 24987
rect 23299 24698 23366 24987
rect 22966 24650 23366 24698
rect 23543 24987 23943 25050
rect 23543 24698 23602 24987
rect 23876 24698 23943 24987
rect 23543 24650 23943 24698
rect 24120 24987 24520 25050
rect 24120 24698 24179 24987
rect 24453 24698 24520 24987
rect 24120 24650 24520 24698
rect 24697 24987 25097 25050
rect 24697 24698 24756 24987
rect 25030 24698 25097 24987
rect 24697 24650 25097 24698
rect 25274 24987 25674 25050
rect 25274 24698 25333 24987
rect 25607 24698 25674 24987
rect 25274 24650 25674 24698
rect 25851 24987 26251 25050
rect 25851 24698 25910 24987
rect 26184 24698 26251 24987
rect 25851 24650 26251 24698
rect 26428 24987 26828 25050
rect 26428 24698 26487 24987
rect 26761 24698 26828 24987
rect 26428 24650 26828 24698
rect 27005 24987 27405 25050
rect 27005 24698 27064 24987
rect 27338 24698 27405 24987
rect 27005 24650 27405 24698
rect 27582 24987 27982 25050
rect 27582 24698 27641 24987
rect 27915 24698 27982 24987
rect 27582 24650 27982 24698
rect 28159 24987 28559 25050
rect 28159 24698 28218 24987
rect 28492 24698 28559 24987
rect 28159 24650 28559 24698
rect 28736 24987 29136 25050
rect 28736 24698 28795 24987
rect 29069 24698 29136 24987
rect 28736 24650 29136 24698
rect 29313 24987 29713 25050
rect 29313 24698 29372 24987
rect 29646 24698 29713 24987
rect 29313 24650 29713 24698
rect 29890 24987 30290 25050
rect 29890 24698 29949 24987
rect 30223 24698 30290 24987
rect 29890 24650 30290 24698
rect 30467 24987 30867 25050
rect 30467 24698 30526 24987
rect 30800 24698 30867 24987
rect 30467 24650 30867 24698
rect 31044 24987 31444 25050
rect 31044 24698 31103 24987
rect 31377 24698 31444 24987
rect 31044 24650 31444 24698
rect 31621 24987 32021 25050
rect 31621 24698 31680 24987
rect 31954 24698 32021 24987
rect 31621 24650 32021 24698
rect 32198 24987 32598 25050
rect 32198 24698 32257 24987
rect 32531 24698 32598 24987
rect 32198 24650 32598 24698
rect 32775 24987 33175 25050
rect 32775 24698 32834 24987
rect 33108 24698 33175 24987
rect 32775 24650 33175 24698
rect 33352 24987 33752 25050
rect 33352 24698 33411 24987
rect 33685 24698 33752 24987
rect 33352 24650 33752 24698
rect 33929 24987 34329 25050
rect 33929 24698 33988 24987
rect 34262 24698 34329 24987
rect 33929 24650 34329 24698
rect 34506 24987 34906 25050
rect 34506 24698 34565 24987
rect 34839 24698 34906 24987
rect 34506 24650 34906 24698
rect 35083 24987 35483 25050
rect 35083 24698 35142 24987
rect 35416 24698 35483 24987
rect 35083 24650 35483 24698
rect 35660 24987 36060 25050
rect 35660 24698 35719 24987
rect 35993 24698 36060 24987
rect 35660 24650 36060 24698
rect 36237 24987 36637 25050
rect 36237 24698 36296 24987
rect 36570 24698 36637 24987
rect 36237 24650 36637 24698
rect 36814 24987 37214 25050
rect 36814 24698 36873 24987
rect 37147 24698 37214 24987
rect 36814 24650 37214 24698
rect 37391 24987 37791 25050
rect 37391 24698 37450 24987
rect 37724 24698 37791 24987
rect 37391 24650 37791 24698
rect 37968 24987 38368 25050
rect 37968 24698 38027 24987
rect 38301 24698 38368 24987
rect 37968 24650 38368 24698
rect 38545 24987 38945 25050
rect 38545 24698 38604 24987
rect 38878 24698 38945 24987
rect 38545 24650 38945 24698
rect 39122 24987 39522 25050
rect 39122 24698 39181 24987
rect 39455 24698 39522 24987
rect 39122 24650 39522 24698
rect 39699 24987 40099 25050
rect 39699 24698 39758 24987
rect 40032 24698 40099 24987
rect 39699 24650 40099 24698
rect 40276 24987 40676 25050
rect 40276 24698 40335 24987
rect 40609 24698 40676 24987
rect 40276 24650 40676 24698
rect 40853 24987 41253 25050
rect 40853 24698 40912 24987
rect 41186 24698 41253 24987
rect 40853 24650 41253 24698
rect 41430 24987 41830 25050
rect 41430 24698 41489 24987
rect 41763 24698 41830 24987
rect 41430 24650 41830 24698
rect 42007 24987 42407 25050
rect 42007 24698 42066 24987
rect 42340 24698 42407 24987
rect 42007 24650 42407 24698
rect 42584 24987 42984 25050
rect 42584 24698 42643 24987
rect 42917 24698 42984 24987
rect 42584 24650 42984 24698
rect 43161 24987 43561 25050
rect 43161 24698 43220 24987
rect 43494 24698 43561 24987
rect 43161 24650 43561 24698
rect 43738 24987 44138 25050
rect 43738 24698 43797 24987
rect 44071 24698 44138 24987
rect 43738 24650 44138 24698
rect 44315 24987 44715 25050
rect 44315 24698 44374 24987
rect 44648 24698 44715 24987
rect 44315 24650 44715 24698
rect 44892 24987 45292 25050
rect 44892 24698 44951 24987
rect 45225 24698 45292 24987
rect 44892 24650 45292 24698
rect 45469 24987 45869 25050
rect 45469 24698 45528 24987
rect 45802 24698 45869 24987
rect 45469 24650 45869 24698
rect 46046 24987 46446 25050
rect 46046 24698 46105 24987
rect 46379 24698 46446 24987
rect 46046 24650 46446 24698
rect 46623 24987 47023 25050
rect 46623 24698 46682 24987
rect 46956 24698 47023 24987
rect 46623 24650 47023 24698
rect 47200 24987 47600 25050
rect 47200 24698 47259 24987
rect 47533 24698 47600 24987
rect 47200 24650 47600 24698
rect 47777 24987 48177 25050
rect 47777 24698 47836 24987
rect 48110 24698 48177 24987
rect 47777 24650 48177 24698
rect 48354 24987 48754 25050
rect 48354 24698 48413 24987
rect 48687 24698 48754 24987
rect 48354 24650 48754 24698
rect 48931 24987 49331 25050
rect 48931 24698 48990 24987
rect 49264 24698 49331 24987
rect 48931 24650 49331 24698
rect 49508 24987 49908 25050
rect 49508 24698 49567 24987
rect 49841 24698 49908 24987
rect 49508 24650 49908 24698
rect 50085 24987 50485 25050
rect 50085 24698 50144 24987
rect 50418 24698 50485 24987
rect 50085 24650 50485 24698
rect 50662 24987 51062 25050
rect 50662 24698 50721 24987
rect 50995 24698 51062 24987
rect 50662 24650 51062 24698
rect 51239 24987 51639 25050
rect 51239 24698 51298 24987
rect 51572 24698 51639 24987
rect 51239 24650 51639 24698
rect 51816 24987 52216 25050
rect 51816 24698 51875 24987
rect 52149 24698 52216 24987
rect 51816 24650 52216 24698
rect 52393 24987 52793 25050
rect 52393 24698 52452 24987
rect 52726 24698 52793 24987
rect 52393 24650 52793 24698
rect 52970 24987 53370 25050
rect 52970 24698 53029 24987
rect 53303 24698 53370 24987
rect 52970 24650 53370 24698
rect 53547 24987 53947 25050
rect 53547 24698 53606 24987
rect 53880 24698 53947 24987
rect 53547 24650 53947 24698
rect 54124 24987 54524 25050
rect 54124 24698 54183 24987
rect 54457 24698 54524 24987
rect 54124 24650 54524 24698
rect 54701 24987 55101 25050
rect 54701 24698 54760 24987
rect 55034 24698 55101 24987
rect 54701 24650 55101 24698
rect 55278 24987 55678 25050
rect 55278 24698 55337 24987
rect 55611 24698 55678 24987
rect 55278 24650 55678 24698
rect 55855 24987 56255 25050
rect 55855 24698 55914 24987
rect 56188 24698 56255 24987
rect 55855 24650 56255 24698
rect -54929 24429 -54529 24492
rect -54929 24140 -54870 24429
rect -54596 24140 -54529 24429
rect -54929 24092 -54529 24140
rect -54352 24429 -53952 24492
rect -54352 24140 -54293 24429
rect -54019 24140 -53952 24429
rect -54352 24092 -53952 24140
rect -53775 24429 -53375 24492
rect -53775 24140 -53716 24429
rect -53442 24140 -53375 24429
rect -53775 24092 -53375 24140
rect -53198 24429 -52798 24492
rect -53198 24140 -53139 24429
rect -52865 24140 -52798 24429
rect -53198 24092 -52798 24140
rect -52621 24429 -52221 24492
rect -52621 24140 -52562 24429
rect -52288 24140 -52221 24429
rect -52621 24092 -52221 24140
rect -52044 24429 -51644 24492
rect -52044 24140 -51985 24429
rect -51711 24140 -51644 24429
rect -52044 24092 -51644 24140
rect -51467 24429 -51067 24492
rect -51467 24140 -51408 24429
rect -51134 24140 -51067 24429
rect -51467 24092 -51067 24140
rect -50890 24429 -50490 24492
rect -50890 24140 -50831 24429
rect -50557 24140 -50490 24429
rect -50890 24092 -50490 24140
rect -50313 24429 -49913 24492
rect -50313 24140 -50254 24429
rect -49980 24140 -49913 24429
rect -50313 24092 -49913 24140
rect -49736 24429 -49336 24492
rect -49736 24140 -49677 24429
rect -49403 24140 -49336 24429
rect -49736 24092 -49336 24140
rect -49159 24429 -48759 24492
rect -49159 24140 -49100 24429
rect -48826 24140 -48759 24429
rect -49159 24092 -48759 24140
rect -48582 24429 -48182 24492
rect -48582 24140 -48523 24429
rect -48249 24140 -48182 24429
rect -48582 24092 -48182 24140
rect -48005 24429 -47605 24492
rect -48005 24140 -47946 24429
rect -47672 24140 -47605 24429
rect -48005 24092 -47605 24140
rect -47428 24429 -47028 24492
rect -47428 24140 -47369 24429
rect -47095 24140 -47028 24429
rect -47428 24092 -47028 24140
rect -46851 24429 -46451 24492
rect -46851 24140 -46792 24429
rect -46518 24140 -46451 24429
rect -46851 24092 -46451 24140
rect -46274 24429 -45874 24492
rect -46274 24140 -46215 24429
rect -45941 24140 -45874 24429
rect -46274 24092 -45874 24140
rect -45697 24429 -45297 24492
rect -45697 24140 -45638 24429
rect -45364 24140 -45297 24429
rect -45697 24092 -45297 24140
rect -45120 24429 -44720 24492
rect -45120 24140 -45061 24429
rect -44787 24140 -44720 24429
rect -45120 24092 -44720 24140
rect -44543 24429 -44143 24492
rect -44543 24140 -44484 24429
rect -44210 24140 -44143 24429
rect -44543 24092 -44143 24140
rect -43966 24429 -43566 24492
rect -43966 24140 -43907 24429
rect -43633 24140 -43566 24429
rect -43966 24092 -43566 24140
rect -43389 24429 -42989 24492
rect -43389 24140 -43330 24429
rect -43056 24140 -42989 24429
rect -43389 24092 -42989 24140
rect -42812 24429 -42412 24492
rect -42812 24140 -42753 24429
rect -42479 24140 -42412 24429
rect -42812 24092 -42412 24140
rect -42235 24429 -41835 24492
rect -42235 24140 -42176 24429
rect -41902 24140 -41835 24429
rect -42235 24092 -41835 24140
rect -41658 24429 -41258 24492
rect -41658 24140 -41599 24429
rect -41325 24140 -41258 24429
rect -41658 24092 -41258 24140
rect -41081 24429 -40681 24492
rect -41081 24140 -41022 24429
rect -40748 24140 -40681 24429
rect -41081 24092 -40681 24140
rect -40504 24429 -40104 24492
rect -40504 24140 -40445 24429
rect -40171 24140 -40104 24429
rect -40504 24092 -40104 24140
rect -39927 24429 -39527 24492
rect -39927 24140 -39868 24429
rect -39594 24140 -39527 24429
rect -39927 24092 -39527 24140
rect -39350 24429 -38950 24492
rect -39350 24140 -39291 24429
rect -39017 24140 -38950 24429
rect -39350 24092 -38950 24140
rect -38773 24429 -38373 24492
rect -38773 24140 -38714 24429
rect -38440 24140 -38373 24429
rect -38773 24092 -38373 24140
rect -38196 24429 -37796 24492
rect -38196 24140 -38137 24429
rect -37863 24140 -37796 24429
rect -38196 24092 -37796 24140
rect -37619 24429 -37219 24492
rect -37619 24140 -37560 24429
rect -37286 24140 -37219 24429
rect -37619 24092 -37219 24140
rect -37042 24429 -36642 24492
rect -37042 24140 -36983 24429
rect -36709 24140 -36642 24429
rect -37042 24092 -36642 24140
rect -36465 24429 -36065 24492
rect -36465 24140 -36406 24429
rect -36132 24140 -36065 24429
rect -36465 24092 -36065 24140
rect -35888 24429 -35488 24492
rect -35888 24140 -35829 24429
rect -35555 24140 -35488 24429
rect -35888 24092 -35488 24140
rect -35311 24429 -34911 24492
rect -35311 24140 -35252 24429
rect -34978 24140 -34911 24429
rect -35311 24092 -34911 24140
rect -34734 24429 -34334 24492
rect -34734 24140 -34675 24429
rect -34401 24140 -34334 24429
rect -34734 24092 -34334 24140
rect -34157 24429 -33757 24492
rect -34157 24140 -34098 24429
rect -33824 24140 -33757 24429
rect -34157 24092 -33757 24140
rect -33580 24429 -33180 24492
rect -33580 24140 -33521 24429
rect -33247 24140 -33180 24429
rect -33580 24092 -33180 24140
rect -33003 24429 -32603 24492
rect -33003 24140 -32944 24429
rect -32670 24140 -32603 24429
rect -33003 24092 -32603 24140
rect -32426 24429 -32026 24492
rect -32426 24140 -32367 24429
rect -32093 24140 -32026 24429
rect -32426 24092 -32026 24140
rect -31849 24429 -31449 24492
rect -31849 24140 -31790 24429
rect -31516 24140 -31449 24429
rect -31849 24092 -31449 24140
rect -31272 24429 -30872 24492
rect -31272 24140 -31213 24429
rect -30939 24140 -30872 24429
rect -31272 24092 -30872 24140
rect -30695 24429 -30295 24492
rect -30695 24140 -30636 24429
rect -30362 24140 -30295 24429
rect -30695 24092 -30295 24140
rect -30118 24429 -29718 24492
rect -30118 24140 -30059 24429
rect -29785 24140 -29718 24429
rect -30118 24092 -29718 24140
rect -29541 24429 -29141 24492
rect -29541 24140 -29482 24429
rect -29208 24140 -29141 24429
rect -29541 24092 -29141 24140
rect -28964 24429 -28564 24492
rect -28964 24140 -28905 24429
rect -28631 24140 -28564 24429
rect -28964 24092 -28564 24140
rect -28387 24429 -27987 24492
rect -28387 24140 -28328 24429
rect -28054 24140 -27987 24429
rect -28387 24092 -27987 24140
rect -27810 24429 -27410 24492
rect -27810 24140 -27751 24429
rect -27477 24140 -27410 24429
rect -27810 24092 -27410 24140
rect -27233 24429 -26833 24492
rect -27233 24140 -27174 24429
rect -26900 24140 -26833 24429
rect -27233 24092 -26833 24140
rect -26656 24429 -26256 24492
rect -26656 24140 -26597 24429
rect -26323 24140 -26256 24429
rect -26656 24092 -26256 24140
rect -26079 24429 -25679 24492
rect -26079 24140 -26020 24429
rect -25746 24140 -25679 24429
rect -26079 24092 -25679 24140
rect -25502 24429 -25102 24492
rect -25502 24140 -25443 24429
rect -25169 24140 -25102 24429
rect -25502 24092 -25102 24140
rect -24925 24429 -24525 24492
rect -24925 24140 -24866 24429
rect -24592 24140 -24525 24429
rect -24925 24092 -24525 24140
rect -24348 24429 -23948 24492
rect -24348 24140 -24289 24429
rect -24015 24140 -23948 24429
rect -24348 24092 -23948 24140
rect -23771 24429 -23371 24492
rect -23771 24140 -23712 24429
rect -23438 24140 -23371 24429
rect -23771 24092 -23371 24140
rect -23194 24429 -22794 24492
rect -23194 24140 -23135 24429
rect -22861 24140 -22794 24429
rect -23194 24092 -22794 24140
rect -22617 24429 -22217 24492
rect -22617 24140 -22558 24429
rect -22284 24140 -22217 24429
rect -22617 24092 -22217 24140
rect -22040 24429 -21640 24492
rect -22040 24140 -21981 24429
rect -21707 24140 -21640 24429
rect -22040 24092 -21640 24140
rect -21463 24429 -21063 24492
rect -21463 24140 -21404 24429
rect -21130 24140 -21063 24429
rect -21463 24092 -21063 24140
rect -20886 24429 -20486 24492
rect -20886 24140 -20827 24429
rect -20553 24140 -20486 24429
rect -20886 24092 -20486 24140
rect -20309 24429 -19909 24492
rect -20309 24140 -20250 24429
rect -19976 24140 -19909 24429
rect -20309 24092 -19909 24140
rect -19732 24429 -19332 24492
rect -19732 24140 -19673 24429
rect -19399 24140 -19332 24429
rect -19732 24092 -19332 24140
rect -19155 24429 -18755 24492
rect -19155 24140 -19096 24429
rect -18822 24140 -18755 24429
rect -19155 24092 -18755 24140
rect -18578 24429 -18178 24492
rect -18578 24140 -18519 24429
rect -18245 24140 -18178 24429
rect -18578 24092 -18178 24140
rect -18001 24429 -17601 24492
rect -18001 24140 -17942 24429
rect -17668 24140 -17601 24429
rect -18001 24092 -17601 24140
rect -17424 24429 -17024 24492
rect -17424 24140 -17365 24429
rect -17091 24140 -17024 24429
rect -17424 24092 -17024 24140
rect -16847 24429 -16447 24492
rect -16847 24140 -16788 24429
rect -16514 24140 -16447 24429
rect -16847 24092 -16447 24140
rect -16270 24429 -15870 24492
rect -16270 24140 -16211 24429
rect -15937 24140 -15870 24429
rect -16270 24092 -15870 24140
rect -15693 24429 -15293 24492
rect -15693 24140 -15634 24429
rect -15360 24140 -15293 24429
rect -15693 24092 -15293 24140
rect -15116 24429 -14716 24492
rect -15116 24140 -15057 24429
rect -14783 24140 -14716 24429
rect -15116 24092 -14716 24140
rect -14539 24429 -14139 24492
rect -14539 24140 -14480 24429
rect -14206 24140 -14139 24429
rect -14539 24092 -14139 24140
rect -13962 24429 -13562 24492
rect -13962 24140 -13903 24429
rect -13629 24140 -13562 24429
rect -13962 24092 -13562 24140
rect -13385 24429 -12985 24492
rect -13385 24140 -13326 24429
rect -13052 24140 -12985 24429
rect -13385 24092 -12985 24140
rect -12808 24429 -12408 24492
rect -12808 24140 -12749 24429
rect -12475 24140 -12408 24429
rect -12808 24092 -12408 24140
rect -12231 24429 -11831 24492
rect -12231 24140 -12172 24429
rect -11898 24140 -11831 24429
rect -12231 24092 -11831 24140
rect -11654 24429 -11254 24492
rect -11654 24140 -11595 24429
rect -11321 24140 -11254 24429
rect -11654 24092 -11254 24140
rect -11077 24429 -10677 24492
rect -11077 24140 -11018 24429
rect -10744 24140 -10677 24429
rect -11077 24092 -10677 24140
rect -10500 24429 -10100 24492
rect -10500 24140 -10441 24429
rect -10167 24140 -10100 24429
rect -10500 24092 -10100 24140
rect -9923 24429 -9523 24492
rect -9923 24140 -9864 24429
rect -9590 24140 -9523 24429
rect -9923 24092 -9523 24140
rect -9346 24429 -8946 24492
rect -9346 24140 -9287 24429
rect -9013 24140 -8946 24429
rect -9346 24092 -8946 24140
rect -8769 24429 -8369 24492
rect -8769 24140 -8710 24429
rect -8436 24140 -8369 24429
rect -8769 24092 -8369 24140
rect -8192 24429 -7792 24492
rect -8192 24140 -8133 24429
rect -7859 24140 -7792 24429
rect -8192 24092 -7792 24140
rect -7615 24429 -7215 24492
rect -7615 24140 -7556 24429
rect -7282 24140 -7215 24429
rect -7615 24092 -7215 24140
rect -7038 24429 -6638 24492
rect -7038 24140 -6979 24429
rect -6705 24140 -6638 24429
rect -7038 24092 -6638 24140
rect -6461 24429 -6061 24492
rect -6461 24140 -6402 24429
rect -6128 24140 -6061 24429
rect -6461 24092 -6061 24140
rect -5884 24429 -5484 24492
rect -5884 24140 -5825 24429
rect -5551 24140 -5484 24429
rect -5884 24092 -5484 24140
rect -5307 24429 -4907 24492
rect -5307 24140 -5248 24429
rect -4974 24140 -4907 24429
rect -5307 24092 -4907 24140
rect -4730 24429 -4330 24492
rect -4730 24140 -4671 24429
rect -4397 24140 -4330 24429
rect -4730 24092 -4330 24140
rect -4153 24429 -3753 24492
rect -4153 24140 -4094 24429
rect -3820 24140 -3753 24429
rect -4153 24092 -3753 24140
rect -3576 24429 -3176 24492
rect -3576 24140 -3517 24429
rect -3243 24140 -3176 24429
rect -3576 24092 -3176 24140
rect -2999 24429 -2599 24492
rect -2999 24140 -2940 24429
rect -2666 24140 -2599 24429
rect -2999 24092 -2599 24140
rect -2422 24429 -2022 24492
rect -2422 24140 -2363 24429
rect -2089 24140 -2022 24429
rect -2422 24092 -2022 24140
rect -1845 24429 -1445 24492
rect -1845 24140 -1786 24429
rect -1512 24140 -1445 24429
rect -1845 24092 -1445 24140
rect -1268 24429 -868 24492
rect -1268 24140 -1209 24429
rect -935 24140 -868 24429
rect -1268 24092 -868 24140
rect -691 24429 -291 24492
rect -691 24140 -632 24429
rect -358 24140 -291 24429
rect -691 24092 -291 24140
rect -114 24429 286 24492
rect -114 24140 -55 24429
rect 219 24140 286 24429
rect -114 24092 286 24140
rect 463 24429 863 24492
rect 463 24140 522 24429
rect 796 24140 863 24429
rect 463 24092 863 24140
rect 1040 24429 1440 24492
rect 1040 24140 1099 24429
rect 1373 24140 1440 24429
rect 1040 24092 1440 24140
rect 1617 24429 2017 24492
rect 1617 24140 1676 24429
rect 1950 24140 2017 24429
rect 1617 24092 2017 24140
rect 2194 24429 2594 24492
rect 2194 24140 2253 24429
rect 2527 24140 2594 24429
rect 2194 24092 2594 24140
rect 2771 24429 3171 24492
rect 2771 24140 2830 24429
rect 3104 24140 3171 24429
rect 2771 24092 3171 24140
rect 3348 24429 3748 24492
rect 3348 24140 3407 24429
rect 3681 24140 3748 24429
rect 3348 24092 3748 24140
rect 3925 24429 4325 24492
rect 3925 24140 3984 24429
rect 4258 24140 4325 24429
rect 3925 24092 4325 24140
rect 4502 24429 4902 24492
rect 4502 24140 4561 24429
rect 4835 24140 4902 24429
rect 4502 24092 4902 24140
rect 5079 24429 5479 24492
rect 5079 24140 5138 24429
rect 5412 24140 5479 24429
rect 5079 24092 5479 24140
rect 5656 24429 6056 24492
rect 5656 24140 5715 24429
rect 5989 24140 6056 24429
rect 5656 24092 6056 24140
rect 6233 24429 6633 24492
rect 6233 24140 6292 24429
rect 6566 24140 6633 24429
rect 6233 24092 6633 24140
rect 6810 24429 7210 24492
rect 6810 24140 6869 24429
rect 7143 24140 7210 24429
rect 6810 24092 7210 24140
rect 7387 24429 7787 24492
rect 7387 24140 7446 24429
rect 7720 24140 7787 24429
rect 7387 24092 7787 24140
rect 7964 24429 8364 24492
rect 7964 24140 8023 24429
rect 8297 24140 8364 24429
rect 7964 24092 8364 24140
rect 8541 24429 8941 24492
rect 8541 24140 8600 24429
rect 8874 24140 8941 24429
rect 8541 24092 8941 24140
rect 9118 24429 9518 24492
rect 9118 24140 9177 24429
rect 9451 24140 9518 24429
rect 9118 24092 9518 24140
rect 9695 24429 10095 24492
rect 9695 24140 9754 24429
rect 10028 24140 10095 24429
rect 9695 24092 10095 24140
rect 10272 24429 10672 24492
rect 10272 24140 10331 24429
rect 10605 24140 10672 24429
rect 10272 24092 10672 24140
rect 10849 24429 11249 24492
rect 10849 24140 10908 24429
rect 11182 24140 11249 24429
rect 10849 24092 11249 24140
rect 11426 24429 11826 24492
rect 11426 24140 11485 24429
rect 11759 24140 11826 24429
rect 11426 24092 11826 24140
rect 12003 24429 12403 24492
rect 12003 24140 12062 24429
rect 12336 24140 12403 24429
rect 12003 24092 12403 24140
rect 12580 24429 12980 24492
rect 12580 24140 12639 24429
rect 12913 24140 12980 24429
rect 12580 24092 12980 24140
rect 13157 24429 13557 24492
rect 13157 24140 13216 24429
rect 13490 24140 13557 24429
rect 13157 24092 13557 24140
rect 13734 24429 14134 24492
rect 13734 24140 13793 24429
rect 14067 24140 14134 24429
rect 13734 24092 14134 24140
rect 14311 24429 14711 24492
rect 14311 24140 14370 24429
rect 14644 24140 14711 24429
rect 14311 24092 14711 24140
rect 14888 24429 15288 24492
rect 14888 24140 14947 24429
rect 15221 24140 15288 24429
rect 14888 24092 15288 24140
rect 15465 24429 15865 24492
rect 15465 24140 15524 24429
rect 15798 24140 15865 24429
rect 15465 24092 15865 24140
rect 16042 24429 16442 24492
rect 16042 24140 16101 24429
rect 16375 24140 16442 24429
rect 16042 24092 16442 24140
rect 16619 24429 17019 24492
rect 16619 24140 16678 24429
rect 16952 24140 17019 24429
rect 16619 24092 17019 24140
rect 17196 24429 17596 24492
rect 17196 24140 17255 24429
rect 17529 24140 17596 24429
rect 17196 24092 17596 24140
rect 17773 24429 18173 24492
rect 17773 24140 17832 24429
rect 18106 24140 18173 24429
rect 17773 24092 18173 24140
rect 18350 24429 18750 24492
rect 18350 24140 18409 24429
rect 18683 24140 18750 24429
rect 18350 24092 18750 24140
rect 18927 24429 19327 24492
rect 18927 24140 18986 24429
rect 19260 24140 19327 24429
rect 18927 24092 19327 24140
rect 19504 24429 19904 24492
rect 19504 24140 19563 24429
rect 19837 24140 19904 24429
rect 19504 24092 19904 24140
rect 20081 24429 20481 24492
rect 20081 24140 20140 24429
rect 20414 24140 20481 24429
rect 20081 24092 20481 24140
rect 20658 24429 21058 24492
rect 20658 24140 20717 24429
rect 20991 24140 21058 24429
rect 20658 24092 21058 24140
rect 21235 24429 21635 24492
rect 21235 24140 21294 24429
rect 21568 24140 21635 24429
rect 21235 24092 21635 24140
rect 21812 24429 22212 24492
rect 21812 24140 21871 24429
rect 22145 24140 22212 24429
rect 21812 24092 22212 24140
rect 22389 24429 22789 24492
rect 22389 24140 22448 24429
rect 22722 24140 22789 24429
rect 22389 24092 22789 24140
rect 22966 24429 23366 24492
rect 22966 24140 23025 24429
rect 23299 24140 23366 24429
rect 22966 24092 23366 24140
rect 23543 24429 23943 24492
rect 23543 24140 23602 24429
rect 23876 24140 23943 24429
rect 23543 24092 23943 24140
rect 24120 24429 24520 24492
rect 24120 24140 24179 24429
rect 24453 24140 24520 24429
rect 24120 24092 24520 24140
rect 24697 24429 25097 24492
rect 24697 24140 24756 24429
rect 25030 24140 25097 24429
rect 24697 24092 25097 24140
rect 25274 24429 25674 24492
rect 25274 24140 25333 24429
rect 25607 24140 25674 24429
rect 25274 24092 25674 24140
rect 25851 24429 26251 24492
rect 25851 24140 25910 24429
rect 26184 24140 26251 24429
rect 25851 24092 26251 24140
rect 26428 24429 26828 24492
rect 26428 24140 26487 24429
rect 26761 24140 26828 24429
rect 26428 24092 26828 24140
rect 27005 24429 27405 24492
rect 27005 24140 27064 24429
rect 27338 24140 27405 24429
rect 27005 24092 27405 24140
rect 27582 24429 27982 24492
rect 27582 24140 27641 24429
rect 27915 24140 27982 24429
rect 27582 24092 27982 24140
rect 28159 24429 28559 24492
rect 28159 24140 28218 24429
rect 28492 24140 28559 24429
rect 28159 24092 28559 24140
rect 28736 24429 29136 24492
rect 28736 24140 28795 24429
rect 29069 24140 29136 24429
rect 28736 24092 29136 24140
rect 29313 24429 29713 24492
rect 29313 24140 29372 24429
rect 29646 24140 29713 24429
rect 29313 24092 29713 24140
rect 29890 24429 30290 24492
rect 29890 24140 29949 24429
rect 30223 24140 30290 24429
rect 29890 24092 30290 24140
rect 30467 24429 30867 24492
rect 30467 24140 30526 24429
rect 30800 24140 30867 24429
rect 30467 24092 30867 24140
rect 31044 24429 31444 24492
rect 31044 24140 31103 24429
rect 31377 24140 31444 24429
rect 31044 24092 31444 24140
rect 31621 24429 32021 24492
rect 31621 24140 31680 24429
rect 31954 24140 32021 24429
rect 31621 24092 32021 24140
rect 32198 24429 32598 24492
rect 32198 24140 32257 24429
rect 32531 24140 32598 24429
rect 32198 24092 32598 24140
rect 32775 24429 33175 24492
rect 32775 24140 32834 24429
rect 33108 24140 33175 24429
rect 32775 24092 33175 24140
rect 33352 24429 33752 24492
rect 33352 24140 33411 24429
rect 33685 24140 33752 24429
rect 33352 24092 33752 24140
rect 33929 24429 34329 24492
rect 33929 24140 33988 24429
rect 34262 24140 34329 24429
rect 33929 24092 34329 24140
rect 34506 24429 34906 24492
rect 34506 24140 34565 24429
rect 34839 24140 34906 24429
rect 34506 24092 34906 24140
rect 35083 24429 35483 24492
rect 35083 24140 35142 24429
rect 35416 24140 35483 24429
rect 35083 24092 35483 24140
rect 35660 24429 36060 24492
rect 35660 24140 35719 24429
rect 35993 24140 36060 24429
rect 35660 24092 36060 24140
rect 36237 24429 36637 24492
rect 36237 24140 36296 24429
rect 36570 24140 36637 24429
rect 36237 24092 36637 24140
rect 36814 24429 37214 24492
rect 36814 24140 36873 24429
rect 37147 24140 37214 24429
rect 36814 24092 37214 24140
rect 37391 24429 37791 24492
rect 37391 24140 37450 24429
rect 37724 24140 37791 24429
rect 37391 24092 37791 24140
rect 37968 24429 38368 24492
rect 37968 24140 38027 24429
rect 38301 24140 38368 24429
rect 37968 24092 38368 24140
rect 38545 24429 38945 24492
rect 38545 24140 38604 24429
rect 38878 24140 38945 24429
rect 38545 24092 38945 24140
rect 39122 24429 39522 24492
rect 39122 24140 39181 24429
rect 39455 24140 39522 24429
rect 39122 24092 39522 24140
rect 39699 24429 40099 24492
rect 39699 24140 39758 24429
rect 40032 24140 40099 24429
rect 39699 24092 40099 24140
rect 40276 24429 40676 24492
rect 40276 24140 40335 24429
rect 40609 24140 40676 24429
rect 40276 24092 40676 24140
rect 40853 24429 41253 24492
rect 40853 24140 40912 24429
rect 41186 24140 41253 24429
rect 40853 24092 41253 24140
rect 41430 24429 41830 24492
rect 41430 24140 41489 24429
rect 41763 24140 41830 24429
rect 41430 24092 41830 24140
rect 42007 24429 42407 24492
rect 42007 24140 42066 24429
rect 42340 24140 42407 24429
rect 42007 24092 42407 24140
rect 42584 24429 42984 24492
rect 42584 24140 42643 24429
rect 42917 24140 42984 24429
rect 42584 24092 42984 24140
rect 43161 24429 43561 24492
rect 43161 24140 43220 24429
rect 43494 24140 43561 24429
rect 43161 24092 43561 24140
rect 43738 24429 44138 24492
rect 43738 24140 43797 24429
rect 44071 24140 44138 24429
rect 43738 24092 44138 24140
rect 44315 24429 44715 24492
rect 44315 24140 44374 24429
rect 44648 24140 44715 24429
rect 44315 24092 44715 24140
rect 44892 24429 45292 24492
rect 44892 24140 44951 24429
rect 45225 24140 45292 24429
rect 44892 24092 45292 24140
rect 45469 24429 45869 24492
rect 45469 24140 45528 24429
rect 45802 24140 45869 24429
rect 45469 24092 45869 24140
rect 46046 24429 46446 24492
rect 46046 24140 46105 24429
rect 46379 24140 46446 24429
rect 46046 24092 46446 24140
rect 46623 24429 47023 24492
rect 46623 24140 46682 24429
rect 46956 24140 47023 24429
rect 46623 24092 47023 24140
rect 47200 24429 47600 24492
rect 47200 24140 47259 24429
rect 47533 24140 47600 24429
rect 47200 24092 47600 24140
rect 47777 24429 48177 24492
rect 47777 24140 47836 24429
rect 48110 24140 48177 24429
rect 47777 24092 48177 24140
rect 48354 24429 48754 24492
rect 48354 24140 48413 24429
rect 48687 24140 48754 24429
rect 48354 24092 48754 24140
rect 48931 24429 49331 24492
rect 48931 24140 48990 24429
rect 49264 24140 49331 24429
rect 48931 24092 49331 24140
rect 49508 24429 49908 24492
rect 49508 24140 49567 24429
rect 49841 24140 49908 24429
rect 49508 24092 49908 24140
rect 50085 24429 50485 24492
rect 50085 24140 50144 24429
rect 50418 24140 50485 24429
rect 50662 24429 51062 24492
rect 50662 24163 50721 24429
rect 50085 24093 50485 24140
rect 50663 24140 50721 24163
rect 50995 24140 51062 24429
rect 50085 24092 50432 24093
rect 50663 24092 51062 24140
rect 51239 24429 51639 24492
rect 51239 24140 51298 24429
rect 51572 24140 51639 24429
rect 51239 24092 51639 24140
rect 51816 24429 52216 24492
rect 51816 24140 51875 24429
rect 52149 24140 52216 24429
rect 51816 24092 52216 24140
rect 52393 24429 52793 24492
rect 52393 24140 52452 24429
rect 52726 24140 52793 24429
rect 52393 24092 52793 24140
rect 52970 24429 53370 24492
rect 52970 24140 53029 24429
rect 53303 24140 53370 24429
rect 52970 24092 53370 24140
rect 53547 24429 53947 24492
rect 53547 24140 53606 24429
rect 53880 24140 53947 24429
rect 53547 24092 53947 24140
rect 54124 24429 54524 24492
rect 54124 24140 54183 24429
rect 54457 24140 54524 24429
rect 54124 24092 54524 24140
rect 54701 24429 55101 24492
rect 54701 24140 54760 24429
rect 55034 24140 55101 24429
rect 54701 24092 55101 24140
rect 55278 24429 55678 24492
rect 55278 24140 55337 24429
rect 55611 24140 55678 24429
rect 55278 24092 55678 24140
rect 55855 24429 56255 24492
rect 55855 24140 55914 24429
rect 56188 24140 56255 24429
rect 55855 24092 56255 24140
rect 42549 9113 42618 9393
rect -2635 -8286 1484 -8234
rect 833 -9773 3727 -9690
rect 8336 -21029 8590 -21020
rect 5973 -21454 6890 -21380
rect -2764 -22117 -2751 -22079
rect -2764 -22148 -2516 -22117
rect -2849 -22263 -2310 -22148
rect -2849 -22264 -2280 -22263
rect -2849 -22335 -1927 -22264
rect -2849 -22425 -2310 -22335
rect -1932 -22425 -1927 -22335
rect 11456 -22354 11610 -22347
rect 11453 -22373 11610 -22354
rect 11457 -22386 11610 -22373
rect 11439 -22393 11610 -22386
rect 11439 -22405 11606 -22393
rect 11457 -22430 11601 -22405
<< psubdiffcont >>
rect -55497 -29952 -55172 -29624
rect -55002 -29952 -54677 -29624
rect -54507 -29952 -54182 -29624
rect -54012 -29952 -53687 -29624
rect -53517 -29952 -53192 -29624
rect -53022 -29952 -52697 -29624
rect -52527 -29952 -52202 -29624
rect -52032 -29952 -51707 -29624
rect -51537 -29952 -51212 -29624
rect -51042 -29952 -50717 -29624
rect -50547 -29952 -50222 -29624
rect -50052 -29952 -49727 -29624
rect -49557 -29952 -49232 -29624
rect -49062 -29952 -48737 -29624
rect -48567 -29952 -48242 -29624
rect -48072 -29952 -47747 -29624
rect -47577 -29952 -47252 -29624
rect -47082 -29952 -46757 -29624
rect -46587 -29952 -46262 -29624
rect -46092 -29952 -45767 -29624
rect -45597 -29952 -45272 -29624
rect -45102 -29952 -44777 -29624
rect -44607 -29952 -44282 -29624
rect -44112 -29952 -43787 -29624
rect -43617 -29952 -43292 -29624
rect -43122 -29952 -42797 -29624
rect -42627 -29952 -42302 -29624
rect -42132 -29952 -41807 -29624
rect -41637 -29952 -41312 -29624
rect -41142 -29952 -40817 -29624
rect -40647 -29952 -40322 -29624
rect -40152 -29952 -39827 -29624
rect -39657 -29952 -39332 -29624
rect -39162 -29952 -38837 -29624
rect -38667 -29952 -38342 -29624
rect -38172 -29952 -37847 -29624
rect -37677 -29952 -37352 -29624
rect -37182 -29952 -36857 -29624
rect -36687 -29952 -36362 -29624
rect -36192 -29952 -35867 -29624
rect -35697 -29952 -35372 -29624
rect -35202 -29952 -34877 -29624
rect -34707 -29952 -34382 -29624
rect -34212 -29952 -33887 -29624
rect -33717 -29952 -33392 -29624
rect -33222 -29952 -32897 -29624
rect -32727 -29952 -32402 -29624
rect -32232 -29952 -31907 -29624
rect -31737 -29952 -31412 -29624
rect -31242 -29952 -30917 -29624
rect -30747 -29952 -30422 -29624
rect -30252 -29952 -29927 -29624
rect -29757 -29952 -29432 -29624
rect -29262 -29952 -28937 -29624
rect -28767 -29952 -28442 -29624
rect -28272 -29952 -27947 -29624
rect -27777 -29952 -27452 -29624
rect -27282 -29952 -26957 -29624
rect -26787 -29952 -26462 -29624
rect -26292 -29952 -25967 -29624
rect -25797 -29952 -25472 -29624
rect -25302 -29952 -24977 -29624
rect -24807 -29952 -24482 -29624
rect -24312 -29952 -23987 -29624
rect -23817 -29952 -23492 -29624
rect -23322 -29952 -22997 -29624
rect -22827 -29952 -22502 -29624
rect -22332 -29952 -22007 -29624
rect -21837 -29952 -21512 -29624
rect -21342 -29952 -21017 -29624
rect -20847 -29952 -20522 -29624
rect -20352 -29952 -20027 -29624
rect -19857 -29952 -19532 -29624
rect -19362 -29952 -19037 -29624
rect -18867 -29952 -18542 -29624
rect -18372 -29952 -18047 -29624
rect -17877 -29952 -17552 -29624
rect -17382 -29952 -17057 -29624
rect -16887 -29952 -16562 -29624
rect -16392 -29952 -16067 -29624
rect -15897 -29952 -15572 -29624
rect -15402 -29952 -15077 -29624
rect -14907 -29952 -14582 -29624
rect -14412 -29952 -14087 -29624
rect -13917 -29952 -13592 -29624
rect -13422 -29952 -13097 -29624
rect -12927 -29952 -12602 -29624
rect -12432 -29952 -12107 -29624
rect -11937 -29952 -11612 -29624
rect -11442 -29952 -11117 -29624
rect -10947 -29952 -10622 -29624
rect -10452 -29952 -10127 -29624
rect -9957 -29952 -9632 -29624
rect -9462 -29952 -9137 -29624
rect -8967 -29952 -8642 -29624
rect -8472 -29952 -8147 -29624
rect -7977 -29952 -7652 -29624
rect -7482 -29952 -7157 -29624
rect -6987 -29952 -6662 -29624
rect -6492 -29952 -6167 -29624
rect -5997 -29952 -5672 -29624
rect -5502 -29952 -5177 -29624
rect -5007 -29952 -4682 -29624
rect -4512 -29952 -4187 -29624
rect -4017 -29952 -3692 -29624
rect -3522 -29952 -3197 -29624
rect -3027 -29952 -2702 -29624
rect -2532 -29952 -2207 -29624
rect -2037 -29952 -1712 -29624
rect -1542 -29952 -1217 -29624
rect -1047 -29952 -722 -29624
rect -552 -29952 -227 -29624
rect -57 -29952 268 -29624
rect 438 -29952 763 -29624
rect 933 -29952 1258 -29624
rect 1428 -29952 1753 -29624
rect 1923 -29952 2248 -29624
rect 2418 -29952 2743 -29624
rect 2913 -29952 3238 -29624
rect 3408 -29952 3733 -29624
rect 3903 -29952 4228 -29624
rect 4398 -29952 4723 -29624
rect 4893 -29952 5218 -29624
rect 5388 -29952 5713 -29624
rect 5883 -29952 6208 -29624
rect 6378 -29952 6703 -29624
rect 6873 -29952 7198 -29624
rect 7368 -29952 7693 -29624
rect 7863 -29952 8188 -29624
rect 8358 -29952 8683 -29624
rect 8853 -29952 9178 -29624
rect 9348 -29952 9673 -29624
rect 9843 -29952 10168 -29624
rect 10338 -29952 10663 -29624
rect 10833 -29952 11158 -29624
rect 11328 -29952 11653 -29624
rect 11823 -29952 12148 -29624
rect 12318 -29952 12643 -29624
rect 12813 -29952 13138 -29624
rect 13308 -29952 13633 -29624
rect 13803 -29952 14128 -29624
rect 14298 -29952 14623 -29624
rect 14793 -29952 15118 -29624
rect 15288 -29952 15613 -29624
rect 15783 -29952 16108 -29624
rect 16278 -29952 16603 -29624
rect 16773 -29952 17098 -29624
rect 17268 -29952 17593 -29624
rect 17763 -29952 18088 -29624
rect 18258 -29952 18583 -29624
rect 18753 -29952 19078 -29624
rect 19248 -29952 19573 -29624
rect 19743 -29952 20068 -29624
rect 20238 -29952 20563 -29624
rect 20733 -29952 21058 -29624
rect 21228 -29952 21553 -29624
rect 21723 -29952 22048 -29624
rect 22218 -29952 22543 -29624
rect 22713 -29952 23038 -29624
rect 23208 -29952 23533 -29624
rect 23703 -29952 24028 -29624
rect 24198 -29952 24523 -29624
rect 24693 -29952 25018 -29624
rect 25188 -29952 25513 -29624
rect 25683 -29952 26008 -29624
rect 26178 -29952 26503 -29624
rect 26673 -29952 26998 -29624
rect 27168 -29952 27493 -29624
rect 27663 -29952 27988 -29624
rect 28158 -29952 28483 -29624
rect 28653 -29952 28978 -29624
rect 29148 -29952 29473 -29624
rect 29643 -29952 29968 -29624
rect 30138 -29952 30463 -29624
rect 30633 -29952 30958 -29624
rect 31128 -29952 31453 -29624
rect 31623 -29952 31948 -29624
rect 32118 -29952 32443 -29624
rect 32613 -29952 32938 -29624
rect 33108 -29952 33433 -29624
rect 33603 -29952 33928 -29624
rect 34098 -29952 34423 -29624
rect 34593 -29952 34918 -29624
rect 35088 -29952 35413 -29624
rect 35583 -29952 35908 -29624
rect 36078 -29952 36403 -29624
rect 36573 -29952 36898 -29624
rect 37068 -29952 37393 -29624
rect 37563 -29952 37888 -29624
rect 38058 -29952 38383 -29624
rect 38553 -29952 38878 -29624
rect 39048 -29952 39373 -29624
rect 39543 -29952 39868 -29624
rect 40038 -29952 40363 -29624
rect 40533 -29952 40858 -29624
rect 41028 -29952 41353 -29624
rect 41523 -29952 41848 -29624
rect 42018 -29952 42343 -29624
rect 42513 -29952 42838 -29624
rect 43008 -29952 43333 -29624
rect 43503 -29952 43828 -29624
rect 43998 -29952 44323 -29624
rect 44493 -29952 44818 -29624
rect 44988 -29952 45313 -29624
rect 45483 -29952 45808 -29624
rect 45978 -29952 46303 -29624
rect 46473 -29952 46798 -29624
rect 46968 -29952 47293 -29624
rect 47463 -29952 47788 -29624
rect 47958 -29952 48283 -29624
rect 48453 -29952 48778 -29624
rect 48948 -29952 49273 -29624
rect 49443 -29952 49768 -29624
rect 49938 -29952 50263 -29624
rect 50433 -29952 50758 -29624
rect 50928 -29952 51253 -29624
rect 51423 -29952 51748 -29624
rect 51918 -29952 52243 -29624
rect 52413 -29952 52738 -29624
rect 52908 -29952 53233 -29624
rect 53403 -29952 53728 -29624
rect 53898 -29952 54223 -29624
rect -55497 -30428 -55172 -30100
rect -55002 -30428 -54677 -30100
rect -54507 -30428 -54182 -30100
rect -54012 -30428 -53687 -30100
rect -53517 -30428 -53192 -30100
rect -53022 -30428 -52697 -30100
rect -52527 -30428 -52202 -30100
rect -52032 -30428 -51707 -30100
rect -51537 -30428 -51212 -30100
rect -51042 -30428 -50717 -30100
rect -50547 -30428 -50222 -30100
rect -50052 -30428 -49727 -30100
rect -49557 -30428 -49232 -30100
rect -49062 -30428 -48737 -30100
rect -48567 -30428 -48242 -30100
rect -48072 -30428 -47747 -30100
rect -47577 -30428 -47252 -30100
rect -47082 -30428 -46757 -30100
rect -46587 -30428 -46262 -30100
rect -46092 -30428 -45767 -30100
rect -45597 -30428 -45272 -30100
rect -45102 -30428 -44777 -30100
rect -44607 -30428 -44282 -30100
rect -44112 -30428 -43787 -30100
rect -43617 -30428 -43292 -30100
rect -43122 -30428 -42797 -30100
rect -42627 -30428 -42302 -30100
rect -42132 -30428 -41807 -30100
rect -41637 -30428 -41312 -30100
rect -41142 -30428 -40817 -30100
rect -40647 -30428 -40322 -30100
rect -40152 -30428 -39827 -30100
rect -39657 -30428 -39332 -30100
rect -39162 -30428 -38837 -30100
rect -38667 -30428 -38342 -30100
rect -38172 -30428 -37847 -30100
rect -37677 -30428 -37352 -30100
rect -37182 -30428 -36857 -30100
rect -36687 -30428 -36362 -30100
rect -36192 -30428 -35867 -30100
rect -35697 -30428 -35372 -30100
rect -35202 -30428 -34877 -30100
rect -34707 -30428 -34382 -30100
rect -34212 -30428 -33887 -30100
rect -33717 -30428 -33392 -30100
rect -33222 -30428 -32897 -30100
rect -32727 -30428 -32402 -30100
rect -32232 -30428 -31907 -30100
rect -31737 -30428 -31412 -30100
rect -31242 -30428 -30917 -30100
rect -30747 -30428 -30422 -30100
rect -30252 -30428 -29927 -30100
rect -29757 -30428 -29432 -30100
rect -29262 -30428 -28937 -30100
rect -28767 -30428 -28442 -30100
rect -28272 -30428 -27947 -30100
rect -27777 -30428 -27452 -30100
rect -27282 -30428 -26957 -30100
rect -26787 -30428 -26462 -30100
rect -26292 -30428 -25967 -30100
rect -25797 -30428 -25472 -30100
rect -25302 -30428 -24977 -30100
rect -24807 -30428 -24482 -30100
rect -24312 -30428 -23987 -30100
rect -23817 -30428 -23492 -30100
rect -23322 -30428 -22997 -30100
rect -22827 -30428 -22502 -30100
rect -22332 -30428 -22007 -30100
rect -21837 -30428 -21512 -30100
rect -21342 -30428 -21017 -30100
rect -20847 -30428 -20522 -30100
rect -20352 -30428 -20027 -30100
rect -19857 -30428 -19532 -30100
rect -19362 -30428 -19037 -30100
rect -18867 -30428 -18542 -30100
rect -18372 -30428 -18047 -30100
rect -17877 -30428 -17552 -30100
rect -17382 -30428 -17057 -30100
rect -16887 -30428 -16562 -30100
rect -16392 -30428 -16067 -30100
rect -15897 -30428 -15572 -30100
rect -15402 -30428 -15077 -30100
rect -14907 -30428 -14582 -30100
rect -14412 -30428 -14087 -30100
rect -13917 -30428 -13592 -30100
rect -13422 -30428 -13097 -30100
rect -12927 -30428 -12602 -30100
rect -12432 -30428 -12107 -30100
rect -11937 -30428 -11612 -30100
rect -11442 -30428 -11117 -30100
rect -10947 -30428 -10622 -30100
rect -10452 -30428 -10127 -30100
rect -9957 -30428 -9632 -30100
rect -9462 -30428 -9137 -30100
rect -8967 -30428 -8642 -30100
rect -8472 -30428 -8147 -30100
rect -7977 -30428 -7652 -30100
rect -7482 -30428 -7157 -30100
rect -6987 -30428 -6662 -30100
rect -6492 -30428 -6167 -30100
rect -5997 -30428 -5672 -30100
rect -5502 -30428 -5177 -30100
rect -5007 -30428 -4682 -30100
rect -4512 -30428 -4187 -30100
rect -4017 -30428 -3692 -30100
rect -3522 -30428 -3197 -30100
rect -3027 -30428 -2702 -30100
rect -2532 -30428 -2207 -30100
rect -2037 -30428 -1712 -30100
rect -1542 -30428 -1217 -30100
rect -1047 -30428 -722 -30100
rect -552 -30428 -227 -30100
rect -57 -30428 268 -30100
rect 438 -30428 763 -30100
rect 933 -30428 1258 -30100
rect 1428 -30428 1753 -30100
rect 1923 -30428 2248 -30100
rect 2418 -30428 2743 -30100
rect 2913 -30428 3238 -30100
rect 3408 -30428 3733 -30100
rect 3903 -30428 4228 -30100
rect 4398 -30428 4723 -30100
rect 4893 -30428 5218 -30100
rect 5388 -30428 5713 -30100
rect 5883 -30428 6208 -30100
rect 6378 -30428 6703 -30100
rect 6873 -30428 7198 -30100
rect 7368 -30428 7693 -30100
rect 7863 -30428 8188 -30100
rect 8358 -30428 8683 -30100
rect 8853 -30428 9178 -30100
rect 9348 -30428 9673 -30100
rect 9843 -30428 10168 -30100
rect 10338 -30428 10663 -30100
rect 10833 -30428 11158 -30100
rect 11328 -30428 11653 -30100
rect 11823 -30428 12148 -30100
rect 12318 -30428 12643 -30100
rect 12813 -30428 13138 -30100
rect 13308 -30428 13633 -30100
rect 13803 -30428 14128 -30100
rect 14298 -30428 14623 -30100
rect 14793 -30428 15118 -30100
rect 15288 -30428 15613 -30100
rect 15783 -30428 16108 -30100
rect 16278 -30428 16603 -30100
rect 16773 -30428 17098 -30100
rect 17268 -30428 17593 -30100
rect 17763 -30428 18088 -30100
rect 18258 -30428 18583 -30100
rect 18753 -30428 19078 -30100
rect 19248 -30428 19573 -30100
rect 19743 -30428 20068 -30100
rect 20238 -30428 20563 -30100
rect 20733 -30428 21058 -30100
rect 21228 -30428 21553 -30100
rect 21723 -30428 22048 -30100
rect 22218 -30428 22543 -30100
rect 22713 -30428 23038 -30100
rect 23208 -30428 23533 -30100
rect 23703 -30428 24028 -30100
rect 24198 -30428 24523 -30100
rect 24693 -30428 25018 -30100
rect 25188 -30428 25513 -30100
rect 25683 -30428 26008 -30100
rect 26178 -30428 26503 -30100
rect 26673 -30428 26998 -30100
rect 27168 -30428 27493 -30100
rect 27663 -30428 27988 -30100
rect 28158 -30428 28483 -30100
rect 28653 -30428 28978 -30100
rect 29148 -30428 29473 -30100
rect 29643 -30428 29968 -30100
rect 30138 -30428 30463 -30100
rect 30633 -30428 30958 -30100
rect 31128 -30428 31453 -30100
rect 31623 -30428 31948 -30100
rect 32118 -30428 32443 -30100
rect 32613 -30428 32938 -30100
rect 33108 -30428 33433 -30100
rect 33603 -30428 33928 -30100
rect 34098 -30428 34423 -30100
rect 34593 -30428 34918 -30100
rect 35088 -30428 35413 -30100
rect 35583 -30428 35908 -30100
rect 36078 -30428 36403 -30100
rect 36573 -30428 36898 -30100
rect 37068 -30428 37393 -30100
rect 37563 -30428 37888 -30100
rect 38058 -30428 38383 -30100
rect 38553 -30428 38878 -30100
rect 39048 -30428 39373 -30100
rect 39543 -30428 39868 -30100
rect 40038 -30428 40363 -30100
rect 40533 -30428 40858 -30100
rect 41028 -30428 41353 -30100
rect 41523 -30428 41848 -30100
rect 42018 -30428 42343 -30100
rect 42513 -30428 42838 -30100
rect 43008 -30428 43333 -30100
rect 43503 -30428 43828 -30100
rect 43998 -30428 44323 -30100
rect 44493 -30428 44818 -30100
rect 44988 -30428 45313 -30100
rect 45483 -30428 45808 -30100
rect 45978 -30428 46303 -30100
rect 46473 -30428 46798 -30100
rect 46968 -30428 47293 -30100
rect 47463 -30428 47788 -30100
rect 47958 -30428 48283 -30100
rect 48453 -30428 48778 -30100
rect 48948 -30428 49273 -30100
rect 49443 -30428 49768 -30100
rect 49938 -30428 50263 -30100
rect 50433 -30428 50758 -30100
rect 50928 -30428 51253 -30100
rect 51423 -30428 51748 -30100
rect 51918 -30428 52243 -30100
rect 52413 -30428 52738 -30100
rect 52908 -30428 53233 -30100
rect 53403 -30428 53728 -30100
rect 53898 -30428 54223 -30100
rect -55497 -30904 -55172 -30576
rect -55002 -30904 -54677 -30576
rect -54507 -30904 -54182 -30576
rect -54012 -30904 -53687 -30576
rect -53517 -30904 -53192 -30576
rect -53022 -30904 -52697 -30576
rect -52527 -30904 -52202 -30576
rect -52032 -30904 -51707 -30576
rect -51537 -30904 -51212 -30576
rect -51042 -30904 -50717 -30576
rect -50547 -30904 -50222 -30576
rect -50052 -30904 -49727 -30576
rect -49557 -30904 -49232 -30576
rect -49062 -30904 -48737 -30576
rect -48567 -30904 -48242 -30576
rect -48072 -30904 -47747 -30576
rect -47577 -30904 -47252 -30576
rect -47082 -30904 -46757 -30576
rect -46587 -30904 -46262 -30576
rect -46092 -30904 -45767 -30576
rect -45597 -30904 -45272 -30576
rect -45102 -30904 -44777 -30576
rect -44607 -30904 -44282 -30576
rect -44112 -30904 -43787 -30576
rect -43617 -30904 -43292 -30576
rect -43122 -30904 -42797 -30576
rect -42627 -30904 -42302 -30576
rect -42132 -30904 -41807 -30576
rect -41637 -30904 -41312 -30576
rect -41142 -30904 -40817 -30576
rect -40647 -30904 -40322 -30576
rect -40152 -30904 -39827 -30576
rect -39657 -30904 -39332 -30576
rect -39162 -30904 -38837 -30576
rect -38667 -30904 -38342 -30576
rect -38172 -30904 -37847 -30576
rect -37677 -30904 -37352 -30576
rect -37182 -30904 -36857 -30576
rect -36687 -30904 -36362 -30576
rect -36192 -30904 -35867 -30576
rect -35697 -30904 -35372 -30576
rect -35202 -30904 -34877 -30576
rect -34707 -30904 -34382 -30576
rect -34212 -30904 -33887 -30576
rect -33717 -30904 -33392 -30576
rect -33222 -30904 -32897 -30576
rect -32727 -30904 -32402 -30576
rect -32232 -30904 -31907 -30576
rect -31737 -30904 -31412 -30576
rect -31242 -30904 -30917 -30576
rect -30747 -30904 -30422 -30576
rect -30252 -30904 -29927 -30576
rect -29757 -30904 -29432 -30576
rect -29262 -30904 -28937 -30576
rect -28767 -30904 -28442 -30576
rect -28272 -30904 -27947 -30576
rect -27777 -30904 -27452 -30576
rect -27282 -30904 -26957 -30576
rect -26787 -30904 -26462 -30576
rect -26292 -30904 -25967 -30576
rect -25797 -30904 -25472 -30576
rect -25302 -30904 -24977 -30576
rect -24807 -30904 -24482 -30576
rect -24312 -30904 -23987 -30576
rect -23817 -30904 -23492 -30576
rect -23322 -30904 -22997 -30576
rect -22827 -30904 -22502 -30576
rect -22332 -30904 -22007 -30576
rect -21837 -30904 -21512 -30576
rect -21342 -30904 -21017 -30576
rect -20847 -30904 -20522 -30576
rect -20352 -30904 -20027 -30576
rect -19857 -30904 -19532 -30576
rect -19362 -30904 -19037 -30576
rect -18867 -30904 -18542 -30576
rect -18372 -30904 -18047 -30576
rect -17877 -30904 -17552 -30576
rect -17382 -30904 -17057 -30576
rect -16887 -30904 -16562 -30576
rect -16392 -30904 -16067 -30576
rect -15897 -30904 -15572 -30576
rect -15402 -30904 -15077 -30576
rect -14907 -30904 -14582 -30576
rect -14412 -30904 -14087 -30576
rect -13917 -30904 -13592 -30576
rect -13422 -30904 -13097 -30576
rect -12927 -30904 -12602 -30576
rect -12432 -30904 -12107 -30576
rect -11937 -30904 -11612 -30576
rect -11442 -30904 -11117 -30576
rect -10947 -30904 -10622 -30576
rect -10452 -30904 -10127 -30576
rect -9957 -30904 -9632 -30576
rect -9462 -30904 -9137 -30576
rect -8967 -30904 -8642 -30576
rect -8472 -30904 -8147 -30576
rect -7977 -30904 -7652 -30576
rect -7482 -30904 -7157 -30576
rect -6987 -30904 -6662 -30576
rect -6492 -30904 -6167 -30576
rect -5997 -30904 -5672 -30576
rect -5502 -30904 -5177 -30576
rect -5007 -30904 -4682 -30576
rect -4512 -30904 -4187 -30576
rect -4017 -30904 -3692 -30576
rect -3522 -30904 -3197 -30576
rect -3027 -30904 -2702 -30576
rect -2532 -30904 -2207 -30576
rect -2037 -30904 -1712 -30576
rect -1542 -30904 -1217 -30576
rect -1047 -30904 -722 -30576
rect -552 -30904 -227 -30576
rect -57 -30904 268 -30576
rect 438 -30904 763 -30576
rect 933 -30904 1258 -30576
rect 1428 -30904 1753 -30576
rect 1923 -30904 2248 -30576
rect 2418 -30904 2743 -30576
rect 2913 -30904 3238 -30576
rect 3408 -30904 3733 -30576
rect 3903 -30904 4228 -30576
rect 4398 -30904 4723 -30576
rect 4893 -30904 5218 -30576
rect 5388 -30904 5713 -30576
rect 5883 -30904 6208 -30576
rect 6378 -30904 6703 -30576
rect 6873 -30904 7198 -30576
rect 7368 -30904 7693 -30576
rect 7863 -30904 8188 -30576
rect 8358 -30904 8683 -30576
rect 8853 -30904 9178 -30576
rect 9348 -30904 9673 -30576
rect 9843 -30904 10168 -30576
rect 10338 -30904 10663 -30576
rect 10833 -30904 11158 -30576
rect 11328 -30904 11653 -30576
rect 11823 -30904 12148 -30576
rect 12318 -30904 12643 -30576
rect 12813 -30904 13138 -30576
rect 13308 -30904 13633 -30576
rect 13803 -30904 14128 -30576
rect 14298 -30904 14623 -30576
rect 14793 -30904 15118 -30576
rect 15288 -30904 15613 -30576
rect 15783 -30904 16108 -30576
rect 16278 -30904 16603 -30576
rect 16773 -30904 17098 -30576
rect 17268 -30904 17593 -30576
rect 17763 -30904 18088 -30576
rect 18258 -30904 18583 -30576
rect 18753 -30904 19078 -30576
rect 19248 -30904 19573 -30576
rect 19743 -30904 20068 -30576
rect 20238 -30904 20563 -30576
rect 20733 -30904 21058 -30576
rect 21228 -30904 21553 -30576
rect 21723 -30904 22048 -30576
rect 22218 -30904 22543 -30576
rect 22713 -30904 23038 -30576
rect 23208 -30904 23533 -30576
rect 23703 -30904 24028 -30576
rect 24198 -30904 24523 -30576
rect 24693 -30904 25018 -30576
rect 25188 -30904 25513 -30576
rect 25683 -30904 26008 -30576
rect 26178 -30904 26503 -30576
rect 26673 -30904 26998 -30576
rect 27168 -30904 27493 -30576
rect 27663 -30904 27988 -30576
rect 28158 -30904 28483 -30576
rect 28653 -30904 28978 -30576
rect 29148 -30904 29473 -30576
rect 29643 -30904 29968 -30576
rect 30138 -30904 30463 -30576
rect 30633 -30904 30958 -30576
rect 31128 -30904 31453 -30576
rect 31623 -30904 31948 -30576
rect 32118 -30904 32443 -30576
rect 32613 -30904 32938 -30576
rect 33108 -30904 33433 -30576
rect 33603 -30904 33928 -30576
rect 34098 -30904 34423 -30576
rect 34593 -30904 34918 -30576
rect 35088 -30904 35413 -30576
rect 35583 -30904 35908 -30576
rect 36078 -30904 36403 -30576
rect 36573 -30904 36898 -30576
rect 37068 -30904 37393 -30576
rect 37563 -30904 37888 -30576
rect 38058 -30904 38383 -30576
rect 38553 -30904 38878 -30576
rect 39048 -30904 39373 -30576
rect 39543 -30904 39868 -30576
rect 40038 -30904 40363 -30576
rect 40533 -30904 40858 -30576
rect 41028 -30904 41353 -30576
rect 41523 -30904 41848 -30576
rect 42018 -30904 42343 -30576
rect 42513 -30904 42838 -30576
rect 43008 -30904 43333 -30576
rect 43503 -30904 43828 -30576
rect 43998 -30904 44323 -30576
rect 44493 -30904 44818 -30576
rect 44988 -30904 45313 -30576
rect 45483 -30904 45808 -30576
rect 45978 -30904 46303 -30576
rect 46473 -30904 46798 -30576
rect 46968 -30904 47293 -30576
rect 47463 -30904 47788 -30576
rect 47958 -30904 48283 -30576
rect 48453 -30904 48778 -30576
rect 48948 -30904 49273 -30576
rect 49443 -30904 49768 -30576
rect 49938 -30904 50263 -30576
rect 50433 -30904 50758 -30576
rect 50928 -30904 51253 -30576
rect 51423 -30904 51748 -30576
rect 51918 -30904 52243 -30576
rect 52413 -30904 52738 -30576
rect 52908 -30904 53233 -30576
rect 53403 -30904 53728 -30576
rect 53898 -30904 54223 -30576
rect -55497 -31380 -55172 -31052
rect -55002 -31380 -54677 -31052
rect -54507 -31380 -54182 -31052
rect -54012 -31380 -53687 -31052
rect -53517 -31380 -53192 -31052
rect -53022 -31380 -52697 -31052
rect -52527 -31380 -52202 -31052
rect -52032 -31380 -51707 -31052
rect -51537 -31380 -51212 -31052
rect -51042 -31380 -50717 -31052
rect -50547 -31380 -50222 -31052
rect -50052 -31380 -49727 -31052
rect -49557 -31380 -49232 -31052
rect -49062 -31380 -48737 -31052
rect -48567 -31380 -48242 -31052
rect -48072 -31380 -47747 -31052
rect -47577 -31380 -47252 -31052
rect -47082 -31380 -46757 -31052
rect -46587 -31380 -46262 -31052
rect -46092 -31380 -45767 -31052
rect -45597 -31380 -45272 -31052
rect -45102 -31380 -44777 -31052
rect -44607 -31380 -44282 -31052
rect -44112 -31380 -43787 -31052
rect -43617 -31380 -43292 -31052
rect -43122 -31380 -42797 -31052
rect -42627 -31380 -42302 -31052
rect -42132 -31380 -41807 -31052
rect -41637 -31380 -41312 -31052
rect -41142 -31380 -40817 -31052
rect -40647 -31380 -40322 -31052
rect -40152 -31380 -39827 -31052
rect -39657 -31380 -39332 -31052
rect -39162 -31380 -38837 -31052
rect -38667 -31380 -38342 -31052
rect -38172 -31380 -37847 -31052
rect -37677 -31380 -37352 -31052
rect -37182 -31380 -36857 -31052
rect -36687 -31380 -36362 -31052
rect -36192 -31380 -35867 -31052
rect -35697 -31380 -35372 -31052
rect -35202 -31380 -34877 -31052
rect -34707 -31380 -34382 -31052
rect -34212 -31380 -33887 -31052
rect -33717 -31380 -33392 -31052
rect -33222 -31380 -32897 -31052
rect -32727 -31380 -32402 -31052
rect -32232 -31380 -31907 -31052
rect -31737 -31380 -31412 -31052
rect -31242 -31380 -30917 -31052
rect -30747 -31380 -30422 -31052
rect -30252 -31380 -29927 -31052
rect -29757 -31380 -29432 -31052
rect -29262 -31380 -28937 -31052
rect -28767 -31380 -28442 -31052
rect -28272 -31380 -27947 -31052
rect -27777 -31380 -27452 -31052
rect -27282 -31380 -26957 -31052
rect -26787 -31380 -26462 -31052
rect -26292 -31380 -25967 -31052
rect -25797 -31380 -25472 -31052
rect -25302 -31380 -24977 -31052
rect -24807 -31380 -24482 -31052
rect -24312 -31380 -23987 -31052
rect -23817 -31380 -23492 -31052
rect -23322 -31380 -22997 -31052
rect -22827 -31380 -22502 -31052
rect -22332 -31380 -22007 -31052
rect -21837 -31380 -21512 -31052
rect -21342 -31380 -21017 -31052
rect -20847 -31380 -20522 -31052
rect -20352 -31380 -20027 -31052
rect -19857 -31380 -19532 -31052
rect -19362 -31380 -19037 -31052
rect -18867 -31380 -18542 -31052
rect -18372 -31380 -18047 -31052
rect -17877 -31380 -17552 -31052
rect -17382 -31380 -17057 -31052
rect -16887 -31380 -16562 -31052
rect -16392 -31380 -16067 -31052
rect -15897 -31380 -15572 -31052
rect -15402 -31380 -15077 -31052
rect -14907 -31380 -14582 -31052
rect -14412 -31380 -14087 -31052
rect -13917 -31380 -13592 -31052
rect -13422 -31380 -13097 -31052
rect -12927 -31380 -12602 -31052
rect -12432 -31380 -12107 -31052
rect -11937 -31380 -11612 -31052
rect -11442 -31380 -11117 -31052
rect -10947 -31380 -10622 -31052
rect -10452 -31380 -10127 -31052
rect -9957 -31380 -9632 -31052
rect -9462 -31380 -9137 -31052
rect -8967 -31380 -8642 -31052
rect -8472 -31380 -8147 -31052
rect -7977 -31380 -7652 -31052
rect -7482 -31380 -7157 -31052
rect -6987 -31380 -6662 -31052
rect -6492 -31380 -6167 -31052
rect -5997 -31380 -5672 -31052
rect -5502 -31380 -5177 -31052
rect -5007 -31380 -4682 -31052
rect -4512 -31380 -4187 -31052
rect -4017 -31380 -3692 -31052
rect -3522 -31380 -3197 -31052
rect -3027 -31380 -2702 -31052
rect -2532 -31380 -2207 -31052
rect -2037 -31380 -1712 -31052
rect -1542 -31380 -1217 -31052
rect -1047 -31380 -722 -31052
rect -552 -31380 -227 -31052
rect -57 -31380 268 -31052
rect 438 -31380 763 -31052
rect 933 -31380 1258 -31052
rect 1428 -31380 1753 -31052
rect 1923 -31380 2248 -31052
rect 2418 -31380 2743 -31052
rect 2913 -31380 3238 -31052
rect 3408 -31380 3733 -31052
rect 3903 -31380 4228 -31052
rect 4398 -31380 4723 -31052
rect 4893 -31380 5218 -31052
rect 5388 -31380 5713 -31052
rect 5883 -31380 6208 -31052
rect 6378 -31380 6703 -31052
rect 6873 -31380 7198 -31052
rect 7368 -31380 7693 -31052
rect 7863 -31380 8188 -31052
rect 8358 -31380 8683 -31052
rect 8853 -31380 9178 -31052
rect 9348 -31380 9673 -31052
rect 9843 -31380 10168 -31052
rect 10338 -31380 10663 -31052
rect 10833 -31380 11158 -31052
rect 11328 -31380 11653 -31052
rect 11823 -31380 12148 -31052
rect 12318 -31380 12643 -31052
rect 12813 -31380 13138 -31052
rect 13308 -31380 13633 -31052
rect 13803 -31380 14128 -31052
rect 14298 -31380 14623 -31052
rect 14793 -31380 15118 -31052
rect 15288 -31380 15613 -31052
rect 15783 -31380 16108 -31052
rect 16278 -31380 16603 -31052
rect 16773 -31380 17098 -31052
rect 17268 -31380 17593 -31052
rect 17763 -31380 18088 -31052
rect 18258 -31380 18583 -31052
rect 18753 -31380 19078 -31052
rect 19248 -31380 19573 -31052
rect 19743 -31380 20068 -31052
rect 20238 -31380 20563 -31052
rect 20733 -31380 21058 -31052
rect 21228 -31380 21553 -31052
rect 21723 -31380 22048 -31052
rect 22218 -31380 22543 -31052
rect 22713 -31380 23038 -31052
rect 23208 -31380 23533 -31052
rect 23703 -31380 24028 -31052
rect 24198 -31380 24523 -31052
rect 24693 -31380 25018 -31052
rect 25188 -31380 25513 -31052
rect 25683 -31380 26008 -31052
rect 26178 -31380 26503 -31052
rect 26673 -31380 26998 -31052
rect 27168 -31380 27493 -31052
rect 27663 -31380 27988 -31052
rect 28158 -31380 28483 -31052
rect 28653 -31380 28978 -31052
rect 29148 -31380 29473 -31052
rect 29643 -31380 29968 -31052
rect 30138 -31380 30463 -31052
rect 30633 -31380 30958 -31052
rect 31128 -31380 31453 -31052
rect 31623 -31380 31948 -31052
rect 32118 -31380 32443 -31052
rect 32613 -31380 32938 -31052
rect 33108 -31380 33433 -31052
rect 33603 -31380 33928 -31052
rect 34098 -31380 34423 -31052
rect 34593 -31380 34918 -31052
rect 35088 -31380 35413 -31052
rect 35583 -31380 35908 -31052
rect 36078 -31380 36403 -31052
rect 36573 -31380 36898 -31052
rect 37068 -31380 37393 -31052
rect 37563 -31380 37888 -31052
rect 38058 -31380 38383 -31052
rect 38553 -31380 38878 -31052
rect 39048 -31380 39373 -31052
rect 39543 -31380 39868 -31052
rect 40038 -31380 40363 -31052
rect 40533 -31380 40858 -31052
rect 41028 -31380 41353 -31052
rect 41523 -31380 41848 -31052
rect 42018 -31380 42343 -31052
rect 42513 -31380 42838 -31052
rect 43008 -31380 43333 -31052
rect 43503 -31380 43828 -31052
rect 43998 -31380 44323 -31052
rect 44493 -31380 44818 -31052
rect 44988 -31380 45313 -31052
rect 45483 -31380 45808 -31052
rect 45978 -31380 46303 -31052
rect 46473 -31380 46798 -31052
rect 46968 -31380 47293 -31052
rect 47463 -31380 47788 -31052
rect 47958 -31380 48283 -31052
rect 48453 -31380 48778 -31052
rect 48948 -31380 49273 -31052
rect 49443 -31380 49768 -31052
rect 49938 -31380 50263 -31052
rect 50433 -31380 50758 -31052
rect 50928 -31380 51253 -31052
rect 51423 -31380 51748 -31052
rect 51918 -31380 52243 -31052
rect 52413 -31380 52738 -31052
rect 52908 -31380 53233 -31052
rect 53403 -31380 53728 -31052
rect 53898 -31380 54223 -31052
rect -55497 -31856 -55172 -31528
rect -55002 -31856 -54677 -31528
rect -54507 -31856 -54182 -31528
rect -54012 -31856 -53687 -31528
rect -53517 -31856 -53192 -31528
rect -53022 -31856 -52697 -31528
rect -52527 -31856 -52202 -31528
rect -52032 -31856 -51707 -31528
rect -51537 -31856 -51212 -31528
rect -51042 -31856 -50717 -31528
rect -50547 -31856 -50222 -31528
rect -50052 -31856 -49727 -31528
rect -49557 -31856 -49232 -31528
rect -49062 -31856 -48737 -31528
rect -48567 -31856 -48242 -31528
rect -48072 -31856 -47747 -31528
rect -47577 -31856 -47252 -31528
rect -47082 -31856 -46757 -31528
rect -46587 -31856 -46262 -31528
rect -46092 -31856 -45767 -31528
rect -45597 -31856 -45272 -31528
rect -45102 -31856 -44777 -31528
rect -44607 -31856 -44282 -31528
rect -44112 -31856 -43787 -31528
rect -43617 -31856 -43292 -31528
rect -43122 -31856 -42797 -31528
rect -42627 -31856 -42302 -31528
rect -42132 -31856 -41807 -31528
rect -41637 -31856 -41312 -31528
rect -41142 -31856 -40817 -31528
rect -40647 -31856 -40322 -31528
rect -40152 -31856 -39827 -31528
rect -39657 -31856 -39332 -31528
rect -39162 -31856 -38837 -31528
rect -38667 -31856 -38342 -31528
rect -38172 -31856 -37847 -31528
rect -37677 -31856 -37352 -31528
rect -37182 -31856 -36857 -31528
rect -36687 -31856 -36362 -31528
rect -36192 -31856 -35867 -31528
rect -35697 -31856 -35372 -31528
rect -35202 -31856 -34877 -31528
rect -34707 -31856 -34382 -31528
rect -34212 -31856 -33887 -31528
rect -33717 -31856 -33392 -31528
rect -33222 -31856 -32897 -31528
rect -32727 -31856 -32402 -31528
rect -32232 -31856 -31907 -31528
rect -31737 -31856 -31412 -31528
rect -31242 -31856 -30917 -31528
rect -30747 -31856 -30422 -31528
rect -30252 -31856 -29927 -31528
rect -29757 -31856 -29432 -31528
rect -29262 -31856 -28937 -31528
rect -28767 -31856 -28442 -31528
rect -28272 -31856 -27947 -31528
rect -27777 -31856 -27452 -31528
rect -27282 -31856 -26957 -31528
rect -26787 -31856 -26462 -31528
rect -26292 -31856 -25967 -31528
rect -25797 -31856 -25472 -31528
rect -25302 -31856 -24977 -31528
rect -24807 -31856 -24482 -31528
rect -24312 -31856 -23987 -31528
rect -23817 -31856 -23492 -31528
rect -23322 -31856 -22997 -31528
rect -22827 -31856 -22502 -31528
rect -22332 -31856 -22007 -31528
rect -21837 -31856 -21512 -31528
rect -21342 -31856 -21017 -31528
rect -20847 -31856 -20522 -31528
rect -20352 -31856 -20027 -31528
rect -19857 -31856 -19532 -31528
rect -19362 -31856 -19037 -31528
rect -18867 -31856 -18542 -31528
rect -18372 -31856 -18047 -31528
rect -17877 -31856 -17552 -31528
rect -17382 -31856 -17057 -31528
rect -16887 -31856 -16562 -31528
rect -16392 -31856 -16067 -31528
rect -15897 -31856 -15572 -31528
rect -15402 -31856 -15077 -31528
rect -14907 -31856 -14582 -31528
rect -14412 -31856 -14087 -31528
rect -13917 -31856 -13592 -31528
rect -13422 -31856 -13097 -31528
rect -12927 -31856 -12602 -31528
rect -12432 -31856 -12107 -31528
rect -11937 -31856 -11612 -31528
rect -11442 -31856 -11117 -31528
rect -10947 -31856 -10622 -31528
rect -10452 -31856 -10127 -31528
rect -9957 -31856 -9632 -31528
rect -9462 -31856 -9137 -31528
rect -8967 -31856 -8642 -31528
rect -8472 -31856 -8147 -31528
rect -7977 -31856 -7652 -31528
rect -7482 -31856 -7157 -31528
rect -6987 -31856 -6662 -31528
rect -6492 -31856 -6167 -31528
rect -5997 -31856 -5672 -31528
rect -5502 -31856 -5177 -31528
rect -5007 -31856 -4682 -31528
rect -4512 -31856 -4187 -31528
rect -4017 -31856 -3692 -31528
rect -3522 -31856 -3197 -31528
rect -3027 -31856 -2702 -31528
rect -2532 -31856 -2207 -31528
rect -2037 -31856 -1712 -31528
rect -1542 -31856 -1217 -31528
rect -1047 -31856 -722 -31528
rect -552 -31856 -227 -31528
rect -57 -31856 268 -31528
rect 438 -31856 763 -31528
rect 933 -31856 1258 -31528
rect 1428 -31856 1753 -31528
rect 1923 -31856 2248 -31528
rect 2418 -31856 2743 -31528
rect 2913 -31856 3238 -31528
rect 3408 -31856 3733 -31528
rect 3903 -31856 4228 -31528
rect 4398 -31856 4723 -31528
rect 4893 -31856 5218 -31528
rect 5388 -31856 5713 -31528
rect 5883 -31856 6208 -31528
rect 6378 -31856 6703 -31528
rect 6873 -31856 7198 -31528
rect 7368 -31856 7693 -31528
rect 7863 -31856 8188 -31528
rect 8358 -31856 8683 -31528
rect 8853 -31856 9178 -31528
rect 9348 -31856 9673 -31528
rect 9843 -31856 10168 -31528
rect 10338 -31856 10663 -31528
rect 10833 -31856 11158 -31528
rect 11328 -31856 11653 -31528
rect 11823 -31856 12148 -31528
rect 12318 -31856 12643 -31528
rect 12813 -31856 13138 -31528
rect 13308 -31856 13633 -31528
rect 13803 -31856 14128 -31528
rect 14298 -31856 14623 -31528
rect 14793 -31856 15118 -31528
rect 15288 -31856 15613 -31528
rect 15783 -31856 16108 -31528
rect 16278 -31856 16603 -31528
rect 16773 -31856 17098 -31528
rect 17268 -31856 17593 -31528
rect 17763 -31856 18088 -31528
rect 18258 -31856 18583 -31528
rect 18753 -31856 19078 -31528
rect 19248 -31856 19573 -31528
rect 19743 -31856 20068 -31528
rect 20238 -31856 20563 -31528
rect 20733 -31856 21058 -31528
rect 21228 -31856 21553 -31528
rect 21723 -31856 22048 -31528
rect 22218 -31856 22543 -31528
rect 22713 -31856 23038 -31528
rect 23208 -31856 23533 -31528
rect 23703 -31856 24028 -31528
rect 24198 -31856 24523 -31528
rect 24693 -31856 25018 -31528
rect 25188 -31856 25513 -31528
rect 25683 -31856 26008 -31528
rect 26178 -31856 26503 -31528
rect 26673 -31856 26998 -31528
rect 27168 -31856 27493 -31528
rect 27663 -31856 27988 -31528
rect 28158 -31856 28483 -31528
rect 28653 -31856 28978 -31528
rect 29148 -31856 29473 -31528
rect 29643 -31856 29968 -31528
rect 30138 -31856 30463 -31528
rect 30633 -31856 30958 -31528
rect 31128 -31856 31453 -31528
rect 31623 -31856 31948 -31528
rect 32118 -31856 32443 -31528
rect 32613 -31856 32938 -31528
rect 33108 -31856 33433 -31528
rect 33603 -31856 33928 -31528
rect 34098 -31856 34423 -31528
rect 34593 -31856 34918 -31528
rect 35088 -31856 35413 -31528
rect 35583 -31856 35908 -31528
rect 36078 -31856 36403 -31528
rect 36573 -31856 36898 -31528
rect 37068 -31856 37393 -31528
rect 37563 -31856 37888 -31528
rect 38058 -31856 38383 -31528
rect 38553 -31856 38878 -31528
rect 39048 -31856 39373 -31528
rect 39543 -31856 39868 -31528
rect 40038 -31856 40363 -31528
rect 40533 -31856 40858 -31528
rect 41028 -31856 41353 -31528
rect 41523 -31856 41848 -31528
rect 42018 -31856 42343 -31528
rect 42513 -31856 42838 -31528
rect 43008 -31856 43333 -31528
rect 43503 -31856 43828 -31528
rect 43998 -31856 44323 -31528
rect 44493 -31856 44818 -31528
rect 44988 -31856 45313 -31528
rect 45483 -31856 45808 -31528
rect 45978 -31856 46303 -31528
rect 46473 -31856 46798 -31528
rect 46968 -31856 47293 -31528
rect 47463 -31856 47788 -31528
rect 47958 -31856 48283 -31528
rect 48453 -31856 48778 -31528
rect 48948 -31856 49273 -31528
rect 49443 -31856 49768 -31528
rect 49938 -31856 50263 -31528
rect 50433 -31856 50758 -31528
rect 50928 -31856 51253 -31528
rect 51423 -31856 51748 -31528
rect 51918 -31856 52243 -31528
rect 52413 -31856 52738 -31528
rect 52908 -31856 53233 -31528
rect 53403 -31856 53728 -31528
rect 53898 -31856 54223 -31528
<< nsubdiffcont >>
rect -54870 25814 -54596 26103
rect -54293 25814 -54019 26103
rect -53716 25814 -53442 26103
rect -53139 25814 -52865 26103
rect -52562 25814 -52288 26103
rect -51985 25814 -51711 26103
rect -51408 25814 -51134 26103
rect -50831 25814 -50557 26103
rect -50254 25814 -49980 26103
rect -49677 25814 -49403 26103
rect -49100 25814 -48826 26103
rect -48523 25814 -48249 26103
rect -47946 25814 -47672 26103
rect -47369 25814 -47095 26103
rect -46792 25814 -46518 26103
rect -46215 25814 -45941 26103
rect -45638 25814 -45364 26103
rect -45061 25814 -44787 26103
rect -44484 25814 -44210 26103
rect -43907 25814 -43633 26103
rect -43330 25814 -43056 26103
rect -42753 25814 -42479 26103
rect -42176 25814 -41902 26103
rect -41599 25814 -41325 26103
rect -41022 25814 -40748 26103
rect -40445 25814 -40171 26103
rect -39868 25814 -39594 26103
rect -39291 25814 -39017 26103
rect -38714 25814 -38440 26103
rect -38137 25814 -37863 26103
rect -37560 25814 -37286 26103
rect -36983 25814 -36709 26103
rect -36406 25814 -36132 26103
rect -35829 25814 -35555 26103
rect -35252 25814 -34978 26103
rect -34675 25814 -34401 26103
rect -34098 25814 -33824 26103
rect -33521 25814 -33247 26103
rect -32944 25814 -32670 26103
rect -32367 25814 -32093 26103
rect -31790 25814 -31516 26103
rect -31213 25814 -30939 26103
rect -30636 25814 -30362 26103
rect -30059 25814 -29785 26103
rect -29482 25814 -29208 26103
rect -28905 25814 -28631 26103
rect -28328 25814 -28054 26103
rect -27751 25814 -27477 26103
rect -27174 25814 -26900 26103
rect -26597 25814 -26323 26103
rect -26020 25814 -25746 26103
rect -25443 25814 -25169 26103
rect -24866 25814 -24592 26103
rect -24289 25814 -24015 26103
rect -23712 25814 -23438 26103
rect -23135 25814 -22861 26103
rect -22558 25814 -22284 26103
rect -21981 25814 -21707 26103
rect -21404 25814 -21130 26103
rect -20827 25814 -20553 26103
rect -20250 25814 -19976 26103
rect -19673 25814 -19399 26103
rect -19096 25814 -18822 26103
rect -18519 25814 -18245 26103
rect -17942 25814 -17668 26103
rect -17365 25814 -17091 26103
rect -16788 25814 -16514 26103
rect -16211 25814 -15937 26103
rect -15634 25814 -15360 26103
rect -15057 25814 -14783 26103
rect -14480 25814 -14206 26103
rect -13903 25814 -13629 26103
rect -13326 25814 -13052 26103
rect -12749 25814 -12475 26103
rect -12172 25814 -11898 26103
rect -11595 25814 -11321 26103
rect -11018 25814 -10744 26103
rect -10441 25814 -10167 26103
rect -9864 25814 -9590 26103
rect -9287 25814 -9013 26103
rect -8710 25814 -8436 26103
rect -8133 25814 -7859 26103
rect -7556 25814 -7282 26103
rect -6979 25814 -6705 26103
rect -6402 25814 -6128 26103
rect -5825 25814 -5551 26103
rect -5248 25814 -4974 26103
rect -4671 25814 -4397 26103
rect -4094 25814 -3820 26103
rect -3517 25814 -3243 26103
rect -2940 25814 -2666 26103
rect -2363 25814 -2089 26103
rect -1786 25814 -1512 26103
rect -1209 25814 -935 26103
rect -632 25814 -358 26103
rect -55 25814 219 26103
rect 522 25814 796 26103
rect 1099 25814 1373 26103
rect 1676 25814 1950 26103
rect 2253 25814 2527 26103
rect 2830 25814 3104 26103
rect 3407 25814 3681 26103
rect 3984 25814 4258 26103
rect 4561 25814 4835 26103
rect 5138 25814 5412 26103
rect 5715 25814 5989 26103
rect 6292 25814 6566 26103
rect 6869 25814 7143 26103
rect 7446 25814 7720 26103
rect 8023 25814 8297 26103
rect 8600 25814 8874 26103
rect 9177 25814 9451 26103
rect 9754 25814 10028 26103
rect 10331 25814 10605 26103
rect 10908 25814 11182 26103
rect 11485 25814 11759 26103
rect 12062 25814 12336 26103
rect 12639 25814 12913 26103
rect 13216 25814 13490 26103
rect 13793 25814 14067 26103
rect 14370 25814 14644 26103
rect 14947 25814 15221 26103
rect 15524 25814 15798 26103
rect 16101 25814 16375 26103
rect 16678 25814 16952 26103
rect 17255 25814 17529 26103
rect 17832 25814 18106 26103
rect 18409 25814 18683 26103
rect 18986 25814 19260 26103
rect 19563 25814 19837 26103
rect 20140 25814 20414 26103
rect 20717 25814 20991 26103
rect 21294 25814 21568 26103
rect 21871 25814 22145 26103
rect 22448 25814 22722 26103
rect 23025 25814 23299 26103
rect 23602 25814 23876 26103
rect 24179 25814 24453 26103
rect 24756 25814 25030 26103
rect 25333 25814 25607 26103
rect 25910 25814 26184 26103
rect 26487 25814 26761 26103
rect 27064 25814 27338 26103
rect 27641 25814 27915 26103
rect 28218 25814 28492 26103
rect 28795 25814 29069 26103
rect 29372 25814 29646 26103
rect 29949 25814 30223 26103
rect 30526 25814 30800 26103
rect 31103 25814 31377 26103
rect 31680 25814 31954 26103
rect 32257 25814 32531 26103
rect 32834 25814 33108 26103
rect 33411 25814 33685 26103
rect 33988 25814 34262 26103
rect 34565 25814 34839 26103
rect 35142 25814 35416 26103
rect 35719 25814 35993 26103
rect 36296 25814 36570 26103
rect 36873 25814 37147 26103
rect 37450 25814 37724 26103
rect 38027 25814 38301 26103
rect 38604 25814 38878 26103
rect 39181 25814 39455 26103
rect 39758 25814 40032 26103
rect 40335 25814 40609 26103
rect 40912 25814 41186 26103
rect 41489 25814 41763 26103
rect 42066 25814 42340 26103
rect 42643 25814 42917 26103
rect 43220 25814 43494 26103
rect 43797 25814 44071 26103
rect 44374 25814 44648 26103
rect 44951 25814 45225 26103
rect 45528 25814 45802 26103
rect 46105 25814 46379 26103
rect 46682 25814 46956 26103
rect 47259 25814 47533 26103
rect 47836 25814 48110 26103
rect 48413 25814 48687 26103
rect 48990 25814 49264 26103
rect 49567 25814 49841 26103
rect 50144 25814 50418 26103
rect 50721 25814 50995 26103
rect 51298 25814 51572 26103
rect 51875 25814 52149 26103
rect 52452 25814 52726 26103
rect 53029 25814 53303 26103
rect 53606 25814 53880 26103
rect 54183 25814 54457 26103
rect 54760 25814 55034 26103
rect 55337 25814 55611 26103
rect 55914 25814 56188 26103
rect -54870 25256 -54596 25545
rect -54293 25256 -54019 25545
rect -53716 25256 -53442 25545
rect -53139 25256 -52865 25545
rect -52562 25256 -52288 25545
rect -51985 25256 -51711 25545
rect -51408 25256 -51134 25545
rect -50831 25256 -50557 25545
rect -50254 25256 -49980 25545
rect -49677 25256 -49403 25545
rect -49100 25256 -48826 25545
rect -48523 25256 -48249 25545
rect -47946 25256 -47672 25545
rect -47369 25256 -47095 25545
rect -46792 25256 -46518 25545
rect -46215 25256 -45941 25545
rect -45638 25256 -45364 25545
rect -45061 25256 -44787 25545
rect -44484 25256 -44210 25545
rect -43907 25256 -43633 25545
rect -43330 25256 -43056 25545
rect -42753 25256 -42479 25545
rect -42176 25256 -41902 25545
rect -41599 25256 -41325 25545
rect -41022 25256 -40748 25545
rect -40445 25256 -40171 25545
rect -39868 25256 -39594 25545
rect -39291 25256 -39017 25545
rect -38714 25256 -38440 25545
rect -38137 25256 -37863 25545
rect -37560 25256 -37286 25545
rect -36983 25256 -36709 25545
rect -36406 25256 -36132 25545
rect -35829 25256 -35555 25545
rect -35252 25256 -34978 25545
rect -34675 25256 -34401 25545
rect -34098 25256 -33824 25545
rect -33521 25256 -33247 25545
rect -32944 25256 -32670 25545
rect -32367 25256 -32093 25545
rect -31790 25256 -31516 25545
rect -31213 25256 -30939 25545
rect -30636 25256 -30362 25545
rect -30059 25256 -29785 25545
rect -29482 25256 -29208 25545
rect -28905 25256 -28631 25545
rect -28328 25256 -28054 25545
rect -27751 25256 -27477 25545
rect -27174 25256 -26900 25545
rect -26597 25256 -26323 25545
rect -26020 25256 -25746 25545
rect -25443 25256 -25169 25545
rect -24866 25256 -24592 25545
rect -24289 25256 -24015 25545
rect -23712 25256 -23438 25545
rect -23135 25256 -22861 25545
rect -22558 25256 -22284 25545
rect -21981 25256 -21707 25545
rect -21404 25256 -21130 25545
rect -20827 25256 -20553 25545
rect -20250 25256 -19976 25545
rect -19673 25256 -19399 25545
rect -19096 25256 -18822 25545
rect -18519 25256 -18245 25545
rect -17942 25256 -17668 25545
rect -17365 25256 -17091 25545
rect -16788 25256 -16514 25545
rect -16211 25256 -15937 25545
rect -15634 25256 -15360 25545
rect -15057 25256 -14783 25545
rect -14480 25256 -14206 25545
rect -13903 25256 -13629 25545
rect -13326 25256 -13052 25545
rect -12749 25256 -12475 25545
rect -12172 25256 -11898 25545
rect -11595 25256 -11321 25545
rect -11018 25256 -10744 25545
rect -10441 25256 -10167 25545
rect -9864 25256 -9590 25545
rect -9287 25256 -9013 25545
rect -8710 25256 -8436 25545
rect -8133 25256 -7859 25545
rect -7556 25256 -7282 25545
rect -6979 25256 -6705 25545
rect -6402 25256 -6128 25545
rect -5825 25256 -5551 25545
rect -5248 25256 -4974 25545
rect -4671 25256 -4397 25545
rect -4094 25256 -3820 25545
rect -3517 25256 -3243 25545
rect -2940 25256 -2666 25545
rect -2363 25256 -2089 25545
rect -1786 25256 -1512 25545
rect -1209 25256 -935 25545
rect -632 25256 -358 25545
rect -55 25256 219 25545
rect 522 25256 796 25545
rect 1099 25256 1373 25545
rect 1676 25256 1950 25545
rect 2253 25256 2527 25545
rect 2830 25256 3104 25545
rect 3407 25256 3681 25545
rect 3984 25256 4258 25545
rect 4561 25256 4835 25545
rect 5138 25256 5412 25545
rect 5715 25256 5989 25545
rect 6292 25256 6566 25545
rect 6869 25256 7143 25545
rect 7446 25256 7720 25545
rect 8023 25256 8297 25545
rect 8600 25256 8874 25545
rect 9177 25256 9451 25545
rect 9754 25256 10028 25545
rect 10331 25256 10605 25545
rect 10908 25256 11182 25545
rect 11485 25256 11759 25545
rect 12062 25256 12336 25545
rect 12639 25256 12913 25545
rect 13216 25256 13490 25545
rect 13793 25256 14067 25545
rect 14370 25256 14644 25545
rect 14947 25256 15221 25545
rect 15524 25256 15798 25545
rect 16101 25256 16375 25545
rect 16678 25256 16952 25545
rect 17255 25256 17529 25545
rect 17832 25256 18106 25545
rect 18409 25256 18683 25545
rect 18986 25256 19260 25545
rect 19563 25256 19837 25545
rect 20140 25256 20414 25545
rect 20717 25256 20991 25545
rect 21294 25256 21568 25545
rect 21871 25256 22145 25545
rect 22448 25256 22722 25545
rect 23025 25256 23299 25545
rect 23602 25256 23876 25545
rect 24179 25256 24453 25545
rect 24756 25256 25030 25545
rect 25333 25256 25607 25545
rect 25910 25256 26184 25545
rect 26487 25256 26761 25545
rect 27064 25256 27338 25545
rect 27641 25256 27915 25545
rect 28218 25256 28492 25545
rect 28795 25256 29069 25545
rect 29372 25256 29646 25545
rect 29949 25256 30223 25545
rect 30526 25256 30800 25545
rect 31103 25256 31377 25545
rect 31680 25256 31954 25545
rect 32257 25256 32531 25545
rect 32834 25256 33108 25545
rect 33411 25256 33685 25545
rect 33988 25256 34262 25545
rect 34565 25256 34839 25545
rect 35142 25256 35416 25545
rect 35719 25256 35993 25545
rect 36296 25256 36570 25545
rect 36873 25256 37147 25545
rect 37450 25256 37724 25545
rect 38027 25256 38301 25545
rect 38604 25256 38878 25545
rect 39181 25256 39455 25545
rect 39758 25256 40032 25545
rect 40335 25256 40609 25545
rect 40912 25256 41186 25545
rect 41489 25256 41763 25545
rect 42066 25256 42340 25545
rect 42643 25256 42917 25545
rect 43220 25256 43494 25545
rect 43797 25256 44071 25545
rect 44374 25256 44648 25545
rect 44951 25256 45225 25545
rect 45528 25256 45802 25545
rect 46105 25256 46379 25545
rect 46682 25256 46956 25545
rect 47259 25256 47533 25545
rect 47836 25256 48110 25545
rect 48413 25256 48687 25545
rect 48990 25256 49264 25545
rect 49567 25256 49841 25545
rect 50144 25256 50418 25545
rect 50721 25256 50995 25545
rect 51298 25256 51572 25545
rect 51875 25256 52149 25545
rect 52452 25256 52726 25545
rect 53029 25256 53303 25545
rect 53606 25256 53880 25545
rect 54183 25256 54457 25545
rect 54760 25256 55034 25545
rect 55337 25256 55611 25545
rect 55914 25256 56188 25545
rect -54870 24698 -54596 24987
rect -54293 24698 -54019 24987
rect -53716 24698 -53442 24987
rect -53139 24698 -52865 24987
rect -52562 24698 -52288 24987
rect -51985 24698 -51711 24987
rect -51408 24698 -51134 24987
rect -50831 24698 -50557 24987
rect -50254 24698 -49980 24987
rect -49677 24698 -49403 24987
rect -49100 24698 -48826 24987
rect -48523 24698 -48249 24987
rect -47946 24698 -47672 24987
rect -47369 24698 -47095 24987
rect -46792 24698 -46518 24987
rect -46215 24698 -45941 24987
rect -45638 24698 -45364 24987
rect -45061 24698 -44787 24987
rect -44484 24698 -44210 24987
rect -43907 24698 -43633 24987
rect -43330 24698 -43056 24987
rect -42753 24698 -42479 24987
rect -42176 24698 -41902 24987
rect -41599 24698 -41325 24987
rect -41022 24698 -40748 24987
rect -40445 24698 -40171 24987
rect -39868 24698 -39594 24987
rect -39291 24698 -39017 24987
rect -38714 24698 -38440 24987
rect -38137 24698 -37863 24987
rect -37560 24698 -37286 24987
rect -36983 24698 -36709 24987
rect -36406 24698 -36132 24987
rect -35829 24698 -35555 24987
rect -35252 24698 -34978 24987
rect -34675 24698 -34401 24987
rect -34098 24698 -33824 24987
rect -33521 24698 -33247 24987
rect -32944 24698 -32670 24987
rect -32367 24698 -32093 24987
rect -31790 24698 -31516 24987
rect -31213 24698 -30939 24987
rect -30636 24698 -30362 24987
rect -30059 24698 -29785 24987
rect -29482 24698 -29208 24987
rect -28905 24698 -28631 24987
rect -28328 24698 -28054 24987
rect -27751 24698 -27477 24987
rect -27174 24698 -26900 24987
rect -26597 24698 -26323 24987
rect -26020 24698 -25746 24987
rect -25443 24698 -25169 24987
rect -24866 24698 -24592 24987
rect -24289 24698 -24015 24987
rect -23712 24698 -23438 24987
rect -23135 24698 -22861 24987
rect -22558 24698 -22284 24987
rect -21981 24698 -21707 24987
rect -21404 24698 -21130 24987
rect -20827 24698 -20553 24987
rect -20250 24698 -19976 24987
rect -19673 24698 -19399 24987
rect -19096 24698 -18822 24987
rect -18519 24698 -18245 24987
rect -17942 24698 -17668 24987
rect -17365 24698 -17091 24987
rect -16788 24698 -16514 24987
rect -16211 24698 -15937 24987
rect -15634 24698 -15360 24987
rect -15057 24698 -14783 24987
rect -14480 24698 -14206 24987
rect -13903 24698 -13629 24987
rect -13326 24698 -13052 24987
rect -12749 24698 -12475 24987
rect -12172 24698 -11898 24987
rect -11595 24698 -11321 24987
rect -11018 24698 -10744 24987
rect -10441 24698 -10167 24987
rect -9864 24698 -9590 24987
rect -9287 24698 -9013 24987
rect -8710 24698 -8436 24987
rect -8133 24698 -7859 24987
rect -7556 24698 -7282 24987
rect -6979 24698 -6705 24987
rect -6402 24698 -6128 24987
rect -5825 24698 -5551 24987
rect -5248 24698 -4974 24987
rect -4671 24698 -4397 24987
rect -4094 24698 -3820 24987
rect -3517 24698 -3243 24987
rect -2940 24698 -2666 24987
rect -2363 24698 -2089 24987
rect -1786 24698 -1512 24987
rect -1209 24698 -935 24987
rect -632 24698 -358 24987
rect -55 24698 219 24987
rect 522 24698 796 24987
rect 1099 24698 1373 24987
rect 1676 24698 1950 24987
rect 2253 24698 2527 24987
rect 2830 24698 3104 24987
rect 3407 24698 3681 24987
rect 3984 24698 4258 24987
rect 4561 24698 4835 24987
rect 5138 24698 5412 24987
rect 5715 24698 5989 24987
rect 6292 24698 6566 24987
rect 6869 24698 7143 24987
rect 7446 24698 7720 24987
rect 8023 24698 8297 24987
rect 8600 24698 8874 24987
rect 9177 24698 9451 24987
rect 9754 24698 10028 24987
rect 10331 24698 10605 24987
rect 10908 24698 11182 24987
rect 11485 24698 11759 24987
rect 12062 24698 12336 24987
rect 12639 24698 12913 24987
rect 13216 24698 13490 24987
rect 13793 24698 14067 24987
rect 14370 24698 14644 24987
rect 14947 24698 15221 24987
rect 15524 24698 15798 24987
rect 16101 24698 16375 24987
rect 16678 24698 16952 24987
rect 17255 24698 17529 24987
rect 17832 24698 18106 24987
rect 18409 24698 18683 24987
rect 18986 24698 19260 24987
rect 19563 24698 19837 24987
rect 20140 24698 20414 24987
rect 20717 24698 20991 24987
rect 21294 24698 21568 24987
rect 21871 24698 22145 24987
rect 22448 24698 22722 24987
rect 23025 24698 23299 24987
rect 23602 24698 23876 24987
rect 24179 24698 24453 24987
rect 24756 24698 25030 24987
rect 25333 24698 25607 24987
rect 25910 24698 26184 24987
rect 26487 24698 26761 24987
rect 27064 24698 27338 24987
rect 27641 24698 27915 24987
rect 28218 24698 28492 24987
rect 28795 24698 29069 24987
rect 29372 24698 29646 24987
rect 29949 24698 30223 24987
rect 30526 24698 30800 24987
rect 31103 24698 31377 24987
rect 31680 24698 31954 24987
rect 32257 24698 32531 24987
rect 32834 24698 33108 24987
rect 33411 24698 33685 24987
rect 33988 24698 34262 24987
rect 34565 24698 34839 24987
rect 35142 24698 35416 24987
rect 35719 24698 35993 24987
rect 36296 24698 36570 24987
rect 36873 24698 37147 24987
rect 37450 24698 37724 24987
rect 38027 24698 38301 24987
rect 38604 24698 38878 24987
rect 39181 24698 39455 24987
rect 39758 24698 40032 24987
rect 40335 24698 40609 24987
rect 40912 24698 41186 24987
rect 41489 24698 41763 24987
rect 42066 24698 42340 24987
rect 42643 24698 42917 24987
rect 43220 24698 43494 24987
rect 43797 24698 44071 24987
rect 44374 24698 44648 24987
rect 44951 24698 45225 24987
rect 45528 24698 45802 24987
rect 46105 24698 46379 24987
rect 46682 24698 46956 24987
rect 47259 24698 47533 24987
rect 47836 24698 48110 24987
rect 48413 24698 48687 24987
rect 48990 24698 49264 24987
rect 49567 24698 49841 24987
rect 50144 24698 50418 24987
rect 50721 24698 50995 24987
rect 51298 24698 51572 24987
rect 51875 24698 52149 24987
rect 52452 24698 52726 24987
rect 53029 24698 53303 24987
rect 53606 24698 53880 24987
rect 54183 24698 54457 24987
rect 54760 24698 55034 24987
rect 55337 24698 55611 24987
rect 55914 24698 56188 24987
rect -54870 24140 -54596 24429
rect -54293 24140 -54019 24429
rect -53716 24140 -53442 24429
rect -53139 24140 -52865 24429
rect -52562 24140 -52288 24429
rect -51985 24140 -51711 24429
rect -51408 24140 -51134 24429
rect -50831 24140 -50557 24429
rect -50254 24140 -49980 24429
rect -49677 24140 -49403 24429
rect -49100 24140 -48826 24429
rect -48523 24140 -48249 24429
rect -47946 24140 -47672 24429
rect -47369 24140 -47095 24429
rect -46792 24140 -46518 24429
rect -46215 24140 -45941 24429
rect -45638 24140 -45364 24429
rect -45061 24140 -44787 24429
rect -44484 24140 -44210 24429
rect -43907 24140 -43633 24429
rect -43330 24140 -43056 24429
rect -42753 24140 -42479 24429
rect -42176 24140 -41902 24429
rect -41599 24140 -41325 24429
rect -41022 24140 -40748 24429
rect -40445 24140 -40171 24429
rect -39868 24140 -39594 24429
rect -39291 24140 -39017 24429
rect -38714 24140 -38440 24429
rect -38137 24140 -37863 24429
rect -37560 24140 -37286 24429
rect -36983 24140 -36709 24429
rect -36406 24140 -36132 24429
rect -35829 24140 -35555 24429
rect -35252 24140 -34978 24429
rect -34675 24140 -34401 24429
rect -34098 24140 -33824 24429
rect -33521 24140 -33247 24429
rect -32944 24140 -32670 24429
rect -32367 24140 -32093 24429
rect -31790 24140 -31516 24429
rect -31213 24140 -30939 24429
rect -30636 24140 -30362 24429
rect -30059 24140 -29785 24429
rect -29482 24140 -29208 24429
rect -28905 24140 -28631 24429
rect -28328 24140 -28054 24429
rect -27751 24140 -27477 24429
rect -27174 24140 -26900 24429
rect -26597 24140 -26323 24429
rect -26020 24140 -25746 24429
rect -25443 24140 -25169 24429
rect -24866 24140 -24592 24429
rect -24289 24140 -24015 24429
rect -23712 24140 -23438 24429
rect -23135 24140 -22861 24429
rect -22558 24140 -22284 24429
rect -21981 24140 -21707 24429
rect -21404 24140 -21130 24429
rect -20827 24140 -20553 24429
rect -20250 24140 -19976 24429
rect -19673 24140 -19399 24429
rect -19096 24140 -18822 24429
rect -18519 24140 -18245 24429
rect -17942 24140 -17668 24429
rect -17365 24140 -17091 24429
rect -16788 24140 -16514 24429
rect -16211 24140 -15937 24429
rect -15634 24140 -15360 24429
rect -15057 24140 -14783 24429
rect -14480 24140 -14206 24429
rect -13903 24140 -13629 24429
rect -13326 24140 -13052 24429
rect -12749 24140 -12475 24429
rect -12172 24140 -11898 24429
rect -11595 24140 -11321 24429
rect -11018 24140 -10744 24429
rect -10441 24140 -10167 24429
rect -9864 24140 -9590 24429
rect -9287 24140 -9013 24429
rect -8710 24140 -8436 24429
rect -8133 24140 -7859 24429
rect -7556 24140 -7282 24429
rect -6979 24140 -6705 24429
rect -6402 24140 -6128 24429
rect -5825 24140 -5551 24429
rect -5248 24140 -4974 24429
rect -4671 24140 -4397 24429
rect -4094 24140 -3820 24429
rect -3517 24140 -3243 24429
rect -2940 24140 -2666 24429
rect -2363 24140 -2089 24429
rect -1786 24140 -1512 24429
rect -1209 24140 -935 24429
rect -632 24140 -358 24429
rect -55 24140 219 24429
rect 522 24140 796 24429
rect 1099 24140 1373 24429
rect 1676 24140 1950 24429
rect 2253 24140 2527 24429
rect 2830 24140 3104 24429
rect 3407 24140 3681 24429
rect 3984 24140 4258 24429
rect 4561 24140 4835 24429
rect 5138 24140 5412 24429
rect 5715 24140 5989 24429
rect 6292 24140 6566 24429
rect 6869 24140 7143 24429
rect 7446 24140 7720 24429
rect 8023 24140 8297 24429
rect 8600 24140 8874 24429
rect 9177 24140 9451 24429
rect 9754 24140 10028 24429
rect 10331 24140 10605 24429
rect 10908 24140 11182 24429
rect 11485 24140 11759 24429
rect 12062 24140 12336 24429
rect 12639 24140 12913 24429
rect 13216 24140 13490 24429
rect 13793 24140 14067 24429
rect 14370 24140 14644 24429
rect 14947 24140 15221 24429
rect 15524 24140 15798 24429
rect 16101 24140 16375 24429
rect 16678 24140 16952 24429
rect 17255 24140 17529 24429
rect 17832 24140 18106 24429
rect 18409 24140 18683 24429
rect 18986 24140 19260 24429
rect 19563 24140 19837 24429
rect 20140 24140 20414 24429
rect 20717 24140 20991 24429
rect 21294 24140 21568 24429
rect 21871 24140 22145 24429
rect 22448 24140 22722 24429
rect 23025 24140 23299 24429
rect 23602 24140 23876 24429
rect 24179 24140 24453 24429
rect 24756 24140 25030 24429
rect 25333 24140 25607 24429
rect 25910 24140 26184 24429
rect 26487 24140 26761 24429
rect 27064 24140 27338 24429
rect 27641 24140 27915 24429
rect 28218 24140 28492 24429
rect 28795 24140 29069 24429
rect 29372 24140 29646 24429
rect 29949 24140 30223 24429
rect 30526 24140 30800 24429
rect 31103 24140 31377 24429
rect 31680 24140 31954 24429
rect 32257 24140 32531 24429
rect 32834 24140 33108 24429
rect 33411 24140 33685 24429
rect 33988 24140 34262 24429
rect 34565 24140 34839 24429
rect 35142 24140 35416 24429
rect 35719 24140 35993 24429
rect 36296 24140 36570 24429
rect 36873 24140 37147 24429
rect 37450 24140 37724 24429
rect 38027 24140 38301 24429
rect 38604 24140 38878 24429
rect 39181 24140 39455 24429
rect 39758 24140 40032 24429
rect 40335 24140 40609 24429
rect 40912 24140 41186 24429
rect 41489 24140 41763 24429
rect 42066 24140 42340 24429
rect 42643 24140 42917 24429
rect 43220 24140 43494 24429
rect 43797 24140 44071 24429
rect 44374 24140 44648 24429
rect 44951 24140 45225 24429
rect 45528 24140 45802 24429
rect 46105 24140 46379 24429
rect 46682 24140 46956 24429
rect 47259 24140 47533 24429
rect 47836 24140 48110 24429
rect 48413 24140 48687 24429
rect 48990 24140 49264 24429
rect 49567 24140 49841 24429
rect 50144 24140 50418 24429
rect 50721 24140 50995 24429
rect 51298 24140 51572 24429
rect 51875 24140 52149 24429
rect 52452 24140 52726 24429
rect 53029 24140 53303 24429
rect 53606 24140 53880 24429
rect 54183 24140 54457 24429
rect 54760 24140 55034 24429
rect 55337 24140 55611 24429
rect 55914 24140 56188 24429
<< metal1 >>
rect -55208 26103 56994 26259
rect -55208 25814 -54870 26103
rect -54596 25814 -54293 26103
rect -54019 25814 -53716 26103
rect -53442 25814 -53139 26103
rect -52865 25814 -52562 26103
rect -52288 25814 -51985 26103
rect -51711 25814 -51408 26103
rect -51134 25814 -50831 26103
rect -50557 25814 -50254 26103
rect -49980 25814 -49677 26103
rect -49403 25814 -49100 26103
rect -48826 25814 -48523 26103
rect -48249 25814 -47946 26103
rect -47672 25814 -47369 26103
rect -47095 25814 -46792 26103
rect -46518 25814 -46215 26103
rect -45941 25814 -45638 26103
rect -45364 25814 -45061 26103
rect -44787 25814 -44484 26103
rect -44210 25814 -43907 26103
rect -43633 25814 -43330 26103
rect -43056 25814 -42753 26103
rect -42479 25814 -42176 26103
rect -41902 25814 -41599 26103
rect -41325 25814 -41022 26103
rect -40748 25814 -40445 26103
rect -40171 25814 -39868 26103
rect -39594 25814 -39291 26103
rect -39017 25814 -38714 26103
rect -38440 25814 -38137 26103
rect -37863 25814 -37560 26103
rect -37286 25814 -36983 26103
rect -36709 25814 -36406 26103
rect -36132 25814 -35829 26103
rect -35555 25814 -35252 26103
rect -34978 25814 -34675 26103
rect -34401 25814 -34098 26103
rect -33824 25814 -33521 26103
rect -33247 25814 -32944 26103
rect -32670 25814 -32367 26103
rect -32093 25814 -31790 26103
rect -31516 25814 -31213 26103
rect -30939 25814 -30636 26103
rect -30362 25814 -30059 26103
rect -29785 25814 -29482 26103
rect -29208 25814 -28905 26103
rect -28631 25814 -28328 26103
rect -28054 25814 -27751 26103
rect -27477 25814 -27174 26103
rect -26900 25814 -26597 26103
rect -26323 25814 -26020 26103
rect -25746 25814 -25443 26103
rect -25169 25814 -24866 26103
rect -24592 25814 -24289 26103
rect -24015 25814 -23712 26103
rect -23438 25814 -23135 26103
rect -22861 25814 -22558 26103
rect -22284 25814 -21981 26103
rect -21707 25814 -21404 26103
rect -21130 25814 -20827 26103
rect -20553 25814 -20250 26103
rect -19976 25814 -19673 26103
rect -19399 25814 -19096 26103
rect -18822 25814 -18519 26103
rect -18245 25814 -17942 26103
rect -17668 25814 -17365 26103
rect -17091 25814 -16788 26103
rect -16514 25814 -16211 26103
rect -15937 25814 -15634 26103
rect -15360 25814 -15057 26103
rect -14783 25814 -14480 26103
rect -14206 25814 -13903 26103
rect -13629 25814 -13326 26103
rect -13052 25814 -12749 26103
rect -12475 25814 -12172 26103
rect -11898 25814 -11595 26103
rect -11321 25814 -11018 26103
rect -10744 25814 -10441 26103
rect -10167 25814 -9864 26103
rect -9590 25814 -9287 26103
rect -9013 25814 -8710 26103
rect -8436 25814 -8133 26103
rect -7859 25814 -7556 26103
rect -7282 25814 -6979 26103
rect -6705 25814 -6402 26103
rect -6128 25814 -5825 26103
rect -5551 25814 -5248 26103
rect -4974 25814 -4671 26103
rect -4397 25814 -4094 26103
rect -3820 25814 -3517 26103
rect -3243 25814 -2940 26103
rect -2666 25814 -2363 26103
rect -2089 25814 -1786 26103
rect -1512 25814 -1209 26103
rect -935 25814 -632 26103
rect -358 25814 -55 26103
rect 219 25814 522 26103
rect 796 25814 1099 26103
rect 1373 25814 1676 26103
rect 1950 25814 2253 26103
rect 2527 25814 2830 26103
rect 3104 25814 3407 26103
rect 3681 25814 3984 26103
rect 4258 25814 4561 26103
rect 4835 25814 5138 26103
rect 5412 25814 5715 26103
rect 5989 25814 6292 26103
rect 6566 25814 6869 26103
rect 7143 25814 7446 26103
rect 7720 25814 8023 26103
rect 8297 25814 8600 26103
rect 8874 25814 9177 26103
rect 9451 25814 9754 26103
rect 10028 25814 10331 26103
rect 10605 25814 10908 26103
rect 11182 25814 11485 26103
rect 11759 25814 12062 26103
rect 12336 25814 12639 26103
rect 12913 25814 13216 26103
rect 13490 25814 13793 26103
rect 14067 25814 14370 26103
rect 14644 25814 14947 26103
rect 15221 25814 15524 26103
rect 15798 25814 16101 26103
rect 16375 25814 16678 26103
rect 16952 25814 17255 26103
rect 17529 25814 17832 26103
rect 18106 25814 18409 26103
rect 18683 25814 18986 26103
rect 19260 25814 19563 26103
rect 19837 25814 20140 26103
rect 20414 25814 20717 26103
rect 20991 25814 21294 26103
rect 21568 25814 21871 26103
rect 22145 25814 22448 26103
rect 22722 25814 23025 26103
rect 23299 25814 23602 26103
rect 23876 25814 24179 26103
rect 24453 25814 24756 26103
rect 25030 25814 25333 26103
rect 25607 25814 25910 26103
rect 26184 25814 26487 26103
rect 26761 25814 27064 26103
rect 27338 25814 27641 26103
rect 27915 25814 28218 26103
rect 28492 25814 28795 26103
rect 29069 25814 29372 26103
rect 29646 25814 29949 26103
rect 30223 25814 30526 26103
rect 30800 25814 31103 26103
rect 31377 25814 31680 26103
rect 31954 25814 32257 26103
rect 32531 25814 32834 26103
rect 33108 25814 33411 26103
rect 33685 25814 33988 26103
rect 34262 25814 34565 26103
rect 34839 25814 35142 26103
rect 35416 25814 35719 26103
rect 35993 25814 36296 26103
rect 36570 25814 36873 26103
rect 37147 25814 37450 26103
rect 37724 25814 38027 26103
rect 38301 25814 38604 26103
rect 38878 25814 39181 26103
rect 39455 25814 39758 26103
rect 40032 25814 40335 26103
rect 40609 25814 40912 26103
rect 41186 25814 41489 26103
rect 41763 25814 42066 26103
rect 42340 25814 42643 26103
rect 42917 25814 43220 26103
rect 43494 25814 43797 26103
rect 44071 25814 44374 26103
rect 44648 25814 44951 26103
rect 45225 25814 45528 26103
rect 45802 25814 46105 26103
rect 46379 25814 46682 26103
rect 46956 25814 47259 26103
rect 47533 25814 47836 26103
rect 48110 25814 48413 26103
rect 48687 25814 48990 26103
rect 49264 25814 49567 26103
rect 49841 25814 50144 26103
rect 50418 25814 50721 26103
rect 50995 25814 51298 26103
rect 51572 25814 51875 26103
rect 52149 25814 52452 26103
rect 52726 25814 53029 26103
rect 53303 25814 53606 26103
rect 53880 25814 54183 26103
rect 54457 25814 54760 26103
rect 55034 25814 55337 26103
rect 55611 25814 55914 26103
rect 56188 25814 56994 26103
rect -55208 25545 56994 25814
rect -55208 25256 -54870 25545
rect -54596 25256 -54293 25545
rect -54019 25256 -53716 25545
rect -53442 25256 -53139 25545
rect -52865 25256 -52562 25545
rect -52288 25256 -51985 25545
rect -51711 25256 -51408 25545
rect -51134 25256 -50831 25545
rect -50557 25256 -50254 25545
rect -49980 25256 -49677 25545
rect -49403 25256 -49100 25545
rect -48826 25256 -48523 25545
rect -48249 25256 -47946 25545
rect -47672 25256 -47369 25545
rect -47095 25256 -46792 25545
rect -46518 25256 -46215 25545
rect -45941 25256 -45638 25545
rect -45364 25256 -45061 25545
rect -44787 25256 -44484 25545
rect -44210 25256 -43907 25545
rect -43633 25256 -43330 25545
rect -43056 25256 -42753 25545
rect -42479 25256 -42176 25545
rect -41902 25256 -41599 25545
rect -41325 25256 -41022 25545
rect -40748 25256 -40445 25545
rect -40171 25256 -39868 25545
rect -39594 25256 -39291 25545
rect -39017 25256 -38714 25545
rect -38440 25256 -38137 25545
rect -37863 25256 -37560 25545
rect -37286 25256 -36983 25545
rect -36709 25256 -36406 25545
rect -36132 25256 -35829 25545
rect -35555 25256 -35252 25545
rect -34978 25256 -34675 25545
rect -34401 25256 -34098 25545
rect -33824 25256 -33521 25545
rect -33247 25256 -32944 25545
rect -32670 25256 -32367 25545
rect -32093 25256 -31790 25545
rect -31516 25256 -31213 25545
rect -30939 25256 -30636 25545
rect -30362 25256 -30059 25545
rect -29785 25256 -29482 25545
rect -29208 25256 -28905 25545
rect -28631 25256 -28328 25545
rect -28054 25256 -27751 25545
rect -27477 25256 -27174 25545
rect -26900 25256 -26597 25545
rect -26323 25256 -26020 25545
rect -25746 25256 -25443 25545
rect -25169 25256 -24866 25545
rect -24592 25256 -24289 25545
rect -24015 25256 -23712 25545
rect -23438 25256 -23135 25545
rect -22861 25256 -22558 25545
rect -22284 25256 -21981 25545
rect -21707 25256 -21404 25545
rect -21130 25256 -20827 25545
rect -20553 25256 -20250 25545
rect -19976 25256 -19673 25545
rect -19399 25256 -19096 25545
rect -18822 25256 -18519 25545
rect -18245 25256 -17942 25545
rect -17668 25256 -17365 25545
rect -17091 25256 -16788 25545
rect -16514 25256 -16211 25545
rect -15937 25256 -15634 25545
rect -15360 25256 -15057 25545
rect -14783 25256 -14480 25545
rect -14206 25256 -13903 25545
rect -13629 25256 -13326 25545
rect -13052 25256 -12749 25545
rect -12475 25256 -12172 25545
rect -11898 25256 -11595 25545
rect -11321 25256 -11018 25545
rect -10744 25256 -10441 25545
rect -10167 25256 -9864 25545
rect -9590 25256 -9287 25545
rect -9013 25256 -8710 25545
rect -8436 25256 -8133 25545
rect -7859 25256 -7556 25545
rect -7282 25256 -6979 25545
rect -6705 25256 -6402 25545
rect -6128 25256 -5825 25545
rect -5551 25256 -5248 25545
rect -4974 25256 -4671 25545
rect -4397 25256 -4094 25545
rect -3820 25256 -3517 25545
rect -3243 25256 -2940 25545
rect -2666 25256 -2363 25545
rect -2089 25256 -1786 25545
rect -1512 25256 -1209 25545
rect -935 25256 -632 25545
rect -358 25256 -55 25545
rect 219 25256 522 25545
rect 796 25256 1099 25545
rect 1373 25256 1676 25545
rect 1950 25256 2253 25545
rect 2527 25256 2830 25545
rect 3104 25256 3407 25545
rect 3681 25256 3984 25545
rect 4258 25256 4561 25545
rect 4835 25256 5138 25545
rect 5412 25256 5715 25545
rect 5989 25256 6292 25545
rect 6566 25256 6869 25545
rect 7143 25256 7446 25545
rect 7720 25256 8023 25545
rect 8297 25256 8600 25545
rect 8874 25256 9177 25545
rect 9451 25256 9754 25545
rect 10028 25256 10331 25545
rect 10605 25256 10908 25545
rect 11182 25256 11485 25545
rect 11759 25256 12062 25545
rect 12336 25256 12639 25545
rect 12913 25256 13216 25545
rect 13490 25256 13793 25545
rect 14067 25256 14370 25545
rect 14644 25256 14947 25545
rect 15221 25256 15524 25545
rect 15798 25256 16101 25545
rect 16375 25256 16678 25545
rect 16952 25256 17255 25545
rect 17529 25256 17832 25545
rect 18106 25256 18409 25545
rect 18683 25256 18986 25545
rect 19260 25256 19563 25545
rect 19837 25256 20140 25545
rect 20414 25256 20717 25545
rect 20991 25256 21294 25545
rect 21568 25256 21871 25545
rect 22145 25256 22448 25545
rect 22722 25256 23025 25545
rect 23299 25256 23602 25545
rect 23876 25256 24179 25545
rect 24453 25256 24756 25545
rect 25030 25256 25333 25545
rect 25607 25256 25910 25545
rect 26184 25256 26487 25545
rect 26761 25256 27064 25545
rect 27338 25256 27641 25545
rect 27915 25256 28218 25545
rect 28492 25256 28795 25545
rect 29069 25256 29372 25545
rect 29646 25256 29949 25545
rect 30223 25256 30526 25545
rect 30800 25256 31103 25545
rect 31377 25256 31680 25545
rect 31954 25256 32257 25545
rect 32531 25256 32834 25545
rect 33108 25256 33411 25545
rect 33685 25256 33988 25545
rect 34262 25256 34565 25545
rect 34839 25256 35142 25545
rect 35416 25256 35719 25545
rect 35993 25256 36296 25545
rect 36570 25256 36873 25545
rect 37147 25256 37450 25545
rect 37724 25256 38027 25545
rect 38301 25256 38604 25545
rect 38878 25256 39181 25545
rect 39455 25256 39758 25545
rect 40032 25256 40335 25545
rect 40609 25256 40912 25545
rect 41186 25256 41489 25545
rect 41763 25256 42066 25545
rect 42340 25256 42643 25545
rect 42917 25256 43220 25545
rect 43494 25256 43797 25545
rect 44071 25256 44374 25545
rect 44648 25256 44951 25545
rect 45225 25256 45528 25545
rect 45802 25256 46105 25545
rect 46379 25256 46682 25545
rect 46956 25256 47259 25545
rect 47533 25256 47836 25545
rect 48110 25256 48413 25545
rect 48687 25256 48990 25545
rect 49264 25256 49567 25545
rect 49841 25256 50144 25545
rect 50418 25256 50721 25545
rect 50995 25256 51298 25545
rect 51572 25256 51875 25545
rect 52149 25256 52452 25545
rect 52726 25256 53029 25545
rect 53303 25256 53606 25545
rect 53880 25256 54183 25545
rect 54457 25256 54760 25545
rect 55034 25256 55337 25545
rect 55611 25256 55914 25545
rect 56188 25256 56994 25545
rect -55208 24987 56994 25256
rect -55208 24698 -54870 24987
rect -54596 24698 -54293 24987
rect -54019 24698 -53716 24987
rect -53442 24698 -53139 24987
rect -52865 24698 -52562 24987
rect -52288 24698 -51985 24987
rect -51711 24698 -51408 24987
rect -51134 24698 -50831 24987
rect -50557 24698 -50254 24987
rect -49980 24698 -49677 24987
rect -49403 24698 -49100 24987
rect -48826 24698 -48523 24987
rect -48249 24698 -47946 24987
rect -47672 24698 -47369 24987
rect -47095 24698 -46792 24987
rect -46518 24698 -46215 24987
rect -45941 24698 -45638 24987
rect -45364 24698 -45061 24987
rect -44787 24698 -44484 24987
rect -44210 24698 -43907 24987
rect -43633 24698 -43330 24987
rect -43056 24698 -42753 24987
rect -42479 24698 -42176 24987
rect -41902 24698 -41599 24987
rect -41325 24698 -41022 24987
rect -40748 24698 -40445 24987
rect -40171 24698 -39868 24987
rect -39594 24698 -39291 24987
rect -39017 24698 -38714 24987
rect -38440 24698 -38137 24987
rect -37863 24698 -37560 24987
rect -37286 24698 -36983 24987
rect -36709 24698 -36406 24987
rect -36132 24698 -35829 24987
rect -35555 24698 -35252 24987
rect -34978 24698 -34675 24987
rect -34401 24698 -34098 24987
rect -33824 24698 -33521 24987
rect -33247 24698 -32944 24987
rect -32670 24698 -32367 24987
rect -32093 24698 -31790 24987
rect -31516 24698 -31213 24987
rect -30939 24698 -30636 24987
rect -30362 24698 -30059 24987
rect -29785 24698 -29482 24987
rect -29208 24698 -28905 24987
rect -28631 24698 -28328 24987
rect -28054 24698 -27751 24987
rect -27477 24698 -27174 24987
rect -26900 24698 -26597 24987
rect -26323 24698 -26020 24987
rect -25746 24698 -25443 24987
rect -25169 24698 -24866 24987
rect -24592 24698 -24289 24987
rect -24015 24698 -23712 24987
rect -23438 24698 -23135 24987
rect -22861 24698 -22558 24987
rect -22284 24698 -21981 24987
rect -21707 24698 -21404 24987
rect -21130 24698 -20827 24987
rect -20553 24698 -20250 24987
rect -19976 24698 -19673 24987
rect -19399 24698 -19096 24987
rect -18822 24698 -18519 24987
rect -18245 24698 -17942 24987
rect -17668 24698 -17365 24987
rect -17091 24698 -16788 24987
rect -16514 24698 -16211 24987
rect -15937 24698 -15634 24987
rect -15360 24698 -15057 24987
rect -14783 24698 -14480 24987
rect -14206 24698 -13903 24987
rect -13629 24698 -13326 24987
rect -13052 24698 -12749 24987
rect -12475 24698 -12172 24987
rect -11898 24698 -11595 24987
rect -11321 24698 -11018 24987
rect -10744 24698 -10441 24987
rect -10167 24698 -9864 24987
rect -9590 24698 -9287 24987
rect -9013 24698 -8710 24987
rect -8436 24698 -8133 24987
rect -7859 24698 -7556 24987
rect -7282 24698 -6979 24987
rect -6705 24698 -6402 24987
rect -6128 24698 -5825 24987
rect -5551 24698 -5248 24987
rect -4974 24698 -4671 24987
rect -4397 24698 -4094 24987
rect -3820 24698 -3517 24987
rect -3243 24698 -2940 24987
rect -2666 24698 -2363 24987
rect -2089 24698 -1786 24987
rect -1512 24698 -1209 24987
rect -935 24698 -632 24987
rect -358 24698 -55 24987
rect 219 24698 522 24987
rect 796 24698 1099 24987
rect 1373 24698 1676 24987
rect 1950 24698 2253 24987
rect 2527 24698 2830 24987
rect 3104 24698 3407 24987
rect 3681 24698 3984 24987
rect 4258 24698 4561 24987
rect 4835 24698 5138 24987
rect 5412 24698 5715 24987
rect 5989 24698 6292 24987
rect 6566 24698 6869 24987
rect 7143 24698 7446 24987
rect 7720 24698 8023 24987
rect 8297 24698 8600 24987
rect 8874 24698 9177 24987
rect 9451 24698 9754 24987
rect 10028 24698 10331 24987
rect 10605 24698 10908 24987
rect 11182 24698 11485 24987
rect 11759 24698 12062 24987
rect 12336 24698 12639 24987
rect 12913 24698 13216 24987
rect 13490 24698 13793 24987
rect 14067 24698 14370 24987
rect 14644 24698 14947 24987
rect 15221 24698 15524 24987
rect 15798 24698 16101 24987
rect 16375 24698 16678 24987
rect 16952 24698 17255 24987
rect 17529 24698 17832 24987
rect 18106 24698 18409 24987
rect 18683 24698 18986 24987
rect 19260 24698 19563 24987
rect 19837 24698 20140 24987
rect 20414 24698 20717 24987
rect 20991 24698 21294 24987
rect 21568 24698 21871 24987
rect 22145 24698 22448 24987
rect 22722 24698 23025 24987
rect 23299 24698 23602 24987
rect 23876 24698 24179 24987
rect 24453 24698 24756 24987
rect 25030 24698 25333 24987
rect 25607 24698 25910 24987
rect 26184 24698 26487 24987
rect 26761 24698 27064 24987
rect 27338 24698 27641 24987
rect 27915 24698 28218 24987
rect 28492 24698 28795 24987
rect 29069 24698 29372 24987
rect 29646 24698 29949 24987
rect 30223 24698 30526 24987
rect 30800 24698 31103 24987
rect 31377 24698 31680 24987
rect 31954 24698 32257 24987
rect 32531 24698 32834 24987
rect 33108 24698 33411 24987
rect 33685 24698 33988 24987
rect 34262 24698 34565 24987
rect 34839 24698 35142 24987
rect 35416 24698 35719 24987
rect 35993 24698 36296 24987
rect 36570 24698 36873 24987
rect 37147 24698 37450 24987
rect 37724 24698 38027 24987
rect 38301 24698 38604 24987
rect 38878 24698 39181 24987
rect 39455 24698 39758 24987
rect 40032 24698 40335 24987
rect 40609 24698 40912 24987
rect 41186 24698 41489 24987
rect 41763 24698 42066 24987
rect 42340 24698 42643 24987
rect 42917 24698 43220 24987
rect 43494 24698 43797 24987
rect 44071 24698 44374 24987
rect 44648 24698 44951 24987
rect 45225 24698 45528 24987
rect 45802 24698 46105 24987
rect 46379 24698 46682 24987
rect 46956 24698 47259 24987
rect 47533 24698 47836 24987
rect 48110 24698 48413 24987
rect 48687 24698 48990 24987
rect 49264 24698 49567 24987
rect 49841 24698 50144 24987
rect 50418 24698 50721 24987
rect 50995 24698 51298 24987
rect 51572 24698 51875 24987
rect 52149 24698 52452 24987
rect 52726 24698 53029 24987
rect 53303 24698 53606 24987
rect 53880 24698 54183 24987
rect 54457 24698 54760 24987
rect 55034 24698 55337 24987
rect 55611 24698 55914 24987
rect 56188 24698 56994 24987
rect -55208 24429 56994 24698
rect -55208 24140 -54870 24429
rect -54596 24140 -54293 24429
rect -54019 24140 -53716 24429
rect -53442 24140 -53139 24429
rect -52865 24140 -52562 24429
rect -52288 24140 -51985 24429
rect -51711 24140 -51408 24429
rect -51134 24140 -50831 24429
rect -50557 24140 -50254 24429
rect -49980 24140 -49677 24429
rect -49403 24140 -49100 24429
rect -48826 24140 -48523 24429
rect -48249 24140 -47946 24429
rect -47672 24140 -47369 24429
rect -47095 24140 -46792 24429
rect -46518 24140 -46215 24429
rect -45941 24140 -45638 24429
rect -45364 24140 -45061 24429
rect -44787 24140 -44484 24429
rect -44210 24140 -43907 24429
rect -43633 24140 -43330 24429
rect -43056 24140 -42753 24429
rect -42479 24140 -42176 24429
rect -41902 24140 -41599 24429
rect -41325 24140 -41022 24429
rect -40748 24140 -40445 24429
rect -40171 24140 -39868 24429
rect -39594 24140 -39291 24429
rect -39017 24140 -38714 24429
rect -38440 24140 -38137 24429
rect -37863 24140 -37560 24429
rect -37286 24140 -36983 24429
rect -36709 24140 -36406 24429
rect -36132 24140 -35829 24429
rect -35555 24140 -35252 24429
rect -34978 24140 -34675 24429
rect -34401 24140 -34098 24429
rect -33824 24140 -33521 24429
rect -33247 24140 -32944 24429
rect -32670 24140 -32367 24429
rect -32093 24140 -31790 24429
rect -31516 24140 -31213 24429
rect -30939 24140 -30636 24429
rect -30362 24140 -30059 24429
rect -29785 24140 -29482 24429
rect -29208 24140 -28905 24429
rect -28631 24140 -28328 24429
rect -28054 24140 -27751 24429
rect -27477 24140 -27174 24429
rect -26900 24140 -26597 24429
rect -26323 24140 -26020 24429
rect -25746 24140 -25443 24429
rect -25169 24140 -24866 24429
rect -24592 24140 -24289 24429
rect -24015 24140 -23712 24429
rect -23438 24140 -23135 24429
rect -22861 24140 -22558 24429
rect -22284 24140 -21981 24429
rect -21707 24140 -21404 24429
rect -21130 24140 -20827 24429
rect -20553 24140 -20250 24429
rect -19976 24140 -19673 24429
rect -19399 24140 -19096 24429
rect -18822 24140 -18519 24429
rect -18245 24140 -17942 24429
rect -17668 24140 -17365 24429
rect -17091 24140 -16788 24429
rect -16514 24140 -16211 24429
rect -15937 24140 -15634 24429
rect -15360 24140 -15057 24429
rect -14783 24140 -14480 24429
rect -14206 24140 -13903 24429
rect -13629 24140 -13326 24429
rect -13052 24140 -12749 24429
rect -12475 24140 -12172 24429
rect -11898 24140 -11595 24429
rect -11321 24140 -11018 24429
rect -10744 24140 -10441 24429
rect -10167 24140 -9864 24429
rect -9590 24140 -9287 24429
rect -9013 24140 -8710 24429
rect -8436 24140 -8133 24429
rect -7859 24140 -7556 24429
rect -7282 24140 -6979 24429
rect -6705 24140 -6402 24429
rect -6128 24352 -5825 24429
rect -6128 24339 -5922 24352
rect -6128 24257 -6106 24339
rect -6013 24270 -5922 24339
rect -5829 24270 -5825 24352
rect -6013 24257 -5825 24270
rect -6128 24169 -5825 24257
rect -6128 24156 -5932 24169
rect -6128 24140 -6113 24156
rect -55208 24074 -6113 24140
rect -6020 24087 -5932 24156
rect -5839 24140 -5825 24169
rect -5551 24140 -5248 24429
rect -4974 24140 -4671 24429
rect -4397 24140 -4094 24429
rect -3820 24140 -3517 24429
rect -3243 24140 -2940 24429
rect -2666 24140 -2363 24429
rect -2089 24140 -1786 24429
rect -1512 24140 -1209 24429
rect -935 24140 -632 24429
rect -358 24140 -55 24429
rect 219 24140 522 24429
rect 796 24140 1099 24429
rect 1373 24140 1676 24429
rect 1950 24140 2253 24429
rect 2527 24140 2830 24429
rect 3104 24140 3407 24429
rect 3681 24140 3984 24429
rect 4258 24140 4561 24429
rect 4835 24140 5138 24429
rect 5412 24140 5715 24429
rect 5989 24140 6292 24429
rect 6566 24140 6869 24429
rect 7143 24140 7446 24429
rect 7720 24140 8023 24429
rect 8297 24140 8600 24429
rect 8874 24140 9177 24429
rect 9451 24140 9754 24429
rect 10028 24140 10331 24429
rect 10605 24140 10908 24429
rect 11182 24140 11485 24429
rect 11759 24140 12062 24429
rect 12336 24140 12639 24429
rect 12913 24140 13216 24429
rect 13490 24140 13793 24429
rect 14067 24140 14370 24429
rect 14644 24140 14947 24429
rect 15221 24140 15524 24429
rect 15798 24140 16101 24429
rect 16375 24140 16678 24429
rect 16952 24140 17255 24429
rect 17529 24140 17832 24429
rect 18106 24140 18409 24429
rect 18683 24140 18986 24429
rect 19260 24140 19563 24429
rect 19837 24140 20140 24429
rect 20414 24140 20717 24429
rect 20991 24140 21294 24429
rect 21568 24140 21871 24429
rect 22145 24140 22448 24429
rect 22722 24140 23025 24429
rect 23299 24140 23602 24429
rect 23876 24140 24179 24429
rect 24453 24140 24756 24429
rect 25030 24140 25333 24429
rect 25607 24140 25910 24429
rect 26184 24140 26487 24429
rect 26761 24140 27064 24429
rect 27338 24140 27641 24429
rect 27915 24140 28218 24429
rect 28492 24140 28795 24429
rect 29069 24140 29372 24429
rect 29646 24140 29949 24429
rect 30223 24140 30526 24429
rect 30800 24140 31103 24429
rect 31377 24140 31680 24429
rect 31954 24140 32257 24429
rect 32531 24140 32834 24429
rect 33108 24140 33411 24429
rect 33685 24140 33988 24429
rect 34262 24140 34565 24429
rect 34839 24140 35142 24429
rect 35416 24140 35719 24429
rect 35993 24140 36296 24429
rect 36570 24140 36873 24429
rect 37147 24140 37450 24429
rect 37724 24140 38027 24429
rect 38301 24140 38604 24429
rect 38878 24140 39181 24429
rect 39455 24140 39758 24429
rect 40032 24140 40335 24429
rect 40609 24140 40912 24429
rect 41186 24140 41489 24429
rect 41763 24140 42066 24429
rect 42340 24140 42643 24429
rect 42917 24140 43220 24429
rect 43494 24140 43797 24429
rect 44071 24140 44374 24429
rect 44648 24140 44951 24429
rect 45225 24140 45528 24429
rect 45802 24140 46105 24429
rect 46379 24140 46682 24429
rect 46956 24140 47259 24429
rect 47533 24140 47836 24429
rect 48110 24140 48413 24429
rect 48687 24140 48990 24429
rect 49264 24140 49567 24429
rect 49841 24140 50144 24429
rect 50418 24140 50721 24429
rect 50995 24140 51298 24429
rect 51572 24140 51875 24429
rect 52149 24140 52452 24429
rect 52726 24140 53029 24429
rect 53303 24140 53606 24429
rect 53880 24140 54183 24429
rect 54457 24140 54760 24429
rect 55034 24140 55337 24429
rect 55611 24140 55914 24429
rect 56188 24140 56994 24429
rect -5839 24138 48787 24140
rect -5839 24134 48680 24138
rect -5839 24096 48564 24134
rect -5839 24088 26429 24096
rect -5839 24087 26300 24088
rect -6020 24074 26160 24087
rect -55208 24070 26160 24074
rect -55208 24067 530 24070
rect -55208 24066 418 24067
rect -55208 24007 198 24066
rect 250 24007 307 24066
rect 359 24008 418 24066
rect 470 24011 530 24067
rect 582 24067 1562 24070
rect 582 24066 1450 24067
rect 582 24011 1230 24066
rect 470 24008 1230 24011
rect 359 24007 1230 24008
rect 1282 24007 1339 24066
rect 1391 24008 1450 24066
rect 1502 24011 1562 24067
rect 1614 24017 26160 24070
rect 26233 24018 26300 24087
rect 26373 24026 26429 24088
rect 26502 24084 48564 24096
rect 26502 24082 27850 24084
rect 26502 24077 27699 24082
rect 26502 24026 27546 24077
rect 26373 24018 27546 24026
rect 26233 24017 27546 24018
rect 1614 24011 27546 24017
rect 1502 24009 27546 24011
rect 1502 24008 25018 24009
rect 1391 24007 25018 24008
rect -55208 24002 25018 24007
rect -55208 23996 24864 24002
rect -55208 23984 24725 23996
rect -55208 23979 -5934 23984
rect -55208 23897 -6128 23979
rect -6035 23902 -5934 23979
rect -5841 23956 24725 23984
rect -5841 23955 529 23956
rect -5841 23902 199 23955
rect -6035 23897 199 23902
rect -55208 23896 199 23897
rect 251 23896 308 23955
rect 360 23896 420 23955
rect 472 23897 529 23955
rect 581 23955 1561 23956
rect 581 23897 1231 23955
rect 472 23896 1231 23897
rect 1283 23896 1340 23955
rect 1392 23896 1452 23955
rect 1504 23897 1561 23955
rect 1613 23926 24725 23956
rect 24798 23932 24864 23996
rect 24937 23939 25018 24002
rect 25091 24007 27546 24009
rect 27619 24012 27699 24077
rect 27772 24014 27850 24082
rect 27923 24081 48564 24084
rect 48616 24084 48680 24134
rect 48735 24086 48787 24138
rect 48842 24086 56994 24140
rect 48735 24084 56994 24086
rect 48616 24081 56994 24084
rect 27923 24031 56994 24081
rect 27923 24023 48679 24031
rect 27923 24014 48560 24023
rect 27772 24012 48560 24014
rect 27619 24007 48560 24012
rect 25091 23970 48560 24007
rect 48612 23978 48679 24023
rect 48731 24027 56994 24031
rect 48731 23978 48786 24027
rect 48612 23974 48786 23978
rect 48838 23974 56994 24027
rect 48612 23970 56994 23974
rect 25091 23962 56994 23970
rect 25091 23959 26437 23962
rect 25091 23958 26302 23959
rect 25091 23939 26157 23958
rect 24937 23932 26157 23939
rect 24798 23926 26157 23932
rect 1613 23897 26157 23926
rect 1504 23896 26157 23897
rect -55208 23888 26157 23896
rect 26230 23889 26302 23958
rect 26375 23892 26437 23959
rect 26510 23961 56994 23962
rect 26510 23959 27853 23961
rect 26510 23950 27699 23959
rect 26510 23892 27544 23950
rect 26375 23889 27544 23892
rect 26230 23888 27544 23889
rect -55208 23880 27544 23888
rect 27617 23889 27699 23950
rect 27772 23891 27853 23959
rect 27926 23919 56994 23961
rect 27926 23912 48744 23919
rect 27926 23891 48615 23912
rect 27772 23889 48615 23891
rect 27617 23880 48615 23889
rect -55208 23857 48615 23880
rect 48677 23864 48744 23912
rect 48806 23864 56994 23919
rect 48677 23857 56994 23864
rect -55208 23853 56994 23857
rect 22905 23415 56994 23438
rect 22905 23308 22923 23415
rect 23021 23308 56994 23415
rect 22905 23293 56994 23308
rect 23166 23182 56994 23194
rect 23166 23075 23184 23182
rect 23282 23075 56994 23182
rect 23166 23049 56994 23075
rect 23505 22881 56994 22894
rect 23505 22774 23521 22881
rect 23619 22774 56994 22881
rect 23505 22753 56994 22774
rect -4282 22512 56994 22536
rect -4282 22403 -4271 22512
rect -4129 22403 56994 22512
rect -4282 22395 56994 22403
rect -3601 22330 -3537 22331
rect -3601 22319 56994 22330
rect -3601 22197 -3590 22319
rect -3536 22197 56994 22319
rect -3601 22191 56994 22197
rect -3592 22189 56994 22191
rect 29670 22115 30080 22130
rect 4582 22092 30080 22115
rect 4582 22091 5008 22092
rect 4582 21969 4621 22091
rect 4724 21969 4808 22091
rect 4911 21970 5008 22091
rect 5111 21970 30080 22092
rect 4911 21969 30080 21970
rect 4582 21892 30080 21969
rect 4582 21770 4624 21892
rect 4727 21890 5007 21892
rect 4727 21770 4814 21890
rect 4582 21768 4814 21770
rect 4917 21770 5007 21890
rect 5110 21770 30080 21892
rect 4917 21768 30080 21770
rect 4582 21705 30080 21768
rect 29670 20290 30080 21705
rect -7756 17393 -7534 17403
rect 42596 16872 42621 16920
rect 32263 15615 32288 15663
rect -6188 14854 -5946 14895
rect -6188 14851 -6045 14854
rect -6188 14826 -6169 14851
rect -6692 14782 -6169 14826
rect -6108 14785 -6045 14851
rect -5984 14785 -5946 14854
rect -6108 14782 -5946 14785
rect -6692 14762 -5946 14782
rect -6697 14749 -5946 14762
rect -9915 14728 -5946 14749
rect -9915 14723 -6042 14728
rect -9915 14654 -6171 14723
rect -6110 14659 -6042 14723
rect -5981 14659 -5946 14728
rect -6110 14654 -5946 14659
rect -9915 14646 -5946 14654
rect -6188 14625 -5946 14646
rect -10401 -16877 -10002 13532
rect 42484 9484 42514 9533
rect 32153 8241 32176 8290
rect 49908 -378 50473 -255
rect 56028 -275 56994 -255
rect 56028 -327 56382 -275
rect 56434 -327 56501 -275
rect 56553 -327 56994 -275
rect 56028 -378 56994 -327
rect 49908 -1437 50031 -378
rect 56356 -379 56595 -378
rect 56356 -381 56496 -379
rect 56356 -433 56379 -381
rect 56431 -431 56496 -381
rect 56548 -431 56595 -379
rect 56431 -433 56595 -431
rect 56356 -444 56595 -433
rect 56361 -446 56595 -444
rect 56363 -447 56594 -446
rect 47175 -1923 47489 -1873
rect 47175 -1992 47198 -1923
rect 47271 -1929 47489 -1923
rect 47271 -1992 47373 -1929
rect 47175 -1998 47373 -1992
rect 47446 -1997 47489 -1929
rect 47446 -1998 49164 -1997
rect 47175 -2069 49164 -1998
rect 50037 -2014 50234 -1968
rect 47175 -2088 48944 -2069
rect 47175 -2157 47197 -2088
rect 47270 -2091 48944 -2088
rect 47270 -2157 47370 -2091
rect 47175 -2160 47370 -2157
rect 47443 -2150 48944 -2091
rect 47443 -2160 47489 -2150
rect 47175 -2182 47489 -2160
rect -2662 -2316 -2506 -2307
rect -8299 -2317 -2506 -2316
rect -8459 -2345 -2506 -2317
rect -8459 -2354 -2628 -2345
rect -8459 -2446 -8415 -2354
rect -8338 -2440 -2628 -2354
rect -2537 -2440 -2506 -2345
rect -8338 -2446 -2506 -2440
rect -8459 -2474 -2506 -2446
rect -8459 -2480 -8297 -2474
rect -2662 -2482 -2506 -2474
rect 160 -2532 606 -2516
rect 160 -2535 443 -2532
rect 160 -2631 224 -2535
rect -3347 -2652 224 -2631
rect 341 -2649 443 -2535
rect 560 -2649 606 -2532
rect 341 -2652 606 -2649
rect -3347 -2711 606 -2652
rect -3347 -2720 440 -2711
rect -3347 -2786 221 -2720
rect 160 -2837 221 -2786
rect 338 -2828 440 -2720
rect 557 -2828 606 -2711
rect 338 -2837 606 -2828
rect 160 -2901 606 -2837
rect -6450 -3169 -6259 -3162
rect -6450 -3216 -5955 -3169
rect -6450 -3274 -6441 -3216
rect -6385 -3218 -5955 -3216
rect -6385 -3274 -6333 -3218
rect -6450 -3276 -6333 -3274
rect -6277 -3255 -5955 -3218
rect -4924 -3176 -4822 -3160
rect -4924 -3243 -4906 -3176
rect -4843 -3243 -4822 -3176
rect -2657 -3161 -2500 -3136
rect -2657 -3180 -2624 -3161
rect -2866 -3223 -2624 -3180
rect -2542 -3223 -2500 -3161
rect -2866 -3229 -2500 -3223
rect -6277 -3276 -6259 -3255
rect -4924 -3257 -4822 -3243
rect -2657 -3247 -2500 -3229
rect -6450 -3291 -6259 -3276
rect -8856 -3801 -6006 -3645
rect 49363 -4142 49615 -4114
rect 49363 -4143 49506 -4142
rect 49363 -4205 49385 -4143
rect 49451 -4201 49506 -4143
rect 49569 -4176 49615 -4142
rect 49924 -4176 50015 -2351
rect 56114 -2640 56994 -2569
rect 49569 -4201 50420 -4176
rect 49451 -4205 50420 -4201
rect -5190 -4234 -5133 -4230
rect -3889 -4231 -3795 -4223
rect -5190 -4286 -5187 -4234
rect -5135 -4286 -5133 -4234
rect -5190 -4288 -5133 -4286
rect -3995 -4233 -3795 -4231
rect -3995 -4288 -3876 -4233
rect -3810 -4288 -3795 -4233
rect -3889 -4307 -3795 -4288
rect 49363 -4256 50420 -4205
rect 49363 -4261 49514 -4256
rect 49363 -4323 49380 -4261
rect 49446 -4315 49514 -4261
rect 49577 -4267 50420 -4256
rect 49577 -4315 49615 -4267
rect 49446 -4323 49615 -4315
rect 49363 -4338 49615 -4323
rect 5232 -4959 5370 -4933
rect -5211 -4962 5370 -4959
rect -5218 -4981 5370 -4962
rect -5218 -5003 5255 -4981
rect -5218 -5010 -5077 -5003
rect -5218 -5068 -5193 -5010
rect -5131 -5061 -5077 -5010
rect -5015 -5051 5255 -5003
rect 5326 -5051 5370 -4981
rect 56353 -4961 56587 -4942
rect 56353 -5007 56374 -4961
rect -5015 -5061 5370 -5051
rect -5131 -5068 5370 -5061
rect -5218 -5121 5370 -5068
rect -5218 -5127 5253 -5121
rect -5218 -5185 -5193 -5127
rect -5131 -5185 -5075 -5127
rect -5013 -5185 5253 -5127
rect -5218 -5191 5253 -5185
rect 5324 -5191 5370 -5121
rect -5218 -5204 5370 -5191
rect -5211 -5206 5370 -5204
rect -5078 -5207 5370 -5206
rect 5232 -5220 5370 -5207
rect 50039 -5130 50512 -5007
rect 56161 -5013 56374 -5007
rect 56426 -5013 56493 -4961
rect 56545 -5013 56587 -4961
rect 56161 -5065 56587 -5013
rect 56161 -5067 56488 -5065
rect 56161 -5119 56371 -5067
rect 56423 -5117 56488 -5067
rect 56540 -5117 56587 -5065
rect 56423 -5119 56587 -5117
rect 56161 -5130 56587 -5119
rect 5444 -5401 5564 -5387
rect -6450 -5427 5564 -5401
rect -6450 -5446 5466 -5427
rect -6450 -5504 -6423 -5446
rect -6367 -5492 5466 -5446
rect -6367 -5504 -6315 -5492
rect -6450 -5550 -6315 -5504
rect -6259 -5498 5466 -5492
rect 5531 -5498 5564 -5427
rect -6259 -5550 5564 -5498
rect -6450 -5562 5564 -5550
rect -6450 -5620 -6423 -5562
rect -6367 -5620 5468 -5562
rect -6450 -5633 5468 -5620
rect 5533 -5633 5564 -5562
rect -6450 -5647 5564 -5633
rect -6201 -5649 5564 -5647
rect 5444 -5664 5564 -5649
rect 50039 -6125 50162 -5130
rect 56353 -5132 56587 -5130
rect 56355 -5133 56586 -5132
rect 47766 -6601 48144 -6585
rect 47766 -6681 47793 -6601
rect 47871 -6604 48144 -6601
rect 47871 -6681 47971 -6604
rect 47766 -6684 47971 -6681
rect 48049 -6684 48144 -6604
rect 50137 -6606 50256 -6603
rect 50137 -6659 50281 -6606
rect 47766 -6688 48144 -6684
rect 50092 -6675 50281 -6659
rect 47766 -6736 49174 -6688
rect 50092 -6705 50256 -6675
rect 47766 -6738 47966 -6736
rect 47766 -6818 47792 -6738
rect 47870 -6816 47966 -6738
rect 48044 -6760 49174 -6736
rect 48044 -6816 48144 -6760
rect 50137 -6816 50256 -6705
rect 47870 -6818 48144 -6816
rect 47766 -6877 48144 -6818
rect -7866 -7621 -7591 -7609
rect -7866 -7716 -7693 -7621
rect -7609 -7638 -7591 -7621
rect 3194 -7636 3334 -7626
rect 3194 -7638 3215 -7636
rect -7609 -7703 3215 -7638
rect 3304 -7703 3334 -7636
rect -7609 -7716 3334 -7703
rect -7866 -7730 3334 -7716
rect -7866 -7825 -7836 -7730
rect -7752 -7755 3334 -7730
rect -7752 -7822 3214 -7755
rect 3303 -7822 3334 -7755
rect -7752 -7825 3334 -7822
rect -7866 -7842 3334 -7825
rect -7866 -7850 -7591 -7842
rect 3194 -7858 3334 -7842
rect 49859 -8219 49950 -7083
rect 56182 -7392 56994 -7321
rect 43745 -8605 49950 -8219
rect 49859 -8939 49950 -8605
rect 49859 -9030 50457 -8939
rect 55816 -9255 56994 -9252
rect 55816 -9352 55881 -9255
rect 56139 -9352 56994 -9255
rect 55816 -9356 56994 -9352
rect -6020 -9492 -3288 -9481
rect -6020 -9553 -6009 -9492
rect -5941 -9553 -3288 -9492
rect -6020 -9561 -3288 -9553
rect -6020 -9571 -2701 -9561
rect -3378 -9651 -2701 -9571
rect 4097 -10186 4258 -10174
rect 4097 -10238 4110 -10186
rect 4176 -10238 4258 -10186
rect 4097 -10297 4258 -10238
rect 4097 -10349 4138 -10297
rect 4233 -10349 4258 -10297
rect 4097 -10366 4258 -10349
rect 701 -11602 1077 -11595
rect 701 -11659 1083 -11602
rect 701 -11661 882 -11659
rect 701 -11722 750 -11661
rect 809 -11720 882 -11661
rect 941 -11720 1083 -11659
rect 809 -11722 1083 -11720
rect 701 -11749 1083 -11722
rect 47761 -13575 48160 -13488
rect 8292 -13576 8620 -13575
rect 8292 -13582 25628 -13576
rect 8292 -13591 25459 -13582
rect 8292 -13593 8518 -13591
rect 8292 -13682 8337 -13593
rect 8414 -13680 8518 -13593
rect 8595 -13649 25459 -13591
rect 25555 -13649 25628 -13582
rect 8595 -13680 25628 -13649
rect 8414 -13682 25628 -13680
rect 8292 -13706 25628 -13682
rect 8292 -13736 25453 -13706
rect 8292 -13825 8340 -13736
rect 8417 -13825 8518 -13736
rect 8595 -13805 25453 -13736
rect 25552 -13805 25628 -13706
rect 8595 -13825 25628 -13805
rect 8292 -13873 25628 -13825
rect 42743 -13592 43028 -13576
rect 47761 -13592 47809 -13575
rect 42743 -13603 47809 -13592
rect 42743 -13683 42760 -13603
rect 42838 -13606 47809 -13603
rect 42838 -13683 42938 -13606
rect 42743 -13686 42938 -13683
rect 43016 -13655 47809 -13606
rect 47887 -13578 48160 -13575
rect 47887 -13655 47987 -13578
rect 43016 -13658 47987 -13655
rect 48065 -13658 48160 -13578
rect 43016 -13686 48160 -13658
rect 42743 -13710 48160 -13686
rect 42743 -13712 47982 -13710
rect 42743 -13738 47808 -13712
rect 42743 -13740 42933 -13738
rect 42743 -13820 42759 -13740
rect 42837 -13818 42933 -13740
rect 43011 -13792 47808 -13738
rect 47886 -13790 47982 -13712
rect 48060 -13790 48160 -13710
rect 47886 -13792 48160 -13790
rect 43011 -13805 48160 -13792
rect 43011 -13813 43071 -13805
rect 43011 -13818 43028 -13813
rect 42837 -13820 43028 -13818
rect 42743 -13835 43028 -13820
rect 47761 -13851 48160 -13805
rect 8292 -13897 25452 -13873
rect 8292 -13986 8340 -13897
rect 8417 -13986 8516 -13897
rect 8593 -13972 25452 -13897
rect 25551 -13972 25628 -13873
rect 8593 -13986 25628 -13972
rect 8292 -14013 25628 -13986
rect 8641 -14014 25628 -14013
rect 25393 -14016 25628 -14014
rect 43894 -14201 50243 -14190
rect 43894 -14203 49513 -14201
rect 43894 -14257 49382 -14203
rect 49460 -14255 49513 -14203
rect 49591 -14255 50243 -14201
rect 49460 -14257 50243 -14255
rect 43894 -14308 50243 -14257
rect 43894 -14313 49516 -14308
rect 43894 -14389 49384 -14313
rect 49453 -14384 49516 -14313
rect 49585 -14384 50243 -14308
rect 49453 -14389 50243 -14384
rect 43894 -14452 50243 -14389
rect 43894 -14457 49514 -14452
rect 43894 -14533 49381 -14457
rect 49450 -14528 49514 -14457
rect 49583 -14528 50243 -14452
rect 49450 -14533 50243 -14528
rect 43894 -14550 50243 -14533
rect 49394 -14755 49740 -14739
rect 49394 -14761 49618 -14755
rect -6856 -14805 -6689 -14783
rect -6856 -14889 -6830 -14805
rect -6723 -14889 -6689 -14805
rect -6856 -14908 -6689 -14889
rect 49394 -14839 49422 -14761
rect 49506 -14833 49618 -14761
rect 49702 -14833 49740 -14755
rect 49506 -14839 49740 -14833
rect 49394 -14842 49740 -14839
rect 49394 -14900 50076 -14842
rect 49394 -14908 49616 -14900
rect 49394 -14986 49424 -14908
rect 49508 -14978 49616 -14908
rect 49700 -14968 50084 -14900
rect 49700 -14978 49740 -14968
rect 49508 -14986 49740 -14978
rect 49394 -15006 49740 -14986
rect 9490 -16192 9985 -15247
rect 13232 -15685 13507 -15668
rect 13232 -15767 13245 -15685
rect 13319 -15689 13507 -15685
rect 13319 -15767 13391 -15689
rect 13232 -15771 13391 -15767
rect 13465 -15715 13507 -15689
rect 13465 -15771 50027 -15715
rect 13232 -15772 50027 -15771
rect 13232 -15832 50029 -15772
rect 13232 -15845 13396 -15832
rect 13232 -15927 13244 -15845
rect 13318 -15914 13396 -15845
rect 13470 -15914 50029 -15832
rect 13318 -15927 50029 -15914
rect 13232 -15940 50029 -15927
rect 13232 -15945 13507 -15940
rect 13641 -16090 13920 -16086
rect -15 -16328 9985 -16192
rect 13639 -16092 49616 -16090
rect 13639 -16096 13815 -16092
rect 13639 -16172 13660 -16096
rect 13742 -16168 13815 -16096
rect 13897 -16120 49616 -16092
rect 13897 -16168 49440 -16120
rect 13742 -16172 49440 -16168
rect 13639 -16228 49440 -16172
rect 13639 -16237 13813 -16228
rect 13639 -16313 13662 -16237
rect 13744 -16304 13813 -16237
rect 13895 -16290 49440 -16228
rect 49580 -16290 49616 -16120
rect 13895 -16304 49616 -16290
rect 13744 -16313 49616 -16304
rect 49932 -16306 50029 -15940
rect 13639 -16315 49616 -16313
rect -6069 -16463 -5812 -16406
rect -6069 -16517 -6045 -16463
rect -5991 -16517 -5923 -16463
rect -5869 -16517 -5812 -16463
rect -6069 -16541 -5812 -16517
rect -383 -16541 9985 -16328
rect 13641 -16334 13920 -16315
rect 47139 -16476 47501 -16438
rect 47139 -16480 47356 -16476
rect 47139 -16554 47214 -16480
rect 47292 -16550 47356 -16480
rect 47434 -16550 47501 -16476
rect 47292 -16554 47501 -16550
rect 47139 -16555 47501 -16554
rect 47139 -16607 47941 -16555
rect 47139 -16618 47357 -16607
rect 47139 -16692 47224 -16618
rect 47302 -16681 47357 -16618
rect 47435 -16681 47941 -16607
rect 47302 -16692 47941 -16681
rect 47139 -16734 47941 -16692
rect 14370 -16789 14736 -16761
rect 47139 -16766 47501 -16734
rect 14370 -16793 14539 -16789
rect 14370 -16868 14391 -16793
rect 14455 -16864 14539 -16793
rect 14603 -16864 14669 -16789
rect 14733 -16864 14736 -16789
rect 14455 -16868 14736 -16864
rect -10434 -16924 -9984 -16877
rect -10434 -16929 -10159 -16924
rect -10434 -17050 -10386 -16929
rect -10278 -17045 -10159 -16929
rect -10051 -17045 -9984 -16924
rect -10278 -17050 -9984 -17045
rect -10434 -17140 -9984 -17050
rect -10434 -17144 -10159 -17140
rect -10434 -17265 -10386 -17144
rect -10278 -17261 -10159 -17144
rect -10051 -17261 -9984 -17140
rect -8334 -16895 -8027 -16886
rect 14370 -16895 14736 -16868
rect -8334 -16902 14736 -16895
rect -8334 -16903 -8130 -16902
rect -8334 -17000 -8300 -16903
rect -8210 -16999 -8130 -16903
rect -8040 -16942 14736 -16902
rect -8040 -16943 14669 -16942
rect -8040 -16946 14537 -16943
rect -8040 -16999 14391 -16946
rect -8210 -17000 14391 -16999
rect -8334 -17021 14391 -17000
rect 14455 -17018 14537 -16946
rect 14601 -17017 14669 -16943
rect 14733 -17017 14736 -16942
rect 14601 -17018 14736 -17017
rect 14455 -17021 14736 -17018
rect -8334 -17067 14736 -17021
rect -8334 -17070 -8130 -17067
rect -8334 -17167 -8300 -17070
rect -8210 -17164 -8130 -17070
rect -8040 -17107 14736 -17067
rect -8040 -17164 14391 -17107
rect -8210 -17167 14391 -17164
rect -8334 -17182 14391 -17167
rect 14455 -17182 14530 -17107
rect 14594 -17182 14669 -17107
rect 14733 -17182 14736 -17107
rect -8334 -17197 14736 -17182
rect -8334 -17207 -8027 -17197
rect 14370 -17203 14736 -17197
rect 32750 -17006 43850 -16974
rect 32750 -17128 43704 -17006
rect 43788 -17128 43850 -17006
rect 47762 -17031 47941 -16734
rect 49648 -17009 49898 -16985
rect 49648 -17013 49814 -17009
rect 49648 -17031 49672 -17013
rect 32750 -17151 43850 -17128
rect -10278 -17265 -9984 -17261
rect -10434 -17309 -9984 -17265
rect -3235 -17514 -2995 -17492
rect 4082 -17514 4272 -17505
rect -3235 -17518 4272 -17514
rect -3235 -17676 -3210 -17518
rect -3022 -17532 4272 -17518
rect -3022 -17676 4113 -17532
rect -3235 -17682 4113 -17676
rect 4249 -17682 4272 -17532
rect -3235 -17707 4272 -17682
rect -3235 -17720 -2995 -17707
rect 4082 -17720 4272 -17707
rect 12048 -17976 15387 -17948
rect 12048 -18045 15178 -17976
rect 12049 -18099 15178 -18045
rect 15340 -18099 15387 -17976
rect 32750 -18019 32923 -17151
rect 44085 -17240 47549 -17085
rect 47762 -17087 49672 -17031
rect 49750 -17083 49814 -17013
rect 49892 -17083 49898 -17009
rect 49750 -17087 49898 -17083
rect 47762 -17140 49898 -17087
rect 47762 -17151 49815 -17140
rect 47762 -17210 49682 -17151
rect 44085 -17252 44240 -17240
rect 37186 -17388 37322 -17362
rect 37186 -17492 37209 -17388
rect 37308 -17492 37322 -17388
rect 37186 -17516 37322 -17492
rect 40451 -17407 44240 -17252
rect 40451 -17540 40606 -17407
rect 47394 -17475 47549 -17240
rect 49648 -17225 49682 -17210
rect 49760 -17214 49815 -17151
rect 49893 -17214 49898 -17140
rect 49760 -17225 49898 -17214
rect 49648 -17255 49898 -17225
rect 50389 -17373 50538 -16916
rect 50757 -17408 50906 -16916
rect 51167 -17418 51316 -16926
rect 51546 -17392 51695 -16900
rect -3766 -18108 -3503 -18106
rect -3766 -18136 5129 -18108
rect 12049 -18131 15387 -18099
rect -3766 -18245 -3731 -18136
rect -3599 -18167 5129 -18136
rect -3599 -18168 4918 -18167
rect -3599 -18245 4591 -18168
rect -3766 -18262 4591 -18245
rect 4670 -18170 4918 -18168
rect 4670 -18262 4752 -18170
rect -3766 -18264 4752 -18262
rect 4831 -18261 4918 -18170
rect 4997 -18236 5129 -18167
rect 4997 -18261 5053 -18236
rect 4831 -18264 5053 -18261
rect -3766 -18321 5053 -18264
rect -3766 -18430 -3731 -18321
rect -3599 -18330 5053 -18321
rect 5121 -18330 5129 -18236
rect -3599 -18332 5129 -18330
rect -3599 -18426 4593 -18332
rect 4672 -18426 4753 -18332
rect 4832 -18426 4919 -18332
rect 4998 -18426 5129 -18332
rect -3599 -18430 5129 -18426
rect -3766 -18445 5129 -18430
rect -3737 -18446 5129 -18445
rect 29262 -18381 29419 -18360
rect 29262 -18455 29284 -18381
rect 29359 -18455 29419 -18381
rect 29262 -18466 29419 -18455
rect 31078 -18485 31554 -18459
rect 31078 -18546 31466 -18485
rect 31528 -18546 31554 -18485
rect 31078 -18565 31554 -18546
rect 31818 -18565 32237 -18459
rect 49884 -18633 50008 -18627
rect 49884 -18690 49905 -18633
rect 49979 -18690 50008 -18633
rect 5027 -18723 8565 -18702
rect 5027 -18724 8452 -18723
rect 5027 -18796 8344 -18724
rect 8398 -18795 8452 -18724
rect 8508 -18795 8565 -18723
rect 8398 -18796 8565 -18795
rect 5027 -18974 8565 -18796
rect 11737 -18733 11815 -18700
rect 11737 -18796 11747 -18733
rect 11802 -18796 11815 -18733
rect 49884 -18719 50008 -18690
rect 11737 -18814 11815 -18796
rect 5027 -19081 8375 -18974
rect 8467 -19081 8565 -18974
rect 5027 -19129 8565 -19081
rect 6166 -19469 6449 -19129
rect 42756 -19290 43047 -19224
rect 42756 -19292 42935 -19290
rect 42756 -19364 42792 -19292
rect 42860 -19362 42935 -19292
rect 43003 -19362 43047 -19290
rect 54327 -19320 54506 -19286
rect 42860 -19364 43047 -19362
rect 42756 -19366 43047 -19364
rect 42474 -19414 43047 -19366
rect 54146 -19359 54506 -19320
rect 54146 -19361 54444 -19359
rect 54146 -19368 54340 -19361
rect 42755 -19456 43047 -19414
rect 54327 -19414 54340 -19368
rect 54392 -19412 54444 -19361
rect 54496 -19412 54506 -19359
rect 54392 -19414 54506 -19412
rect 54327 -19426 54506 -19414
rect 6166 -19484 6264 -19469
rect 6166 -19500 6210 -19484
rect 42755 -19528 42789 -19456
rect 42857 -19457 43047 -19456
rect 42857 -19528 42933 -19457
rect 42755 -19529 42933 -19528
rect 43001 -19529 43047 -19457
rect 42755 -19559 43047 -19529
rect 7340 -19753 7460 -19743
rect 7340 -19760 7352 -19753
rect 6903 -19817 7352 -19760
rect 7439 -19761 7460 -19753
rect 7340 -19830 7352 -19817
rect 7441 -19830 7460 -19761
rect 7340 -19844 7460 -19830
rect 14284 -20049 16488 -19898
rect 26336 -20146 27026 -20008
rect -1911 -20279 -1494 -20199
rect -1911 -20381 -1493 -20279
rect 6945 -20325 10177 -20235
rect -1613 -20461 -1493 -20381
rect -3222 -20727 -2992 -20700
rect -3222 -20813 -3171 -20727
rect -3026 -20736 -2992 -20727
rect -3026 -20812 -2750 -20736
rect -1910 -20748 -1861 -20747
rect -1910 -20783 -1551 -20748
rect -3026 -20813 -2992 -20812
rect -3222 -20845 -2992 -20813
rect -1926 -20828 -1551 -20783
rect 5248 -20807 5379 -20785
rect -1459 -20828 -1323 -20827
rect -1926 -20832 -1323 -20828
rect -1607 -20912 -1323 -20832
rect 5248 -20868 5276 -20807
rect 5347 -20828 5379 -20807
rect 7081 -20812 7166 -20797
rect 7081 -20819 7091 -20812
rect 5347 -20868 6027 -20828
rect 6893 -20868 7091 -20819
rect 5248 -20880 6027 -20868
rect 7081 -20878 7091 -20868
rect 7148 -20878 7166 -20812
rect 5248 -20899 5379 -20880
rect 7081 -20893 7166 -20878
rect -1989 -21301 -1372 -21141
rect 10635 -21221 10790 -20541
rect 14868 -20567 15206 -20526
rect 13699 -20573 15206 -20567
rect 13699 -20699 14892 -20573
rect 14868 -20737 14892 -20699
rect 14980 -20737 15064 -20573
rect 15152 -20737 15206 -20573
rect 15918 -20527 16134 -20512
rect 17288 -20527 17469 -20507
rect 15918 -20543 17469 -20527
rect 27339 -20540 27441 -20289
rect 15918 -20638 15936 -20543
rect 15988 -20544 17469 -20543
rect 15988 -20545 17299 -20544
rect 15988 -20638 16040 -20545
rect 15918 -20640 16040 -20638
rect 16092 -20598 17299 -20545
rect 17353 -20545 17469 -20544
rect 17353 -20598 17405 -20545
rect 16092 -20599 17405 -20598
rect 17459 -20599 17469 -20545
rect 25624 -20554 31711 -20540
rect 25624 -20577 26645 -20554
rect 16092 -20610 17469 -20599
rect 16092 -20640 16134 -20610
rect 17288 -20623 17469 -20610
rect 25558 -20580 26645 -20577
rect 15918 -20668 16134 -20640
rect 25558 -20632 25572 -20580
rect 25624 -20627 26645 -20580
rect 26723 -20627 31711 -20554
rect 25624 -20632 31711 -20627
rect 25558 -20642 31711 -20632
rect 14868 -20758 15206 -20737
rect 21126 -20750 21230 -20738
rect 21126 -20815 21142 -20750
rect 21213 -20815 21230 -20750
rect 21126 -20827 21230 -20815
rect 22484 -20753 22562 -20742
rect 22484 -20825 22493 -20753
rect 22553 -20825 22562 -20753
rect 22484 -20836 22562 -20825
rect 13689 -21221 13842 -21215
rect 10588 -21245 13842 -21221
rect 10588 -21350 13712 -21245
rect 13814 -21350 13842 -21245
rect 10588 -21376 13842 -21350
rect 7083 -21406 7183 -21394
rect 13689 -21398 13842 -21376
rect 7083 -21417 8200 -21406
rect 7083 -21489 7104 -21417
rect 7163 -21489 8200 -21417
rect 7083 -21506 8200 -21489
rect 7083 -21510 7183 -21506
rect -3099 -21563 -2985 -21548
rect -3099 -21572 -2604 -21563
rect -3099 -21667 -3084 -21572
rect -3009 -21652 -2604 -21572
rect -3009 -21667 -2985 -21652
rect -3099 -21688 -2985 -21667
rect -1914 -21808 -1721 -21799
rect -1914 -21856 -1789 -21808
rect -1802 -21861 -1789 -21856
rect -1734 -21861 -1721 -21808
rect -1802 -21869 -1721 -21861
rect 7070 -21906 8159 -21817
rect 5743 -21966 5829 -21953
rect 5743 -22022 5753 -21966
rect 5813 -21970 5829 -21966
rect 5813 -22022 6061 -21970
rect 7070 -21985 7165 -21906
rect 5743 -22035 5829 -22022
rect 6846 -22040 7166 -21985
rect 6884 -22053 7166 -22040
rect 14122 -22024 14252 -21991
rect 14122 -22025 14157 -22024
rect 13767 -22090 14157 -22025
rect 14225 -22090 14252 -22024
rect 13767 -22093 14252 -22090
rect -2958 -22114 -2788 -22108
rect -2958 -22362 -1818 -22114
rect 14122 -22128 14252 -22093
rect -2958 -22365 -2450 -22362
rect -1858 -22365 -1818 -22362
rect -2958 -22453 -1818 -22365
rect 26125 -22396 26235 -22364
rect 26125 -22456 26152 -22396
rect 26205 -22456 26235 -22396
rect 11710 -22480 11840 -22460
rect 11327 -22495 11638 -22493
rect 7592 -22524 11638 -22495
rect 7592 -22582 7609 -22524
rect 7664 -22582 11638 -22524
rect 7592 -22596 11638 -22582
rect 11710 -22580 11730 -22480
rect 11830 -22580 11840 -22480
rect 26125 -22483 26235 -22456
rect 7592 -22598 11450 -22596
rect 7592 -22599 7696 -22598
rect 11710 -22600 11840 -22580
rect -1659 -22747 -1504 -22697
rect -1659 -22751 -1563 -22747
rect -3765 -22835 -3504 -22817
rect -3765 -22836 -3461 -22835
rect -3765 -22847 -2790 -22836
rect -1659 -22847 -1586 -22751
rect -3765 -22909 -3725 -22847
rect -3665 -22848 -2790 -22847
rect -3665 -22909 -3602 -22848
rect -3765 -22910 -3602 -22909
rect -3542 -22872 -2790 -22848
rect -3542 -22910 -2759 -22872
rect -1910 -22877 -1586 -22847
rect 38254 -22791 39138 -22773
rect 38254 -22811 39032 -22791
rect 5742 -22871 5828 -22857
rect 5742 -22877 5756 -22871
rect -3765 -22919 -2759 -22910
rect -3765 -22925 -3504 -22919
rect -1949 -22927 -1586 -22877
rect 5359 -22926 5756 -22877
rect 5813 -22926 5828 -22871
rect 14425 -22909 14516 -22862
rect 5359 -22929 5828 -22926
rect 5742 -22939 5828 -22929
rect 13793 -22918 14516 -22909
rect 14622 -22918 14693 -22862
rect 13793 -22972 14693 -22918
rect 38254 -22894 38275 -22811
rect 38353 -22894 39032 -22811
rect 38254 -22895 39032 -22894
rect 39121 -22895 39138 -22791
rect 38254 -22922 39138 -22895
rect 49878 -22850 50019 -22841
rect 49878 -22879 50644 -22850
rect 13793 -22983 14445 -22972
rect 7095 -23012 7210 -22992
rect 7095 -23017 7120 -23012
rect 6903 -23072 7120 -23017
rect 7191 -23072 7210 -23012
rect 13791 -23051 14445 -22983
rect 6903 -23074 7210 -23072
rect 7095 -23089 7210 -23074
rect 14425 -23061 14445 -23051
rect 14521 -23061 14604 -22972
rect 14680 -23061 14693 -22972
rect 49878 -22989 49907 -22879
rect 49996 -22880 50644 -22879
rect 49996 -22989 50534 -22880
rect 49878 -22990 50534 -22989
rect 50623 -22990 50644 -22880
rect 49878 -23017 50644 -22990
rect 49878 -23019 50019 -23017
rect 14425 -23079 14693 -23061
rect -1877 -23387 -1414 -23376
rect -1877 -23447 -1488 -23387
rect -1429 -23447 -1414 -23387
rect -1877 -23457 -1414 -23447
rect 6931 -23403 7695 -23388
rect 6931 -23476 7611 -23403
rect 7680 -23476 7695 -23403
rect 6931 -23491 7695 -23476
rect 6154 -23650 6256 -23646
rect 6154 -23702 6169 -23650
rect 6238 -23651 6256 -23650
rect 6238 -23692 15433 -23651
rect 6238 -23702 10766 -23692
rect 6154 -23755 10766 -23702
rect 6154 -23807 6171 -23755
rect 6240 -23792 10766 -23755
rect 10818 -23792 15433 -23692
rect 6240 -23807 15433 -23792
rect 6154 -23817 15433 -23807
rect 6154 -23823 6256 -23817
rect -1644 -23897 -1570 -23888
rect -1644 -23898 -1635 -23897
rect -1931 -23955 -1635 -23898
rect -1644 -23959 -1635 -23955
rect -1579 -23959 -1570 -23897
rect -1644 -23971 -1570 -23959
rect 5082 -24041 13790 -24027
rect 5082 -24074 8694 -24041
rect 5082 -24141 5895 -24074
rect 5996 -24116 8694 -24074
rect 8777 -24066 13790 -24041
rect 8777 -24116 10918 -24066
rect 5996 -24138 10918 -24116
rect 11078 -24138 13790 -24066
rect 5996 -24141 13790 -24138
rect 5082 -24205 13790 -24141
rect 5082 -24248 10920 -24205
rect 5082 -24250 9412 -24248
rect 5082 -24267 9210 -24250
rect 5082 -24279 5333 -24267
rect 5082 -24393 5131 -24279
rect 5233 -24381 5333 -24279
rect 5435 -24364 9210 -24267
rect 9312 -24362 9412 -24250
rect 9514 -24362 9605 -24248
rect 9707 -24272 10920 -24248
rect 11070 -24268 13790 -24205
rect 11070 -24272 12403 -24268
rect 9707 -24275 12403 -24272
rect 9707 -24328 12251 -24275
rect 9707 -24362 10919 -24328
rect 9312 -24364 10919 -24362
rect 5435 -24381 10919 -24364
rect 5233 -24393 10919 -24381
rect 5082 -24395 10919 -24393
rect 11069 -24365 12251 -24328
rect 12319 -24358 12403 -24275
rect 12471 -24270 12715 -24268
rect 12471 -24358 12555 -24270
rect 12319 -24360 12555 -24358
rect 12623 -24358 12715 -24270
rect 12783 -24358 13790 -24268
rect 12623 -24360 13790 -24358
rect 12319 -24365 13790 -24360
rect 11069 -24395 13790 -24365
rect 5082 -24416 13790 -24395
rect 10881 -24422 11105 -24416
rect -6855 -24460 -1721 -24446
rect -6855 -24463 -6744 -24460
rect -6855 -24519 -6849 -24463
rect -6796 -24518 -6744 -24463
rect -6691 -24462 -1721 -24460
rect -6691 -24518 -1789 -24462
rect -1735 -24518 -1721 -24462
rect -6796 -24519 -1721 -24518
rect -6855 -24530 -1721 -24519
rect 15267 -24447 15433 -23817
rect 21702 -24028 21943 -23975
rect 21702 -24096 21729 -24028
rect 21790 -24029 21943 -24028
rect 21790 -24096 21843 -24029
rect 21702 -24097 21843 -24096
rect 21902 -24097 21943 -24029
rect 21702 -24107 21943 -24097
rect 28151 -24445 28391 -24405
rect 28151 -24447 28195 -24445
rect -6855 -24531 -1822 -24530
rect 15267 -24606 28195 -24447
rect 28352 -24606 28391 -24445
rect 6160 -24630 6290 -24610
rect 15267 -24613 28391 -24606
rect -2650 -24650 6290 -24630
rect 28151 -24639 28391 -24613
rect -2650 -24670 6180 -24650
rect -2650 -24740 -2630 -24670
rect -2570 -24740 6180 -24670
rect -2650 -24750 6180 -24740
rect 6270 -24750 6290 -24650
rect -2650 -24770 6290 -24750
rect 6160 -24780 6290 -24770
rect -1684 -24844 -1540 -24826
rect 4331 -24837 4422 -24827
rect 4331 -24844 4356 -24837
rect -1684 -24846 4356 -24844
rect -1684 -24909 -1652 -24846
rect -1570 -24896 4356 -24846
rect 4413 -24896 4422 -24837
rect -1570 -24901 4422 -24896
rect -1570 -24909 -1540 -24901
rect -1684 -24923 -1540 -24909
rect 4331 -24919 4422 -24901
rect 4536 -25003 4621 -25002
rect -3085 -25014 4621 -25003
rect -3085 -25016 4546 -25014
rect -3085 -25069 -3075 -25016
rect -3017 -25069 4546 -25016
rect -3085 -25084 4546 -25069
rect 4540 -25085 4546 -25084
rect 4608 -25085 4621 -25014
rect 4540 -25098 4621 -25085
rect 32062 -25305 32222 -25063
rect 43671 -25305 43831 -25016
rect 500 -25309 780 -25308
rect -6336 -25449 -5286 -25309
rect 284 -25432 780 -25309
rect -19549 -26481 -19442 -26475
rect -6336 -26534 -6196 -25449
rect -6773 -26651 -6196 -26534
rect -6773 -26657 -6213 -26651
rect 486 -27060 780 -25432
rect 32062 -25334 32223 -25305
rect 32062 -25447 32080 -25334
rect 32192 -25447 32223 -25334
rect 32062 -25471 32223 -25447
rect 43669 -25320 43831 -25305
rect 43669 -25445 43698 -25320
rect 43816 -25445 43831 -25320
rect 43669 -25473 43831 -25445
rect 43671 -25502 43831 -25473
rect 6500 -25730 6620 -25710
rect 6500 -25800 6520 -25730
rect 6590 -25738 6620 -25730
rect 11310 -25738 11420 -25720
rect 6590 -25740 11420 -25738
rect 6590 -25800 11330 -25740
rect 11400 -25800 11420 -25740
rect 6500 -25830 6620 -25800
rect 11310 -25820 11420 -25800
rect 486 -27061 56686 -27060
rect 486 -27101 56938 -27061
rect 486 -27103 56846 -27101
rect -8456 -27177 -7667 -27156
rect -8456 -27183 -8446 -27177
rect -8460 -27301 -8446 -27183
rect -8317 -27219 -7667 -27177
rect -6577 -27190 -5597 -27156
rect -8317 -27291 -7546 -27219
rect -6659 -27225 -5597 -27190
rect 486 -27173 56683 -27103
rect 56771 -27171 56846 -27103
rect 56934 -27171 56938 -27101
rect 56771 -27173 56938 -27171
rect -6659 -27236 -5638 -27225
rect 486 -27232 56938 -27173
rect -6577 -27249 -5638 -27236
rect 500 -27239 56938 -27232
rect 500 -27244 56840 -27239
rect -8317 -27301 -7667 -27291
rect -8460 -27312 -7667 -27301
rect -8456 -27318 -7667 -27312
rect -6577 -27318 -5625 -27249
rect 500 -27314 56680 -27244
rect 56768 -27309 56840 -27244
rect 56928 -27309 56938 -27239
rect 56768 -27314 56938 -27309
rect 500 -27328 56938 -27314
rect 500 -27340 56729 -27328
rect 55845 -27341 56047 -27340
rect 446 -27623 604 -27622
rect -7255 -29213 -7164 -27637
rect 371 -27670 56994 -27623
rect 99 -27720 56994 -27670
rect 446 -27867 56994 -27720
rect -6460 -29213 -6369 -29212
rect -7256 -29283 -5421 -29213
rect -7257 -29304 -5421 -29283
rect -7257 -29479 -5427 -29304
rect -55858 -29579 54839 -29479
rect -55858 -29583 38125 -29579
rect -55858 -29624 38004 -29583
rect 38064 -29624 38125 -29583
rect 38185 -29624 54839 -29579
rect -55858 -29952 -55497 -29624
rect -55172 -29952 -55002 -29624
rect -54677 -29952 -54507 -29624
rect -54182 -29952 -54012 -29624
rect -53687 -29952 -53517 -29624
rect -53192 -29952 -53022 -29624
rect -52697 -29952 -52527 -29624
rect -52202 -29952 -52032 -29624
rect -51707 -29952 -51537 -29624
rect -51212 -29952 -51042 -29624
rect -50717 -29952 -50547 -29624
rect -50222 -29952 -50052 -29624
rect -49727 -29952 -49557 -29624
rect -49232 -29952 -49062 -29624
rect -48737 -29952 -48567 -29624
rect -48242 -29952 -48072 -29624
rect -47747 -29952 -47577 -29624
rect -47252 -29952 -47082 -29624
rect -46757 -29952 -46587 -29624
rect -46262 -29952 -46092 -29624
rect -45767 -29952 -45597 -29624
rect -45272 -29952 -45102 -29624
rect -44777 -29952 -44607 -29624
rect -44282 -29952 -44112 -29624
rect -43787 -29952 -43617 -29624
rect -43292 -29952 -43122 -29624
rect -42797 -29952 -42627 -29624
rect -42302 -29952 -42132 -29624
rect -41807 -29952 -41637 -29624
rect -41312 -29952 -41142 -29624
rect -40817 -29952 -40647 -29624
rect -40322 -29952 -40152 -29624
rect -39827 -29952 -39657 -29624
rect -39332 -29952 -39162 -29624
rect -38837 -29952 -38667 -29624
rect -38342 -29952 -38172 -29624
rect -37847 -29952 -37677 -29624
rect -37352 -29952 -37182 -29624
rect -36857 -29952 -36687 -29624
rect -36362 -29952 -36192 -29624
rect -35867 -29952 -35697 -29624
rect -35372 -29952 -35202 -29624
rect -34877 -29952 -34707 -29624
rect -34382 -29952 -34212 -29624
rect -33887 -29952 -33717 -29624
rect -33392 -29952 -33222 -29624
rect -32897 -29952 -32727 -29624
rect -32402 -29952 -32232 -29624
rect -31907 -29952 -31737 -29624
rect -31412 -29952 -31242 -29624
rect -30917 -29952 -30747 -29624
rect -30422 -29952 -30252 -29624
rect -29927 -29952 -29757 -29624
rect -29432 -29952 -29262 -29624
rect -28937 -29952 -28767 -29624
rect -28442 -29952 -28272 -29624
rect -27947 -29952 -27777 -29624
rect -27452 -29821 -27282 -29624
rect -26957 -29816 -26787 -29624
rect -27452 -29921 -27343 -29821
rect -26911 -29916 -26787 -29816
rect -27452 -29952 -27282 -29921
rect -26957 -29952 -26787 -29916
rect -26462 -29952 -26292 -29624
rect -25967 -29952 -25797 -29624
rect -25472 -29952 -25302 -29624
rect -24977 -29798 -24807 -29624
rect -24482 -29778 -24312 -29624
rect -24977 -29898 -24934 -29798
rect -24851 -29898 -24807 -29798
rect -24459 -29878 -24312 -29778
rect -24977 -29952 -24807 -29898
rect -24482 -29952 -24312 -29878
rect -23987 -29952 -23817 -29624
rect -23492 -29952 -23322 -29624
rect -22997 -29952 -22827 -29624
rect -22502 -29793 -22332 -29624
rect -22007 -29788 -21837 -29624
rect -22502 -29893 -22352 -29793
rect -22007 -29888 -21972 -29788
rect -21889 -29888 -21837 -29788
rect -22502 -29952 -22332 -29893
rect -22007 -29952 -21837 -29888
rect -21512 -29952 -21342 -29624
rect -21017 -29952 -20847 -29624
rect -20522 -29952 -20352 -29624
rect -20027 -29952 -19857 -29624
rect -19532 -29787 -19362 -29624
rect -19532 -29796 -19407 -29787
rect -19515 -29887 -19407 -29796
rect -19515 -29896 -19362 -29887
rect -19532 -29952 -19362 -29896
rect -19037 -29952 -18867 -29624
rect -18542 -29952 -18372 -29624
rect -18047 -29952 -17877 -29624
rect -17552 -29952 -17382 -29624
rect -17057 -29778 -16887 -29624
rect -17035 -29878 -16929 -29778
rect -17057 -29952 -16887 -29878
rect -16562 -29952 -16392 -29624
rect -16067 -29952 -15897 -29624
rect -15572 -29952 -15402 -29624
rect -15077 -29952 -14907 -29624
rect -14582 -29952 -14412 -29624
rect -14087 -29784 -13917 -29624
rect -14087 -29884 -14030 -29784
rect -13947 -29884 -13917 -29784
rect -14087 -29952 -13917 -29884
rect -13592 -29952 -13422 -29624
rect -13097 -29952 -12927 -29624
rect -12602 -29952 -12432 -29624
rect -12107 -29784 -11937 -29624
rect -11612 -29778 -11442 -29624
rect -12107 -29884 -11942 -29784
rect -11612 -29878 -11552 -29778
rect -11469 -29878 -11442 -29778
rect -12107 -29952 -11937 -29884
rect -11612 -29952 -11442 -29878
rect -11117 -29952 -10947 -29624
rect -10622 -29952 -10452 -29624
rect -10127 -29952 -9957 -29624
rect -9632 -29952 -9462 -29624
rect -9137 -29952 -8967 -29624
rect -8642 -29952 -8472 -29624
rect -8147 -29952 -7977 -29624
rect -7652 -29952 -7482 -29624
rect -7157 -29952 -6987 -29624
rect -6662 -29952 -6492 -29624
rect -6167 -29816 -5997 -29624
rect -6167 -29881 -6034 -29816
rect -6167 -29948 -5997 -29881
rect -6167 -29952 -6034 -29948
rect -5672 -29952 -5502 -29624
rect -5177 -29952 -5007 -29624
rect -4682 -29952 -4512 -29624
rect -4187 -29952 -4017 -29624
rect -3692 -29952 -3522 -29624
rect -3197 -29952 -3027 -29624
rect -2702 -29952 -2532 -29624
rect -2207 -29952 -2037 -29624
rect -1712 -29952 -1542 -29624
rect -1217 -29952 -1047 -29624
rect -722 -29952 -552 -29624
rect -227 -29952 -57 -29624
rect 268 -29952 438 -29624
rect 763 -29874 933 -29624
rect 763 -29882 929 -29874
rect -55858 -29969 -6034 -29952
rect -55858 -29971 -11559 -29969
rect -55858 -29974 -21978 -29971
rect -55858 -29980 -24537 -29974
rect -55858 -29994 -24738 -29980
rect -55858 -30008 -24929 -29994
rect -55858 -30019 -26978 -30008
rect -55858 -30021 -27170 -30019
rect -55858 -30080 -27348 -30021
rect -27265 -30080 -27170 -30021
rect -27087 -30080 -26978 -30019
rect -26895 -30080 -24929 -30008
rect -24846 -30080 -24738 -29994
rect -24655 -30074 -24537 -29980
rect -24454 -29976 -21978 -29974
rect -24454 -30074 -22358 -29976
rect -24655 -30076 -22358 -30074
rect -22275 -30076 -22171 -29976
rect -22088 -30071 -21978 -29976
rect -21895 -29974 -14025 -29971
rect -21895 -29976 -19411 -29974
rect -21895 -29992 -19603 -29976
rect -21895 -30071 -19821 -29992
rect -22088 -30076 -19821 -30071
rect -24655 -30080 -19821 -30076
rect -19738 -30076 -19603 -29992
rect -19520 -30074 -19411 -29976
rect -19328 -29980 -14203 -29974
rect -19328 -29985 -14383 -29980
rect -19328 -30074 -17303 -29985
rect -19520 -30076 -17303 -30074
rect -19738 -30080 -17303 -30076
rect -17220 -29987 -16918 -29985
rect -17220 -30080 -17116 -29987
rect -17033 -30080 -16918 -29987
rect -16835 -30080 -14383 -29985
rect -14300 -30074 -14203 -29980
rect -14120 -30071 -14025 -29974
rect -13942 -29978 -11559 -29971
rect -13942 -29990 -11734 -29978
rect -13942 -30071 -11949 -29990
rect -14120 -30074 -11949 -30071
rect -14300 -30080 -11949 -30074
rect -11866 -30078 -11734 -29990
rect -11651 -30069 -11559 -29978
rect -11476 -30013 -6034 -29969
rect -5973 -30013 -5906 -29952
rect -5845 -29996 750 -29952
rect 852 -29988 929 -29882
rect 1258 -29952 1428 -29624
rect 1753 -29952 1923 -29624
rect 2248 -29952 2418 -29624
rect 2743 -29952 2913 -29624
rect 3238 -29952 3408 -29624
rect 3733 -29952 3903 -29624
rect 4228 -29952 4398 -29624
rect 4723 -29952 4893 -29624
rect 5218 -29812 5388 -29624
rect 5218 -29925 5287 -29812
rect 5381 -29925 5388 -29812
rect 5218 -29952 5388 -29925
rect 5713 -29952 5883 -29624
rect 6208 -29952 6378 -29624
rect 6703 -29952 6873 -29624
rect 7198 -29952 7368 -29624
rect 7693 -29952 7863 -29624
rect 8188 -29952 8358 -29624
rect 8683 -29952 8853 -29624
rect 9178 -29854 9348 -29624
rect 9178 -29952 9213 -29854
rect 1031 -29988 1105 -29952
rect 852 -29996 1105 -29988
rect 1207 -29964 9213 -29952
rect 9298 -29952 9348 -29854
rect 9673 -29952 9843 -29624
rect 10168 -29952 10338 -29624
rect 10663 -29952 10833 -29624
rect 11158 -29952 11328 -29624
rect 11653 -29952 11823 -29624
rect 12148 -29781 12318 -29624
rect 12148 -29871 12243 -29781
rect 12311 -29871 12318 -29781
rect 12643 -29775 12813 -29624
rect 12643 -29865 12700 -29775
rect 12768 -29865 12813 -29775
rect 12148 -29952 12318 -29871
rect 12643 -29952 12813 -29865
rect 13138 -29952 13308 -29624
rect 13633 -29952 13803 -29624
rect 14128 -29952 14298 -29624
rect 14623 -29952 14793 -29624
rect 15118 -29952 15288 -29624
rect 15613 -29952 15783 -29624
rect 16108 -29952 16278 -29624
rect 16603 -29952 16773 -29624
rect 17098 -29952 17268 -29624
rect 17593 -29952 17763 -29624
rect 18088 -29952 18258 -29624
rect 18583 -29952 18753 -29624
rect 19078 -29952 19248 -29624
rect 19573 -29952 19743 -29624
rect 20068 -29952 20238 -29624
rect 20563 -29937 20733 -29624
rect 20572 -29952 20733 -29937
rect 21058 -29759 21228 -29624
rect 21058 -29827 21109 -29759
rect 21170 -29827 21228 -29759
rect 21058 -29892 21228 -29827
rect 21553 -29869 21723 -29624
rect 21058 -29952 21107 -29892
rect 9298 -29964 9372 -29952
rect 1207 -29966 9372 -29964
rect 9457 -29964 9539 -29952
rect 9624 -29964 12229 -29952
rect 9457 -29966 12229 -29964
rect 1207 -29996 12229 -29966
rect -5845 -30013 12229 -29996
rect -11476 -30019 12229 -30013
rect -11476 -30021 5287 -30019
rect -11476 -30026 5100 -30021
rect -11476 -30069 4921 -30026
rect -11651 -30078 4921 -30069
rect -11866 -30080 4921 -30078
rect 5015 -30080 5100 -30026
rect 5194 -30080 5287 -30021
rect 5381 -30042 12229 -30019
rect 12297 -30031 12383 -29952
rect 12451 -30031 12545 -29952
rect 12297 -30036 12545 -30031
rect 12613 -29954 20376 -29952
rect 12613 -30036 12708 -29954
rect 12297 -30042 12708 -30036
rect 5381 -30044 12708 -30042
rect 12776 -30008 20376 -29954
rect 20441 -30006 20507 -29952
rect 20572 -29960 21107 -29952
rect 21168 -29952 21228 -29892
rect 21553 -29937 21717 -29869
rect 21553 -29952 21723 -29937
rect 22048 -29952 22218 -29624
rect 22543 -29952 22713 -29624
rect 23038 -29952 23208 -29624
rect 23533 -29952 23703 -29624
rect 24028 -29952 24198 -29624
rect 24523 -29952 24693 -29624
rect 25018 -29952 25188 -29624
rect 25513 -29952 25683 -29624
rect 26008 -29952 26178 -29624
rect 26503 -29952 26673 -29624
rect 26998 -29952 27168 -29624
rect 27493 -29952 27663 -29624
rect 27988 -29952 28158 -29624
rect 28483 -29952 28653 -29624
rect 28978 -29952 29148 -29624
rect 29473 -29952 29643 -29624
rect 29968 -29952 30138 -29624
rect 30463 -29952 30633 -29624
rect 30958 -29952 31128 -29624
rect 31453 -29952 31623 -29624
rect 31948 -29952 32118 -29624
rect 32443 -29952 32613 -29624
rect 32938 -29952 33108 -29624
rect 33433 -29952 33603 -29624
rect 33928 -29805 34098 -29624
rect 33939 -29863 34098 -29805
rect 33928 -29952 34098 -29863
rect 34423 -29952 34593 -29624
rect 34918 -29952 35088 -29624
rect 35413 -29952 35583 -29624
rect 35908 -29952 36078 -29624
rect 36403 -29809 36573 -29624
rect 36403 -29867 36560 -29809
rect 36403 -29952 36573 -29867
rect 36898 -29952 37068 -29624
rect 37393 -29952 37563 -29624
rect 37888 -29642 38004 -29624
rect 37888 -29694 38058 -29642
rect 37888 -29753 38005 -29694
rect 37888 -29807 38058 -29753
rect 37888 -29866 38007 -29807
rect 37888 -29952 38058 -29866
rect 38383 -29952 38553 -29624
rect 38878 -29952 39048 -29624
rect 39373 -29952 39543 -29624
rect 39868 -29952 40038 -29624
rect 40363 -29952 40533 -29624
rect 40858 -29952 41028 -29624
rect 41353 -29952 41523 -29624
rect 41848 -29952 42018 -29624
rect 42343 -29952 42513 -29624
rect 42838 -29952 43008 -29624
rect 43333 -29952 43503 -29624
rect 43828 -29952 43998 -29624
rect 44323 -29952 44493 -29624
rect 44818 -29952 44988 -29624
rect 45313 -29952 45483 -29624
rect 45808 -29793 45978 -29624
rect 45808 -29810 45839 -29793
rect 45893 -29794 45978 -29793
rect 45808 -29873 45820 -29810
rect 45893 -29851 45946 -29794
rect 45874 -29852 45946 -29851
rect 45874 -29870 45960 -29852
rect 45874 -29873 45978 -29870
rect 45808 -29952 45978 -29873
rect 46303 -29952 46473 -29624
rect 46798 -29792 46968 -29624
rect 46798 -29860 46955 -29792
rect 46798 -29952 46968 -29860
rect 47293 -29952 47463 -29624
rect 47788 -29770 47958 -29624
rect 47788 -29833 47957 -29770
rect 47788 -29952 47958 -29833
rect 48283 -29952 48453 -29624
rect 48778 -29952 48948 -29624
rect 49273 -29801 49443 -29624
rect 49315 -29864 49377 -29801
rect 49431 -29864 49443 -29801
rect 49273 -29952 49443 -29864
rect 49768 -29952 49938 -29624
rect 50263 -29952 50433 -29624
rect 50758 -29952 50928 -29624
rect 51253 -29952 51423 -29624
rect 51748 -29952 51918 -29624
rect 52243 -29952 52413 -29624
rect 52738 -29952 52908 -29624
rect 53233 -29952 53403 -29624
rect 53728 -29952 53898 -29624
rect 54223 -29952 54839 -29624
rect 21168 -29956 21249 -29952
rect 21310 -29956 54839 -29952
rect 21168 -29960 54839 -29956
rect 20572 -30006 54839 -29960
rect 20441 -30008 54839 -30006
rect 12776 -30044 54839 -30008
rect 5381 -30080 54839 -30044
rect -55858 -30100 54839 -30080
rect -55858 -30428 -55497 -30100
rect -55172 -30428 -55002 -30100
rect -54677 -30428 -54507 -30100
rect -54182 -30428 -54012 -30100
rect -53687 -30428 -53517 -30100
rect -53192 -30428 -53022 -30100
rect -52697 -30428 -52527 -30100
rect -52202 -30428 -52032 -30100
rect -51707 -30428 -51537 -30100
rect -51212 -30428 -51042 -30100
rect -50717 -30428 -50547 -30100
rect -50222 -30428 -50052 -30100
rect -49727 -30428 -49557 -30100
rect -49232 -30428 -49062 -30100
rect -48737 -30428 -48567 -30100
rect -48242 -30428 -48072 -30100
rect -47747 -30428 -47577 -30100
rect -47252 -30428 -47082 -30100
rect -46757 -30428 -46587 -30100
rect -46262 -30428 -46092 -30100
rect -45767 -30428 -45597 -30100
rect -45272 -30428 -45102 -30100
rect -44777 -30428 -44607 -30100
rect -44282 -30428 -44112 -30100
rect -43787 -30428 -43617 -30100
rect -43292 -30428 -43122 -30100
rect -42797 -30428 -42627 -30100
rect -42302 -30428 -42132 -30100
rect -41807 -30428 -41637 -30100
rect -41312 -30428 -41142 -30100
rect -40817 -30428 -40647 -30100
rect -40322 -30428 -40152 -30100
rect -39827 -30428 -39657 -30100
rect -39332 -30428 -39162 -30100
rect -38837 -30428 -38667 -30100
rect -38342 -30428 -38172 -30100
rect -37847 -30428 -37677 -30100
rect -37352 -30428 -37182 -30100
rect -36857 -30428 -36687 -30100
rect -36362 -30428 -36192 -30100
rect -35867 -30428 -35697 -30100
rect -35372 -30428 -35202 -30100
rect -34877 -30428 -34707 -30100
rect -34382 -30428 -34212 -30100
rect -33887 -30428 -33717 -30100
rect -33392 -30428 -33222 -30100
rect -32897 -30428 -32727 -30100
rect -32402 -30428 -32232 -30100
rect -31907 -30428 -31737 -30100
rect -31412 -30428 -31242 -30100
rect -30917 -30428 -30747 -30100
rect -30422 -30428 -30252 -30100
rect -29927 -30428 -29757 -30100
rect -29432 -30428 -29262 -30100
rect -28937 -30428 -28767 -30100
rect -28442 -30428 -28272 -30100
rect -27947 -30428 -27777 -30100
rect -27452 -30428 -27282 -30100
rect -26957 -30428 -26787 -30100
rect -26462 -30428 -26292 -30100
rect -25967 -30428 -25797 -30100
rect -25472 -30428 -25302 -30100
rect -24977 -30428 -24807 -30100
rect -24482 -30428 -24312 -30100
rect -23987 -30428 -23817 -30100
rect -23492 -30428 -23322 -30100
rect -22997 -30428 -22827 -30100
rect -22502 -30428 -22332 -30100
rect -22007 -30428 -21837 -30100
rect -21512 -30428 -21342 -30100
rect -21017 -30428 -20847 -30100
rect -20522 -30428 -20352 -30100
rect -20027 -30428 -19857 -30100
rect -19532 -30428 -19362 -30100
rect -19037 -30428 -18867 -30100
rect -18542 -30428 -18372 -30100
rect -18047 -30428 -17877 -30100
rect -17552 -30428 -17382 -30100
rect -17057 -30428 -16887 -30100
rect -16562 -30428 -16392 -30100
rect -16067 -30428 -15897 -30100
rect -15572 -30428 -15402 -30100
rect -15077 -30428 -14907 -30100
rect -14582 -30428 -14412 -30100
rect -14087 -30428 -13917 -30100
rect -13592 -30428 -13422 -30100
rect -13097 -30428 -12927 -30100
rect -12602 -30428 -12432 -30100
rect -12107 -30428 -11937 -30100
rect -11612 -30428 -11442 -30100
rect -11117 -30428 -10947 -30100
rect -10622 -30428 -10452 -30100
rect -10127 -30428 -9957 -30100
rect -9632 -30428 -9462 -30100
rect -9137 -30428 -8967 -30100
rect -8642 -30428 -8472 -30100
rect -8147 -30428 -7977 -30100
rect -7652 -30428 -7482 -30100
rect -7157 -30428 -6987 -30100
rect -6662 -30428 -6492 -30100
rect -6167 -30428 -5997 -30100
rect -5672 -30428 -5502 -30100
rect -5177 -30428 -5007 -30100
rect -4682 -30428 -4512 -30100
rect -4187 -30428 -4017 -30100
rect -3692 -30428 -3522 -30100
rect -3197 -30428 -3027 -30100
rect -2702 -30428 -2532 -30100
rect -2207 -30428 -2037 -30100
rect -1712 -30428 -1542 -30100
rect -1217 -30428 -1047 -30100
rect -722 -30428 -552 -30100
rect -227 -30428 -57 -30100
rect 268 -30428 438 -30100
rect 763 -30428 933 -30100
rect 1258 -30428 1428 -30100
rect 1753 -30428 1923 -30100
rect 2248 -30428 2418 -30100
rect 2743 -30428 2913 -30100
rect 3238 -30428 3408 -30100
rect 3733 -30428 3903 -30100
rect 4228 -30428 4398 -30100
rect 4723 -30428 4893 -30100
rect 5218 -30428 5388 -30100
rect 5713 -30428 5883 -30100
rect 6208 -30428 6378 -30100
rect 6703 -30428 6873 -30100
rect 7198 -30428 7368 -30100
rect 7693 -30428 7863 -30100
rect 8188 -30428 8358 -30100
rect 8683 -30428 8853 -30100
rect 9178 -30428 9348 -30100
rect 9673 -30428 9843 -30100
rect 10168 -30428 10338 -30100
rect 10663 -30428 10833 -30100
rect 11158 -30428 11328 -30100
rect 11653 -30428 11823 -30100
rect 12148 -30428 12318 -30100
rect 12643 -30428 12813 -30100
rect 13138 -30428 13308 -30100
rect 13633 -30428 13803 -30100
rect 14128 -30428 14298 -30100
rect 14623 -30428 14793 -30100
rect 15118 -30428 15288 -30100
rect 15613 -30428 15783 -30100
rect 16108 -30428 16278 -30100
rect 16603 -30428 16773 -30100
rect 17098 -30428 17268 -30100
rect 17593 -30428 17763 -30100
rect 18088 -30428 18258 -30100
rect 18583 -30428 18753 -30100
rect 19078 -30428 19248 -30100
rect 19573 -30428 19743 -30100
rect 20068 -30428 20238 -30100
rect 20563 -30428 20733 -30100
rect 21058 -30428 21228 -30100
rect 21553 -30428 21723 -30100
rect 22048 -30428 22218 -30100
rect 22543 -30428 22713 -30100
rect 23038 -30428 23208 -30100
rect 23533 -30428 23703 -30100
rect 24028 -30428 24198 -30100
rect 24523 -30428 24693 -30100
rect 25018 -30428 25188 -30100
rect 25513 -30428 25683 -30100
rect 26008 -30428 26178 -30100
rect 26503 -30428 26673 -30100
rect 26998 -30428 27168 -30100
rect 27493 -30428 27663 -30100
rect 27988 -30428 28158 -30100
rect 28483 -30428 28653 -30100
rect 28978 -30428 29148 -30100
rect 29473 -30428 29643 -30100
rect 29968 -30428 30138 -30100
rect 30463 -30428 30633 -30100
rect 30958 -30428 31128 -30100
rect 31453 -30428 31623 -30100
rect 31948 -30428 32118 -30100
rect 32443 -30428 32613 -30100
rect 32938 -30428 33108 -30100
rect 33433 -30428 33603 -30100
rect 33928 -30428 34098 -30100
rect 34423 -30428 34593 -30100
rect 34918 -30428 35088 -30100
rect 35413 -30428 35583 -30100
rect 35908 -30428 36078 -30100
rect 36403 -30428 36573 -30100
rect 36898 -30428 37068 -30100
rect 37393 -30428 37563 -30100
rect 37888 -30428 38058 -30100
rect 38383 -30428 38553 -30100
rect 38878 -30428 39048 -30100
rect 39373 -30428 39543 -30100
rect 39868 -30428 40038 -30100
rect 40363 -30428 40533 -30100
rect 40858 -30428 41028 -30100
rect 41353 -30428 41523 -30100
rect 41848 -30428 42018 -30100
rect 42343 -30428 42513 -30100
rect 42838 -30428 43008 -30100
rect 43333 -30428 43503 -30100
rect 43828 -30428 43998 -30100
rect 44323 -30428 44493 -30100
rect 44818 -30428 44988 -30100
rect 45313 -30428 45483 -30100
rect 45808 -30428 45978 -30100
rect 46303 -30428 46473 -30100
rect 46798 -30428 46968 -30100
rect 47293 -30428 47463 -30100
rect 47788 -30428 47958 -30100
rect 48283 -30428 48453 -30100
rect 48778 -30428 48948 -30100
rect 49273 -30428 49443 -30100
rect 49768 -30428 49938 -30100
rect 50263 -30428 50433 -30100
rect 50758 -30428 50928 -30100
rect 51253 -30428 51423 -30100
rect 51748 -30428 51918 -30100
rect 52243 -30428 52413 -30100
rect 52738 -30428 52908 -30100
rect 53233 -30428 53403 -30100
rect 53728 -30428 53898 -30100
rect 54223 -30320 54839 -30100
rect 54223 -30428 54840 -30320
rect -55858 -30576 54840 -30428
rect -55858 -30904 -55497 -30576
rect -55172 -30904 -55002 -30576
rect -54677 -30904 -54507 -30576
rect -54182 -30904 -54012 -30576
rect -53687 -30904 -53517 -30576
rect -53192 -30904 -53022 -30576
rect -52697 -30904 -52527 -30576
rect -52202 -30904 -52032 -30576
rect -51707 -30904 -51537 -30576
rect -51212 -30904 -51042 -30576
rect -50717 -30904 -50547 -30576
rect -50222 -30904 -50052 -30576
rect -49727 -30904 -49557 -30576
rect -49232 -30904 -49062 -30576
rect -48737 -30904 -48567 -30576
rect -48242 -30904 -48072 -30576
rect -47747 -30904 -47577 -30576
rect -47252 -30904 -47082 -30576
rect -46757 -30904 -46587 -30576
rect -46262 -30904 -46092 -30576
rect -45767 -30904 -45597 -30576
rect -45272 -30904 -45102 -30576
rect -44777 -30904 -44607 -30576
rect -44282 -30904 -44112 -30576
rect -43787 -30904 -43617 -30576
rect -43292 -30904 -43122 -30576
rect -42797 -30904 -42627 -30576
rect -42302 -30904 -42132 -30576
rect -41807 -30904 -41637 -30576
rect -41312 -30904 -41142 -30576
rect -40817 -30904 -40647 -30576
rect -40322 -30904 -40152 -30576
rect -39827 -30904 -39657 -30576
rect -39332 -30904 -39162 -30576
rect -38837 -30904 -38667 -30576
rect -38342 -30904 -38172 -30576
rect -37847 -30904 -37677 -30576
rect -37352 -30904 -37182 -30576
rect -36857 -30904 -36687 -30576
rect -36362 -30904 -36192 -30576
rect -35867 -30904 -35697 -30576
rect -35372 -30904 -35202 -30576
rect -34877 -30904 -34707 -30576
rect -34382 -30904 -34212 -30576
rect -33887 -30904 -33717 -30576
rect -33392 -30904 -33222 -30576
rect -32897 -30904 -32727 -30576
rect -32402 -30904 -32232 -30576
rect -31907 -30904 -31737 -30576
rect -31412 -30904 -31242 -30576
rect -30917 -30904 -30747 -30576
rect -30422 -30904 -30252 -30576
rect -29927 -30904 -29757 -30576
rect -29432 -30904 -29262 -30576
rect -28937 -30904 -28767 -30576
rect -28442 -30904 -28272 -30576
rect -27947 -30904 -27777 -30576
rect -27452 -30904 -27282 -30576
rect -26957 -30904 -26787 -30576
rect -26462 -30904 -26292 -30576
rect -25967 -30904 -25797 -30576
rect -25472 -30904 -25302 -30576
rect -24977 -30904 -24807 -30576
rect -24482 -30904 -24312 -30576
rect -23987 -30904 -23817 -30576
rect -23492 -30904 -23322 -30576
rect -22997 -30904 -22827 -30576
rect -22502 -30904 -22332 -30576
rect -22007 -30904 -21837 -30576
rect -21512 -30904 -21342 -30576
rect -21017 -30904 -20847 -30576
rect -20522 -30904 -20352 -30576
rect -20027 -30904 -19857 -30576
rect -19532 -30904 -19362 -30576
rect -19037 -30904 -18867 -30576
rect -18542 -30904 -18372 -30576
rect -18047 -30904 -17877 -30576
rect -17552 -30904 -17382 -30576
rect -17057 -30904 -16887 -30576
rect -16562 -30904 -16392 -30576
rect -16067 -30904 -15897 -30576
rect -15572 -30904 -15402 -30576
rect -15077 -30904 -14907 -30576
rect -14582 -30904 -14412 -30576
rect -14087 -30904 -13917 -30576
rect -13592 -30904 -13422 -30576
rect -13097 -30904 -12927 -30576
rect -12602 -30904 -12432 -30576
rect -12107 -30904 -11937 -30576
rect -11612 -30904 -11442 -30576
rect -11117 -30904 -10947 -30576
rect -10622 -30904 -10452 -30576
rect -10127 -30904 -9957 -30576
rect -9632 -30904 -9462 -30576
rect -9137 -30904 -8967 -30576
rect -8642 -30904 -8472 -30576
rect -8147 -30904 -7977 -30576
rect -7652 -30904 -7482 -30576
rect -7157 -30904 -6987 -30576
rect -6662 -30904 -6492 -30576
rect -6167 -30904 -5997 -30576
rect -5672 -30904 -5502 -30576
rect -5177 -30904 -5007 -30576
rect -4682 -30904 -4512 -30576
rect -4187 -30904 -4017 -30576
rect -3692 -30904 -3522 -30576
rect -3197 -30904 -3027 -30576
rect -2702 -30904 -2532 -30576
rect -2207 -30904 -2037 -30576
rect -1712 -30904 -1542 -30576
rect -1217 -30904 -1047 -30576
rect -722 -30904 -552 -30576
rect -227 -30904 -57 -30576
rect 268 -30904 438 -30576
rect 763 -30904 933 -30576
rect 1258 -30904 1428 -30576
rect 1753 -30904 1923 -30576
rect 2248 -30904 2418 -30576
rect 2743 -30904 2913 -30576
rect 3238 -30904 3408 -30576
rect 3733 -30904 3903 -30576
rect 4228 -30904 4398 -30576
rect 4723 -30904 4893 -30576
rect 5218 -30904 5388 -30576
rect 5713 -30904 5883 -30576
rect 6208 -30904 6378 -30576
rect 6703 -30904 6873 -30576
rect 7198 -30904 7368 -30576
rect 7693 -30904 7863 -30576
rect 8188 -30904 8358 -30576
rect 8683 -30904 8853 -30576
rect 9178 -30904 9348 -30576
rect 9673 -30904 9843 -30576
rect 10168 -30904 10338 -30576
rect 10663 -30904 10833 -30576
rect 11158 -30904 11328 -30576
rect 11653 -30904 11823 -30576
rect 12148 -30904 12318 -30576
rect 12643 -30904 12813 -30576
rect 13138 -30904 13308 -30576
rect 13633 -30904 13803 -30576
rect 14128 -30904 14298 -30576
rect 14623 -30904 14793 -30576
rect 15118 -30904 15288 -30576
rect 15613 -30904 15783 -30576
rect 16108 -30904 16278 -30576
rect 16603 -30904 16773 -30576
rect 17098 -30904 17268 -30576
rect 17593 -30904 17763 -30576
rect 18088 -30904 18258 -30576
rect 18583 -30904 18753 -30576
rect 19078 -30904 19248 -30576
rect 19573 -30904 19743 -30576
rect 20068 -30904 20238 -30576
rect 20563 -30904 20733 -30576
rect 21058 -30904 21228 -30576
rect 21553 -30904 21723 -30576
rect 22048 -30904 22218 -30576
rect 22543 -30904 22713 -30576
rect 23038 -30904 23208 -30576
rect 23533 -30904 23703 -30576
rect 24028 -30904 24198 -30576
rect 24523 -30904 24693 -30576
rect 25018 -30904 25188 -30576
rect 25513 -30904 25683 -30576
rect 26008 -30904 26178 -30576
rect 26503 -30904 26673 -30576
rect 26998 -30904 27168 -30576
rect 27493 -30904 27663 -30576
rect 27988 -30904 28158 -30576
rect 28483 -30904 28653 -30576
rect 28978 -30904 29148 -30576
rect 29473 -30904 29643 -30576
rect 29968 -30904 30138 -30576
rect 30463 -30904 30633 -30576
rect 30958 -30904 31128 -30576
rect 31453 -30904 31623 -30576
rect 31948 -30904 32118 -30576
rect 32443 -30904 32613 -30576
rect 32938 -30904 33108 -30576
rect 33433 -30904 33603 -30576
rect 33928 -30904 34098 -30576
rect 34423 -30904 34593 -30576
rect 34918 -30904 35088 -30576
rect 35413 -30904 35583 -30576
rect 35908 -30904 36078 -30576
rect 36403 -30904 36573 -30576
rect 36898 -30904 37068 -30576
rect 37393 -30904 37563 -30576
rect 37888 -30904 38058 -30576
rect 38383 -30904 38553 -30576
rect 38878 -30904 39048 -30576
rect 39373 -30904 39543 -30576
rect 39868 -30904 40038 -30576
rect 40363 -30904 40533 -30576
rect 40858 -30904 41028 -30576
rect 41353 -30904 41523 -30576
rect 41848 -30904 42018 -30576
rect 42343 -30904 42513 -30576
rect 42838 -30904 43008 -30576
rect 43333 -30904 43503 -30576
rect 43828 -30904 43998 -30576
rect 44323 -30904 44493 -30576
rect 44818 -30904 44988 -30576
rect 45313 -30904 45483 -30576
rect 45808 -30904 45978 -30576
rect 46303 -30904 46473 -30576
rect 46798 -30904 46968 -30576
rect 47293 -30904 47463 -30576
rect 47788 -30904 47958 -30576
rect 48283 -30904 48453 -30576
rect 48778 -30904 48948 -30576
rect 49273 -30904 49443 -30576
rect 49768 -30904 49938 -30576
rect 50263 -30904 50433 -30576
rect 50758 -30904 50928 -30576
rect 51253 -30904 51423 -30576
rect 51748 -30904 51918 -30576
rect 52243 -30904 52413 -30576
rect 52738 -30904 52908 -30576
rect 53233 -30904 53403 -30576
rect 53728 -30904 53898 -30576
rect 54223 -30904 54840 -30576
rect -55858 -31052 54840 -30904
rect -55858 -31380 -55497 -31052
rect -55172 -31380 -55002 -31052
rect -54677 -31380 -54507 -31052
rect -54182 -31380 -54012 -31052
rect -53687 -31380 -53517 -31052
rect -53192 -31380 -53022 -31052
rect -52697 -31380 -52527 -31052
rect -52202 -31380 -52032 -31052
rect -51707 -31380 -51537 -31052
rect -51212 -31380 -51042 -31052
rect -50717 -31380 -50547 -31052
rect -50222 -31380 -50052 -31052
rect -49727 -31380 -49557 -31052
rect -49232 -31380 -49062 -31052
rect -48737 -31380 -48567 -31052
rect -48242 -31380 -48072 -31052
rect -47747 -31380 -47577 -31052
rect -47252 -31380 -47082 -31052
rect -46757 -31380 -46587 -31052
rect -46262 -31380 -46092 -31052
rect -45767 -31380 -45597 -31052
rect -45272 -31380 -45102 -31052
rect -44777 -31380 -44607 -31052
rect -44282 -31380 -44112 -31052
rect -43787 -31380 -43617 -31052
rect -43292 -31380 -43122 -31052
rect -42797 -31380 -42627 -31052
rect -42302 -31380 -42132 -31052
rect -41807 -31380 -41637 -31052
rect -41312 -31380 -41142 -31052
rect -40817 -31380 -40647 -31052
rect -40322 -31380 -40152 -31052
rect -39827 -31380 -39657 -31052
rect -39332 -31380 -39162 -31052
rect -38837 -31380 -38667 -31052
rect -38342 -31380 -38172 -31052
rect -37847 -31380 -37677 -31052
rect -37352 -31380 -37182 -31052
rect -36857 -31380 -36687 -31052
rect -36362 -31380 -36192 -31052
rect -35867 -31380 -35697 -31052
rect -35372 -31380 -35202 -31052
rect -34877 -31380 -34707 -31052
rect -34382 -31380 -34212 -31052
rect -33887 -31380 -33717 -31052
rect -33392 -31380 -33222 -31052
rect -32897 -31380 -32727 -31052
rect -32402 -31380 -32232 -31052
rect -31907 -31380 -31737 -31052
rect -31412 -31380 -31242 -31052
rect -30917 -31380 -30747 -31052
rect -30422 -31380 -30252 -31052
rect -29927 -31380 -29757 -31052
rect -29432 -31380 -29262 -31052
rect -28937 -31380 -28767 -31052
rect -28442 -31380 -28272 -31052
rect -27947 -31380 -27777 -31052
rect -27452 -31380 -27282 -31052
rect -26957 -31380 -26787 -31052
rect -26462 -31380 -26292 -31052
rect -25967 -31380 -25797 -31052
rect -25472 -31380 -25302 -31052
rect -24977 -31380 -24807 -31052
rect -24482 -31380 -24312 -31052
rect -23987 -31380 -23817 -31052
rect -23492 -31380 -23322 -31052
rect -22997 -31380 -22827 -31052
rect -22502 -31380 -22332 -31052
rect -22007 -31380 -21837 -31052
rect -21512 -31380 -21342 -31052
rect -21017 -31380 -20847 -31052
rect -20522 -31380 -20352 -31052
rect -20027 -31380 -19857 -31052
rect -19532 -31380 -19362 -31052
rect -19037 -31380 -18867 -31052
rect -18542 -31380 -18372 -31052
rect -18047 -31380 -17877 -31052
rect -17552 -31380 -17382 -31052
rect -17057 -31380 -16887 -31052
rect -16562 -31380 -16392 -31052
rect -16067 -31380 -15897 -31052
rect -15572 -31380 -15402 -31052
rect -15077 -31380 -14907 -31052
rect -14582 -31380 -14412 -31052
rect -14087 -31380 -13917 -31052
rect -13592 -31380 -13422 -31052
rect -13097 -31380 -12927 -31052
rect -12602 -31380 -12432 -31052
rect -12107 -31380 -11937 -31052
rect -11612 -31380 -11442 -31052
rect -11117 -31380 -10947 -31052
rect -10622 -31380 -10452 -31052
rect -10127 -31380 -9957 -31052
rect -9632 -31380 -9462 -31052
rect -9137 -31380 -8967 -31052
rect -8642 -31380 -8472 -31052
rect -8147 -31380 -7977 -31052
rect -7652 -31380 -7482 -31052
rect -7157 -31380 -6987 -31052
rect -6662 -31380 -6492 -31052
rect -6167 -31380 -5997 -31052
rect -5672 -31380 -5502 -31052
rect -5177 -31380 -5007 -31052
rect -4682 -31380 -4512 -31052
rect -4187 -31380 -4017 -31052
rect -3692 -31380 -3522 -31052
rect -3197 -31380 -3027 -31052
rect -2702 -31380 -2532 -31052
rect -2207 -31380 -2037 -31052
rect -1712 -31380 -1542 -31052
rect -1217 -31380 -1047 -31052
rect -722 -31380 -552 -31052
rect -227 -31380 -57 -31052
rect 268 -31380 438 -31052
rect 763 -31380 933 -31052
rect 1258 -31380 1428 -31052
rect 1753 -31380 1923 -31052
rect 2248 -31380 2418 -31052
rect 2743 -31380 2913 -31052
rect 3238 -31380 3408 -31052
rect 3733 -31380 3903 -31052
rect 4228 -31380 4398 -31052
rect 4723 -31380 4893 -31052
rect 5218 -31380 5388 -31052
rect 5713 -31380 5883 -31052
rect 6208 -31380 6378 -31052
rect 6703 -31380 6873 -31052
rect 7198 -31380 7368 -31052
rect 7693 -31380 7863 -31052
rect 8188 -31380 8358 -31052
rect 8683 -31380 8853 -31052
rect 9178 -31380 9348 -31052
rect 9673 -31380 9843 -31052
rect 10168 -31380 10338 -31052
rect 10663 -31380 10833 -31052
rect 11158 -31380 11328 -31052
rect 11653 -31380 11823 -31052
rect 12148 -31380 12318 -31052
rect 12643 -31380 12813 -31052
rect 13138 -31380 13308 -31052
rect 13633 -31380 13803 -31052
rect 14128 -31380 14298 -31052
rect 14623 -31380 14793 -31052
rect 15118 -31380 15288 -31052
rect 15613 -31380 15783 -31052
rect 16108 -31380 16278 -31052
rect 16603 -31380 16773 -31052
rect 17098 -31380 17268 -31052
rect 17593 -31380 17763 -31052
rect 18088 -31380 18258 -31052
rect 18583 -31380 18753 -31052
rect 19078 -31380 19248 -31052
rect 19573 -31380 19743 -31052
rect 20068 -31380 20238 -31052
rect 20563 -31380 20733 -31052
rect 21058 -31380 21228 -31052
rect 21553 -31380 21723 -31052
rect 22048 -31380 22218 -31052
rect 22543 -31380 22713 -31052
rect 23038 -31380 23208 -31052
rect 23533 -31380 23703 -31052
rect 24028 -31380 24198 -31052
rect 24523 -31380 24693 -31052
rect 25018 -31380 25188 -31052
rect 25513 -31380 25683 -31052
rect 26008 -31380 26178 -31052
rect 26503 -31380 26673 -31052
rect 26998 -31380 27168 -31052
rect 27493 -31380 27663 -31052
rect 27988 -31380 28158 -31052
rect 28483 -31380 28653 -31052
rect 28978 -31380 29148 -31052
rect 29473 -31380 29643 -31052
rect 29968 -31380 30138 -31052
rect 30463 -31380 30633 -31052
rect 30958 -31380 31128 -31052
rect 31453 -31380 31623 -31052
rect 31948 -31380 32118 -31052
rect 32443 -31380 32613 -31052
rect 32938 -31380 33108 -31052
rect 33433 -31380 33603 -31052
rect 33928 -31380 34098 -31052
rect 34423 -31380 34593 -31052
rect 34918 -31380 35088 -31052
rect 35413 -31380 35583 -31052
rect 35908 -31380 36078 -31052
rect 36403 -31380 36573 -31052
rect 36898 -31380 37068 -31052
rect 37393 -31380 37563 -31052
rect 37888 -31380 38058 -31052
rect 38383 -31380 38553 -31052
rect 38878 -31380 39048 -31052
rect 39373 -31380 39543 -31052
rect 39868 -31380 40038 -31052
rect 40363 -31380 40533 -31052
rect 40858 -31380 41028 -31052
rect 41353 -31380 41523 -31052
rect 41848 -31380 42018 -31052
rect 42343 -31380 42513 -31052
rect 42838 -31380 43008 -31052
rect 43333 -31380 43503 -31052
rect 43828 -31380 43998 -31052
rect 44323 -31380 44493 -31052
rect 44818 -31380 44988 -31052
rect 45313 -31380 45483 -31052
rect 45808 -31380 45978 -31052
rect 46303 -31380 46473 -31052
rect 46798 -31380 46968 -31052
rect 47293 -31380 47463 -31052
rect 47788 -31380 47958 -31052
rect 48283 -31380 48453 -31052
rect 48778 -31380 48948 -31052
rect 49273 -31380 49443 -31052
rect 49768 -31380 49938 -31052
rect 50263 -31380 50433 -31052
rect 50758 -31380 50928 -31052
rect 51253 -31380 51423 -31052
rect 51748 -31380 51918 -31052
rect 52243 -31380 52413 -31052
rect 52738 -31380 52908 -31052
rect 53233 -31380 53403 -31052
rect 53728 -31380 53898 -31052
rect 54223 -31380 54840 -31052
rect -55858 -31528 54840 -31380
rect -55858 -31856 -55497 -31528
rect -55172 -31856 -55002 -31528
rect -54677 -31856 -54507 -31528
rect -54182 -31856 -54012 -31528
rect -53687 -31856 -53517 -31528
rect -53192 -31856 -53022 -31528
rect -52697 -31856 -52527 -31528
rect -52202 -31856 -52032 -31528
rect -51707 -31856 -51537 -31528
rect -51212 -31856 -51042 -31528
rect -50717 -31856 -50547 -31528
rect -50222 -31856 -50052 -31528
rect -49727 -31856 -49557 -31528
rect -49232 -31856 -49062 -31528
rect -48737 -31856 -48567 -31528
rect -48242 -31856 -48072 -31528
rect -47747 -31856 -47577 -31528
rect -47252 -31856 -47082 -31528
rect -46757 -31856 -46587 -31528
rect -46262 -31856 -46092 -31528
rect -45767 -31856 -45597 -31528
rect -45272 -31856 -45102 -31528
rect -44777 -31856 -44607 -31528
rect -44282 -31856 -44112 -31528
rect -43787 -31856 -43617 -31528
rect -43292 -31856 -43122 -31528
rect -42797 -31856 -42627 -31528
rect -42302 -31856 -42132 -31528
rect -41807 -31856 -41637 -31528
rect -41312 -31856 -41142 -31528
rect -40817 -31856 -40647 -31528
rect -40322 -31856 -40152 -31528
rect -39827 -31856 -39657 -31528
rect -39332 -31856 -39162 -31528
rect -38837 -31856 -38667 -31528
rect -38342 -31856 -38172 -31528
rect -37847 -31856 -37677 -31528
rect -37352 -31856 -37182 -31528
rect -36857 -31856 -36687 -31528
rect -36362 -31856 -36192 -31528
rect -35867 -31856 -35697 -31528
rect -35372 -31856 -35202 -31528
rect -34877 -31856 -34707 -31528
rect -34382 -31856 -34212 -31528
rect -33887 -31856 -33717 -31528
rect -33392 -31856 -33222 -31528
rect -32897 -31856 -32727 -31528
rect -32402 -31856 -32232 -31528
rect -31907 -31856 -31737 -31528
rect -31412 -31856 -31242 -31528
rect -30917 -31856 -30747 -31528
rect -30422 -31856 -30252 -31528
rect -29927 -31856 -29757 -31528
rect -29432 -31856 -29262 -31528
rect -28937 -31856 -28767 -31528
rect -28442 -31856 -28272 -31528
rect -27947 -31856 -27777 -31528
rect -27452 -31856 -27282 -31528
rect -26957 -31856 -26787 -31528
rect -26462 -31856 -26292 -31528
rect -25967 -31856 -25797 -31528
rect -25472 -31856 -25302 -31528
rect -24977 -31856 -24807 -31528
rect -24482 -31856 -24312 -31528
rect -23987 -31856 -23817 -31528
rect -23492 -31856 -23322 -31528
rect -22997 -31856 -22827 -31528
rect -22502 -31856 -22332 -31528
rect -22007 -31856 -21837 -31528
rect -21512 -31856 -21342 -31528
rect -21017 -31856 -20847 -31528
rect -20522 -31856 -20352 -31528
rect -20027 -31856 -19857 -31528
rect -19532 -31856 -19362 -31528
rect -19037 -31856 -18867 -31528
rect -18542 -31856 -18372 -31528
rect -18047 -31856 -17877 -31528
rect -17552 -31856 -17382 -31528
rect -17057 -31856 -16887 -31528
rect -16562 -31856 -16392 -31528
rect -16067 -31856 -15897 -31528
rect -15572 -31856 -15402 -31528
rect -15077 -31856 -14907 -31528
rect -14582 -31856 -14412 -31528
rect -14087 -31856 -13917 -31528
rect -13592 -31856 -13422 -31528
rect -13097 -31856 -12927 -31528
rect -12602 -31856 -12432 -31528
rect -12107 -31856 -11937 -31528
rect -11612 -31856 -11442 -31528
rect -11117 -31856 -10947 -31528
rect -10622 -31856 -10452 -31528
rect -10127 -31856 -9957 -31528
rect -9632 -31856 -9462 -31528
rect -9137 -31856 -8967 -31528
rect -8642 -31856 -8472 -31528
rect -8147 -31856 -7977 -31528
rect -7652 -31856 -7482 -31528
rect -7157 -31856 -6987 -31528
rect -6662 -31856 -6492 -31528
rect -6167 -31856 -5997 -31528
rect -5672 -31856 -5502 -31528
rect -5177 -31856 -5007 -31528
rect -4682 -31856 -4512 -31528
rect -4187 -31856 -4017 -31528
rect -3692 -31856 -3522 -31528
rect -3197 -31856 -3027 -31528
rect -2702 -31856 -2532 -31528
rect -2207 -31856 -2037 -31528
rect -1712 -31856 -1542 -31528
rect -1217 -31856 -1047 -31528
rect -722 -31856 -552 -31528
rect -227 -31856 -57 -31528
rect 268 -31856 438 -31528
rect 763 -31856 933 -31528
rect 1258 -31856 1428 -31528
rect 1753 -31856 1923 -31528
rect 2248 -31856 2418 -31528
rect 2743 -31856 2913 -31528
rect 3238 -31856 3408 -31528
rect 3733 -31856 3903 -31528
rect 4228 -31856 4398 -31528
rect 4723 -31856 4893 -31528
rect 5218 -31856 5388 -31528
rect 5713 -31856 5883 -31528
rect 6208 -31856 6378 -31528
rect 6703 -31856 6873 -31528
rect 7198 -31856 7368 -31528
rect 7693 -31856 7863 -31528
rect 8188 -31856 8358 -31528
rect 8683 -31856 8853 -31528
rect 9178 -31856 9348 -31528
rect 9673 -31856 9843 -31528
rect 10168 -31856 10338 -31528
rect 10663 -31856 10833 -31528
rect 11158 -31856 11328 -31528
rect 11653 -31856 11823 -31528
rect 12148 -31856 12318 -31528
rect 12643 -31856 12813 -31528
rect 13138 -31856 13308 -31528
rect 13633 -31856 13803 -31528
rect 14128 -31856 14298 -31528
rect 14623 -31856 14793 -31528
rect 15118 -31856 15288 -31528
rect 15613 -31856 15783 -31528
rect 16108 -31856 16278 -31528
rect 16603 -31856 16773 -31528
rect 17098 -31856 17268 -31528
rect 17593 -31856 17763 -31528
rect 18088 -31856 18258 -31528
rect 18583 -31856 18753 -31528
rect 19078 -31856 19248 -31528
rect 19573 -31856 19743 -31528
rect 20068 -31856 20238 -31528
rect 20563 -31856 20733 -31528
rect 21058 -31856 21228 -31528
rect 21553 -31856 21723 -31528
rect 22048 -31856 22218 -31528
rect 22543 -31856 22713 -31528
rect 23038 -31856 23208 -31528
rect 23533 -31856 23703 -31528
rect 24028 -31856 24198 -31528
rect 24523 -31856 24693 -31528
rect 25018 -31856 25188 -31528
rect 25513 -31856 25683 -31528
rect 26008 -31856 26178 -31528
rect 26503 -31856 26673 -31528
rect 26998 -31856 27168 -31528
rect 27493 -31856 27663 -31528
rect 27988 -31856 28158 -31528
rect 28483 -31856 28653 -31528
rect 28978 -31856 29148 -31528
rect 29473 -31856 29643 -31528
rect 29968 -31856 30138 -31528
rect 30463 -31856 30633 -31528
rect 30958 -31856 31128 -31528
rect 31453 -31856 31623 -31528
rect 31948 -31856 32118 -31528
rect 32443 -31856 32613 -31528
rect 32938 -31856 33108 -31528
rect 33433 -31856 33603 -31528
rect 33928 -31856 34098 -31528
rect 34423 -31856 34593 -31528
rect 34918 -31856 35088 -31528
rect 35413 -31856 35583 -31528
rect 35908 -31856 36078 -31528
rect 36403 -31856 36573 -31528
rect 36898 -31856 37068 -31528
rect 37393 -31856 37563 -31528
rect 37888 -31856 38058 -31528
rect 38383 -31856 38553 -31528
rect 38878 -31856 39048 -31528
rect 39373 -31856 39543 -31528
rect 39868 -31856 40038 -31528
rect 40363 -31856 40533 -31528
rect 40858 -31856 41028 -31528
rect 41353 -31856 41523 -31528
rect 41848 -31856 42018 -31528
rect 42343 -31856 42513 -31528
rect 42838 -31856 43008 -31528
rect 43333 -31856 43503 -31528
rect 43828 -31856 43998 -31528
rect 44323 -31856 44493 -31528
rect 44818 -31856 44988 -31528
rect 45313 -31856 45483 -31528
rect 45808 -31856 45978 -31528
rect 46303 -31856 46473 -31528
rect 46798 -31856 46968 -31528
rect 47293 -31856 47463 -31528
rect 47788 -31856 47958 -31528
rect 48283 -31856 48453 -31528
rect 48778 -31856 48948 -31528
rect 49273 -31856 49443 -31528
rect 49768 -31856 49938 -31528
rect 50263 -31856 50433 -31528
rect 50758 -31856 50928 -31528
rect 51253 -31856 51423 -31528
rect 51748 -31856 51918 -31528
rect 52243 -31856 52413 -31528
rect 52738 -31856 52908 -31528
rect 53233 -31856 53403 -31528
rect 53728 -31856 53898 -31528
rect 54223 -31856 54840 -31528
rect -55858 -32147 54840 -31856
rect -55274 -32154 -53816 -32147
<< via1 >>
rect -6106 24257 -6013 24339
rect -5922 24270 -5829 24352
rect -6113 24074 -6020 24156
rect -5932 24087 -5839 24169
rect 198 24007 250 24066
rect 307 24007 359 24066
rect 418 24008 470 24067
rect 530 24011 582 24070
rect 1230 24007 1282 24066
rect 1339 24007 1391 24066
rect 1450 24008 1502 24067
rect 1562 24011 1614 24070
rect 26160 24017 26233 24087
rect 26300 24018 26373 24088
rect 26429 24026 26502 24096
rect -6128 23897 -6035 23979
rect -5934 23902 -5841 23984
rect 199 23896 251 23955
rect 308 23896 360 23955
rect 420 23896 472 23955
rect 529 23897 581 23956
rect 1231 23896 1283 23955
rect 1340 23896 1392 23955
rect 1452 23896 1504 23955
rect 1561 23897 1613 23956
rect 24725 23926 24798 23996
rect 24864 23932 24937 24002
rect 25018 23939 25091 24009
rect 27546 24007 27619 24077
rect 27699 24012 27772 24082
rect 27850 24014 27923 24084
rect 48564 24081 48616 24134
rect 48680 24084 48735 24138
rect 48787 24086 48842 24140
rect 48560 23970 48612 24023
rect 48679 23978 48731 24031
rect 48786 23974 48838 24027
rect 26157 23888 26230 23958
rect 26302 23889 26375 23959
rect 26437 23892 26510 23962
rect 27544 23880 27617 23950
rect 27699 23889 27772 23959
rect 27853 23891 27926 23961
rect 48615 23857 48677 23912
rect 48744 23864 48806 23919
rect 22923 23308 23021 23415
rect 23184 23075 23282 23182
rect 23521 22774 23619 22881
rect -4271 22403 -4129 22512
rect -3590 22197 -3536 22319
rect 4621 21969 4724 22091
rect 4808 21969 4911 22091
rect 5008 21970 5111 22092
rect 4624 21770 4727 21892
rect 4814 21768 4917 21890
rect 5007 21770 5110 21892
rect 24736 19970 24809 20040
rect 24887 19973 24960 20043
rect 25037 19979 25110 20049
rect 26155 19989 26228 20059
rect 26302 19993 26375 20063
rect 26444 20001 26517 20071
rect 27557 19989 27630 20059
rect 27694 19993 27767 20063
rect 27836 20003 27909 20073
rect -6169 14782 -6108 14851
rect -6045 14785 -5984 14854
rect -6171 14654 -6110 14723
rect -6042 14659 -5981 14728
rect 56382 -327 56434 -275
rect 56501 -327 56553 -275
rect 56379 -433 56431 -381
rect 56496 -431 56548 -379
rect 47198 -1992 47271 -1923
rect 47373 -1998 47446 -1929
rect 47197 -2157 47270 -2088
rect 47370 -2160 47443 -2091
rect -8415 -2446 -8338 -2354
rect -2628 -2440 -2537 -2345
rect 224 -2652 341 -2535
rect 443 -2649 560 -2532
rect 221 -2837 338 -2720
rect 440 -2828 557 -2711
rect -6441 -3274 -6385 -3216
rect -6333 -3276 -6277 -3218
rect -4906 -3243 -4843 -3176
rect -2624 -3223 -2542 -3161
rect 49385 -4205 49451 -4143
rect 49506 -4201 49569 -4142
rect -5187 -4286 -5135 -4234
rect -3876 -4288 -3810 -4233
rect 49380 -4323 49446 -4261
rect 49514 -4315 49577 -4256
rect -5193 -5068 -5131 -5010
rect -5077 -5061 -5015 -5003
rect 5255 -5051 5326 -4981
rect -5193 -5185 -5131 -5127
rect -5075 -5185 -5013 -5127
rect 5253 -5191 5324 -5121
rect 56374 -5013 56426 -4961
rect 56493 -5013 56545 -4961
rect 56371 -5119 56423 -5067
rect 56488 -5117 56540 -5065
rect -6423 -5504 -6367 -5446
rect -6315 -5550 -6259 -5492
rect 5466 -5498 5531 -5427
rect -6423 -5620 -6367 -5562
rect 5468 -5633 5533 -5562
rect 47793 -6681 47871 -6601
rect 47971 -6684 48049 -6604
rect 47792 -6818 47870 -6738
rect 47966 -6816 48044 -6736
rect -7693 -7716 -7609 -7621
rect 3215 -7703 3304 -7636
rect -7836 -7825 -7752 -7730
rect 3214 -7822 3303 -7755
rect 218 -8275 270 -8216
rect 323 -8275 375 -8216
rect 437 -8274 489 -8215
rect 545 -8270 597 -8211
rect 1227 -8268 1279 -8209
rect 1346 -8267 1398 -8208
rect 1473 -8264 1525 -8205
rect 1584 -8262 1636 -8203
rect 55881 -9352 56139 -9255
rect -6009 -9553 -5941 -9492
rect 4110 -10238 4176 -10186
rect 4138 -10349 4233 -10297
rect 750 -11722 809 -11661
rect 882 -11720 941 -11659
rect 8337 -13682 8414 -13593
rect 8518 -13680 8595 -13591
rect 25459 -13649 25555 -13582
rect 8340 -13825 8417 -13736
rect 8518 -13825 8595 -13736
rect 25453 -13805 25552 -13706
rect 42760 -13683 42838 -13603
rect 42938 -13686 43016 -13606
rect 47809 -13655 47887 -13575
rect 47987 -13658 48065 -13578
rect 42759 -13820 42837 -13740
rect 42933 -13818 43011 -13738
rect 47808 -13792 47886 -13712
rect 47982 -13790 48060 -13710
rect 8340 -13986 8417 -13897
rect 8516 -13986 8593 -13897
rect 25452 -13972 25551 -13873
rect 49382 -14257 49460 -14203
rect 49513 -14255 49591 -14201
rect 49384 -14389 49453 -14313
rect 49516 -14384 49585 -14308
rect 49381 -14533 49450 -14457
rect 49514 -14528 49583 -14452
rect -6830 -14889 -6723 -14805
rect 49422 -14839 49506 -14761
rect 49618 -14833 49702 -14755
rect 49424 -14986 49508 -14908
rect 49616 -14978 49700 -14900
rect 13245 -15767 13319 -15685
rect 13391 -15771 13465 -15689
rect 13244 -15927 13318 -15845
rect 13396 -15914 13470 -15832
rect 13660 -16172 13742 -16096
rect 13815 -16168 13897 -16092
rect 13662 -16313 13744 -16237
rect 13813 -16304 13895 -16228
rect 49440 -16290 49580 -16120
rect -6045 -16517 -5991 -16463
rect -5923 -16517 -5869 -16463
rect 47214 -16554 47292 -16480
rect 47356 -16550 47434 -16476
rect 47224 -16692 47302 -16618
rect 47357 -16681 47435 -16607
rect 14391 -16868 14455 -16793
rect 14539 -16864 14603 -16789
rect 14669 -16864 14733 -16789
rect -10386 -17050 -10278 -16929
rect -10159 -17045 -10051 -16924
rect -10386 -17265 -10278 -17144
rect -10159 -17261 -10051 -17140
rect -8300 -17000 -8210 -16903
rect -8130 -16999 -8040 -16902
rect 14391 -17021 14455 -16946
rect 14537 -17018 14601 -16943
rect 14669 -17017 14733 -16942
rect -8300 -17167 -8210 -17070
rect -8130 -17164 -8040 -17067
rect 14391 -17182 14455 -17107
rect 14530 -17182 14594 -17107
rect 14669 -17182 14733 -17107
rect 43704 -17128 43788 -17006
rect -3210 -17676 -3022 -17518
rect 4113 -17682 4249 -17532
rect 15178 -18099 15340 -17976
rect 49672 -17087 49750 -17013
rect 49814 -17083 49892 -17009
rect 37209 -17492 37308 -17388
rect 49682 -17225 49760 -17151
rect 49815 -17214 49893 -17140
rect 48511 -17387 48563 -17334
rect 48622 -17385 48674 -17332
rect 48728 -17384 48780 -17331
rect 48846 -17385 48898 -17332
rect 43687 -17946 43839 -17879
rect -3731 -18245 -3599 -18136
rect 4591 -18262 4670 -18168
rect 4752 -18264 4831 -18170
rect 4918 -18261 4997 -18167
rect -3731 -18430 -3599 -18321
rect 5053 -18330 5121 -18236
rect 4593 -18426 4672 -18332
rect 4753 -18426 4832 -18332
rect 4919 -18426 4998 -18332
rect 29284 -18455 29359 -18381
rect 31466 -18546 31528 -18485
rect 49905 -18690 49979 -18633
rect 303 -18812 370 -18754
rect 444 -18810 511 -18752
rect 8344 -18796 8398 -18724
rect 8452 -18795 8508 -18723
rect 301 -18939 368 -18881
rect 445 -18933 512 -18875
rect 11747 -18796 11802 -18733
rect 38290 -18746 38343 -18693
rect 8375 -19081 8467 -18974
rect 42792 -19364 42860 -19292
rect 42935 -19362 43003 -19290
rect 54340 -19414 54392 -19361
rect 54444 -19412 54496 -19359
rect 42789 -19528 42857 -19456
rect 42933 -19529 43001 -19457
rect 7352 -19761 7439 -19753
rect 7352 -19830 7441 -19761
rect -3171 -20813 -3026 -20727
rect 5276 -20868 5347 -20807
rect 7091 -20878 7148 -20812
rect 8365 -20972 8457 -20913
rect 14892 -20737 14980 -20573
rect 15064 -20737 15152 -20573
rect 15936 -20638 15988 -20543
rect 16040 -20640 16092 -20545
rect 17299 -20598 17353 -20544
rect 17405 -20599 17459 -20545
rect 25572 -20632 25624 -20580
rect 26645 -20627 26723 -20554
rect 21142 -20815 21213 -20750
rect 22493 -20825 22553 -20753
rect 13712 -21350 13814 -21245
rect 7104 -21489 7163 -21417
rect -3084 -21667 -3009 -21572
rect -1789 -21861 -1734 -21808
rect 5753 -22022 5813 -21966
rect 8699 -22053 8770 -21984
rect 14157 -22090 14225 -22024
rect 26152 -22456 26205 -22396
rect 5909 -22558 5981 -22505
rect 7609 -22582 7664 -22524
rect 11730 -22580 11830 -22480
rect -3725 -22909 -3665 -22847
rect -3602 -22910 -3542 -22848
rect 5756 -22926 5813 -22871
rect 14516 -22918 14622 -22862
rect 38275 -22894 38353 -22811
rect 39032 -22895 39121 -22791
rect 7120 -23072 7191 -23012
rect 14445 -23061 14521 -22972
rect 14604 -23061 14680 -22972
rect 49907 -22989 49996 -22879
rect 50534 -22990 50623 -22880
rect -1488 -23447 -1429 -23387
rect 7611 -23476 7680 -23403
rect 6169 -23702 6238 -23650
rect 6171 -23807 6240 -23755
rect 10766 -23792 10818 -23692
rect -1635 -23959 -1579 -23897
rect 5895 -24141 5996 -24074
rect 8694 -24116 8777 -24041
rect 10918 -24138 11078 -24066
rect 764 -24387 866 -24273
rect 949 -24381 1051 -24267
rect 1128 -24379 1230 -24265
rect 4937 -24401 5039 -24287
rect 5131 -24393 5233 -24279
rect 5333 -24381 5435 -24267
rect 9210 -24364 9312 -24250
rect 9412 -24362 9514 -24248
rect 9605 -24362 9707 -24248
rect 10920 -24272 11070 -24205
rect 10919 -24395 11069 -24328
rect 12251 -24365 12319 -24275
rect 12403 -24358 12471 -24268
rect 12555 -24360 12623 -24270
rect 12715 -24358 12783 -24268
rect -6849 -24519 -6796 -24463
rect -6744 -24518 -6691 -24460
rect -1789 -24518 -1735 -24462
rect 20383 -24089 20444 -24021
rect 20505 -24085 20566 -24017
rect 21110 -24091 21171 -24023
rect 21244 -24088 21305 -24020
rect 21729 -24096 21790 -24028
rect 21843 -24097 21902 -24029
rect 28195 -24606 28352 -24445
rect -2630 -24740 -2570 -24670
rect 6180 -24750 6270 -24650
rect -1652 -24909 -1570 -24846
rect 4356 -24896 4413 -24837
rect -3075 -25069 -3017 -25016
rect 4546 -25085 4608 -25014
rect -27358 -26438 -27265 -26333
rect -27172 -26432 -27079 -26327
rect -26953 -26432 -26860 -26327
rect -24900 -26447 -24807 -26342
rect -24699 -26432 -24606 -26327
rect -24510 -26438 -24417 -26333
rect -22310 -26482 -22217 -26377
rect -22057 -26479 -21964 -26374
rect -19777 -26479 -19684 -26374
rect -19547 -26475 -19454 -26374
rect -17292 -26464 -17199 -26359
rect -17089 -26464 -16996 -26359
rect -16934 -26458 -16841 -26353
rect -14372 -26479 -14279 -26374
rect -14159 -26467 -14066 -26362
rect -13993 -26455 -13900 -26350
rect -11963 -26470 -11870 -26365
rect -11780 -26467 -11687 -26362
rect -11570 -26464 -11477 -26359
rect -27352 -26633 -27259 -26528
rect -27166 -26627 -27073 -26522
rect -26965 -26621 -26872 -26516
rect -24914 -26650 -24821 -26545
rect -24693 -26636 -24600 -26531
rect -24516 -26627 -24423 -26522
rect -22372 -26656 -22279 -26551
rect -22150 -26650 -22057 -26545
rect -21958 -26647 -21865 -26542
rect -19823 -26659 -19730 -26554
rect -19628 -26647 -19535 -26542
rect -19442 -26633 -19349 -26528
rect -17310 -26645 -17217 -26540
rect -17121 -26647 -17028 -26542
rect -16920 -26639 -16827 -26534
rect -14372 -26636 -14279 -26531
rect -14162 -26636 -14069 -26531
rect -13982 -26624 -13889 -26519
rect -11972 -26647 -11879 -26542
rect -11797 -26639 -11704 -26534
rect -11582 -26630 -11489 -26525
rect 32080 -25447 32192 -25334
rect 43698 -25445 43816 -25320
rect 44605 -25602 44659 -25539
rect 44715 -25603 44769 -25540
rect 33766 -25685 33819 -25631
rect 33889 -25685 33942 -25631
rect 35210 -25692 35263 -25638
rect 35352 -25689 35405 -25635
rect 36586 -25671 36639 -25617
rect 36703 -25672 36756 -25618
rect 37992 -25674 38045 -25620
rect 38117 -25672 38170 -25618
rect 45823 -25619 45877 -25556
rect 45954 -25619 46008 -25556
rect 46948 -25626 47002 -25563
rect 47077 -25619 47131 -25556
rect 47967 -25623 48021 -25560
rect 48100 -25620 48154 -25557
rect 49256 -25623 49310 -25560
rect 49394 -25622 49448 -25559
rect 6520 -25800 6590 -25730
rect 11330 -25800 11400 -25740
rect -8446 -27301 -8317 -27177
rect 56683 -27173 56771 -27103
rect 56846 -27171 56934 -27101
rect 56680 -27314 56768 -27244
rect 56840 -27309 56928 -27239
rect 38004 -29624 38064 -29583
rect 38125 -29624 38185 -29579
rect -27343 -29921 -27282 -29821
rect -27282 -29921 -27260 -29821
rect -27172 -29921 -27089 -29821
rect -26994 -29916 -26957 -29816
rect -26957 -29916 -26911 -29816
rect -24934 -29898 -24851 -29798
rect -24751 -29889 -24668 -29789
rect -24542 -29878 -24482 -29778
rect -24482 -29878 -24459 -29778
rect -22352 -29893 -22332 -29793
rect -22332 -29893 -22269 -29793
rect -22165 -29893 -22082 -29793
rect -21972 -29888 -21889 -29788
rect -19805 -29898 -19722 -29798
rect -19598 -29896 -19532 -29796
rect -19532 -29896 -19515 -29796
rect -19407 -29887 -19362 -29787
rect -19362 -29887 -19324 -29787
rect -17294 -29882 -17211 -29782
rect -17118 -29878 -17057 -29778
rect -17057 -29878 -17035 -29778
rect -16929 -29878 -16887 -29778
rect -16887 -29878 -16846 -29778
rect -14376 -29889 -14293 -29789
rect -14203 -29884 -14120 -29784
rect -14030 -29884 -13947 -29784
rect -11942 -29884 -11937 -29784
rect -11937 -29884 -11859 -29784
rect -11741 -29882 -11658 -29782
rect -11552 -29878 -11469 -29778
rect -6034 -29881 -5997 -29816
rect -5997 -29881 -5973 -29816
rect -5902 -29873 -5841 -29808
rect -6034 -29952 -5997 -29948
rect -5997 -29952 -5973 -29948
rect -5906 -29952 -5845 -29948
rect 750 -29952 763 -29882
rect 763 -29952 852 -29882
rect -27348 -30080 -27265 -30021
rect -27170 -30080 -27087 -30019
rect -26978 -30080 -26895 -30008
rect -24929 -30080 -24846 -29994
rect -24738 -30080 -24655 -29980
rect -24537 -30074 -24454 -29974
rect -22358 -30076 -22275 -29976
rect -22171 -30076 -22088 -29976
rect -21978 -30071 -21895 -29971
rect -19821 -30080 -19738 -29992
rect -19603 -30076 -19520 -29976
rect -19411 -30074 -19328 -29974
rect -17303 -30080 -17220 -29985
rect -17116 -30080 -17033 -29987
rect -16918 -30080 -16835 -29985
rect -14383 -30080 -14300 -29980
rect -14203 -30074 -14120 -29974
rect -14025 -30071 -13942 -29971
rect -11949 -30080 -11866 -29990
rect -11734 -30078 -11651 -29978
rect -11559 -30069 -11476 -29969
rect -6034 -30013 -5973 -29952
rect -5906 -30013 -5845 -29952
rect 750 -29996 852 -29952
rect 929 -29952 933 -29874
rect 933 -29952 1031 -29874
rect 1105 -29952 1207 -29882
rect 4925 -29929 5019 -29816
rect 5098 -29931 5192 -29818
rect 5287 -29925 5381 -29812
rect 929 -29988 1031 -29952
rect 1105 -29996 1207 -29952
rect 9213 -29964 9298 -29854
rect 9372 -29952 9457 -29856
rect 9539 -29952 9624 -29854
rect 12243 -29871 12311 -29781
rect 12389 -29860 12457 -29770
rect 12543 -29865 12611 -29775
rect 12700 -29865 12768 -29775
rect 12383 -29952 12451 -29941
rect 12545 -29952 12613 -29946
rect 20376 -29952 20441 -29939
rect 20507 -29952 20563 -29937
rect 20563 -29952 20572 -29937
rect 21109 -29827 21170 -29759
rect 21249 -29823 21310 -29755
rect 21790 -29815 21853 -29748
rect 9372 -29966 9457 -29952
rect 9539 -29964 9624 -29952
rect 4921 -30080 5015 -30026
rect 5100 -30080 5194 -30021
rect 5287 -30080 5381 -30019
rect 12229 -30042 12297 -29952
rect 12383 -30031 12451 -29952
rect 12545 -30036 12613 -29952
rect 12708 -30044 12776 -29954
rect 20376 -30008 20441 -29952
rect 20507 -30006 20572 -29952
rect 21107 -29960 21168 -29892
rect 21249 -29952 21310 -29888
rect 21717 -29937 21723 -29869
rect 21723 -29937 21778 -29869
rect 21865 -29935 21926 -29867
rect 33774 -29864 33828 -29806
rect 33885 -29863 33928 -29805
rect 33928 -29863 33939 -29805
rect 35213 -29851 35267 -29793
rect 35320 -29852 35374 -29794
rect 36560 -29867 36573 -29809
rect 36573 -29867 36614 -29809
rect 36706 -29867 36760 -29809
rect 38004 -29642 38058 -29624
rect 38058 -29642 38064 -29624
rect 38125 -29638 38185 -29624
rect 38005 -29753 38058 -29694
rect 38058 -29753 38065 -29694
rect 38129 -29754 38189 -29695
rect 38007 -29866 38058 -29807
rect 38058 -29866 38067 -29807
rect 38130 -29866 38184 -29808
rect 44612 -29864 44666 -29801
rect 44746 -29867 44800 -29804
rect 45839 -29810 45893 -29793
rect 45820 -29851 45893 -29810
rect 45820 -29873 45874 -29851
rect 45946 -29852 45978 -29794
rect 45978 -29807 46000 -29794
rect 45960 -29870 45978 -29852
rect 45978 -29870 46014 -29807
rect 46955 -29860 46968 -29792
rect 46968 -29860 47010 -29792
rect 47082 -29859 47136 -29796
rect 47957 -29833 47958 -29770
rect 47958 -29833 48011 -29770
rect 48094 -29833 48148 -29770
rect 49261 -29864 49273 -29801
rect 49273 -29864 49315 -29801
rect 49377 -29864 49431 -29801
rect 21249 -29956 21310 -29952
<< metal2 >>
rect -6162 24352 -5746 24354
rect -6162 24339 -5922 24352
rect -6162 24257 -6106 24339
rect -6013 24270 -5922 24339
rect -5829 24270 -5746 24352
rect -6013 24257 -5746 24270
rect -6162 24169 -5746 24257
rect -6162 24156 -5932 24169
rect -6162 24074 -6113 24156
rect -6020 24087 -5932 24156
rect -5839 24087 -5746 24169
rect 48489 24140 48958 24157
rect 48489 24138 48787 24140
rect 48489 24134 48680 24138
rect -6020 24074 -5746 24087
rect -6162 23984 -5746 24074
rect -6162 23979 -5934 23984
rect -6162 23897 -6128 23979
rect -6035 23902 -5934 23979
rect -5841 23902 -5746 23984
rect -6035 23897 -5746 23902
rect -6162 23854 -5746 23897
rect 165 24070 606 24083
rect 165 24067 530 24070
rect 165 24066 418 24067
rect 165 24007 198 24066
rect 250 24007 307 24066
rect 359 24008 418 24066
rect 470 24011 530 24067
rect 582 24011 606 24070
rect 470 24008 606 24011
rect 359 24007 606 24008
rect 165 23956 606 24007
rect 165 23955 529 23956
rect 165 23896 199 23955
rect 251 23896 308 23955
rect 360 23896 420 23955
rect 472 23897 529 23955
rect 581 23897 606 23956
rect 472 23896 606 23897
rect -6162 14895 -5982 23854
rect -4282 22512 -4099 22537
rect -4282 22403 -4271 22512
rect -4129 22403 -4099 22512
rect -6188 14854 -5946 14895
rect -6188 14851 -6045 14854
rect -6188 14782 -6169 14851
rect -6108 14785 -6045 14851
rect -5984 14785 -5946 14854
rect -6108 14782 -5946 14785
rect -6188 14728 -5946 14782
rect -6188 14723 -6042 14728
rect -6188 14654 -6171 14723
rect -6110 14659 -6042 14723
rect -5981 14659 -5946 14728
rect -6110 14654 -5946 14659
rect -6188 14625 -5946 14654
rect -4282 -1164 -4099 22403
rect -3601 22330 -3537 22331
rect -3601 22319 -3528 22330
rect -3601 22197 -3590 22319
rect -3536 22197 -3528 22319
rect -3601 22191 -3528 22197
rect -5987 -1168 -4099 -1164
rect -6368 -1347 -4099 -1168
rect -8457 -2317 -8299 -2316
rect -8459 -2354 -8297 -2317
rect -8459 -2446 -8415 -2354
rect -8338 -2446 -8297 -2354
rect -8459 -2480 -8297 -2446
rect -8457 -15490 -8299 -2480
rect -6368 -2839 -6185 -1347
rect -3599 -2531 -3528 22191
rect -2662 -2345 -2506 -2307
rect -2662 -2440 -2628 -2345
rect -2537 -2440 -2506 -2345
rect -2662 -2482 -2506 -2440
rect -6368 -2895 -5602 -2839
rect -6334 -2898 -5602 -2895
rect -6450 -3216 -6257 -3162
rect -6450 -3274 -6441 -3216
rect -6385 -3218 -6257 -3216
rect -6385 -3274 -6333 -3218
rect -6450 -3276 -6333 -3274
rect -6277 -3276 -6257 -3218
rect -4924 -3176 -4822 -3160
rect -3596 -3161 -3533 -2531
rect -2655 -3136 -2511 -2482
rect 165 -2516 606 23896
rect 160 -2532 606 -2516
rect 160 -2535 443 -2532
rect 160 -2652 224 -2535
rect 341 -2649 443 -2535
rect 560 -2649 606 -2532
rect 341 -2652 606 -2649
rect 160 -2711 606 -2652
rect 160 -2720 440 -2711
rect 160 -2837 221 -2720
rect 338 -2828 440 -2720
rect 557 -2828 606 -2711
rect 338 -2837 606 -2828
rect 160 -2901 606 -2837
rect -2657 -3161 -2500 -3136
rect -4924 -3243 -4906 -3176
rect -4843 -3243 -4822 -3176
rect -4924 -3257 -4822 -3243
rect -2657 -3223 -2624 -3161
rect -2542 -3223 -2500 -3161
rect -2657 -3247 -2500 -3223
rect -6450 -3291 -6257 -3276
rect -6448 -5446 -6257 -3291
rect -5197 -4234 -5129 -4222
rect -5197 -4286 -5187 -4234
rect -5135 -4286 -5129 -4234
rect -5197 -4292 -5129 -4286
rect -3889 -4231 -3795 -4223
rect -3889 -4288 -3876 -4231
rect -3809 -4288 -3795 -4231
rect -5190 -4962 -5133 -4292
rect -3889 -4307 -3795 -4288
rect -5218 -5003 -5009 -4962
rect -5218 -5010 -5077 -5003
rect -5218 -5068 -5193 -5010
rect -5131 -5061 -5077 -5010
rect -5015 -5061 -5009 -5003
rect -5131 -5068 -5009 -5061
rect -5218 -5127 -5009 -5068
rect -5218 -5185 -5193 -5127
rect -5131 -5185 -5075 -5127
rect -5013 -5185 -5009 -5127
rect -5218 -5204 -5009 -5185
rect -5190 -5206 -5133 -5204
rect -6448 -5504 -6423 -5446
rect -6367 -5492 -6257 -5446
rect -6367 -5504 -6315 -5492
rect -6448 -5550 -6315 -5504
rect -6259 -5550 -6257 -5492
rect -6448 -5562 -6257 -5550
rect -6448 -5620 -6423 -5562
rect -6367 -5620 -6257 -5562
rect -6448 -5647 -6257 -5620
rect -7866 -7621 -7591 -7609
rect -7866 -7716 -7693 -7621
rect -7609 -7716 -7591 -7621
rect -7866 -7730 -7591 -7716
rect -7866 -7825 -7836 -7730
rect -7752 -7825 -7591 -7730
rect -7866 -7850 -7591 -7825
rect -8457 -15562 -8417 -15490
rect -8351 -15562 -8299 -15490
rect -8457 -15576 -8299 -15562
rect -10434 -16894 -9984 -16877
rect -8334 -16894 -8027 -16886
rect -10434 -16902 -8027 -16894
rect -10434 -16903 -8130 -16902
rect -10434 -16924 -8300 -16903
rect -10434 -16929 -10159 -16924
rect -10434 -17050 -10386 -16929
rect -10278 -17045 -10159 -16929
rect -10051 -17000 -8300 -16924
rect -8210 -16999 -8130 -16903
rect -8040 -16999 -8027 -16902
rect -8210 -17000 -8027 -16999
rect -10051 -17045 -8027 -17000
rect -10278 -17050 -8027 -17045
rect -10434 -17067 -8027 -17050
rect -10434 -17070 -8130 -17067
rect -10434 -17140 -8300 -17070
rect -10434 -17144 -10159 -17140
rect -10434 -17265 -10386 -17144
rect -10278 -17261 -10159 -17144
rect -10051 -17167 -8300 -17140
rect -8210 -17164 -8130 -17070
rect -8040 -17164 -8027 -17067
rect -8210 -17167 -8027 -17164
rect -10051 -17202 -8027 -17167
rect -10051 -17261 -9984 -17202
rect -8334 -17207 -8027 -17202
rect -10278 -17265 -9984 -17261
rect -10434 -17309 -9984 -17265
rect -8460 -18001 -8294 -17969
rect -8460 -18073 -8411 -18001
rect -8345 -18073 -8294 -18001
rect -27398 -26327 -26825 -26289
rect -27398 -26333 -27172 -26327
rect -27398 -26438 -27358 -26333
rect -27265 -26432 -27172 -26333
rect -27079 -26432 -26953 -26327
rect -26860 -26432 -26825 -26327
rect -27265 -26438 -26825 -26432
rect -27398 -26516 -26825 -26438
rect -27398 -26522 -26965 -26516
rect -27398 -26528 -27166 -26522
rect -27398 -26633 -27352 -26528
rect -27259 -26627 -27166 -26528
rect -27073 -26621 -26965 -26522
rect -26872 -26621 -26825 -26516
rect -27073 -26627 -26825 -26621
rect -27259 -26633 -26825 -26627
rect -27398 -29816 -26825 -26633
rect -27398 -29821 -26994 -29816
rect -27398 -29921 -27343 -29821
rect -27260 -29921 -27172 -29821
rect -27089 -29916 -26994 -29821
rect -26911 -29916 -26825 -29816
rect -27089 -29921 -26825 -29916
rect -27398 -30008 -26825 -29921
rect -27398 -30019 -26978 -30008
rect -27398 -30021 -27170 -30019
rect -27398 -30080 -27348 -30021
rect -27265 -30080 -27170 -30021
rect -27087 -30080 -26978 -30019
rect -26895 -30080 -26825 -30008
rect -27398 -30125 -26825 -30080
rect -24972 -26327 -24399 -26306
rect -24972 -26342 -24699 -26327
rect -24972 -26447 -24900 -26342
rect -24807 -26432 -24699 -26342
rect -24606 -26333 -24399 -26327
rect -24606 -26432 -24510 -26333
rect -24807 -26438 -24510 -26432
rect -24417 -26438 -24399 -26333
rect -24807 -26447 -24399 -26438
rect -24972 -26522 -24399 -26447
rect -24972 -26531 -24516 -26522
rect -24972 -26545 -24693 -26531
rect -24972 -26650 -24914 -26545
rect -24821 -26636 -24693 -26545
rect -24600 -26627 -24516 -26531
rect -24423 -26627 -24399 -26522
rect -24600 -26636 -24399 -26627
rect -24821 -26650 -24399 -26636
rect -24972 -29778 -24399 -26650
rect -24972 -29789 -24542 -29778
rect -24972 -29798 -24751 -29789
rect -24972 -29898 -24934 -29798
rect -24851 -29889 -24751 -29798
rect -24668 -29878 -24542 -29789
rect -24459 -29878 -24399 -29778
rect -24668 -29889 -24399 -29878
rect -24851 -29898 -24399 -29889
rect -24972 -29974 -24399 -29898
rect -24972 -29980 -24537 -29974
rect -24972 -29994 -24738 -29980
rect -24972 -30080 -24929 -29994
rect -24846 -30080 -24738 -29994
rect -24655 -30074 -24537 -29980
rect -24454 -30074 -24399 -29974
rect -24655 -30080 -24399 -30074
rect -24972 -30147 -24399 -30080
rect -22412 -26374 -21839 -26318
rect -22412 -26377 -22057 -26374
rect -22412 -26482 -22310 -26377
rect -22217 -26479 -22057 -26377
rect -21964 -26479 -21839 -26374
rect -22217 -26482 -21839 -26479
rect -22412 -26542 -21839 -26482
rect -22412 -26545 -21958 -26542
rect -22412 -26551 -22150 -26545
rect -22412 -26656 -22372 -26551
rect -22279 -26650 -22150 -26551
rect -22057 -26647 -21958 -26545
rect -21865 -26647 -21839 -26542
rect -22057 -26650 -21839 -26647
rect -22279 -26656 -21839 -26650
rect -22412 -29788 -21839 -26656
rect -22412 -29793 -21972 -29788
rect -22412 -29893 -22352 -29793
rect -22269 -29893 -22165 -29793
rect -22082 -29888 -21972 -29793
rect -21889 -29888 -21839 -29788
rect -22082 -29893 -21839 -29888
rect -22412 -29971 -21839 -29893
rect -22412 -29976 -21978 -29971
rect -22412 -30076 -22358 -29976
rect -22275 -30076 -22171 -29976
rect -22088 -30071 -21978 -29976
rect -21895 -30071 -21839 -29971
rect -22088 -30076 -21839 -30071
rect -22412 -30107 -21839 -30076
rect -19876 -26374 -19303 -26329
rect -19876 -26479 -19777 -26374
rect -19684 -26475 -19547 -26374
rect -19454 -26475 -19303 -26374
rect -19684 -26479 -19303 -26475
rect -19876 -26528 -19303 -26479
rect -19876 -26542 -19442 -26528
rect -19876 -26554 -19628 -26542
rect -19876 -26659 -19823 -26554
rect -19730 -26647 -19628 -26554
rect -19535 -26633 -19442 -26542
rect -19349 -26633 -19303 -26528
rect -19535 -26647 -19303 -26633
rect -19730 -26659 -19303 -26647
rect -19876 -29787 -19303 -26659
rect -19876 -29796 -19407 -29787
rect -19876 -29798 -19598 -29796
rect -19876 -29898 -19805 -29798
rect -19722 -29896 -19598 -29798
rect -19515 -29887 -19407 -29796
rect -19324 -29887 -19303 -29787
rect -19515 -29896 -19303 -29887
rect -19722 -29898 -19303 -29896
rect -19876 -29974 -19303 -29898
rect -19876 -29976 -19411 -29974
rect -19876 -29992 -19603 -29976
rect -19876 -30080 -19821 -29992
rect -19738 -30076 -19603 -29992
rect -19520 -30074 -19411 -29976
rect -19328 -30074 -19303 -29974
rect -19520 -30076 -19303 -30074
rect -19738 -30080 -19303 -30076
rect -19876 -30117 -19303 -30080
rect -17362 -26353 -16789 -26295
rect -17362 -26359 -16934 -26353
rect -17362 -26464 -17292 -26359
rect -17199 -26464 -17089 -26359
rect -16996 -26458 -16934 -26359
rect -16841 -26458 -16789 -26353
rect -16996 -26464 -16789 -26458
rect -17362 -26534 -16789 -26464
rect -17362 -26540 -16920 -26534
rect -17362 -26645 -17310 -26540
rect -17217 -26542 -16920 -26540
rect -17217 -26645 -17121 -26542
rect -17362 -26647 -17121 -26645
rect -17028 -26639 -16920 -26542
rect -16827 -26639 -16789 -26534
rect -17028 -26647 -16789 -26639
rect -17362 -29778 -16789 -26647
rect -17362 -29782 -17118 -29778
rect -17362 -29882 -17294 -29782
rect -17211 -29878 -17118 -29782
rect -17035 -29878 -16929 -29778
rect -16846 -29878 -16789 -29778
rect -17211 -29882 -16789 -29878
rect -17362 -29985 -16789 -29882
rect -17362 -30080 -17303 -29985
rect -17220 -29987 -16918 -29985
rect -17220 -30080 -17116 -29987
rect -17033 -30080 -16918 -29987
rect -16835 -30080 -16789 -29985
rect -17362 -30114 -16789 -30080
rect -14443 -26350 -13870 -26306
rect -14443 -26362 -13993 -26350
rect -14443 -26374 -14159 -26362
rect -14443 -26479 -14372 -26374
rect -14279 -26467 -14159 -26374
rect -14066 -26455 -13993 -26362
rect -13900 -26455 -13870 -26350
rect -14066 -26467 -13870 -26455
rect -14279 -26479 -13870 -26467
rect -14443 -26519 -13870 -26479
rect -14443 -26531 -13982 -26519
rect -14443 -26636 -14372 -26531
rect -14279 -26636 -14162 -26531
rect -14069 -26624 -13982 -26531
rect -13889 -26624 -13870 -26519
rect -14069 -26636 -13870 -26624
rect -14443 -29784 -13870 -26636
rect -14443 -29789 -14203 -29784
rect -14443 -29889 -14376 -29789
rect -14293 -29884 -14203 -29789
rect -14120 -29884 -14030 -29784
rect -13947 -29884 -13870 -29784
rect -14293 -29889 -13870 -29884
rect -14443 -29971 -13870 -29889
rect -14443 -29974 -14025 -29971
rect -14443 -29980 -14203 -29974
rect -14443 -30080 -14383 -29980
rect -14300 -30074 -14203 -29980
rect -14120 -30071 -14025 -29974
rect -13942 -30071 -13870 -29971
rect -14120 -30074 -13870 -30071
rect -14300 -30080 -13870 -30074
rect -14443 -30118 -13870 -30080
rect -12011 -26359 -11438 -26329
rect -12011 -26362 -11570 -26359
rect -12011 -26365 -11780 -26362
rect -12011 -26470 -11963 -26365
rect -11870 -26467 -11780 -26365
rect -11687 -26464 -11570 -26362
rect -11477 -26464 -11438 -26359
rect -11687 -26467 -11438 -26464
rect -11870 -26470 -11438 -26467
rect -12011 -26525 -11438 -26470
rect -12011 -26534 -11582 -26525
rect -12011 -26542 -11797 -26534
rect -12011 -26647 -11972 -26542
rect -11879 -26639 -11797 -26542
rect -11704 -26630 -11582 -26534
rect -11489 -26630 -11438 -26525
rect -11704 -26639 -11438 -26630
rect -11879 -26647 -11438 -26639
rect -12011 -29778 -11438 -26647
rect -8460 -27177 -8294 -18073
rect -8460 -27301 -8446 -27177
rect -8317 -27301 -8294 -27177
rect -8460 -27312 -8294 -27301
rect -12011 -29782 -11552 -29778
rect -12011 -29784 -11741 -29782
rect -12011 -29884 -11942 -29784
rect -11859 -29882 -11741 -29784
rect -11658 -29878 -11552 -29782
rect -11469 -29878 -11438 -29778
rect -11658 -29882 -11438 -29878
rect -11859 -29884 -11438 -29882
rect -12011 -29969 -11438 -29884
rect -12011 -29978 -11559 -29969
rect -12011 -29990 -11734 -29978
rect -12011 -30080 -11949 -29990
rect -11866 -30078 -11734 -29990
rect -11651 -30069 -11559 -29978
rect -11476 -30069 -11438 -29969
rect -11651 -30078 -11438 -30069
rect -11866 -30080 -11438 -30078
rect -12011 -30122 -11438 -30080
rect -7849 -32424 -7601 -7850
rect 165 -8211 606 -2901
rect 165 -8215 545 -8211
rect 165 -8216 437 -8215
rect 165 -8275 218 -8216
rect 270 -8275 323 -8216
rect 375 -8274 437 -8216
rect 489 -8270 545 -8215
rect 597 -8270 606 -8211
rect 489 -8274 606 -8270
rect 375 -8275 606 -8274
rect 165 -8298 606 -8275
rect 1197 24070 1638 24083
rect 1197 24067 1562 24070
rect 1197 24066 1450 24067
rect 1197 24007 1230 24066
rect 1282 24007 1339 24066
rect 1391 24008 1450 24066
rect 1502 24011 1562 24067
rect 1614 24011 1638 24070
rect 1502 24008 1638 24011
rect 1391 24007 1638 24008
rect 1197 23956 1638 24007
rect 1197 23955 1561 23956
rect 1197 23896 1231 23955
rect 1283 23896 1340 23955
rect 1392 23896 1452 23955
rect 1504 23897 1561 23955
rect 1613 23897 1638 23956
rect 1504 23896 1638 23897
rect 1197 -8203 1638 23896
rect 24705 24009 25123 24125
rect 24705 24002 25018 24009
rect 24705 23996 24864 24002
rect 24705 23926 24725 23996
rect 24798 23932 24864 23996
rect 24937 23939 25018 24002
rect 25091 23939 25123 24009
rect 24937 23932 25123 23939
rect 24798 23926 25123 23932
rect 22905 23415 23050 23438
rect 22905 23308 22923 23415
rect 23021 23308 23050 23415
rect 4558 22092 5130 22110
rect 4558 22091 5008 22092
rect 4558 21969 4621 22091
rect 4724 21969 4808 22091
rect 4911 21970 5008 22091
rect 5111 21970 5130 22092
rect 4911 21969 5130 21970
rect 4558 21892 5130 21969
rect 4558 21770 4624 21892
rect 4727 21890 5007 21892
rect 4727 21770 4814 21890
rect 4558 21768 4814 21770
rect 4917 21770 5007 21890
rect 5110 21770 5130 21892
rect 4917 21768 5130 21770
rect 4558 -4703 5130 21768
rect 22905 20322 23050 23308
rect 23166 23182 23311 23194
rect 23166 23075 23184 23182
rect 23282 23075 23311 23182
rect 23166 20279 23311 23075
rect 23505 22881 23646 22894
rect 23505 22774 23521 22881
rect 23619 22774 23646 22881
rect 23505 20281 23646 22774
rect 24705 20049 25123 23926
rect 24705 20043 25037 20049
rect 24705 20040 24887 20043
rect 24705 19970 24736 20040
rect 24809 19973 24887 20040
rect 24960 19979 25037 20043
rect 25110 19979 25123 20049
rect 24960 19973 25123 19979
rect 24809 19970 25123 19973
rect 24705 19903 25123 19970
rect 26123 24096 26541 24106
rect 26123 24088 26429 24096
rect 26123 24087 26300 24088
rect 26123 24017 26160 24087
rect 26233 24018 26300 24087
rect 26373 24026 26429 24088
rect 26502 24026 26541 24096
rect 26373 24018 26541 24026
rect 26233 24017 26541 24018
rect 26123 23962 26541 24017
rect 26123 23959 26437 23962
rect 26123 23958 26302 23959
rect 26123 23888 26157 23958
rect 26230 23889 26302 23958
rect 26375 23892 26437 23959
rect 26510 23892 26541 23962
rect 26375 23889 26541 23892
rect 26230 23888 26541 23889
rect 26123 20071 26541 23888
rect 26123 20063 26444 20071
rect 26123 20059 26302 20063
rect 26123 19989 26155 20059
rect 26228 19993 26302 20059
rect 26375 20001 26444 20063
rect 26517 20001 26541 20071
rect 26375 19993 26541 20001
rect 26228 19989 26541 19993
rect 26123 19960 26541 19989
rect 27528 24084 27946 24087
rect 27528 24082 27850 24084
rect 27528 24077 27699 24082
rect 27528 24007 27546 24077
rect 27619 24012 27699 24077
rect 27772 24014 27850 24082
rect 27923 24014 27946 24084
rect 27772 24012 27946 24014
rect 27619 24007 27946 24012
rect 27528 23961 27946 24007
rect 27528 23959 27853 23961
rect 27528 23950 27699 23959
rect 27528 23880 27544 23950
rect 27617 23889 27699 23950
rect 27772 23891 27853 23959
rect 27926 23891 27946 23961
rect 27772 23889 27946 23891
rect 27617 23880 27946 23889
rect 27528 20073 27946 23880
rect 27528 20063 27836 20073
rect 27528 20059 27694 20063
rect 27528 19989 27557 20059
rect 27630 19993 27694 20059
rect 27767 20003 27836 20063
rect 27909 20003 27946 20073
rect 27767 19993 27946 20003
rect 27630 19989 27946 19993
rect 27528 19941 27946 19989
rect 48489 24081 48564 24134
rect 48616 24084 48680 24134
rect 48735 24086 48787 24138
rect 48842 24086 48958 24140
rect 48735 24084 48958 24086
rect 48616 24081 48958 24084
rect 48489 24031 48958 24081
rect 48489 24023 48679 24031
rect 48489 23970 48560 24023
rect 48612 23978 48679 24023
rect 48731 24027 48958 24031
rect 48731 23978 48786 24027
rect 48612 23974 48786 23978
rect 48838 23974 48958 24027
rect 48612 23970 48958 23974
rect 48489 23919 48958 23970
rect 48489 23912 48744 23919
rect 48489 23857 48615 23912
rect 48677 23864 48744 23912
rect 48806 23864 48958 23919
rect 48677 23857 48958 23864
rect 47175 -1923 47489 -1873
rect 47175 -1953 47198 -1923
rect 47173 -1992 47198 -1953
rect 47271 -1929 47489 -1923
rect 47271 -1992 47373 -1929
rect 47173 -1998 47373 -1992
rect 47446 -1998 47489 -1929
rect 47173 -2088 47489 -1998
rect 47173 -2157 47197 -2088
rect 47270 -2091 47489 -2088
rect 47270 -2157 47370 -2091
rect 47173 -2160 47370 -2157
rect 47443 -2160 47489 -2091
rect 47173 -2182 47489 -2160
rect 8335 -4129 8569 -4093
rect 8335 -4130 8483 -4129
rect 8335 -4205 8348 -4130
rect 8422 -4204 8483 -4130
rect 8557 -4204 8569 -4129
rect 8422 -4205 8569 -4204
rect 8335 -4288 8569 -4205
rect 8335 -4289 8482 -4288
rect 8335 -4364 8346 -4289
rect 8420 -4363 8482 -4289
rect 8556 -4363 8569 -4288
rect 8420 -4364 8569 -4363
rect 8335 -4376 8569 -4364
rect 4558 -4815 4886 -4703
rect 4988 -4815 5130 -4703
rect 3194 -7636 3334 -7626
rect 3194 -7703 3215 -7636
rect 3304 -7703 3334 -7636
rect 3194 -7755 3334 -7703
rect 3194 -7822 3214 -7755
rect 3303 -7822 3334 -7755
rect 3194 -7858 3334 -7822
rect 1197 -8205 1584 -8203
rect 1197 -8208 1473 -8205
rect 1197 -8209 1346 -8208
rect 1197 -8268 1227 -8209
rect 1279 -8267 1346 -8209
rect 1398 -8264 1473 -8208
rect 1525 -8262 1584 -8205
rect 1636 -8262 1638 -8203
rect 1525 -8264 1638 -8262
rect 1398 -8267 1638 -8264
rect 1279 -8268 1638 -8267
rect 1197 -8286 1638 -8268
rect -7298 -9191 -5924 -9027
rect -7298 -12428 -7124 -9191
rect -6020 -9492 -5925 -9191
rect -6020 -9553 -6009 -9492
rect -5941 -9553 -5925 -9492
rect 3207 -9508 3282 -7858
rect -6020 -9571 -5925 -9553
rect 4097 -10186 4258 -10174
rect 4097 -10238 4110 -10186
rect 4176 -10238 4258 -10186
rect 4097 -10297 4258 -10238
rect 4097 -10349 4138 -10297
rect 4233 -10349 4258 -10297
rect 4097 -10366 4258 -10349
rect -7296 -32424 -7124 -12428
rect 702 -11659 962 -11569
rect 702 -11661 882 -11659
rect 702 -11722 750 -11661
rect 809 -11720 882 -11661
rect 941 -11720 962 -11659
rect 809 -11722 962 -11720
rect -6856 -14805 -6689 -14783
rect -6856 -14889 -6830 -14805
rect -6723 -14889 -6689 -14805
rect -6856 -14908 -6689 -14889
rect -6855 -24446 -6691 -14908
rect -6070 -16463 -5812 -16403
rect -6070 -16517 -6045 -16463
rect -5991 -16517 -5923 -16463
rect -5869 -16517 -5812 -16463
rect -6070 -18553 -5812 -16517
rect -3235 -17518 -2995 -17492
rect -3235 -17676 -3210 -17518
rect -3022 -17676 -2995 -17518
rect -3235 -17720 -2995 -17676
rect -3766 -18136 -3503 -18106
rect -3766 -18245 -3731 -18136
rect -3599 -18245 -3503 -18136
rect -3766 -18321 -3503 -18245
rect -3766 -18430 -3731 -18321
rect -3599 -18430 -3503 -18321
rect -3766 -18445 -3503 -18430
rect -6855 -24460 -6688 -24446
rect -6855 -24463 -6744 -24460
rect -6855 -24519 -6849 -24463
rect -6796 -24518 -6744 -24463
rect -6691 -24518 -6688 -24460
rect -6796 -24519 -6688 -24518
rect -6855 -24531 -6688 -24519
rect -6855 -32424 -6691 -24531
rect -6068 -29808 -5813 -18553
rect -3765 -22847 -3504 -18445
rect -3220 -20700 -3000 -17720
rect 702 -18690 962 -11722
rect 4104 -17505 4251 -10366
rect 4082 -17532 4272 -17505
rect 4082 -17682 4113 -17532
rect 4249 -17682 4272 -17532
rect 4082 -17720 4272 -17682
rect 4558 -18108 5130 -4815
rect 5232 -4981 5370 -4933
rect 5232 -5051 5255 -4981
rect 5326 -5051 5370 -4981
rect 5232 -5121 5370 -5051
rect 5232 -5191 5253 -5121
rect 5324 -5191 5370 -5121
rect 5232 -5220 5370 -5191
rect 4557 -18167 5130 -18108
rect 4557 -18168 4918 -18167
rect 4557 -18262 4591 -18168
rect 4670 -18170 4918 -18168
rect 4670 -18262 4752 -18170
rect 4557 -18264 4752 -18262
rect 4831 -18261 4918 -18170
rect 4997 -18236 5130 -18167
rect 4997 -18261 5053 -18236
rect 4831 -18264 5053 -18261
rect 4557 -18330 5053 -18264
rect 5121 -18307 5130 -18236
rect 5121 -18330 5129 -18307
rect 4557 -18332 5129 -18330
rect 4557 -18426 4593 -18332
rect 4672 -18426 4753 -18332
rect 4832 -18426 4919 -18332
rect 4998 -18426 5129 -18332
rect 4557 -18446 5129 -18426
rect 264 -18752 962 -18690
rect 264 -18754 444 -18752
rect 264 -18812 303 -18754
rect 370 -18810 444 -18754
rect 511 -18810 962 -18752
rect 370 -18812 962 -18810
rect 264 -18875 962 -18812
rect 264 -18881 445 -18875
rect 264 -18939 301 -18881
rect 368 -18933 445 -18881
rect 512 -18933 962 -18875
rect 368 -18939 962 -18933
rect 264 -18959 962 -18939
rect 274 -18961 534 -18959
rect -3222 -20727 -2992 -20700
rect -3222 -20813 -3171 -20727
rect -3026 -20813 -2992 -20727
rect 5252 -20785 5369 -5220
rect 5444 -5427 5564 -5387
rect 5444 -5498 5466 -5427
rect 5531 -5498 5564 -5427
rect 5444 -5562 5564 -5498
rect 5444 -5633 5468 -5562
rect 5533 -5633 5564 -5562
rect 5444 -5664 5564 -5633
rect 5457 -20569 5526 -5664
rect 7183 -6820 7485 -6777
rect 7183 -6997 7245 -6820
rect 7439 -6997 7485 -6820
rect 7183 -7086 7485 -6997
rect 8364 -13575 8534 -4376
rect 28896 -13122 29195 -13054
rect 28896 -13299 28957 -13122
rect 29123 -13299 29195 -13122
rect 8292 -13591 8620 -13575
rect 8292 -13593 8518 -13591
rect 8292 -13682 8337 -13593
rect 8414 -13680 8518 -13593
rect 8595 -13680 8620 -13591
rect 8414 -13682 8620 -13680
rect 8292 -13736 8620 -13682
rect 8292 -13825 8340 -13736
rect 8417 -13825 8518 -13736
rect 8595 -13825 8620 -13736
rect 8292 -13897 8620 -13825
rect 8292 -13986 8340 -13897
rect 8417 -13986 8516 -13897
rect 8593 -13986 8620 -13897
rect 8292 -14013 8620 -13986
rect 25393 -13582 25628 -13576
rect 25393 -13649 25459 -13582
rect 25555 -13649 25628 -13582
rect 25393 -13706 25628 -13649
rect 25393 -13805 25453 -13706
rect 25552 -13805 25628 -13706
rect 25393 -13873 25628 -13805
rect 25393 -13972 25452 -13873
rect 25551 -13972 25628 -13873
rect 25393 -14016 25628 -13972
rect 13232 -15685 13507 -15668
rect 13232 -15767 13245 -15685
rect 13319 -15689 13507 -15685
rect 13319 -15767 13391 -15689
rect 13232 -15771 13391 -15767
rect 13465 -15771 13507 -15689
rect 13232 -15832 13507 -15771
rect 13232 -15845 13396 -15832
rect 13232 -15927 13244 -15845
rect 13318 -15914 13396 -15845
rect 13470 -15914 13507 -15832
rect 13318 -15927 13507 -15914
rect 13232 -15945 13507 -15927
rect 13280 -17273 13487 -15945
rect 13641 -16092 13920 -16086
rect 13641 -16096 13815 -16092
rect 13641 -16172 13660 -16096
rect 13742 -16168 13815 -16096
rect 13897 -16168 13920 -16092
rect 13742 -16172 13920 -16168
rect 13641 -16228 13920 -16172
rect 13641 -16237 13813 -16228
rect 13641 -16313 13662 -16237
rect 13744 -16304 13813 -16237
rect 13895 -16304 13920 -16228
rect 13744 -16313 13920 -16304
rect 13641 -16334 13920 -16313
rect 25469 -16331 25573 -14016
rect 7854 -17431 13487 -17273
rect 7340 -19753 7460 -19743
rect 7340 -19830 7352 -19753
rect 7439 -19761 7460 -19753
rect 7441 -19830 7460 -19761
rect 7340 -19844 7460 -19830
rect 5457 -20636 5819 -20569
rect -3222 -20845 -2992 -20813
rect 5248 -20807 5379 -20785
rect 5248 -20868 5276 -20807
rect 5347 -20868 5379 -20807
rect 5248 -20899 5379 -20868
rect -3099 -21572 -2985 -21548
rect -3099 -21667 -3084 -21572
rect -3009 -21667 -2985 -21572
rect -3099 -21688 -2985 -21667
rect -3765 -22909 -3725 -22847
rect -3665 -22848 -3504 -22847
rect -3665 -22909 -3602 -22848
rect -3765 -22910 -3602 -22909
rect -3542 -22910 -3504 -22848
rect -3765 -22925 -3504 -22910
rect -3085 -25016 -3004 -21688
rect -1802 -21808 -1721 -21799
rect -1802 -21861 -1789 -21808
rect -1734 -21861 -1721 -21808
rect -2646 -24630 -2583 -23587
rect -1802 -24462 -1721 -21861
rect 5752 -21953 5819 -20636
rect 7081 -20812 7166 -20797
rect 7081 -20878 7091 -20812
rect 7148 -20878 7166 -20812
rect 7081 -20893 7166 -20878
rect 6176 -21922 6239 -20915
rect 7093 -21394 7161 -20893
rect 7083 -21417 7183 -21394
rect 7083 -21489 7104 -21417
rect 7163 -21489 7183 -21417
rect 7083 -21510 7183 -21489
rect 5743 -21966 5829 -21953
rect 5743 -22022 5753 -21966
rect 5813 -22022 5829 -21966
rect 5743 -22035 5829 -22022
rect 5752 -22857 5819 -22035
rect 5882 -22505 6003 -22493
rect 5882 -22558 5909 -22505
rect 5981 -22558 6003 -22505
rect 5882 -22570 6003 -22558
rect 5742 -22871 5828 -22857
rect 5742 -22926 5756 -22871
rect 5813 -22926 5828 -22871
rect 5742 -22939 5828 -22926
rect -1644 -23897 -1570 -23888
rect -1644 -23959 -1635 -23897
rect -1579 -23959 -1570 -23897
rect -1644 -23971 -1570 -23959
rect -1802 -24518 -1789 -24462
rect -1735 -24518 -1721 -24462
rect -1802 -24530 -1721 -24518
rect -2650 -24670 -2540 -24630
rect -2650 -24740 -2630 -24670
rect -2570 -24740 -2540 -24670
rect -2650 -24770 -2540 -24740
rect -1635 -24826 -1578 -23971
rect 5898 -24056 5996 -22570
rect 6176 -23646 6239 -22613
rect 7095 -23012 7210 -22992
rect 7095 -23072 7120 -23012
rect 7191 -23072 7210 -23012
rect 7095 -23089 7210 -23072
rect 6154 -23650 6256 -23646
rect 6154 -23702 6169 -23650
rect 6238 -23702 6256 -23650
rect 6154 -23755 6256 -23702
rect 6154 -23807 6171 -23755
rect 6240 -23807 6256 -23755
rect 6154 -23823 6256 -23807
rect 5875 -24074 6025 -24056
rect 5875 -24141 5895 -24074
rect 5996 -24141 6025 -24074
rect 5875 -24161 6025 -24141
rect 697 -24265 1283 -24222
rect 697 -24267 1128 -24265
rect 697 -24273 949 -24267
rect 697 -24387 764 -24273
rect 866 -24381 949 -24273
rect 1051 -24379 1128 -24267
rect 1230 -24379 1283 -24265
rect 1051 -24381 1283 -24379
rect 866 -24387 1283 -24381
rect -1684 -24846 -1540 -24826
rect -1684 -24909 -1652 -24846
rect -1570 -24909 -1540 -24846
rect -1684 -24923 -1540 -24909
rect -3085 -25069 -3075 -25016
rect -3017 -25069 -3004 -25016
rect -3085 -25084 -3004 -25069
rect -6068 -29816 -5902 -29808
rect -6068 -29881 -6034 -29816
rect -5973 -29873 -5902 -29816
rect -5841 -29873 -5813 -29808
rect -5973 -29881 -5813 -29873
rect -6068 -29948 -5813 -29881
rect -6068 -30013 -6034 -29948
rect -5973 -30013 -5906 -29948
rect -5845 -30013 -5813 -29948
rect -6068 -30049 -5813 -30013
rect 697 -29874 1283 -24387
rect 4889 -24267 5497 -24245
rect 4889 -24279 5333 -24267
rect 4889 -24287 5131 -24279
rect 4889 -24401 4937 -24287
rect 5039 -24393 5131 -24287
rect 5233 -24381 5333 -24279
rect 5435 -24381 5497 -24267
rect 5233 -24393 5497 -24381
rect 5039 -24401 5497 -24393
rect 4331 -24837 4422 -24827
rect 4331 -24896 4356 -24837
rect 4413 -24896 4422 -24837
rect 4331 -24919 4422 -24896
rect 697 -29882 929 -29874
rect 697 -29996 750 -29882
rect 852 -29988 929 -29882
rect 1031 -29882 1283 -29874
rect 1031 -29988 1105 -29882
rect 852 -29996 1105 -29988
rect 1207 -29996 1283 -29882
rect 697 -30080 1283 -29996
rect 4351 -32424 4408 -24919
rect 4540 -25014 4621 -25002
rect 4540 -25085 4546 -25014
rect 4608 -25085 4621 -25014
rect 4540 -32424 4621 -25085
rect 4889 -29812 5497 -24401
rect 6176 -24610 6239 -23823
rect 6160 -24650 6290 -24610
rect 6160 -24750 6180 -24650
rect 6270 -24750 6290 -24650
rect 6160 -24780 6290 -24750
rect 4889 -29816 5287 -29812
rect 4889 -29929 4925 -29816
rect 5019 -29818 5287 -29816
rect 5019 -29929 5098 -29818
rect 4889 -29931 5098 -29929
rect 5192 -29925 5287 -29818
rect 5381 -29925 5497 -29812
rect 5192 -29931 5497 -29925
rect 4889 -30019 5497 -29931
rect 4889 -30021 5287 -30019
rect 4889 -30026 5100 -30021
rect 4889 -30080 4921 -30026
rect 5015 -30080 5100 -30026
rect 5194 -30080 5287 -30021
rect 5381 -30080 5497 -30019
rect 4889 -30154 5497 -30080
rect 6176 -32424 6239 -24780
rect 6500 -25730 6620 -25710
rect 6500 -25800 6520 -25730
rect 6590 -25800 6620 -25730
rect 6500 -25830 6620 -25800
rect 6519 -32424 6581 -25830
rect 7104 -32424 7197 -23089
rect 7362 -32424 7448 -19844
rect 7854 -21654 7934 -17431
rect 13673 -17523 13856 -16334
rect 25469 -16435 26737 -16331
rect 14370 -16789 14736 -16761
rect 14370 -16793 14539 -16789
rect 14370 -16868 14391 -16793
rect 14455 -16864 14539 -16793
rect 14603 -16864 14669 -16789
rect 14733 -16864 14736 -16789
rect 14455 -16868 14736 -16864
rect 14370 -16942 14736 -16868
rect 14370 -16943 14669 -16942
rect 14370 -16946 14537 -16943
rect 14370 -17021 14391 -16946
rect 14455 -17018 14537 -16946
rect 14601 -17017 14669 -16943
rect 14733 -17017 14736 -16942
rect 14601 -17018 14736 -17017
rect 14455 -17021 14736 -17018
rect 14370 -17107 14736 -17021
rect 14370 -17182 14391 -17107
rect 14455 -17182 14530 -17107
rect 14594 -17182 14669 -17107
rect 14733 -17182 14736 -17107
rect 14370 -17203 14736 -17182
rect 8083 -17706 13856 -17523
rect 8083 -21228 8177 -17706
rect 8328 -18723 8565 -18703
rect 8328 -18724 8452 -18723
rect 8328 -18796 8343 -18724
rect 8399 -18795 8452 -18724
rect 8508 -18795 8565 -18723
rect 8399 -18796 8565 -18795
rect 8328 -18814 8565 -18796
rect 11737 -18729 11815 -18700
rect 11737 -18800 11743 -18729
rect 11806 -18800 11815 -18729
rect 11737 -18814 11815 -18800
rect 8326 -18974 8509 -18943
rect 8326 -19081 8375 -18974
rect 8467 -19081 8509 -18974
rect 8326 -20913 8509 -19081
rect 11292 -20748 11358 -20587
rect 8326 -20972 8365 -20913
rect 8457 -20972 8509 -20913
rect 8326 -20996 8509 -20972
rect 10761 -20814 11358 -20748
rect 8083 -21322 8283 -21228
rect 10501 -21300 10641 -21299
rect 10501 -21371 10693 -21300
rect 7854 -21734 8280 -21654
rect 8678 -21984 8793 -21974
rect 8678 -22053 8699 -21984
rect 8770 -22053 8793 -21984
rect 7592 -22524 7696 -22495
rect 7592 -22582 7609 -22524
rect 7664 -22582 7696 -22524
rect 7592 -22599 7696 -22582
rect 7592 -23403 7695 -22599
rect 7592 -23476 7611 -23403
rect 7680 -23476 7695 -23403
rect 7592 -23491 7695 -23476
rect 8678 -24041 8793 -22053
rect 8678 -24116 8694 -24041
rect 8777 -24116 8793 -24041
rect 8678 -24138 8793 -24116
rect 9148 -24248 9756 -24177
rect 9148 -24250 9412 -24248
rect 9148 -24364 9210 -24250
rect 9312 -24362 9412 -24250
rect 9514 -24362 9605 -24248
rect 9707 -24362 9756 -24248
rect 9312 -24364 9756 -24362
rect 9148 -29854 9756 -24364
rect 9148 -29964 9213 -29854
rect 9298 -29856 9539 -29854
rect 9298 -29964 9372 -29856
rect 9148 -29966 9372 -29964
rect 9457 -29964 9539 -29856
rect 9624 -29964 9756 -29854
rect 9457 -29966 9756 -29964
rect 9148 -30006 9756 -29966
rect 10594 -32424 10693 -21371
rect 10761 -23692 10827 -20814
rect 13689 -21245 13842 -21215
rect 13689 -21350 13712 -21245
rect 13814 -21350 13842 -21245
rect 13689 -21398 13842 -21350
rect 13704 -21934 13823 -21398
rect 14122 -22024 14252 -21991
rect 14122 -22090 14157 -22024
rect 14225 -22090 14252 -22024
rect 11710 -22480 11840 -22460
rect 11710 -22580 11730 -22480
rect 11830 -22580 11840 -22480
rect 11710 -22600 11840 -22580
rect 10761 -23772 10766 -23692
rect 10762 -23792 10766 -23772
rect 10818 -23772 10827 -23692
rect 10818 -23792 10825 -23772
rect 10762 -23815 10825 -23792
rect 10924 -24031 11053 -23534
rect 10881 -24066 11105 -24031
rect 10881 -24138 10918 -24066
rect 11078 -24138 11105 -24066
rect 10881 -24205 11105 -24138
rect 10881 -24272 10920 -24205
rect 11070 -24272 11105 -24205
rect 10881 -24328 11105 -24272
rect 10881 -24395 10919 -24328
rect 11069 -24395 11105 -24328
rect 10881 -24422 11105 -24395
rect 11322 -25720 11384 -23094
rect 12213 -24268 12821 -24177
rect 12213 -24275 12403 -24268
rect 12213 -24365 12251 -24275
rect 12319 -24358 12403 -24275
rect 12471 -24270 12715 -24268
rect 12471 -24358 12555 -24270
rect 12319 -24360 12555 -24358
rect 12623 -24358 12715 -24270
rect 12783 -24358 12821 -24268
rect 12623 -24360 12821 -24358
rect 12319 -24365 12821 -24360
rect 11310 -25740 11420 -25720
rect 11310 -25800 11330 -25740
rect 11400 -25800 11420 -25740
rect 11310 -25820 11420 -25800
rect 12213 -29770 12821 -24365
rect 12213 -29781 12389 -29770
rect 12213 -29871 12243 -29781
rect 12311 -29860 12389 -29781
rect 12457 -29775 12821 -29770
rect 12457 -29860 12543 -29775
rect 12311 -29865 12543 -29860
rect 12611 -29865 12700 -29775
rect 12768 -29865 12821 -29775
rect 12311 -29871 12821 -29865
rect 12213 -29941 12821 -29871
rect 12213 -29952 12383 -29941
rect 12213 -30042 12229 -29952
rect 12297 -30031 12383 -29952
rect 12451 -29946 12821 -29941
rect 12451 -30031 12545 -29946
rect 12297 -30036 12545 -30031
rect 12613 -29954 12821 -29946
rect 12613 -30036 12708 -29954
rect 12297 -30042 12708 -30036
rect 12213 -30044 12708 -30042
rect 12776 -30044 12821 -29954
rect 12213 -30080 12821 -30044
rect 14122 -32424 14252 -22090
rect 14434 -22862 14676 -17203
rect 15134 -17976 15387 -17946
rect 15134 -18099 15178 -17976
rect 15340 -18099 15387 -17976
rect 15134 -18695 15387 -18099
rect 15133 -18731 15387 -18695
rect 15133 -18854 15177 -18731
rect 15339 -18854 15387 -18731
rect 15133 -18878 15387 -18854
rect 14868 -20573 15206 -20526
rect 14868 -20737 14892 -20573
rect 14980 -20737 15064 -20573
rect 15152 -20737 15206 -20573
rect 15918 -20543 16134 -20512
rect 15918 -20638 15936 -20543
rect 15988 -20545 16134 -20543
rect 15988 -20638 16040 -20545
rect 15918 -20640 16040 -20638
rect 16092 -20640 16134 -20545
rect 17288 -20543 17469 -20507
rect 17288 -20599 17299 -20543
rect 17355 -20599 17405 -20543
rect 17461 -20599 17469 -20543
rect 26633 -20554 26737 -16435
rect 28896 -17834 29195 -13299
rect 42743 -13603 43028 -13576
rect 42743 -13683 42760 -13603
rect 42838 -13606 43028 -13603
rect 42838 -13683 42938 -13606
rect 42743 -13686 42938 -13683
rect 43016 -13686 43028 -13606
rect 42743 -13738 43028 -13686
rect 42743 -13740 42933 -13738
rect 42743 -13820 42759 -13740
rect 42837 -13818 42933 -13740
rect 43011 -13818 43028 -13738
rect 42837 -13820 43028 -13818
rect 42743 -13835 43028 -13820
rect 37186 -17379 37322 -17362
rect 37186 -17498 37198 -17379
rect 37313 -17498 37322 -17379
rect 37186 -17516 37322 -17498
rect 29262 -18374 29419 -18360
rect 29262 -18461 29275 -18374
rect 29368 -18461 29419 -18374
rect 29262 -18466 29419 -18461
rect 31439 -18485 31925 -18462
rect 31439 -18546 31466 -18485
rect 31528 -18546 31925 -18485
rect 31439 -18568 31925 -18546
rect 31819 -18681 31925 -18568
rect 38254 -18693 38379 -18678
rect 38254 -18746 38290 -18693
rect 38343 -18746 38379 -18693
rect 17288 -20623 17469 -20599
rect 25555 -20579 25636 -20577
rect 15918 -20668 16134 -20640
rect 25555 -20635 25568 -20579
rect 25624 -20635 25636 -20579
rect 25555 -20661 25636 -20635
rect 26633 -20627 26645 -20554
rect 26723 -20627 26737 -20554
rect 14868 -20758 15206 -20737
rect 14425 -22918 14516 -22862
rect 14622 -22918 14693 -22862
rect 14425 -22972 14693 -22918
rect 14425 -23061 14445 -22972
rect 14521 -23061 14604 -22972
rect 14680 -23061 14693 -22972
rect 14425 -23079 14693 -23061
rect 14895 -32424 15156 -20758
rect 15922 -26190 16129 -20668
rect 21126 -20747 21230 -20738
rect 21126 -20815 21142 -20747
rect 21216 -20815 21230 -20747
rect 21126 -20827 21230 -20815
rect 22484 -20753 22562 -20742
rect 22484 -20825 22493 -20753
rect 22553 -20825 22562 -20753
rect 22484 -20836 22562 -20825
rect 26125 -22387 26235 -22364
rect 26125 -22459 26145 -22387
rect 26210 -22459 26235 -22387
rect 26125 -22483 26235 -22459
rect 20366 -24017 20607 -23975
rect 20366 -24021 20505 -24017
rect 20366 -24089 20383 -24021
rect 20444 -24085 20505 -24021
rect 20566 -24085 20607 -24017
rect 20444 -24089 20607 -24085
rect 20366 -29937 20607 -24089
rect 20366 -29939 20507 -29937
rect 20366 -30008 20376 -29939
rect 20441 -30006 20507 -29939
rect 20572 -30006 20607 -29937
rect 21089 -24020 21330 -23976
rect 21089 -24023 21244 -24020
rect 21089 -24091 21110 -24023
rect 21171 -24088 21244 -24023
rect 21305 -24088 21330 -24020
rect 21171 -24091 21330 -24088
rect 21089 -29755 21330 -24091
rect 21089 -29759 21249 -29755
rect 21089 -29827 21109 -29759
rect 21170 -29823 21249 -29759
rect 21310 -29823 21330 -29755
rect 21170 -29827 21330 -29823
rect 21089 -29888 21330 -29827
rect 21089 -29892 21249 -29888
rect 21089 -29960 21107 -29892
rect 21168 -29956 21249 -29892
rect 21310 -29956 21330 -29888
rect 21168 -29960 21330 -29956
rect 21089 -29986 21330 -29960
rect 21702 -24028 21943 -23975
rect 21702 -24096 21729 -24028
rect 21790 -24029 21943 -24028
rect 21790 -24096 21843 -24029
rect 21702 -24097 21843 -24096
rect 21902 -24097 21943 -24029
rect 21702 -29748 21943 -24097
rect 26633 -25295 26737 -20627
rect 27332 -22384 27485 -22362
rect 27332 -22449 27375 -22384
rect 27448 -22449 27485 -22384
rect 21702 -29815 21790 -29748
rect 21853 -29815 21943 -29748
rect 21702 -29867 21943 -29815
rect 21702 -29869 21865 -29867
rect 21702 -29937 21717 -29869
rect 21778 -29935 21865 -29869
rect 21926 -29935 21943 -29867
rect 21778 -29937 21943 -29935
rect 21702 -29968 21943 -29937
rect 20441 -30008 20607 -30006
rect 20366 -30029 20607 -30008
rect 27332 -32424 27485 -22449
rect 28180 -24405 28351 -20250
rect 30936 -20285 31027 -20180
rect 28151 -24445 28391 -24405
rect 28151 -24606 28195 -24445
rect 28352 -24606 28391 -24445
rect 28151 -24639 28391 -24606
rect 30865 -32424 31027 -20285
rect 38254 -22811 38379 -18746
rect 42786 -19224 42999 -13835
rect 43657 -17006 43871 -16967
rect 43657 -17128 43704 -17006
rect 43788 -17128 43871 -17006
rect 43657 -17879 43871 -17128
rect 43657 -17946 43687 -17879
rect 43839 -17946 43871 -17879
rect 43657 -17973 43871 -17946
rect 45110 -18087 45368 -12457
rect 47173 -16438 47482 -2182
rect 47766 -6601 48171 -6585
rect 47766 -6681 47793 -6601
rect 47871 -6604 48171 -6601
rect 47871 -6681 47971 -6604
rect 47766 -6684 47971 -6681
rect 48049 -6684 48171 -6604
rect 47766 -6736 48171 -6684
rect 47766 -6738 47966 -6736
rect 47766 -6818 47792 -6738
rect 47870 -6816 47966 -6738
rect 48044 -6816 48171 -6736
rect 47870 -6818 48171 -6816
rect 47766 -6880 48171 -6818
rect 47769 -13488 48171 -6880
rect 47761 -13575 48171 -13488
rect 47761 -13655 47809 -13575
rect 47887 -13578 48171 -13575
rect 47887 -13655 47987 -13578
rect 47761 -13658 47987 -13655
rect 48065 -13658 48171 -13578
rect 47761 -13710 48171 -13658
rect 47761 -13712 47982 -13710
rect 47761 -13792 47808 -13712
rect 47886 -13790 47982 -13712
rect 48060 -13790 48171 -13710
rect 47886 -13792 48171 -13790
rect 47761 -13851 48171 -13792
rect 47769 -13854 48171 -13851
rect 47835 -13863 48048 -13854
rect 47139 -16476 47501 -16438
rect 47139 -16480 47356 -16476
rect 47139 -16554 47214 -16480
rect 47292 -16550 47356 -16480
rect 47434 -16550 47501 -16476
rect 47292 -16554 47501 -16550
rect 47139 -16607 47501 -16554
rect 47139 -16618 47357 -16607
rect 47139 -16692 47224 -16618
rect 47302 -16681 47357 -16618
rect 47435 -16681 47501 -16607
rect 47302 -16692 47501 -16681
rect 47139 -16766 47501 -16692
rect 48489 -17331 48958 23857
rect 56364 -244 56594 -229
rect 56356 -256 56594 -244
rect 56356 -275 56595 -256
rect 56356 -327 56382 -275
rect 56434 -327 56501 -275
rect 56553 -327 56595 -275
rect 56356 -379 56595 -327
rect 56356 -381 56496 -379
rect 56356 -433 56379 -381
rect 56431 -431 56496 -381
rect 56548 -431 56595 -379
rect 56431 -433 56595 -431
rect 56356 -446 56595 -433
rect 56356 -447 56594 -446
rect 49363 -4142 49615 -4114
rect 49363 -4143 49506 -4142
rect 49363 -4205 49385 -4143
rect 49451 -4201 49506 -4143
rect 49569 -4201 49615 -4142
rect 49451 -4205 49615 -4201
rect 49363 -4256 49615 -4205
rect 49363 -4261 49514 -4256
rect 49363 -4323 49380 -4261
rect 49446 -4315 49514 -4261
rect 49577 -4315 49615 -4256
rect 49446 -4323 49615 -4315
rect 49363 -4338 49615 -4323
rect 49366 -14201 49597 -4338
rect 56356 -4873 56586 -447
rect 56356 -4942 56930 -4873
rect 56353 -4961 56930 -4942
rect 56353 -5013 56374 -4961
rect 56426 -5013 56493 -4961
rect 56545 -5013 56930 -4961
rect 56353 -5065 56930 -5013
rect 56353 -5067 56488 -5065
rect 56353 -5119 56371 -5067
rect 56423 -5117 56488 -5067
rect 56540 -5103 56930 -5065
rect 56540 -5117 56587 -5103
rect 56423 -5119 56587 -5117
rect 56353 -5132 56587 -5119
rect 56355 -5133 56586 -5132
rect 51603 -9255 56191 -9252
rect 51603 -9352 55881 -9255
rect 56139 -9352 56191 -9255
rect 51603 -9356 56191 -9352
rect 51603 -9970 51676 -9356
rect 51603 -9973 51743 -9970
rect 51603 -9997 51764 -9973
rect 51603 -10070 51887 -9997
rect 49366 -14203 49513 -14201
rect 49366 -14257 49382 -14203
rect 49460 -14255 49513 -14203
rect 49591 -14255 49597 -14201
rect 49460 -14257 49597 -14255
rect 49366 -14308 49597 -14257
rect 49366 -14313 49516 -14308
rect 49366 -14389 49384 -14313
rect 49453 -14384 49516 -14313
rect 49585 -14384 49597 -14308
rect 49453 -14389 49597 -14384
rect 49366 -14452 49597 -14389
rect 49366 -14457 49514 -14452
rect 49366 -14533 49381 -14457
rect 49450 -14528 49514 -14457
rect 49583 -14528 49597 -14452
rect 49450 -14533 49597 -14528
rect 49366 -14547 49597 -14533
rect 49394 -14755 49740 -14739
rect 49394 -14761 49618 -14755
rect 49394 -14839 49422 -14761
rect 49506 -14833 49618 -14761
rect 49702 -14833 49740 -14755
rect 49506 -14839 49740 -14833
rect 49394 -14900 49740 -14839
rect 49394 -14908 49616 -14900
rect 49394 -14986 49424 -14908
rect 49508 -14978 49616 -14908
rect 49700 -14978 49740 -14900
rect 49508 -14986 49740 -14978
rect 49394 -15006 49740 -14986
rect 49422 -16120 49680 -15006
rect 49422 -16290 49440 -16120
rect 49580 -16290 49680 -16120
rect 49422 -16333 49680 -16290
rect 49648 -17009 49898 -16985
rect 49648 -17013 49814 -17009
rect 49648 -17087 49672 -17013
rect 49750 -17083 49814 -17013
rect 49892 -17031 49898 -17009
rect 49892 -17083 54506 -17031
rect 49750 -17087 54506 -17083
rect 49648 -17140 54506 -17087
rect 49648 -17151 49815 -17140
rect 49648 -17225 49682 -17151
rect 49760 -17214 49815 -17151
rect 49893 -17210 54506 -17140
rect 49893 -17214 49898 -17210
rect 49760 -17225 49898 -17214
rect 49648 -17255 49898 -17225
rect 48489 -17332 48728 -17331
rect 48489 -17334 48622 -17332
rect 48489 -17387 48511 -17334
rect 48563 -17385 48622 -17334
rect 48674 -17384 48728 -17332
rect 48780 -17332 48958 -17331
rect 48780 -17384 48846 -17332
rect 48674 -17385 48846 -17384
rect 48898 -17369 48958 -17332
rect 48898 -17385 48957 -17369
rect 48563 -17387 48957 -17385
rect 48489 -17403 48957 -17387
rect 45110 -18229 45164 -18087
rect 45316 -18229 45368 -18087
rect 45110 -18250 45368 -18229
rect 49884 -18633 50008 -18627
rect 49884 -18690 49905 -18633
rect 49979 -18690 50008 -18633
rect 49884 -18719 50008 -18690
rect 42756 -19290 43047 -19224
rect 42756 -19292 42935 -19290
rect 42756 -19364 42792 -19292
rect 42860 -19362 42935 -19292
rect 43003 -19362 43047 -19290
rect 42860 -19364 43047 -19362
rect 42756 -19400 43047 -19364
rect 42755 -19456 43047 -19400
rect 42755 -19528 42789 -19456
rect 42857 -19457 43047 -19456
rect 42857 -19528 42933 -19457
rect 42755 -19529 42933 -19528
rect 43001 -19529 43047 -19457
rect 42755 -19559 43047 -19529
rect 41604 -21120 41733 -21098
rect 41604 -21182 41640 -21120
rect 41702 -21182 41733 -21120
rect 38254 -22894 38275 -22811
rect 38353 -22894 38379 -22811
rect 38254 -22920 38379 -22894
rect 39010 -22791 39138 -22773
rect 39010 -22895 39032 -22791
rect 39121 -22895 39138 -22791
rect 32062 -25334 32223 -25305
rect 32062 -25447 32080 -25334
rect 32192 -25447 32223 -25334
rect 32062 -25471 32223 -25447
rect 32067 -32424 32219 -25471
rect 33741 -25631 33977 -25593
rect 33741 -25685 33766 -25631
rect 33819 -25685 33889 -25631
rect 33942 -25685 33977 -25631
rect 33741 -29805 33977 -25685
rect 33741 -29806 33885 -29805
rect 33741 -29864 33774 -29806
rect 33828 -29863 33885 -29806
rect 33939 -29863 33977 -29805
rect 33828 -29864 33977 -29863
rect 33741 -29893 33977 -29864
rect 35196 -25635 35432 -25581
rect 35196 -25638 35352 -25635
rect 35196 -25692 35210 -25638
rect 35263 -25689 35352 -25638
rect 35405 -25689 35432 -25635
rect 35263 -25692 35432 -25689
rect 35196 -29793 35432 -25692
rect 35196 -29851 35213 -29793
rect 35267 -29794 35432 -29793
rect 35267 -29851 35320 -29794
rect 35196 -29852 35320 -29851
rect 35374 -29852 35432 -29794
rect 35196 -29881 35432 -29852
rect 36549 -25617 36785 -25605
rect 36549 -25671 36586 -25617
rect 36639 -25618 36785 -25617
rect 36639 -25671 36703 -25618
rect 36549 -25672 36703 -25671
rect 36756 -25672 36785 -25618
rect 36549 -29809 36785 -25672
rect 36549 -29867 36560 -29809
rect 36614 -29867 36706 -29809
rect 36760 -29867 36785 -29809
rect 36549 -29905 36785 -29867
rect 37983 -25618 38219 -25599
rect 37983 -25620 38117 -25618
rect 37983 -25674 37992 -25620
rect 38045 -25672 38117 -25620
rect 38170 -25672 38219 -25618
rect 38045 -25674 38219 -25672
rect 37983 -29579 38219 -25674
rect 37983 -29583 38125 -29579
rect 37983 -29642 38004 -29583
rect 38064 -29638 38125 -29583
rect 38185 -29638 38219 -29579
rect 38064 -29642 38219 -29638
rect 37983 -29694 38219 -29642
rect 37983 -29753 38005 -29694
rect 38065 -29695 38219 -29694
rect 38065 -29753 38129 -29695
rect 37983 -29754 38129 -29753
rect 38189 -29754 38219 -29695
rect 37983 -29807 38219 -29754
rect 37983 -29866 38007 -29807
rect 38067 -29808 38219 -29807
rect 38067 -29866 38130 -29808
rect 38184 -29866 38219 -29808
rect 37983 -29908 38219 -29866
rect 39010 -32424 39138 -22895
rect 41604 -32424 41733 -21182
rect 49884 -22841 50006 -18719
rect 54327 -19359 54506 -17210
rect 54327 -19361 54444 -19359
rect 54327 -19414 54340 -19361
rect 54392 -19412 54444 -19361
rect 54496 -19412 54506 -19359
rect 54392 -19414 54506 -19412
rect 54327 -19427 54506 -19414
rect 53211 -21056 53348 -21047
rect 53211 -21119 53259 -21056
rect 53321 -21119 53348 -21056
rect 49878 -22879 50019 -22841
rect 49878 -22989 49907 -22879
rect 49996 -22989 50019 -22879
rect 49878 -23019 50019 -22989
rect 50505 -22880 50644 -22850
rect 50505 -22990 50534 -22880
rect 50623 -22990 50644 -22880
rect 43669 -25319 43830 -25305
rect 43669 -25456 43694 -25319
rect 43819 -25456 43830 -25319
rect 43669 -25473 43830 -25456
rect 44584 -25539 44820 -25520
rect 44584 -25602 44605 -25539
rect 44659 -25540 44820 -25539
rect 44659 -25602 44715 -25540
rect 44584 -25603 44715 -25602
rect 44769 -25603 44820 -25540
rect 44584 -29801 44820 -25603
rect 44584 -29864 44612 -29801
rect 44666 -29804 44820 -29801
rect 44666 -29864 44746 -29804
rect 44584 -29867 44746 -29864
rect 44800 -29867 44820 -29804
rect 44584 -29906 44820 -29867
rect 45800 -25556 46036 -25535
rect 45800 -25619 45823 -25556
rect 45877 -25619 45954 -25556
rect 46008 -25619 46036 -25556
rect 45800 -29793 46036 -25619
rect 45800 -29810 45839 -29793
rect 45893 -29794 46036 -29793
rect 45800 -29873 45820 -29810
rect 45893 -29851 45946 -29794
rect 46000 -29807 46036 -29794
rect 45874 -29852 45946 -29851
rect 45874 -29870 45960 -29852
rect 46014 -29870 46036 -29807
rect 45874 -29873 46036 -29870
rect 45800 -29921 46036 -29873
rect 46930 -25556 47166 -25523
rect 46930 -25563 47077 -25556
rect 46930 -25626 46948 -25563
rect 47002 -25619 47077 -25563
rect 47131 -25619 47166 -25556
rect 47002 -25626 47166 -25619
rect 46930 -29792 47166 -25626
rect 46930 -29860 46955 -29792
rect 47010 -29796 47166 -29792
rect 47010 -29859 47082 -29796
rect 47136 -29859 47166 -29796
rect 47010 -29860 47166 -29859
rect 46930 -29914 47166 -29860
rect 47939 -25557 48175 -25475
rect 47939 -25560 48100 -25557
rect 47939 -25623 47967 -25560
rect 48021 -25620 48100 -25560
rect 48154 -25620 48175 -25557
rect 48021 -25623 48175 -25620
rect 47939 -29770 48175 -25623
rect 47939 -29833 47957 -29770
rect 48011 -29833 48094 -29770
rect 48148 -29833 48175 -29770
rect 47939 -29861 48175 -29833
rect 49228 -25559 49464 -25511
rect 49228 -25560 49394 -25559
rect 49228 -25623 49256 -25560
rect 49310 -25622 49394 -25560
rect 49448 -25622 49464 -25559
rect 49310 -25623 49464 -25622
rect 49228 -29801 49464 -25623
rect 49228 -29864 49261 -29801
rect 49315 -29864 49377 -29801
rect 49431 -29864 49464 -29801
rect 49228 -29897 49464 -29864
rect 50505 -32424 50644 -22990
rect 53211 -32424 53348 -21119
rect 56702 -27061 56928 -5103
rect 56665 -27101 56938 -27061
rect 56665 -27103 56846 -27101
rect 56665 -27173 56683 -27103
rect 56771 -27171 56846 -27103
rect 56934 -27171 56938 -27101
rect 56771 -27173 56938 -27171
rect 56665 -27239 56938 -27173
rect 56665 -27244 56840 -27239
rect 56665 -27314 56680 -27244
rect 56768 -27309 56840 -27244
rect 56928 -27309 56938 -27239
rect 56768 -27314 56938 -27309
rect 56665 -27328 56938 -27314
rect 56702 -27330 56928 -27328
<< via2 >>
rect -4906 -3243 -4843 -3176
rect -3876 -4233 -3809 -4231
rect -3876 -4288 -3810 -4233
rect -3810 -4288 -3809 -4233
rect -8417 -15562 -8351 -15490
rect -8411 -18073 -8345 -18001
rect 8348 -4205 8422 -4130
rect 8483 -4204 8557 -4129
rect 8346 -4364 8420 -4289
rect 8482 -4363 8556 -4288
rect 4886 -4815 4988 -4703
rect 7245 -6997 7439 -6820
rect 28957 -13299 29123 -13122
rect 8343 -18796 8344 -18724
rect 8344 -18796 8398 -18724
rect 8398 -18796 8399 -18724
rect 8452 -18795 8508 -18723
rect 11743 -18733 11806 -18729
rect 11743 -18796 11747 -18733
rect 11747 -18796 11802 -18733
rect 11802 -18796 11806 -18733
rect 11743 -18800 11806 -18796
rect 11730 -22580 11830 -22480
rect 15177 -18854 15339 -18731
rect 17299 -20544 17355 -20543
rect 17299 -20598 17353 -20544
rect 17353 -20598 17355 -20544
rect 17299 -20599 17355 -20598
rect 17405 -20545 17461 -20543
rect 17405 -20599 17459 -20545
rect 17459 -20599 17461 -20545
rect 37198 -17388 37313 -17379
rect 37198 -17492 37209 -17388
rect 37209 -17492 37308 -17388
rect 37308 -17492 37313 -17388
rect 37198 -17498 37313 -17492
rect 29275 -18381 29368 -18374
rect 29275 -18455 29284 -18381
rect 29284 -18455 29359 -18381
rect 29359 -18455 29368 -18381
rect 29275 -18461 29368 -18455
rect 25568 -20580 25624 -20579
rect 25568 -20632 25572 -20580
rect 25572 -20632 25624 -20580
rect 25568 -20635 25624 -20632
rect 21142 -20750 21216 -20747
rect 21142 -20815 21213 -20750
rect 21213 -20815 21216 -20750
rect 22493 -20825 22553 -20753
rect 26145 -22396 26210 -22387
rect 26145 -22456 26152 -22396
rect 26152 -22456 26205 -22396
rect 26205 -22456 26210 -22396
rect 26145 -22459 26210 -22456
rect 27375 -22449 27448 -22384
rect 45164 -18229 45316 -18087
rect 41648 -19304 41707 -19244
rect 41640 -21182 41702 -21120
rect 32080 -25447 32192 -25334
rect 53259 -19256 53315 -19199
rect 53259 -21119 53321 -21056
rect 43694 -25320 43819 -25319
rect 43694 -25445 43698 -25320
rect 43698 -25445 43816 -25320
rect 43816 -25445 43819 -25320
rect 43694 -25456 43819 -25445
<< metal3 >>
rect -4924 -3176 -4822 -3160
rect -4924 -3243 -4906 -3176
rect -4843 -3243 -4822 -3176
rect -4924 -3257 -4822 -3243
rect -4924 -4743 -4823 -3257
rect 8335 -4129 8569 -4093
rect 8335 -4130 8483 -4129
rect 8335 -4144 8348 -4130
rect -2768 -4205 8348 -4144
rect 8422 -4204 8483 -4130
rect 8557 -4204 8569 -4129
rect 8422 -4205 8569 -4204
rect -3889 -4227 -3795 -4223
rect -2768 -4227 8569 -4205
rect -3889 -4231 8569 -4227
rect -3889 -4288 -3876 -4231
rect -3809 -4288 8569 -4231
rect -3889 -4289 8482 -4288
rect -3889 -4307 8346 -4289
rect -3886 -4314 8346 -4307
rect 8335 -4364 8346 -4314
rect 8420 -4363 8482 -4289
rect 8556 -4363 8569 -4288
rect 8420 -4364 8569 -4363
rect 8335 -4376 8569 -4364
rect 4832 -4703 5040 -4657
rect 4832 -4743 4886 -4703
rect -4924 -4815 4886 -4743
rect 4988 -4815 5040 -4703
rect -4924 -4844 5040 -4815
rect -4924 -4848 -4823 -4844
rect 4832 -4878 5040 -4844
rect 7183 -6820 7485 -6777
rect 7183 -6827 7245 -6820
rect -6357 -6997 7245 -6827
rect 7439 -6997 7485 -6820
rect -6357 -7018 7485 -6997
rect -6357 -11485 -6275 -7018
rect 7183 -7086 7485 -7018
rect -8459 -15490 -8278 -15482
rect -8459 -15562 -8417 -15490
rect -8351 -15562 -8278 -15490
rect -8459 -18001 -8278 -15562
rect 29261 -17379 37323 -17362
rect 29261 -17498 37198 -17379
rect 37313 -17498 37323 -17379
rect 29261 -17517 37323 -17498
rect -8459 -18073 -8411 -18001
rect -8345 -18073 -8278 -18001
rect -8459 -18108 -8278 -18073
rect 29262 -18360 29417 -17517
rect 45110 -18087 45368 -18073
rect 45110 -18106 45164 -18087
rect 43674 -18229 45164 -18106
rect 45316 -18229 45368 -18087
rect 43674 -18249 45368 -18229
rect 29262 -18374 29419 -18360
rect 29262 -18461 29275 -18374
rect 29368 -18461 29419 -18374
rect 29262 -18466 29419 -18461
rect 8328 -18723 11815 -18700
rect 8328 -18724 8452 -18723
rect 8328 -18796 8343 -18724
rect 8399 -18795 8452 -18724
rect 8508 -18729 11815 -18723
rect 8508 -18795 11743 -18729
rect 8399 -18796 11743 -18795
rect 8328 -18800 11743 -18796
rect 11806 -18800 11815 -18729
rect 8328 -18814 11815 -18800
rect 15133 -18731 15384 -18695
rect 15133 -18854 15177 -18731
rect 15339 -18740 15384 -18731
rect 15339 -18854 19551 -18740
rect 15133 -18874 19551 -18854
rect 15133 -18878 15384 -18874
rect 41628 -19244 41718 -19237
rect 41628 -19304 41648 -19244
rect 41707 -19304 41718 -19244
rect 17288 -20525 17469 -20507
rect 20068 -20525 20157 -20524
rect 17288 -20543 20157 -20525
rect 17288 -20599 17299 -20543
rect 17355 -20599 17405 -20543
rect 17461 -20599 20157 -20543
rect 25555 -20579 25636 -20577
rect 25555 -20580 25568 -20579
rect 17288 -20614 20157 -20599
rect 17288 -20623 17469 -20614
rect 20068 -20738 20157 -20614
rect 23255 -20635 25568 -20580
rect 25624 -20635 25636 -20579
rect 23255 -20661 25636 -20635
rect 20068 -20747 21230 -20738
rect 23255 -20742 23336 -20661
rect 20068 -20815 21142 -20747
rect 21216 -20815 21230 -20747
rect 20068 -20827 21230 -20815
rect 22424 -20753 23336 -20742
rect 22424 -20823 22493 -20753
rect 22484 -20825 22493 -20823
rect 22553 -20823 23336 -20753
rect 22553 -20825 22562 -20823
rect 22484 -20836 22562 -20825
rect 41628 -21120 41718 -19304
rect 43674 -20502 43756 -18249
rect 45110 -18250 45368 -18249
rect 53238 -19199 53328 -19187
rect 53238 -19256 53259 -19199
rect 53315 -19256 53328 -19199
rect 53238 -19271 53328 -19256
rect 41628 -21182 41640 -21120
rect 41702 -21182 41718 -21120
rect 53244 -21056 53328 -19271
rect 53244 -21119 53259 -21056
rect 53321 -21119 53328 -21056
rect 53244 -21139 53328 -21119
rect 41628 -21209 41718 -21182
rect 27332 -22364 27485 -22362
rect 26125 -22384 27485 -22364
rect 26125 -22387 27375 -22384
rect 26125 -22459 26145 -22387
rect 26210 -22449 27375 -22387
rect 27448 -22449 27485 -22384
rect 26210 -22459 27485 -22449
rect 11710 -22463 11840 -22460
rect 11710 -22480 17158 -22463
rect 11710 -22580 11730 -22480
rect 11830 -22580 17158 -22480
rect 26125 -22482 27485 -22459
rect 26125 -22483 27452 -22482
rect 11710 -22597 17158 -22580
rect 11710 -22600 11840 -22597
rect 32062 -25319 43832 -25305
rect 32062 -25334 43694 -25319
rect 32062 -25447 32080 -25334
rect 32192 -25447 43694 -25334
rect 32062 -25456 43694 -25447
rect 43819 -25456 43832 -25319
rect 32062 -25471 43832 -25456
rect 43669 -25474 43830 -25471
<< metal4 >>
rect -27683 6835 -27616 6959
<< metal5 >>
rect -33413 6835 -33201 7200
use a2x1mux_mag  a2x1mux_mag_0
timestamp 1714554054
transform 1 0 11521 0 1 -22420
box -615 -1160 2414 924
use A_MUX_mag  A_MUX_mag_0
timestamp 1714138925
transform 1 0 10363 0 1 -20243
box -285 -452 3979 2227
use A_MUX_mag  A_MUX_mag_1
timestamp 1714138925
transform 1 0 27205 0 1 -19948
box -285 -452 3979 2227
use CP_mag  CP_mag_0
timestamp 1714559806
transform 1 0 8022 0 1 -22735
box 76 665 2629 1839
use Current_Mirror_Top  Current_Mirror_Top_0
timestamp 1714139039
transform 1 0 51904 0 -1 -9894
box -1992 -209 4486 7070
use Feedback_Divider_mag  Feedback_Divider_mag_0
timestamp 1714559211
transform 1 0 -12035 0 1 8548
box 17773 -23960 58979 12279
use INV_2  INV_2_0
timestamp 1714126980
transform 1 0 -7671 0 1 -27192
box 21 -485 1081 648
use INV_2  INV_2_1
timestamp 1714126980
transform 1 0 49067 0 1 -6661
box 21 -485 1081 648
use INV_2  INV_2_2
timestamp 1714126980
transform 1 0 49014 0 1 -1970
box 21 -485 1081 648
use LF_mag  LF_mag_0
timestamp 1714558529
transform 1 0 -55438 0 1 -26725
box -85 43 54977 46220
use mux_2x1_ibr  mux_2x1_ibr_0
timestamp 1714558529
transform 1 0 5862 0 1 -22468
box 0 -1051 1135 1051
use mux_2x1_ibr  mux_2x1_ibr_1
timestamp 1714558529
transform 1 0 5862 0 -1 -20366
box 0 -1051 1135 1051
use mux_2x1_ibr  mux_2x1_ibr_3
timestamp 1714558529
transform 1 0 -2960 0 1 -23349
box 0 -1051 1135 1051
use mux_2x1_ibr  mux_2x1_ibr_4
timestamp 1714558529
transform 1 0 -2955 0 1 -21250
box 0 -1051 1135 1051
use mux_4x1_ibr  mux_4x1_ibr_0
timestamp 1714558529
transform 1 0 -4968 0 1 -4738
box -1194 5 2193 2107
use Output_Div_Mag  Output_Div_Mag_0
timestamp 1714558796
transform 1 0 32258 0 1 -18132
box -638 -7578 10327 786
use Output_Div_Mag  Output_Div_Mag_1
timestamp 1714558796
transform 1 0 43867 0 1 -18086
box -638 -7578 10327 786
use PFD_layout  PFD_layout_0
timestamp 1714557138
transform 1 0 -1040 0 1 -24269
box -555 -148 6587 5567
use pre_div_mag  pre_div_mag_0
timestamp 1714558796
transform 1 0 -6164 0 1 -8963
box -638 -7578 10327 786
use Tappered_Buffer  Tappered_Buffer_0
timestamp 1714490790
transform 1 0 50329 0 1 -1131
box -161 -3147 5956 950
use Tappered_Buffer  Tappered_Buffer_1
timestamp 1714490790
transform 1 0 -5513 0 1 -26185
box -161 -3147 5956 950
use Tappered_Buffer  Tappered_Buffer_2
timestamp 1714490790
transform 1 0 50366 0 1 -5883
box -161 -3147 5956 950
use VCO_mag  VCO_mag_0
timestamp 1714543819
transform 1 0 16391 0 1 -20374
box -5 -3738 10083 3421
<< labels >>
flabel via1 56133 -9304 56133 -9304 0 FreeSans 1600 0 0 0 Iref
port 47 nsew
flabel metal2 8123 -20623 8123 -20623 0 FreeSans 960 0 0 0 IPD_
port 10 nsew
flabel metal1 -714 -31035 -714 -31035 0 FreeSans 2400 0 0 0 VSS
port 44 nsew
flabel metal1 -3118 24923 -3118 24923 0 FreeSans 2400 0 0 0 VDD
port 45 nsew
flabel metal2 7884 -20465 7884 -20465 0 FreeSans 960 0 0 0 IPD+
port 9 nsew
flabel metal2 15994 -25870 15994 -25870 0 FreeSans 1600 0 0 0 VCO_op_bar
port 22 nsew
flabel space -55858 -32154 56977 26259 0 FreeSans 1600 0 0 0 Test_output
port 48 nsew
flabel metal1 56473 -7353 56473 -7353 0 FreeSans 1600 0 0 0 Output1
port 50 nsew
flabel metal1 56617 -2611 56617 -2611 0 FreeSans 1600 0 0 0 Output2
port 51 nsew
flabel metal1 56798 -318 56798 -318 0 FreeSans 1600 0 0 0 VDD_BUFF
port 52 nsew
flabel metal1 56594 23367 56594 23367 0 FreeSans 1600 0 0 0 F2
port 53 nsew
flabel metal1 56594 23129 56594 23129 0 FreeSans 1600 0 0 0 F1
port 54 nsew
flabel metal1 56566 22830 56566 22830 0 FreeSans 1600 0 0 0 F0
port 55 nsew
flabel metal1 56569 22449 56569 22449 0 FreeSans 1600 0 0 0 T0
port 56 nsew
flabel metal1 56543 22249 56543 22249 0 FreeSans 1600 0 0 0 T1
port 57 nsew
flabel metal1 -10170 5390 -10170 5390 0 FreeSans 1600 0 0 0 LP_RES_CAP_INT
port 58 nsew
flabel metal1 10850 21920 10850 21920 0 FreeSans 1600 0 0 0 Vdiv_FB_MUX_INT
port 59 nsew
flabel metal3 15702 -18824 15702 -18824 0 FreeSans 1600 0 0 0 VCNT_MUX_INT
port 60 nsew
flabel metal1 7251 -16421 7251 -16421 0 FreeSans 1600 0 0 0 VSS_INT_1
port 61 nsew
flabel metal1 45658 -14304 45658 -14304 0 FreeSans 1600 0 0 0 VSS_INT_2
port 62 nsew
flabel metal1 49954 -858 49954 -858 0 FreeSans 1600 0 0 0 VDD_BUFF_INT_1
port 63 nsew
flabel metal1 50126 -5696 50126 -5696 0 FreeSans 1600 0 0 0 VDD_BUFF_INT_2
port 64 nsew
flabel metal1 -5662 -25395 -5662 -25395 0 FreeSans 1600 0 0 0 VDD_BUFF_INT_3
port 65 nsew
flabel metal1 -6237 -27229 -6237 -27229 0 FreeSans 1600 0 0 0 INV_BUFF_INT_3
port 66 nsew
flabel metal1 50187 -6711 50187 -6711 0 FreeSans 1600 0 0 0 INV_BUFF_INT_2
port 67 nsew
flabel metal1 50144 -1987 50144 -1987 0 FreeSans 1600 0 0 0 INV_BUFF_INT_1
port 68 nsew
flabel metal1 49787 -8432 49787 -8432 0 FreeSans 1600 0 0 0 VSS_BUFF_INT_5
port 69 nsew
flabel metal1 44684 -17157 44684 -17157 0 FreeSans 1600 0 0 0 VDD_INT_5
port 70 nsew
flabel metal1 47842 -2099 47842 -2099 0 FreeSans 1600 0 0 0 Output_2_INT
port 71 nsew
flabel metal2 47863 -7237 47863 -7237 0 FreeSans 1600 0 0 0 Output_1_INT
port 72 nsew
flabel metal2 -8402 -24118 -8402 -24118 0 FreeSans 1600 0 0 0 Test_Output_INT
port 73 nsew
flabel metal2 -3143 -19495 -3143 -19495 0 FreeSans 1600 0 0 0 PRE_DIV_OP_INT
port 74 nsew
flabel metal1 -1694 -22894 -1694 -22894 0 FreeSans 1600 0 0 0 PFD_Vdiv_IN_INT
port 78 nsew
flabel metal1 -1688 -23411 -1688 -23411 0 FreeSans 1600 0 0 0 VSS_INT_8
port 80 nsew
flabel metal2 769 -15584 769 -15584 0 FreeSans 1600 0 0 0 VDD_INT_8
port 81 nsew
flabel metal1 6755 -18872 6755 -18872 0 FreeSans 1600 0 0 0 VDD_INT_9
port 82 nsew
flabel metal1 5488 -20853 5488 -20853 0 FreeSans 1600 0 0 0 PU_INT
port 83 nsew
flabel metal1 5651 -22897 5651 -22897 0 FreeSans 1600 0 0 0 PD_INT
port 84 nsew
flabel metal1 7276 -21443 7276 -21443 0 FreeSans 1600 0 0 0 PU_MUX_OP_INT
port 86 nsew
flabel metal1 7192 -21874 7192 -21874 0 FreeSans 1600 0 0 0 PD_MUX_OP_INT
port 87 nsew
flabel metal1 7983 -22576 7983 -22576 0 FreeSans 1600 0 0 0 VDD_INT_10
port 88 nsew
flabel metal1 31338 -18537 31338 -18537 0 FreeSans 1600 0 0 0 VSS_INT_11
port 89 nsew
flabel metal3 30164 -17424 30164 -17424 0 FreeSans 1600 0 0 0 VDD_INT_13
port 90 nsew
flabel metal2 26682 -24928 26682 -24928 0 FreeSans 1600 0 0 0 VCO_op
port 21 nsew
flabel metal2 29022 -13843 29022 -13843 0 FreeSans 1600 0 0 0 CLK_FB_IN_INT
flabel metal2 -7762 -32291 -7762 -32291 0 FreeSans 1600 0 0 0 P1
port 91 nsew
flabel metal2 -7216 -32322 -7216 -32322 0 FreeSans 1600 0 0 0 P0
port 94 nsew
flabel metal2 -6778 -32322 -6778 -32322 0 FreeSans 1600 0 0 0 Vref
port 95 nsew
flabel metal2 4375 -32388 4375 -32388 0 FreeSans 1600 0 0 0 Vdiv_test
port 96 nsew
flabel metal2 4568 -32244 4568 -32244 0 FreeSans 1600 0 0 0 S0
port 97 nsew
flabel metal2 6217 -32391 6217 -32391 0 FreeSans 1600 0 0 0 S1
port 98 nsew
flabel metal2 6557 -32335 6557 -32335 0 FreeSans 1600 0 0 0 S2
port 99 nsew
flabel metal2 7138 -32063 7138 -32063 0 FreeSans 1600 0 0 0 PD_test
port 100 nsew
flabel metal2 7382 -32414 7382 -32414 0 FreeSans 1600 0 0 0 PU_test
port 101 nsew
flabel metal2 10639 -32356 10639 -32356 0 FreeSans 1600 0 0 0 LP_op_test
port 102 nsew
flabel metal2 14182 -32334 14182 -32334 0 FreeSans 1600 0 0 0 LP_ext
port 103 nsew
flabel metal2 14983 -32048 14983 -32048 0 FreeSans 1600 0 0 0 vcntl_test
port 104 nsew
flabel metal2 27401 -32380 27401 -32380 0 FreeSans 1600 0 0 0 VDD_VCO
port 105 nsew
flabel metal2 30946 -32323 30946 -32323 0 FreeSans 1600 0 0 0 Vo_test
port 106 nsew
flabel metal2 32147 -32345 32147 -32345 0 FreeSans 1600 0 0 0 RST_DIV
port 107 nsew
flabel metal2 39088 -32345 39088 -32345 0 FreeSans 1600 0 0 0 OPA0
port 108 nsew
flabel metal2 41661 -32334 41661 -32334 0 FreeSans 1600 0 0 0 OPA1
port 109 nsew
flabel metal2 50558 -32351 50558 -32351 0 FreeSans 1600 0 0 0 OPB0
port 110 nsew
flabel metal2 53248 -32305 53248 -32305 0 FreeSans 1600 0 0 0 OPB1
port 111 nsew
flabel metal1 56943 -27772 56943 -27772 0 FreeSans 1600 0 0 0 Test_output
port 112 nsew
flabel metal1 -1686 -20341 -1686 -20341 0 FreeSans 1600 0 0 0 VDD_INT_7
port 75 nsew
flabel metal1 -1664 -21246 -1664 -21246 0 FreeSans 1600 0 0 0 VSS_INT_7
port 76 nsew
flabel metal1 -2526 -22248 -2526 -22248 0 FreeSans 1600 0 0 0 VDD_INT_8
port 77 nsew
flabel metal1 -1776 -20782 -1776 -20782 0 FreeSans 1600 0 0 0 PFD_Vref_IN_INT
port 79 nsew
<< end >>
