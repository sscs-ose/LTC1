magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -3643 2045 3643
<< psubdiff >>
rect -45 1621 45 1643
rect -45 -1621 -23 1621
rect 23 -1621 45 1621
rect -45 -1643 45 -1621
<< psubdiffcont >>
rect -23 -1621 23 1621
<< metal1 >>
rect -34 1621 34 1632
rect -34 -1621 -23 1621
rect 23 -1621 34 1621
rect -34 -1632 34 -1621
<< end >>
