magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1097 -1045 1097 1045
<< metal1 >>
rect -97 39 97 45
rect -97 -39 -91 39
rect 91 -39 97 39
rect -97 -45 97 -39
<< via1 >>
rect -91 -39 91 39
<< metal2 >>
rect -97 39 97 45
rect -97 -39 -91 39
rect 91 -39 97 39
rect -97 -45 97 -39
<< end >>
