* NGSPICE file created from Filter_magic_flat.ext - technology: gf180mcuC

.subckt Filter_magic_flat VIN_N1 VDD VSS VCM1 VIN_P1 VOUT_OPAMP_P VOUT_OPAMP_N VOUT_P
+ VOUT_N
X0 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t36 VOUT_N.t37 VSS.t75 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1 VDD.t396 VDD.t395 VDD.t396 VDD.t208 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X2 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t122 VDD.t790 VDD.t710 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X3 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t123 VDD.t1385 VDD.t1119 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X4 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t124 VOUT_P.t195 VDD.t1030 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X5 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t2 Folded_Diff_Op_Amp_Layout_0.VCD.t14 VSS.t280 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t37 VSS.t196 VSS.t185 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X7 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t115 VDD.t789 VDD.t729 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X8 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.t28 Folded_Diff_Op_Amp_Layout_0.IB2.t16 VDD.t572 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X9 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t12 VDD.t20 VDD.t9 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X10 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB2.t34 Folded_Diff_Op_Amp_Layout_0.OUT2.t32 VDD.t574 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X11 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2.t35 Folded_Diff_Op_Amp_Layout_0.VPD.t30 VDD.t575 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X12 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t126 VDD.t1388 VDD.t776 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X13 VDD.t394 VDD.t393 VDD.t394 VDD.t162 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X14 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB2.t36 Folded_Diff_Op_Amp_Layout_0.OUT1.t20 VDD.t576 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X15 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t36 VOUT_P.t198 VSS.t72 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X16 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t37 VOUT_P.t199 VSS.t84 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X17 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t127 VOUT_P.t193 VDD.t673 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X18 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t128 VOUT_N.t253 VDD.t907 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X19 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t129 VOUT_N.t254 VDD.t1048 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X20 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t130 VDD.t1395 VDD.t1205 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X21 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t131 VOUT_P.t192 VDD.t835 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X22 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t3 Folded_Diff_Op_Amp_Layout_0.VCD.t13 VSS.t263 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X23 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t113 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t114 VDD.t636 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X24 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t0 Folded_Diff_Op_Amp_Layout_0.VCD.t30 VSS.t260 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X25 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t132 VDD.t1319 VDD.t910 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X26 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS4.t5 Folded_Diff_Op_Amp_Layout_0.IB4.t17 VDD.t519 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X27 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.t4 Folded_Diff_Op_Amp_Layout_0.IB2.t15 VDD.t561 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X28 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t38 VSS.t573 VSS.t87 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X29 a_25284_4817.t1 a_24108_3715.t0 VDD.t48 ppolyf_u r_width=1u r_length=5u
X30 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IVS.t76 VSS.t15 VSS.t14 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X31 Folded_Diff_Op_Amp_Layout_0.IBS Folded_Diff_Op_Amp_Layout_0.IBS.t5 VSS.t36 VSS.t35 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X32 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t133 VDD.t1320 VDD.t910 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X33 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t134 VDD.t1321 VDD.t1053 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X34 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t135 VOUT_P.t189 VDD.t773 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X35 a_24836_4817.t1 a_26012_3715.t1 VDD.t478 ppolyf_u r_width=1u r_length=5u
X36 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IB4.t8 VSS.t528 VSS.t527 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X37 VSS Folded_Diff_Op_Amp_Layout_0.VBIASN.t5 Folded_Diff_Op_Amp_Layout_0.VB2.t32 VSS.t514 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X38 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t136 VDD.t1324 VDD.t806 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X39 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t137 VOUT_P.t188 VDD.t626 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X40 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t138 VDD.t1298 VDD.t914 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X41 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t1 Folded_Diff_Op_Amp_Layout_0.VCD.t31 VSS.t261 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X42 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t39 VOUT_P.t201 VSS.t116 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X43 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t139 VOUT_N.t228 VDD.t1201 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X44 VSS.t488 VSS.t487 VSS.t488 VSS.t299 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X45 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t140 VOUT_P.t186 VDD.t919 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X46 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS1.t2 Folded_Diff_Op_Amp_Layout_0.IBS.t8 VDD.t536 pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
X47 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t38 VSS.t195 VSS.t78 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X48 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t141 VDD.t1303 VDD.t914 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X49 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t13 VDD.t22 VDD.t9 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X50 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t40 VSS.t576 VSS.t78 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X51 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t142 VDD.t1304 VDD.t826 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X52 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t143 VDD.t1305 VDD.t831 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X53 VIN_N1.t0 a_n5986_5540.t1 VDD.t49 ppolyf_u r_width=1u r_length=2.3u
X54 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t111 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t112 VDD.t646 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X55 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t144 VDD.t1306 VDD.t1094 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X56 a_29734_1647.t1 VOUT_N.t1 cap_mim_2f0_m4m5_noshield c_width=21u c_length=21u
X57 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t4 Folded_Diff_Op_Amp_Layout_0.VCD.t12 VSS.t279 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X58 VDD.t392 VDD.t391 VDD.t392 VDD.t327 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X59 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t41 VOUT_P.t203 VSS.t136 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X60 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t145 VOUT_N.t232 VDD.t835 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X61 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t42 VSS.t579 VSS.t113 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X62 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t146 VOUT_N.t261 VDD.t778 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X63 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t147 VDD.t1417 VDD.t838 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X64 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t2 Folded_Diff_Op_Amp_Layout_0.VBM.t27 VSS.t262 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X65 a_n5706_9350.t0 a_n6266_8788.t0 VDD.t44 ppolyf_u r_width=1u r_length=2.3u
X66 VDD.t36 VDD.t37 VDD.t35 ppolyf_u r_width=1u r_length=2.3u
X67 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IVS.t56 VSS.t547 VSS.t545 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X68 VDD.t390 VDD.t389 VDD.t390 VDD.t268 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X69 VSS.t486 VSS.t485 VSS.t486 VSS.t299 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X70 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t14 VDD.t8 VDD.t7 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X71 VDD.t388 VDD.t387 VDD.t388 VDD.t265 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X72 filter_res_magic_0.R7_R8_R10_C a_n6826_5540.t1 VDD.t118 ppolyf_u r_width=1u r_length=2.3u
X73 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t32 VSS.t229 VSS.t56 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X74 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t43 VSS.t580 VSS.t108 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X75 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t44 VSS.t581 VSS.t149 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X76 Folded_Diff_Op_Amp_Layout_0.IBS Folded_Diff_Op_Amp_Layout_0.IBIAS1.t3 VDD.t508 VDD.t507 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X77 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB2.t38 Folded_Diff_Op_Amp_Layout_0.OUT1.t21 VDD.t577 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X78 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t39 VSS.t194 VSS.t156 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X79 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t148 VOUT_P.t183 VDD.t844 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X80 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t149 VDD.t1420 VDD.t1098 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X81 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB2.t39 Folded_Diff_Op_Amp_Layout_0.OUT2.t31 VDD.t578 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X82 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t150 VOUT_N.t263 VDD.t1100 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X83 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t5 Folded_Diff_Op_Amp_Layout_0.VB1.t26 VSS.t281 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X84 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t40 VOUT_N.t36 VSS.t92 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X85 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.VB2.t22 Folded_Diff_Op_Amp_Layout_0.VB2.t23 VDD.t570 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X86 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t109 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t110 VDD.t721 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X87 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t107 VDD.t735 VDD.t657 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X88 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t152 VDD.t1423 VDD.t1035 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X89 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t153 VDD.t1424 VDD.t1098 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X90 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t45 VSS.t582 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X91 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t34 Folded_Diff_Op_Amp_Layout_0.VPD.t15 VDD.t943 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X92 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS1.t4 Folded_Diff_Op_Amp_Layout_0.VBIASN.t0 VDD.t481 pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
X93 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t7 Folded_Diff_Op_Amp_Layout_0.IPD.t23 VDD.t500 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X94 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t154 VOUT_P.t180 VDD.t882 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X95 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t155 VDD.t1204 VDD.t885 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X96 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t15 Folded_Diff_Op_Amp_Layout_0.BD.t28 VDD.t11 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X97 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t46 VOUT_P.t208 VSS.t100 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X98 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t7 Folded_Diff_Op_Amp_Layout_0.BD.t44 VDD.t498 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X99 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.IB5.t6 Folded_Diff_Op_Amp_Layout_0.IB5.t7 VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X100 VSS.t484 VSS.t483 VSS.t484 VSS.t293 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X101 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t41 VOUT_N.t35 VSS.t182 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X102 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t156 VDD.t1206 VDD.t1205 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X103 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t157 VOUT_P.t179 VDD.t828 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X104 Folded_Diff_Op_Amp_Layout_0.OUT1.t4 a_29734_1647.t1 VDD.t411 ppolyf_u r_width=1u r_length=6.2u
X105 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IB4.t19 VSS.t616 VSS.t14 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X106 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1.t35 VDD.t947 VDD.t946 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X107 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t36 Folded_Diff_Op_Amp_Layout_0.VND.t15 VDD.t948 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X108 VDD.t386 VDD.t385 VDD.t386 VDD.t257 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X109 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t3 Folded_Diff_Op_Amp_Layout_0.VCD.t33 VSS.t263 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X110 VSS.t482 VSS.t481 VSS.t482 VSS.t314 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X111 VDD.t384 VDD.t383 VDD.t384 VDD.t314 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X112 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t47 VSS.t585 VSS.t156 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X113 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t158 VOUT_N.t205 VDD.t922 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X114 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t105 VDD.t734 VDD.t719 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X115 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t33 Folded_Diff_Op_Amp_Layout_0.IND.t32 VSS.t0 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X116 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t160 VDD.t1211 VDD.t925 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X117 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t48 VOUT_P.t210 VSS.t140 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X118 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t8 Folded_Diff_Op_Amp_Layout_0.IPD.t22 VDD.t501 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X119 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t42 VOUT_N.t34 VSS.t140 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X120 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t49 VSS.t588 VSS.t80 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X121 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t103 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t104 VDD.t726 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X122 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2.t40 Folded_Diff_Op_Amp_Layout_0.VND.t29 VDD.t575 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X123 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t161 VOUT_P.t178 VDD.t895 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X124 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t101 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t102 VDD.t714 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X125 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB2.t41 Folded_Diff_Op_Amp_Layout_0.OUT2.t30 VDD.t576 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X126 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2.t42 Folded_Diff_Op_Amp_Layout_0.VPD.t27 VDD.t579 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X127 a_29734_3659.t4 VOUT_P.t225 cap_mim_2f0_m4m5_noshield c_width=21u c_length=21u
X128 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t16 Folded_Diff_Op_Amp_Layout_0.BD.t27 VDD.t11 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X129 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t8 Folded_Diff_Op_Amp_Layout_0.IND.t47 VDD.t461 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X130 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t162 VDD.t1214 VDD.t900 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X131 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t9 Folded_Diff_Op_Amp_Layout_0.BD.t40 VDD.t467 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X132 a_n5986_9350.t0 VIN_P1.t0 VDD.t49 ppolyf_u r_width=1u r_length=2.3u
X133 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t17 VDD.t14 VDD.t7 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X134 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t163 VDD.t1215 VDD.t885 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X135 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t164 VDD.t694 VDD.t693 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X136 VSS.t480 VSS.t479 VSS.t480 VSS.t317 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X137 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t165 VOUT_P.t175 VDD.t695 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X138 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t166 VOUT_P.t174 VDD.t698 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X139 a_n7106_6102.t1 a_n5986_5540.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X140 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t167 VDD.t702 VDD.t701 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X141 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1.t37 VDD.t952 VDD.t951 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X142 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t99 VDD.t1312 VDD.t719 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X143 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3.t16 Folded_Diff_Op_Amp_Layout_0.IND.t0 VSS.t27 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X144 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t169 VOUT_P.t173 VDD.t602 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X145 VDD.t502 VDD.t503 VDD.t35 ppolyf_u r_width=1u r_length=2.3u
X146 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t34 Folded_Diff_Op_Amp_Layout_0.IPD.t55 VSS.t0 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X147 VDD.t382 VDD.t381 VDD.t382 VDD.t144 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X148 Folded_Diff_Op_Amp_Layout_0.IB5 Folded_Diff_Op_Amp_Layout_0.IB5.t4 Folded_Diff_Op_Amp_Layout_0.VB4.t1 VSS.t59 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X149 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t170 VDD.t706 VDD.t705 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X150 a_24556_2845.t0 a_24836_1743.t0 VDD.t410 ppolyf_u r_width=1u r_length=5u
X151 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t35 Folded_Diff_Op_Amp_Layout_0.IND.t31 VSS.t8 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X152 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t36 VSS.t214 VSS.t3 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X153 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t171 VOUT_N.t94 VDD.t707 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X154 a_n6826_9350.t0 a_n7106_8433.t2 VDD.t118 ppolyf_u r_width=1u r_length=2.3u
X155 a_n6546_6102.t1 a_n5426_5540.t0 VDD.t89 ppolyf_u r_width=1u r_length=2.3u
X156 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t172 VDD.t711 VDD.t710 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X157 VDD.t380 VDD.t379 VDD.t380 VDD.t226 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X158 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.t2 Folded_Diff_Op_Amp_Layout_0.IB2.t13 VDD.t560 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X159 VSS.t478 VSS.t477 VSS.t478 VSS.t311 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X160 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1.t38 VDD.t953 VDD.t946 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X161 VSS.t476 VSS.t475 VSS.t476 VSS.t302 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X162 VDD.t378 VDD.t377 VDD.t378 VDD.t159 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X163 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3.t17 Folded_Diff_Op_Amp_Layout_0.IND.t1 VSS.t28 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X164 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t173 VDD.t1222 VDD.t1044 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X165 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t174 VDD.t1223 VDD.t1041 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X166 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t30 Folded_Diff_Op_Amp_Layout_0.VB4.t31 VSS.t226 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X167 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t10 Folded_Diff_Op_Amp_Layout_0.BD.t41 VDD.t468 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X168 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t37 VSS.t215 VSS.t204 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X169 VDD Folded_Diff_Op_Amp_Layout_0.VB2.t44 Folded_Diff_Op_Amp_Layout_0.IB2.t0 VDD.t580 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=1u
X170 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IVS.t54 VSS.t546 VSS.t545 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X171 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t97 VDD.t1311 VDD.t712 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X172 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t176 VDD.t1224 VDD.t597 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X173 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t177 VDD.t1225 VDD.t1119 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X174 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t178 VOUT_N.t207 VDD.t1030 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X175 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t95 VDD.t1310 VDD.t729 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X176 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t9 Folded_Diff_Op_Amp_Layout_0.BD.t46 VDD.t462 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X177 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB2.t45 Folded_Diff_Op_Amp_Layout_0.OUT1.t23 VDD.t578 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X178 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t180 VOUT_N.t208 VDD.t623 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X179 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t181 VOUT_P.t167 VDD.t1048 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X180 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t182 VOUT_P.t166 VDD.t907 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X181 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t52 Folded_Diff_Op_Amp_Layout_0.IVS.t53 VSS.t540 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X182 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t183 VDD.t904 VDD.t900 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X183 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t38 VSS.t216 VSS.t3 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X184 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t184 VOUT_P.t164 VDD.t594 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X185 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t185 VOUT_P.t163 VDD.t907 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X186 a_26292_4817.t0 a_26012_3715.t0 VDD.t32 ppolyf_u r_width=1u r_length=5u
X187 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t39 Folded_Diff_Op_Amp_Layout_0.IPD.t53 VSS.t49 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X188 a_26740_4817.t0 a_27020_3715.t1 VDD.t33 ppolyf_u r_width=1u r_length=5u
X189 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t186 VDD.t911 VDD.t910 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X190 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t21 Folded_Diff_Op_Amp_Layout_0.IVS.t66 VDD.t135 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X191 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t11 Folded_Diff_Op_Amp_Layout_0.BD.t42 VDD.t469 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X192 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB2.t46 Folded_Diff_Op_Amp_Layout_0.OUT2.t29 VDD.t574 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X193 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t187 VOUT_N.t131 VDD.t773 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X194 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t188 VDD.t915 VDD.t914 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X195 a_n6266_10267.t1 a_n5706_9705.t1 VDD.t44 ppolyf_u r_width=1u r_length=2.3u
X196 VDD.t376 VDD.t375 VDD.t376 VDD.t162 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X197 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t189 VOUT_N.t133 VDD.t797 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X198 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t190 VDD.t918 VDD.t815 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X199 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t10 Folded_Diff_Op_Amp_Layout_0.IND.t49 VDD.t463 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X200 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t191 VOUT_N.t135 VDD.t919 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X201 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t43 VSS.t187 VSS.t98 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X202 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t192 VDD.t1087 VDD.t898 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X203 VSS.t474 VSS.t472 VSS.t474 VSS.t473 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X204 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t6 Folded_Diff_Op_Amp_Layout_0.VCD.t11 VSS.t263 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X205 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t193 VDD.t1088 VDD.t914 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X206 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t194 VOUT_N.t167 VDD.t866 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X207 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t195 VOUT_N.t168 VDD.t919 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X208 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t196 VDD.t1093 VDD.t664 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X209 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t39 Folded_Diff_Op_Amp_Layout_0.VPD.t12 VDD.t954 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X210 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t197 VDD.t1095 VDD.t1094 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X211 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t40 Folded_Diff_Op_Amp_Layout_0.IPD.t52 VSS.t5 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X212 VDD.t374 VDD.t373 VDD.t374 VDD.t314 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X213 Folded_Diff_Op_Amp_Layout_0.OUT1.t5 a_29734_1647.t1 VDD.t412 ppolyf_u r_width=1u r_length=6.2u
X214 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3.t18 Folded_Diff_Op_Amp_Layout_0.IPD.t63 VSS.t250 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X215 VSS.t471 VSS.t470 VSS.t471 VSS.t419 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X216 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t198 VOUT_P.t160 VDD.t778 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X217 a_n5986_9350.t1 a_n7106_8788.t1 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X218 a_n5146_6102.t1 a_n4866_5185.t1 VDD.t114 ppolyf_u r_width=1u r_length=2.3u
X219 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t44 VSS.t186 VSS.t185 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X220 Folded_Diff_Op_Amp_Layout_0.OUT1.t2 a_29734_1647.t0 VDD.t66 ppolyf_u r_width=1u r_length=6.2u
X221 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t41 Folded_Diff_Op_Amp_Layout_0.IND.t28 VSS.t0 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X222 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t40 Folded_Diff_Op_Amp_Layout_0.VPD.t11 VDD.t954 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X223 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t42 VSS.t491 VSS.t56 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X224 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2.t47 Folded_Diff_Op_Amp_Layout_0.VND.t27 VDD.t579 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X225 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t11 Folded_Diff_Op_Amp_Layout_0.IND.t50 VDD.t499 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X226 a_n5426_9350.t1 a_n6546_8788.t1 VDD.t89 ppolyf_u r_width=1u r_length=2.3u
X227 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t199 VDD.t1099 VDD.t1098 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X228 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB4.t28 VSS.t225 VSS.t224 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X229 VSS.t469 VSS.t468 VSS.t469 VSS.t340 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X230 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t200 VOUT_P.t158 VDD.t1100 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X231 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IB4.t6 VSS.t564 VSS.t545 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X232 a_n6546_6102.t0 filter_res_magic_0.R7_R8_R10_C VDD.t34 ppolyf_u r_width=1u r_length=2.3u
X233 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t201 VDD.t1234 VDD.t597 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X234 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS4.t2 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t3 VDD.t50 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X235 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t93 VDD.t1309 VDD.t657 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X236 VSS Folded_Diff_Op_Amp_Layout_0.VBIASN.t3 Folded_Diff_Op_Amp_Layout_0.VBIASN.t4 VSS.t255 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X237 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t203 VDD.t1235 VDD.t1035 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X238 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t204 VOUT_P.t157 VDD.t599 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X239 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t205 VDD.t1238 VDD.t1098 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X240 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t22 VDD.t541 VDD.t403 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X241 VDD.t372 VDD.t371 VDD.t372 VDD.t162 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X242 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t206 VOUT_N.t212 VDD.t609 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X243 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB4.t26 VSS.t45 VSS.t44 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X244 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t12 Folded_Diff_Op_Amp_Layout_0.IND.t51 VDD.t456 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X245 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB2.t48 Folded_Diff_Op_Amp_Layout_0.OUT1.t25 VDD.t577 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X246 VSS.t467 VSS.t466 VSS.t467 VSS.t305 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X247 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t45 VOUT_N.t33 VSS.t182 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X248 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t207 VDD.t1241 VDD.t607 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X249 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t23 VDD.t542 VDD.t93 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X250 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t79 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t1 VSS.t16 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X251 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3.t19 Folded_Diff_Op_Amp_Layout_0.OUT2.t9 VSS.t248 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X252 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t4 Folded_Diff_Op_Amp_Layout_0.VBM.t25 VSS.t264 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X253 VDD.t370 VDD.t369 VDD.t370 VDD.t202 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.56u
X254 VSS.t465 VSS.t464 VSS.t465 VSS.t302 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X255 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t208 VOUT_P.t156 VDD.t1152 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X256 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t50 VSS.t589 VSS.t87 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X257 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t209 VDD.t1244 VDD.t1205 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X258 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t210 VOUT_N.t214 VDD.t828 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X259 a_24108_2845.t1 VOUT_P.t197 VDD.t491 ppolyf_u r_width=1u r_length=5u
X260 Folded_Diff_Op_Amp_Layout_0.IB3 Folded_Diff_Op_Amp_Layout_0.VB3.t6 Folded_Diff_Op_Amp_Layout_0.VB3.t7 VSS.t23 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X261 VDD.t368 VDD.t367 VDD.t368 VDD.t257 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X262 a_n5426_10267.t1 a_n4866_9705.t1 VDD.t49 ppolyf_u r_width=1u r_length=2.3u
X263 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t211 VOUT_P.t154 VDD.t922 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X264 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t12 Folded_Diff_Op_Amp_Layout_0.IPD.t18 VDD.t470 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X265 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t212 VDD.t926 VDD.t925 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X266 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t7 Folded_Diff_Op_Amp_Layout_0.VB1.t24 VSS.t278 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X267 VSS.t463 VSS.t462 VSS.t463 VSS.t314 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X268 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t91 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t92 VDD.t661 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X269 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t213 VDD.t927 VDD.t671 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X270 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3.t20 Folded_Diff_Op_Amp_Layout_0.IPD.t65 VSS.t27 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X271 VDD.t64 VDD.t65 VDD.t35 ppolyf_u r_width=1u r_length=2.3u
X272 VDD.t366 VDD.t365 VDD.t366 VDD.t218 pfet_03v3 ad=0.814p pd=3.65u as=0 ps=0 w=3.13u l=0.56u
X273 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3.t21 Folded_Diff_Op_Amp_Layout_0.OUT1.t12 VSS.t251 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X274 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t89 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t90 VDD.t726 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X275 a_n7106_9350.t1 a_n6826_9705.t1 VDD.t118 ppolyf_u r_width=1u r_length=2.3u
X276 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t13 Folded_Diff_Op_Amp_Layout_0.BD.t36 VDD.t460 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X277 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t214 VDD.t928 VDD.t847 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X278 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t50 Folded_Diff_Op_Amp_Layout_0.IVS.t51 VSS.t540 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X279 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2.t49 Folded_Diff_Op_Amp_Layout_0.VND.t25 VDD.t583 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X280 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t215 VOUT_P.t150 VDD.t929 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X281 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t24 Folded_Diff_Op_Amp_Layout_0.IVS.t69 VDD.t135 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X282 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t216 VDD.t932 VDD.t680 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X283 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3.t22 Folded_Diff_Op_Amp_Layout_0.IPD.t66 VSS.t28 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X284 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t87 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t88 VDD.t721 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X285 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t217 VOUT_N.t137 VDD.t695 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X286 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t25 Folded_Diff_Op_Amp_Layout_0.IVS.t70 VDD.t135 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X287 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t218 VOUT_N.t138 VDD.t698 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X288 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t45 VSS.t492 VSS.t204 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X289 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t219 VDD.t937 VDD.t701 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X290 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t85 VDD.t1396 VDD.t650 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X291 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t24 Folded_Diff_Op_Amp_Layout_0.VB4.t25 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X292 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t13 Folded_Diff_Op_Amp_Layout_0.BD.t50 VDD.t458 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X293 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t14 Folded_Diff_Op_Amp_Layout_0.BD.t51 VDD.t457 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X294 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t221 VOUT_N.t170 VDD.t762 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X295 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t83 VDD.t1221 VDD.t719 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X296 VDD.t364 VDD.t363 VDD.t364 VDD.t231 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X297 a_n4866_9705.t0 a_n5146_8788.t1 VDD.t114 ppolyf_u r_width=1u r_length=2.3u
X298 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t46 VSS.t493 VSS.t56 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X299 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2.t50 Folded_Diff_Op_Amp_Layout_0.VND.t24 VDD.t575 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X300 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t223 VOUT_N.t171 VDD.t602 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X301 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t26 Folded_Diff_Op_Amp_Layout_0.IVS.t71 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X302 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.t26 Folded_Diff_Op_Amp_Layout_0.IB2.t12 VDD.t171 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X303 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB2.t52 Folded_Diff_Op_Amp_Layout_0.OUT2.t28 VDD.t576 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X304 VSS.t461 VSS.t460 VSS.t461 VSS.t320 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X305 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t224 VDD.t1107 VDD.t705 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X306 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t225 VOUT_N.t172 VDD.t599 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X307 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t47 Folded_Diff_Op_Amp_Layout_0.IPD.t49 VSS.t8 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X308 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t226 VOUT_P.t147 VDD.t707 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X309 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VB3.t0 Folded_Diff_Op_Amp_Layout_0.IB3.t5 VSS.t284 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X310 VSS.t459 VSS.t458 VSS.t459 VSS.t320 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X311 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t227 VDD.t1112 VDD.t710 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X312 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t228 VDD.t1113 VDD.t1094 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X313 VDD.t362 VDD.t361 VDD.t362 VDD.t226 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X314 VDD.t360 VDD.t359 VDD.t360 VDD.t218 pfet_03v3 ad=0.814p pd=3.65u as=0 ps=0 w=3.13u l=0.56u
X315 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t27 Folded_Diff_Op_Amp_Layout_0.IVS.t72 VDD.t67 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X316 a_24556_2845.t1 VOUT_N.t75 VDD.t488 ppolyf_u r_width=1u r_length=5u
X317 VDD.t358 VDD.t357 VDD.t358 VDD.t202 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.56u
X318 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t48 VSS.t496 VSS.t206 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X319 VDD.t356 VDD.t355 VDD.t356 VDD.t159 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X320 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t229 VDD.t1114 VDD.t1041 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X321 Folded_Diff_Op_Amp_Layout_0.VBIASN Folded_Diff_Op_Amp_Layout_0.VBIASN.t1 VSS.t254 VSS.t253 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X322 a_n7106_8433.t0 a_n6546_8788.t0 VDD.t34 ppolyf_u r_width=1u r_length=2.3u
X323 a_n5146_6102.t0 a_n5706_5540.t1 VDD.t55 ppolyf_u r_width=1u r_length=2.3u
X324 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t230 VDD.t1403 VDD.t838 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X325 VDD.t354 VDD.t353 VDD.t354 VDD.t254 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X326 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t231 VOUT_N.t256 VDD.t1152 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X327 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t232 VDD.t1406 VDD.t597 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X328 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS4.t6 Folded_Diff_Op_Amp_Layout_0.IB4.t16 VDD.t519 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X329 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t81 VDD.t1220 VDD.t712 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X330 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t15 Folded_Diff_Op_Amp_Layout_0.IND.t54 VDD.t459 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X331 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t46 VOUT_N.t32 VSS.t175 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X332 Folded_Diff_Op_Amp_Layout_0.IB5 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t5 VDD.t472 VDD.t471 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X333 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t41 Folded_Diff_Op_Amp_Layout_0.VND.t13 VDD.t954 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X334 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t28 VDD.t551 VDD.t403 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X335 a_n7106_6102.t0 filter_res_magic_0.R3_R7.t1 VDD.t90 ppolyf_u r_width=1u r_length=2.3u
X336 VSS.t457 VSS.t456 VSS.t457 VSS.t302 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X337 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t234 VOUT_P.t144 VDD.t623 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X338 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t51 VOUT_P.t213 VSS.t67 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X339 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t52 VSS.t592 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X340 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t8 Folded_Diff_Op_Amp_Layout_0.VCD.t10 VSS.t280 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X341 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t235 VDD.t1409 VDD.t1051 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X342 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t236 VOUT_N.t258 VDD.t594 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X343 VDD.t352 VDD.t351 VDD.t352 VDD.t271 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X344 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t29 VDD.t552 VDD.t93 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X345 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t30 VDD.t553 VDD.t403 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X346 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t237 VDD.t1412 VDD.t900 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X347 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t238 VOUT_N.t260 VDD.t907 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X348 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t239 VDD.t1427 VDD.t676 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X349 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3.t24 Folded_Diff_Op_Amp_Layout_0.IND.t41 VSS.t250 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X350 VSS.t455 VSS.t453 VSS.t455 VSS.t454 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X351 a_n6546_10267.t0 a_n5986_9705.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X352 VDD.t350 VDD.t349 VDD.t350 VDD.t208 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X353 VSS.t452 VSS.t451 VSS.t452 VSS.t419 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X354 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t47 VOUT_N.t31 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X355 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t31 VDD.t94 VDD.t93 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X356 VSS Folded_Diff_Op_Amp_Layout_0.IB4.t4 Folded_Diff_Op_Amp_Layout_0.IB4.t5 VSS.t540 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X357 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t80 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t117 VSS.t16 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X358 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t240 VOUT_N.t265 VDD.t685 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X359 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t241 VDD.t1430 VDD.t813 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X360 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB2.t53 Folded_Diff_Op_Amp_Layout_0.OUT1.t28 VDD.t574 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X361 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t53 VSS.t593 VSS.t87 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X362 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t5 Folded_Diff_Op_Amp_Layout_0.VCD.t35 VSS.t260 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X363 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t18 Folded_Diff_Op_Amp_Layout_0.BD.t25 VDD.t4 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X364 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t49 VSS.t46 VSS.t3 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X365 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB2.t54 Folded_Diff_Op_Amp_Layout_0.OUT1.t29 VDD.t578 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X366 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t242 VDD.t1431 VDD.t815 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X367 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t243 VOUT_P.t141 VDD.t797 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X368 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t244 VDD.t1434 VDD.t815 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X369 a_n5426_10267.t0 a_n5986_9705.t1 VDD.t89 ppolyf_u r_width=1u r_length=2.3u
X370 VDD.t348 VDD.t347 VDD.t348 VDD.t168 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X371 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t245 VDD.t1435 VDD.t898 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X372 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t32 VDD.t95 VDD.t78 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X373 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t54 VOUT_P.t216 VSS.t72 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X374 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t246 VDD.t1436 VDD.t664 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X375 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t247 VOUT_P.t137 VDD.t866 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X376 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t248 VOUT_P.t136 VDD.t919 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X377 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB4.t22 VSS.t40 VSS.t39 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X378 VDD Folded_Diff_Op_Amp_Layout_0.VBM.t32 Folded_Diff_Op_Amp_Layout_0.VBM.t33 VDD.t56 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X379 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t48 VOUT_N.t30 VSS.t175 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X380 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t249 VOUT_N.t215 VDD.t629 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X381 VDD.t494 VDD.t495 VDD.t473 ppolyf_u r_width=1u r_length=6.2u
X382 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t33 VDD.t96 VDD.t80 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X383 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB2.t55 Folded_Diff_Op_Amp_Layout_0.OUT2.t27 VDD.t577 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X384 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t55 VSS.t596 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X385 VSS.t450 VSS.t449 VSS.t450 VSS.t293 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X386 VSS.t448 VSS.t447 VSS.t448 VSS.t290 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X387 Folded_Diff_Op_Amp_Layout_0.OUT1.t3 a_29734_1647.t1 VDD.t139 ppolyf_u r_width=1u r_length=6.2u
X388 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t250 VOUT_P.t135 VDD.t682 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X389 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t251 VDD.t1264 VDD.t1005 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X390 VDD.t431 VDD.t432 VDD.t430 ppolyf_u r_width=1u r_length=6.2u
X391 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB4.t20 VSS.t38 VSS.t37 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X392 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t48 Folded_Diff_Op_Amp_Layout_0.IVS.t49 VSS.t535 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X393 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t252 VOUT_P.t133 VDD.t746 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X394 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t79 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t80 VDD.t726 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X395 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.VB2.t20 Folded_Diff_Op_Amp_Layout_0.VB2.t21 VDD.t569 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X396 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2.t56 Folded_Diff_Op_Amp_Layout_0.VPD.t23 VDD.t583 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X397 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t49 VOUT_N.t29 VSS.t84 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X398 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t6 Folded_Diff_Op_Amp_Layout_0.VBM.t23 VSS.t262 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X399 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t19 Folded_Diff_Op_Amp_Layout_0.BD.t24 VDD.t4 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X400 VDD.t346 VDD.t345 VDD.t346 VDD.t314 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X401 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t34 Folded_Diff_Op_Amp_Layout_0.IVS.t12 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X402 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t253 VDD.t1267 VDD.t822 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X403 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t254 VDD.t1268 VDD.t791 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X404 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t255 VDD.t593 VDD.t592 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X405 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t8 Folded_Diff_Op_Amp_Layout_0.IBIAS.t9 VDD.t1 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X406 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t256 VOUT_N.t77 VDD.t594 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X407 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t257 VDD.t598 VDD.t597 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X408 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t9 Folded_Diff_Op_Amp_Layout_0.VB1.t22 VSS.t277 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X409 a_n5706_9350.t1 a_n5146_8788.t0 VDD.t55 ppolyf_u r_width=1u r_length=2.3u
X410 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t50 VSS.t172 VSS.t113 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X411 VSS.t446 VSS.t445 VSS.t446 VSS.t320 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X412 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t7 VDD.t525 VDD.t524 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X413 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t35 Folded_Diff_Op_Amp_Layout_0.IVS.t13 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X414 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t258 VOUT_N.t78 VDD.t599 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X415 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t10 Folded_Diff_Op_Amp_Layout_0.VB1.t21 VSS.t281 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X416 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t259 VOUT_N.t79 VDD.t602 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X417 VDD.t344 VDD.t343 VDD.t344 VDD.t268 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X418 a_n6266_6102.t1 a_n6826_5540.t0 VDD.t43 ppolyf_u r_width=1u r_length=2.3u
X419 VDD.t342 VDD.t341 VDD.t342 VDD.t240 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X420 VDD.t340 VDD.t339 VDD.t340 VDD.t265 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X421 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2.t57 Folded_Diff_Op_Amp_Layout_0.VND.t21 VDD.t579 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X422 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t260 VDD.t606 VDD.t605 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X423 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t261 VDD.t608 VDD.t607 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X424 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t262 VOUT_P.t129 VDD.t609 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X425 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t11 Folded_Diff_Op_Amp_Layout_0.VB1.t20 VSS.t264 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X426 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS1.t6 Folded_Diff_Op_Amp_Layout_0.IB5.t10 VDD.t436 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X427 VOUT_N.t272 VOUT_OPAMP_P.t1 cap_mim_2f0_m4m5_noshield c_width=15.2u c_length=16u
X428 VDD.t338 VDD.t337 VDD.t338 VDD.t223 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X429 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1.t42 VDD.t962 VDD.t961 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X430 VDD.t336 VDD.t335 VDD.t336 VDD.t289 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X431 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t263 VOUT_N.t235 VDD.t1152 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X432 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t56 VSS.t597 VSS.t185 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X433 a_n7106_9350.t0 a_n7106_8788.t0 VDD.t90 ppolyf_u r_width=1u r_length=2.3u
X434 filter_res_magic_0.R7_R8_R10_C.t0 a_n7106_8433.t4 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X435 Folded_Diff_Op_Amp_Layout_0.VBM Folded_Diff_Op_Amp_Layout_0.VBM.t30 VDD.t92 VDD.t91 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X436 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t52 Folded_Diff_Op_Amp_Layout_0.IND.t25 VSS.t5 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X437 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t53 Folded_Diff_Op_Amp_Layout_0.IPD.t47 VSS.t49 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X438 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t51 VSS.t171 VSS.t80 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X439 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t52 VOUT_N.t28 VSS.t84 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X440 VDD.t484 VDD.t485 VDD.t86 ppolyf_u r_width=1u r_length=5u
X441 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS4.t8 Folded_Diff_Op_Amp_Layout_0.IB4.t14 VDD.t519 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X442 VSS Folded_Diff_Op_Amp_Layout_0.IB4.t21 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t19 VSS.t16 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X443 a_n5986_7019.t1 a_n5706_6457.t0 VDD.t44 ppolyf_u r_width=1u r_length=2.3u
X444 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2.t58 Folded_Diff_Op_Amp_Layout_0.VPD.t22 VDD.t579 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X445 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t7 Folded_Diff_Op_Amp_Layout_0.VBM.t22 VSS.t278 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X446 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t77 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t78 VDD.t661 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X447 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS4.t9 Folded_Diff_Op_Amp_Layout_0.IB4.t13 VDD.t519 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X448 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t8 Folded_Diff_Op_Amp_Layout_0.VCD.t49 VSS.t261 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X449 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t264 VDD.t1329 VDD.t671 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X450 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t265 VDD.t1330 VDD.t765 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X451 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t266 VOUT_P.t127 VDD.t612 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X452 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t16 Folded_Diff_Op_Amp_Layout_0.IND.t55 VDD.t500 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X453 a_n5146_10267.t1 a_n5426_9350.t0 VDD.t114 ppolyf_u r_width=1u r_length=2.3u
X454 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t9 Folded_Diff_Op_Amp_Layout_0.VCD.t50 VSS.t263 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X455 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.t30 Folded_Diff_Op_Amp_Layout_0.IB2.t10 VDD.t573 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X456 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t54 Folded_Diff_Op_Amp_Layout_0.IPD.t46 VSS.t8 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X457 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t53 VOUT_N.t27 VSS.t75 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X458 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t267 VOUT_P.t126 VDD.t623 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X459 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t268 VDD.t1335 VDD.t847 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X460 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t269 VOUT_N.t238 VDD.t929 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X461 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t270 VOUT_P.t125 VDD.t626 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X462 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t12 Folded_Diff_Op_Amp_Layout_0.VCD.t9 VSS.t279 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X463 a_n5706_5185.t1 a_n6266_4623.t0 VDD.t44 ppolyf_u r_width=1u r_length=2.3u
X464 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t271 VDD.t1161 VDD.t680 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X465 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t75 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t76 VDD.t721 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X466 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t272 VDD.t1162 VDD.t632 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X467 a_n6546_10267.t1 a_n7106_9705.t0 VDD.t34 ppolyf_u r_width=1u r_length=2.3u
X468 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t54 VSS.t166 VSS.t78 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X469 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t14 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t15 VDD.t446 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X470 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t55 Folded_Diff_Op_Amp_Layout_0.IND.t24 VSS.t49 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X471 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t73 VDD.t731 VDD.t650 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X472 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t17 Folded_Diff_Op_Amp_Layout_0.IND.t56 VDD.t501 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X473 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t57 VSS.t598 VSS.t98 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X474 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t274 VOUT_P.t123 VDD.t762 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X475 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t275 VDD.t1165 VDD.t634 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X476 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t276 VDD.t1166 VDD.t791 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X477 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t55 VOUT_N.t26 VSS.t136 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X478 VDD.t334 VDD.t333 VDD.t334 VDD.t231 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X479 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t56 VSS.t57 VSS.t56 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X480 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t56 VSS.t163 VSS.t113 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X481 VSS.t444 VSS.t443 VSS.t444 VSS.t308 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X482 VSS.t442 VSS.t441 VSS.t442 VSS.t317 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X483 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t277 VOUT_P.t121 VDD.t794 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X484 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t278 VOUT_P.t120 VDD.t599 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X485 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t81 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t4 VSS.t30 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X486 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS1.t7 Folded_Diff_Op_Amp_Layout_0.IBS.t0 VDD.t433 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X487 VSS.t440 VSS.t439 VSS.t440 VSS.t340 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X488 VDD.t116 VDD.t117 VDD.t115 ppolyf_u r_width=1u r_length=5u
X489 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t58 VOUT_P.t220 VSS.t116 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X490 VSS.t438 VSS.t437 VSS.t438 VSS.t365 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X491 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t14 Folded_Diff_Op_Amp_Layout_0.IPD.t16 VDD.t461 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X492 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t57 VSS.t162 VSS.t149 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X493 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t279 VDD.t1171 VDD.t1094 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X494 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t280 VDD.t1148 VDD.t1044 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X495 a_25564_2845.t1 a_25284_1743.t1 VDD.t53 ppolyf_u r_width=1u r_length=5u
X496 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t18 Folded_Diff_Op_Amp_Layout_0.BD.t55 VDD.t467 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X497 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t59 VSS.t601 VSS.t156 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X498 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t58 VSS.t161 VSS.t70 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X499 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t10 Folded_Diff_Op_Amp_Layout_0.VBM.t19 VSS.t277 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X500 VSS.t436 VSS.t435 VSS.t436 VSS.t340 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X501 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1.t43 VDD.t964 VDD.t963 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X502 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t59 VOUT_N.t25 VSS.t67 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X503 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t281 VDD.t1149 VDD.t838 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X504 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t20 Folded_Diff_Op_Amp_Layout_0.BD.t23 VDD.t17 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X505 VSS.t434 VSS.t433 VSS.t434 VSS.t293 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X506 VDD.t332 VDD.t331 VDD.t332 VDD.t254 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X507 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t282 VOUT_P.t118 VDD.t1012 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X508 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t283 VOUT_P.t117 VDD.t1152 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X509 VSS.t432 VSS.t431 VSS.t432 VSS.t311 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X510 VDD.t330 VDD.t329 VDD.t330 VDD.t165 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X511 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t46 Folded_Diff_Op_Amp_Layout_0.IVS.t47 VSS.t535 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X512 VDD.t328 VDD.t326 VDD.t328 VDD.t327 pfet_03v3 ad=0.13p pd=1.02u as=0 ps=0 w=0.5u l=0.28u
X513 a_n6826_9350.t1 a_n6266_8788.t1 VDD.t43 ppolyf_u r_width=1u r_length=2.3u
X514 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t60 VSS.t158 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X515 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t284 VOUT_P.t116 VDD.t1048 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X516 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.IBS.t10 VSS.t286 VSS.t285 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=1u
X517 VOUT_OPAMP_N.t3 VOUT_OPAMP_N.t4 VDD.t49 ppolyf_u r_width=1u r_length=2.3u
X518 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t57 VSS.t200 VSS.t3 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X519 VDD.t489 VDD.t490 VDD.t40 ppolyf_u r_width=1u r_length=2.3u
X520 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t58 VSS.t201 VSS.t56 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X521 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t285 VDD.t1157 VDD.t765 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X522 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t286 VOUT_N.t188 VDD.t770 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X523 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t11 Folded_Diff_Op_Amp_Layout_0.VCD.t52 VSS.t280 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X524 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t59 Folded_Diff_Op_Amp_Layout_0.IND.t22 VSS.t8 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X525 VSS.t430 VSS.t429 VSS.t430 VSS.t314 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X526 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t60 VOUT_P.t222 VSS.t182 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X527 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t287 VDD.t1160 VDD.t1051 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X528 VDD.t325 VDD.t324 VDD.t325 VDD.t245 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X529 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t71 VDD.t730 VDD.t729 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X530 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t19 Folded_Diff_Op_Amp_Layout_0.BD.t56 VDD.t468 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X531 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3.t25 Folded_Diff_Op_Amp_Layout_0.IND.t42 VSS.t27 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X532 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t21 VDD.t27 VDD.t26 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X533 VDD.t442 VDD.t443 VDD.t35 ppolyf_u r_width=1u r_length=2.3u
X534 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t289 VDD.t809 VDD.t783 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X535 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t290 VDD.t810 VDD.t676 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X536 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2.t60 Folded_Diff_Op_Amp_Layout_0.VND.t20 VDD.t584 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X537 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t61 VSS.t157 VSS.t156 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X538 a_n7106_7019.t0 a_n6826_6457.t0 VDD.t118 ppolyf_u r_width=1u r_length=2.3u
X539 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t44 Folded_Diff_Op_Amp_Layout_0.VND.t11 VDD.t954 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X540 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t13 Folded_Diff_Op_Amp_Layout_0.VCD.t8 VSS.t261 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X541 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t14 Folded_Diff_Op_Amp_Layout_0.VCD.t7 VSS.t260 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X542 a_n4866_5185.t0 a_n5426_4623.t0 VDD.t49 ppolyf_u r_width=1u r_length=2.3u
X543 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3.t26 Folded_Diff_Op_Amp_Layout_0.OUT1.t15 VSS.t248 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X544 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t62 VOUT_N.t24 VSS.t140 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X545 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t61 VSS.t604 VSS.t87 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X546 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t291 VOUT_P.t113 VDD.t685 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X547 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t292 VDD.t814 VDD.t813 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X548 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.IB5.t2 Folded_Diff_Op_Amp_Layout_0.IB5.t3 VSS.t58 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X549 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t15 Folded_Diff_Op_Amp_Layout_0.BD.t38 VDD.t462 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X550 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t45 Folded_Diff_Op_Amp_Layout_0.VND.t10 VDD.t943 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X551 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t293 VDD.t816 VDD.t815 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X552 a_27020_3715.t0 a_26292_1743.t1 VDD.t413 ppolyf_u r_width=1u r_length=5u
X553 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3.t27 Folded_Diff_Op_Amp_Layout_0.IND.t44 VSS.t28 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X554 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t63 VSS.t153 VSS.t80 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X555 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t64 VOUT_N.t23 VSS.t84 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X556 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t65 VSS.t150 VSS.t149 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X557 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t294 VOUT_N.t109 VDD.t817 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X558 VDD.t323 VDD.t322 VDD.t323 VDD.t168 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X559 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.VB2.t18 Folded_Diff_Op_Amp_Layout_0.VB2.t19 VDD.t568 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X560 VDD.t321 VDD.t320 VDD.t321 VDD.t289 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X561 a_n5706_8433.t0 a_n5986_7871.t1 VDD.t44 ppolyf_u r_width=1u r_length=2.3u
X562 VDD.t496 VDD.t497 VDD.t35 ppolyf_u r_width=1u r_length=2.3u
X563 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t60 VSS.t205 VSS.t204 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X564 VSS.t428 VSS.t427 VSS.t428 VSS.t299 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X565 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t12 Folded_Diff_Op_Amp_Layout_0.VCD.t53 VSS.t279 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X566 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t295 VOUT_P.t111 VDD.t629 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X567 a_25564_2845.t0 a_26740_1743.t1 VDD.t54 ppolyf_u r_width=1u r_length=5u
X568 a_n5146_10267.t0 a_n5706_9705.t0 VDD.t55 ppolyf_u r_width=1u r_length=2.3u
X569 a_n6826_5185.t0 filter_res_magic_0.R3_R7.t0 VDD.t118 ppolyf_u r_width=1u r_length=2.3u
X570 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3.t28 Folded_Diff_Op_Amp_Layout_0.OUT1.t17 VSS.t249 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X571 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t296 VDD.t823 VDD.t822 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X572 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t22 Folded_Diff_Op_Amp_Layout_0.BD.t21 VDD.t23 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X573 VSS.t426 VSS.t425 VSS.t426 VSS.t314 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X574 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t62 VSS.t605 VSS.t70 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X575 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS4.t0 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t1 VDD.t50 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X576 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.VB2.t16 Folded_Diff_Op_Amp_Layout_0.VB2.t17 VDD.t567 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X577 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t23 VDD.t526 VDD.t26 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X578 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t24 Folded_Diff_Op_Amp_Layout_0.BD.t19 VDD.t17 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X579 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t297 VOUT_N.t110 VDD.t682 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X580 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t298 VDD.t1190 VDD.t1005 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X581 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t299 VOUT_P.t109 VDD.t1100 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X582 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t16 Folded_Diff_Op_Amp_Layout_0.IPD.t14 VDD.t463 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X583 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t300 VOUT_N.t200 VDD.t746 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X584 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t15 Folded_Diff_Op_Amp_Layout_0.VB1.t16 VSS.t262 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X585 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t61 VSS.t207 VSS.t206 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X586 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t69 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t70 VDD.t726 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X587 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t63 VSS.t629 VSS.t108 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X588 VOUT_N.t74 a_n7106_9705.t1 VDD.t90 ppolyf_u r_width=1u r_length=2.3u
X589 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t301 VDD.t1195 VDD.t822 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X590 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t302 VDD.t1196 VDD.t592 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X591 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t303 VOUT_N.t201 VDD.t698 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X592 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t304 VOUT_P.t106 VDD.t594 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X593 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t305 VOUT_N.t202 VDD.t1201 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X594 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t306 VDD.t792 VDD.t791 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X595 VSS Folded_Diff_Op_Amp_Layout_0.IB4.t2 Folded_Diff_Op_Amp_Layout_0.IB4.t3 VSS.t535 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X596 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t307 VDD.t793 VDD.t781 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X597 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t308 VOUT_N.t104 VDD.t794 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X598 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t25 VDD.t852 VDD.t15 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X599 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t62 VSS.t208 VSS.t204 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X600 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t309 VOUT_P.t103 VDD.t797 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X601 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t67 VDD.t725 VDD.t650 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X602 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t13 Folded_Diff_Op_Amp_Layout_0.VBM.t16 VSS.t281 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X603 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t66 VSS.t148 VSS.t113 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X604 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t64 VOUT_P.t228 VSS.t92 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X605 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t67 VOUT_N.t22 VSS.t92 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X606 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t311 VOUT_P.t102 VDD.t800 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X607 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t82 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t3 VSS.t30 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X608 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t312 VOUT_P.t101 VDD.t602 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X609 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2.t61 Folded_Diff_Op_Amp_Layout_0.VPD.t21 VDD.t583 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X610 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t313 VDD.t805 VDD.t605 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X611 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t314 VDD.t807 VDD.t806 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X612 VDD.t319 VDD.t318 VDD.t319 VDD.t240 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X613 Folded_Diff_Op_Amp_Layout_0.IB5 Folded_Diff_Op_Amp_Layout_0.IB5.t0 Folded_Diff_Op_Amp_Layout_0.VB4.t3 VSS.t199 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X614 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3.t29 Folded_Diff_Op_Amp_Layout_0.OUT2.t12 VSS.t251 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X615 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t65 VSS.t632 VSS.t156 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X616 VDD.t317 VDD.t316 VDD.t317 VDD.t289 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X617 VDD.t585 VDD.t586 VDD.t40 ppolyf_u r_width=1u r_length=2.3u
X618 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t66 VOUT_P.t230 VSS.t100 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X619 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t16 Folded_Diff_Op_Amp_Layout_0.VB1.t15 VSS.t277 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X620 a_n5986_7019.t0 a_n6266_6457.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X621 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3.t30 Folded_Diff_Op_Amp_Layout_0.IPD.t68 VSS.t250 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X622 VSS.t424 VSS.t423 VSS.t424 VSS.t419 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X623 VSS.t422 VSS.t421 VSS.t422 VSS.t293 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X624 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t63 Folded_Diff_Op_Amp_Layout_0.IPD.t41 VSS.t0 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X625 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3.t31 Folded_Diff_Op_Amp_Layout_0.OUT2.t1 VSS.t247 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X626 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t315 VDD.t808 VDD.t765 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X627 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t17 Folded_Diff_Op_Amp_Layout_0.IPD.t13 VDD.t456 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X628 a_n5426_7019.t1 a_n5706_6457.t1 VDD.t89 ppolyf_u r_width=1u r_length=2.3u
X629 VSS.t420 VSS.t418 VSS.t420 VSS.t419 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X630 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t316 VOUT_N.t80 VDD.t612 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X631 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t317 VDD.t616 VDD.t615 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X632 VOUT_OPAMP_P.t2 VOUT_OPAMP_P.t3 VDD.t49 ppolyf_u r_width=1u r_length=2.3u
X633 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t26 Folded_Diff_Op_Amp_Layout_0.BD.t17 VDD.t23 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X634 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t318 VOUT_N.t82 VDD.t617 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X635 a_n5986_5185.t0 a_n6546_4623.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X636 VDD.t315 VDD.t313 VDD.t315 VDD.t314 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X637 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1.t46 VDD.t969 VDD.t963 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X638 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t68 VOUT_N.t21 VSS.t140 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X639 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t69 VSS.t143 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X640 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t65 VDD.t724 VDD.t639 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X641 VDD.t312 VDD.t311 VDD.t312 VDD.t257 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X642 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t320 VOUT_N.t83 VDD.t620 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X643 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t321 VOUT_N.t84 VDD.t623 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X644 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t322 VOUT_N.t85 VDD.t626 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X645 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t18 Folded_Diff_Op_Amp_Layout_0.VB4.t19 VSS.t502 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X646 VDD.t45 VDD.t46 VDD.t35 ppolyf_u r_width=1u r_length=2.3u
X647 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t67 VSS.t635 VSS.t98 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X648 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t323 VOUT_P.t100 VDD.t629 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X649 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t324 VDD.t633 VDD.t632 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X650 VDD.t310 VDD.t309 VDD.t310 VDD.t254 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X651 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t20 Folded_Diff_Op_Amp_Layout_0.IND.t59 VDD.t470 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X652 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t70 VOUT_N.t20 VSS.t140 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X653 VSS.t417 VSS.t416 VSS.t417 VSS.t340 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X654 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t14 Folded_Diff_Op_Amp_Layout_0.VCD.t36 VSS.t261 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X655 a_n6826_8433.t0 a_n7106_7871.t1 VDD.t118 ppolyf_u r_width=1u r_length=2.3u
X656 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t27 VDD.t10 VDD.t9 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X657 a_n5986_5185.t1 a_n5426_4623.t1 VDD.t89 ppolyf_u r_width=1u r_length=2.3u
X658 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2.t62 Folded_Diff_Op_Amp_Layout_0.VPD.t20 VDD.t584 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X659 VDD.t308 VDD.t307 VDD.t308 VDD.t223 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X660 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t325 VDD.t635 VDD.t634 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X661 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t36 Folded_Diff_Op_Amp_Layout_0.IVS.t14 VDD.t67 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X662 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VB3.t12 Folded_Diff_Op_Amp_Layout_0.IB3.t4 VSS.t26 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X663 VSS.t415 VSS.t414 VSS.t415 VSS.t317 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X664 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t326 VDD.t1038 VDD.t791 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X665 a_n6266_10267.t0 a_n6826_9705.t0 VDD.t43 ppolyf_u r_width=1u r_length=2.3u
X666 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t21 Folded_Diff_Op_Amp_Layout_0.BD.t58 VDD.t460 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X667 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t28 VDD.t16 VDD.t15 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X668 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t71 VSS.t139 VSS.t80 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X669 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t327 VOUT_N.t151 VDD.t794 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X670 VDD.t306 VDD.t305 VDD.t306 VDD.t147 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X671 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t328 VDD.t1042 VDD.t1041 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X672 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t64 VSS.t4 VSS.t3 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X673 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2.t63 Folded_Diff_Op_Amp_Layout_0.VND.t19 VDD.t583 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X674 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t68 VSS.t636 VSS.t185 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X675 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t17 Folded_Diff_Op_Amp_Layout_0.VCD.t6 VSS.t279 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X676 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t329 VDD.t1043 VDD.t615 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X677 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t330 VDD.t1045 VDD.t1044 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X678 VDD.t304 VDD.t303 VDD.t304 VDD.t50 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X679 VSS Folded_Diff_Op_Amp_Layout_0.IB4.t22 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t18 VSS.t30 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X680 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t18 Folded_Diff_Op_Amp_Layout_0.BD.t33 VDD.t457 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X681 a_24108_2845.t0 a_25284_1743.t0 VDD.t48 ppolyf_u r_width=1u r_length=5u
X682 VDD.t302 VDD.t301 VDD.t302 VDD.t50 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X683 VSS.t413 VSS.t412 VSS.t413 VSS.t311 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X684 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t19 Folded_Diff_Op_Amp_Layout_0.BD.t34 VDD.t458 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X685 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t69 VOUT_P.t233 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X686 VSS.t411 VSS.t410 VSS.t411 VSS.t290 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X687 VDD.t300 VDD.t299 VDD.t300 VDD.t245 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X688 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t331 VOUT_N.t154 VDD.t1012 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X689 a_26012_2845.t1 a_24836_1743.t1 VDD.t478 ppolyf_u r_width=1u r_length=5u
X690 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t63 VDD.t1297 VDD.t644 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X691 VDD.t298 VDD.t297 VDD.t298 VDD.t271 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X692 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t61 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t62 VDD.t646 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X693 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3.t33 Folded_Diff_Op_Amp_Layout_0.OUT2.t2 VSS.t248 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X694 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t333 VOUT_N.t155 VDD.t1048 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X695 VDD.t296 VDD.t295 VDD.t296 VDD.t141 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X696 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t47 Folded_Diff_Op_Amp_Layout_0.VND.t9 VDD.t970 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X697 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t334 VDD.t1052 VDD.t1051 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X698 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t65 Folded_Diff_Op_Amp_Layout_0.IPD.t39 VSS.t5 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X699 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t72 VOUT_N.t19 VSS.t136 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X700 VSS.t409 VSS.t408 VSS.t409 VSS.t305 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X701 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t70 VOUT_P.t234 VSS.t182 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X702 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t335 VDD.t766 VDD.t765 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X703 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t336 VOUT_N.t100 VDD.t767 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X704 VDD.t294 VDD.t293 VDD.t294 VDD.t240 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X705 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t337 VOUT_P.t95 VDD.t770 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X706 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t338 VOUT_N.t101 VDD.t773 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X707 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB4.t16 VSS.t501 VSS.t500 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X708 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t339 VDD.t777 VDD.t776 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X709 VOUT_OPAMP_N.t1 VOUT_OPAMP_N.t2 VDD.t114 ppolyf_u r_width=1u r_length=2.3u
X710 VDD.t292 VDD.t291 VDD.t292 VDD.t245 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X711 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t340 VOUT_P.t93 VDD.t778 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X712 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t59 VDD.t1294 VDD.t729 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X713 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t57 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t58 VDD.t641 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X714 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t37 VDD.t104 VDD.t78 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X715 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3.t34 Folded_Diff_Op_Amp_Layout_0.OUT2.t3 VSS.t249 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X716 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t342 VDD.t782 VDD.t781 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X717 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t343 VDD.t784 VDD.t783 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X718 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t344 VOUT_P.t92 VDD.t767 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X719 Folded_Diff_Op_Amp_Layout_0.IB3 Folded_Diff_Op_Amp_Layout_0.VB3.t4 Folded_Diff_Op_Amp_Layout_0.VB3.t5 VSS.t22 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X720 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t345 VOUT_P.t91 VDD.t1022 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X721 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t346 VDD.t1439 VDD.t666 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X722 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t20 Folded_Diff_Op_Amp_Layout_0.IPD.t10 VDD.t459 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X723 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t67 Folded_Diff_Op_Amp_Layout_0.IND.t20 VSS.t8 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X724 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t38 VDD.t105 VDD.t80 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X725 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t29 VDD.t47 VDD.t9 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X726 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3.t35 Folded_Diff_Op_Amp_Layout_0.IPD.t59 VSS.t28 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X727 VSS.t407 VSS.t406 VSS.t407 VSS.t352 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X728 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t347 VOUT_N.t268 VDD.t1030 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X729 a_n6546_7019.t1 a_n6826_6457.t1 VDD.t34 ppolyf_u r_width=1u r_length=2.3u
X730 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t348 VOUT_P.t90 VDD.t817 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X731 Folded_Diff_Op_Amp_Layout_0.IB3 Folded_Diff_Op_Amp_Layout_0.VB3.t2 Folded_Diff_Op_Amp_Layout_0.VB3.t3 VSS.t21 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X732 a_n6266_8433.t0 a_n5986_7871.t0 VDD.t0 ppolyf_u r_width=1u r_length=2.3u
X733 a_n5426_5540.t1 a_n5146_4623.t1 VDD.t114 ppolyf_u r_width=1u r_length=2.3u
X734 a_n7106_9350.t2 filter_res_magic_0.R3_R7.t7 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X735 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t48 Folded_Diff_Op_Amp_Layout_0.VPD.t8 VDD.t948 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X736 VDD.t290 VDD.t288 VDD.t290 VDD.t289 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X737 VSS Folded_Diff_Op_Amp_Layout_0.IBS.t3 Folded_Diff_Op_Amp_Layout_0.IBS.t4 VSS.t221 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X738 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t349 VDD.t1444 VDD.t822 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X739 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t30 Folded_Diff_Op_Amp_Layout_0.BD.t13 VDD.t11 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X740 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t73 VSS.t135 VSS.t108 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X741 a_n5706_8433.t1 a_n5426_7871.t1 VDD.t89 ppolyf_u r_width=1u r_length=2.3u
X742 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t55 VDD.t1291 VDD.t639 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X743 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VBIASN.t7 VSS.t518 VSS.t517 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X744 VDD.t287 VDD.t286 VDD.t287 VDD.t213 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X745 VDD.t285 VDD.t284 VDD.t285 VDD.t231 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X746 a_n7106_5185.t0 a_n6546_4623.t1 VDD.t34 ppolyf_u r_width=1u r_length=2.3u
X747 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3.t36 Folded_Diff_Op_Amp_Layout_0.IND.t34 VSS.t250 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X748 a_n7106_9350.t2 filter_res_magic_0.R3_R7.t6 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X749 VDD.t283 VDD.t281 VDD.t283 VDD.t282 pfet_03v3 ad=1.04p pd=4.52u as=0 ps=0 w=4u l=0.28u
X750 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t351 VOUT_N.t270 VDD.t1100 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X751 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t22 Folded_Diff_Op_Amp_Layout_0.BD.t59 VDD.t498 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X752 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3.t37 Folded_Diff_Op_Amp_Layout_0.OUT1.t7 VSS.t251 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X753 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t352 VDD.t1447 VDD.t1035 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X754 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t353 VDD.t1448 VDD.t925 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X755 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t10 VDD.t859 VDD.t524 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X756 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1.t49 VDD.t975 VDD.t963 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X757 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t39 Folded_Diff_Op_Amp_Layout_0.IVS.t0 VDD.t67 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X758 VDD.t479 VDD.t480 VDD.t40 ppolyf_u r_width=1u r_length=2.3u
X759 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t354 VOUT_P.t88 VDD.t817 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X760 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t53 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t54 VDD.t661 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X761 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t355 VOUT_P.t87 VDD.t698 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X762 VSS.t405 VSS.t404 VSS.t405 VSS.t320 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X763 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t356 VOUT_P.t86 VDD.t1201 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X764 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t357 VOUT_P.t85 VDD.t794 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X765 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t40 Folded_Diff_Op_Amp_Layout_0.IVS.t1 VDD.t67 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X766 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t358 VOUT_N.t239 VDD.t797 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X767 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t359 VDD.t1348 VDD.t781 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X768 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t51 VDD.t651 VDD.t650 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X769 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t361 VDD.t1349 VDD.t607 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X770 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3.t38 Folded_Diff_Op_Amp_Layout_0.OUT1.t8 VSS.t247 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X771 VDD.t280 VDD.t279 VDD.t280 VDD.t223 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X772 VSS.t403 VSS.t402 VSS.t403 VSS.t305 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X773 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t362 VOUT_N.t241 VDD.t800 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X774 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t68 VSS.t11 VSS.t3 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X775 VDD.t278 VDD.t277 VDD.t278 VDD.t226 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X776 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t71 VSS.t641 VSS.t185 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X777 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t74 VOUT_N.t18 VSS.t100 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X778 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t363 VDD.t1352 VDD.t806 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X779 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t364 VOUT_P.t82 VDD.t882 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X780 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t69 Folded_Diff_Op_Amp_Layout_0.IND.t18 VSS.t8 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X781 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t70 Folded_Diff_Op_Amp_Layout_0.IND.t17 VSS.t49 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X782 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t365 VOUT_P.t81 VDD.t866 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X783 VDD.t276 VDD.t275 VDD.t276 VDD.t179 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X784 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t72 VOUT_P.t236 VSS.t175 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X785 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t366 VDD.t869 VDD.t605 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X786 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1.t50 VDD.t976 VDD.t961 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X787 VDD.t274 VDD.t273 VDD.t274 VDD.t271 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X788 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t41 Folded_Diff_Op_Amp_Layout_0.IVS.t2 VDD.t72 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X789 VSS.t401 VSS.t400 VSS.t401 VSS.t302 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X790 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t14 Folded_Diff_Op_Amp_Layout_0.VB4.t15 VSS.t497 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X791 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t75 VOUT_N.t17 VSS.t67 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X792 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t76 VSS.t130 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X793 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t367 VDD.t871 VDD.t870 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X794 VDD.t272 VDD.t270 VDD.t272 VDD.t271 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X795 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t42 Folded_Diff_Op_Amp_Layout_0.IVS.t3 VDD.t75 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X796 VDD.t269 VDD.t267 VDD.t269 VDD.t268 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X797 VDD.t266 VDD.t264 VDD.t266 VDD.t265 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X798 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t368 VDD.t872 VDD.t615 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X799 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t12 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t13 VDD.t446 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X800 VDD.t263 VDD.t261 VDD.t263 VDD.t262 pfet_03v3 ad=1.04p pd=4.52u as=0 ps=0 w=4u l=0.28u
X801 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t51 Folded_Diff_Op_Amp_Layout_0.VPD.t7 VDD.t970 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X802 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t73 VOUT_P.t237 VSS.t182 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X803 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t369 VOUT_N.t119 VDD.t800 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X804 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t31 Folded_Diff_Op_Amp_Layout_0.BD.t12 VDD.t11 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X805 VDD.t260 VDD.t259 VDD.t260 VDD.t150 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X806 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t370 VOUT_P.t79 VDD.t617 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X807 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t43 VDD.t79 VDD.t78 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X808 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t12 Folded_Diff_Op_Amp_Layout_0.VB4.t13 VSS.t209 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X809 VSS.t399 VSS.t398 VSS.t399 VSS.t376 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X810 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t32 VDD.t466 VDD.t7 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X811 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3.t39 Folded_Diff_Op_Amp_Layout_0.IPD.t60 VSS.t252 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X812 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t49 VDD.t649 VDD.t639 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X813 VDD.t258 VDD.t256 VDD.t258 VDD.t257 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X814 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t372 VOUT_P.t78 VDD.t620 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X815 a_n5426_7019.t0 VOUT_OPAMP_N.t0 VDD.t55 ppolyf_u r_width=1u r_length=2.3u
X816 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t373 VDD.t879 VDD.t592 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X817 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t15 Folded_Diff_Op_Amp_Layout_0.VCD.t37 VSS.t263 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X818 VOUT_OPAMP_P.t5 VOUT_OPAMP_P.t6 VDD.t114 ppolyf_u r_width=1u r_length=2.3u
X819 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t44 VDD.t81 VDD.t80 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X820 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t45 VDD.t82 VDD.t78 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X821 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t71 Folded_Diff_Op_Amp_Layout_0.IPD.t38 VSS.t8 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X822 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t374 VOUT_N.t120 VDD.t629 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X823 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t375 VOUT_P.t76 VDD.t740 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X824 VDD.t255 VDD.t253 VDD.t255 VDD.t254 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X825 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t376 VDD.t1073 VDD.t693 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X826 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t21 Folded_Diff_Op_Amp_Layout_0.IPD.t9 VDD.t500 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X827 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t74 VOUT_P.t238 VSS.t175 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X828 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t377 VOUT_N.t163 VDD.t746 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X829 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t46 VDD.t83 VDD.t80 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X830 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t378 VOUT_N.t164 VDD.t695 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X831 VSS Folded_Diff_Op_Amp_Layout_0.VBIASN.t8 Folded_Diff_Op_Amp_Layout_0.VCD.t45 VSS.t519 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X832 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t72 VSS.t610 VSS.t206 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X833 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t83 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t120 VSS.t64 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X834 VDD.t252 VDD.t251 VDD.t252 VDD.t156 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X835 a_n6826_8433.t1 a_n6546_7871.t0 VDD.t34 ppolyf_u r_width=1u r_length=2.3u
X836 a_n7106_7019.t1 filter_res_magic_0.R7_R8_R10_C VDD.t90 ppolyf_u r_width=1u r_length=2.3u
X837 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t379 VOUT_P.t75 VDD.t755 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X838 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t380 VDD.t1080 VDD.t678 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X839 VDD.t250 VDD.t249 VDD.t250 VDD.t147 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X840 a_n5706_5185.t0 a_n5146_4623.t0 VDD.t55 ppolyf_u r_width=1u r_length=2.3u
X841 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t77 VSS.t128 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X842 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t381 VDD.t1081 VDD.t1041 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X843 VDD.t248 VDD.t247 VDD.t248 VDD.t213 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X844 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t382 VDD.t1082 VDD.t615 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X845 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t383 VOUT_P.t72 VDD.t620 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X846 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t75 VOUT_P.t239 VSS.t84 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X847 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t76 VOUT_P.t240 VSS.t75 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X848 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t384 VOUT_P.t71 VDD.t762 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X849 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t33 VDD.t865 VDD.t7 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X850 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2.t64 Folded_Diff_Op_Amp_Layout_0.VPD.t19 VDD.t584 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X851 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t47 VDD.t85 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X852 a_n7106_9350.t2 filter_res_magic_0.R3_R7.t5 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X853 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t11 VDD.t860 VDD.t524 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X854 a_26012_2845.t0 a_26292_1743.t0 VDD.t32 ppolyf_u r_width=1u r_length=5u
X855 a_27020_2845.t0 a_26740_1743.t0 VDD.t33 ppolyf_u r_width=1u r_length=5u
X856 a_n7106_9350.t3 filter_res_magic_0.R3_R7.t4 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X857 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.IBIAS.t6 VDD.t531 VDD.t530 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X858 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t22 Folded_Diff_Op_Amp_Layout_0.BD.t69 VDD.t469 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X859 VDD.t246 VDD.t244 VDD.t246 VDD.t245 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X860 a_n7106_5185.t1 VOUT_P.t0 VDD.t90 ppolyf_u r_width=1u r_length=2.3u
X861 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t12 VDD.t861 VDD.t524 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X862 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t18 Folded_Diff_Op_Amp_Layout_0.VB1.t13 VSS.t264 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X863 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t47 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t48 VDD.t646 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X864 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t45 VDD.t645 VDD.t644 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X865 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t386 VOUT_N.t175 VDD.t740 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X866 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t78 VOUT_N.t16 VSS.t72 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X867 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t387 VOUT_P.t70 VDD.t844 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X868 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t388 VDD.t1120 VDD.t1119 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X869 VDD.t243 VDD.t242 VDD.t243 VDD.t141 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X870 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t16 Folded_Diff_Op_Amp_Layout_0.VBM.t13 VSS.t277 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X871 VSS.t397 VSS.t396 VSS.t397 VSS.t352 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X872 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t389 VDD.t1121 VDD.t1051 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X873 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t48 VDD.t416 VDD.t398 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X874 VSS Folded_Diff_Op_Amp_Layout_0.IBS.t11 Folded_Diff_Op_Amp_Layout_0.IBIAS.t10 VSS.t61 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=1u
X875 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.VB2.t14 Folded_Diff_Op_Amp_Layout_0.VB2.t15 VDD.t566 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X876 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t390 VOUT_P.t67 VDD.t767 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X877 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t23 Folded_Diff_Op_Amp_Layout_0.BD.t70 VDD.t467 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X878 VDD.t241 VDD.t239 VDD.t241 VDD.t240 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X879 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t391 VDD.t1124 VDD.t1059 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X880 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t392 VOUT_P.t66 VDD.t773 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X881 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t393 VDD.t1127 VDD.t632 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X882 VSS.t395 VSS.t394 VSS.t395 VSS.t340 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X883 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t394 VDD.t1128 VDD.t776 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X884 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t395 VDD.t1129 VDD.t705 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X885 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t49 VDD.t417 VDD.t121 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X886 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t17 Folded_Diff_Op_Amp_Layout_0.VBM.t12 VSS.t278 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X887 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t73 Folded_Diff_Op_Amp_Layout_0.IND.t15 VSS.t0 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X888 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t396 VOUT_N.t178 VDD.t778 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X889 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t43 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t44 VDD.t641 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X890 Folded_Diff_Op_Amp_Layout_0.IB5 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t8 VDD.t465 VDD.t464 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X891 VDD.t238 VDD.t237 VDD.t238 VDD.t165 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X892 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t77 VSS.t652 VSS.t80 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X893 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t397 VDD.t1019 VDD.t781 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X894 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t398 VOUT_N.t146 VDD.t767 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X895 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t10 VDD.t451 VDD.t428 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X896 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t79 VOUT_N.t15 VSS.t116 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X897 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t399 VOUT_N.t147 VDD.t1022 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X898 a_24836_4817.t0 a_24556_3715.t0 VDD.t410 ppolyf_u r_width=1u r_length=5u
X899 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t400 VDD.t1025 VDD.t666 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X900 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t401 VOUT_P.t61 VDD.t922 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X901 VSS Folded_Diff_Op_Amp_Layout_0.VBIASN.t9 Folded_Diff_Op_Amp_Layout_0.VCD.t63 VSS.t622 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X902 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t78 VOUT_P.t242 VSS.t175 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X903 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t79 VSS.t655 VSS.t78 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X904 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t402 VOUT_N.t148 VDD.t1022 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X905 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t80 VOUT_N.t14 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X906 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IVS.t44 VSS.t534 VSS.t245 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X907 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t403 VOUT_P.t60 VDD.t1030 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X908 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t23 Folded_Diff_Op_Amp_Layout_0.IND.t64 VDD.t499 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X909 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t404 VOUT_P.t59 VDD.t609 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X910 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t19 Folded_Diff_Op_Amp_Layout_0.VCD.t5 VSS.t261 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X911 VSS.t393 VSS.t392 VSS.t393 VSS.t340 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X912 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1.t52 VDD.t979 VDD.t961 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X913 VDD.t236 VDD.t235 VDD.t236 VDD.t176 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X914 VSS.t391 VSS.t389 VSS.t391 VSS.t390 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X915 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t81 VOUT_N.t13 VSS.t67 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X916 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t80 VOUT_P.t244 VSS.t75 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X917 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t8 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t9 VDD.t446 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X918 a_n6546_7019.t0 a_n6266_6457.t1 VDD.t43 ppolyf_u r_width=1u r_length=2.3u
X919 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t81 VOUT_P.t245 VSS.t72 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X920 VSS.t388 VSS.t387 VSS.t388 VSS.t299 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X921 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t6 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t7 VDD.t446 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X922 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t41 VDD.t640 VDD.t639 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X923 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t18 Folded_Diff_Op_Amp_Layout_0.VCD.t40 VSS.t279 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X924 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t74 VSS.t613 VSS.t3 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X925 VDD.t234 VDD.t233 VDD.t234 VDD.t213 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X926 VDD.t232 VDD.t230 VDD.t232 VDD.t231 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X927 a_29734_1647.t1 VOUT_N.t0 cap_mim_2f0_m4m5_noshield c_width=21u c_length=21u
X928 VSS.t386 VSS.t385 VSS.t386 VSS.t376 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X929 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t82 VSS.t119 VSS.t98 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X930 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.t24 Folded_Diff_Op_Amp_Layout_0.IB2.t6 VDD.t571 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X931 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t82 VOUT_P.t246 VSS.t136 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X932 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t406 VDD.t1036 VDD.t1035 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X933 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t407 VDD.t1037 VDD.t925 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X934 VOUT_OPAMP_P.t4 a_n5426_7871.t0 VDD.t55 ppolyf_u r_width=1u r_length=2.3u
X935 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t75 Folded_Diff_Op_Amp_Layout_0.IND.t13 VSS.t49 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X936 VSS.t384 VSS.t383 VSS.t384 VSS.t290 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X937 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t39 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t40 VDD.t636 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X938 Folded_Diff_Op_Amp_Layout_0.IBIAS1 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t0 VDD.t510 VDD.t61 pfet_03v3 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.56u
X939 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t408 VOUT_N.t179 VDD.t817 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X940 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t51 Folded_Diff_Op_Amp_Layout_0.IVS.t60 VDD.t106 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X941 Folded_Diff_Op_Amp_Layout_0.IBS Folded_Diff_Op_Amp_Layout_0.IBIAS1.t10 VDD.t477 VDD.t476 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X942 a_n6826_5185.t1 a_n6266_4623.t1 VDD.t43 ppolyf_u r_width=1u r_length=2.3u
X943 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t37 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t38 VDD.t661 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X944 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t409 VDD.t1134 VDD.t1053 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X945 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t83 VOUT_N.t12 VSS.t116 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X946 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t410 VOUT_N.t181 VDD.t668 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X947 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t52 Folded_Diff_Op_Amp_Layout_0.IVS.t61 VDD.t109 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X948 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t83 VSS.t662 VSS.t149 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X949 Folded_Diff_Op_Amp_Layout_0.OUT2.t19 a_29734_3659.t3 VDD.t411 ppolyf_u r_width=1u r_length=6.2u
X950 VDD.t229 VDD.t228 VDD.t229 VDD.t218 pfet_03v3 ad=0.814p pd=3.65u as=0 ps=0 w=3.13u l=0.56u
X951 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3.t40 Folded_Diff_Op_Amp_Layout_0.OUT1.t9 VSS.t248 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X952 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t411 VOUT_N.t182 VDD.t929 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X953 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t412 VDD.t1139 VDD.t607 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X954 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t84 VSS.t663 VSS.t70 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X955 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t413 VDD.t1140 VDD.t870 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X956 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t414 VDD.t1141 VDD.t1059 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X957 a_n7106_8433.t1 a_n7106_7871.t0 VDD.t90 ppolyf_u r_width=1u r_length=2.3u
X958 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t85 VOUT_P.t249 VSS.t67 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X959 VDD.t227 VDD.t225 VDD.t227 VDD.t226 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X960 VSS Folded_Diff_Op_Amp_Layout_0.IVS.t85 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t119 VSS.t64 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X961 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t84 VSS.t115 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X962 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1.t53 VDD.t980 VDD.t963 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X963 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t85 VSS.t114 VSS.t113 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X964 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t19 Folded_Diff_Op_Amp_Layout_0.VBM.t10 VSS.t264 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X965 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t415 VOUT_N.t184 VDD.t882 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X966 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t416 VOUT_N.t185 VDD.t866 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X967 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t417 VOUT_P.t55 VDD.t770 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X968 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t418 VOUT_N.t248 VDD.t759 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X969 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t20 Folded_Diff_Op_Amp_Layout_0.VCD.t42 VSS.t280 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X970 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3.t41 Folded_Diff_Op_Amp_Layout_0.IND.t38 VSS.t252 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X971 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t419 VDD.t1374 VDD.t605 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X972 VSS.t382 VSS.t380 VSS.t382 VSS.t381 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X973 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3.t42 Folded_Diff_Op_Amp_Layout_0.OUT1.t11 VSS.t249 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X974 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t76 Folded_Diff_Op_Amp_Layout_0.IND.t12 VSS.t49 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X975 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t77 VSS.t236 VSS.t206 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X976 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.t6 Folded_Diff_Op_Amp_Layout_0.IB2.t5 VDD.t562 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X977 VDD.t224 VDD.t222 VDD.t224 VDD.t223 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X978 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t86 VSS.t666 VSS.t185 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X979 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t20 Folded_Diff_Op_Amp_Layout_0.VB1.t11 VSS.t278 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X980 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t420 VDD.t1375 VDD.t870 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X981 VSS.t379 VSS.t378 VSS.t379 VSS.t343 nfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=1u
X982 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t35 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t36 VDD.t641 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X983 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t21 Folded_Diff_Op_Amp_Layout_0.VCD.t4 VSS.t260 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X984 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t421 VDD.t1376 VDD.t664 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X985 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VBIASN.t10 VSS.t626 VSS.t625 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X986 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t78 VSS.t237 VSS.t206 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X987 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t87 VSS.t667 VSS.t156 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X988 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t422 VDD.t1377 VDD.t671 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X989 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t423 VOUT_P.t51 VDD.t673 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X990 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t424 VOUT_P.t50 VDD.t800 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X991 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t32 Folded_Diff_Op_Amp_Layout_0.VB1.t33 VDD.t940 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X992 VDD.t221 VDD.t220 VDD.t221 VDD.t150 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X993 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t425 VDD.t1382 VDD.t676 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X994 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t86 VSS.t112 VSS.t87 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X995 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t426 VDD.t1383 VDD.t678 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X996 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t22 Folded_Diff_Op_Amp_Layout_0.VCD.t3 VSS.t263 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X997 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t427 VDD.t1384 VDD.t592 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X998 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t88 VSS.t668 VSS.t149 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X999 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t428 VOUT_N.t95 VDD.t740 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1000 VSS.t377 VSS.t375 VSS.t377 VSS.t376 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X1001 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t429 VDD.t743 VDD.t693 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1002 VSS.t374 VSS.t373 VSS.t374 VSS.t299 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1003 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t430 VOUT_N.t96 VDD.t688 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1004 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t4 Folded_Diff_Op_Amp_Layout_0.IBIAS.t5 VDD.t862 pfet_03v3 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.56u
X1005 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t54 Folded_Diff_Op_Amp_Layout_0.VPD.t5 VDD.t970 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X1006 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t431 VOUT_P.t47 VDD.t746 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1007 VDD.t59 VDD.t60 VDD.t40 ppolyf_u r_width=1u r_length=2.3u
X1008 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3.t43 Folded_Diff_Op_Amp_Layout_0.OUT2.t6 VSS.t251 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X1009 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t87 VSS.t111 VSS.t78 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1010 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t432 VOUT_P.t46 VDD.t695 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1011 a_29734_3659.t5 VOUT_P.t226 cap_mim_2f0_m4m5_noshield c_width=21u c_length=21u
X1012 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IVS.t42 VSS.t533 VSS.t245 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X1013 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t79 VSS.t238 VSS.t56 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1014 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t88 VSS.t110 VSS.t70 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1015 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t433 VOUT_P.t45 VDD.t688 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1016 VDD.t219 VDD.t217 VDD.t219 VDD.t218 pfet_03v3 ad=0.814p pd=3.65u as=0 ps=0 w=3.13u l=0.56u
X1017 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t434 VOUT_P.t44 VDD.t707 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1018 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t435 VOUT_N.t97 VDD.t755 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1019 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t436 VDD.t758 VDD.t678 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1020 Folded_Diff_Op_Amp_Layout_0.VOUT.t1 a_24108_3715.t1 VDD.t491 ppolyf_u r_width=1u r_length=5u
X1021 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t23 Folded_Diff_Op_Amp_Layout_0.VB1.t8 VSS.t262 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1022 VDD.t216 VDD.t215 VDD.t216 VDD.t202 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.56u
X1023 VDD.t214 VDD.t212 VDD.t214 VDD.t213 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1024 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.VB2.t12 Folded_Diff_Op_Amp_Layout_0.VB2.t13 VDD.t565 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1025 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3.t44 Folded_Diff_Op_Amp_Layout_0.OUT2.t7 VSS.t249 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1026 VDD.t211 VDD.t210 VDD.t211 VDD.t176 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1027 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t437 VOUT_P.t43 VDD.t759 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1028 a_n6266_8433.t1 a_n6546_7871.t1 VDD.t43 ppolyf_u r_width=1u r_length=2.3u
X1029 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t438 VOUT_N.t99 VDD.t762 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1030 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t439 VOUT_N.t218 VDD.t620 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1031 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t440 VDD.t1271 VDD.t1005 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1032 VSS Folded_Diff_Op_Amp_Layout_0.IB4.t23 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t17 VSS.t64 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X1033 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3.t45 Folded_Diff_Op_Amp_Layout_0.OUT2.t16 VSS.t247 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1034 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t89 VSS.t109 VSS.t108 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1035 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t441 VDD.t1272 VDD.t813 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1036 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t33 VDD.t658 VDD.t657 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1037 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t21 Folded_Diff_Op_Amp_Layout_0.VBM.t8 VSS.t281 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1038 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t35 Folded_Diff_Op_Amp_Layout_0.BD.t9 VDD.t4 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1039 VDD.t209 VDD.t207 VDD.t209 VDD.t208 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X1040 VDD.t414 VDD.t415 VDD.t40 ppolyf_u r_width=1u r_length=2.3u
X1041 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t90 VSS.t107 VSS.t98 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1042 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t443 VOUT_P.t41 VDD.t740 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1043 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t444 VOUT_N.t220 VDD.t849 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1044 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t24 Folded_Diff_Op_Amp_Layout_0.BD.t71 VDD.t460 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1045 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t91 VOUT_N.t11 VSS.t92 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1046 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t89 VOUT_P.t253 VSS.t92 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1047 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t445 VOUT_N.t221 VDD.t844 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1048 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t446 VDD.t1279 VDD.t1119 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1049 VDD.t206 VDD.t204 VDD.t206 VDD.t205 pfet_03v3 ad=1.04p pd=4.52u as=0 ps=0 w=4u l=0.28u
X1050 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2.t67 Folded_Diff_Op_Amp_Layout_0.VND.t18 VDD.t584 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X1051 VOUT_N.t273 VOUT_OPAMP_P.t0 cap_mim_2f0_m4m5_noshield c_width=15.2u c_length=16u
X1052 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t24 Folded_Diff_Op_Amp_Layout_0.VCD.t2 VSS.t280 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1053 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3.t46 Folded_Diff_Op_Amp_Layout_0.OUT1.t18 VSS.t247 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1054 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t92 VSS.t104 VSS.t103 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1055 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t447 VDD.t1280 VDD.t1059 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1056 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t448 VOUT_N.t223 VDD.t1012 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1057 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t449 VDD.t1283 VDD.t632 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1058 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t450 VDD.t1284 VDD.t705 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1059 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t451 VDD.t1172 VDD.t1016 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1060 VDD.t203 VDD.t201 VDD.t203 VDD.t202 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.56u
X1061 VSS.t372 VSS.t371 VSS.t372 VSS.t314 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1062 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t452 VDD.t1173 VDD.t701 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1063 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t24 Folded_Diff_Op_Amp_Layout_0.BD.t61 VDD.t458 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X1064 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t25 Folded_Diff_Op_Amp_Layout_0.BD.t62 VDD.t457 pfet_03v3 ad=1.65p pd=8.38u as=0.975p ps=4.27u w=3.75u l=0.28u
X1065 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB2.t68 Folded_Diff_Op_Amp_Layout_0.OUT1.t34 VDD.t576 pfet_03v3 ad=1.38p pd=7.14u as=1.38p ps=7.14u w=3.13u l=0.28u
X1066 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t93 VOUT_N.t10 VSS.t100 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1067 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t31 VDD.t656 VDD.t644 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1068 filter_res_magic_0.R7_R8_R10_C.t0 a_n7106_8433.t3 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X1069 VSS.t370 VSS.t369 VSS.t370 VSS.t293 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1070 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t90 VOUT_P.t254 VSS.t182 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1071 Folded_Diff_Op_Amp_Layout_0.OUT2.t0 a_29734_3659.t0 VDD.t412 ppolyf_u r_width=1u r_length=6.2u
X1072 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t25 Folded_Diff_Op_Amp_Layout_0.VB1.t6 VSS.t264 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1073 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t22 Folded_Diff_Op_Amp_Layout_0.VCD.t55 VSS.t260 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1074 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t454 VOUT_P.t37 VDD.t1022 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1075 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t455 VOUT_N.t193 VDD.t922 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1076 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t456 VDD.t1178 VDD.t831 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1077 Folded_Diff_Op_Amp_Layout_0.VOUT.t0 a_24556_3715.t1 VDD.t488 ppolyf_u r_width=1u r_length=5u
X1078 VDD.t200 VDD.t199 VDD.t200 VDD.t144 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1079 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t457 VOUT_N.t195 VDD.t609 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1080 Folded_Diff_Op_Amp_Layout_0.OUT2.t14 a_29734_3659.t1 VDD.t66 ppolyf_u r_width=1u r_length=6.2u
X1081 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t23 Folded_Diff_Op_Amp_Layout_0.VBM.t6 VSS.t278 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1082 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t80 VSS.t239 VSS.t204 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1083 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t81 Folded_Diff_Op_Amp_Layout_0.IPD.t35 VSS.t5 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1084 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t91 VOUT_P.t255 VSS.t140 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1085 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t92 VSS.t675 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1086 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB2.t69 Folded_Diff_Op_Amp_Layout_0.OUT2.t26 VDD.t578 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1087 VDD.t198 VDD.t197 VDD.t198 VDD.t168 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1088 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IB4.t0 VSS.t246 VSS.t245 nfet_03v3 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=1u
X1089 VSS.t368 VSS.t367 VSS.t368 VSS.t343 nfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=1u
X1090 VSS.t366 VSS.t364 VSS.t366 VSS.t365 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X1091 VSS.t363 VSS.t362 VSS.t363 VSS.t352 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1092 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t94 VSS.t99 VSS.t98 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1093 VSS.t361 VSS.t360 VSS.t361 VSS.t317 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X1094 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t26 Folded_Diff_Op_Amp_Layout_0.IND.t67 VDD.t459 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1095 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t458 VDD.t1181 VDD.t1016 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1096 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t459 VOUT_P.t36 VDD.t895 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1097 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t36 Folded_Diff_Op_Amp_Layout_0.BD.t8 VDD.t4 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1098 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1.t55 VDD.t983 VDD.t961 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1099 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t460 VOUT_N.t197 VDD.t828 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1100 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t24 Folded_Diff_Op_Amp_Layout_0.VBM.t5 VSS.t262 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1101 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t93 VSS.t676 VSS.t149 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1102 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t29 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t30 VDD.t636 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1103 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t461 VOUT_N.t198 VDD.t612 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1104 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t10 Folded_Diff_Op_Amp_Layout_0.VB4.t11 VSS.t265 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1105 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t462 VOUT_P.t35 VDD.t668 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1106 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t463 VDD.t1054 VDD.t1053 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1107 VDD.t196 VDD.t195 VDD.t196 VDD.t179 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1108 VSS.t359 VSS.t358 VSS.t359 VSS.t311 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X1109 VSS.t357 VSS.t356 VSS.t357 VSS.t314 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1110 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t464 VOUT_P.t33 VDD.t929 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1111 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t465 VDD.t1057 VDD.t826 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1112 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t53 Folded_Diff_Op_Amp_Layout_0.IVS.t62 VDD.t72 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1113 VSS.t355 VSS.t354 VSS.t355 VSS.t327 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X1114 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t26 Folded_Diff_Op_Amp_Layout_0.VB1.t5 VSS.t281 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1115 VDD.t41 VDD.t42 VDD.t40 ppolyf_u r_width=1u r_length=2.3u
X1116 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t95 VSS.t97 VSS.t70 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1117 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t466 VDD.t1058 VDD.t870 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1118 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t467 VDD.t1060 VDD.t1059 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1119 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VB3.t10 Folded_Diff_Op_Amp_Layout_0.IB3.t1 VSS.t25 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1120 VSS.t353 VSS.t351 VSS.t353 VSS.t352 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1121 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t468 VOUT_P.t31 VDD.t617 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1122 VSS.t350 VSS.t349 VSS.t350 VSS.t302 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1123 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t96 VOUT_N.t9 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1124 VSS.t348 VSS.t347 VSS.t348 VSS.t290 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1125 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t25 Folded_Diff_Op_Amp_Layout_0.BD.t72 VDD.t498 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1126 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t469 VDD.t1063 VDD.t783 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1127 VDD.t194 VDD.t193 VDD.t194 VDD.t159 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1128 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t54 Folded_Diff_Op_Amp_Layout_0.IVS.t63 VDD.t75 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1129 VSS.t346 VSS.t345 VSS.t346 VSS.t340 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1130 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t470 VOUT_N.t160 VDD.t770 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1131 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t471 VOUT_P.t30 VDD.t759 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1132 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t472 VDD.t1068 VDD.t847 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1133 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t94 VOUT_P.t258 VSS.t136 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1134 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t473 VOUT_P.t29 VDD.t849 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1135 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t27 Folded_Diff_Op_Amp_Layout_0.IND.t68 VDD.t501 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X1136 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t97 VOUT_N.t8 VSS.t92 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1137 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t27 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t28 VDD.t641 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1138 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t474 VDD.t665 VDD.t664 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1139 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t475 VDD.t667 VDD.t666 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1140 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t476 VOUT_P.t27 VDD.t668 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1141 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t477 VDD.t672 VDD.t671 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1142 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t478 VOUT_N.t87 VDD.t673 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1143 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t25 Folded_Diff_Op_Amp_Layout_0.VCD.t58 VSS.t280 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1144 VDD.t513 VDD.t514 VDD.t115 ppolyf_u r_width=1u r_length=5u
X1145 VSS.t344 VSS.t342 VSS.t344 VSS.t343 nfet_03v3 ad=0.52p pd=2.52u as=0 ps=0 w=2u l=1u
X1146 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t479 VDD.t677 VDD.t676 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1147 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t480 VDD.t679 VDD.t678 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1148 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t481 VDD.t681 VDD.t680 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1149 VDD.t192 VDD.t191 VDD.t192 VDD.t150 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1150 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t482 VOUT_N.t89 VDD.t682 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1151 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t483 VOUT_P.t23 VDD.t685 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1152 a_n7106_9350.t3 filter_res_magic_0.R3_R7.t3 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X1153 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB4.t8 VSS.t259 VSS.t258 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1154 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t26 Folded_Diff_Op_Amp_Layout_0.IPD.t4 VDD.t461 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1155 VSS.t341 VSS.t339 VSS.t341 VSS.t340 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1156 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t25 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t26 VDD.t714 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1157 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t27 Folded_Diff_Op_Amp_Layout_0.VCD.t1 VSS.t260 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1158 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t83 VSS.t505 VSS.t204 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1159 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2.t70 Folded_Diff_Op_Amp_Layout_0.VPD.t17 VDD.t575 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X1160 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t484 VOUT_P.t22 VDD.t688 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1161 VSS.t338 VSS.t337 VSS.t338 VSS.t317 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X1162 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t56 Folded_Diff_Op_Amp_Layout_0.VND.t5 VDD.t943 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1163 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t84 Folded_Diff_Op_Amp_Layout_0.IPD.t33 VSS.t49 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1164 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t95 VSS.t679 VSS.t108 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1165 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t485 VOUT_N.t90 VDD.t688 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1166 VDD.t190 VDD.t189 VDD.t190 VDD.t147 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1167 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t23 VDD.t1253 VDD.t712 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1168 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t55 VDD.t426 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1169 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IVS.t87 VSS.t559 VSS.t19 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1170 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t487 VOUT_N.t139 VDD.t707 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1171 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t488 VDD.t1001 VDD.t898 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1172 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t96 VSS.t680 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1173 VDD.t87 VDD.t88 VDD.t86 ppolyf_u r_width=1u r_length=5u
X1174 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t37 VDD.t509 VDD.t26 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1175 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t489 VOUT_N.t140 VDD.t759 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1176 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t57 Folded_Diff_Op_Amp_Layout_0.VPD.t3 VDD.t948 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1177 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t56 VDD.t427 VDD.t398 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1178 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t28 Folded_Diff_Op_Amp_Layout_0.BD.t65 VDD.t468 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1179 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t490 VDD.t1004 VDD.t813 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1180 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t21 VDD.t1252 VDD.t657 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1181 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t492 VDD.t1006 VDD.t1005 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1182 VSS.t336 VSS.t335 VSS.t336 VSS.t311 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X1183 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB4.t6 VSS.t568 VSS.t567 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1184 VSS.t334 VSS.t333 VSS.t334 VSS.t320 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1185 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t493 VOUT_N.t142 VDD.t755 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1186 Folded_Diff_Op_Amp_Layout_0.IB3 Folded_Diff_Op_Amp_Layout_0.VB3.t48 VSS.t288 VSS.t287 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X1187 VDD.t188 VDD.t187 VDD.t188 VDD.t141 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1188 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t57 VDD.t122 VDD.t121 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1189 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t28 Folded_Diff_Op_Amp_Layout_0.VB1.t3 VSS.t262 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1190 VDD.t186 VDD.t185 VDD.t186 VDD.t156 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X1191 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t494 VOUT_P.t19 VDD.t849 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1192 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3.t49 Folded_Diff_Op_Amp_Layout_0.IPD.t70 VSS.t252 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X1193 VSS.t332 VSS.t331 VSS.t332 VSS.t305 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1194 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t495 VDD.t1011 VDD.t634 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1195 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t4 VDD.t445 VDD.t428 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1196 VDD.t184 VDD.t183 VDD.t184 VDD.t179 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1197 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P.t27 Folded_Diff_Op_Amp_Layout_0.BD.t74 VDD.t462 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1198 VDD.t182 VDD.t181 VDD.t182 VDD.t176 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1199 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t86 Folded_Diff_Op_Amp_Layout_0.IPD.t32 VSS.t49 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1200 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t87 VSS.t510 VSS.t206 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1201 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t97 VOUT_P.t261 VSS.t100 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1202 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t59 Folded_Diff_Op_Amp_Layout_0.IVS.t21 VDD.t72 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1203 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t11 VDD.t120 VDD.t119 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1204 VDD.t180 VDD.t178 VDD.t180 VDD.t179 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1205 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t496 VOUT_P.t17 VDD.t1012 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1206 VSS.t330 VSS.t329 VSS.t330 VSS.t305 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1207 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t497 VDD.t1015 VDD.t701 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1208 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t498 VDD.t1017 VDD.t1016 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1209 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t60 Folded_Diff_Op_Amp_Layout_0.IVS.t22 VDD.t72 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1210 VSS.t328 VSS.t326 VSS.t328 VSS.t327 nfet_03v3 ad=0.88p pd=4.88u as=0 ps=0 w=2u l=1u
X1211 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t26 Folded_Diff_Op_Amp_Layout_0.VBM.t3 VSS.t281 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1212 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t27 Folded_Diff_Op_Amp_Layout_0.VBM.t2 VSS.t277 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1213 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t88 Folded_Diff_Op_Amp_Layout_0.IND.t9 VSS.t5 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1214 VOUT_P.t272 VOUT_OPAMP_N.t6 cap_mim_2f0_m4m5_noshield c_width=15.2u c_length=16u
X1215 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t61 Folded_Diff_Op_Amp_Layout_0.IVS.t23 VDD.t75 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1216 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N.t29 Folded_Diff_Op_Amp_Layout_0.BD.t66 VDD.t469 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1217 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t19 VDD.t1251 VDD.t644 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1218 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t500 VDD.t1018 VDD.t710 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1219 VDD.t474 VDD.t475 VDD.t473 ppolyf_u r_width=1u r_length=6.2u
X1220 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t89 VSS.t513 VSS.t206 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1221 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1.t58 VDD.t988 VDD.t951 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1222 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t98 VOUT_N.t7 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1223 VSS.t325 VSS.t324 VSS.t325 VSS.t290 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1224 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t99 VSS.t88 VSS.t87 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1225 VDD.t177 VDD.t175 VDD.t177 VDD.t176 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1226 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t98 VSS.t683 VSS.t129 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1227 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t501 VDD.t1355 VDD.t776 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1228 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t62 Folded_Diff_Op_Amp_Layout_0.IVS.t24 VDD.t75 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1229 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t502 VOUT_N.t243 VDD.t673 pfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1230 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t28 Folded_Diff_Op_Amp_Layout_0.IPD.t2 VDD.t463 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1231 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t503 VDD.t1358 VDD.t831 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1232 a_25284_4817.t0 a_25564_3715.t0 VDD.t53 ppolyf_u r_width=1u r_length=5u
X1233 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IVS.t40 VSS.t532 VSS.t527 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1234 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t99 VOUT_P.t263 VSS.t136 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1235 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t90 Folded_Diff_Op_Amp_Layout_0.IPD.t29 VSS.t0 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1236 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t504 VDD.t1359 VDD.t1205 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1237 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t505 VOUT_N.t244 VDD.t835 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1238 Folded_Diff_Op_Amp_Layout_0.OUT2.t15 a_29734_3659.t2 VDD.t139 ppolyf_u r_width=1u r_length=6.2u
X1239 VDD.t492 VDD.t493 VDD.t430 ppolyf_u r_width=1u r_length=6.2u
X1240 VDD.t174 VDD.t173 VDD.t174 VDD.t144 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1241 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t17 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t18 VDD.t636 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1242 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1.t59 VDD.t989 VDD.t946 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1243 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t506 VDD.t1362 VDD.t910 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1244 VDD.t172 VDD.t170 VDD.t172 VDD.t171 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X1245 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t91 VSS.t550 VSS.t206 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1246 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t507 VDD.t1363 VDD.t1053 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1247 VDD.t169 VDD.t167 VDD.t169 VDD.t168 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1248 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t508 VDD.t1364 VDD.t806 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1249 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t509 VOUT_N.t246 VDD.t626 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1250 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t4 Folded_Diff_Op_Amp_Layout_0.VB4.t5 VSS.t242 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1251 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS1.t12 Folded_Diff_Op_Amp_Layout_0.VB3.t14 VDD.t504 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1252 VDD.t166 VDD.t164 VDD.t166 VDD.t165 pfet_03v3 ad=1.65p pd=8.38u as=0 ps=0 w=3.75u l=0.28u
X1253 VSS.t323 VSS.t322 VSS.t323 VSS.t314 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1254 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t63 Folded_Diff_Op_Amp_Layout_0.IVS.t25 VDD.t106 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1255 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.t0 Folded_Diff_Op_Amp_Layout_0.IB2.t3 VDD.t559 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1256 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t38 VDD.t558 VDD.t26 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1257 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t92 VSS.t551 VSS.t56 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1258 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t93 Folded_Diff_Op_Amp_Layout_0.IND.t7 VSS.t0 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1259 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT.t29 Folded_Diff_Op_Amp_Layout_0.VCD.t0 VSS.t261 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1260 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t39 Folded_Diff_Op_Amp_Layout_0.BD.t5 VDD.t17 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1261 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t510 VOUT_P.t12 VDD.t1201 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1262 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t511 VDD.t1369 VDD.t1016 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1263 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t64 Folded_Diff_Op_Amp_Layout_0.IVS.t26 VDD.t109 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1264 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VB3.t8 Folded_Diff_Op_Amp_Layout_0.IB3.t0 VSS.t24 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1265 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t512 VOUT_N.t247 VDD.t895 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1266 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t513 VDD.t827 VDD.t826 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1267 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3.t51 Folded_Diff_Op_Amp_Layout_0.IND.t62 VSS.t252 nfet_03v3 ad=1.27p pd=6.64u as=1.27p ps=6.64u w=2.88u l=0.28u
X1268 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t514 VOUT_P.t10 VDD.t828 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1269 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t515 VDD.t832 VDD.t831 pfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1270 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t29 Folded_Diff_Op_Amp_Layout_0.IPD.t1 VDD.t499 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1271 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t15 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t16 VDD.t646 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1272 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t65 Folded_Diff_Op_Amp_Layout_0.IVS.t27 VDD.t135 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1273 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t516 VOUT_P.t8 VDD.t612 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1274 Folded_Diff_Op_Amp_Layout_0.VBM VCM1.t28 Folded_Diff_Op_Amp_Layout_0.VCD.t61 VSS.t279 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1275 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t60 Folded_Diff_Op_Amp_Layout_0.VND.t3 VDD.t970 pfet_03v3 ad=0.814p pd=3.65u as=1.38p ps=7.14u w=3.13u l=0.28u
X1276 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t517 VOUT_P.t7 VDD.t835 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1277 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t66 VDD.t138 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1278 VSS.t321 VSS.t319 VSS.t321 VSS.t320 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1279 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t518 VDD.t839 VDD.t838 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1280 a_n7106_9350.t2 filter_res_magic_0.R3_R7.t2 cap_mim_2f0_m4m5_noshield c_width=16.2u c_length=15u
X1281 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VBIASN.t11 VSS.t628 VSS.t627 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X1282 VSS.t318 VSS.t316 VSS.t318 VSS.t317 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X1283 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t100 VSS.t686 VSS.t108 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1284 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t100 VOUT_N.t6 VSS.t84 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1285 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t101 VOUT_N.t5 VSS.t75 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1286 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t519 VDD.t840 VDD.t826 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1287 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t67 VDD.t397 VDD.t84 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1288 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P.t30 Folded_Diff_Op_Amp_Layout_0.IPD.t0 VDD.t456 pfet_03v3 ad=0.975p pd=4.27u as=0.975p ps=4.27u w=3.75u l=0.28u
X1289 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t61 Folded_Diff_Op_Amp_Layout_0.VPD.t1 VDD.t943 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1290 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB2.t72 Folded_Diff_Op_Amp_Layout_0.OUT1.t35 VDD.t574 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1291 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t520 VOUT_N.t114 VDD.t617 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1292 a_26292_4817.t1 a_27020_2845.t1 VDD.t413 ppolyf_u r_width=1u r_length=5u
X1293 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IVS.t89 VSS.t20 VSS.t19 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1294 VDD.t163 VDD.t161 VDD.t163 VDD.t162 pfet_03v3 ad=1.38p pd=7.14u as=0 ps=0 w=3.13u l=0.28u
X1295 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t68 VDD.t399 VDD.t398 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1296 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t521 VDD.t843 VDD.t783 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1297 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t522 VOUT_N.t115 VDD.t844 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1298 VDD.t160 VDD.t158 VDD.t160 VDD.t159 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1299 VSS Folded_Diff_Op_Amp_Layout_0.VBIASN.t12 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t4 VSS.t327 nfet_03v3 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=1u
X1300 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t40 Folded_Diff_Op_Amp_Layout_0.BD.t4 VDD.t17 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1301 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS1.t13 Folded_Diff_Op_Amp_Layout_0.IB5.t8 VDD.t61 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1302 VSS.t315 VSS.t313 VSS.t315 VSS.t314 nfet_03v3 ad=1.27p pd=6.64u as=0 ps=0 w=2.88u l=0.28u
X1303 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t94 Folded_Diff_Op_Amp_Layout_0.IPD.t27 VSS.t8 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1304 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t95 VSS.t556 VSS.t3 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1305 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t101 VOUT_P.t265 VSS.t72 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1306 a_26740_4817.t1 a_25564_3715.t1 VDD.t54 ppolyf_u r_width=1u r_length=5u
X1307 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t69 VDD.t400 VDD.t121 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1308 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t70 VDD.t401 VDD.t398 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1309 VDD.t157 VDD.t155 VDD.t157 VDD.t156 pfet_03v3 ad=0.22p pd=1.88u as=0 ps=0 w=0.5u l=0.28u
X1310 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t2 Folded_Diff_Op_Amp_Layout_0.IBIAS.t3 VDD.t587 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1311 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t523 VDD.t848 VDD.t847 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1312 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t13 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t14 VDD.t721 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1313 Folded_Diff_Op_Amp_Layout_0.VCD VCM1.t29 Folded_Diff_Op_Amp_Layout_0.VBM.t0 VSS.t264 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1314 VDD Folded_Diff_Op_Amp_Layout_0.VB1.t62 Folded_Diff_Op_Amp_Layout_0.VND.t2 VDD.t948 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1315 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t524 VOUT_N.t116 VDD.t849 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1316 VSS.t312 VSS.t310 VSS.t312 VSS.t311 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X1317 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N.t30 Folded_Diff_Op_Amp_Layout_0.IND.t71 VDD.t470 pfet_03v3 ad=0.975p pd=4.27u as=1.65p ps=8.38u w=3.75u l=0.28u
X1318 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t2 VDD.t444 VDD.t428 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1319 VSS.t309 VSS.t307 VSS.t309 VSS.t308 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.28u
X1320 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.VB2.t10 Folded_Diff_Op_Amp_Layout_0.VB2.t11 VDD.t564 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1321 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t72 VDD.t402 VDD.t121 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1322 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IVS.t90 VSS.t617 VSS.t14 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1323 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4.t96 VSS.t268 VSS.t204 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1324 VSS.t306 VSS.t304 VSS.t306 VSS.t305 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1325 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t525 VOUT_N.t121 VDD.t882 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1326 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t526 VDD.t886 VDD.t885 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1327 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t97 VSS.t269 VSS.t56 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1328 VSS.t303 VSS.t301 VSS.t303 VSS.t302 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1329 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t527 VDD.t887 VDD.t666 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1330 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t0 VDD.t429 VDD.t428 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1331 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t41 Folded_Diff_Op_Amp_Layout_0.BD.t3 VDD.t23 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1332 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1.t63 VDD.t996 VDD.t951 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1333 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t102 VSS.t81 VSS.t80 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1334 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t528 VOUT_N.t123 VDD.t668 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1335 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t30 Folded_Diff_Op_Amp_Layout_0.VB1.t1 VSS.t278 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1336 VDD.t154 VDD.t152 VDD.t154 VDD.t153 pfet_03v3 ad=1.76p pd=8.88u as=0 ps=0 w=4u l=0.28u
X1337 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t102 VOUT_P.t266 VSS.t116 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1338 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t103 VOUT_P.t267 VSS.t100 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1339 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t74 VDD.t404 VDD.t403 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1340 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.VB2.t8 Folded_Diff_Op_Amp_Layout_0.VB2.t9 VDD.t563 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X1341 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4.t98 VSS.t270 VSS.t204 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1342 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t99 Folded_Diff_Op_Amp_Layout_0.IPD.t25 VSS.t5 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1343 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t103 VSS.t79 VSS.t78 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1344 VDD.t151 VDD.t149 VDD.t151 VDD.t150 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1345 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t529 VOUT_P.t3 VDD.t682 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1346 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t530 VOUT_N.t124 VDD.t685 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1347 VOUT_P.t273 VOUT_OPAMP_N.t5 cap_mim_2f0_m4m5_noshield c_width=15.2u c_length=16u
X1348 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t104 VOUT_P.t268 VSS.t89 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1349 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t531 VDD.t894 VDD.t680 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1350 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t11 VDD.t720 VDD.t719 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1351 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IBIAS3.t75 VDD.t405 VDD.t93 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1352 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t9 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t10 VDD.t714 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1353 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t104 VOUT_N.t4 VSS.t75 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1354 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1.t64 VDD.t997 VDD.t951 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1355 VSS Folded_Diff_Op_Amp_Layout_0.VBIASN.t13 Folded_Diff_Op_Amp_Layout_0.VCD.t46 VSS.t524 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X1356 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t42 VDD.t527 VDD.t15 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1357 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t105 VOUT_N.t3 VSS.t72 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1358 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t533 VOUT_N.t126 VDD.t895 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1359 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t7 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t8 VDD.t714 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1360 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IVS.t38 VSS.t531 VSS.t527 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1361 VSS.t300 VSS.t298 VSS.t300 VSS.t299 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1362 VDD.t148 VDD.t146 VDD.t148 VDD.t147 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1363 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t5 VDD.t713 VDD.t712 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1364 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB2.t73 Folded_Diff_Op_Amp_Layout_0.OUT2.t25 VDD.t577 pfet_03v3 ad=1.38p pd=7.14u as=0.814p ps=3.65u w=3.13u l=0.28u
X1365 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t105 VOUT_P.t269 VSS.t175 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1366 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS.t43 Folded_Diff_Op_Amp_Layout_0.BD.t1 VDD.t23 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1367 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t535 VDD.t899 VDD.t898 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1368 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t536 VDD.t901 VDD.t900 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1369 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t76 Folded_Diff_Op_Amp_Layout_0.IVS.t36 VDD.t106 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1370 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t537 VDD.t902 VDD.t885 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1371 VOUT_P Folded_Diff_Op_Amp_Layout_0.IBIAS2.t538 VDD.t903 VDD.t693 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1372 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1.t65 VDD.t998 VDD.t946 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.28u
X1373 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t77 Folded_Diff_Op_Amp_Layout_0.IVS.t37 VDD.t109 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1374 VSS.t297 VSS.t295 VSS.t297 VSS.t296 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.28u
X1375 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t100 Folded_Diff_Op_Amp_Layout_0.IND.t3 VSS.t5 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1376 VSS.t294 VSS.t292 VSS.t294 VSS.t293 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1377 VSS.t291 VSS.t289 VSS.t291 VSS.t290 nfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1378 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t78 Folded_Diff_Op_Amp_Layout_0.IVS.t17 VDD.t106 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1379 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t101 Folded_Diff_Op_Amp_Layout_0.IND.t2 VSS.t5 nfet_03v3 ad=0.749p pd=3.4u as=1.27p ps=6.64u w=2.88u l=0.28u
X1380 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IB4.t25 VSS.t29 VSS.t19 nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=1u
X1381 a_n6266_6102.t0 a_n5706_5540.t0 VDD.t44 ppolyf_u r_width=1u r_length=2.3u
X1382 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3.t52 Folded_Diff_Op_Amp_Layout_0.IPD.t71 VSS.t27 nfet_03v3 ad=1.27p pd=6.64u as=0.749p ps=3.4u w=2.88u l=0.28u
X1383 VSS Folded_Diff_Op_Amp_Layout_0.OUT2.t106 VOUT_P.t270 VSS.t116 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1384 VDD.t145 VDD.t143 VDD.t145 VDD.t144 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1385 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t79 Folded_Diff_Op_Amp_Layout_0.IVS.t18 VDD.t109 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1386 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS2.t539 VOUT_P.t1 VDD.t755 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1387 VDD.t142 VDD.t140 VDD.t142 VDD.t141 pfet_03v3 ad=1.32p pd=6.88u as=0 ps=0 w=3u l=0.28u
X1388 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS1.t14 Folded_Diff_Op_Amp_Layout_0.IBS.t1 VDD.t439 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1389 VOUT_N Folded_Diff_Op_Amp_Layout_0.OUT1.t106 VSS.t71 VSS.t70 nfet_03v3 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.28u
X1390 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t540 VDD.t1287 VDD.t634 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1391 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS.t44 VDD.t21 VDD.t15 pfet_03v3 ad=0.814p pd=3.65u as=0.814p ps=3.65u w=3.13u l=0.56u
X1392 VSS Folded_Diff_Op_Amp_Layout_0.VB4.t102 Folded_Diff_Op_Amp_Layout_0.IPD.t24 VSS.t0 nfet_03v3 ad=0.749p pd=3.4u as=0.749p ps=3.4u w=2.88u l=0.28u
X1393 VSS Folded_Diff_Op_Amp_Layout_0.OUT1.t107 VOUT_N.t2 VSS.t67 nfet_03v3 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.28u
X1394 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VB1.t30 VDD.t939 VDD.t938 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.28u
X1395 VOUT_P Folded_Diff_Op_Amp_Layout_0.OUT2.t107 VSS.t699 VSS.t113 nfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1396 VDD Folded_Diff_Op_Amp_Layout_0.IBIAS3.t80 Folded_Diff_Op_Amp_Layout_0.IVS.t19 VDD.t97 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1397 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.IBIAS.t0 VDD.t39 VDD.t38 pfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.56u
X1398 VOUT_N Folded_Diff_Op_Amp_Layout_0.IBIAS2.t541 VDD.t1288 VDD.t1044 pfet_03v3 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.28u
X1399 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VOUT.t31 Folded_Diff_Op_Amp_Layout_0.VB1.t0 VSS.t277 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
R0 Folded_Diff_Op_Amp_Layout_0.OUT1.t75 Folded_Diff_Op_Amp_Layout_0.OUT1.t59 122.014
R1 Folded_Diff_Op_Amp_Layout_0.OUT1.t77 Folded_Diff_Op_Amp_Layout_0.OUT1.t92 122.014
R2 Folded_Diff_Op_Amp_Layout_0.OUT1.t62 Folded_Diff_Op_Amp_Layout_0.OUT1.t68 122.014
R3 Folded_Diff_Op_Amp_Layout_0.OUT1.t63 Folded_Diff_Op_Amp_Layout_0.OUT1.t51 122.014
R4 Folded_Diff_Op_Amp_Layout_0.OUT1.t101 Folded_Diff_Op_Amp_Layout_0.OUT1.t53 122.014
R5 Folded_Diff_Op_Amp_Layout_0.OUT1.t103 Folded_Diff_Op_Amp_Layout_0.OUT1.t87 122.014
R6 Folded_Diff_Op_Amp_Layout_0.OUT1.t91 Folded_Diff_Op_Amp_Layout_0.OUT1.t67 122.014
R7 Folded_Diff_Op_Amp_Layout_0.OUT1.t82 Folded_Diff_Op_Amp_Layout_0.OUT1.t43 122.014
R8 Folded_Diff_Op_Amp_Layout_0.OUT1.t88 Folded_Diff_Op_Amp_Layout_0.OUT1.t58 122.014
R9 Folded_Diff_Op_Amp_Layout_0.OUT1.t96 Folded_Diff_Op_Amp_Layout_0.OUT1.t80 122.014
R10 Folded_Diff_Op_Amp_Layout_0.OUT1.t56 Folded_Diff_Op_Amp_Layout_0.OUT1.t85 122.014
R11 Folded_Diff_Op_Amp_Layout_0.OUT1.t52 Folded_Diff_Op_Amp_Layout_0.OUT1.t49 122.014
R12 Folded_Diff_Op_Amp_Layout_0.OUT1.n22 Folded_Diff_Op_Amp_Layout_0.OUT1.t90 68.0848
R13 Folded_Diff_Op_Amp_Layout_0.OUT1.n56 Folded_Diff_Op_Amp_Layout_0.OUT1.t95 65.7181
R14 Folded_Diff_Op_Amp_Layout_0.OUT1.n60 Folded_Diff_Op_Amp_Layout_0.OUT1.t71 65.7181
R15 Folded_Diff_Op_Amp_Layout_0.OUT1.n23 Folded_Diff_Op_Amp_Layout_0.OUT1.t36 65.7179
R16 Folded_Diff_Op_Amp_Layout_0.OUT1.n59 Folded_Diff_Op_Amp_Layout_0.OUT1.t64 65.7179
R17 Folded_Diff_Op_Amp_Layout_0.OUT1.n63 Folded_Diff_Op_Amp_Layout_0.OUT1.t81 65.7179
R18 Folded_Diff_Op_Amp_Layout_0.OUT1.n72 Folded_Diff_Op_Amp_Layout_0.OUT1.t102 63.548
R19 Folded_Diff_Op_Amp_Layout_0.OUT1.n65 Folded_Diff_Op_Amp_Layout_0.OUT1.t63 63.548
R20 Folded_Diff_Op_Amp_Layout_0.OUT1.n40 Folded_Diff_Op_Amp_Layout_0.OUT1.t94 63.548
R21 Folded_Diff_Op_Amp_Layout_0.OUT1.n49 Folded_Diff_Op_Amp_Layout_0.OUT1.t100 63.548
R22 Folded_Diff_Op_Amp_Layout_0.OUT1.n25 Folded_Diff_Op_Amp_Layout_0.OUT1.t82 63.548
R23 Folded_Diff_Op_Amp_Layout_0.OUT1.n34 Folded_Diff_Op_Amp_Layout_0.OUT1.t52 63.548
R24 Folded_Diff_Op_Amp_Layout_0.OUT1.n75 Folded_Diff_Op_Amp_Layout_0.OUT1.t55 62.5719
R25 Folded_Diff_Op_Amp_Layout_0.OUT1.n73 Folded_Diff_Op_Amp_Layout_0.OUT1.t42 62.5719
R26 Folded_Diff_Op_Amp_Layout_0.OUT1.n71 Folded_Diff_Op_Amp_Layout_0.OUT1.t83 62.5719
R27 Folded_Diff_Op_Amp_Layout_0.OUT1.n68 Folded_Diff_Op_Amp_Layout_0.OUT1.t72 62.5719
R28 Folded_Diff_Op_Amp_Layout_0.OUT1.n66 Folded_Diff_Op_Amp_Layout_0.OUT1.t62 62.5719
R29 Folded_Diff_Op_Amp_Layout_0.OUT1.n64 Folded_Diff_Op_Amp_Layout_0.OUT1.t79 62.5719
R30 Folded_Diff_Op_Amp_Layout_0.OUT1.n61 Folded_Diff_Op_Amp_Layout_0.OUT1.t70 62.5719
R31 Folded_Diff_Op_Amp_Layout_0.OUT1.n57 Folded_Diff_Op_Amp_Layout_0.OUT1.t66 62.5719
R32 Folded_Diff_Op_Amp_Layout_0.OUT1.n43 Folded_Diff_Op_Amp_Layout_0.OUT1.t41 62.5719
R33 Folded_Diff_Op_Amp_Layout_0.OUT1.n41 Folded_Diff_Op_Amp_Layout_0.OUT1.t40 62.5719
R34 Folded_Diff_Op_Amp_Layout_0.OUT1.n39 Folded_Diff_Op_Amp_Layout_0.OUT1.t93 62.5719
R35 Folded_Diff_Op_Amp_Layout_0.OUT1.n46 Folded_Diff_Op_Amp_Layout_0.OUT1.t37 62.5719
R36 Folded_Diff_Op_Amp_Layout_0.OUT1.n47 Folded_Diff_Op_Amp_Layout_0.OUT1.t50 62.5719
R37 Folded_Diff_Op_Amp_Layout_0.OUT1.n48 Folded_Diff_Op_Amp_Layout_0.OUT1.t76 62.5719
R38 Folded_Diff_Op_Amp_Layout_0.OUT1.n28 Folded_Diff_Op_Amp_Layout_0.OUT1.t45 62.5719
R39 Folded_Diff_Op_Amp_Layout_0.OUT1.n26 Folded_Diff_Op_Amp_Layout_0.OUT1.t91 62.5719
R40 Folded_Diff_Op_Amp_Layout_0.OUT1.n24 Folded_Diff_Op_Amp_Layout_0.OUT1.t74 62.5719
R41 Folded_Diff_Op_Amp_Layout_0.OUT1.n31 Folded_Diff_Op_Amp_Layout_0.OUT1.t44 62.5719
R42 Folded_Diff_Op_Amp_Layout_0.OUT1.n32 Folded_Diff_Op_Amp_Layout_0.OUT1.t56 62.5719
R43 Folded_Diff_Op_Amp_Layout_0.OUT1.n33 Folded_Diff_Op_Amp_Layout_0.OUT1.t69 62.5719
R44 Folded_Diff_Op_Amp_Layout_0.OUT1.n21 Folded_Diff_Op_Amp_Layout_0.OUT1.t97 62.5719
R45 Folded_Diff_Op_Amp_Layout_0.OUT1.n52 Folded_Diff_Op_Amp_Layout_0.OUT1.t106 61.8074
R46 Folded_Diff_Op_Amp_Layout_0.OUT1.n37 Folded_Diff_Op_Amp_Layout_0.OUT1.t88 61.8074
R47 Folded_Diff_Op_Amp_Layout_0.OUT1.n77 Folded_Diff_Op_Amp_Layout_0.OUT1.t107 61.8072
R48 Folded_Diff_Op_Amp_Layout_0.OUT1.n70 Folded_Diff_Op_Amp_Layout_0.OUT1.t75 61.8072
R49 Folded_Diff_Op_Amp_Layout_0.OUT1.n45 Folded_Diff_Op_Amp_Layout_0.OUT1.t104 61.8072
R50 Folded_Diff_Op_Amp_Layout_0.OUT1.n30 Folded_Diff_Op_Amp_Layout_0.OUT1.t101 61.8072
R51 Folded_Diff_Op_Amp_Layout_0.OUT1.n75 Folded_Diff_Op_Amp_Layout_0.OUT1.t61 41.7148
R52 Folded_Diff_Op_Amp_Layout_0.OUT1.n73 Folded_Diff_Op_Amp_Layout_0.OUT1.t60 41.7148
R53 Folded_Diff_Op_Amp_Layout_0.OUT1.n71 Folded_Diff_Op_Amp_Layout_0.OUT1.t89 41.7148
R54 Folded_Diff_Op_Amp_Layout_0.OUT1.n68 Folded_Diff_Op_Amp_Layout_0.OUT1.t39 41.7148
R55 Folded_Diff_Op_Amp_Layout_0.OUT1.n66 Folded_Diff_Op_Amp_Layout_0.OUT1.t77 41.7148
R56 Folded_Diff_Op_Amp_Layout_0.OUT1.n64 Folded_Diff_Op_Amp_Layout_0.OUT1.t73 41.7148
R57 Folded_Diff_Op_Amp_Layout_0.OUT1.n61 Folded_Diff_Op_Amp_Layout_0.OUT1.t84 41.7148
R58 Folded_Diff_Op_Amp_Layout_0.OUT1.n57 Folded_Diff_Op_Amp_Layout_0.OUT1.t98 41.7148
R59 Folded_Diff_Op_Amp_Layout_0.OUT1.n43 Folded_Diff_Op_Amp_Layout_0.OUT1.t57 41.7148
R60 Folded_Diff_Op_Amp_Layout_0.OUT1.n41 Folded_Diff_Op_Amp_Layout_0.OUT1.t54 41.7148
R61 Folded_Diff_Op_Amp_Layout_0.OUT1.n39 Folded_Diff_Op_Amp_Layout_0.OUT1.t86 41.7148
R62 Folded_Diff_Op_Amp_Layout_0.OUT1.n46 Folded_Diff_Op_Amp_Layout_0.OUT1.t105 41.7148
R63 Folded_Diff_Op_Amp_Layout_0.OUT1.n47 Folded_Diff_Op_Amp_Layout_0.OUT1.t47 41.7148
R64 Folded_Diff_Op_Amp_Layout_0.OUT1.n48 Folded_Diff_Op_Amp_Layout_0.OUT1.t48 41.7148
R65 Folded_Diff_Op_Amp_Layout_0.OUT1.n28 Folded_Diff_Op_Amp_Layout_0.OUT1.t65 41.7148
R66 Folded_Diff_Op_Amp_Layout_0.OUT1.n26 Folded_Diff_Op_Amp_Layout_0.OUT1.t103 41.7148
R67 Folded_Diff_Op_Amp_Layout_0.OUT1.n24 Folded_Diff_Op_Amp_Layout_0.OUT1.t99 41.7148
R68 Folded_Diff_Op_Amp_Layout_0.OUT1.n31 Folded_Diff_Op_Amp_Layout_0.OUT1.t78 41.7148
R69 Folded_Diff_Op_Amp_Layout_0.OUT1.n32 Folded_Diff_Op_Amp_Layout_0.OUT1.t96 41.7148
R70 Folded_Diff_Op_Amp_Layout_0.OUT1.n33 Folded_Diff_Op_Amp_Layout_0.OUT1.t46 41.7148
R71 Folded_Diff_Op_Amp_Layout_0.OUT1.n21 Folded_Diff_Op_Amp_Layout_0.OUT1.t38 41.7148
R72 Folded_Diff_Op_Amp_Layout_0.OUT1.n62 Folded_Diff_Op_Amp_Layout_0.OUT1.n61 17.8184
R73 Folded_Diff_Op_Amp_Layout_0.OUT1.n58 Folded_Diff_Op_Amp_Layout_0.OUT1.n57 17.8184
R74 Folded_Diff_Op_Amp_Layout_0.OUT1.n22 Folded_Diff_Op_Amp_Layout_0.OUT1.n21 17.8184
R75 Folded_Diff_Op_Amp_Layout_0.OUT1.n76 Folded_Diff_Op_Amp_Layout_0.OUT1.n75 15.9934
R76 Folded_Diff_Op_Amp_Layout_0.OUT1.n72 Folded_Diff_Op_Amp_Layout_0.OUT1.n71 15.9934
R77 Folded_Diff_Op_Amp_Layout_0.OUT1.n69 Folded_Diff_Op_Amp_Layout_0.OUT1.n68 15.9934
R78 Folded_Diff_Op_Amp_Layout_0.OUT1.n65 Folded_Diff_Op_Amp_Layout_0.OUT1.n64 15.9934
R79 Folded_Diff_Op_Amp_Layout_0.OUT1.n44 Folded_Diff_Op_Amp_Layout_0.OUT1.n43 15.9934
R80 Folded_Diff_Op_Amp_Layout_0.OUT1.n40 Folded_Diff_Op_Amp_Layout_0.OUT1.n39 15.9934
R81 Folded_Diff_Op_Amp_Layout_0.OUT1.n51 Folded_Diff_Op_Amp_Layout_0.OUT1.n46 15.9934
R82 Folded_Diff_Op_Amp_Layout_0.OUT1.n49 Folded_Diff_Op_Amp_Layout_0.OUT1.n48 15.9934
R83 Folded_Diff_Op_Amp_Layout_0.OUT1.n29 Folded_Diff_Op_Amp_Layout_0.OUT1.n28 15.9934
R84 Folded_Diff_Op_Amp_Layout_0.OUT1.n25 Folded_Diff_Op_Amp_Layout_0.OUT1.n24 15.9934
R85 Folded_Diff_Op_Amp_Layout_0.OUT1.n36 Folded_Diff_Op_Amp_Layout_0.OUT1.n31 15.9934
R86 Folded_Diff_Op_Amp_Layout_0.OUT1.n34 Folded_Diff_Op_Amp_Layout_0.OUT1.n33 15.9934
R87 Folded_Diff_Op_Amp_Layout_0.OUT1.n74 Folded_Diff_Op_Amp_Layout_0.OUT1.n73 13.9076
R88 Folded_Diff_Op_Amp_Layout_0.OUT1.n67 Folded_Diff_Op_Amp_Layout_0.OUT1.n66 13.9076
R89 Folded_Diff_Op_Amp_Layout_0.OUT1.n42 Folded_Diff_Op_Amp_Layout_0.OUT1.n41 13.9076
R90 Folded_Diff_Op_Amp_Layout_0.OUT1.n50 Folded_Diff_Op_Amp_Layout_0.OUT1.n47 13.9076
R91 Folded_Diff_Op_Amp_Layout_0.OUT1.n27 Folded_Diff_Op_Amp_Layout_0.OUT1.n26 13.9076
R92 Folded_Diff_Op_Amp_Layout_0.OUT1.n35 Folded_Diff_Op_Amp_Layout_0.OUT1.n32 13.9076
R93 Folded_Diff_Op_Amp_Layout_0.OUT1.n19 Folded_Diff_Op_Amp_Layout_0.OUT1.n79 8.881
R94 Folded_Diff_Op_Amp_Layout_0.OUT1.n78 Folded_Diff_Op_Amp_Layout_0.OUT1.n77 8.79758
R95 Folded_Diff_Op_Amp_Layout_0.OUT1.n60 Folded_Diff_Op_Amp_Layout_0.OUT1.n59 7.75675
R96 Folded_Diff_Op_Amp_Layout_0.OUT1.n111 Folded_Diff_Op_Amp_Layout_0.OUT1.n176 6.80551
R97 Folded_Diff_Op_Amp_Layout_0.OUT1.n185 Folded_Diff_Op_Amp_Layout_0.OUT1.t5 6.49823
R98 Folded_Diff_Op_Amp_Layout_0.OUT1.n185 Folded_Diff_Op_Amp_Layout_0.OUT1.t3 6.4095
R99 Folded_Diff_Op_Amp_Layout_0.OUT1.n54 Folded_Diff_Op_Amp_Layout_0.OUT1.n53 5.6201
R100 Folded_Diff_Op_Amp_Layout_0.OUT1.n95 Folded_Diff_Op_Amp_Layout_0.OUT1.n94 5.52316
R101 Folded_Diff_Op_Amp_Layout_0.OUT1.n82 Folded_Diff_Op_Amp_Layout_0.OUT1.n81 5.49577
R102 Folded_Diff_Op_Amp_Layout_0.OUT1.n78 Folded_Diff_Op_Amp_Layout_0.OUT1.n70 5.42798
R103 Folded_Diff_Op_Amp_Layout_0.OUT1.n98 Folded_Diff_Op_Amp_Layout_0.OUT1.t15 5.40577
R104 Folded_Diff_Op_Amp_Layout_0.OUT1.n101 Folded_Diff_Op_Amp_Layout_0.OUT1.n99 5.40577
R105 Folded_Diff_Op_Amp_Layout_0.OUT1.n102 Folded_Diff_Op_Amp_Layout_0.OUT1.t17 5.40577
R106 Folded_Diff_Op_Amp_Layout_0.OUT1.n151 Folded_Diff_Op_Amp_Layout_0.OUT1.n150 4.67186
R107 Folded_Diff_Op_Amp_Layout_0.OUT1.n97 Folded_Diff_Op_Amp_Layout_0.OUT1.t7 4.64664
R108 Folded_Diff_Op_Amp_Layout_0.OUT1.n159 Folded_Diff_Op_Amp_Layout_0.OUT1.n158 4.54551
R109 Folded_Diff_Op_Amp_Layout_0.OUT1.n79 Folded_Diff_Op_Amp_Layout_0.OUT1.n78 4.5329
R110 Folded_Diff_Op_Amp_Layout_0.OUT1.n55 Folded_Diff_Op_Amp_Layout_0.OUT1.n54 4.5329
R111 Folded_Diff_Op_Amp_Layout_0.OUT1.n95 Folded_Diff_Op_Amp_Layout_0.OUT1.t8 4.39621
R112 Folded_Diff_Op_Amp_Layout_0.OUT1.n96 Folded_Diff_Op_Amp_Layout_0.OUT1.n93 4.39621
R113 Folded_Diff_Op_Amp_Layout_0.OUT1.n82 Folded_Diff_Op_Amp_Layout_0.OUT1.t18 4.36882
R114 Folded_Diff_Op_Amp_Layout_0.OUT1.n83 Folded_Diff_Op_Amp_Layout_0.OUT1.n80 4.36882
R115 Folded_Diff_Op_Amp_Layout_0.OUT1.n140 Folded_Diff_Op_Amp_Layout_0.OUT1.n139 4.08047
R116 Folded_Diff_Op_Amp_Layout_0.OUT1.n139 Folded_Diff_Op_Amp_Layout_0.OUT1.n138 3.8345
R117 Folded_Diff_Op_Amp_Layout_0.OUT1.n98 Folded_Diff_Op_Amp_Layout_0.OUT1.t9 3.71925
R118 Folded_Diff_Op_Amp_Layout_0.OUT1.n101 Folded_Diff_Op_Amp_Layout_0.OUT1.n100 3.71925
R119 Folded_Diff_Op_Amp_Layout_0.OUT1.n102 Folded_Diff_Op_Amp_Layout_0.OUT1.t11 3.71925
R120 Folded_Diff_Op_Amp_Layout_0.OUT1.n53 Folded_Diff_Op_Amp_Layout_0.OUT1.n45 3.17917
R121 Folded_Diff_Op_Amp_Layout_0.OUT1.n38 Folded_Diff_Op_Amp_Layout_0.OUT1.n30 3.17917
R122 Folded_Diff_Op_Amp_Layout_0.OUT1.n55 Folded_Diff_Op_Amp_Layout_0.OUT1.n23 3.17917
R123 Folded_Diff_Op_Amp_Layout_0.OUT1.n53 Folded_Diff_Op_Amp_Layout_0.OUT1.n52 3.17779
R124 Folded_Diff_Op_Amp_Layout_0.OUT1.n38 Folded_Diff_Op_Amp_Layout_0.OUT1.n37 3.17779
R125 Folded_Diff_Op_Amp_Layout_0.OUT1.n79 Folded_Diff_Op_Amp_Layout_0.OUT1.n63 3.17736
R126 Folded_Diff_Op_Amp_Layout_0.OUT1.n56 Folded_Diff_Op_Amp_Layout_0.OUT1.n55 3.17716
R127 Folded_Diff_Op_Amp_Layout_0.OUT1.n108 Folded_Diff_Op_Amp_Layout_0.OUT1.n107 2.61464
R128 Folded_Diff_Op_Amp_Layout_0.OUT1.n183 Folded_Diff_Op_Amp_Layout_0.OUT1.t4 2.4095
R129 Folded_Diff_Op_Amp_Layout_0.OUT1.n188 Folded_Diff_Op_Amp_Layout_0.OUT1.t2 2.4095
R130 Folded_Diff_Op_Amp_Layout_0.OUT1.n54 Folded_Diff_Op_Amp_Layout_0.OUT1.n38 2.2505
R131 Folded_Diff_Op_Amp_Layout_0.OUT1.n88 Folded_Diff_Op_Amp_Layout_0.OUT1.n87 1.84515
R132 Folded_Diff_Op_Amp_Layout_0.OUT1.n18 Folded_Diff_Op_Amp_Layout_0.OUT1.n5 1.84461
R133 Folded_Diff_Op_Amp_Layout_0.OUT1.n84 Folded_Diff_Op_Amp_Layout_0.OUT1.n83 1.80781
R134 Folded_Diff_Op_Amp_Layout_0.OUT1.n147 Folded_Diff_Op_Amp_Layout_0.OUT1.n146 1.63933
R135 Folded_Diff_Op_Amp_Layout_0.OUT1.n138 Folded_Diff_Op_Amp_Layout_0.OUT1.n178 1.6657
R136 Folded_Diff_Op_Amp_Layout_0.OUT1.n20 Folded_Diff_Op_Amp_Layout_0.OUT1.n174 1.51151
R137 Folded_Diff_Op_Amp_Layout_0.OUT1.n140 Folded_Diff_Op_Amp_Layout_0.OUT1.n136 1.48953
R138 Folded_Diff_Op_Amp_Layout_0.OUT1.n141 Folded_Diff_Op_Amp_Layout_0.OUT1.n135 1.48953
R139 Folded_Diff_Op_Amp_Layout_0.OUT1.n186 Folded_Diff_Op_Amp_Layout_0.OUT1.n188 1.43397
R140 Folded_Diff_Op_Amp_Layout_0.OUT1.n125 Folded_Diff_Op_Amp_Layout_0.OUT1.n124 1.40904
R141 Folded_Diff_Op_Amp_Layout_0.OUT1.n131 Folded_Diff_Op_Amp_Layout_0.OUT1.t20 1.40877
R142 Folded_Diff_Op_Amp_Layout_0.OUT1.n14 Folded_Diff_Op_Amp_Layout_0.OUT1.n13 1.40609
R143 Folded_Diff_Op_Amp_Layout_0.OUT1.n2 Folded_Diff_Op_Amp_Layout_0.OUT1.t34 1.40609
R144 Folded_Diff_Op_Amp_Layout_0.OUT1.n103 Folded_Diff_Op_Amp_Layout_0.OUT1.n102 1.27615
R145 Folded_Diff_Op_Amp_Layout_0.OUT1.n59 Folded_Diff_Op_Amp_Layout_0.OUT1.n58 1.21895
R146 Folded_Diff_Op_Amp_Layout_0.OUT1.n62 Folded_Diff_Op_Amp_Layout_0.OUT1.n60 1.21875
R147 Folded_Diff_Op_Amp_Layout_0.OUT1.n143 Folded_Diff_Op_Amp_Layout_0.OUT1.n112 1.20171
R148 Folded_Diff_Op_Amp_Layout_0.OUT1.n132 Folded_Diff_Op_Amp_Layout_0.OUT1.n131 1.19492
R149 Folded_Diff_Op_Amp_Layout_0.OUT1.n126 Folded_Diff_Op_Amp_Layout_0.OUT1.n125 1.19459
R150 Folded_Diff_Op_Amp_Layout_0.OUT1.n15 Folded_Diff_Op_Amp_Layout_0.OUT1.n14 1.19451
R151 Folded_Diff_Op_Amp_Layout_0.OUT1.n3 Folded_Diff_Op_Amp_Layout_0.OUT1.n2 1.19451
R152 Folded_Diff_Op_Amp_Layout_0.OUT1.n164 Folded_Diff_Op_Amp_Layout_0.OUT1.n163 1.18237
R153 Folded_Diff_Op_Amp_Layout_0.OUT1.n119 Folded_Diff_Op_Amp_Layout_0.OUT1.n118 1.17925
R154 Folded_Diff_Op_Amp_Layout_0.OUT1.n10 Folded_Diff_Op_Amp_Layout_0.OUT1.n9 1.17901
R155 Folded_Diff_Op_Amp_Layout_0.OUT1.n165 Folded_Diff_Op_Amp_Layout_0.OUT1.n164 1.17275
R156 Folded_Diff_Op_Amp_Layout_0.OUT1.n172 Folded_Diff_Op_Amp_Layout_0.OUT1.n92 1.1515
R157 Folded_Diff_Op_Amp_Layout_0.OUT1.n148 Folded_Diff_Op_Amp_Layout_0.OUT1.n147 1.14574
R158 Folded_Diff_Op_Amp_Layout_0.OUT1.n89 Folded_Diff_Op_Amp_Layout_0.OUT1.n88 1.14438
R159 Folded_Diff_Op_Amp_Layout_0.OUT1.n104 Folded_Diff_Op_Amp_Layout_0.OUT1.n103 1.12746
R160 Folded_Diff_Op_Amp_Layout_0.OUT1.n110 Folded_Diff_Op_Amp_Layout_0.OUT1.n109 1.1255
R161 Folded_Diff_Op_Amp_Layout_0.OUT1.n86 Folded_Diff_Op_Amp_Layout_0.OUT1.n85 1.1255
R162 Folded_Diff_Op_Amp_Layout_0.OUT1.n153 Folded_Diff_Op_Amp_Layout_0.OUT1.n152 1.1255
R163 Folded_Diff_Op_Amp_Layout_0.OUT1.n161 Folded_Diff_Op_Amp_Layout_0.OUT1.n160 1.1255
R164 Folded_Diff_Op_Amp_Layout_0.OUT1.n175 Folded_Diff_Op_Amp_Layout_0.OUT1.n20 1.1255
R165 Folded_Diff_Op_Amp_Layout_0.OUT1.n171 Folded_Diff_Op_Amp_Layout_0.OUT1.n170 1.1255
R166 Folded_Diff_Op_Amp_Layout_0.OUT1.n178 Folded_Diff_Op_Amp_Layout_0.OUT1.n179 1.12145
R167 Folded_Diff_Op_Amp_Layout_0.OUT1.n63 Folded_Diff_Op_Amp_Layout_0.OUT1.n62 0.905911
R168 Folded_Diff_Op_Amp_Layout_0.OUT1.n23 Folded_Diff_Op_Amp_Layout_0.OUT1.n22 0.90591
R169 Folded_Diff_Op_Amp_Layout_0.OUT1.n58 Folded_Diff_Op_Amp_Layout_0.OUT1.n56 0.905703
R170 Folded_Diff_Op_Amp_Layout_0.OUT1.n97 Folded_Diff_Op_Amp_Layout_0.OUT1.n96 0.877022
R171 Folded_Diff_Op_Amp_Layout_0.OUT1.n144 Folded_Diff_Op_Amp_Layout_0.OUT1.n143 0.873064
R172 Folded_Diff_Op_Amp_Layout_0.OUT1.n118 Folded_Diff_Op_Amp_Layout_0.OUT1.n117 0.827253
R173 Folded_Diff_Op_Amp_Layout_0.OUT1.n9 Folded_Diff_Op_Amp_Layout_0.OUT1.n8 0.824332
R174 Folded_Diff_Op_Amp_Layout_0.OUT1.n167 Folded_Diff_Op_Amp_Layout_0.OUT1.n166 0.743266
R175 Folded_Diff_Op_Amp_Layout_0.OUT1.n0 Folded_Diff_Op_Amp_Layout_0.OUT1.n11 0.727104
R176 Folded_Diff_Op_Amp_Layout_0.OUT1.n122 Folded_Diff_Op_Amp_Layout_0.OUT1.n120 0.727104
R177 Folded_Diff_Op_Amp_Layout_0.OUT1.n104 Folded_Diff_Op_Amp_Layout_0.OUT1.n98 0.650065
R178 Folded_Diff_Op_Amp_Layout_0.OUT1.n103 Folded_Diff_Op_Amp_Layout_0.OUT1.n101 0.650065
R179 Folded_Diff_Op_Amp_Layout_0.OUT1.n112 Folded_Diff_Op_Amp_Layout_0.OUT1.n111 0.632941
R180 Folded_Diff_Op_Amp_Layout_0.OUT1.n91 Folded_Diff_Op_Amp_Layout_0.OUT1.n90 0.632941
R181 Folded_Diff_Op_Amp_Layout_0.OUT1.n128 Folded_Diff_Op_Amp_Layout_0.OUT1.n127 0.631966
R182 Folded_Diff_Op_Amp_Layout_0.OUT1.n96 Folded_Diff_Op_Amp_Layout_0.OUT1.n95 0.626587
R183 Folded_Diff_Op_Amp_Layout_0.OUT1.n105 Folded_Diff_Op_Amp_Layout_0.OUT1.n104 0.626587
R184 Folded_Diff_Op_Amp_Layout_0.OUT1.n83 Folded_Diff_Op_Amp_Layout_0.OUT1.n82 0.626587
R185 Folded_Diff_Op_Amp_Layout_0.OUT1.n74 Folded_Diff_Op_Amp_Layout_0.OUT1.n72 0.626587
R186 Folded_Diff_Op_Amp_Layout_0.OUT1.n76 Folded_Diff_Op_Amp_Layout_0.OUT1.n74 0.626587
R187 Folded_Diff_Op_Amp_Layout_0.OUT1.n67 Folded_Diff_Op_Amp_Layout_0.OUT1.n65 0.626587
R188 Folded_Diff_Op_Amp_Layout_0.OUT1.n69 Folded_Diff_Op_Amp_Layout_0.OUT1.n67 0.626587
R189 Folded_Diff_Op_Amp_Layout_0.OUT1.n42 Folded_Diff_Op_Amp_Layout_0.OUT1.n40 0.626587
R190 Folded_Diff_Op_Amp_Layout_0.OUT1.n44 Folded_Diff_Op_Amp_Layout_0.OUT1.n42 0.626587
R191 Folded_Diff_Op_Amp_Layout_0.OUT1.n51 Folded_Diff_Op_Amp_Layout_0.OUT1.n50 0.626587
R192 Folded_Diff_Op_Amp_Layout_0.OUT1.n50 Folded_Diff_Op_Amp_Layout_0.OUT1.n49 0.626587
R193 Folded_Diff_Op_Amp_Layout_0.OUT1.n27 Folded_Diff_Op_Amp_Layout_0.OUT1.n25 0.626587
R194 Folded_Diff_Op_Amp_Layout_0.OUT1.n29 Folded_Diff_Op_Amp_Layout_0.OUT1.n27 0.626587
R195 Folded_Diff_Op_Amp_Layout_0.OUT1.n36 Folded_Diff_Op_Amp_Layout_0.OUT1.n35 0.626587
R196 Folded_Diff_Op_Amp_Layout_0.OUT1.n35 Folded_Diff_Op_Amp_Layout_0.OUT1.n34 0.626587
R197 Folded_Diff_Op_Amp_Layout_0.OUT1.n114 Folded_Diff_Op_Amp_Layout_0.OUT1.n133 0.616779
R198 Folded_Diff_Op_Amp_Layout_0.OUT1.n156 Folded_Diff_Op_Amp_Layout_0.OUT1.n154 0.616779
R199 Folded_Diff_Op_Amp_Layout_0.OUT1.n17 Folded_Diff_Op_Amp_Layout_0.OUT1.n16 0.631966
R200 Folded_Diff_Op_Amp_Layout_0.OUT1.n5 Folded_Diff_Op_Amp_Layout_0.OUT1.n4 0.616779
R201 Folded_Diff_Op_Amp_Layout_0.OUT1.n117 Folded_Diff_Op_Amp_Layout_0.OUT1.t35 0.58197
R202 Folded_Diff_Op_Amp_Layout_0.OUT1.n117 Folded_Diff_Op_Amp_Layout_0.OUT1.n116 0.58197
R203 Folded_Diff_Op_Amp_Layout_0.OUT1.n163 Folded_Diff_Op_Amp_Layout_0.OUT1.t25 0.58197
R204 Folded_Diff_Op_Amp_Layout_0.OUT1.n163 Folded_Diff_Op_Amp_Layout_0.OUT1.n162 0.58197
R205 Folded_Diff_Op_Amp_Layout_0.OUT1.n158 Folded_Diff_Op_Amp_Layout_0.OUT1.t21 0.58197
R206 Folded_Diff_Op_Amp_Layout_0.OUT1.n158 Folded_Diff_Op_Amp_Layout_0.OUT1.n157 0.58197
R207 Folded_Diff_Op_Amp_Layout_0.OUT1.n146 Folded_Diff_Op_Amp_Layout_0.OUT1.t29 0.58197
R208 Folded_Diff_Op_Amp_Layout_0.OUT1.n146 Folded_Diff_Op_Amp_Layout_0.OUT1.n145 0.58197
R209 Folded_Diff_Op_Amp_Layout_0.OUT1.n150 Folded_Diff_Op_Amp_Layout_0.OUT1.t23 0.58197
R210 Folded_Diff_Op_Amp_Layout_0.OUT1.n150 Folded_Diff_Op_Amp_Layout_0.OUT1.n149 0.58197
R211 Folded_Diff_Op_Amp_Layout_0.OUT1.n8 Folded_Diff_Op_Amp_Layout_0.OUT1.t28 0.58197
R212 Folded_Diff_Op_Amp_Layout_0.OUT1.n8 Folded_Diff_Op_Amp_Layout_0.OUT1.n7 0.58197
R213 Folded_Diff_Op_Amp_Layout_0.OUT1.n107 Folded_Diff_Op_Amp_Layout_0.OUT1.n106 0.56925
R214 Folded_Diff_Op_Amp_Layout_0.OUT1.n87 Folded_Diff_Op_Amp_Layout_0.OUT1.t12 0.56925
R215 Folded_Diff_Op_Amp_Layout_0.OUT1.n169 Folded_Diff_Op_Amp_Layout_0.OUT1.n168 0.5585
R216 Folded_Diff_Op_Amp_Layout_0.OUT1.n92 Folded_Diff_Op_Amp_Layout_0.OUT1.n91 0.54725
R217 Folded_Diff_Op_Amp_Layout_0.OUT1.n155 Folded_Diff_Op_Amp_Layout_0.OUT1.n167 0.474125
R218 Folded_Diff_Op_Amp_Layout_0.OUT1.n121 Folded_Diff_Op_Amp_Layout_0.OUT1.n128 0.474125
R219 Folded_Diff_Op_Amp_Layout_0.OUT1.n113 Folded_Diff_Op_Amp_Layout_0.OUT1.n129 0.474125
R220 Folded_Diff_Op_Amp_Layout_0.OUT1.n143 Folded_Diff_Op_Amp_Layout_0.OUT1.n142 0.459221
R221 Folded_Diff_Op_Amp_Layout_0.OUT1.n160 Folded_Diff_Op_Amp_Layout_0.OUT1.n159 0.366599
R222 Folded_Diff_Op_Amp_Layout_0.OUT1.n135 Folded_Diff_Op_Amp_Layout_0.OUT1.n134 0.3255
R223 Folded_Diff_Op_Amp_Layout_0.OUT1.n77 Folded_Diff_Op_Amp_Layout_0.OUT1.n76 0.279823
R224 Folded_Diff_Op_Amp_Layout_0.OUT1.n70 Folded_Diff_Op_Amp_Layout_0.OUT1.n69 0.279823
R225 Folded_Diff_Op_Amp_Layout_0.OUT1.n45 Folded_Diff_Op_Amp_Layout_0.OUT1.n44 0.279823
R226 Folded_Diff_Op_Amp_Layout_0.OUT1.n30 Folded_Diff_Op_Amp_Layout_0.OUT1.n29 0.279823
R227 Folded_Diff_Op_Amp_Layout_0.OUT1.n52 Folded_Diff_Op_Amp_Layout_0.OUT1.n51 0.279615
R228 Folded_Diff_Op_Amp_Layout_0.OUT1.n37 Folded_Diff_Op_Amp_Layout_0.OUT1.n36 0.279615
R229 Folded_Diff_Op_Amp_Layout_0.OUT1.n152 Folded_Diff_Op_Amp_Layout_0.OUT1.n151 0.223214
R230 Folded_Diff_Op_Amp_Layout_0.OUT1.n173 Folded_Diff_Op_Amp_Layout_0.OUT1.n172 0.221875
R231 Folded_Diff_Op_Amp_Layout_0.OUT1.n105 Folded_Diff_Op_Amp_Layout_0.OUT1.n97 0.1805
R232 Folded_Diff_Op_Amp_Layout_0.OUT1.n85 Folded_Diff_Op_Amp_Layout_0.OUT1.n84 0.171378
R233 Folded_Diff_Op_Amp_Layout_0.OUT1.n108 Folded_Diff_Op_Amp_Layout_0.OUT1.n105 0.163273
R234 Folded_Diff_Op_Amp_Layout_0.OUT1.n138 Folded_Diff_Op_Amp_Layout_0.OUT1.n137 0.119218
R235 Folded_Diff_Op_Amp_Layout_0.OUT1.n120 Folded_Diff_Op_Amp_Layout_0.OUT1.n115 0.0823987
R236 Folded_Diff_Op_Amp_Layout_0.OUT1.n166 Folded_Diff_Op_Amp_Layout_0.OUT1.n161 0.0823987
R237 Folded_Diff_Op_Amp_Layout_0.OUT1.n11 Folded_Diff_Op_Amp_Layout_0.OUT1.n6 0.0823987
R238 Folded_Diff_Op_Amp_Layout_0.OUT1.n90 Folded_Diff_Op_Amp_Layout_0.OUT1.n86 0.0712285
R239 Folded_Diff_Op_Amp_Layout_0.OUT1.n154 Folded_Diff_Op_Amp_Layout_0.OUT1.n148 0.0712285
R240 Folded_Diff_Op_Amp_Layout_0.OUT1.n4 Folded_Diff_Op_Amp_Layout_0.OUT1.n1 0.0712285
R241 Folded_Diff_Op_Amp_Layout_0.OUT1.n16 Folded_Diff_Op_Amp_Layout_0.OUT1.n12 0.0712285
R242 Folded_Diff_Op_Amp_Layout_0.OUT1.n127 Folded_Diff_Op_Amp_Layout_0.OUT1.n123 0.0712285
R243 Folded_Diff_Op_Amp_Layout_0.OUT1.n133 Folded_Diff_Op_Amp_Layout_0.OUT1.n130 0.0712285
R244 Folded_Diff_Op_Amp_Layout_0.OUT1.n182 Folded_Diff_Op_Amp_Layout_0.OUT1.n185 0.0607113
R245 Folded_Diff_Op_Amp_Layout_0.OUT1.n111 Folded_Diff_Op_Amp_Layout_0.OUT1.n110 0.0534597
R246 Folded_Diff_Op_Amp_Layout_0.OUT1.n90 Folded_Diff_Op_Amp_Layout_0.OUT1.n89 0.0534597
R247 Folded_Diff_Op_Amp_Layout_0.OUT1.n154 Folded_Diff_Op_Amp_Layout_0.OUT1.n153 0.0534597
R248 Folded_Diff_Op_Amp_Layout_0.OUT1.n16 Folded_Diff_Op_Amp_Layout_0.OUT1.n15 0.0534597
R249 Folded_Diff_Op_Amp_Layout_0.OUT1.n4 Folded_Diff_Op_Amp_Layout_0.OUT1.n3 0.0534597
R250 Folded_Diff_Op_Amp_Layout_0.OUT1.n127 Folded_Diff_Op_Amp_Layout_0.OUT1.n126 0.0534597
R251 Folded_Diff_Op_Amp_Layout_0.OUT1.n133 Folded_Diff_Op_Amp_Layout_0.OUT1.n132 0.0534597
R252 Folded_Diff_Op_Amp_Layout_0.OUT1.n172 Folded_Diff_Op_Amp_Layout_0.OUT1.n171 0.0525
R253 Folded_Diff_Op_Amp_Layout_0.OUT1.n171 Folded_Diff_Op_Amp_Layout_0.OUT1.n144 0.0525
R254 Folded_Diff_Op_Amp_Layout_0.OUT1.n20 Folded_Diff_Op_Amp_Layout_0.OUT1.n18 0.0494128
R255 Folded_Diff_Op_Amp_Layout_0.OUT1.n166 Folded_Diff_Op_Amp_Layout_0.OUT1.n165 0.0415773
R256 Folded_Diff_Op_Amp_Layout_0.OUT1.n11 Folded_Diff_Op_Amp_Layout_0.OUT1.n10 0.0415773
R257 Folded_Diff_Op_Amp_Layout_0.OUT1.n120 Folded_Diff_Op_Amp_Layout_0.OUT1.n119 0.0415773
R258 Folded_Diff_Op_Amp_Layout_0.OUT1.n141 Folded_Diff_Op_Amp_Layout_0.OUT1.n140 0.0354016
R259 Folded_Diff_Op_Amp_Layout_0.OUT1.n175 Folded_Diff_Op_Amp_Layout_0.OUT1 0.0296408
R260 Folded_Diff_Op_Amp_Layout_0.OUT1.n170 Folded_Diff_Op_Amp_Layout_0.OUT1.n169 0.0265
R261 Folded_Diff_Op_Amp_Layout_0.OUT1.n184 Folded_Diff_Op_Amp_Layout_0.OUT1.n180 0.0214155
R262 Folded_Diff_Op_Amp_Layout_0.OUT1.n180 Folded_Diff_Op_Amp_Layout_0.OUT1.n187 0.0210986
R263 Folded_Diff_Op_Amp_Layout_0.OUT1.n109 Folded_Diff_Op_Amp_Layout_0.OUT1.n108 0.0204805
R264 Folded_Diff_Op_Amp_Layout_0.OUT1.n186 Folded_Diff_Op_Amp_Layout_0.OUT1.n182 0.0277051
R265 Folded_Diff_Op_Amp_Layout_0.OUT1.n142 Folded_Diff_Op_Amp_Layout_0.OUT1.n141 0.0182008
R266 Folded_Diff_Op_Amp_Layout_0.OUT1.n179 Folded_Diff_Op_Amp_Layout_0.OUT1.n183 1.4506
R267 Folded_Diff_Op_Amp_Layout_0.OUT1.n20 Folded_Diff_Op_Amp_Layout_0.OUT1.n19 0.0199708
R268 Folded_Diff_Op_Amp_Layout_0.OUT1.n181 Folded_Diff_Op_Amp_Layout_0.OUT1.n186 0.0171032
R269 Folded_Diff_Op_Amp_Layout_0.OUT1.n129 Folded_Diff_Op_Amp_Layout_0.OUT1.n122 0.016662
R270 Folded_Diff_Op_Amp_Layout_0.OUT1.n114 Folded_Diff_Op_Amp_Layout_0.OUT1.n113 0.016662
R271 Folded_Diff_Op_Amp_Layout_0.OUT1.n156 Folded_Diff_Op_Amp_Layout_0.OUT1.n155 0.016662
R272 Folded_Diff_Op_Amp_Layout_0.OUT1.n122 Folded_Diff_Op_Amp_Layout_0.OUT1.n121 0.0166619
R273 Folded_Diff_Op_Amp_Layout_0.OUT1.n168 Folded_Diff_Op_Amp_Layout_0.OUT1.n156 0.0156875
R274 Folded_Diff_Op_Amp_Layout_0.OUT1.n134 Folded_Diff_Op_Amp_Layout_0.OUT1.n114 0.0156875
R275 Folded_Diff_Op_Amp_Layout_0.OUT1.n18 Folded_Diff_Op_Amp_Layout_0.OUT1.n173 0.014
R276 Folded_Diff_Op_Amp_Layout_0.OUT1.n187 Folded_Diff_Op_Amp_Layout_0.OUT1.n181 0.0128592
R277 Folded_Diff_Op_Amp_Layout_0.OUT1.n179 Folded_Diff_Op_Amp_Layout_0.OUT1.n184 0.0125423
R278 Folded_Diff_Op_Amp_Layout_0.OUT1.n178 Folded_Diff_Op_Amp_Layout_0.OUT1.n177 0.010845
R279 Folded_Diff_Op_Amp_Layout_0.OUT1.n0 Folded_Diff_Op_Amp_Layout_0.OUT1.n5 0.506449
R280 Folded_Diff_Op_Amp_Layout_0.OUT1.n0 Folded_Diff_Op_Amp_Layout_0.OUT1.n17 0.490287
R281 VOUT_N.n176 VOUT_N.t75 7.30465
R282 VOUT_N.n2026 VOUT_N.n2025 7.04823
R283 VOUT_N VOUT_N.t74 4.20265
R284 VOUT_N.n170 VOUT_N.n169 4.07744
R285 VOUT_N.n179 VOUT_N.n178 2.40958
R286 VOUT_N.n2024 VOUT_N.t273 2.38651
R287 VOUT_N.n2024 VOUT_N.t272 2.2505
R288 VOUT_N.n2025 VOUT_N.n2024 2.20377
R289 VOUT_N.n1909 VOUT_N.n1908 1.84464
R290 VOUT_N.n1896 VOUT_N.n1895 1.84464
R291 VOUT_N.n169 VOUT_N.n168 1.52554
R292 VOUT_N.n2153 VOUT_N.n2152 1.50509
R293 VOUT_N.n2159 VOUT_N.n2158 1.50275
R294 VOUT_N.n145 VOUT_N.n144 1.50001
R295 VOUT_N.n131 VOUT_N.n126 1.50001
R296 VOUT_N.n131 VOUT_N.n130 1.50001
R297 VOUT_N.n167 VOUT_N.n166 1.50001
R298 VOUT_N.n66 VOUT_N.n65 1.50001
R299 VOUT_N.n92 VOUT_N.n91 1.50001
R300 VOUT_N.n104 VOUT_N.n103 1.4999
R301 VOUT_N.n2050 VOUT_N.n2049 1.49371
R302 VOUT_N.n2173 VOUT_N.n2172 1.49371
R303 VOUT_N.n1631 VOUT_N.n1349 1.49371
R304 VOUT_N.n1630 VOUT_N.n1351 1.49371
R305 VOUT_N.n2204 VOUT_N.n2203 1.49371
R306 VOUT_N.n1672 VOUT_N.n1671 1.49371
R307 VOUT_N.n1300 VOUT_N.n1299 1.49371
R308 VOUT_N.n942 VOUT_N.n941 1.49371
R309 VOUT_N.n2154 VOUT_N.n2149 1.48107
R310 VOUT_N.n1939 VOUT_N.n1938 1.47979
R311 VOUT_N.n2146 VOUT_N.n2145 1.47979
R312 VOUT_N.n1708 VOUT_N.n1707 1.47979
R313 VOUT_N.n551 VOUT_N.t2 1.46987
R314 VOUT_N.n541 VOUT_N.n540 1.46987
R315 VOUT_N.n532 VOUT_N.t6 1.46987
R316 VOUT_N.n522 VOUT_N.n521 1.46987
R317 VOUT_N.n517 VOUT_N.t4 1.46987
R318 VOUT_N.n507 VOUT_N.n506 1.46987
R319 VOUT_N.n1823 VOUT_N.n1822 1.46987
R320 VOUT_N.n1833 VOUT_N.t37 1.46987
R321 VOUT_N.n1838 VOUT_N.n1837 1.46987
R322 VOUT_N.n1848 VOUT_N.t23 1.46987
R323 VOUT_N.n2011 VOUT_N.n2010 1.46987
R324 VOUT_N.n2021 VOUT_N.t13 1.46959
R325 VOUT_N.n326 VOUT_N.n325 1.43193
R326 VOUT_N.n1454 VOUT_N.n1453 1.43193
R327 VOUT_N.n1437 VOUT_N.t171 1.43193
R328 VOUT_N.n1433 VOUT_N.n1432 1.43193
R329 VOUT_N.n1416 VOUT_N.t87 1.43193
R330 VOUT_N.n1412 VOUT_N.n1411 1.43193
R331 VOUT_N.n1395 VOUT_N.t241 1.43193
R332 VOUT_N.n1391 VOUT_N.n1390 1.43193
R333 VOUT_N.n1374 VOUT_N.t135 1.43193
R334 VOUT_N.n1370 VOUT_N.n1369 1.43193
R335 VOUT_N.n1306 VOUT_N.t90 1.43193
R336 VOUT_N.n1323 VOUT_N.n1322 1.43193
R337 VOUT_N.n1327 VOUT_N.t151 1.43193
R338 VOUT_N.n1344 VOUT_N.n1343 1.43193
R339 VOUT_N.n1353 VOUT_N.t195 1.43193
R340 VOUT_N.n309 VOUT_N.t79 1.43193
R341 VOUT_N.n305 VOUT_N.n304 1.43193
R342 VOUT_N.n288 VOUT_N.t243 1.43193
R343 VOUT_N.n284 VOUT_N.n283 1.43193
R344 VOUT_N.n267 VOUT_N.t119 1.43193
R345 VOUT_N.n263 VOUT_N.n262 1.43193
R346 VOUT_N.n246 VOUT_N.t168 1.43193
R347 VOUT_N.n242 VOUT_N.n241 1.43193
R348 VOUT_N.n225 VOUT_N.t212 1.43193
R349 VOUT_N.n221 VOUT_N.n220 1.43193
R350 VOUT_N.n204 VOUT_N.t104 1.43193
R351 VOUT_N.n200 VOUT_N.n199 1.43193
R352 VOUT_N.n183 VOUT_N.t96 1.43193
R353 VOUT_N.n1903 VOUT_N.n1902 1.28777
R354 VOUT_N.n2068 VOUT_N.n2067 1.28777
R355 VOUT_N.n2061 VOUT_N.n2060 1.28777
R356 VOUT_N.n2078 VOUT_N.n2077 1.28777
R357 VOUT_N.n1778 VOUT_N.n1777 1.28777
R358 VOUT_N.n1786 VOUT_N.n1785 1.28777
R359 VOUT_N.n1770 VOUT_N.n1769 1.28777
R360 VOUT_N.n2181 VOUT_N.n2178 1.1949
R361 VOUT_N.n2191 VOUT_N.n2190 1.1949
R362 VOUT_N.n1981 VOUT_N.n1980 1.1949
R363 VOUT_N.n1988 VOUT_N.n1985 1.1949
R364 VOUT_N.n11 VOUT_N.n10 1.1949
R365 VOUT_N.n18 VOUT_N.n15 1.1949
R366 VOUT_N.n1740 VOUT_N.n1739 1.1949
R367 VOUT_N.n1747 VOUT_N.n1744 1.1949
R368 VOUT_N.n783 VOUT_N.n782 1.1948
R369 VOUT_N.n771 VOUT_N.n770 1.1948
R370 VOUT_N.n759 VOUT_N.n758 1.1948
R371 VOUT_N.n747 VOUT_N.n746 1.1948
R372 VOUT_N.n735 VOUT_N.n734 1.1948
R373 VOUT_N.n723 VOUT_N.n722 1.1948
R374 VOUT_N.n627 VOUT_N.n626 1.1948
R375 VOUT_N.n639 VOUT_N.n638 1.1948
R376 VOUT_N.n651 VOUT_N.n650 1.1948
R377 VOUT_N.n663 VOUT_N.n662 1.1948
R378 VOUT_N.n675 VOUT_N.n674 1.1948
R379 VOUT_N.n687 VOUT_N.n686 1.1948
R380 VOUT_N.n699 VOUT_N.n698 1.1948
R381 VOUT_N.n711 VOUT_N.n710 1.1948
R382 VOUT_N.n1118 VOUT_N.n1117 1.1948
R383 VOUT_N.n1106 VOUT_N.n1105 1.1948
R384 VOUT_N.n1094 VOUT_N.n1093 1.1948
R385 VOUT_N.n1082 VOUT_N.n1081 1.1948
R386 VOUT_N.n1070 VOUT_N.n1069 1.1948
R387 VOUT_N.n1058 VOUT_N.n1057 1.1948
R388 VOUT_N.n1046 VOUT_N.n1045 1.1948
R389 VOUT_N.n1034 VOUT_N.n1033 1.1948
R390 VOUT_N.n1022 VOUT_N.n1021 1.1948
R391 VOUT_N.n1010 VOUT_N.n1009 1.1948
R392 VOUT_N.n956 VOUT_N.n955 1.1948
R393 VOUT_N.n968 VOUT_N.n967 1.1948
R394 VOUT_N.n980 VOUT_N.n979 1.1948
R395 VOUT_N.n992 VOUT_N.n991 1.1948
R396 VOUT_N.n1438 VOUT_N.n1437 1.19473
R397 VOUT_N.n1417 VOUT_N.n1416 1.19473
R398 VOUT_N.n1396 VOUT_N.n1395 1.19473
R399 VOUT_N.n1375 VOUT_N.n1374 1.19473
R400 VOUT_N.n1307 VOUT_N.n1306 1.19473
R401 VOUT_N.n1328 VOUT_N.n1327 1.19473
R402 VOUT_N.n1354 VOUT_N.n1353 1.19473
R403 VOUT_N.n310 VOUT_N.n309 1.19473
R404 VOUT_N.n289 VOUT_N.n288 1.19473
R405 VOUT_N.n268 VOUT_N.n267 1.19473
R406 VOUT_N.n247 VOUT_N.n246 1.19473
R407 VOUT_N.n226 VOUT_N.n225 1.19473
R408 VOUT_N.n205 VOUT_N.n204 1.19473
R409 VOUT_N.n184 VOUT_N.n183 1.19473
R410 VOUT_N.n2109 VOUT_N.n2108 1.19461
R411 VOUT_N.n1866 VOUT_N.n1865 1.19461
R412 VOUT_N.n552 VOUT_N.n551 1.19458
R413 VOUT_N.n542 VOUT_N.n541 1.19458
R414 VOUT_N.n518 VOUT_N.n517 1.19458
R415 VOUT_N.n508 VOUT_N.n507 1.19458
R416 VOUT_N.n1839 VOUT_N.n1838 1.19458
R417 VOUT_N.n1849 VOUT_N.n1848 1.19458
R418 VOUT_N.n322 VOUT_N.n321 1.19445
R419 VOUT_N.n1450 VOUT_N.n1449 1.19445
R420 VOUT_N.n1429 VOUT_N.n1428 1.19445
R421 VOUT_N.n1408 VOUT_N.n1407 1.19445
R422 VOUT_N.n1387 VOUT_N.n1386 1.19445
R423 VOUT_N.n1366 VOUT_N.n1365 1.19445
R424 VOUT_N.n1319 VOUT_N.n1318 1.19445
R425 VOUT_N.n1340 VOUT_N.n1339 1.19445
R426 VOUT_N.n301 VOUT_N.n300 1.19445
R427 VOUT_N.n280 VOUT_N.n279 1.19445
R428 VOUT_N.n259 VOUT_N.n258 1.19445
R429 VOUT_N.n238 VOUT_N.n237 1.19445
R430 VOUT_N.n217 VOUT_N.n216 1.19445
R431 VOUT_N.n196 VOUT_N.n195 1.19445
R432 VOUT_N.n529 VOUT_N.n528 1.19426
R433 VOUT_N.n1830 VOUT_N.n1829 1.19426
R434 VOUT_N.n2018 VOUT_N.n2017 1.19426
R435 VOUT_N.n548 VOUT_N.n547 1.17959
R436 VOUT_N.n514 VOUT_N.n513 1.17959
R437 VOUT_N.n1845 VOUT_N.n1844 1.17959
R438 VOUT_N.n533 VOUT_N.n532 1.1793
R439 VOUT_N.n523 VOUT_N.n522 1.1793
R440 VOUT_N.n1824 VOUT_N.n1823 1.1793
R441 VOUT_N.n1834 VOUT_N.n1833 1.1793
R442 VOUT_N.n2012 VOUT_N.n2011 1.1793
R443 VOUT_N.n316 VOUT_N.n315 1.1791
R444 VOUT_N.n1444 VOUT_N.n1443 1.1791
R445 VOUT_N.n1423 VOUT_N.n1422 1.1791
R446 VOUT_N.n1402 VOUT_N.n1401 1.1791
R447 VOUT_N.n1381 VOUT_N.n1380 1.1791
R448 VOUT_N.n1360 VOUT_N.n1359 1.1791
R449 VOUT_N.n1313 VOUT_N.n1312 1.1791
R450 VOUT_N.n1334 VOUT_N.n1333 1.1791
R451 VOUT_N.n295 VOUT_N.n294 1.1791
R452 VOUT_N.n274 VOUT_N.n273 1.1791
R453 VOUT_N.n253 VOUT_N.n252 1.1791
R454 VOUT_N.n232 VOUT_N.n231 1.1791
R455 VOUT_N.n211 VOUT_N.n210 1.1791
R456 VOUT_N.n190 VOUT_N.n189 1.1791
R457 VOUT_N.n1872 VOUT_N.n1871 1.17896
R458 VOUT_N.n2103 VOUT_N.n2102 1.17896
R459 VOUT_N.n2022 VOUT_N.n2021 1.17896
R460 VOUT_N.n327 VOUT_N.n326 1.17884
R461 VOUT_N.n1455 VOUT_N.n1454 1.17884
R462 VOUT_N.n1434 VOUT_N.n1433 1.17884
R463 VOUT_N.n1413 VOUT_N.n1412 1.17884
R464 VOUT_N.n1392 VOUT_N.n1391 1.17884
R465 VOUT_N.n1371 VOUT_N.n1370 1.17884
R466 VOUT_N.n1324 VOUT_N.n1323 1.17884
R467 VOUT_N.n1345 VOUT_N.n1344 1.17884
R468 VOUT_N.n306 VOUT_N.n305 1.17884
R469 VOUT_N.n285 VOUT_N.n284 1.17884
R470 VOUT_N.n264 VOUT_N.n263 1.17884
R471 VOUT_N.n243 VOUT_N.n242 1.17884
R472 VOUT_N.n222 VOUT_N.n221 1.17884
R473 VOUT_N.n201 VOUT_N.n200 1.17884
R474 VOUT_N.n777 VOUT_N.n776 1.17849
R475 VOUT_N.n765 VOUT_N.n764 1.17849
R476 VOUT_N.n753 VOUT_N.n752 1.17849
R477 VOUT_N.n741 VOUT_N.n740 1.17849
R478 VOUT_N.n729 VOUT_N.n728 1.17849
R479 VOUT_N.n621 VOUT_N.n620 1.17849
R480 VOUT_N.n633 VOUT_N.n632 1.17849
R481 VOUT_N.n645 VOUT_N.n644 1.17849
R482 VOUT_N.n657 VOUT_N.n656 1.17849
R483 VOUT_N.n669 VOUT_N.n668 1.17849
R484 VOUT_N.n681 VOUT_N.n680 1.17849
R485 VOUT_N.n693 VOUT_N.n692 1.17849
R486 VOUT_N.n705 VOUT_N.n704 1.17849
R487 VOUT_N.n717 VOUT_N.n716 1.17849
R488 VOUT_N.n1112 VOUT_N.n1111 1.17849
R489 VOUT_N.n1100 VOUT_N.n1099 1.17849
R490 VOUT_N.n1088 VOUT_N.n1087 1.17849
R491 VOUT_N.n1076 VOUT_N.n1075 1.17849
R492 VOUT_N.n1064 VOUT_N.n1063 1.17849
R493 VOUT_N.n1052 VOUT_N.n1051 1.17849
R494 VOUT_N.n1040 VOUT_N.n1039 1.17849
R495 VOUT_N.n1028 VOUT_N.n1027 1.17849
R496 VOUT_N.n1016 VOUT_N.n1015 1.17849
R497 VOUT_N.n950 VOUT_N.n949 1.17849
R498 VOUT_N.n962 VOUT_N.n961 1.17849
R499 VOUT_N.n974 VOUT_N.n973 1.17849
R500 VOUT_N.n986 VOUT_N.n985 1.17849
R501 VOUT_N.n1004 VOUT_N.n1003 1.17849
R502 VOUT_N.n2062 VOUT_N.n2061 1.1742
R503 VOUT_N.n2079 VOUT_N.n2078 1.1742
R504 VOUT_N.n2158 VOUT_N.n2157 1.16696
R505 VOUT_N.n1944 VOUT_N.n1943 1.16696
R506 VOUT_N.n1966 VOUT_N.n1965 1.16696
R507 VOUT_N.n2139 VOUT_N.n2138 1.16696
R508 VOUT_N.n1699 VOUT_N.n1698 1.16696
R509 VOUT_N.n1720 VOUT_N.n1719 1.16696
R510 VOUT_N.n1897 VOUT_N.n1896 1.14437
R511 VOUT_N.n1940 VOUT_N.n1939 1.14073
R512 VOUT_N.n2147 VOUT_N.n2146 1.14073
R513 VOUT_N.n1709 VOUT_N.n1708 1.14073
R514 VOUT_N.n1686 VOUT_N.n1685 1.1353
R515 VOUT_N.n1734 VOUT_N.n1733 1.12925
R516 VOUT_N.n1764 VOUT_N.n1763 1.12925
R517 VOUT_N.n2182 VOUT_N.n2181 1.12829
R518 VOUT_N.n1914 VOUT_N.n1913 1.12829
R519 VOUT_N.n1700 VOUT_N.n1699 1.12829
R520 VOUT_N.n1989 VOUT_N.n1988 1.12795
R521 VOUT_N.n19 VOUT_N.n18 1.12795
R522 VOUT_N.n1789 VOUT_N.n1788 1.12795
R523 VOUT_N.n1748 VOUT_N.n1747 1.12795
R524 VOUT_N.n1710 VOUT_N.n1709 1.12695
R525 VOUT_N.n1947 VOUT_N.n1946 1.1255
R526 VOUT_N.n1913 VOUT_N.n1910 1.1255
R527 VOUT_N.n1962 VOUT_N.n1961 1.1255
R528 VOUT_N.n1893 VOUT_N.n1892 1.1255
R529 VOUT_N.n1905 VOUT_N.n1904 1.1255
R530 VOUT_N.n2070 VOUT_N.n2069 1.1255
R531 VOUT_N.n2059 VOUT_N.n2058 1.1255
R532 VOUT_N.n2075 VOUT_N.n2074 1.1255
R533 VOUT_N.n2152 VOUT_N.n2151 1.1255
R534 VOUT_N.n2143 VOUT_N.n2142 1.1255
R535 VOUT_N.n2136 VOUT_N.n2135 1.1255
R536 VOUT_N.n1936 VOUT_N.n1935 1.1255
R537 VOUT_N.n1780 VOUT_N.n1779 1.1255
R538 VOUT_N.n1691 VOUT_N.n1690 1.1255
R539 VOUT_N.n1788 VOUT_N.n1787 1.1255
R540 VOUT_N.n1716 VOUT_N.n1715 1.1255
R541 VOUT_N.n1772 VOUT_N.n1771 1.1255
R542 VOUT_N.n2025 VOUT_N 1.1216
R543 VOUT_N.n2000 VOUT_N.n1999 1.11801
R544 VOUT_N.n1928 VOUT_N.n1927 1.11801
R545 VOUT_N.n1884 VOUT_N.n1883 1.11801
R546 VOUT_N.n2129 VOUT_N.n2095 1.11801
R547 VOUT_N.n2199 VOUT_N.n2056 1.11801
R548 VOUT_N.n1244 VOUT_N.n999 1.11801
R549 VOUT_N.n1540 VOUT_N.n1539 1.11801
R550 VOUT_N.n1620 VOUT_N.n1619 1.11801
R551 VOUT_N.n1628 VOUT_N.n1627 1.11801
R552 VOUT_N.n1579 VOUT_N.n1578 1.11801
R553 VOUT_N.n1559 VOUT_N.n1558 1.11801
R554 VOUT_N.n1147 VOUT_N.n1146 1.11801
R555 VOUT_N.n1499 VOUT_N.n1498 1.11801
R556 VOUT_N.n1158 VOUT_N.n1157 1.11801
R557 VOUT_N.n574 VOUT_N.n538 1.11801
R558 VOUT_N.n575 VOUT_N.n536 1.11801
R559 VOUT_N.n466 VOUT_N.n465 1.11801
R560 VOUT_N.n454 VOUT_N.n453 1.11801
R561 VOUT_N.n413 VOUT_N.n412 1.11801
R562 VOUT_N.n410 VOUT_N.n409 1.11801
R563 VOUT_N.n364 VOUT_N.n363 1.11801
R564 VOUT_N.n355 VOUT_N.n354 1.11801
R565 VOUT_N.n457 VOUT_N.n456 1.11801
R566 VOUT_N.n1759 VOUT_N.n1758 1.11801
R567 VOUT_N.n1810 VOUT_N.n1725 1.11801
R568 VOUT_N.n2047 VOUT_N.n2046 1.11801
R569 VOUT_N.n2239 VOUT_N.n2238 1.11801
R570 VOUT_N.n2236 VOUT_N.n1820 1.11801
R571 VOUT_N.n2043 VOUT_N.n2008 1.11801
R572 VOUT_N.n611 VOUT_N.n610 1.11801
R573 VOUT_N.n1678 VOUT_N.n33 1.11801
R574 VOUT_N.n178 VOUT_N.n171 1.11801
R575 VOUT_N.n1976 VOUT_N.n1975 1.11782
R576 VOUT_N.n1971 VOUT_N.n1970 1.11782
R577 VOUT_N.n2004 VOUT_N.n2003 1.11782
R578 VOUT_N.n1885 VOUT_N.n1854 1.11782
R579 VOUT_N.n2121 VOUT_N.n2120 1.11782
R580 VOUT_N.n2125 VOUT_N.n2124 1.11782
R581 VOUT_N.n2198 VOUT_N.n2197 1.11782
R582 VOUT_N.n1257 VOUT_N.n1256 1.11782
R583 VOUT_N.n1486 VOUT_N.n1485 1.11782
R584 VOUT_N.n361 VOUT_N.n360 1.11782
R585 VOUT_N.n463 VOUT_N.n462 1.11782
R586 VOUT_N.n1805 VOUT_N.n1804 1.11782
R587 VOUT_N.n1809 VOUT_N.n1808 1.11782
R588 VOUT_N.n2242 VOUT_N.n2241 1.11782
R589 VOUT_N.n1677 VOUT_N.n1676 1.11782
R590 VOUT_N.n177 VOUT_N.n176 1.11782
R591 VOUT_N.n2244 VOUT_N.n2243 1.11782
R592 VOUT_N.n1705 VOUT_N.n1692 1.10737
R593 VOUT_N.n1943 VOUT_N.n1942 1.09451
R594 VOUT_N.n1965 VOUT_N.n1964 1.09451
R595 VOUT_N.n2138 VOUT_N.n2137 1.09451
R596 VOUT_N.n2157 VOUT_N.n2156 1.09451
R597 VOUT_N.n1698 VOUT_N.n1695 1.09451
R598 VOUT_N.n1719 VOUT_N.n1718 1.09451
R599 VOUT_N.n2108 VOUT_N.n2107 0.923611
R600 VOUT_N.n1865 VOUT_N.n1864 0.923611
R601 VOUT_N.n1871 VOUT_N.n1870 0.923589
R602 VOUT_N.n2102 VOUT_N.n2101 0.923589
R603 VOUT_N.n2178 VOUT_N.n2177 0.923589
R604 VOUT_N.n2190 VOUT_N.n2189 0.923589
R605 VOUT_N.n1980 VOUT_N.n1979 0.923589
R606 VOUT_N.n1985 VOUT_N.n1984 0.923589
R607 VOUT_N.n10 VOUT_N.n9 0.923589
R608 VOUT_N.n15 VOUT_N.n14 0.923589
R609 VOUT_N.n1739 VOUT_N.n1738 0.923589
R610 VOUT_N.n1744 VOUT_N.n1743 0.923589
R611 VOUT_N.n547 VOUT_N.n546 0.923538
R612 VOUT_N.n528 VOUT_N.n527 0.923538
R613 VOUT_N.n513 VOUT_N.n512 0.923538
R614 VOUT_N.n1829 VOUT_N.n1828 0.923538
R615 VOUT_N.n1844 VOUT_N.n1843 0.923538
R616 VOUT_N.n2017 VOUT_N.n2016 0.923538
R617 VOUT_N.n1995 VOUT_N.n1982 0.885703
R618 VOUT_N.n2193 VOUT_N.n2192 0.885703
R619 VOUT_N.n25 VOUT_N.n12 0.885703
R620 VOUT_N.n1722 VOUT_N.n1721 0.885703
R621 VOUT_N.n1754 VOUT_N.n1741 0.885703
R622 VOUT_N.n590 VOUT_N.n589 0.835535
R623 VOUT_N.n2219 VOUT_N.n2218 0.835535
R624 VOUT_N.n782 VOUT_N.n781 0.824999
R625 VOUT_N.n770 VOUT_N.n769 0.824999
R626 VOUT_N.n758 VOUT_N.n757 0.824999
R627 VOUT_N.n746 VOUT_N.n745 0.824999
R628 VOUT_N.n734 VOUT_N.n733 0.824999
R629 VOUT_N.n722 VOUT_N.n721 0.824999
R630 VOUT_N.n626 VOUT_N.n625 0.824999
R631 VOUT_N.n638 VOUT_N.n637 0.824999
R632 VOUT_N.n650 VOUT_N.n649 0.824999
R633 VOUT_N.n662 VOUT_N.n661 0.824999
R634 VOUT_N.n674 VOUT_N.n673 0.824999
R635 VOUT_N.n686 VOUT_N.n685 0.824999
R636 VOUT_N.n698 VOUT_N.n697 0.824999
R637 VOUT_N.n710 VOUT_N.n709 0.824999
R638 VOUT_N.n1117 VOUT_N.n1116 0.824999
R639 VOUT_N.n1105 VOUT_N.n1104 0.824999
R640 VOUT_N.n1093 VOUT_N.n1092 0.824999
R641 VOUT_N.n1081 VOUT_N.n1080 0.824999
R642 VOUT_N.n1069 VOUT_N.n1068 0.824999
R643 VOUT_N.n1057 VOUT_N.n1056 0.824999
R644 VOUT_N.n1045 VOUT_N.n1044 0.824999
R645 VOUT_N.n1033 VOUT_N.n1032 0.824999
R646 VOUT_N.n1021 VOUT_N.n1020 0.824999
R647 VOUT_N.n1009 VOUT_N.n1008 0.824999
R648 VOUT_N.n955 VOUT_N.n954 0.824999
R649 VOUT_N.n967 VOUT_N.n966 0.824999
R650 VOUT_N.n979 VOUT_N.n978 0.824999
R651 VOUT_N.n991 VOUT_N.n990 0.824999
R652 VOUT_N.n776 VOUT_N.n775 0.824997
R653 VOUT_N.n764 VOUT_N.n763 0.824997
R654 VOUT_N.n752 VOUT_N.n751 0.824997
R655 VOUT_N.n740 VOUT_N.n739 0.824997
R656 VOUT_N.n728 VOUT_N.n727 0.824997
R657 VOUT_N.n620 VOUT_N.n619 0.824997
R658 VOUT_N.n632 VOUT_N.n631 0.824997
R659 VOUT_N.n644 VOUT_N.n643 0.824997
R660 VOUT_N.n656 VOUT_N.n655 0.824997
R661 VOUT_N.n668 VOUT_N.n667 0.824997
R662 VOUT_N.n680 VOUT_N.n679 0.824997
R663 VOUT_N.n692 VOUT_N.n691 0.824997
R664 VOUT_N.n704 VOUT_N.n703 0.824997
R665 VOUT_N.n716 VOUT_N.n715 0.824997
R666 VOUT_N.n1111 VOUT_N.n1110 0.824997
R667 VOUT_N.n1099 VOUT_N.n1098 0.824997
R668 VOUT_N.n1087 VOUT_N.n1086 0.824997
R669 VOUT_N.n1075 VOUT_N.n1074 0.824997
R670 VOUT_N.n1063 VOUT_N.n1062 0.824997
R671 VOUT_N.n1051 VOUT_N.n1050 0.824997
R672 VOUT_N.n1039 VOUT_N.n1038 0.824997
R673 VOUT_N.n1027 VOUT_N.n1026 0.824997
R674 VOUT_N.n1015 VOUT_N.n1014 0.824997
R675 VOUT_N.n949 VOUT_N.n948 0.824997
R676 VOUT_N.n961 VOUT_N.n960 0.824997
R677 VOUT_N.n973 VOUT_N.n972 0.824997
R678 VOUT_N.n985 VOUT_N.n984 0.824997
R679 VOUT_N.n1003 VOUT_N.n1002 0.824997
R680 VOUT_N.n321 VOUT_N.n320 0.82495
R681 VOUT_N.n315 VOUT_N.n314 0.82495
R682 VOUT_N.n1449 VOUT_N.n1448 0.82495
R683 VOUT_N.n1443 VOUT_N.n1442 0.82495
R684 VOUT_N.n1428 VOUT_N.n1427 0.82495
R685 VOUT_N.n1422 VOUT_N.n1421 0.82495
R686 VOUT_N.n1407 VOUT_N.n1406 0.82495
R687 VOUT_N.n1401 VOUT_N.n1400 0.82495
R688 VOUT_N.n1386 VOUT_N.n1385 0.82495
R689 VOUT_N.n1380 VOUT_N.n1379 0.82495
R690 VOUT_N.n1365 VOUT_N.n1364 0.82495
R691 VOUT_N.n1359 VOUT_N.n1358 0.82495
R692 VOUT_N.n1312 VOUT_N.n1311 0.82495
R693 VOUT_N.n1318 VOUT_N.n1317 0.82495
R694 VOUT_N.n1333 VOUT_N.n1332 0.82495
R695 VOUT_N.n1339 VOUT_N.n1338 0.82495
R696 VOUT_N.n300 VOUT_N.n299 0.82495
R697 VOUT_N.n294 VOUT_N.n293 0.82495
R698 VOUT_N.n279 VOUT_N.n278 0.82495
R699 VOUT_N.n273 VOUT_N.n272 0.82495
R700 VOUT_N.n258 VOUT_N.n257 0.82495
R701 VOUT_N.n252 VOUT_N.n251 0.82495
R702 VOUT_N.n237 VOUT_N.n236 0.82495
R703 VOUT_N.n231 VOUT_N.n230 0.82495
R704 VOUT_N.n216 VOUT_N.n215 0.82495
R705 VOUT_N.n210 VOUT_N.n209 0.82495
R706 VOUT_N.n195 VOUT_N.n194 0.82495
R707 VOUT_N.n189 VOUT_N.n188 0.82495
R708 VOUT_N.n102 VOUT_N.n101 0.736598
R709 VOUT_N.n2085 VOUT_N.n2071 0.727104
R710 VOUT_N.n2163 VOUT_N.n2148 0.727104
R711 VOUT_N.n2168 VOUT_N.n2140 0.727104
R712 VOUT_N.n1955 VOUT_N.n1941 0.727104
R713 VOUT_N.n1880 VOUT_N.n1867 0.727104
R714 VOUT_N.n2112 VOUT_N.n2110 0.727104
R715 VOUT_N.n1290 VOUT_N.n957 0.727104
R716 VOUT_N.n1281 VOUT_N.n969 0.727104
R717 VOUT_N.n1272 VOUT_N.n981 0.727104
R718 VOUT_N.n1263 VOUT_N.n993 0.727104
R719 VOUT_N.n1121 VOUT_N.n1119 0.727104
R720 VOUT_N.n1130 VOUT_N.n1107 0.727104
R721 VOUT_N.n1161 VOUT_N.n1095 0.727104
R722 VOUT_N.n1170 VOUT_N.n1083 0.727104
R723 VOUT_N.n1179 VOUT_N.n1071 0.727104
R724 VOUT_N.n1188 VOUT_N.n1059 0.727104
R725 VOUT_N.n1207 VOUT_N.n1047 0.727104
R726 VOUT_N.n1216 VOUT_N.n1035 0.727104
R727 VOUT_N.n1225 VOUT_N.n1023 0.727104
R728 VOUT_N.n1234 VOUT_N.n1011 0.727104
R729 VOUT_N.n1662 VOUT_N.n1314 0.727104
R730 VOUT_N.n1653 VOUT_N.n1325 0.727104
R731 VOUT_N.n1644 VOUT_N.n1335 0.727104
R732 VOUT_N.n1635 VOUT_N.n1346 0.727104
R733 VOUT_N.n1458 VOUT_N.n1456 0.727104
R734 VOUT_N.n1467 VOUT_N.n1445 0.727104
R735 VOUT_N.n1502 VOUT_N.n1435 0.727104
R736 VOUT_N.n1511 VOUT_N.n1424 0.727104
R737 VOUT_N.n1520 VOUT_N.n1414 0.727104
R738 VOUT_N.n1529 VOUT_N.n1403 0.727104
R739 VOUT_N.n1582 VOUT_N.n1393 0.727104
R740 VOUT_N.n1591 VOUT_N.n1382 0.727104
R741 VOUT_N.n1600 VOUT_N.n1372 0.727104
R742 VOUT_N.n1609 VOUT_N.n1361 0.727104
R743 VOUT_N.n931 VOUT_N.n628 0.727104
R744 VOUT_N.n922 VOUT_N.n640 0.727104
R745 VOUT_N.n913 VOUT_N.n652 0.727104
R746 VOUT_N.n904 VOUT_N.n664 0.727104
R747 VOUT_N.n885 VOUT_N.n676 0.727104
R748 VOUT_N.n876 VOUT_N.n688 0.727104
R749 VOUT_N.n867 VOUT_N.n700 0.727104
R750 VOUT_N.n858 VOUT_N.n712 0.727104
R751 VOUT_N.n786 VOUT_N.n784 0.727104
R752 VOUT_N.n795 VOUT_N.n772 0.727104
R753 VOUT_N.n814 VOUT_N.n760 0.727104
R754 VOUT_N.n823 VOUT_N.n748 0.727104
R755 VOUT_N.n832 VOUT_N.n736 0.727104
R756 VOUT_N.n841 VOUT_N.n724 0.727104
R757 VOUT_N.n560 VOUT_N.n549 0.727104
R758 VOUT_N.n578 VOUT_N.n534 0.727104
R759 VOUT_N.n587 VOUT_N.n524 0.727104
R760 VOUT_N.n596 VOUT_N.n515 0.727104
R761 VOUT_N.n330 VOUT_N.n328 0.727104
R762 VOUT_N.n339 VOUT_N.n317 0.727104
R763 VOUT_N.n367 VOUT_N.n307 0.727104
R764 VOUT_N.n376 VOUT_N.n296 0.727104
R765 VOUT_N.n385 VOUT_N.n286 0.727104
R766 VOUT_N.n394 VOUT_N.n275 0.727104
R767 VOUT_N.n416 VOUT_N.n265 0.727104
R768 VOUT_N.n425 VOUT_N.n254 0.727104
R769 VOUT_N.n434 VOUT_N.n244 0.727104
R770 VOUT_N.n443 VOUT_N.n233 0.727104
R771 VOUT_N.n469 VOUT_N.n223 0.727104
R772 VOUT_N.n478 VOUT_N.n212 0.727104
R773 VOUT_N.n487 VOUT_N.n202 0.727104
R774 VOUT_N.n496 VOUT_N.n191 0.727104
R775 VOUT_N.n1795 VOUT_N.n1781 0.727104
R776 VOUT_N.n2230 VOUT_N.n1825 0.727104
R777 VOUT_N.n2221 VOUT_N.n1835 0.727104
R778 VOUT_N.n2212 VOUT_N.n1846 0.727104
R779 VOUT_N.n2037 VOUT_N.n2013 0.727104
R780 VOUT_N.n1919 VOUT_N.n1906 0.726858
R781 VOUT_N.n1800 VOUT_N.n1773 0.726858
R782 VOUT_N.n2028 VOUT_N.n2023 0.726858
R783 VOUT_N.n1177 VOUT_N.n1176 0.685007
R784 VOUT_N.n1223 VOUT_N.n1222 0.685007
R785 VOUT_N.n1279 VOUT_N.n1278 0.685007
R786 VOUT_N.n830 VOUT_N.n829 0.685007
R787 VOUT_N.n874 VOUT_N.n873 0.685007
R788 VOUT_N.n920 VOUT_N.n919 0.685007
R789 VOUT_N.n2243 VOUT_N.n2242 0.659441
R790 VOUT_N.n1968 VOUT_N.n1967 0.617177
R791 VOUT_N.n335 VOUT_N.n323 0.616779
R792 VOUT_N.n555 VOUT_N.n553 0.616779
R793 VOUT_N.n564 VOUT_N.n543 0.616779
R794 VOUT_N.n1875 VOUT_N.n1873 0.616779
R795 VOUT_N.n2117 VOUT_N.n2104 0.616779
R796 VOUT_N.n1950 VOUT_N.n1948 0.616779
R797 VOUT_N.n1923 VOUT_N.n1898 0.616779
R798 VOUT_N.n2081 VOUT_N.n2080 0.616779
R799 VOUT_N.n2090 VOUT_N.n2063 0.616779
R800 VOUT_N.n582 VOUT_N.n530 0.616779
R801 VOUT_N.n591 VOUT_N.n519 0.616779
R802 VOUT_N.n600 VOUT_N.n509 0.616779
R803 VOUT_N.n791 VOUT_N.n778 0.616779
R804 VOUT_N.n800 VOUT_N.n766 0.616779
R805 VOUT_N.n819 VOUT_N.n754 0.616779
R806 VOUT_N.n828 VOUT_N.n742 0.616779
R807 VOUT_N.n837 VOUT_N.n730 0.616779
R808 VOUT_N.n936 VOUT_N.n622 0.616779
R809 VOUT_N.n927 VOUT_N.n634 0.616779
R810 VOUT_N.n918 VOUT_N.n646 0.616779
R811 VOUT_N.n909 VOUT_N.n658 0.616779
R812 VOUT_N.n890 VOUT_N.n670 0.616779
R813 VOUT_N.n881 VOUT_N.n682 0.616779
R814 VOUT_N.n872 VOUT_N.n694 0.616779
R815 VOUT_N.n863 VOUT_N.n706 0.616779
R816 VOUT_N.n846 VOUT_N.n718 0.616779
R817 VOUT_N.n1463 VOUT_N.n1451 0.616779
R818 VOUT_N.n1472 VOUT_N.n1439 0.616779
R819 VOUT_N.n1507 VOUT_N.n1430 0.616779
R820 VOUT_N.n1516 VOUT_N.n1418 0.616779
R821 VOUT_N.n1525 VOUT_N.n1409 0.616779
R822 VOUT_N.n1534 VOUT_N.n1397 0.616779
R823 VOUT_N.n1587 VOUT_N.n1388 0.616779
R824 VOUT_N.n1596 VOUT_N.n1376 0.616779
R825 VOUT_N.n1605 VOUT_N.n1367 0.616779
R826 VOUT_N.n1667 VOUT_N.n1308 0.616779
R827 VOUT_N.n1658 VOUT_N.n1320 0.616779
R828 VOUT_N.n1649 VOUT_N.n1329 0.616779
R829 VOUT_N.n1640 VOUT_N.n1341 0.616779
R830 VOUT_N.n1614 VOUT_N.n1355 0.616779
R831 VOUT_N.n1126 VOUT_N.n1113 0.616779
R832 VOUT_N.n1135 VOUT_N.n1101 0.616779
R833 VOUT_N.n1166 VOUT_N.n1089 0.616779
R834 VOUT_N.n1175 VOUT_N.n1077 0.616779
R835 VOUT_N.n1184 VOUT_N.n1065 0.616779
R836 VOUT_N.n1193 VOUT_N.n1053 0.616779
R837 VOUT_N.n1212 VOUT_N.n1041 0.616779
R838 VOUT_N.n1221 VOUT_N.n1029 0.616779
R839 VOUT_N.n1230 VOUT_N.n1017 0.616779
R840 VOUT_N.n1295 VOUT_N.n951 0.616779
R841 VOUT_N.n1286 VOUT_N.n963 0.616779
R842 VOUT_N.n1277 VOUT_N.n975 0.616779
R843 VOUT_N.n1268 VOUT_N.n987 0.616779
R844 VOUT_N.n1239 VOUT_N.n1005 0.616779
R845 VOUT_N.n344 VOUT_N.n311 0.616779
R846 VOUT_N.n372 VOUT_N.n302 0.616779
R847 VOUT_N.n381 VOUT_N.n290 0.616779
R848 VOUT_N.n390 VOUT_N.n281 0.616779
R849 VOUT_N.n399 VOUT_N.n269 0.616779
R850 VOUT_N.n421 VOUT_N.n260 0.616779
R851 VOUT_N.n430 VOUT_N.n248 0.616779
R852 VOUT_N.n439 VOUT_N.n239 0.616779
R853 VOUT_N.n448 VOUT_N.n227 0.616779
R854 VOUT_N.n474 VOUT_N.n218 0.616779
R855 VOUT_N.n483 VOUT_N.n206 0.616779
R856 VOUT_N.n492 VOUT_N.n197 0.616779
R857 VOUT_N.n501 VOUT_N.n185 0.616779
R858 VOUT_N.n2225 VOUT_N.n1831 0.616779
R859 VOUT_N.n2216 VOUT_N.n1840 0.616779
R860 VOUT_N.n2207 VOUT_N.n1850 0.616779
R861 VOUT_N.n2032 VOUT_N.n2019 0.616779
R862 VOUT_N.n320 VOUT_N.t268 0.607167
R863 VOUT_N.n320 VOUT_N.n319 0.607167
R864 VOUT_N.n314 VOUT_N.t220 0.607167
R865 VOUT_N.n314 VOUT_N.n313 0.607167
R866 VOUT_N.n781 VOUT_N.t235 0.607167
R867 VOUT_N.n781 VOUT_N.n780 0.607167
R868 VOUT_N.n775 VOUT_N.t138 0.607167
R869 VOUT_N.n775 VOUT_N.n774 0.607167
R870 VOUT_N.n769 VOUT_N.t270 0.607167
R871 VOUT_N.n769 VOUT_N.n768 0.607167
R872 VOUT_N.n763 VOUT_N.t140 0.607167
R873 VOUT_N.n763 VOUT_N.n762 0.607167
R874 VOUT_N.n757 VOUT_N.t131 0.607167
R875 VOUT_N.n757 VOUT_N.n756 0.607167
R876 VOUT_N.n751 VOUT_N.t84 0.607167
R877 VOUT_N.n751 VOUT_N.n750 0.607167
R878 VOUT_N.n745 VOUT_N.t228 0.607167
R879 VOUT_N.n745 VOUT_N.n744 0.607167
R880 VOUT_N.n739 VOUT_N.t184 0.607167
R881 VOUT_N.n739 VOUT_N.n738 0.607167
R882 VOUT_N.n733 VOUT_N.t114 0.607167
R883 VOUT_N.n733 VOUT_N.n732 0.607167
R884 VOUT_N.n727 VOUT_N.t154 0.607167
R885 VOUT_N.n727 VOUT_N.n726 0.607167
R886 VOUT_N.n721 VOUT_N.t160 0.607167
R887 VOUT_N.n721 VOUT_N.n720 0.607167
R888 VOUT_N.n619 VOUT_N.t258 0.607167
R889 VOUT_N.n619 VOUT_N.n618 0.607167
R890 VOUT_N.n625 VOUT_N.t123 0.607167
R891 VOUT_N.n625 VOUT_N.n624 0.607167
R892 VOUT_N.n631 VOUT_N.t178 0.607167
R893 VOUT_N.n631 VOUT_N.n630 0.607167
R894 VOUT_N.n637 VOUT_N.t97 0.607167
R895 VOUT_N.n637 VOUT_N.n636 0.607167
R896 VOUT_N.n643 VOUT_N.t137 0.607167
R897 VOUT_N.n643 VOUT_N.n642 0.607167
R898 VOUT_N.n649 VOUT_N.t247 0.607167
R899 VOUT_N.n649 VOUT_N.n648 0.607167
R900 VOUT_N.n655 VOUT_N.t238 0.607167
R901 VOUT_N.n655 VOUT_N.n654 0.607167
R902 VOUT_N.n661 VOUT_N.t185 0.607167
R903 VOUT_N.n661 VOUT_N.n660 0.607167
R904 VOUT_N.n667 VOUT_N.t99 0.607167
R905 VOUT_N.n667 VOUT_N.n666 0.607167
R906 VOUT_N.n673 VOUT_N.t200 0.607167
R907 VOUT_N.n673 VOUT_N.n672 0.607167
R908 VOUT_N.n679 VOUT_N.t193 0.607167
R909 VOUT_N.n679 VOUT_N.n678 0.607167
R910 VOUT_N.n685 VOUT_N.t214 0.607167
R911 VOUT_N.n685 VOUT_N.n684 0.607167
R912 VOUT_N.n691 VOUT_N.t124 0.607167
R913 VOUT_N.n691 VOUT_N.n690 0.607167
R914 VOUT_N.n697 VOUT_N.t147 0.607167
R915 VOUT_N.n697 VOUT_N.n696 0.607167
R916 VOUT_N.n703 VOUT_N.t218 0.607167
R917 VOUT_N.n703 VOUT_N.n702 0.607167
R918 VOUT_N.n709 VOUT_N.t110 0.607167
R919 VOUT_N.n709 VOUT_N.n708 0.607167
R920 VOUT_N.n715 VOUT_N.t85 0.607167
R921 VOUT_N.n715 VOUT_N.n714 0.607167
R922 VOUT_N.n1448 VOUT_N.t207 0.607167
R923 VOUT_N.n1448 VOUT_N.n1447 0.607167
R924 VOUT_N.n1442 VOUT_N.t116 0.607167
R925 VOUT_N.n1442 VOUT_N.n1441 0.607167
R926 VOUT_N.n1427 VOUT_N.t155 0.607167
R927 VOUT_N.n1427 VOUT_N.n1426 0.607167
R928 VOUT_N.n1421 VOUT_N.t78 0.607167
R929 VOUT_N.n1421 VOUT_N.n1420 0.607167
R930 VOUT_N.n1406 VOUT_N.t80 0.607167
R931 VOUT_N.n1406 VOUT_N.n1405 0.607167
R932 VOUT_N.n1400 VOUT_N.t260 0.607167
R933 VOUT_N.n1400 VOUT_N.n1399 0.607167
R934 VOUT_N.n1385 VOUT_N.t95 0.607167
R935 VOUT_N.n1385 VOUT_N.n1384 0.607167
R936 VOUT_N.n1379 VOUT_N.t146 0.607167
R937 VOUT_N.n1379 VOUT_N.n1378 0.607167
R938 VOUT_N.n1364 VOUT_N.t179 0.607167
R939 VOUT_N.n1364 VOUT_N.n1363 0.607167
R940 VOUT_N.n1358 VOUT_N.t120 0.607167
R941 VOUT_N.n1358 VOUT_N.n1357 0.607167
R942 VOUT_N.n1311 VOUT_N.t239 0.607167
R943 VOUT_N.n1311 VOUT_N.n1310 0.607167
R944 VOUT_N.n1317 VOUT_N.t221 0.607167
R945 VOUT_N.n1317 VOUT_N.n1316 0.607167
R946 VOUT_N.n1332 VOUT_N.t139 0.607167
R947 VOUT_N.n1332 VOUT_N.n1331 0.607167
R948 VOUT_N.n1338 VOUT_N.t232 0.607167
R949 VOUT_N.n1338 VOUT_N.n1337 0.607167
R950 VOUT_N.n1116 VOUT_N.t256 0.607167
R951 VOUT_N.n1116 VOUT_N.n1115 0.607167
R952 VOUT_N.n1110 VOUT_N.t201 0.607167
R953 VOUT_N.n1110 VOUT_N.n1109 0.607167
R954 VOUT_N.n1104 VOUT_N.t263 0.607167
R955 VOUT_N.n1104 VOUT_N.n1103 0.607167
R956 VOUT_N.n1098 VOUT_N.t248 0.607167
R957 VOUT_N.n1098 VOUT_N.n1097 0.607167
R958 VOUT_N.n1092 VOUT_N.t101 0.607167
R959 VOUT_N.n1092 VOUT_N.n1091 0.607167
R960 VOUT_N.n1086 VOUT_N.t208 0.607167
R961 VOUT_N.n1086 VOUT_N.n1085 0.607167
R962 VOUT_N.n1080 VOUT_N.t202 0.607167
R963 VOUT_N.n1080 VOUT_N.n1079 0.607167
R964 VOUT_N.n1074 VOUT_N.t121 0.607167
R965 VOUT_N.n1074 VOUT_N.n1073 0.607167
R966 VOUT_N.n1068 VOUT_N.t82 0.607167
R967 VOUT_N.n1068 VOUT_N.n1067 0.607167
R968 VOUT_N.n1062 VOUT_N.t223 0.607167
R969 VOUT_N.n1062 VOUT_N.n1061 0.607167
R970 VOUT_N.n1056 VOUT_N.t188 0.607167
R971 VOUT_N.n1056 VOUT_N.n1055 0.607167
R972 VOUT_N.n1050 VOUT_N.t246 0.607167
R973 VOUT_N.n1050 VOUT_N.n1049 0.607167
R974 VOUT_N.n1044 VOUT_N.t89 0.607167
R975 VOUT_N.n1044 VOUT_N.n1043 0.607167
R976 VOUT_N.n1038 VOUT_N.t83 0.607167
R977 VOUT_N.n1038 VOUT_N.n1037 0.607167
R978 VOUT_N.n1032 VOUT_N.t148 0.607167
R979 VOUT_N.n1032 VOUT_N.n1031 0.607167
R980 VOUT_N.n1026 VOUT_N.t265 0.607167
R981 VOUT_N.n1026 VOUT_N.n1025 0.607167
R982 VOUT_N.n1020 VOUT_N.t197 0.607167
R983 VOUT_N.n1020 VOUT_N.n1019 0.607167
R984 VOUT_N.n1014 VOUT_N.t205 0.607167
R985 VOUT_N.n1014 VOUT_N.n1013 0.607167
R986 VOUT_N.n1008 VOUT_N.t163 0.607167
R987 VOUT_N.n1008 VOUT_N.n1007 0.607167
R988 VOUT_N.n948 VOUT_N.t77 0.607167
R989 VOUT_N.n948 VOUT_N.n947 0.607167
R990 VOUT_N.n954 VOUT_N.t181 0.607167
R991 VOUT_N.n954 VOUT_N.n953 0.607167
R992 VOUT_N.n960 VOUT_N.t261 0.607167
R993 VOUT_N.n960 VOUT_N.n959 0.607167
R994 VOUT_N.n966 VOUT_N.t142 0.607167
R995 VOUT_N.n966 VOUT_N.n965 0.607167
R996 VOUT_N.n972 VOUT_N.t164 0.607167
R997 VOUT_N.n972 VOUT_N.n971 0.607167
R998 VOUT_N.n978 VOUT_N.t126 0.607167
R999 VOUT_N.n978 VOUT_N.n977 0.607167
R1000 VOUT_N.n984 VOUT_N.t182 0.607167
R1001 VOUT_N.n984 VOUT_N.n983 0.607167
R1002 VOUT_N.n990 VOUT_N.t167 0.607167
R1003 VOUT_N.n990 VOUT_N.n989 0.607167
R1004 VOUT_N.n1002 VOUT_N.t170 0.607167
R1005 VOUT_N.n1002 VOUT_N.n1001 0.607167
R1006 VOUT_N.n299 VOUT_N.t254 0.607167
R1007 VOUT_N.n299 VOUT_N.n298 0.607167
R1008 VOUT_N.n293 VOUT_N.t172 0.607167
R1009 VOUT_N.n293 VOUT_N.n292 0.607167
R1010 VOUT_N.n278 VOUT_N.t198 0.607167
R1011 VOUT_N.n278 VOUT_N.n277 0.607167
R1012 VOUT_N.n272 VOUT_N.t253 0.607167
R1013 VOUT_N.n272 VOUT_N.n271 0.607167
R1014 VOUT_N.n257 VOUT_N.t175 0.607167
R1015 VOUT_N.n257 VOUT_N.n256 0.607167
R1016 VOUT_N.n251 VOUT_N.t100 0.607167
R1017 VOUT_N.n251 VOUT_N.n250 0.607167
R1018 VOUT_N.n236 VOUT_N.t109 0.607167
R1019 VOUT_N.n236 VOUT_N.n235 0.607167
R1020 VOUT_N.n230 VOUT_N.t215 0.607167
R1021 VOUT_N.n230 VOUT_N.n229 0.607167
R1022 VOUT_N.n215 VOUT_N.t244 0.607167
R1023 VOUT_N.n215 VOUT_N.n214 0.607167
R1024 VOUT_N.n209 VOUT_N.t94 0.607167
R1025 VOUT_N.n209 VOUT_N.n208 0.607167
R1026 VOUT_N.n194 VOUT_N.t115 0.607167
R1027 VOUT_N.n194 VOUT_N.n193 0.607167
R1028 VOUT_N.n188 VOUT_N.t133 0.607167
R1029 VOUT_N.n188 VOUT_N.n187 0.607167
R1030 VOUT_N.n546 VOUT_N.t34 0.5465
R1031 VOUT_N.n546 VOUT_N.n545 0.5465
R1032 VOUT_N.n2107 VOUT_N.t3 0.5465
R1033 VOUT_N.n2107 VOUT_N.n2106 0.5465
R1034 VOUT_N.n1870 VOUT_N.t26 0.5465
R1035 VOUT_N.n1870 VOUT_N.n1869 0.5465
R1036 VOUT_N.n1864 VOUT_N.t12 0.5465
R1037 VOUT_N.n1864 VOUT_N.n1863 0.5465
R1038 VOUT_N.n2101 VOUT_N.t30 0.5465
R1039 VOUT_N.n2101 VOUT_N.n2100 0.5465
R1040 VOUT_N.n2156 VOUT_N.n2155 0.5465
R1041 VOUT_N.n2077 VOUT_N.n2076 0.5465
R1042 VOUT_N.n1908 VOUT_N.t25 0.5465
R1043 VOUT_N.n1942 VOUT_N.t17 0.5465
R1044 VOUT_N.n1895 VOUT_N.n1894 0.5465
R1045 VOUT_N.n1964 VOUT_N.n1963 0.5465
R1046 VOUT_N.n1902 VOUT_N.t21 0.5465
R1047 VOUT_N.n1902 VOUT_N.n1901 0.5465
R1048 VOUT_N.n1938 VOUT_N.t24 0.5465
R1049 VOUT_N.n1938 VOUT_N.n1937 0.5465
R1050 VOUT_N.n2067 VOUT_N.t14 0.5465
R1051 VOUT_N.n2067 VOUT_N.n2066 0.5465
R1052 VOUT_N.n2145 VOUT_N.t9 0.5465
R1053 VOUT_N.n2145 VOUT_N.n2144 0.5465
R1054 VOUT_N.n2060 VOUT_N.t29 0.5465
R1055 VOUT_N.n2137 VOUT_N.t28 0.5465
R1056 VOUT_N.n2177 VOUT_N.t16 0.5465
R1057 VOUT_N.n2177 VOUT_N.n2176 0.5465
R1058 VOUT_N.n2189 VOUT_N.t32 0.5465
R1059 VOUT_N.n2189 VOUT_N.n2188 0.5465
R1060 VOUT_N.n1979 VOUT_N.t15 0.5465
R1061 VOUT_N.n1979 VOUT_N.n1978 0.5465
R1062 VOUT_N.n1984 VOUT_N.t19 0.5465
R1063 VOUT_N.n1984 VOUT_N.n1983 0.5465
R1064 VOUT_N.n527 VOUT_N.t31 0.5465
R1065 VOUT_N.n527 VOUT_N.n526 0.5465
R1066 VOUT_N.n512 VOUT_N.t36 0.5465
R1067 VOUT_N.n512 VOUT_N.n511 0.5465
R1068 VOUT_N.n9 VOUT_N.t18 0.5465
R1069 VOUT_N.n9 VOUT_N.n8 0.5465
R1070 VOUT_N.n14 VOUT_N.t33 0.5465
R1071 VOUT_N.n14 VOUT_N.n13 0.5465
R1072 VOUT_N.n1769 VOUT_N.n1768 0.5465
R1073 VOUT_N.n1707 VOUT_N.t11 0.5465
R1074 VOUT_N.n1707 VOUT_N.n1706 0.5465
R1075 VOUT_N.n1777 VOUT_N.t22 0.5465
R1076 VOUT_N.n1777 VOUT_N.n1776 0.5465
R1077 VOUT_N.n1695 VOUT_N.t5 0.5465
R1078 VOUT_N.n1785 VOUT_N.t27 0.5465
R1079 VOUT_N.n1718 VOUT_N.n1717 0.5465
R1080 VOUT_N.n1738 VOUT_N.t10 0.5465
R1081 VOUT_N.n1738 VOUT_N.n1737 0.5465
R1082 VOUT_N.n1743 VOUT_N.t35 0.5465
R1083 VOUT_N.n1743 VOUT_N.n1742 0.5465
R1084 VOUT_N.n1828 VOUT_N.t8 0.5465
R1085 VOUT_N.n1828 VOUT_N.n1827 0.5465
R1086 VOUT_N.n1843 VOUT_N.t7 0.5465
R1087 VOUT_N.n1843 VOUT_N.n1842 0.5465
R1088 VOUT_N.n2016 VOUT_N.t20 0.5465
R1089 VOUT_N.n2016 VOUT_N.n2015 0.5465
R1090 VOUT_N.n1518 VOUT_N.n1517 0.482824
R1091 VOUT_N.n1598 VOUT_N.n1597 0.482824
R1092 VOUT_N.n1651 VOUT_N.n1650 0.482824
R1093 VOUT_N.n383 VOUT_N.n382 0.482824
R1094 VOUT_N.n432 VOUT_N.n431 0.482824
R1095 VOUT_N.n485 VOUT_N.n484 0.482824
R1096 VOUT_N.n151 VOUT_N.n150 0.469524
R1097 VOUT_N.n92 VOUT_N.n71 0.469524
R1098 VOUT_N.n2196 VOUT_N.n2195 0.468246
R1099 VOUT_N.n1998 VOUT_N.n1997 0.468246
R1100 VOUT_N.n2120 VOUT_N.n2118 0.468246
R1101 VOUT_N.n1883 VOUT_N.n1882 0.468246
R1102 VOUT_N.n28 VOUT_N.n27 0.468246
R1103 VOUT_N.n1757 VOUT_N.n1756 0.468246
R1104 VOUT_N.n103 VOUT_N.n102 0.4505
R1105 VOUT_N.n84 VOUT_N.n75 0.4505
R1106 VOUT_N.n90 VOUT_N.n74 0.4505
R1107 VOUT_N.n65 VOUT_N.n62 0.4505
R1108 VOUT_N.n1297 VOUT_N.n1296 0.43212
R1109 VOUT_N.n938 VOUT_N.n937 0.43212
R1110 VOUT_N.n1195 VOUT_N.n1194 0.431486
R1111 VOUT_N.n848 VOUT_N.n847 0.431486
R1112 VOUT_N.n1241 VOUT_N.n1240 0.428951
R1113 VOUT_N.n892 VOUT_N.n891 0.428951
R1114 VOUT_N.n608 VOUT_N.n607 0.428
R1115 VOUT_N.n33 VOUT_N.n32 0.428
R1116 VOUT_N.n2240 VOUT_N.n2239 0.428
R1117 VOUT_N.n1137 VOUT_N.n1136 0.415007
R1118 VOUT_N.n1159 VOUT_N.n1158 0.415007
R1119 VOUT_N.n1261 VOUT_N.n1260 0.415007
R1120 VOUT_N.n802 VOUT_N.n801 0.415007
R1121 VOUT_N.n812 VOUT_N.n811 0.415007
R1122 VOUT_N.n902 VOUT_N.n901 0.415007
R1123 VOUT_N.n1205 VOUT_N.n1204 0.408669
R1124 VOUT_N.n856 VOUT_N.n855 0.408669
R1125 VOUT_N.n1547 VOUT_N.n1546 0.395359
R1126 VOUT_N.n613 VOUT_N.n612 0.395359
R1127 VOUT_N.n1465 VOUT_N.n1464 0.389021
R1128 VOUT_N.n1509 VOUT_N.n1508 0.389021
R1129 VOUT_N.n1527 VOUT_N.n1526 0.389021
R1130 VOUT_N.n1589 VOUT_N.n1588 0.389021
R1131 VOUT_N.n1607 VOUT_N.n1606 0.389021
R1132 VOUT_N.n1642 VOUT_N.n1641 0.389021
R1133 VOUT_N.n1660 VOUT_N.n1659 0.389021
R1134 VOUT_N.n337 VOUT_N.n336 0.389021
R1135 VOUT_N.n374 VOUT_N.n373 0.389021
R1136 VOUT_N.n392 VOUT_N.n391 0.389021
R1137 VOUT_N.n423 VOUT_N.n422 0.389021
R1138 VOUT_N.n441 VOUT_N.n440 0.389021
R1139 VOUT_N.n476 VOUT_N.n475 0.389021
R1140 VOUT_N.n494 VOUT_N.n493 0.389021
R1141 VOUT_N.n2092 VOUT_N.n2091 0.366838
R1142 VOUT_N.n1926 VOUT_N.n1925 0.366838
R1143 VOUT_N.n2171 VOUT_N.n2170 0.366838
R1144 VOUT_N.n1970 VOUT_N.n1969 0.366838
R1145 VOUT_N.n603 VOUT_N.n602 0.366838
R1146 VOUT_N.n576 VOUT_N.n575 0.366838
R1147 VOUT_N.n567 VOUT_N.n566 0.366838
R1148 VOUT_N.n1725 VOUT_N.n1724 0.366838
R1149 VOUT_N.n1803 VOUT_N.n1802 0.366838
R1150 VOUT_N.n2233 VOUT_N.n2232 0.366838
R1151 VOUT_N.n2206 VOUT_N.n2205 0.366838
R1152 VOUT_N.n2040 VOUT_N.n2039 0.366838
R1153 VOUT_N.n2000 VOUT_N.n1976 0.356063
R1154 VOUT_N.n1859 VOUT_N.n1858 0.356063
R1155 VOUT_N.n2198 VOUT_N.n2174 0.356063
R1156 VOUT_N.n1814 VOUT_N.n1813 0.356063
R1157 VOUT_N.n1730 VOUT_N.n1729 0.356063
R1158 VOUT_N.n1974 VOUT_N.n1973 0.345923
R1159 VOUT_N.n572 VOUT_N.n571 0.345923
R1160 VOUT_N.n2048 VOUT_N.n2047 0.345923
R1161 VOUT_N.n1904 VOUT_N.n1900 0.336464
R1162 VOUT_N.n2069 VOUT_N.n2065 0.336464
R1163 VOUT_N.n2058 VOUT_N.n2057 0.336464
R1164 VOUT_N.n2074 VOUT_N.n2073 0.336464
R1165 VOUT_N.n1779 VOUT_N.n1775 0.336464
R1166 VOUT_N.n1787 VOUT_N.n1784 0.336464
R1167 VOUT_N.n1771 VOUT_N.n1767 0.336464
R1168 VOUT_N.n1669 VOUT_N.n1668 0.330394
R1169 VOUT_N.n503 VOUT_N.n502 0.330394
R1170 VOUT_N.n1536 VOUT_N.n1535 0.329761
R1171 VOUT_N.n401 VOUT_N.n400 0.329761
R1172 VOUT_N.n1616 VOUT_N.n1615 0.327225
R1173 VOUT_N.n450 VOUT_N.n449 0.327225
R1174 VOUT_N.n1474 VOUT_N.n1473 0.313282
R1175 VOUT_N.n1500 VOUT_N.n1499 0.313282
R1176 VOUT_N.n1633 VOUT_N.n1632 0.313282
R1177 VOUT_N.n346 VOUT_N.n345 0.313282
R1178 VOUT_N.n365 VOUT_N.n364 0.313282
R1179 VOUT_N.n467 VOUT_N.n466 0.313282
R1180 VOUT_N.n1580 VOUT_N.n1579 0.306944
R1181 VOUT_N.n414 VOUT_N.n413 0.306944
R1182 VOUT_N.n999 VOUT_N.n998 0.2705
R1183 VOUT_N.n1256 VOUT_N.n1255 0.2705
R1184 VOUT_N.n1552 VOUT_N.n1551 0.2705
R1185 VOUT_N.n1569 VOUT_N.n1568 0.2705
R1186 VOUT_N.n1145 VOUT_N.n1144 0.2705
R1187 VOUT_N.n1156 VOUT_N.n1155 0.2705
R1188 VOUT_N.n943 VOUT_N.n942 0.2705
R1189 VOUT_N.n1677 VOUT_N.n1673 0.238176
R1190 VOUT_N.n1930 VOUT_N.n1929 0.231204
R1191 VOUT_N.n2131 VOUT_N.n2130 0.231204
R1192 VOUT_N.n1809 VOUT_N.n1805 0.231204
R1193 VOUT_N.n1910 VOUT_N.n1907 0.191654
R1194 VOUT_N.n1892 VOUT_N.n1891 0.191654
R1195 VOUT_N.n2083 VOUT_N.n2082 0.186204
R1196 VOUT_N.n2088 VOUT_N.n2087 0.186204
R1197 VOUT_N.n1922 VOUT_N.n1921 0.186204
R1198 VOUT_N.n1917 VOUT_N.n1916 0.186204
R1199 VOUT_N.n2161 VOUT_N.n2160 0.186204
R1200 VOUT_N.n2166 VOUT_N.n2165 0.186204
R1201 VOUT_N.n1958 VOUT_N.n1957 0.186204
R1202 VOUT_N.n1953 VOUT_N.n1952 0.186204
R1203 VOUT_N.n2185 VOUT_N.n2184 0.186204
R1204 VOUT_N.n1993 VOUT_N.n1992 0.186204
R1205 VOUT_N.n2115 VOUT_N.n2114 0.186204
R1206 VOUT_N.n1878 VOUT_N.n1877 0.186204
R1207 VOUT_N.n1124 VOUT_N.n1123 0.186204
R1208 VOUT_N.n1128 VOUT_N.n1127 0.186204
R1209 VOUT_N.n1133 VOUT_N.n1132 0.186204
R1210 VOUT_N.n1164 VOUT_N.n1163 0.186204
R1211 VOUT_N.n1168 VOUT_N.n1167 0.186204
R1212 VOUT_N.n1173 VOUT_N.n1172 0.186204
R1213 VOUT_N.n1182 VOUT_N.n1181 0.186204
R1214 VOUT_N.n1186 VOUT_N.n1185 0.186204
R1215 VOUT_N.n1191 VOUT_N.n1190 0.186204
R1216 VOUT_N.n1210 VOUT_N.n1209 0.186204
R1217 VOUT_N.n1214 VOUT_N.n1213 0.186204
R1218 VOUT_N.n1219 VOUT_N.n1218 0.186204
R1219 VOUT_N.n1228 VOUT_N.n1227 0.186204
R1220 VOUT_N.n1232 VOUT_N.n1231 0.186204
R1221 VOUT_N.n1237 VOUT_N.n1236 0.186204
R1222 VOUT_N.n1266 VOUT_N.n1265 0.186204
R1223 VOUT_N.n1270 VOUT_N.n1269 0.186204
R1224 VOUT_N.n1275 VOUT_N.n1274 0.186204
R1225 VOUT_N.n1284 VOUT_N.n1283 0.186204
R1226 VOUT_N.n1288 VOUT_N.n1287 0.186204
R1227 VOUT_N.n1293 VOUT_N.n1292 0.186204
R1228 VOUT_N.n1461 VOUT_N.n1460 0.186204
R1229 VOUT_N.n1470 VOUT_N.n1469 0.186204
R1230 VOUT_N.n1505 VOUT_N.n1504 0.186204
R1231 VOUT_N.n1514 VOUT_N.n1513 0.186204
R1232 VOUT_N.n1523 VOUT_N.n1522 0.186204
R1233 VOUT_N.n1532 VOUT_N.n1531 0.186204
R1234 VOUT_N.n1585 VOUT_N.n1584 0.186204
R1235 VOUT_N.n1594 VOUT_N.n1593 0.186204
R1236 VOUT_N.n1603 VOUT_N.n1602 0.186204
R1237 VOUT_N.n1612 VOUT_N.n1611 0.186204
R1238 VOUT_N.n1638 VOUT_N.n1637 0.186204
R1239 VOUT_N.n1647 VOUT_N.n1646 0.186204
R1240 VOUT_N.n1656 VOUT_N.n1655 0.186204
R1241 VOUT_N.n1665 VOUT_N.n1664 0.186204
R1242 VOUT_N.n789 VOUT_N.n788 0.186204
R1243 VOUT_N.n793 VOUT_N.n792 0.186204
R1244 VOUT_N.n798 VOUT_N.n797 0.186204
R1245 VOUT_N.n817 VOUT_N.n816 0.186204
R1246 VOUT_N.n821 VOUT_N.n820 0.186204
R1247 VOUT_N.n826 VOUT_N.n825 0.186204
R1248 VOUT_N.n835 VOUT_N.n834 0.186204
R1249 VOUT_N.n839 VOUT_N.n838 0.186204
R1250 VOUT_N.n844 VOUT_N.n843 0.186204
R1251 VOUT_N.n861 VOUT_N.n860 0.186204
R1252 VOUT_N.n865 VOUT_N.n864 0.186204
R1253 VOUT_N.n870 VOUT_N.n869 0.186204
R1254 VOUT_N.n879 VOUT_N.n878 0.186204
R1255 VOUT_N.n883 VOUT_N.n882 0.186204
R1256 VOUT_N.n888 VOUT_N.n887 0.186204
R1257 VOUT_N.n907 VOUT_N.n906 0.186204
R1258 VOUT_N.n911 VOUT_N.n910 0.186204
R1259 VOUT_N.n916 VOUT_N.n915 0.186204
R1260 VOUT_N.n925 VOUT_N.n924 0.186204
R1261 VOUT_N.n929 VOUT_N.n928 0.186204
R1262 VOUT_N.n934 VOUT_N.n933 0.186204
R1263 VOUT_N.n333 VOUT_N.n332 0.186204
R1264 VOUT_N.n342 VOUT_N.n341 0.186204
R1265 VOUT_N.n370 VOUT_N.n369 0.186204
R1266 VOUT_N.n379 VOUT_N.n378 0.186204
R1267 VOUT_N.n388 VOUT_N.n387 0.186204
R1268 VOUT_N.n397 VOUT_N.n396 0.186204
R1269 VOUT_N.n419 VOUT_N.n418 0.186204
R1270 VOUT_N.n428 VOUT_N.n427 0.186204
R1271 VOUT_N.n437 VOUT_N.n436 0.186204
R1272 VOUT_N.n446 VOUT_N.n445 0.186204
R1273 VOUT_N.n472 VOUT_N.n471 0.186204
R1274 VOUT_N.n481 VOUT_N.n480 0.186204
R1275 VOUT_N.n490 VOUT_N.n489 0.186204
R1276 VOUT_N.n499 VOUT_N.n498 0.186204
R1277 VOUT_N.n599 VOUT_N.n598 0.186204
R1278 VOUT_N.n594 VOUT_N.n593 0.186204
R1279 VOUT_N.n585 VOUT_N.n584 0.186204
R1280 VOUT_N.n581 VOUT_N.n580 0.186204
R1281 VOUT_N.n563 VOUT_N.n562 0.186204
R1282 VOUT_N.n558 VOUT_N.n557 0.186204
R1283 VOUT_N.n23 VOUT_N.n22 0.186204
R1284 VOUT_N.n1712 VOUT_N.n1711 0.186204
R1285 VOUT_N.n1703 VOUT_N.n1702 0.186204
R1286 VOUT_N.n1798 VOUT_N.n1797 0.186204
R1287 VOUT_N.n1793 VOUT_N.n1792 0.186204
R1288 VOUT_N.n1752 VOUT_N.n1751 0.186204
R1289 VOUT_N.n2228 VOUT_N.n2227 0.186204
R1290 VOUT_N.n2224 VOUT_N.n2223 0.186204
R1291 VOUT_N.n2215 VOUT_N.n2214 0.186204
R1292 VOUT_N.n2210 VOUT_N.n2209 0.186204
R1293 VOUT_N.n2035 VOUT_N.n2034 0.186204
R1294 VOUT_N.n2031 VOUT_N.n2030 0.186204
R1295 VOUT_N.n1148 VOUT_N.n1147 0.176697
R1296 VOUT_N.n1487 VOUT_N.n1486 0.176697
R1297 VOUT_N.n807 VOUT_N.n806 0.176697
R1298 VOUT_N.n356 VOUT_N.n355 0.176697
R1299 VOUT_N.n1200 VOUT_N.n1199 0.166556
R1300 VOUT_N.n1560 VOUT_N.n1559 0.166556
R1301 VOUT_N.n853 VOUT_N.n852 0.166556
R1302 VOUT_N.n406 VOUT_N.n405 0.166556
R1303 VOUT_N.n1246 VOUT_N.n1245 0.162754
R1304 VOUT_N.n1629 VOUT_N.n1628 0.162754
R1305 VOUT_N.n897 VOUT_N.n896 0.162754
R1306 VOUT_N.n458 VOUT_N.n457 0.162754
R1307 VOUT_N.n1626 VOUT_N.n1625 0.145641
R1308 VOUT_N.n1557 VOUT_N.n1556 0.145641
R1309 VOUT_N.n1574 VOUT_N.n1573 0.145641
R1310 VOUT_N.n1481 VOUT_N.n1480 0.145641
R1311 VOUT_N.n1497 VOUT_N.n1496 0.145641
R1312 VOUT_N.n1302 VOUT_N.n1301 0.145641
R1313 VOUT_N.n1910 VOUT_N.n1909 0.106363
R1314 VOUT_N.n2008 VOUT_N.n2007 0.106345
R1315 VOUT_N.n1886 VOUT_N.n1885 0.106345
R1316 VOUT_N.n2203 VOUT_N.n2202 0.106345
R1317 VOUT_N.n2126 VOUT_N.n2125 0.106345
R1318 VOUT_N.n1820 VOUT_N.n1818 0.106345
R1319 VOUT_N.n1760 VOUT_N.n1759 0.106345
R1320 VOUT_N.n1682 VOUT_N.n1681 0.106345
R1321 VOUT_N.n169 VOUT_N.n105 0.105505
R1322 VOUT_N.n2192 VOUT_N.n2187 0.0992756
R1323 VOUT_N.n1982 VOUT_N.n1977 0.0992756
R1324 VOUT_N.n12 VOUT_N.n7 0.0992756
R1325 VOUT_N.n1721 VOUT_N.n1716 0.0992756
R1326 VOUT_N.n1741 VOUT_N.n1736 0.0992756
R1327 VOUT_N VOUT_N.n2245 0.0835282
R1328 VOUT_N.n1913 VOUT_N.n1912 0.0832399
R1329 VOUT_N.n1699 VOUT_N.n1694 0.0832399
R1330 VOUT_N.n2181 VOUT_N.n2180 0.0831446
R1331 VOUT_N.n1906 VOUT_N.n1899 0.0824117
R1332 VOUT_N.n1773 VOUT_N.n1766 0.0824117
R1333 VOUT_N.n2023 VOUT_N.n2020 0.0824117
R1334 VOUT_N.n328 VOUT_N.n324 0.0823987
R1335 VOUT_N.n317 VOUT_N.n312 0.0823987
R1336 VOUT_N.n549 VOUT_N.n544 0.0823987
R1337 VOUT_N.n2110 VOUT_N.n2105 0.0823987
R1338 VOUT_N.n1867 VOUT_N.n1862 0.0823987
R1339 VOUT_N.n1941 VOUT_N.n1936 0.0823987
R1340 VOUT_N.n2148 VOUT_N.n2143 0.0823987
R1341 VOUT_N.n2071 VOUT_N.n2064 0.0823987
R1342 VOUT_N.n2140 VOUT_N.n2136 0.0823987
R1343 VOUT_N.n534 VOUT_N.n531 0.0823987
R1344 VOUT_N.n524 VOUT_N.n520 0.0823987
R1345 VOUT_N.n515 VOUT_N.n510 0.0823987
R1346 VOUT_N.n784 VOUT_N.n779 0.0823987
R1347 VOUT_N.n772 VOUT_N.n767 0.0823987
R1348 VOUT_N.n760 VOUT_N.n755 0.0823987
R1349 VOUT_N.n748 VOUT_N.n743 0.0823987
R1350 VOUT_N.n736 VOUT_N.n731 0.0823987
R1351 VOUT_N.n724 VOUT_N.n719 0.0823987
R1352 VOUT_N.n628 VOUT_N.n623 0.0823987
R1353 VOUT_N.n640 VOUT_N.n635 0.0823987
R1354 VOUT_N.n652 VOUT_N.n647 0.0823987
R1355 VOUT_N.n664 VOUT_N.n659 0.0823987
R1356 VOUT_N.n676 VOUT_N.n671 0.0823987
R1357 VOUT_N.n688 VOUT_N.n683 0.0823987
R1358 VOUT_N.n700 VOUT_N.n695 0.0823987
R1359 VOUT_N.n712 VOUT_N.n707 0.0823987
R1360 VOUT_N.n1456 VOUT_N.n1452 0.0823987
R1361 VOUT_N.n1445 VOUT_N.n1440 0.0823987
R1362 VOUT_N.n1435 VOUT_N.n1431 0.0823987
R1363 VOUT_N.n1424 VOUT_N.n1419 0.0823987
R1364 VOUT_N.n1414 VOUT_N.n1410 0.0823987
R1365 VOUT_N.n1403 VOUT_N.n1398 0.0823987
R1366 VOUT_N.n1393 VOUT_N.n1389 0.0823987
R1367 VOUT_N.n1382 VOUT_N.n1377 0.0823987
R1368 VOUT_N.n1372 VOUT_N.n1368 0.0823987
R1369 VOUT_N.n1361 VOUT_N.n1356 0.0823987
R1370 VOUT_N.n1314 VOUT_N.n1309 0.0823987
R1371 VOUT_N.n1325 VOUT_N.n1321 0.0823987
R1372 VOUT_N.n1335 VOUT_N.n1330 0.0823987
R1373 VOUT_N.n1346 VOUT_N.n1342 0.0823987
R1374 VOUT_N.n1119 VOUT_N.n1114 0.0823987
R1375 VOUT_N.n1107 VOUT_N.n1102 0.0823987
R1376 VOUT_N.n1095 VOUT_N.n1090 0.0823987
R1377 VOUT_N.n1083 VOUT_N.n1078 0.0823987
R1378 VOUT_N.n1071 VOUT_N.n1066 0.0823987
R1379 VOUT_N.n1059 VOUT_N.n1054 0.0823987
R1380 VOUT_N.n1047 VOUT_N.n1042 0.0823987
R1381 VOUT_N.n1035 VOUT_N.n1030 0.0823987
R1382 VOUT_N.n1023 VOUT_N.n1018 0.0823987
R1383 VOUT_N.n1011 VOUT_N.n1006 0.0823987
R1384 VOUT_N.n957 VOUT_N.n952 0.0823987
R1385 VOUT_N.n969 VOUT_N.n964 0.0823987
R1386 VOUT_N.n981 VOUT_N.n976 0.0823987
R1387 VOUT_N.n993 VOUT_N.n988 0.0823987
R1388 VOUT_N.n307 VOUT_N.n303 0.0823987
R1389 VOUT_N.n296 VOUT_N.n291 0.0823987
R1390 VOUT_N.n286 VOUT_N.n282 0.0823987
R1391 VOUT_N.n275 VOUT_N.n270 0.0823987
R1392 VOUT_N.n265 VOUT_N.n261 0.0823987
R1393 VOUT_N.n254 VOUT_N.n249 0.0823987
R1394 VOUT_N.n244 VOUT_N.n240 0.0823987
R1395 VOUT_N.n233 VOUT_N.n228 0.0823987
R1396 VOUT_N.n223 VOUT_N.n219 0.0823987
R1397 VOUT_N.n212 VOUT_N.n207 0.0823987
R1398 VOUT_N.n202 VOUT_N.n198 0.0823987
R1399 VOUT_N.n191 VOUT_N.n186 0.0823987
R1400 VOUT_N.n1781 VOUT_N.n1774 0.0823987
R1401 VOUT_N.n1825 VOUT_N.n1821 0.0823987
R1402 VOUT_N.n1835 VOUT_N.n1832 0.0823987
R1403 VOUT_N.n1846 VOUT_N.n1841 0.0823987
R1404 VOUT_N.n2013 VOUT_N.n2009 0.0823987
R1405 VOUT_N.n1698 VOUT_N.n1697 0.0817926
R1406 VOUT_N.n1904 VOUT_N.n1903 0.0748144
R1407 VOUT_N.n2069 VOUT_N.n2068 0.0748144
R1408 VOUT_N.n1779 VOUT_N.n1778 0.0748144
R1409 VOUT_N.n1787 VOUT_N.n1786 0.0748144
R1410 VOUT_N.n1771 VOUT_N.n1770 0.0748144
R1411 VOUT_N.n2063 VOUT_N.n2059 0.0712285
R1412 VOUT_N.n1898 VOUT_N.n1893 0.0712285
R1413 VOUT_N.n2080 VOUT_N.n2075 0.0712285
R1414 VOUT_N.n1948 VOUT_N.n1944 0.0712285
R1415 VOUT_N.n2104 VOUT_N.n2099 0.0712285
R1416 VOUT_N.n1873 VOUT_N.n1868 0.0712285
R1417 VOUT_N.n1005 VOUT_N.n1000 0.0712285
R1418 VOUT_N.n987 VOUT_N.n982 0.0712285
R1419 VOUT_N.n975 VOUT_N.n970 0.0712285
R1420 VOUT_N.n963 VOUT_N.n958 0.0712285
R1421 VOUT_N.n951 VOUT_N.n946 0.0712285
R1422 VOUT_N.n1017 VOUT_N.n1012 0.0712285
R1423 VOUT_N.n1029 VOUT_N.n1024 0.0712285
R1424 VOUT_N.n1041 VOUT_N.n1036 0.0712285
R1425 VOUT_N.n1053 VOUT_N.n1048 0.0712285
R1426 VOUT_N.n1065 VOUT_N.n1060 0.0712285
R1427 VOUT_N.n1077 VOUT_N.n1072 0.0712285
R1428 VOUT_N.n1089 VOUT_N.n1084 0.0712285
R1429 VOUT_N.n1101 VOUT_N.n1096 0.0712285
R1430 VOUT_N.n1113 VOUT_N.n1108 0.0712285
R1431 VOUT_N.n1355 VOUT_N.n1352 0.0712285
R1432 VOUT_N.n1341 VOUT_N.n1336 0.0712285
R1433 VOUT_N.n1329 VOUT_N.n1326 0.0712285
R1434 VOUT_N.n1320 VOUT_N.n1315 0.0712285
R1435 VOUT_N.n1308 VOUT_N.n1305 0.0712285
R1436 VOUT_N.n1367 VOUT_N.n1362 0.0712285
R1437 VOUT_N.n1376 VOUT_N.n1373 0.0712285
R1438 VOUT_N.n1388 VOUT_N.n1383 0.0712285
R1439 VOUT_N.n1397 VOUT_N.n1394 0.0712285
R1440 VOUT_N.n1409 VOUT_N.n1404 0.0712285
R1441 VOUT_N.n1418 VOUT_N.n1415 0.0712285
R1442 VOUT_N.n1430 VOUT_N.n1425 0.0712285
R1443 VOUT_N.n1439 VOUT_N.n1436 0.0712285
R1444 VOUT_N.n1451 VOUT_N.n1446 0.0712285
R1445 VOUT_N.n718 VOUT_N.n713 0.0712285
R1446 VOUT_N.n706 VOUT_N.n701 0.0712285
R1447 VOUT_N.n694 VOUT_N.n689 0.0712285
R1448 VOUT_N.n682 VOUT_N.n677 0.0712285
R1449 VOUT_N.n670 VOUT_N.n665 0.0712285
R1450 VOUT_N.n658 VOUT_N.n653 0.0712285
R1451 VOUT_N.n646 VOUT_N.n641 0.0712285
R1452 VOUT_N.n634 VOUT_N.n629 0.0712285
R1453 VOUT_N.n622 VOUT_N.n617 0.0712285
R1454 VOUT_N.n730 VOUT_N.n725 0.0712285
R1455 VOUT_N.n742 VOUT_N.n737 0.0712285
R1456 VOUT_N.n754 VOUT_N.n749 0.0712285
R1457 VOUT_N.n766 VOUT_N.n761 0.0712285
R1458 VOUT_N.n778 VOUT_N.n773 0.0712285
R1459 VOUT_N.n185 VOUT_N.n182 0.0712285
R1460 VOUT_N.n197 VOUT_N.n192 0.0712285
R1461 VOUT_N.n206 VOUT_N.n203 0.0712285
R1462 VOUT_N.n218 VOUT_N.n213 0.0712285
R1463 VOUT_N.n227 VOUT_N.n224 0.0712285
R1464 VOUT_N.n239 VOUT_N.n234 0.0712285
R1465 VOUT_N.n248 VOUT_N.n245 0.0712285
R1466 VOUT_N.n260 VOUT_N.n255 0.0712285
R1467 VOUT_N.n269 VOUT_N.n266 0.0712285
R1468 VOUT_N.n281 VOUT_N.n276 0.0712285
R1469 VOUT_N.n290 VOUT_N.n287 0.0712285
R1470 VOUT_N.n302 VOUT_N.n297 0.0712285
R1471 VOUT_N.n311 VOUT_N.n308 0.0712285
R1472 VOUT_N.n509 VOUT_N.n505 0.0712285
R1473 VOUT_N.n519 VOUT_N.n516 0.0712285
R1474 VOUT_N.n530 VOUT_N.n525 0.0712285
R1475 VOUT_N.n543 VOUT_N.n539 0.0712285
R1476 VOUT_N.n553 VOUT_N.n550 0.0712285
R1477 VOUT_N.n323 VOUT_N.n318 0.0712285
R1478 VOUT_N.n2019 VOUT_N.n2014 0.0712285
R1479 VOUT_N.n1850 VOUT_N.n1847 0.0712285
R1480 VOUT_N.n1840 VOUT_N.n1836 0.0712285
R1481 VOUT_N.n1831 VOUT_N.n1826 0.0712285
R1482 VOUT_N.n1967 VOUT_N.n1966 0.0709833
R1483 VOUT_N.n147 VOUT_N.n146 0.0707439
R1484 VOUT_N.n68 VOUT_N.n67 0.0707439
R1485 VOUT_N.n1988 VOUT_N.n1987 0.0623855
R1486 VOUT_N.n1987 VOUT_N.n1986 0.0623855
R1487 VOUT_N.n18 VOUT_N.n17 0.0623855
R1488 VOUT_N.n17 VOUT_N.n16 0.0623855
R1489 VOUT_N.n1788 VOUT_N.n1783 0.0623855
R1490 VOUT_N.n1783 VOUT_N.n1782 0.0623855
R1491 VOUT_N.n1747 VOUT_N.n1746 0.0623855
R1492 VOUT_N.n1746 VOUT_N.n1745 0.0623855
R1493 VOUT_N.n1967 VOUT_N.n1962 0.0536862
R1494 VOUT_N.n1898 VOUT_N.n1897 0.0534597
R1495 VOUT_N.n2080 VOUT_N.n2079 0.0534597
R1496 VOUT_N.n2063 VOUT_N.n2062 0.0534597
R1497 VOUT_N.n1948 VOUT_N.n1947 0.0534597
R1498 VOUT_N.n1873 VOUT_N.n1872 0.0534597
R1499 VOUT_N.n2104 VOUT_N.n2103 0.0534597
R1500 VOUT_N.n951 VOUT_N.n950 0.0534597
R1501 VOUT_N.n963 VOUT_N.n962 0.0534597
R1502 VOUT_N.n975 VOUT_N.n974 0.0534597
R1503 VOUT_N.n987 VOUT_N.n986 0.0534597
R1504 VOUT_N.n1113 VOUT_N.n1112 0.0534597
R1505 VOUT_N.n1101 VOUT_N.n1100 0.0534597
R1506 VOUT_N.n1089 VOUT_N.n1088 0.0534597
R1507 VOUT_N.n1077 VOUT_N.n1076 0.0534597
R1508 VOUT_N.n1065 VOUT_N.n1064 0.0534597
R1509 VOUT_N.n1053 VOUT_N.n1052 0.0534597
R1510 VOUT_N.n1041 VOUT_N.n1040 0.0534597
R1511 VOUT_N.n1029 VOUT_N.n1028 0.0534597
R1512 VOUT_N.n1017 VOUT_N.n1016 0.0534597
R1513 VOUT_N.n1005 VOUT_N.n1004 0.0534597
R1514 VOUT_N.n1308 VOUT_N.n1307 0.0534597
R1515 VOUT_N.n1320 VOUT_N.n1319 0.0534597
R1516 VOUT_N.n1329 VOUT_N.n1328 0.0534597
R1517 VOUT_N.n1341 VOUT_N.n1340 0.0534597
R1518 VOUT_N.n1451 VOUT_N.n1450 0.0534597
R1519 VOUT_N.n1439 VOUT_N.n1438 0.0534597
R1520 VOUT_N.n1430 VOUT_N.n1429 0.0534597
R1521 VOUT_N.n1418 VOUT_N.n1417 0.0534597
R1522 VOUT_N.n1409 VOUT_N.n1408 0.0534597
R1523 VOUT_N.n1397 VOUT_N.n1396 0.0534597
R1524 VOUT_N.n1388 VOUT_N.n1387 0.0534597
R1525 VOUT_N.n1376 VOUT_N.n1375 0.0534597
R1526 VOUT_N.n1367 VOUT_N.n1366 0.0534597
R1527 VOUT_N.n1355 VOUT_N.n1354 0.0534597
R1528 VOUT_N.n622 VOUT_N.n621 0.0534597
R1529 VOUT_N.n634 VOUT_N.n633 0.0534597
R1530 VOUT_N.n646 VOUT_N.n645 0.0534597
R1531 VOUT_N.n658 VOUT_N.n657 0.0534597
R1532 VOUT_N.n670 VOUT_N.n669 0.0534597
R1533 VOUT_N.n682 VOUT_N.n681 0.0534597
R1534 VOUT_N.n694 VOUT_N.n693 0.0534597
R1535 VOUT_N.n706 VOUT_N.n705 0.0534597
R1536 VOUT_N.n778 VOUT_N.n777 0.0534597
R1537 VOUT_N.n766 VOUT_N.n765 0.0534597
R1538 VOUT_N.n754 VOUT_N.n753 0.0534597
R1539 VOUT_N.n742 VOUT_N.n741 0.0534597
R1540 VOUT_N.n730 VOUT_N.n729 0.0534597
R1541 VOUT_N.n718 VOUT_N.n717 0.0534597
R1542 VOUT_N.n553 VOUT_N.n552 0.0534597
R1543 VOUT_N.n543 VOUT_N.n542 0.0534597
R1544 VOUT_N.n530 VOUT_N.n529 0.0534597
R1545 VOUT_N.n519 VOUT_N.n518 0.0534597
R1546 VOUT_N.n509 VOUT_N.n508 0.0534597
R1547 VOUT_N.n323 VOUT_N.n322 0.0534597
R1548 VOUT_N.n311 VOUT_N.n310 0.0534597
R1549 VOUT_N.n302 VOUT_N.n301 0.0534597
R1550 VOUT_N.n290 VOUT_N.n289 0.0534597
R1551 VOUT_N.n281 VOUT_N.n280 0.0534597
R1552 VOUT_N.n269 VOUT_N.n268 0.0534597
R1553 VOUT_N.n260 VOUT_N.n259 0.0534597
R1554 VOUT_N.n248 VOUT_N.n247 0.0534597
R1555 VOUT_N.n239 VOUT_N.n238 0.0534597
R1556 VOUT_N.n227 VOUT_N.n226 0.0534597
R1557 VOUT_N.n218 VOUT_N.n217 0.0534597
R1558 VOUT_N.n206 VOUT_N.n205 0.0534597
R1559 VOUT_N.n197 VOUT_N.n196 0.0534597
R1560 VOUT_N.n185 VOUT_N.n184 0.0534597
R1561 VOUT_N.n1831 VOUT_N.n1830 0.0534597
R1562 VOUT_N.n1840 VOUT_N.n1839 0.0534597
R1563 VOUT_N.n1850 VOUT_N.n1849 0.0534597
R1564 VOUT_N.n2019 VOUT_N.n2018 0.0534597
R1565 VOUT_N.n2180 VOUT_N.n2179 0.0420655
R1566 VOUT_N.n1912 VOUT_N.n1911 0.0419676
R1567 VOUT_N.n1694 VOUT_N.n1693 0.0419676
R1568 VOUT_N.n2071 VOUT_N.n2070 0.0415773
R1569 VOUT_N.n1941 VOUT_N.n1940 0.0415773
R1570 VOUT_N.n2148 VOUT_N.n2147 0.0415773
R1571 VOUT_N.n2140 VOUT_N.n2139 0.0415773
R1572 VOUT_N.n1867 VOUT_N.n1866 0.0415773
R1573 VOUT_N.n2110 VOUT_N.n2109 0.0415773
R1574 VOUT_N.n993 VOUT_N.n992 0.0415773
R1575 VOUT_N.n981 VOUT_N.n980 0.0415773
R1576 VOUT_N.n969 VOUT_N.n968 0.0415773
R1577 VOUT_N.n957 VOUT_N.n956 0.0415773
R1578 VOUT_N.n1011 VOUT_N.n1010 0.0415773
R1579 VOUT_N.n1023 VOUT_N.n1022 0.0415773
R1580 VOUT_N.n1035 VOUT_N.n1034 0.0415773
R1581 VOUT_N.n1047 VOUT_N.n1046 0.0415773
R1582 VOUT_N.n1059 VOUT_N.n1058 0.0415773
R1583 VOUT_N.n1071 VOUT_N.n1070 0.0415773
R1584 VOUT_N.n1083 VOUT_N.n1082 0.0415773
R1585 VOUT_N.n1095 VOUT_N.n1094 0.0415773
R1586 VOUT_N.n1107 VOUT_N.n1106 0.0415773
R1587 VOUT_N.n1119 VOUT_N.n1118 0.0415773
R1588 VOUT_N.n1346 VOUT_N.n1345 0.0415773
R1589 VOUT_N.n1335 VOUT_N.n1334 0.0415773
R1590 VOUT_N.n1325 VOUT_N.n1324 0.0415773
R1591 VOUT_N.n1314 VOUT_N.n1313 0.0415773
R1592 VOUT_N.n1361 VOUT_N.n1360 0.0415773
R1593 VOUT_N.n1372 VOUT_N.n1371 0.0415773
R1594 VOUT_N.n1382 VOUT_N.n1381 0.0415773
R1595 VOUT_N.n1393 VOUT_N.n1392 0.0415773
R1596 VOUT_N.n1403 VOUT_N.n1402 0.0415773
R1597 VOUT_N.n1414 VOUT_N.n1413 0.0415773
R1598 VOUT_N.n1424 VOUT_N.n1423 0.0415773
R1599 VOUT_N.n1435 VOUT_N.n1434 0.0415773
R1600 VOUT_N.n1445 VOUT_N.n1444 0.0415773
R1601 VOUT_N.n1456 VOUT_N.n1455 0.0415773
R1602 VOUT_N.n712 VOUT_N.n711 0.0415773
R1603 VOUT_N.n700 VOUT_N.n699 0.0415773
R1604 VOUT_N.n688 VOUT_N.n687 0.0415773
R1605 VOUT_N.n676 VOUT_N.n675 0.0415773
R1606 VOUT_N.n664 VOUT_N.n663 0.0415773
R1607 VOUT_N.n652 VOUT_N.n651 0.0415773
R1608 VOUT_N.n640 VOUT_N.n639 0.0415773
R1609 VOUT_N.n628 VOUT_N.n627 0.0415773
R1610 VOUT_N.n724 VOUT_N.n723 0.0415773
R1611 VOUT_N.n736 VOUT_N.n735 0.0415773
R1612 VOUT_N.n748 VOUT_N.n747 0.0415773
R1613 VOUT_N.n760 VOUT_N.n759 0.0415773
R1614 VOUT_N.n772 VOUT_N.n771 0.0415773
R1615 VOUT_N.n784 VOUT_N.n783 0.0415773
R1616 VOUT_N.n191 VOUT_N.n190 0.0415773
R1617 VOUT_N.n202 VOUT_N.n201 0.0415773
R1618 VOUT_N.n212 VOUT_N.n211 0.0415773
R1619 VOUT_N.n223 VOUT_N.n222 0.0415773
R1620 VOUT_N.n233 VOUT_N.n232 0.0415773
R1621 VOUT_N.n244 VOUT_N.n243 0.0415773
R1622 VOUT_N.n254 VOUT_N.n253 0.0415773
R1623 VOUT_N.n265 VOUT_N.n264 0.0415773
R1624 VOUT_N.n275 VOUT_N.n274 0.0415773
R1625 VOUT_N.n286 VOUT_N.n285 0.0415773
R1626 VOUT_N.n296 VOUT_N.n295 0.0415773
R1627 VOUT_N.n307 VOUT_N.n306 0.0415773
R1628 VOUT_N.n515 VOUT_N.n514 0.0415773
R1629 VOUT_N.n524 VOUT_N.n523 0.0415773
R1630 VOUT_N.n534 VOUT_N.n533 0.0415773
R1631 VOUT_N.n549 VOUT_N.n548 0.0415773
R1632 VOUT_N.n317 VOUT_N.n316 0.0415773
R1633 VOUT_N.n328 VOUT_N.n327 0.0415773
R1634 VOUT_N.n1781 VOUT_N.n1780 0.0415773
R1635 VOUT_N.n2013 VOUT_N.n2012 0.0415773
R1636 VOUT_N.n1846 VOUT_N.n1845 0.0415773
R1637 VOUT_N.n1835 VOUT_N.n1834 0.0415773
R1638 VOUT_N.n1825 VOUT_N.n1824 0.0415773
R1639 VOUT_N.n1906 VOUT_N.n1905 0.0415636
R1640 VOUT_N.n1773 VOUT_N.n1772 0.0415636
R1641 VOUT_N.n2023 VOUT_N.n2022 0.0415636
R1642 VOUT_N.n1946 VOUT_N.n1945 0.0383947
R1643 VOUT_N.n1961 VOUT_N.n1960 0.0383947
R1644 VOUT_N.n2135 VOUT_N.n2134 0.0383947
R1645 VOUT_N.n2151 VOUT_N.n2150 0.0383947
R1646 VOUT_N.n1697 VOUT_N.n1696 0.0383947
R1647 VOUT_N.n1715 VOUT_N.n1714 0.0383947
R1648 VOUT_N.n2095 VOUT_N.n2092 0.0334577
R1649 VOUT_N.n1927 VOUT_N.n1926 0.0334577
R1650 VOUT_N.n2172 VOUT_N.n2171 0.0334577
R1651 VOUT_N.n1147 VOUT_N.n1139 0.0334577
R1652 VOUT_N.n1158 VOUT_N.n1150 0.0334577
R1653 VOUT_N.n1299 VOUT_N.n1297 0.0334577
R1654 VOUT_N.n1299 VOUT_N.n1298 0.0334577
R1655 VOUT_N.n1559 VOUT_N.n1540 0.0334577
R1656 VOUT_N.n1628 VOUT_N.n1620 0.0334577
R1657 VOUT_N.n1632 VOUT_N.n1631 0.0334577
R1658 VOUT_N.n1671 VOUT_N.n1669 0.0334577
R1659 VOUT_N.n1671 VOUT_N.n1670 0.0334577
R1660 VOUT_N.n854 VOUT_N.n853 0.0334577
R1661 VOUT_N.n855 VOUT_N.n854 0.0334577
R1662 VOUT_N.n939 VOUT_N.n938 0.0334577
R1663 VOUT_N.n413 VOUT_N.n410 0.0334577
R1664 VOUT_N.n457 VOUT_N.n454 0.0334577
R1665 VOUT_N.n575 VOUT_N.n574 0.0334577
R1666 VOUT_N.n1727 VOUT_N.n1726 0.0334577
R1667 VOUT_N.n1692 VOUT_N.n1691 0.0319869
R1668 VOUT_N.n67 VOUT_N.t0 0.0306947
R1669 VOUT_N.n146 VOUT_N.t1 0.0285465
R1670 VOUT_N.n1982 VOUT_N.n1981 0.0254881
R1671 VOUT_N.n2192 VOUT_N.n2191 0.0254881
R1672 VOUT_N.n12 VOUT_N.n11 0.0254881
R1673 VOUT_N.n1721 VOUT_N.n1720 0.0254881
R1674 VOUT_N.n1741 VOUT_N.n1740 0.0254881
R1675 VOUT_N.n1931 VOUT_N.n1930 0.0235313
R1676 VOUT_N.n1198 VOUT_N.n1197 0.0235313
R1677 VOUT_N.n1563 VOUT_N.n1562 0.0235313
R1678 VOUT_N.n805 VOUT_N.n804 0.0235313
R1679 VOUT_N.n998 VOUT_N.n997 0.0235313
R1680 VOUT_N.n1490 VOUT_N.n1489 0.0235313
R1681 VOUT_N.n349 VOUT_N.n348 0.0235313
R1682 VOUT_N.n1 VOUT_N.n0 0.0235313
R1683 VOUT_N.n405 VOUT_N.n404 0.0228651
R1684 VOUT_N.n2050 VOUT_N.n2048 0.0228651
R1685 VOUT_N.n2007 VOUT_N.n2006 0.0228651
R1686 VOUT_N.n2002 VOUT_N.n2001 0.0228651
R1687 VOUT_N.n2173 VOUT_N.n2133 0.0228651
R1688 VOUT_N.n2202 VOUT_N.n2201 0.0228651
R1689 VOUT_N.n2133 VOUT_N.n2132 0.0228651
R1690 VOUT_N.n2097 VOUT_N.n2096 0.0228651
R1691 VOUT_N.n1250 VOUT_N.n1249 0.0228651
R1692 VOUT_N.n1249 VOUT_N.n1248 0.0228651
R1693 VOUT_N.n1553 VOUT_N.n1552 0.0228651
R1694 VOUT_N.n1202 VOUT_N.n1201 0.0228651
R1695 VOUT_N.n1570 VOUT_N.n1569 0.0228651
R1696 VOUT_N.n1576 VOUT_N.n1575 0.0228651
R1697 VOUT_N.n1349 VOUT_N.n1347 0.0228651
R1698 VOUT_N.n1631 VOUT_N.n1630 0.0228651
R1699 VOUT_N.n1477 VOUT_N.n1476 0.0228651
R1700 VOUT_N.n1483 VOUT_N.n1482 0.0228651
R1701 VOUT_N.n1566 VOUT_N.n1565 0.0228651
R1702 VOUT_N.n895 VOUT_N.n894 0.0228651
R1703 VOUT_N.n996 VOUT_N.n995 0.0228651
R1704 VOUT_N.n1255 VOUT_N.n1254 0.0228651
R1705 VOUT_N.n900 VOUT_N.n899 0.0228651
R1706 VOUT_N.n893 VOUT_N.n892 0.0228651
R1707 VOUT_N.n851 VOUT_N.n850 0.0228651
R1708 VOUT_N.n1567 VOUT_N.n1566 0.0228651
R1709 VOUT_N.n1141 VOUT_N.n1140 0.0228651
R1710 VOUT_N.n1548 VOUT_N.n1547 0.0228651
R1711 VOUT_N.n809 VOUT_N.n808 0.0228651
R1712 VOUT_N.n1492 VOUT_N.n1491 0.0228651
R1713 VOUT_N.n1152 VOUT_N.n1151 0.0228651
R1714 VOUT_N.n1546 VOUT_N.n1545 0.0228651
R1715 VOUT_N.n352 VOUT_N.n351 0.0228651
R1716 VOUT_N.n1543 VOUT_N.n1542 0.0228651
R1717 VOUT_N.n403 VOUT_N.n402 0.0228651
R1718 VOUT_N.n1731 VOUT_N.n1730 0.0228651
R1719 VOUT_N.n1813 VOUT_N.n1812 0.0228651
R1720 VOUT_N.n1761 VOUT_N.n1760 0.0228651
R1721 VOUT_N.n1815 VOUT_N.n1814 0.0228651
R1722 VOUT_N.n31 VOUT_N.n30 0.0228651
R1723 VOUT_N.n2203 VOUT_N.n2054 0.0228651
R1724 VOUT_N.n2204 VOUT_N.n2051 0.0228651
R1725 VOUT_N.n1304 VOUT_N.n1303 0.0228651
R1726 VOUT_N.n945 VOUT_N.n944 0.0228651
R1727 VOUT_N.n941 VOUT_N.n939 0.0228651
R1728 VOUT_N.n1681 VOUT_N.n1680 0.0228651
R1729 VOUT_N.n610 VOUT_N.n609 0.0228651
R1730 VOUT_N.n615 VOUT_N.n614 0.0228651
R1731 VOUT_N.n1672 VOUT_N.n1304 0.0228651
R1732 VOUT_N.n1300 VOUT_N.n945 0.0228651
R1733 VOUT_N.n180 VOUT_N.n179 0.0228651
R1734 VOUT_N.n173 VOUT_N.n172 0.0228651
R1735 VOUT_N.n3 VOUT_N.n2 0.0228651
R1736 VOUT_N.n99 VOUT_N.n98 0.0195244
R1737 VOUT_N.n100 VOUT_N.n99 0.0195244
R1738 VOUT_N.n101 VOUT_N.n100 0.0195244
R1739 VOUT_N.n148 VOUT_N.n147 0.0195244
R1740 VOUT_N.n149 VOUT_N.n148 0.0195244
R1741 VOUT_N.n150 VOUT_N.n149 0.0195244
R1742 VOUT_N.n69 VOUT_N.n68 0.0195244
R1743 VOUT_N.n70 VOUT_N.n69 0.0195244
R1744 VOUT_N.n71 VOUT_N.n70 0.0195244
R1745 VOUT_N.n1927 VOUT_N.n1890 0.0179841
R1746 VOUT_N.n1929 VOUT_N.n1928 0.0179841
R1747 VOUT_N.n1885 VOUT_N.n1884 0.0179841
R1748 VOUT_N.n1861 VOUT_N.n1860 0.0179841
R1749 VOUT_N.n2128 VOUT_N.n2127 0.0179841
R1750 VOUT_N.n2130 VOUT_N.n2129 0.0179841
R1751 VOUT_N.n2200 VOUT_N.n2199 0.0179841
R1752 VOUT_N.n2095 VOUT_N.n2094 0.0179841
R1753 VOUT_N.n456 VOUT_N.n455 0.0179841
R1754 VOUT_N.n1556 VOUT_N.n1555 0.0179841
R1755 VOUT_N.n1625 VOUT_N.n1624 0.0179841
R1756 VOUT_N.n1245 VOUT_N.n1244 0.0179841
R1757 VOUT_N.n1623 VOUT_N.n1622 0.0179841
R1758 VOUT_N.n1578 VOUT_N.n1574 0.0179841
R1759 VOUT_N.n1627 VOUT_N.n1621 0.0179841
R1760 VOUT_N.n1558 VOUT_N.n1541 0.0179841
R1761 VOUT_N.n1480 VOUT_N.n1479 0.0179841
R1762 VOUT_N.n1138 VOUT_N.n1137 0.0179841
R1763 VOUT_N.n1144 VOUT_N.n1143 0.0179841
R1764 VOUT_N.n1252 VOUT_N.n1251 0.0179841
R1765 VOUT_N.n1551 VOUT_N.n1550 0.0179841
R1766 VOUT_N.n1496 VOUT_N.n1495 0.0179841
R1767 VOUT_N.n1498 VOUT_N.n1493 0.0179841
R1768 VOUT_N.n1149 VOUT_N.n1148 0.0179841
R1769 VOUT_N.n605 VOUT_N.n604 0.0179841
R1770 VOUT_N.n360 VOUT_N.n359 0.0179841
R1771 VOUT_N.n409 VOUT_N.n408 0.0179841
R1772 VOUT_N.n453 VOUT_N.n452 0.0179841
R1773 VOUT_N.n538 VOUT_N.n537 0.0179841
R1774 VOUT_N.n1858 VOUT_N.n1857 0.0179841
R1775 VOUT_N.n569 VOUT_N.n568 0.0179841
R1776 VOUT_N.n1856 VOUT_N.n1855 0.0179841
R1777 VOUT_N.n462 VOUT_N.n461 0.0179841
R1778 VOUT_N.n354 VOUT_N.n350 0.0179841
R1779 VOUT_N.n357 VOUT_N.n356 0.0179841
R1780 VOUT_N.n363 VOUT_N.n362 0.0179841
R1781 VOUT_N.n407 VOUT_N.n406 0.0179841
R1782 VOUT_N.n412 VOUT_N.n411 0.0179841
R1783 VOUT_N.n451 VOUT_N.n450 0.0179841
R1784 VOUT_N.n459 VOUT_N.n458 0.0179841
R1785 VOUT_N.n465 VOUT_N.n464 0.0179841
R1786 VOUT_N.n1758 VOUT_N.n1735 0.0179841
R1787 VOUT_N.n1811 VOUT_N.n1810 0.0179841
R1788 VOUT_N.n30 VOUT_N.n29 0.0179841
R1789 VOUT_N.n606 VOUT_N.n605 0.0179841
R1790 VOUT_N.n1728 VOUT_N.n1727 0.0179841
R1791 VOUT_N.n2239 VOUT_N.n2236 0.0179841
R1792 VOUT_N.n2047 VOUT_N.n2043 0.0179841
R1793 VOUT_N.n2045 VOUT_N.n2044 0.0179841
R1794 VOUT_N.n611 VOUT_N.n181 0.0179841
R1795 VOUT_N.n1679 VOUT_N.n1678 0.0179841
R1796 VOUT_N.n171 VOUT_N.n34 0.0179841
R1797 VOUT_N.n1684 VOUT_N.n1683 0.0179841
R1798 VOUT_N.n2243 VOUT_N.n5 0.0179841
R1799 VOUT_N.n2046 VOUT_N.n2045 0.0177304
R1800 VOUT_N.n1857 VOUT_N.n1856 0.0177304
R1801 VOUT_N.n1999 VOUT_N.n1998 0.0177304
R1802 VOUT_N.n1928 VOUT_N.n1888 0.0177304
R1803 VOUT_N.n1890 VOUT_N.n1889 0.0177304
R1804 VOUT_N.n1853 VOUT_N.n1852 0.0177304
R1805 VOUT_N.n1884 VOUT_N.n1861 0.0177304
R1806 VOUT_N.n1860 VOUT_N.n1859 0.0177304
R1807 VOUT_N.n2094 VOUT_N.n2093 0.0177304
R1808 VOUT_N.n2199 VOUT_N.n2198 0.0177304
R1809 VOUT_N.n2129 VOUT_N.n2128 0.0177304
R1810 VOUT_N.n2127 VOUT_N.n2126 0.0177304
R1811 VOUT_N.n1555 VOUT_N.n1554 0.0177304
R1812 VOUT_N.n1244 VOUT_N.n1243 0.0177304
R1813 VOUT_N.n1624 VOUT_N.n1623 0.0177304
R1814 VOUT_N.n1578 VOUT_N.n1577 0.0177304
R1815 VOUT_N.n1558 VOUT_N.n1557 0.0177304
R1816 VOUT_N.n1627 VOUT_N.n1626 0.0177304
R1817 VOUT_N.n1619 VOUT_N.n1618 0.0177304
R1818 VOUT_N.n1539 VOUT_N.n1538 0.0177304
R1819 VOUT_N.n354 VOUT_N.n353 0.0177304
R1820 VOUT_N.n1139 VOUT_N.n1138 0.0177304
R1821 VOUT_N.n1479 VOUT_N.n1478 0.0177304
R1822 VOUT_N.n1146 VOUT_N.n1145 0.0177304
R1823 VOUT_N.n1143 VOUT_N.n1142 0.0177304
R1824 VOUT_N.n1550 VOUT_N.n1549 0.0177304
R1825 VOUT_N.n1253 VOUT_N.n1252 0.0177304
R1826 VOUT_N.n1150 VOUT_N.n1149 0.0177304
R1827 VOUT_N.n1498 VOUT_N.n1497 0.0177304
R1828 VOUT_N.n1495 VOUT_N.n1494 0.0177304
R1829 VOUT_N.n1157 VOUT_N.n1156 0.0177304
R1830 VOUT_N.n536 VOUT_N.n535 0.0177304
R1831 VOUT_N.n568 VOUT_N.n567 0.0177304
R1832 VOUT_N.n358 VOUT_N.n357 0.0177304
R1833 VOUT_N.n410 VOUT_N.n407 0.0177304
R1834 VOUT_N.n454 VOUT_N.n451 0.0177304
R1835 VOUT_N.n460 VOUT_N.n459 0.0177304
R1836 VOUT_N.n2238 VOUT_N.n2237 0.0177304
R1837 VOUT_N.n1758 VOUT_N.n1757 0.0177304
R1838 VOUT_N.n1810 VOUT_N.n1809 0.0177304
R1839 VOUT_N.n29 VOUT_N.n28 0.0177304
R1840 VOUT_N.n604 VOUT_N.n603 0.0177304
R1841 VOUT_N.n607 VOUT_N.n606 0.0177304
R1842 VOUT_N.n1729 VOUT_N.n1728 0.0177304
R1843 VOUT_N.n2236 VOUT_N.n2235 0.0177304
R1844 VOUT_N.n1820 VOUT_N.n1819 0.0177304
R1845 VOUT_N.n2043 VOUT_N.n2042 0.0177304
R1846 VOUT_N.n1678 VOUT_N.n1677 0.0177304
R1847 VOUT_N.n612 VOUT_N.n611 0.0177304
R1848 VOUT_N.n171 VOUT_N.n170 0.0177304
R1849 VOUT_N.n1683 VOUT_N.n1682 0.0177304
R1850 VOUT_N.n5 VOUT_N.n4 0.0177304
R1851 VOUT_N.n1260 VOUT_N.n1259 0.0174187
R1852 VOUT_N.n1259 VOUT_N.n1258 0.0174187
R1853 VOUT_N.n1351 VOUT_N.n1350 0.0174187
R1854 VOUT_N.n850 VOUT_N.n849 0.0174187
R1855 VOUT_N.n899 VOUT_N.n898 0.0174187
R1856 VOUT_N.n898 VOUT_N.n897 0.0174187
R1857 VOUT_N.n849 VOUT_N.n848 0.0174187
R1858 VOUT_N.n610 VOUT_N.n504 0.0174187
R1859 VOUT_N.n616 VOUT_N.n615 0.0174187
R1860 VOUT_N.n942 VOUT_N.n616 0.0174187
R1861 VOUT_N.n504 VOUT_N.n503 0.0174187
R1862 VOUT_N.n1975 VOUT_N.n1972 0.0173591
R1863 VOUT_N.n2197 VOUT_N.n2175 0.0173591
R1864 VOUT_N.n2004 VOUT_N.n2000 0.0173591
R1865 VOUT_N.n1971 VOUT_N.n1932 0.0173591
R1866 VOUT_N.n1887 VOUT_N.n1886 0.0173591
R1867 VOUT_N.n2005 VOUT_N.n2004 0.0173591
R1868 VOUT_N.n1976 VOUT_N.n1971 0.0173591
R1869 VOUT_N.n1975 VOUT_N.n1974 0.0173591
R1870 VOUT_N.n1888 VOUT_N.n1887 0.0173591
R1871 VOUT_N.n2124 VOUT_N.n2122 0.0173591
R1872 VOUT_N.n1854 VOUT_N.n1851 0.0173591
R1873 VOUT_N.n1854 VOUT_N.n1853 0.0173591
R1874 VOUT_N.n2125 VOUT_N.n2121 0.0173591
R1875 VOUT_N.n2121 VOUT_N.n2098 0.0173591
R1876 VOUT_N.n2124 VOUT_N.n2123 0.0173591
R1877 VOUT_N.n2197 VOUT_N.n2196 0.0173591
R1878 VOUT_N.n1196 VOUT_N.n1195 0.0173591
R1879 VOUT_N.n1203 VOUT_N.n1202 0.0173591
R1880 VOUT_N.n1242 VOUT_N.n1241 0.0173591
R1881 VOUT_N.n1258 VOUT_N.n1257 0.0173591
R1882 VOUT_N.n1197 VOUT_N.n1196 0.0173591
R1883 VOUT_N.n1257 VOUT_N.n1246 0.0173591
R1884 VOUT_N.n1243 VOUT_N.n1242 0.0173591
R1885 VOUT_N.n1573 VOUT_N.n1572 0.0173591
R1886 VOUT_N.n1572 VOUT_N.n1571 0.0173591
R1887 VOUT_N.n1204 VOUT_N.n1203 0.0173591
R1888 VOUT_N.n1476 VOUT_N.n1475 0.0173591
R1889 VOUT_N.n1489 VOUT_N.n1488 0.0173591
R1890 VOUT_N.n1540 VOUT_N.n1537 0.0173591
R1891 VOUT_N.n1562 VOUT_N.n1561 0.0173591
R1892 VOUT_N.n1620 VOUT_N.n1617 0.0173591
R1893 VOUT_N.n1561 VOUT_N.n1560 0.0173591
R1894 VOUT_N.n1537 VOUT_N.n1536 0.0173591
R1895 VOUT_N.n1617 VOUT_N.n1616 0.0173591
R1896 VOUT_N.n1485 VOUT_N.n1481 0.0173591
R1897 VOUT_N.n1485 VOUT_N.n1484 0.0173591
R1898 VOUT_N.n1475 VOUT_N.n1474 0.0173591
R1899 VOUT_N.n803 VOUT_N.n802 0.0173591
R1900 VOUT_N.n810 VOUT_N.n809 0.0173591
R1901 VOUT_N.n804 VOUT_N.n803 0.0173591
R1902 VOUT_N.n1155 VOUT_N.n1154 0.0173591
R1903 VOUT_N.n1154 VOUT_N.n1153 0.0173591
R1904 VOUT_N.n1488 VOUT_N.n1487 0.0173591
R1905 VOUT_N.n811 VOUT_N.n810 0.0173591
R1906 VOUT_N.n348 VOUT_N.n347 0.0173591
R1907 VOUT_N.n364 VOUT_N.n361 0.0173591
R1908 VOUT_N.n463 VOUT_N.n460 0.0173591
R1909 VOUT_N.n573 VOUT_N.n572 0.0173591
R1910 VOUT_N.n570 VOUT_N.n569 0.0173591
R1911 VOUT_N.n361 VOUT_N.n358 0.0173591
R1912 VOUT_N.n574 VOUT_N.n573 0.0173591
R1913 VOUT_N.n571 VOUT_N.n570 0.0173591
R1914 VOUT_N.n466 VOUT_N.n463 0.0173591
R1915 VOUT_N.n347 VOUT_N.n346 0.0173591
R1916 VOUT_N.n1676 VOUT_N.n1674 0.0173591
R1917 VOUT_N.n1808 VOUT_N.n1806 0.0173591
R1918 VOUT_N.n1804 VOUT_N.n1765 0.0173591
R1919 VOUT_N.n1818 VOUT_N.n1817 0.0173591
R1920 VOUT_N.n1805 VOUT_N.n1764 0.0173591
R1921 VOUT_N.n1759 VOUT_N.n1734 0.0173591
R1922 VOUT_N.n1734 VOUT_N.n1732 0.0173591
R1923 VOUT_N.n1764 VOUT_N.n1762 0.0173591
R1924 VOUT_N.n1804 VOUT_N.n1803 0.0173591
R1925 VOUT_N.n1808 VOUT_N.n1807 0.0173591
R1926 VOUT_N.n1817 VOUT_N.n1816 0.0173591
R1927 VOUT_N.n2241 VOUT_N.n1687 0.0173591
R1928 VOUT_N.n2234 VOUT_N.n2233 0.0173591
R1929 VOUT_N.n2042 VOUT_N.n2041 0.0173591
R1930 VOUT_N.n2235 VOUT_N.n2234 0.0173591
R1931 VOUT_N.n2041 VOUT_N.n2040 0.0173591
R1932 VOUT_N.n2242 VOUT_N.n1686 0.0173591
R1933 VOUT_N.n177 VOUT_N.n174 0.0173591
R1934 VOUT_N.n1686 VOUT_N.n1684 0.0173591
R1935 VOUT_N.n2241 VOUT_N.n2240 0.0173591
R1936 VOUT_N.n1676 VOUT_N.n1675 0.0173591
R1937 VOUT_N.n178 VOUT_N.n177 0.0173591
R1938 VOUT_N.n2244 VOUT_N.n1 0.0173591
R1939 VOUT_N.n2245 VOUT_N.n2244 0.0173591
R1940 VOUT_N.n1935 VOUT_N.n1934 0.0167343
R1941 VOUT_N.n2142 VOUT_N.n2141 0.0167343
R1942 VOUT_N.n1690 VOUT_N.n1689 0.0167343
R1943 VOUT_N.n1932 VOUT_N.n1931 0.0122638
R1944 VOUT_N.n2056 VOUT_N.n2055 0.0122638
R1945 VOUT_N.n1199 VOUT_N.n1198 0.0122638
R1946 VOUT_N.n1579 VOUT_N.n1563 0.0122638
R1947 VOUT_N.n806 VOUT_N.n805 0.0122638
R1948 VOUT_N.n997 VOUT_N.n996 0.0122638
R1949 VOUT_N.n1499 VOUT_N.n1490 0.0122638
R1950 VOUT_N.n355 VOUT_N.n349 0.0122638
R1951 VOUT_N.n33 VOUT_N.n6 0.0122638
R1952 VOUT_N.n1725 VOUT_N.n1688 0.0122638
R1953 VOUT_N.n404 VOUT_N.n403 0.0119325
R1954 VOUT_N.n2051 VOUT_N.n2050 0.0119325
R1955 VOUT_N.n176 VOUT_N.n175 0.0119325
R1956 VOUT_N.n1970 VOUT_N.n1933 0.0119325
R1957 VOUT_N.n2003 VOUT_N.n2002 0.0119325
R1958 VOUT_N.n2006 VOUT_N.n2005 0.0119325
R1959 VOUT_N.n2120 VOUT_N.n2119 0.0119325
R1960 VOUT_N.n2053 VOUT_N.n2052 0.0119325
R1961 VOUT_N.n2054 VOUT_N.n2053 0.0119325
R1962 VOUT_N.n2201 VOUT_N.n2200 0.0119325
R1963 VOUT_N.n2174 VOUT_N.n2173 0.0119325
R1964 VOUT_N.n2132 VOUT_N.n2131 0.0119325
R1965 VOUT_N.n2098 VOUT_N.n2097 0.0119325
R1966 VOUT_N.n995 VOUT_N.n994 0.0119325
R1967 VOUT_N.n1349 VOUT_N.n1348 0.0119325
R1968 VOUT_N.n1248 VOUT_N.n1247 0.0119325
R1969 VOUT_N.n1256 VOUT_N.n1250 0.0119325
R1970 VOUT_N.n1254 VOUT_N.n1253 0.0119325
R1971 VOUT_N.n1554 VOUT_N.n1553 0.0119325
R1972 VOUT_N.n1549 VOUT_N.n1548 0.0119325
R1973 VOUT_N.n1545 VOUT_N.n1544 0.0119325
R1974 VOUT_N.n1544 VOUT_N.n1543 0.0119325
R1975 VOUT_N.n1201 VOUT_N.n1200 0.0119325
R1976 VOUT_N.n1577 VOUT_N.n1576 0.0119325
R1977 VOUT_N.n1571 VOUT_N.n1570 0.0119325
R1978 VOUT_N.n1568 VOUT_N.n1567 0.0119325
R1979 VOUT_N.n1565 VOUT_N.n1564 0.0119325
R1980 VOUT_N.n1486 VOUT_N.n1477 0.0119325
R1981 VOUT_N.n1630 VOUT_N.n1629 0.0119325
R1982 VOUT_N.n1484 VOUT_N.n1483 0.0119325
R1983 VOUT_N.n1142 VOUT_N.n1141 0.0119325
R1984 VOUT_N.n353 VOUT_N.n352 0.0119325
R1985 VOUT_N.n808 VOUT_N.n807 0.0119325
R1986 VOUT_N.n852 VOUT_N.n851 0.0119325
R1987 VOUT_N.n894 VOUT_N.n893 0.0119325
R1988 VOUT_N.n896 VOUT_N.n895 0.0119325
R1989 VOUT_N.n901 VOUT_N.n900 0.0119325
R1990 VOUT_N.n941 VOUT_N.n940 0.0119325
R1991 VOUT_N.n1493 VOUT_N.n1492 0.0119325
R1992 VOUT_N.n1153 VOUT_N.n1152 0.0119325
R1993 VOUT_N.n402 VOUT_N.n401 0.0119325
R1994 VOUT_N.n609 VOUT_N.n608 0.0119325
R1995 VOUT_N.n32 VOUT_N.n31 0.0119325
R1996 VOUT_N.n1816 VOUT_N.n1815 0.0119325
R1997 VOUT_N.n1812 VOUT_N.n1811 0.0119325
R1998 VOUT_N.n1762 VOUT_N.n1761 0.0119325
R1999 VOUT_N.n1732 VOUT_N.n1731 0.0119325
R2000 VOUT_N.n2205 VOUT_N.n2204 0.0119325
R2001 VOUT_N.n1680 VOUT_N.n1679 0.0119325
R2002 VOUT_N.n1673 VOUT_N.n1672 0.0119325
R2003 VOUT_N.n1303 VOUT_N.n1302 0.0119325
R2004 VOUT_N.n1301 VOUT_N.n1300 0.0119325
R2005 VOUT_N.n944 VOUT_N.n943 0.0119325
R2006 VOUT_N.n614 VOUT_N.n613 0.0119325
R2007 VOUT_N.n181 VOUT_N.n180 0.0119325
R2008 VOUT_N.n174 VOUT_N.n173 0.0119325
R2009 VOUT_N.n4 VOUT_N.n3 0.0119325
R2010 VOUT_N.n2082 VOUT_N.n2081 0.00905634
R2011 VOUT_N.n2091 VOUT_N.n2090 0.00905634
R2012 VOUT_N.n1923 VOUT_N.n1922 0.00905634
R2013 VOUT_N.n1916 VOUT_N.n1915 0.00905634
R2014 VOUT_N.n1969 VOUT_N.n1968 0.00905634
R2015 VOUT_N.n1950 VOUT_N.n1949 0.00905634
R2016 VOUT_N.n2184 VOUT_N.n2183 0.00905634
R2017 VOUT_N.n2118 VOUT_N.n2117 0.00905634
R2018 VOUT_N.n1875 VOUT_N.n1874 0.00905634
R2019 VOUT_N.n1127 VOUT_N.n1126 0.00905634
R2020 VOUT_N.n1136 VOUT_N.n1135 0.00905634
R2021 VOUT_N.n1167 VOUT_N.n1166 0.00905634
R2022 VOUT_N.n1176 VOUT_N.n1175 0.00905634
R2023 VOUT_N.n1185 VOUT_N.n1184 0.00905634
R2024 VOUT_N.n1194 VOUT_N.n1193 0.00905634
R2025 VOUT_N.n1213 VOUT_N.n1212 0.00905634
R2026 VOUT_N.n1222 VOUT_N.n1221 0.00905634
R2027 VOUT_N.n1231 VOUT_N.n1230 0.00905634
R2028 VOUT_N.n1240 VOUT_N.n1239 0.00905634
R2029 VOUT_N.n1269 VOUT_N.n1268 0.00905634
R2030 VOUT_N.n1278 VOUT_N.n1277 0.00905634
R2031 VOUT_N.n1287 VOUT_N.n1286 0.00905634
R2032 VOUT_N.n1296 VOUT_N.n1295 0.00905634
R2033 VOUT_N.n1464 VOUT_N.n1463 0.00905634
R2034 VOUT_N.n1473 VOUT_N.n1472 0.00905634
R2035 VOUT_N.n1508 VOUT_N.n1507 0.00905634
R2036 VOUT_N.n1517 VOUT_N.n1516 0.00905634
R2037 VOUT_N.n1526 VOUT_N.n1525 0.00905634
R2038 VOUT_N.n1535 VOUT_N.n1534 0.00905634
R2039 VOUT_N.n1588 VOUT_N.n1587 0.00905634
R2040 VOUT_N.n1597 VOUT_N.n1596 0.00905634
R2041 VOUT_N.n1606 VOUT_N.n1605 0.00905634
R2042 VOUT_N.n1615 VOUT_N.n1614 0.00905634
R2043 VOUT_N.n1641 VOUT_N.n1640 0.00905634
R2044 VOUT_N.n1650 VOUT_N.n1649 0.00905634
R2045 VOUT_N.n1659 VOUT_N.n1658 0.00905634
R2046 VOUT_N.n1668 VOUT_N.n1667 0.00905634
R2047 VOUT_N.n792 VOUT_N.n791 0.00905634
R2048 VOUT_N.n801 VOUT_N.n800 0.00905634
R2049 VOUT_N.n820 VOUT_N.n819 0.00905634
R2050 VOUT_N.n829 VOUT_N.n828 0.00905634
R2051 VOUT_N.n838 VOUT_N.n837 0.00905634
R2052 VOUT_N.n847 VOUT_N.n846 0.00905634
R2053 VOUT_N.n864 VOUT_N.n863 0.00905634
R2054 VOUT_N.n873 VOUT_N.n872 0.00905634
R2055 VOUT_N.n882 VOUT_N.n881 0.00905634
R2056 VOUT_N.n891 VOUT_N.n890 0.00905634
R2057 VOUT_N.n910 VOUT_N.n909 0.00905634
R2058 VOUT_N.n919 VOUT_N.n918 0.00905634
R2059 VOUT_N.n928 VOUT_N.n927 0.00905634
R2060 VOUT_N.n937 VOUT_N.n936 0.00905634
R2061 VOUT_N.n336 VOUT_N.n335 0.00905634
R2062 VOUT_N.n345 VOUT_N.n344 0.00905634
R2063 VOUT_N.n373 VOUT_N.n372 0.00905634
R2064 VOUT_N.n382 VOUT_N.n381 0.00905634
R2065 VOUT_N.n391 VOUT_N.n390 0.00905634
R2066 VOUT_N.n400 VOUT_N.n399 0.00905634
R2067 VOUT_N.n422 VOUT_N.n421 0.00905634
R2068 VOUT_N.n431 VOUT_N.n430 0.00905634
R2069 VOUT_N.n440 VOUT_N.n439 0.00905634
R2070 VOUT_N.n449 VOUT_N.n448 0.00905634
R2071 VOUT_N.n475 VOUT_N.n474 0.00905634
R2072 VOUT_N.n484 VOUT_N.n483 0.00905634
R2073 VOUT_N.n493 VOUT_N.n492 0.00905634
R2074 VOUT_N.n502 VOUT_N.n501 0.00905634
R2075 VOUT_N.n600 VOUT_N.n599 0.00905634
R2076 VOUT_N.n591 VOUT_N.n590 0.00905634
R2077 VOUT_N.n582 VOUT_N.n581 0.00905634
R2078 VOUT_N.n564 VOUT_N.n563 0.00905634
R2079 VOUT_N.n555 VOUT_N.n554 0.00905634
R2080 VOUT_N.n1702 VOUT_N.n1701 0.00905634
R2081 VOUT_N.n2225 VOUT_N.n2224 0.00905634
R2082 VOUT_N.n2216 VOUT_N.n2215 0.00905634
R2083 VOUT_N.n2207 VOUT_N.n2206 0.00905634
R2084 VOUT_N.n2032 VOUT_N.n2031 0.00905634
R2085 VOUT_N.n1711 VOUT_N.n1710 0.00740328
R2086 VOUT_N.n2160 VOUT_N.n2159 0.00735609
R2087 VOUT_N.n1992 VOUT_N.n1991 0.00735609
R2088 VOUT_N.n1997 VOUT_N.n1996 0.00735609
R2089 VOUT_N.n2186 VOUT_N.n2185 0.00735609
R2090 VOUT_N.n22 VOUT_N.n21 0.00735609
R2091 VOUT_N.n27 VOUT_N.n26 0.00735609
R2092 VOUT_N.n1724 VOUT_N.n1723 0.00735609
R2093 VOUT_N.n1792 VOUT_N.n1791 0.00735609
R2094 VOUT_N.n1751 VOUT_N.n1750 0.00735609
R2095 VOUT_N.n1756 VOUT_N.n1755 0.00735609
R2096 VOUT_N.n73 VOUT_N.n72 0.00556853
R2097 VOUT_N.n87 VOUT_N.n86 0.00556853
R2098 VOUT_N.n81 VOUT_N.n80 0.00556853
R2099 VOUT_N.n158 VOUT_N.n157 0.00556853
R2100 VOUT_N.n163 VOUT_N.n162 0.00556853
R2101 VOUT_N.n138 VOUT_N.n137 0.00556853
R2102 VOUT_N.n141 VOUT_N.n140 0.00556853
R2103 VOUT_N.n112 VOUT_N.n111 0.00556853
R2104 VOUT_N.n118 VOUT_N.n117 0.00556853
R2105 VOUT_N.n124 VOUT_N.n123 0.00556853
R2106 VOUT_N.n135 VOUT_N.n134 0.00556853
R2107 VOUT_N.n134 VOUT_N.n133 0.00556853
R2108 VOUT_N.n157 VOUT_N.n156 0.00556853
R2109 VOUT_N.n117 VOUT_N.n116 0.00556853
R2110 VOUT_N.n142 VOUT_N.n141 0.00556853
R2111 VOUT_N.n123 VOUT_N.n122 0.00556853
R2112 VOUT_N.n164 VOUT_N.n163 0.00556853
R2113 VOUT_N.n137 VOUT_N.n136 0.00556853
R2114 VOUT_N.n111 VOUT_N.n110 0.00556853
R2115 VOUT_N.n41 VOUT_N.n40 0.00556853
R2116 VOUT_N.n46 VOUT_N.n45 0.00556853
R2117 VOUT_N.n53 VOUT_N.n52 0.00556853
R2118 VOUT_N.n59 VOUT_N.n58 0.00556853
R2119 VOUT_N.n58 VOUT_N.n57 0.00556853
R2120 VOUT_N.n47 VOUT_N.n46 0.00556853
R2121 VOUT_N.n52 VOUT_N.n51 0.00556853
R2122 VOUT_N.n40 VOUT_N.n39 0.00556853
R2123 VOUT_N.n82 VOUT_N.n81 0.00556853
R2124 VOUT_N.n96 VOUT_N.n95 0.00556853
R2125 VOUT_N.n88 VOUT_N.n87 0.00556853
R2126 VOUT_N.n331 VOUT_N.n330 0.00528925
R2127 VOUT_N.n335 VOUT_N.n334 0.00528925
R2128 VOUT_N.n340 VOUT_N.n339 0.00528925
R2129 VOUT_N.n556 VOUT_N.n555 0.00528925
R2130 VOUT_N.n560 VOUT_N.n559 0.00528925
R2131 VOUT_N.n565 VOUT_N.n564 0.00528925
R2132 VOUT_N.n2113 VOUT_N.n2112 0.00528925
R2133 VOUT_N.n1876 VOUT_N.n1875 0.00528925
R2134 VOUT_N.n1880 VOUT_N.n1879 0.00528925
R2135 VOUT_N.n2117 VOUT_N.n2116 0.00528925
R2136 VOUT_N.n1951 VOUT_N.n1950 0.00528925
R2137 VOUT_N.n1924 VOUT_N.n1923 0.00528925
R2138 VOUT_N.n1956 VOUT_N.n1955 0.00528925
R2139 VOUT_N.n2081 VOUT_N.n2072 0.00528925
R2140 VOUT_N.n2163 VOUT_N.n2162 0.00528925
R2141 VOUT_N.n2086 VOUT_N.n2085 0.00528925
R2142 VOUT_N.n2168 VOUT_N.n2167 0.00528925
R2143 VOUT_N.n2090 VOUT_N.n2089 0.00528925
R2144 VOUT_N.n1920 VOUT_N.n1919 0.00528925
R2145 VOUT_N.n578 VOUT_N.n577 0.00528925
R2146 VOUT_N.n583 VOUT_N.n582 0.00528925
R2147 VOUT_N.n587 VOUT_N.n586 0.00528925
R2148 VOUT_N.n592 VOUT_N.n591 0.00528925
R2149 VOUT_N.n596 VOUT_N.n595 0.00528925
R2150 VOUT_N.n601 VOUT_N.n600 0.00528925
R2151 VOUT_N.n787 VOUT_N.n786 0.00528925
R2152 VOUT_N.n791 VOUT_N.n790 0.00528925
R2153 VOUT_N.n796 VOUT_N.n795 0.00528925
R2154 VOUT_N.n800 VOUT_N.n799 0.00528925
R2155 VOUT_N.n815 VOUT_N.n814 0.00528925
R2156 VOUT_N.n819 VOUT_N.n818 0.00528925
R2157 VOUT_N.n824 VOUT_N.n823 0.00528925
R2158 VOUT_N.n828 VOUT_N.n827 0.00528925
R2159 VOUT_N.n833 VOUT_N.n832 0.00528925
R2160 VOUT_N.n837 VOUT_N.n836 0.00528925
R2161 VOUT_N.n842 VOUT_N.n841 0.00528925
R2162 VOUT_N.n936 VOUT_N.n935 0.00528925
R2163 VOUT_N.n932 VOUT_N.n931 0.00528925
R2164 VOUT_N.n927 VOUT_N.n926 0.00528925
R2165 VOUT_N.n923 VOUT_N.n922 0.00528925
R2166 VOUT_N.n918 VOUT_N.n917 0.00528925
R2167 VOUT_N.n914 VOUT_N.n913 0.00528925
R2168 VOUT_N.n909 VOUT_N.n908 0.00528925
R2169 VOUT_N.n905 VOUT_N.n904 0.00528925
R2170 VOUT_N.n890 VOUT_N.n889 0.00528925
R2171 VOUT_N.n886 VOUT_N.n885 0.00528925
R2172 VOUT_N.n881 VOUT_N.n880 0.00528925
R2173 VOUT_N.n877 VOUT_N.n876 0.00528925
R2174 VOUT_N.n872 VOUT_N.n871 0.00528925
R2175 VOUT_N.n868 VOUT_N.n867 0.00528925
R2176 VOUT_N.n863 VOUT_N.n862 0.00528925
R2177 VOUT_N.n859 VOUT_N.n858 0.00528925
R2178 VOUT_N.n846 VOUT_N.n845 0.00528925
R2179 VOUT_N.n1459 VOUT_N.n1458 0.00528925
R2180 VOUT_N.n1463 VOUT_N.n1462 0.00528925
R2181 VOUT_N.n1468 VOUT_N.n1467 0.00528925
R2182 VOUT_N.n1472 VOUT_N.n1471 0.00528925
R2183 VOUT_N.n1503 VOUT_N.n1502 0.00528925
R2184 VOUT_N.n1507 VOUT_N.n1506 0.00528925
R2185 VOUT_N.n1512 VOUT_N.n1511 0.00528925
R2186 VOUT_N.n1516 VOUT_N.n1515 0.00528925
R2187 VOUT_N.n1521 VOUT_N.n1520 0.00528925
R2188 VOUT_N.n1525 VOUT_N.n1524 0.00528925
R2189 VOUT_N.n1530 VOUT_N.n1529 0.00528925
R2190 VOUT_N.n1534 VOUT_N.n1533 0.00528925
R2191 VOUT_N.n1583 VOUT_N.n1582 0.00528925
R2192 VOUT_N.n1587 VOUT_N.n1586 0.00528925
R2193 VOUT_N.n1592 VOUT_N.n1591 0.00528925
R2194 VOUT_N.n1596 VOUT_N.n1595 0.00528925
R2195 VOUT_N.n1601 VOUT_N.n1600 0.00528925
R2196 VOUT_N.n1605 VOUT_N.n1604 0.00528925
R2197 VOUT_N.n1610 VOUT_N.n1609 0.00528925
R2198 VOUT_N.n1667 VOUT_N.n1666 0.00528925
R2199 VOUT_N.n1663 VOUT_N.n1662 0.00528925
R2200 VOUT_N.n1658 VOUT_N.n1657 0.00528925
R2201 VOUT_N.n1654 VOUT_N.n1653 0.00528925
R2202 VOUT_N.n1649 VOUT_N.n1648 0.00528925
R2203 VOUT_N.n1645 VOUT_N.n1644 0.00528925
R2204 VOUT_N.n1640 VOUT_N.n1639 0.00528925
R2205 VOUT_N.n1636 VOUT_N.n1635 0.00528925
R2206 VOUT_N.n1614 VOUT_N.n1613 0.00528925
R2207 VOUT_N.n1122 VOUT_N.n1121 0.00528925
R2208 VOUT_N.n1126 VOUT_N.n1125 0.00528925
R2209 VOUT_N.n1131 VOUT_N.n1130 0.00528925
R2210 VOUT_N.n1135 VOUT_N.n1134 0.00528925
R2211 VOUT_N.n1162 VOUT_N.n1161 0.00528925
R2212 VOUT_N.n1166 VOUT_N.n1165 0.00528925
R2213 VOUT_N.n1171 VOUT_N.n1170 0.00528925
R2214 VOUT_N.n1175 VOUT_N.n1174 0.00528925
R2215 VOUT_N.n1180 VOUT_N.n1179 0.00528925
R2216 VOUT_N.n1184 VOUT_N.n1183 0.00528925
R2217 VOUT_N.n1189 VOUT_N.n1188 0.00528925
R2218 VOUT_N.n1193 VOUT_N.n1192 0.00528925
R2219 VOUT_N.n1208 VOUT_N.n1207 0.00528925
R2220 VOUT_N.n1212 VOUT_N.n1211 0.00528925
R2221 VOUT_N.n1217 VOUT_N.n1216 0.00528925
R2222 VOUT_N.n1221 VOUT_N.n1220 0.00528925
R2223 VOUT_N.n1226 VOUT_N.n1225 0.00528925
R2224 VOUT_N.n1230 VOUT_N.n1229 0.00528925
R2225 VOUT_N.n1235 VOUT_N.n1234 0.00528925
R2226 VOUT_N.n1295 VOUT_N.n1294 0.00528925
R2227 VOUT_N.n1291 VOUT_N.n1290 0.00528925
R2228 VOUT_N.n1286 VOUT_N.n1285 0.00528925
R2229 VOUT_N.n1282 VOUT_N.n1281 0.00528925
R2230 VOUT_N.n1277 VOUT_N.n1276 0.00528925
R2231 VOUT_N.n1273 VOUT_N.n1272 0.00528925
R2232 VOUT_N.n1268 VOUT_N.n1267 0.00528925
R2233 VOUT_N.n1264 VOUT_N.n1263 0.00528925
R2234 VOUT_N.n1239 VOUT_N.n1238 0.00528925
R2235 VOUT_N.n344 VOUT_N.n343 0.00528925
R2236 VOUT_N.n368 VOUT_N.n367 0.00528925
R2237 VOUT_N.n372 VOUT_N.n371 0.00528925
R2238 VOUT_N.n377 VOUT_N.n376 0.00528925
R2239 VOUT_N.n381 VOUT_N.n380 0.00528925
R2240 VOUT_N.n386 VOUT_N.n385 0.00528925
R2241 VOUT_N.n390 VOUT_N.n389 0.00528925
R2242 VOUT_N.n395 VOUT_N.n394 0.00528925
R2243 VOUT_N.n399 VOUT_N.n398 0.00528925
R2244 VOUT_N.n417 VOUT_N.n416 0.00528925
R2245 VOUT_N.n421 VOUT_N.n420 0.00528925
R2246 VOUT_N.n426 VOUT_N.n425 0.00528925
R2247 VOUT_N.n430 VOUT_N.n429 0.00528925
R2248 VOUT_N.n435 VOUT_N.n434 0.00528925
R2249 VOUT_N.n439 VOUT_N.n438 0.00528925
R2250 VOUT_N.n444 VOUT_N.n443 0.00528925
R2251 VOUT_N.n448 VOUT_N.n447 0.00528925
R2252 VOUT_N.n470 VOUT_N.n469 0.00528925
R2253 VOUT_N.n474 VOUT_N.n473 0.00528925
R2254 VOUT_N.n479 VOUT_N.n478 0.00528925
R2255 VOUT_N.n483 VOUT_N.n482 0.00528925
R2256 VOUT_N.n488 VOUT_N.n487 0.00528925
R2257 VOUT_N.n492 VOUT_N.n491 0.00528925
R2258 VOUT_N.n497 VOUT_N.n496 0.00528925
R2259 VOUT_N.n501 VOUT_N.n500 0.00528925
R2260 VOUT_N.n1796 VOUT_N.n1795 0.00528925
R2261 VOUT_N.n1705 VOUT_N.n1704 0.00528925
R2262 VOUT_N.n1801 VOUT_N.n1800 0.00528925
R2263 VOUT_N.n2230 VOUT_N.n2229 0.00528925
R2264 VOUT_N.n2226 VOUT_N.n2225 0.00528925
R2265 VOUT_N.n2221 VOUT_N.n2220 0.00528925
R2266 VOUT_N.n2217 VOUT_N.n2216 0.00528925
R2267 VOUT_N.n2212 VOUT_N.n2211 0.00528925
R2268 VOUT_N.n2208 VOUT_N.n2207 0.00528925
R2269 VOUT_N.n2037 VOUT_N.n2036 0.00528925
R2270 VOUT_N.n2033 VOUT_N.n2032 0.00528925
R2271 VOUT_N.n2029 VOUT_N.n2028 0.00528925
R2272 VOUT_N.n2084 VOUT_N.n2083 0.00527411
R2273 VOUT_N.n1918 VOUT_N.n1917 0.00527411
R2274 VOUT_N.n2085 VOUT_N.n2084 0.00527411
R2275 VOUT_N.n1919 VOUT_N.n1918 0.00527411
R2276 VOUT_N.n2165 VOUT_N.n2164 0.00527411
R2277 VOUT_N.n2170 VOUT_N.n2169 0.00527411
R2278 VOUT_N.n1959 VOUT_N.n1958 0.00527411
R2279 VOUT_N.n1954 VOUT_N.n1953 0.00527411
R2280 VOUT_N.n2164 VOUT_N.n2163 0.00527411
R2281 VOUT_N.n2169 VOUT_N.n2168 0.00527411
R2282 VOUT_N.n1955 VOUT_N.n1954 0.00527411
R2283 VOUT_N.n1968 VOUT_N.n1959 0.00527411
R2284 VOUT_N.n2195 VOUT_N.n2194 0.00527411
R2285 VOUT_N.n1994 VOUT_N.n1993 0.00527411
R2286 VOUT_N.n1995 VOUT_N.n1994 0.00527411
R2287 VOUT_N.n2194 VOUT_N.n2193 0.00527411
R2288 VOUT_N.n1882 VOUT_N.n1881 0.00527411
R2289 VOUT_N.n1881 VOUT_N.n1880 0.00527411
R2290 VOUT_N.n2112 VOUT_N.n2111 0.00527411
R2291 VOUT_N.n1129 VOUT_N.n1128 0.00527411
R2292 VOUT_N.n1160 VOUT_N.n1159 0.00527411
R2293 VOUT_N.n1169 VOUT_N.n1168 0.00527411
R2294 VOUT_N.n1178 VOUT_N.n1177 0.00527411
R2295 VOUT_N.n1187 VOUT_N.n1186 0.00527411
R2296 VOUT_N.n1206 VOUT_N.n1205 0.00527411
R2297 VOUT_N.n1215 VOUT_N.n1214 0.00527411
R2298 VOUT_N.n1224 VOUT_N.n1223 0.00527411
R2299 VOUT_N.n1233 VOUT_N.n1232 0.00527411
R2300 VOUT_N.n1262 VOUT_N.n1261 0.00527411
R2301 VOUT_N.n1271 VOUT_N.n1270 0.00527411
R2302 VOUT_N.n1280 VOUT_N.n1279 0.00527411
R2303 VOUT_N.n1289 VOUT_N.n1288 0.00527411
R2304 VOUT_N.n1263 VOUT_N.n1262 0.00527411
R2305 VOUT_N.n1272 VOUT_N.n1271 0.00527411
R2306 VOUT_N.n1281 VOUT_N.n1280 0.00527411
R2307 VOUT_N.n1290 VOUT_N.n1289 0.00527411
R2308 VOUT_N.n1234 VOUT_N.n1233 0.00527411
R2309 VOUT_N.n1225 VOUT_N.n1224 0.00527411
R2310 VOUT_N.n1216 VOUT_N.n1215 0.00527411
R2311 VOUT_N.n1207 VOUT_N.n1206 0.00527411
R2312 VOUT_N.n1188 VOUT_N.n1187 0.00527411
R2313 VOUT_N.n1179 VOUT_N.n1178 0.00527411
R2314 VOUT_N.n1170 VOUT_N.n1169 0.00527411
R2315 VOUT_N.n1161 VOUT_N.n1160 0.00527411
R2316 VOUT_N.n1130 VOUT_N.n1129 0.00527411
R2317 VOUT_N.n1121 VOUT_N.n1120 0.00527411
R2318 VOUT_N.n1466 VOUT_N.n1465 0.00527411
R2319 VOUT_N.n1501 VOUT_N.n1500 0.00527411
R2320 VOUT_N.n1510 VOUT_N.n1509 0.00527411
R2321 VOUT_N.n1519 VOUT_N.n1518 0.00527411
R2322 VOUT_N.n1528 VOUT_N.n1527 0.00527411
R2323 VOUT_N.n1581 VOUT_N.n1580 0.00527411
R2324 VOUT_N.n1590 VOUT_N.n1589 0.00527411
R2325 VOUT_N.n1599 VOUT_N.n1598 0.00527411
R2326 VOUT_N.n1608 VOUT_N.n1607 0.00527411
R2327 VOUT_N.n1634 VOUT_N.n1633 0.00527411
R2328 VOUT_N.n1643 VOUT_N.n1642 0.00527411
R2329 VOUT_N.n1652 VOUT_N.n1651 0.00527411
R2330 VOUT_N.n1661 VOUT_N.n1660 0.00527411
R2331 VOUT_N.n1635 VOUT_N.n1634 0.00527411
R2332 VOUT_N.n1644 VOUT_N.n1643 0.00527411
R2333 VOUT_N.n1653 VOUT_N.n1652 0.00527411
R2334 VOUT_N.n1662 VOUT_N.n1661 0.00527411
R2335 VOUT_N.n1609 VOUT_N.n1608 0.00527411
R2336 VOUT_N.n1600 VOUT_N.n1599 0.00527411
R2337 VOUT_N.n1591 VOUT_N.n1590 0.00527411
R2338 VOUT_N.n1582 VOUT_N.n1581 0.00527411
R2339 VOUT_N.n1529 VOUT_N.n1528 0.00527411
R2340 VOUT_N.n1520 VOUT_N.n1519 0.00527411
R2341 VOUT_N.n1511 VOUT_N.n1510 0.00527411
R2342 VOUT_N.n1502 VOUT_N.n1501 0.00527411
R2343 VOUT_N.n1467 VOUT_N.n1466 0.00527411
R2344 VOUT_N.n1458 VOUT_N.n1457 0.00527411
R2345 VOUT_N.n794 VOUT_N.n793 0.00527411
R2346 VOUT_N.n813 VOUT_N.n812 0.00527411
R2347 VOUT_N.n822 VOUT_N.n821 0.00527411
R2348 VOUT_N.n831 VOUT_N.n830 0.00527411
R2349 VOUT_N.n840 VOUT_N.n839 0.00527411
R2350 VOUT_N.n857 VOUT_N.n856 0.00527411
R2351 VOUT_N.n866 VOUT_N.n865 0.00527411
R2352 VOUT_N.n875 VOUT_N.n874 0.00527411
R2353 VOUT_N.n884 VOUT_N.n883 0.00527411
R2354 VOUT_N.n903 VOUT_N.n902 0.00527411
R2355 VOUT_N.n912 VOUT_N.n911 0.00527411
R2356 VOUT_N.n921 VOUT_N.n920 0.00527411
R2357 VOUT_N.n930 VOUT_N.n929 0.00527411
R2358 VOUT_N.n858 VOUT_N.n857 0.00527411
R2359 VOUT_N.n867 VOUT_N.n866 0.00527411
R2360 VOUT_N.n876 VOUT_N.n875 0.00527411
R2361 VOUT_N.n885 VOUT_N.n884 0.00527411
R2362 VOUT_N.n904 VOUT_N.n903 0.00527411
R2363 VOUT_N.n913 VOUT_N.n912 0.00527411
R2364 VOUT_N.n922 VOUT_N.n921 0.00527411
R2365 VOUT_N.n931 VOUT_N.n930 0.00527411
R2366 VOUT_N.n841 VOUT_N.n840 0.00527411
R2367 VOUT_N.n832 VOUT_N.n831 0.00527411
R2368 VOUT_N.n823 VOUT_N.n822 0.00527411
R2369 VOUT_N.n814 VOUT_N.n813 0.00527411
R2370 VOUT_N.n795 VOUT_N.n794 0.00527411
R2371 VOUT_N.n786 VOUT_N.n785 0.00527411
R2372 VOUT_N.n338 VOUT_N.n337 0.00527411
R2373 VOUT_N.n366 VOUT_N.n365 0.00527411
R2374 VOUT_N.n375 VOUT_N.n374 0.00527411
R2375 VOUT_N.n384 VOUT_N.n383 0.00527411
R2376 VOUT_N.n393 VOUT_N.n392 0.00527411
R2377 VOUT_N.n415 VOUT_N.n414 0.00527411
R2378 VOUT_N.n424 VOUT_N.n423 0.00527411
R2379 VOUT_N.n433 VOUT_N.n432 0.00527411
R2380 VOUT_N.n442 VOUT_N.n441 0.00527411
R2381 VOUT_N.n468 VOUT_N.n467 0.00527411
R2382 VOUT_N.n477 VOUT_N.n476 0.00527411
R2383 VOUT_N.n486 VOUT_N.n485 0.00527411
R2384 VOUT_N.n495 VOUT_N.n494 0.00527411
R2385 VOUT_N.n598 VOUT_N.n597 0.00527411
R2386 VOUT_N.n589 VOUT_N.n588 0.00527411
R2387 VOUT_N.n580 VOUT_N.n579 0.00527411
R2388 VOUT_N.n562 VOUT_N.n561 0.00527411
R2389 VOUT_N.n496 VOUT_N.n495 0.00527411
R2390 VOUT_N.n487 VOUT_N.n486 0.00527411
R2391 VOUT_N.n478 VOUT_N.n477 0.00527411
R2392 VOUT_N.n469 VOUT_N.n468 0.00527411
R2393 VOUT_N.n443 VOUT_N.n442 0.00527411
R2394 VOUT_N.n434 VOUT_N.n433 0.00527411
R2395 VOUT_N.n425 VOUT_N.n424 0.00527411
R2396 VOUT_N.n416 VOUT_N.n415 0.00527411
R2397 VOUT_N.n394 VOUT_N.n393 0.00527411
R2398 VOUT_N.n385 VOUT_N.n384 0.00527411
R2399 VOUT_N.n376 VOUT_N.n375 0.00527411
R2400 VOUT_N.n367 VOUT_N.n366 0.00527411
R2401 VOUT_N.n597 VOUT_N.n596 0.00527411
R2402 VOUT_N.n588 VOUT_N.n587 0.00527411
R2403 VOUT_N.n579 VOUT_N.n578 0.00527411
R2404 VOUT_N.n561 VOUT_N.n560 0.00527411
R2405 VOUT_N.n339 VOUT_N.n338 0.00527411
R2406 VOUT_N.n330 VOUT_N.n329 0.00527411
R2407 VOUT_N.n24 VOUT_N.n23 0.00527411
R2408 VOUT_N.n25 VOUT_N.n24 0.00527411
R2409 VOUT_N.n1713 VOUT_N.n1712 0.00527411
R2410 VOUT_N.n1722 VOUT_N.n1713 0.00527411
R2411 VOUT_N.n1799 VOUT_N.n1798 0.00527411
R2412 VOUT_N.n1794 VOUT_N.n1793 0.00527411
R2413 VOUT_N.n1795 VOUT_N.n1794 0.00527411
R2414 VOUT_N.n1800 VOUT_N.n1799 0.00527411
R2415 VOUT_N.n1753 VOUT_N.n1752 0.00527411
R2416 VOUT_N.n1754 VOUT_N.n1753 0.00527411
R2417 VOUT_N.n2232 VOUT_N.n2231 0.00527411
R2418 VOUT_N.n2223 VOUT_N.n2222 0.00527411
R2419 VOUT_N.n2214 VOUT_N.n2213 0.00527411
R2420 VOUT_N.n2039 VOUT_N.n2038 0.00527411
R2421 VOUT_N.n2027 VOUT_N.n2026 0.00527411
R2422 VOUT_N.n2038 VOUT_N.n2037 0.00527411
R2423 VOUT_N.n2213 VOUT_N.n2212 0.00527411
R2424 VOUT_N.n2222 VOUT_N.n2221 0.00527411
R2425 VOUT_N.n2231 VOUT_N.n2230 0.00527411
R2426 VOUT_N.n2028 VOUT_N.n2027 0.00527411
R2427 VOUT_N.n2087 VOUT_N.n2086 0.00525899
R2428 VOUT_N.n2089 VOUT_N.n2088 0.00525899
R2429 VOUT_N.n1925 VOUT_N.n1924 0.00525899
R2430 VOUT_N.n1921 VOUT_N.n1920 0.00525899
R2431 VOUT_N.n2162 VOUT_N.n2161 0.00525899
R2432 VOUT_N.n2167 VOUT_N.n2166 0.00525899
R2433 VOUT_N.n1957 VOUT_N.n1956 0.00525899
R2434 VOUT_N.n1952 VOUT_N.n1951 0.00525899
R2435 VOUT_N.n2114 VOUT_N.n2113 0.00525899
R2436 VOUT_N.n2116 VOUT_N.n2115 0.00525899
R2437 VOUT_N.n1879 VOUT_N.n1878 0.00525899
R2438 VOUT_N.n1877 VOUT_N.n1876 0.00525899
R2439 VOUT_N.n1123 VOUT_N.n1122 0.00525899
R2440 VOUT_N.n1125 VOUT_N.n1124 0.00525899
R2441 VOUT_N.n1132 VOUT_N.n1131 0.00525899
R2442 VOUT_N.n1134 VOUT_N.n1133 0.00525899
R2443 VOUT_N.n1163 VOUT_N.n1162 0.00525899
R2444 VOUT_N.n1165 VOUT_N.n1164 0.00525899
R2445 VOUT_N.n1172 VOUT_N.n1171 0.00525899
R2446 VOUT_N.n1174 VOUT_N.n1173 0.00525899
R2447 VOUT_N.n1181 VOUT_N.n1180 0.00525899
R2448 VOUT_N.n1183 VOUT_N.n1182 0.00525899
R2449 VOUT_N.n1190 VOUT_N.n1189 0.00525899
R2450 VOUT_N.n1192 VOUT_N.n1191 0.00525899
R2451 VOUT_N.n1209 VOUT_N.n1208 0.00525899
R2452 VOUT_N.n1211 VOUT_N.n1210 0.00525899
R2453 VOUT_N.n1218 VOUT_N.n1217 0.00525899
R2454 VOUT_N.n1220 VOUT_N.n1219 0.00525899
R2455 VOUT_N.n1227 VOUT_N.n1226 0.00525899
R2456 VOUT_N.n1229 VOUT_N.n1228 0.00525899
R2457 VOUT_N.n1236 VOUT_N.n1235 0.00525899
R2458 VOUT_N.n1238 VOUT_N.n1237 0.00525899
R2459 VOUT_N.n1265 VOUT_N.n1264 0.00525899
R2460 VOUT_N.n1267 VOUT_N.n1266 0.00525899
R2461 VOUT_N.n1274 VOUT_N.n1273 0.00525899
R2462 VOUT_N.n1276 VOUT_N.n1275 0.00525899
R2463 VOUT_N.n1283 VOUT_N.n1282 0.00525899
R2464 VOUT_N.n1285 VOUT_N.n1284 0.00525899
R2465 VOUT_N.n1292 VOUT_N.n1291 0.00525899
R2466 VOUT_N.n1294 VOUT_N.n1293 0.00525899
R2467 VOUT_N.n1460 VOUT_N.n1459 0.00525899
R2468 VOUT_N.n1462 VOUT_N.n1461 0.00525899
R2469 VOUT_N.n1469 VOUT_N.n1468 0.00525899
R2470 VOUT_N.n1471 VOUT_N.n1470 0.00525899
R2471 VOUT_N.n1504 VOUT_N.n1503 0.00525899
R2472 VOUT_N.n1506 VOUT_N.n1505 0.00525899
R2473 VOUT_N.n1513 VOUT_N.n1512 0.00525899
R2474 VOUT_N.n1515 VOUT_N.n1514 0.00525899
R2475 VOUT_N.n1522 VOUT_N.n1521 0.00525899
R2476 VOUT_N.n1524 VOUT_N.n1523 0.00525899
R2477 VOUT_N.n1531 VOUT_N.n1530 0.00525899
R2478 VOUT_N.n1533 VOUT_N.n1532 0.00525899
R2479 VOUT_N.n1584 VOUT_N.n1583 0.00525899
R2480 VOUT_N.n1586 VOUT_N.n1585 0.00525899
R2481 VOUT_N.n1593 VOUT_N.n1592 0.00525899
R2482 VOUT_N.n1595 VOUT_N.n1594 0.00525899
R2483 VOUT_N.n1602 VOUT_N.n1601 0.00525899
R2484 VOUT_N.n1604 VOUT_N.n1603 0.00525899
R2485 VOUT_N.n1611 VOUT_N.n1610 0.00525899
R2486 VOUT_N.n1613 VOUT_N.n1612 0.00525899
R2487 VOUT_N.n1637 VOUT_N.n1636 0.00525899
R2488 VOUT_N.n1639 VOUT_N.n1638 0.00525899
R2489 VOUT_N.n1646 VOUT_N.n1645 0.00525899
R2490 VOUT_N.n1648 VOUT_N.n1647 0.00525899
R2491 VOUT_N.n1655 VOUT_N.n1654 0.00525899
R2492 VOUT_N.n1657 VOUT_N.n1656 0.00525899
R2493 VOUT_N.n1664 VOUT_N.n1663 0.00525899
R2494 VOUT_N.n1666 VOUT_N.n1665 0.00525899
R2495 VOUT_N.n788 VOUT_N.n787 0.00525899
R2496 VOUT_N.n790 VOUT_N.n789 0.00525899
R2497 VOUT_N.n797 VOUT_N.n796 0.00525899
R2498 VOUT_N.n799 VOUT_N.n798 0.00525899
R2499 VOUT_N.n816 VOUT_N.n815 0.00525899
R2500 VOUT_N.n818 VOUT_N.n817 0.00525899
R2501 VOUT_N.n825 VOUT_N.n824 0.00525899
R2502 VOUT_N.n827 VOUT_N.n826 0.00525899
R2503 VOUT_N.n834 VOUT_N.n833 0.00525899
R2504 VOUT_N.n836 VOUT_N.n835 0.00525899
R2505 VOUT_N.n843 VOUT_N.n842 0.00525899
R2506 VOUT_N.n845 VOUT_N.n844 0.00525899
R2507 VOUT_N.n860 VOUT_N.n859 0.00525899
R2508 VOUT_N.n862 VOUT_N.n861 0.00525899
R2509 VOUT_N.n869 VOUT_N.n868 0.00525899
R2510 VOUT_N.n871 VOUT_N.n870 0.00525899
R2511 VOUT_N.n878 VOUT_N.n877 0.00525899
R2512 VOUT_N.n880 VOUT_N.n879 0.00525899
R2513 VOUT_N.n887 VOUT_N.n886 0.00525899
R2514 VOUT_N.n889 VOUT_N.n888 0.00525899
R2515 VOUT_N.n906 VOUT_N.n905 0.00525899
R2516 VOUT_N.n908 VOUT_N.n907 0.00525899
R2517 VOUT_N.n915 VOUT_N.n914 0.00525899
R2518 VOUT_N.n917 VOUT_N.n916 0.00525899
R2519 VOUT_N.n924 VOUT_N.n923 0.00525899
R2520 VOUT_N.n926 VOUT_N.n925 0.00525899
R2521 VOUT_N.n933 VOUT_N.n932 0.00525899
R2522 VOUT_N.n935 VOUT_N.n934 0.00525899
R2523 VOUT_N.n332 VOUT_N.n331 0.00525899
R2524 VOUT_N.n334 VOUT_N.n333 0.00525899
R2525 VOUT_N.n341 VOUT_N.n340 0.00525899
R2526 VOUT_N.n343 VOUT_N.n342 0.00525899
R2527 VOUT_N.n369 VOUT_N.n368 0.00525899
R2528 VOUT_N.n371 VOUT_N.n370 0.00525899
R2529 VOUT_N.n378 VOUT_N.n377 0.00525899
R2530 VOUT_N.n380 VOUT_N.n379 0.00525899
R2531 VOUT_N.n387 VOUT_N.n386 0.00525899
R2532 VOUT_N.n389 VOUT_N.n388 0.00525899
R2533 VOUT_N.n396 VOUT_N.n395 0.00525899
R2534 VOUT_N.n398 VOUT_N.n397 0.00525899
R2535 VOUT_N.n418 VOUT_N.n417 0.00525899
R2536 VOUT_N.n420 VOUT_N.n419 0.00525899
R2537 VOUT_N.n427 VOUT_N.n426 0.00525899
R2538 VOUT_N.n429 VOUT_N.n428 0.00525899
R2539 VOUT_N.n436 VOUT_N.n435 0.00525899
R2540 VOUT_N.n438 VOUT_N.n437 0.00525899
R2541 VOUT_N.n445 VOUT_N.n444 0.00525899
R2542 VOUT_N.n447 VOUT_N.n446 0.00525899
R2543 VOUT_N.n471 VOUT_N.n470 0.00525899
R2544 VOUT_N.n473 VOUT_N.n472 0.00525899
R2545 VOUT_N.n480 VOUT_N.n479 0.00525899
R2546 VOUT_N.n482 VOUT_N.n481 0.00525899
R2547 VOUT_N.n489 VOUT_N.n488 0.00525899
R2548 VOUT_N.n491 VOUT_N.n490 0.00525899
R2549 VOUT_N.n498 VOUT_N.n497 0.00525899
R2550 VOUT_N.n500 VOUT_N.n499 0.00525899
R2551 VOUT_N.n602 VOUT_N.n601 0.00525899
R2552 VOUT_N.n595 VOUT_N.n594 0.00525899
R2553 VOUT_N.n593 VOUT_N.n592 0.00525899
R2554 VOUT_N.n586 VOUT_N.n585 0.00525899
R2555 VOUT_N.n584 VOUT_N.n583 0.00525899
R2556 VOUT_N.n577 VOUT_N.n576 0.00525899
R2557 VOUT_N.n566 VOUT_N.n565 0.00525899
R2558 VOUT_N.n559 VOUT_N.n558 0.00525899
R2559 VOUT_N.n557 VOUT_N.n556 0.00525899
R2560 VOUT_N.n1704 VOUT_N.n1703 0.00525899
R2561 VOUT_N.n1797 VOUT_N.n1796 0.00525899
R2562 VOUT_N.n1802 VOUT_N.n1801 0.00525899
R2563 VOUT_N.n2229 VOUT_N.n2228 0.00525899
R2564 VOUT_N.n2227 VOUT_N.n2226 0.00525899
R2565 VOUT_N.n2220 VOUT_N.n2219 0.00525899
R2566 VOUT_N.n2218 VOUT_N.n2217 0.00525899
R2567 VOUT_N.n2211 VOUT_N.n2210 0.00525899
R2568 VOUT_N.n2209 VOUT_N.n2208 0.00525899
R2569 VOUT_N.n2036 VOUT_N.n2035 0.00525899
R2570 VOUT_N.n2034 VOUT_N.n2033 0.00525899
R2571 VOUT_N.n2030 VOUT_N.n2029 0.00525899
R2572 VOUT_N.n153 VOUT_N.n152 0.00495689
R2573 VOUT_N.n159 VOUT_N.n158 0.00495689
R2574 VOUT_N.n162 VOUT_N.n161 0.00495689
R2575 VOUT_N.n145 VOUT_N.n135 0.00495689
R2576 VOUT_N.n168 VOUT_N.n167 0.00495689
R2577 VOUT_N.n156 VOUT_N.n155 0.00495689
R2578 VOUT_N.n128 VOUT_N.n127 0.00495689
R2579 VOUT_N.n54 VOUT_N.n53 0.00495689
R2580 VOUT_N.n66 VOUT_N.n59 0.00495689
R2581 VOUT_N.n116 VOUT_N.n115 0.00495689
R2582 VOUT_N.n110 VOUT_N.n109 0.00495689
R2583 VOUT_N.n113 VOUT_N.n112 0.00495689
R2584 VOUT_N.n91 VOUT_N.n73 0.00495689
R2585 VOUT_N.n97 VOUT_N.n96 0.00429028
R2586 VOUT_N.n105 VOUT_N.n104 0.00429028
R2587 VOUT_N.n94 VOUT_N.n93 0.00429028
R2588 VOUT_N.n2159 VOUT_N.n2154 0.00418876
R2589 VOUT_N.n2193 VOUT_N.n2186 0.00418876
R2590 VOUT_N.n1996 VOUT_N.n1995 0.00418876
R2591 VOUT_N.n1991 VOUT_N.n1990 0.00418876
R2592 VOUT_N.n26 VOUT_N.n25 0.00418876
R2593 VOUT_N.n21 VOUT_N.n20 0.00418876
R2594 VOUT_N.n1723 VOUT_N.n1722 0.00418876
R2595 VOUT_N.n1791 VOUT_N.n1790 0.00418876
R2596 VOUT_N.n1755 VOUT_N.n1754 0.00418876
R2597 VOUT_N.n1750 VOUT_N.n1749 0.00418876
R2598 VOUT_N.n65 VOUT_N.n61 0.00346816
R2599 VOUT_N.n64 VOUT_N.n63 0.00346816
R2600 VOUT_N.n89 VOUT_N.n88 0.00346816
R2601 VOUT_N.n85 VOUT_N.n84 0.00346816
R2602 VOUT_N.n83 VOUT_N.n82 0.00346816
R2603 VOUT_N.n79 VOUT_N.n78 0.00346816
R2604 VOUT_N.n77 VOUT_N.n76 0.00346816
R2605 VOUT_N.n165 VOUT_N.n164 0.00346816
R2606 VOUT_N.n144 VOUT_N.n139 0.00346816
R2607 VOUT_N.n143 VOUT_N.n142 0.00346816
R2608 VOUT_N.n108 VOUT_N.n107 0.00346816
R2609 VOUT_N.n120 VOUT_N.n119 0.00346816
R2610 VOUT_N.n122 VOUT_N.n121 0.00346816
R2611 VOUT_N.n131 VOUT_N.n125 0.00346816
R2612 VOUT_N.n133 VOUT_N.n132 0.00346816
R2613 VOUT_N.n139 VOUT_N.n138 0.00346816
R2614 VOUT_N.n107 VOUT_N.n106 0.00346816
R2615 VOUT_N.n119 VOUT_N.n118 0.00346816
R2616 VOUT_N.n125 VOUT_N.n124 0.00346816
R2617 VOUT_N.n121 VOUT_N.n120 0.00346816
R2618 VOUT_N.n166 VOUT_N.n165 0.00346816
R2619 VOUT_N.n144 VOUT_N.n143 0.00346816
R2620 VOUT_N.n132 VOUT_N.n131 0.00346816
R2621 VOUT_N.n37 VOUT_N.n36 0.00346816
R2622 VOUT_N.n39 VOUT_N.n38 0.00346816
R2623 VOUT_N.n43 VOUT_N.n42 0.00346816
R2624 VOUT_N.n45 VOUT_N.n44 0.00346816
R2625 VOUT_N.n49 VOUT_N.n48 0.00346816
R2626 VOUT_N.n51 VOUT_N.n50 0.00346816
R2627 VOUT_N.n57 VOUT_N.n56 0.00346816
R2628 VOUT_N.n84 VOUT_N.n83 0.00346816
R2629 VOUT_N.n50 VOUT_N.n49 0.00346816
R2630 VOUT_N.n90 VOUT_N.n89 0.00346816
R2631 VOUT_N.n44 VOUT_N.n43 0.00346816
R2632 VOUT_N.n38 VOUT_N.n37 0.00346816
R2633 VOUT_N.n36 VOUT_N.n35 0.00346816
R2634 VOUT_N.n86 VOUT_N.n85 0.00346816
R2635 VOUT_N.n42 VOUT_N.n41 0.00346816
R2636 VOUT_N.n65 VOUT_N.n64 0.00346816
R2637 VOUT_N.n61 VOUT_N.n60 0.00346816
R2638 VOUT_N.n78 VOUT_N.n77 0.00346816
R2639 VOUT_N.n80 VOUT_N.n79 0.00346816
R2640 VOUT_N.n48 VOUT_N.n47 0.00346816
R2641 VOUT_N.n56 VOUT_N.n55 0.00346816
R2642 VOUT_N.n1710 VOUT_N.n1705 0.00314088
R2643 VOUT_N.n114 VOUT_N.n113 0.00297812
R2644 VOUT_N.n161 VOUT_N.n160 0.00297812
R2645 VOUT_N.n166 VOUT_N.n159 0.00297812
R2646 VOUT_N.n151 VOUT_N.n145 0.00297812
R2647 VOUT_N.n154 VOUT_N.n153 0.00297812
R2648 VOUT_N.n155 VOUT_N.n154 0.00297812
R2649 VOUT_N.n115 VOUT_N.n114 0.00297812
R2650 VOUT_N.n129 VOUT_N.n128 0.00297812
R2651 VOUT_N.n109 VOUT_N.n108 0.00297812
R2652 VOUT_N.n130 VOUT_N.n129 0.00297812
R2653 VOUT_N.n167 VOUT_N.n151 0.00297812
R2654 VOUT_N.n92 VOUT_N.n66 0.00297812
R2655 VOUT_N.n55 VOUT_N.n54 0.00297812
R2656 VOUT_N.n91 VOUT_N.n90 0.00297812
R2657 VOUT_N.n2154 VOUT_N.n2153 0.00284163
R2658 VOUT_N.n103 VOUT_N.n94 0.00264514
R2659 VOUT_N.n104 VOUT_N.n92 0.00264514
R2660 VOUT_N.n103 VOUT_N.n97 0.00264514
R2661 VOUT_N.n1990 VOUT_N.n1989 0.00219433
R2662 VOUT_N.n20 VOUT_N.n19 0.00219433
R2663 VOUT_N.n1790 VOUT_N.n1789 0.00219433
R2664 VOUT_N.n1749 VOUT_N.n1748 0.00219433
R2665 VOUT_N.n1915 VOUT_N.n1914 0.00192237
R2666 VOUT_N.n1701 VOUT_N.n1700 0.00192237
R2667 VOUT_N.n2183 VOUT_N.n2182 0.00192078
R2668 VSS.t319 VSS.t460 122.014
R2669 VSS.t404 VSS.t458 122.014
R2670 VSS.t289 VSS.t383 122.014
R2671 VSS.t410 VSS.t347 122.014
R2672 VSS.t369 VSS.t421 122.014
R2673 VSS.t292 VSS.t449 122.014
R2674 VSS.t466 VSS.t329 122.014
R2675 VSS.t402 VSS.t331 122.014
R2676 VSS.t373 VSS.t427 122.014
R2677 VSS.t387 VSS.t298 122.014
R2678 VSS.t456 VSS.t301 122.014
R2679 VSS.t349 VSS.t475 122.014
R2680 VSS.t406 VSS.t362 112.368
R2681 VSS.t351 VSS.t406 112.368
R2682 VSS.t470 VSS.t418 112.368
R2683 VSS.t423 VSS.t470 112.368
R2684 VSS.t313 VSS.t425 112.368
R2685 VSS.t371 VSS.t313 112.368
R2686 VSS.t429 VSS.t371 112.368
R2687 VSS.t462 VSS.t429 112.368
R2688 VSS.t356 VSS.t462 112.368
R2689 VSS.t481 VSS.t356 112.368
R2690 VSS.t439 VSS.t339 112.368
R2691 VSS.t468 VSS.t439 112.368
R2692 VSS.t345 VSS.t468 112.368
R2693 VSS.t394 VSS.t345 112.368
R2694 VSS.t435 VSS.t394 112.368
R2695 VSS.t392 VSS.t435 112.368
R2696 VSS.t358 VSS.t431 69.8719
R2697 VSS.t477 VSS.t358 69.8719
R2698 VSS.t412 VSS.t477 69.8719
R2699 VSS.t335 VSS.t310 69.8719
R2700 VSS.t360 VSS.t441 69.8719
R2701 VSS.t479 VSS.t360 69.8719
R2702 VSS.t414 VSS.t479 69.8719
R2703 VSS.t337 VSS.t316 69.8719
R2704 VSS.n769 VSS.t445 59.9648
R2705 VSS.n769 VSS.t319 59.9648
R2706 VSS.n1769 VSS.t404 59.9648
R2707 VSS.n1769 VSS.t333 59.9648
R2708 VSS.n759 VSS.t324 59.9648
R2709 VSS.n1675 VSS.t447 59.9648
R2710 VSS.n1675 VSS.t289 59.9648
R2711 VSS.n759 VSS.t410 59.9648
R2712 VSS.n496 VSS.t433 59.9648
R2713 VSS.n1641 VSS.t483 59.9648
R2714 VSS.n1641 VSS.t369 59.9648
R2715 VSS.n496 VSS.t292 59.9648
R2716 VSS.n486 VSS.t304 59.9648
R2717 VSS.n1545 VSS.t408 59.9648
R2718 VSS.n1545 VSS.t466 59.9648
R2719 VSS.n486 VSS.t402 59.9648
R2720 VSS.n81 VSS.t485 59.9648
R2721 VSS.n1511 VSS.t487 59.9648
R2722 VSS.n1511 VSS.t373 59.9648
R2723 VSS.n81 VSS.t387 59.9648
R2724 VSS.n71 VSS.t464 59.9648
R2725 VSS.n1415 VSS.t400 59.9648
R2726 VSS.n1415 VSS.t456 59.9648
R2727 VSS.n71 VSS.t349 59.9648
R2728 VSS.n2430 VSS.t351 55.1416
R2729 VSS.n2430 VSS.t396 55.1416
R2730 VSS.n2300 VSS.t423 55.1416
R2731 VSS.n2300 VSS.t451 55.1416
R2732 VSS.n3536 VSS.t481 55.1416
R2733 VSS.n3536 VSS.t322 55.1416
R2734 VSS.n3473 VSS.t392 55.1416
R2735 VSS.n3473 VSS.t416 55.1416
R2736 VSS.n2562 VSS.t364 40.5416
R2737 VSS.n3945 VSS.t443 40.5416
R2738 VSS.n3945 VSS.t307 40.4112
R2739 VSS.n2557 VSS.t472 36.5005
R2740 VSS.n3774 VSS.t412 33.8934
R2741 VSS.n3774 VSS.t335 33.8934
R2742 VSS.n2467 VSS.t414 33.8434
R2743 VSS.n2467 VSS.t337 33.8434
R2744 VSS.n2165 VSS.n2145 27.2287
R2745 VSS.n2561 VSS.n2560 20.8576
R2746 VSS.n2560 VSS.n2559 20.8576
R2747 VSS.n2559 VSS.n2558 20.8576
R2748 VSS.n2558 VSS.n2557 20.8576
R2749 VSS.n3222 VSS.t245 20.0254
R2750 VSS.n2605 VSS.t365 20.0254
R2751 VSS.n2505 VSS.t37 20.0254
R2752 VSS.n3942 VSS.t308 20.0254
R2753 VSS.t354 VSS.t326 19.5645
R2754 VSS.t367 VSS.t378 19.5645
R2755 VSS.t385 VSS.t398 19.5645
R2756 VSS.n2487 VSS.t25 18.3212
R2757 VSS.n2480 VSS.t287 18.3212
R2758 VSS.n4054 VSS.t622 18.3212
R2759 VSS.n2496 VSS.t281 17.8951
R2760 VSS.n3185 VSS.t30 17.469
R2761 VSS.n3260 VSS.t545 17.469
R2762 VSS.n2562 VSS.n2561 17.4684
R2763 VSS.n3146 VSS.n3145 17.043
R2764 VSS.t473 VSS.t61 17.043
R2765 VSS.n3796 VSS.t41 16.6169
R2766 VSS.n4084 VSS.t3 16.1029
R2767 VSS.n4064 VSS.t0 16.1029
R2768 VSS.n2621 VSS.t296 15.7648
R2769 VSS.n2561 VSS.t437 15.6434
R2770 VSS.n2557 VSS.t453 15.6434
R2771 VSS.n2558 VSS.t295 15.6434
R2772 VSS.n2559 VSS.t380 15.6434
R2773 VSS.n2560 VSS.t389 15.6434
R2774 VSS.n2456 VSS.t248 14.9527
R2775 VSS.n3396 VSS.t28 14.9527
R2776 VSS.n3831 VSS.t226 14.9127
R2777 VSS.n2505 VSS.t284 14.0605
R2778 VSS.n2502 VSS.t21 14.0605
R2779 VSS.t242 VSS.t277 14.0605
R2780 VSS.t224 VSS.t261 14.0605
R2781 VSS.n3805 VSS.t524 14.0605
R2782 VSS.n3814 VSS.t517 14.0605
R2783 VSS.n968 VSS.t87 13.7786
R2784 VSS.n986 VSS.t182 13.7786
R2785 VSS.n1151 VSS.t185 13.7786
R2786 VSS.n1169 VSS.t175 13.7786
R2787 VSS.n1334 VSS.t108 13.7786
R2788 VSS.n1352 VSS.t136 13.7786
R2789 VSS.n2480 VSS.t263 13.6345
R2790 VSS.n2695 VSS.t367 13.542
R2791 VSS.n2697 VSS.t342 13.542
R2792 VSS.n2675 VSS.t385 13.542
R2793 VSS.n2677 VSS.t375 13.542
R2794 VSS.n3197 VSS.t19 13.2084
R2795 VSS.n3274 VSS.t327 13.2084
R2796 VSS.n2515 VSS.t285 13.2084
R2797 VSS.n3834 VSS.t60 13.2084
R2798 VSS.n3273 VSS.t354 12.7007
R2799 VSS.n3384 VSS.t250 12.6524
R2800 VSS.n3387 VSS.t247 12.6524
R2801 VSS.n2624 VSS.t454 12.3563
R2802 VSS.t262 VSS.n2486 12.3563
R2803 VSS.n2483 VSS.t567 12.3563
R2804 VSS.t514 VSS.t199 11.9302
R2805 VSS.n3156 VSS.t343 10.652
R2806 VSS.n3232 VSS.t540 10.652
R2807 VSS.n3288 VSS.t376 10.652
R2808 VSS.n3959 VSS.t58 10.652
R2809 VSS.n2493 VSS.t280 10.226
R2810 VSS.n2519 VSS.t24 9.79992
R2811 VSS.n2490 VSS.t22 9.79992
R2812 VSS.n3793 VSS.t255 9.79992
R2813 VSS.n3828 VSS.t627 9.79992
R2814 VSS.n3799 VSS.t278 9.37386
R2815 VSS.n4087 VSS.t8 9.20187
R2816 VSS.n4061 VSS.t204 9.20187
R2817 VSS.n3818 VSS.t265 8.9478
R2818 VSS.n2425 VSS.t352 8.81848
R2819 VSS.n3421 VSS.t419 8.81848
R2820 VSS.n3175 VSS.t14 8.09568
R2821 VSS.n3251 VSS.t535 8.09568
R2822 VSS.n2609 VSS.t390 8.09568
R2823 VSS.n2621 VSS.t35 8.09568
R2824 VSS.n2499 VSS.t209 8.09568
R2825 VSS.n965 VSS.t100 7.87372
R2826 VSS.n989 VSS.t149 7.87372
R2827 VSS.n1148 VSS.t72 7.87372
R2828 VSS.n1172 VSS.t129 7.87372
R2829 VSS.n1331 VSS.t116 7.87372
R2830 VSS.n1355 VSS.t156 7.87372
R2831 VSS.n3808 VSS.t502 7.24355
R2832 VSS.n3808 VSS.t264 6.81749
R2833 VSS.n2441 VSS.t251 6.51814
R2834 VSS.n3411 VSS.t252 6.51814
R2835 VSS.t23 VSS.t317 6.39143
R2836 VSS.n3962 VSS.t625 6.39143
R2837 VSS.n2502 VSS.t260 5.96537
R2838 VSS.n3773 VSS.t312 5.8372
R2839 VSS.n2466 VSS.t318 5.8372
R2840 VSS.n3956 VSS.t514 5.5393
R2841 VSS.n4077 VSS.t49 5.36797
R2842 VSS.n4071 VSS.t206 5.36797
R2843 VSS.t517 VSS.t500 5.11324
R2844 VSS.n2555 VSS.t286 5.07024
R2845 VSS.n3012 VSS.t328 5.0182
R2846 VSS.n2866 VSS.t438 4.7885
R2847 VSS.n3840 VSS.t309 4.7885
R2848 VSS.n3948 VSS.t444 4.7885
R2849 VSS.n3773 VSS.t336 4.7885
R2850 VSS.n3777 VSS.t413 4.7885
R2851 VSS.n3778 VSS.t478 4.7885
R2852 VSS.n3779 VSS.t359 4.7885
R2853 VSS.n3780 VSS.t432 4.7885
R2854 VSS.n2473 VSS.t442 4.7885
R2855 VSS.n2472 VSS.t361 4.7885
R2856 VSS.n2471 VSS.t480 4.7885
R2857 VSS.n2470 VSS.t415 4.7885
R2858 VSS.n2466 VSS.t338 4.7885
R2859 VSS.n3017 VSS.n3016 4.78615
R2860 VSS.n3802 VSS.t224 4.68718
R2861 VSS.n974 VSS.t92 4.59321
R2862 VSS.n980 VSS.t78 4.59321
R2863 VSS.n1157 VSS.t89 4.59321
R2864 VSS.n1163 VSS.t113 4.59321
R2865 VSS.n1340 VSS.t140 4.59321
R2866 VSS.n1346 VSS.t103 4.59321
R2867 VSS.n2763 VSS.n2694 4.45746
R2868 VSS.n2778 VSS.n2692 4.45746
R2869 VSS.n1694 VSS.n1693 4.44992
R2870 VSS.n1714 VSS.n1713 4.44992
R2871 VSS.n1564 VSS.n1563 4.44992
R2872 VSS.n1584 VSS.n1583 4.44992
R2873 VSS.n1434 VSS.n1433 4.44992
R2874 VSS.n1454 VSS.n1453 4.44992
R2875 VSS.n2450 VSS.t27 4.21779
R2876 VSS.n3402 VSS.t249 4.21779
R2877 VSS.n3035 VSS.n3034 4.1992
R2878 VSS.n3040 VSS.n3039 4.1992
R2879 VSS.n2549 VSS.n2548 4.05833
R2880 VSS.n760 VSS.n759 4.0005
R2881 VSS.n1676 VSS.n1675 4.0005
R2882 VSS.n497 VSS.n496 4.0005
R2883 VSS.n1642 VSS.n1641 4.0005
R2884 VSS.n487 VSS.n486 4.0005
R2885 VSS.n1546 VSS.n1545 4.0005
R2886 VSS.n82 VSS.n81 4.0005
R2887 VSS.n1512 VSS.n1511 4.0005
R2888 VSS.n72 VSS.n71 4.0005
R2889 VSS.n1416 VSS.n1415 4.0005
R2890 VSS.n2301 VSS.n2300 4.0005
R2891 VSS.n3946 VSS.n3945 4.0005
R2892 VSS.n2563 VSS.n2562 4.0005
R2893 VSS.n3775 VSS.n3774 4.0005
R2894 VSS.n2468 VSS.n2467 4.0005
R2895 VSS.n3474 VSS.n3473 4.0005
R2896 VSS.n3537 VSS.n3536 4.0005
R2897 VSS.n2431 VSS.n2430 4.0005
R2898 VSS.n1770 VSS.n1769 4.0005
R2899 VSS.n770 VSS.n769 4.0005
R2900 VSS.n3012 VSS.t355 3.9695
R2901 VSS.n2682 VSS.t377 3.9695
R2902 VSS.n3008 VSS.t386 3.9695
R2903 VSS.n3009 VSS.t399 3.9695
R2904 VSS.n3207 VSS.t64 3.83506
R2905 VSS.n2615 VSS.t381 3.83506
R2906 VSS.n2493 VSS.t39 3.83506
R2907 VSS.n2941 VSS.n2867 3.75898
R2908 VSS.n2938 VSS.n2868 3.75898
R2909 VSS.n2933 VSS.n2869 3.75898
R2910 VSS.n2928 VSS.n2870 3.75898
R2911 VSS.n2892 VSS.n2872 3.75898
R2912 VSS.n2881 VSS.n2874 3.75898
R2913 VSS.n3850 VSS.n3847 3.75898
R2914 VSS.n3861 VSS.n3845 3.75898
R2915 VSS.n3870 VSS.n3843 3.75898
R2916 VSS.n2433 VSS.t397 3.71925
R2917 VSS.n2303 VSS.t452 3.71925
R2918 VSS.n2299 VSS.t424 3.71925
R2919 VSS.n2298 VSS.t471 3.71925
R2920 VSS.n0 VSS.t420 3.71925
R2921 VSS.n3539 VSS.t323 3.71925
R2922 VSS.n3535 VSS.t482 3.71925
R2923 VSS.n3534 VSS.t357 3.71925
R2924 VSS.n3533 VSS.t463 3.71925
R2925 VSS.n3532 VSS.t430 3.71925
R2926 VSS.n308 VSS.t372 3.71925
R2927 VSS.n309 VSS.t315 3.71925
R2928 VSS.n310 VSS.t426 3.71925
R2929 VSS.n3478 VSS.t393 3.71925
R2930 VSS.n3477 VSS.t436 3.71925
R2931 VSS.n3476 VSS.t395 3.71925
R2932 VSS.n3475 VSS.t346 3.71925
R2933 VSS.n245 VSS.t469 3.71925
R2934 VSS.n246 VSS.t440 3.71925
R2935 VSS.n247 VSS.t341 3.71925
R2936 VSS.n3480 VSS.t417 3.71925
R2937 VSS.n2429 VSS.t353 3.71925
R2938 VSS.n2428 VSS.t407 3.71925
R2939 VSS.n2 VSS.t363 3.71925
R2940 VSS.n768 VSS.t321 3.6965
R2941 VSS.n767 VSS.t461 3.6965
R2942 VSS.n1771 VSS.t459 3.6965
R2943 VSS.n1772 VSS.t405 3.6965
R2944 VSS.n1774 VSS.t334 3.6965
R2945 VSS.n1678 VSS.t448 3.6965
R2946 VSS.n758 VSS.t411 3.6965
R2947 VSS.n757 VSS.t348 3.6965
R2948 VSS.n1673 VSS.t384 3.6965
R2949 VSS.n1674 VSS.t291 3.6965
R2950 VSS.n762 VSS.t325 3.6965
R2951 VSS.n1644 VSS.t484 3.6965
R2952 VSS.n495 VSS.t294 3.6965
R2953 VSS.n494 VSS.t450 3.6965
R2954 VSS.n1639 VSS.t422 3.6965
R2955 VSS.n1640 VSS.t370 3.6965
R2956 VSS.n499 VSS.t434 3.6965
R2957 VSS.n1548 VSS.t409 3.6965
R2958 VSS.n485 VSS.t403 3.6965
R2959 VSS.n484 VSS.t332 3.6965
R2960 VSS.n1543 VSS.t330 3.6965
R2961 VSS.n1544 VSS.t467 3.6965
R2962 VSS.n489 VSS.t306 3.6965
R2963 VSS.n1514 VSS.t488 3.6965
R2964 VSS.n80 VSS.t388 3.6965
R2965 VSS.n79 VSS.t300 3.6965
R2966 VSS.n1509 VSS.t428 3.6965
R2967 VSS.n1510 VSS.t374 3.6965
R2968 VSS.n84 VSS.t486 3.6965
R2969 VSS.n1418 VSS.t401 3.6965
R2970 VSS.n70 VSS.t350 3.6965
R2971 VSS.n69 VSS.t476 3.6965
R2972 VSS.n1413 VSS.t303 3.6965
R2973 VSS.n1414 VSS.t457 3.6965
R2974 VSS.n74 VSS.t465 3.6965
R2975 VSS.n772 VSS.t446 3.6965
R2976 VSS.n2556 VSS.n2534 3.43224
R2977 VSS.n2554 VSS.n2536 3.43224
R2978 VSS.n2553 VSS.n2538 3.43224
R2979 VSS.n2552 VSS.n2540 3.43224
R2980 VSS.n2551 VSS.n2542 3.43224
R2981 VSS.n2550 VSS.n2544 3.43224
R2982 VSS.n2549 VSS.n2546 3.43224
R2983 VSS.n2864 VSS.n2862 3.31707
R2984 VSS.n2592 VSS.n2591 3.31707
R2985 VSS.n2670 VSS.n2669 3.31707
R2986 VSS.n2855 VSS.n2853 3.3165
R2987 VSS.n3329 VSS.n3327 3.3165
R2988 VSS.n3329 VSS.n3328 3.3165
R2989 VSS.n2640 VSS.n2638 3.3165
R2990 VSS.n2167 VSS.n2166 3.3165
R2991 VSS.n2665 VSS.n2663 3.3164
R2992 VSS.n2673 VSS.n2671 3.3164
R2993 VSS.n926 VSS.n897 3.31593
R2994 VSS.n2665 VSS.n2664 3.31583
R2995 VSS.n2673 VSS.n2672 3.31583
R2996 VSS.n1747 VSS.n1746 3.1505
R2997 VSS.n1748 VSS.n1742 3.1505
R2998 VSS.n1617 VSS.n1616 3.1505
R2999 VSS.n1618 VSS.n1612 3.1505
R3000 VSS.n1487 VSS.n1486 3.1505
R3001 VSS.n1488 VSS.n1482 3.1505
R3002 VSS.n3017 VSS.n3014 3.1505
R3003 VSS.n3018 VSS.n3013 3.1505
R3004 VSS.n3035 VSS.n3032 3.1505
R3005 VSS.n3040 VSS.n3037 3.1505
R3006 VSS.n3046 VSS.n3042 3.1505
R3007 VSS.n3045 VSS.n3044 3.1505
R3008 VSS.n2704 VSS.n2703 3.1505
R3009 VSS.n3030 VSS.n3026 3.1505
R3010 VSS.n3029 VSS.n3028 3.1505
R3011 VSS.n2690 VSS.n2689 3.1505
R3012 VSS.n3024 VSS.n3020 3.1505
R3013 VSS.n3023 VSS.n3022 3.1505
R3014 VSS.n2687 VSS.n2686 3.1505
R3015 VSS.n2566 VSS.n2532 3.1505
R3016 VSS.n2947 VSS.n2946 3.1505
R3017 VSS.n286 VSS.n279 3.1505
R3018 VSS.n285 VSS.n281 3.1505
R3019 VSS.n284 VSS.n283 3.1505
R3020 VSS.n3756 VSS.n3755 3.1505
R3021 VSS.n3759 VSS.n3758 3.1505
R3022 VSS.n3762 VSS.n3761 3.1505
R3023 VSS.n3765 VSS.n3764 3.1505
R3024 VSS.n3768 VSS.n3767 3.1505
R3025 VSS.n277 VSS.n270 3.1505
R3026 VSS.n276 VSS.n272 3.1505
R3027 VSS.n275 VSS.n274 3.1505
R3028 VSS.n3519 VSS.n3518 3.1505
R3029 VSS.n3522 VSS.n3521 3.1505
R3030 VSS.n3525 VSS.n3524 3.1505
R3031 VSS.n3528 VSS.n3527 3.1505
R3032 VSS.n3531 VSS.n3530 3.1505
R3033 VSS.n268 VSS.n261 3.1505
R3034 VSS.n267 VSS.n263 3.1505
R3035 VSS.n266 VSS.n265 3.1505
R3036 VSS.n3504 VSS.n3503 3.1505
R3037 VSS.n3507 VSS.n3506 3.1505
R3038 VSS.n3510 VSS.n3509 3.1505
R3039 VSS.n3513 VSS.n3512 3.1505
R3040 VSS.n3516 VSS.n3515 3.1505
R3041 VSS.n259 VSS.n252 3.1505
R3042 VSS.n258 VSS.n254 3.1505
R3043 VSS.n257 VSS.n256 3.1505
R3044 VSS.n3489 VSS.n3488 3.1505
R3045 VSS.n3492 VSS.n3491 3.1505
R3046 VSS.n3495 VSS.n3494 3.1505
R3047 VSS.n3498 VSS.n3497 3.1505
R3048 VSS.n3501 VSS.n3500 3.1505
R3049 VSS.n2640 VSS.n2639 3.06217
R3050 VSS.n1395 VSS.n1394 3.06217
R3051 VSS.n1240 VSS.n1239 3.06217
R3052 VSS.n1057 VSS.n1056 3.06217
R3053 VSS.n1292 VSS.n1244 3.0616
R3054 VSS.n1109 VSS.n1061 3.0616
R3055 VSS.n3324 VSS.n3323 3.01258
R3056 VSS.n3128 VSS.n3127 3.01207
R3057 VSS.n1292 VSS.n1291 3.01207
R3058 VSS.n1109 VSS.n1108 3.01207
R3059 VSS.n926 VSS.n925 3.01207
R3060 VSS.n2855 VSS.n2854 3.01202
R3061 VSS.n2592 VSS.n2590 3.01202
R3062 VSS.n1395 VSS.n1393 3.01202
R3063 VSS.n1240 VSS.n1238 3.01202
R3064 VSS.n1057 VSS.n1055 3.01202
R3065 VSS.n2864 VSS.n2863 3.0115
R3066 VSS.n3825 VSS.t258 2.98293
R3067 VSS.n1687 VSS.n1684 2.91104
R3068 VSS.n1707 VSS.n1704 2.91104
R3069 VSS.n1557 VSS.n1554 2.91104
R3070 VSS.n1577 VSS.n1574 2.91104
R3071 VSS.n1427 VSS.n1424 2.91104
R3072 VSS.n1447 VSS.n1444 2.91104
R3073 VSS.n1699 VSS.n1696 2.86846
R3074 VSS.n1719 VSS.n1716 2.86846
R3075 VSS.n1569 VSS.n1566 2.86846
R3076 VSS.n1589 VSS.n1586 2.86846
R3077 VSS.n1439 VSS.n1436 2.86846
R3078 VSS.n1459 VSS.n1456 2.86846
R3079 VSS.n1752 VSS.n1751 2.80979
R3080 VSS.n1622 VSS.n1621 2.80979
R3081 VSS.n1492 VSS.n1491 2.80979
R3082 VSS.n2714 VSS.n2713 2.75023
R3083 VSS.n2699 VSS.n2697 2.65431
R3084 VSS.n2679 VSS.n2677 2.65431
R3085 VSS.n896 VSS.n895 2.6005
R3086 VSS.n1865 VSS.n1864 2.6005
R3087 VSS.n1874 VSS.n1873 2.6005
R3088 VSS.n1943 VSS.n1942 2.6005
R3089 VSS.n1952 VSS.n1951 2.6005
R3090 VSS.n1411 VSS.n1410 2.6005
R3091 VSS.n1403 VSS.n1402 2.6005
R3092 VSS.n1406 VSS.n1405 2.6005
R3093 VSS.n1408 VSS.n1407 2.6005
R3094 VSS.n1400 VSS.n1399 2.6005
R3095 VSS.n1528 VSS.n1527 2.6005
R3096 VSS.n1526 VSS.n1525 2.6005
R3097 VSS.n1524 VSS.n1523 2.6005
R3098 VSS.n1522 VSS.n1521 2.6005
R3099 VSS.n1520 VSS.n1519 2.6005
R3100 VSS.n90 VSS.n89 2.6005
R3101 VSS.n92 VSS.n91 2.6005
R3102 VSS.n94 VSS.n93 2.6005
R3103 VSS.n96 VSS.n95 2.6005
R3104 VSS.n98 VSS.n97 2.6005
R3105 VSS.n100 VSS.n99 2.6005
R3106 VSS.n102 VSS.n101 2.6005
R3107 VSS.n104 VSS.n103 2.6005
R3108 VSS.n106 VSS.n105 2.6005
R3109 VSS.n108 VSS.n107 2.6005
R3110 VSS.n110 VSS.n109 2.6005
R3111 VSS.n112 VSS.n111 2.6005
R3112 VSS.n114 VSS.n113 2.6005
R3113 VSS.n116 VSS.n115 2.6005
R3114 VSS.n118 VSS.n117 2.6005
R3115 VSS.n120 VSS.n119 2.6005
R3116 VSS.n122 VSS.n121 2.6005
R3117 VSS.n124 VSS.n123 2.6005
R3118 VSS.n126 VSS.n125 2.6005
R3119 VSS.n128 VSS.n127 2.6005
R3120 VSS.n130 VSS.n129 2.6005
R3121 VSS.n132 VSS.n131 2.6005
R3122 VSS.n134 VSS.n133 2.6005
R3123 VSS.n136 VSS.n135 2.6005
R3124 VSS.n138 VSS.n137 2.6005
R3125 VSS.n140 VSS.n139 2.6005
R3126 VSS.n142 VSS.n141 2.6005
R3127 VSS.n144 VSS.n143 2.6005
R3128 VSS.n146 VSS.n145 2.6005
R3129 VSS.n148 VSS.n147 2.6005
R3130 VSS.n150 VSS.n149 2.6005
R3131 VSS.n152 VSS.n151 2.6005
R3132 VSS.n154 VSS.n153 2.6005
R3133 VSS.n156 VSS.n155 2.6005
R3134 VSS.n158 VSS.n157 2.6005
R3135 VSS.n160 VSS.n159 2.6005
R3136 VSS.n162 VSS.n161 2.6005
R3137 VSS.n164 VSS.n163 2.6005
R3138 VSS.n166 VSS.n165 2.6005
R3139 VSS.n169 VSS.n168 2.6005
R3140 VSS.n172 VSS.n171 2.6005
R3141 VSS.n175 VSS.n174 2.6005
R3142 VSS.n178 VSS.n177 2.6005
R3143 VSS.n181 VSS.n180 2.6005
R3144 VSS.n184 VSS.n183 2.6005
R3145 VSS.n187 VSS.n186 2.6005
R3146 VSS.n190 VSS.n189 2.6005
R3147 VSS.n193 VSS.n192 2.6005
R3148 VSS.n196 VSS.n195 2.6005
R3149 VSS.n199 VSS.n198 2.6005
R3150 VSS.n202 VSS.n201 2.6005
R3151 VSS.n205 VSS.n204 2.6005
R3152 VSS.n208 VSS.n207 2.6005
R3153 VSS.n211 VSS.n210 2.6005
R3154 VSS.n214 VSS.n213 2.6005
R3155 VSS.n217 VSS.n216 2.6005
R3156 VSS.n220 VSS.n219 2.6005
R3157 VSS.n1530 VSS.n1529 2.6005
R3158 VSS.n481 VSS.n480 2.6005
R3159 VSS.n478 VSS.n477 2.6005
R3160 VSS.n475 VSS.n474 2.6005
R3161 VSS.n473 VSS.n472 2.6005
R3162 VSS.n470 VSS.n469 2.6005
R3163 VSS.n468 VSS.n467 2.6005
R3164 VSS.n465 VSS.n464 2.6005
R3165 VSS.n463 VSS.n462 2.6005
R3166 VSS.n460 VSS.n459 2.6005
R3167 VSS.n458 VSS.n457 2.6005
R3168 VSS.n455 VSS.n454 2.6005
R3169 VSS.n453 VSS.n452 2.6005
R3170 VSS.n451 VSS.n450 2.6005
R3171 VSS.n449 VSS.n448 2.6005
R3172 VSS.n447 VSS.n446 2.6005
R3173 VSS.n445 VSS.n444 2.6005
R3174 VSS.n443 VSS.n442 2.6005
R3175 VSS.n441 VSS.n440 2.6005
R3176 VSS.n439 VSS.n438 2.6005
R3177 VSS.n437 VSS.n436 2.6005
R3178 VSS.n435 VSS.n434 2.6005
R3179 VSS.n433 VSS.n432 2.6005
R3180 VSS.n431 VSS.n430 2.6005
R3181 VSS.n429 VSS.n428 2.6005
R3182 VSS.n427 VSS.n426 2.6005
R3183 VSS.n425 VSS.n424 2.6005
R3184 VSS.n423 VSS.n422 2.6005
R3185 VSS.n421 VSS.n420 2.6005
R3186 VSS.n419 VSS.n418 2.6005
R3187 VSS.n417 VSS.n416 2.6005
R3188 VSS.n415 VSS.n414 2.6005
R3189 VSS.n413 VSS.n412 2.6005
R3190 VSS.n411 VSS.n410 2.6005
R3191 VSS.n409 VSS.n408 2.6005
R3192 VSS.n407 VSS.n406 2.6005
R3193 VSS.n405 VSS.n404 2.6005
R3194 VSS.n403 VSS.n402 2.6005
R3195 VSS.n401 VSS.n400 2.6005
R3196 VSS.n399 VSS.n398 2.6005
R3197 VSS.n397 VSS.n396 2.6005
R3198 VSS.n395 VSS.n394 2.6005
R3199 VSS.n393 VSS.n392 2.6005
R3200 VSS.n391 VSS.n390 2.6005
R3201 VSS.n389 VSS.n388 2.6005
R3202 VSS.n387 VSS.n386 2.6005
R3203 VSS.n385 VSS.n384 2.6005
R3204 VSS.n383 VSS.n382 2.6005
R3205 VSS.n381 VSS.n380 2.6005
R3206 VSS.n379 VSS.n378 2.6005
R3207 VSS.n377 VSS.n376 2.6005
R3208 VSS.n375 VSS.n374 2.6005
R3209 VSS.n373 VSS.n372 2.6005
R3210 VSS.n371 VSS.n370 2.6005
R3211 VSS.n369 VSS.n368 2.6005
R3212 VSS.n367 VSS.n366 2.6005
R3213 VSS.n365 VSS.n364 2.6005
R3214 VSS.n1532 VSS.n1531 2.6005
R3215 VSS.n1534 VSS.n1533 2.6005
R3216 VSS.n1536 VSS.n1535 2.6005
R3217 VSS.n1538 VSS.n1537 2.6005
R3218 VSS.n1540 VSS.n1539 2.6005
R3219 VSS.n1542 VSS.n1541 2.6005
R3220 VSS.n483 VSS.n482 2.6005
R3221 VSS.n1658 VSS.n1657 2.6005
R3222 VSS.n1656 VSS.n1655 2.6005
R3223 VSS.n1654 VSS.n1653 2.6005
R3224 VSS.n1652 VSS.n1651 2.6005
R3225 VSS.n1650 VSS.n1649 2.6005
R3226 VSS.n505 VSS.n504 2.6005
R3227 VSS.n507 VSS.n506 2.6005
R3228 VSS.n509 VSS.n508 2.6005
R3229 VSS.n511 VSS.n510 2.6005
R3230 VSS.n513 VSS.n512 2.6005
R3231 VSS.n515 VSS.n514 2.6005
R3232 VSS.n517 VSS.n516 2.6005
R3233 VSS.n519 VSS.n518 2.6005
R3234 VSS.n521 VSS.n520 2.6005
R3235 VSS.n523 VSS.n522 2.6005
R3236 VSS.n525 VSS.n524 2.6005
R3237 VSS.n527 VSS.n526 2.6005
R3238 VSS.n529 VSS.n528 2.6005
R3239 VSS.n531 VSS.n530 2.6005
R3240 VSS.n533 VSS.n532 2.6005
R3241 VSS.n535 VSS.n534 2.6005
R3242 VSS.n537 VSS.n536 2.6005
R3243 VSS.n539 VSS.n538 2.6005
R3244 VSS.n541 VSS.n540 2.6005
R3245 VSS.n543 VSS.n542 2.6005
R3246 VSS.n545 VSS.n544 2.6005
R3247 VSS.n547 VSS.n546 2.6005
R3248 VSS.n549 VSS.n548 2.6005
R3249 VSS.n551 VSS.n550 2.6005
R3250 VSS.n553 VSS.n552 2.6005
R3251 VSS.n555 VSS.n554 2.6005
R3252 VSS.n557 VSS.n556 2.6005
R3253 VSS.n559 VSS.n558 2.6005
R3254 VSS.n561 VSS.n560 2.6005
R3255 VSS.n563 VSS.n562 2.6005
R3256 VSS.n565 VSS.n564 2.6005
R3257 VSS.n567 VSS.n566 2.6005
R3258 VSS.n569 VSS.n568 2.6005
R3259 VSS.n571 VSS.n570 2.6005
R3260 VSS.n573 VSS.n572 2.6005
R3261 VSS.n575 VSS.n574 2.6005
R3262 VSS.n577 VSS.n576 2.6005
R3263 VSS.n579 VSS.n578 2.6005
R3264 VSS.n581 VSS.n580 2.6005
R3265 VSS.n584 VSS.n583 2.6005
R3266 VSS.n587 VSS.n586 2.6005
R3267 VSS.n590 VSS.n589 2.6005
R3268 VSS.n593 VSS.n592 2.6005
R3269 VSS.n596 VSS.n595 2.6005
R3270 VSS.n599 VSS.n598 2.6005
R3271 VSS.n602 VSS.n601 2.6005
R3272 VSS.n605 VSS.n604 2.6005
R3273 VSS.n608 VSS.n607 2.6005
R3274 VSS.n611 VSS.n610 2.6005
R3275 VSS.n614 VSS.n613 2.6005
R3276 VSS.n617 VSS.n616 2.6005
R3277 VSS.n620 VSS.n619 2.6005
R3278 VSS.n623 VSS.n622 2.6005
R3279 VSS.n626 VSS.n625 2.6005
R3280 VSS.n629 VSS.n628 2.6005
R3281 VSS.n632 VSS.n631 2.6005
R3282 VSS.n635 VSS.n634 2.6005
R3283 VSS.n1660 VSS.n1659 2.6005
R3284 VSS.n754 VSS.n753 2.6005
R3285 VSS.n751 VSS.n750 2.6005
R3286 VSS.n748 VSS.n747 2.6005
R3287 VSS.n746 VSS.n745 2.6005
R3288 VSS.n743 VSS.n742 2.6005
R3289 VSS.n741 VSS.n740 2.6005
R3290 VSS.n738 VSS.n737 2.6005
R3291 VSS.n736 VSS.n735 2.6005
R3292 VSS.n733 VSS.n732 2.6005
R3293 VSS.n731 VSS.n730 2.6005
R3294 VSS.n728 VSS.n727 2.6005
R3295 VSS.n726 VSS.n725 2.6005
R3296 VSS.n724 VSS.n723 2.6005
R3297 VSS.n722 VSS.n721 2.6005
R3298 VSS.n720 VSS.n719 2.6005
R3299 VSS.n718 VSS.n717 2.6005
R3300 VSS.n716 VSS.n715 2.6005
R3301 VSS.n714 VSS.n713 2.6005
R3302 VSS.n712 VSS.n711 2.6005
R3303 VSS.n710 VSS.n709 2.6005
R3304 VSS.n708 VSS.n707 2.6005
R3305 VSS.n706 VSS.n705 2.6005
R3306 VSS.n704 VSS.n703 2.6005
R3307 VSS.n702 VSS.n701 2.6005
R3308 VSS.n700 VSS.n699 2.6005
R3309 VSS.n698 VSS.n697 2.6005
R3310 VSS.n696 VSS.n695 2.6005
R3311 VSS.n694 VSS.n693 2.6005
R3312 VSS.n692 VSS.n691 2.6005
R3313 VSS.n690 VSS.n689 2.6005
R3314 VSS.n688 VSS.n687 2.6005
R3315 VSS.n686 VSS.n685 2.6005
R3316 VSS.n684 VSS.n683 2.6005
R3317 VSS.n682 VSS.n681 2.6005
R3318 VSS.n680 VSS.n679 2.6005
R3319 VSS.n678 VSS.n677 2.6005
R3320 VSS.n676 VSS.n675 2.6005
R3321 VSS.n674 VSS.n673 2.6005
R3322 VSS.n672 VSS.n671 2.6005
R3323 VSS.n670 VSS.n669 2.6005
R3324 VSS.n668 VSS.n667 2.6005
R3325 VSS.n666 VSS.n665 2.6005
R3326 VSS.n664 VSS.n663 2.6005
R3327 VSS.n662 VSS.n661 2.6005
R3328 VSS.n660 VSS.n659 2.6005
R3329 VSS.n658 VSS.n657 2.6005
R3330 VSS.n656 VSS.n655 2.6005
R3331 VSS.n654 VSS.n653 2.6005
R3332 VSS.n652 VSS.n651 2.6005
R3333 VSS.n650 VSS.n649 2.6005
R3334 VSS.n648 VSS.n647 2.6005
R3335 VSS.n646 VSS.n645 2.6005
R3336 VSS.n644 VSS.n643 2.6005
R3337 VSS.n642 VSS.n641 2.6005
R3338 VSS.n640 VSS.n639 2.6005
R3339 VSS.n638 VSS.n637 2.6005
R3340 VSS.n1662 VSS.n1661 2.6005
R3341 VSS.n1664 VSS.n1663 2.6005
R3342 VSS.n1666 VSS.n1665 2.6005
R3343 VSS.n1668 VSS.n1667 2.6005
R3344 VSS.n1670 VSS.n1669 2.6005
R3345 VSS.n1672 VSS.n1671 2.6005
R3346 VSS.n756 VSS.n755 2.6005
R3347 VSS.n894 VSS.n893 2.6005
R3348 VSS.n891 VSS.n890 2.6005
R3349 VSS.n889 VSS.n888 2.6005
R3350 VSS.n886 VSS.n885 2.6005
R3351 VSS.n884 VSS.n883 2.6005
R3352 VSS.n881 VSS.n880 2.6005
R3353 VSS.n879 VSS.n878 2.6005
R3354 VSS.n876 VSS.n875 2.6005
R3355 VSS.n874 VSS.n873 2.6005
R3356 VSS.n871 VSS.n870 2.6005
R3357 VSS.n869 VSS.n868 2.6005
R3358 VSS.n866 VSS.n865 2.6005
R3359 VSS.n864 VSS.n863 2.6005
R3360 VSS.n862 VSS.n861 2.6005
R3361 VSS.n860 VSS.n859 2.6005
R3362 VSS.n858 VSS.n857 2.6005
R3363 VSS.n856 VSS.n855 2.6005
R3364 VSS.n854 VSS.n853 2.6005
R3365 VSS.n852 VSS.n851 2.6005
R3366 VSS.n850 VSS.n849 2.6005
R3367 VSS.n848 VSS.n847 2.6005
R3368 VSS.n846 VSS.n845 2.6005
R3369 VSS.n844 VSS.n843 2.6005
R3370 VSS.n842 VSS.n841 2.6005
R3371 VSS.n840 VSS.n839 2.6005
R3372 VSS.n838 VSS.n837 2.6005
R3373 VSS.n836 VSS.n835 2.6005
R3374 VSS.n834 VSS.n833 2.6005
R3375 VSS.n832 VSS.n831 2.6005
R3376 VSS.n830 VSS.n829 2.6005
R3377 VSS.n828 VSS.n827 2.6005
R3378 VSS.n826 VSS.n825 2.6005
R3379 VSS.n824 VSS.n823 2.6005
R3380 VSS.n822 VSS.n821 2.6005
R3381 VSS.n820 VSS.n819 2.6005
R3382 VSS.n818 VSS.n817 2.6005
R3383 VSS.n816 VSS.n815 2.6005
R3384 VSS.n814 VSS.n813 2.6005
R3385 VSS.n812 VSS.n811 2.6005
R3386 VSS.n810 VSS.n809 2.6005
R3387 VSS.n808 VSS.n807 2.6005
R3388 VSS.n806 VSS.n805 2.6005
R3389 VSS.n804 VSS.n803 2.6005
R3390 VSS.n802 VSS.n801 2.6005
R3391 VSS.n800 VSS.n799 2.6005
R3392 VSS.n798 VSS.n797 2.6005
R3393 VSS.n796 VSS.n795 2.6005
R3394 VSS.n794 VSS.n793 2.6005
R3395 VSS.n792 VSS.n791 2.6005
R3396 VSS.n790 VSS.n789 2.6005
R3397 VSS.n788 VSS.n787 2.6005
R3398 VSS.n786 VSS.n785 2.6005
R3399 VSS.n784 VSS.n783 2.6005
R3400 VSS.n782 VSS.n781 2.6005
R3401 VSS.n780 VSS.n779 2.6005
R3402 VSS.n778 VSS.n777 2.6005
R3403 VSS.n1776 VSS.n1775 2.6005
R3404 VSS.n1778 VSS.n1777 2.6005
R3405 VSS.n1780 VSS.n1779 2.6005
R3406 VSS.n1782 VSS.n1781 2.6005
R3407 VSS.n1784 VSS.n1783 2.6005
R3408 VSS.n1786 VSS.n1785 2.6005
R3409 VSS.n1792 VSS.n1787 2.6005
R3410 VSS.n3144 VSS.n3143 2.6005
R3411 VSS.n3125 VSS.n3124 2.6005
R3412 VSS.n2711 VSS.n2710 2.6005
R3413 VSS.n2708 VSS.n2707 2.6005
R3414 VSS.n2724 VSS.n2723 2.6005
R3415 VSS.n2723 VSS.n2722 2.6005
R3416 VSS.n2721 VSS.n2720 2.6005
R3417 VSS.n2720 VSS.n2719 2.6005
R3418 VSS.n2718 VSS.n2717 2.6005
R3419 VSS.n2717 VSS.n2716 2.6005
R3420 VSS.n3051 VSS.n3050 2.6005
R3421 VSS.n3050 VSS.n3049 2.6005
R3422 VSS.n3054 VSS.n3053 2.6005
R3423 VSS.n3053 VSS.n3052 2.6005
R3424 VSS.n3057 VSS.n3056 2.6005
R3425 VSS.n3056 VSS.n3055 2.6005
R3426 VSS.n3060 VSS.n3059 2.6005
R3427 VSS.n3059 VSS.n3058 2.6005
R3428 VSS.n3063 VSS.n3062 2.6005
R3429 VSS.n3062 VSS.n3061 2.6005
R3430 VSS.n3066 VSS.n3065 2.6005
R3431 VSS.n3065 VSS.n3064 2.6005
R3432 VSS.n3069 VSS.n3068 2.6005
R3433 VSS.n3068 VSS.n3067 2.6005
R3434 VSS.n3072 VSS.n3071 2.6005
R3435 VSS.n3071 VSS.n3070 2.6005
R3436 VSS.n3075 VSS.n3074 2.6005
R3437 VSS.n3074 VSS.n3073 2.6005
R3438 VSS.n3078 VSS.n3077 2.6005
R3439 VSS.n3077 VSS.n3076 2.6005
R3440 VSS.n3081 VSS.n3080 2.6005
R3441 VSS.n3080 VSS.n3079 2.6005
R3442 VSS.n3084 VSS.n3083 2.6005
R3443 VSS.n3083 VSS.n3082 2.6005
R3444 VSS.n3087 VSS.n3086 2.6005
R3445 VSS.n3086 VSS.n3085 2.6005
R3446 VSS.n3090 VSS.n3089 2.6005
R3447 VSS.n3089 VSS.n3088 2.6005
R3448 VSS.n3093 VSS.n3092 2.6005
R3449 VSS.n3092 VSS.n3091 2.6005
R3450 VSS.n3096 VSS.n3095 2.6005
R3451 VSS.n3095 VSS.n3094 2.6005
R3452 VSS.n3099 VSS.n3098 2.6005
R3453 VSS.n3098 VSS.n3097 2.6005
R3454 VSS.n3102 VSS.n3101 2.6005
R3455 VSS.n3101 VSS.n3100 2.6005
R3456 VSS.n3105 VSS.n3104 2.6005
R3457 VSS.n3104 VSS.n3103 2.6005
R3458 VSS.n3108 VSS.n3107 2.6005
R3459 VSS.n3107 VSS.n3106 2.6005
R3460 VSS.n3111 VSS.n3110 2.6005
R3461 VSS.n3110 VSS.n3109 2.6005
R3462 VSS.n3114 VSS.n3113 2.6005
R3463 VSS.n3113 VSS.n3112 2.6005
R3464 VSS.n3117 VSS.n3116 2.6005
R3465 VSS.n3116 VSS.n3115 2.6005
R3466 VSS.n3120 VSS.n3119 2.6005
R3467 VSS.n3119 VSS.n3118 2.6005
R3468 VSS.n3123 VSS.n3122 2.6005
R3469 VSS.n3122 VSS.n3121 2.6005
R3470 VSS.n3131 VSS.n3130 2.6005
R3471 VSS.n3130 VSS.n3129 2.6005
R3472 VSS.n3134 VSS.n3133 2.6005
R3473 VSS.n3136 VSS.n3135 2.6005
R3474 VSS.n3139 VSS.n3138 2.6005
R3475 VSS.n3141 VSS.n3140 2.6005
R3476 VSS.n2738 VSS.n2737 2.6005
R3477 VSS.n2735 VSS.n2734 2.6005
R3478 VSS.n2732 VSS.n2731 2.6005
R3479 VSS.n2730 VSS.n2729 2.6005
R3480 VSS.n2727 VSS.n2726 2.6005
R3481 VSS.n2315 VSS.n2314 2.6005
R3482 VSS.n3557 VSS.n3556 2.6005
R3483 VSS.n3559 VSS.n3558 2.6005
R3484 VSS.n3561 VSS.n3560 2.6005
R3485 VSS.n3563 VSS.n3562 2.6005
R3486 VSS.n3565 VSS.n3564 2.6005
R3487 VSS.n3567 VSS.n3566 2.6005
R3488 VSS.n3569 VSS.n3568 2.6005
R3489 VSS.n3571 VSS.n3570 2.6005
R3490 VSS.n3573 VSS.n3572 2.6005
R3491 VSS.n3575 VSS.n3574 2.6005
R3492 VSS.n3577 VSS.n3576 2.6005
R3493 VSS.n3579 VSS.n3578 2.6005
R3494 VSS.n3581 VSS.n3580 2.6005
R3495 VSS.n3583 VSS.n3582 2.6005
R3496 VSS.n3585 VSS.n3584 2.6005
R3497 VSS.n3587 VSS.n3586 2.6005
R3498 VSS.n3589 VSS.n3588 2.6005
R3499 VSS.n3591 VSS.n3590 2.6005
R3500 VSS.n3593 VSS.n3592 2.6005
R3501 VSS.n3595 VSS.n3594 2.6005
R3502 VSS.n3597 VSS.n3596 2.6005
R3503 VSS.n3599 VSS.n3598 2.6005
R3504 VSS.n3601 VSS.n3600 2.6005
R3505 VSS.n3603 VSS.n3602 2.6005
R3506 VSS.n3605 VSS.n3604 2.6005
R3507 VSS.n3607 VSS.n3606 2.6005
R3508 VSS.n3609 VSS.n3608 2.6005
R3509 VSS.n3611 VSS.n3610 2.6005
R3510 VSS.n3613 VSS.n3612 2.6005
R3511 VSS.n3615 VSS.n3614 2.6005
R3512 VSS.n3617 VSS.n3616 2.6005
R3513 VSS.n3619 VSS.n3618 2.6005
R3514 VSS.n3621 VSS.n3620 2.6005
R3515 VSS.n3623 VSS.n3622 2.6005
R3516 VSS.n3625 VSS.n3624 2.6005
R3517 VSS.n3627 VSS.n3626 2.6005
R3518 VSS.n3629 VSS.n3628 2.6005
R3519 VSS.n3631 VSS.n3630 2.6005
R3520 VSS.n3633 VSS.n3632 2.6005
R3521 VSS.n3635 VSS.n3634 2.6005
R3522 VSS.n3637 VSS.n3636 2.6005
R3523 VSS.n3639 VSS.n3638 2.6005
R3524 VSS.n3641 VSS.n3640 2.6005
R3525 VSS.n3643 VSS.n3642 2.6005
R3526 VSS.n3646 VSS.n3645 2.6005
R3527 VSS.n3648 VSS.n3647 2.6005
R3528 VSS.n3651 VSS.n3650 2.6005
R3529 VSS.n3653 VSS.n3652 2.6005
R3530 VSS.n3656 VSS.n3655 2.6005
R3531 VSS.n3658 VSS.n3657 2.6005
R3532 VSS.n3661 VSS.n3660 2.6005
R3533 VSS.n3663 VSS.n3662 2.6005
R3534 VSS.n3666 VSS.n3665 2.6005
R3535 VSS.n3668 VSS.n3667 2.6005
R3536 VSS.n3671 VSS.n3670 2.6005
R3537 VSS.n3673 VSS.n3672 2.6005
R3538 VSS.n3730 VSS.n3729 2.6005
R3539 VSS.n2317 VSS.n2316 2.6005
R3540 VSS.n2319 VSS.n2318 2.6005
R3541 VSS.n2321 VSS.n2320 2.6005
R3542 VSS.n2323 VSS.n2322 2.6005
R3543 VSS.n2325 VSS.n2324 2.6005
R3544 VSS.n2327 VSS.n2326 2.6005
R3545 VSS.n2329 VSS.n2328 2.6005
R3546 VSS.n2331 VSS.n2330 2.6005
R3547 VSS.n2333 VSS.n2332 2.6005
R3548 VSS.n2335 VSS.n2334 2.6005
R3549 VSS.n2337 VSS.n2336 2.6005
R3550 VSS.n2339 VSS.n2338 2.6005
R3551 VSS.n2341 VSS.n2340 2.6005
R3552 VSS.n2343 VSS.n2342 2.6005
R3553 VSS.n2345 VSS.n2344 2.6005
R3554 VSS.n2347 VSS.n2346 2.6005
R3555 VSS.n2349 VSS.n2348 2.6005
R3556 VSS.n2351 VSS.n2350 2.6005
R3557 VSS.n2353 VSS.n2352 2.6005
R3558 VSS.n2355 VSS.n2354 2.6005
R3559 VSS.n2357 VSS.n2356 2.6005
R3560 VSS.n2359 VSS.n2358 2.6005
R3561 VSS.n2361 VSS.n2360 2.6005
R3562 VSS.n2363 VSS.n2362 2.6005
R3563 VSS.n2365 VSS.n2364 2.6005
R3564 VSS.n2367 VSS.n2366 2.6005
R3565 VSS.n2369 VSS.n2368 2.6005
R3566 VSS.n2371 VSS.n2370 2.6005
R3567 VSS.n2373 VSS.n2372 2.6005
R3568 VSS.n2376 VSS.n2375 2.6005
R3569 VSS.n2378 VSS.n2377 2.6005
R3570 VSS.n2381 VSS.n2380 2.6005
R3571 VSS.n2383 VSS.n2382 2.6005
R3572 VSS.n2386 VSS.n2385 2.6005
R3573 VSS.n2388 VSS.n2387 2.6005
R3574 VSS.n2391 VSS.n2390 2.6005
R3575 VSS.n2393 VSS.n2392 2.6005
R3576 VSS.n2396 VSS.n2395 2.6005
R3577 VSS.n2398 VSS.n2397 2.6005
R3578 VSS.n3892 VSS.n3891 2.6005
R3579 VSS.n2958 VSS.n2865 2.6005
R3580 VSS.n3927 VSS.n3926 2.6005
R3581 VSS.n3925 VSS.n3924 2.6005
R3582 VSS.n3922 VSS.n3921 2.6005
R3583 VSS.n3920 VSS.n3919 2.6005
R3584 VSS.n3917 VSS.n3916 2.6005
R3585 VSS.n3915 VSS.n3914 2.6005
R3586 VSS.n3912 VSS.n3911 2.6005
R3587 VSS.n3910 VSS.n3909 2.6005
R3588 VSS.n3907 VSS.n3906 2.6005
R3589 VSS.n3905 VSS.n3904 2.6005
R3590 VSS.n3902 VSS.n3901 2.6005
R3591 VSS.n3900 VSS.n3899 2.6005
R3592 VSS.n3897 VSS.n3896 2.6005
R3593 VSS.n3895 VSS.n3894 2.6005
R3594 VSS.n2587 VSS.n2586 2.6005
R3595 VSS.n2981 VSS.n2980 2.6005
R3596 VSS.n2979 VSS.n2978 2.6005
R3597 VSS.n2977 VSS.n2976 2.6005
R3598 VSS.n2975 VSS.n2974 2.6005
R3599 VSS.n2973 VSS.n2972 2.6005
R3600 VSS.n2971 VSS.n2970 2.6005
R3601 VSS.n2969 VSS.n2968 2.6005
R3602 VSS.n2967 VSS.n2966 2.6005
R3603 VSS.n2965 VSS.n2964 2.6005
R3604 VSS.n2963 VSS.n2962 2.6005
R3605 VSS.n3148 VSS.n3147 2.6005
R3606 VSS.n3147 VSS.n3146 2.6005
R3607 VSS.n3151 VSS.n3150 2.6005
R3608 VSS.n3150 VSS.n3149 2.6005
R3609 VSS.n3155 VSS.n3154 2.6005
R3610 VSS.n3154 VSS.n3153 2.6005
R3611 VSS.n3158 VSS.n3157 2.6005
R3612 VSS.n3157 VSS.n3156 2.6005
R3613 VSS.n3161 VSS.n3160 2.6005
R3614 VSS.n3160 VSS.n3159 2.6005
R3615 VSS.n3165 VSS.n3164 2.6005
R3616 VSS.n3164 VSS.n3163 2.6005
R3617 VSS.n3168 VSS.n3167 2.6005
R3618 VSS.n3167 VSS.n3166 2.6005
R3619 VSS.n3171 VSS.n3170 2.6005
R3620 VSS.n3170 VSS.n3169 2.6005
R3621 VSS.n3174 VSS.n3173 2.6005
R3622 VSS.n3173 VSS.n3172 2.6005
R3623 VSS.n3177 VSS.n3176 2.6005
R3624 VSS.n3176 VSS.n3175 2.6005
R3625 VSS.n3180 VSS.n3179 2.6005
R3626 VSS.n3179 VSS.n3178 2.6005
R3627 VSS.n3184 VSS.n3183 2.6005
R3628 VSS.n3183 VSS.n3182 2.6005
R3629 VSS.n3187 VSS.n3186 2.6005
R3630 VSS.n3186 VSS.n3185 2.6005
R3631 VSS.n3190 VSS.n3189 2.6005
R3632 VSS.n3189 VSS.n3188 2.6005
R3633 VSS.n3193 VSS.n3192 2.6005
R3634 VSS.n3192 VSS.n3191 2.6005
R3635 VSS.n3196 VSS.n3195 2.6005
R3636 VSS.n3195 VSS.n3194 2.6005
R3637 VSS.n3199 VSS.n3198 2.6005
R3638 VSS.n3198 VSS.n3197 2.6005
R3639 VSS.n3202 VSS.n3201 2.6005
R3640 VSS.n3201 VSS.n3200 2.6005
R3641 VSS.n3206 VSS.n3205 2.6005
R3642 VSS.n3205 VSS.n3204 2.6005
R3643 VSS.n3209 VSS.n3208 2.6005
R3644 VSS.n3208 VSS.n3207 2.6005
R3645 VSS.n3212 VSS.n3211 2.6005
R3646 VSS.n3211 VSS.n3210 2.6005
R3647 VSS.n3215 VSS.n3214 2.6005
R3648 VSS.n3214 VSS.n3213 2.6005
R3649 VSS.n3218 VSS.n3217 2.6005
R3650 VSS.n3217 VSS.n3216 2.6005
R3651 VSS.n3221 VSS.n3220 2.6005
R3652 VSS.n3220 VSS.n3219 2.6005
R3653 VSS.n3224 VSS.n3223 2.6005
R3654 VSS.n3223 VSS.n3222 2.6005
R3655 VSS.n3227 VSS.n3226 2.6005
R3656 VSS.n3226 VSS.n3225 2.6005
R3657 VSS.n3231 VSS.n3230 2.6005
R3658 VSS.n3230 VSS.n3229 2.6005
R3659 VSS.n3234 VSS.n3233 2.6005
R3660 VSS.n3233 VSS.n3232 2.6005
R3661 VSS.n3237 VSS.n3236 2.6005
R3662 VSS.n3236 VSS.n3235 2.6005
R3663 VSS.n3240 VSS.n3239 2.6005
R3664 VSS.n3239 VSS.n3238 2.6005
R3665 VSS.n3243 VSS.n3242 2.6005
R3666 VSS.n3242 VSS.n3241 2.6005
R3667 VSS.n3246 VSS.n3245 2.6005
R3668 VSS.n3245 VSS.n3244 2.6005
R3669 VSS.n3250 VSS.n3249 2.6005
R3670 VSS.n3249 VSS.n3248 2.6005
R3671 VSS.n3253 VSS.n3252 2.6005
R3672 VSS.n3252 VSS.n3251 2.6005
R3673 VSS.n3256 VSS.n3255 2.6005
R3674 VSS.n3255 VSS.n3254 2.6005
R3675 VSS.n3259 VSS.n3258 2.6005
R3676 VSS.n3258 VSS.n3257 2.6005
R3677 VSS.n3262 VSS.n3261 2.6005
R3678 VSS.n3261 VSS.n3260 2.6005
R3679 VSS.n3265 VSS.n3264 2.6005
R3680 VSS.n3264 VSS.n3263 2.6005
R3681 VSS.n3268 VSS.n3267 2.6005
R3682 VSS.n3267 VSS.n3266 2.6005
R3683 VSS.n3272 VSS.n3271 2.6005
R3684 VSS.n3271 VSS.n3270 2.6005
R3685 VSS.n3276 VSS.n3275 2.6005
R3686 VSS.n3275 VSS.n3274 2.6005
R3687 VSS.n3279 VSS.n3278 2.6005
R3688 VSS.n3278 VSS.n3277 2.6005
R3689 VSS.n3283 VSS.n3282 2.6005
R3690 VSS.n3282 VSS.n3281 2.6005
R3691 VSS.n3287 VSS.n3286 2.6005
R3692 VSS.n3286 VSS.n3285 2.6005
R3693 VSS.n3290 VSS.n3289 2.6005
R3694 VSS.n3289 VSS.n3288 2.6005
R3695 VSS.n3293 VSS.n3292 2.6005
R3696 VSS.n3292 VSS.n3291 2.6005
R3697 VSS.n3297 VSS.n3296 2.6005
R3698 VSS.n3296 VSS.n3295 2.6005
R3699 VSS.n3300 VSS.n3299 2.6005
R3700 VSS.n3299 VSS.n3298 2.6005
R3701 VSS.n3303 VSS.n3302 2.6005
R3702 VSS.n3302 VSS.n3301 2.6005
R3703 VSS.n3306 VSS.n3305 2.6005
R3704 VSS.n3305 VSS.n3304 2.6005
R3705 VSS.n3309 VSS.n3308 2.6005
R3706 VSS.n3308 VSS.n3307 2.6005
R3707 VSS.n3312 VSS.n3311 2.6005
R3708 VSS.n3311 VSS.n3310 2.6005
R3709 VSS.n3315 VSS.n3314 2.6005
R3710 VSS.n3314 VSS.n3313 2.6005
R3711 VSS.n3326 VSS.n3325 2.6005
R3712 VSS.n2992 VSS.n2991 2.6005
R3713 VSS.n2995 VSS.n2994 2.6005
R3714 VSS.n2997 VSS.n2996 2.6005
R3715 VSS.n3000 VSS.n2999 2.6005
R3716 VSS.n3002 VSS.n3001 2.6005
R3717 VSS.n3005 VSS.n3004 2.6005
R3718 VSS.n3007 VSS.n3006 2.6005
R3719 VSS.n2668 VSS.n2666 2.6005
R3720 VSS.n2989 VSS.n2988 2.6005
R3721 VSS.n2986 VSS.n2985 2.6005
R3722 VSS.n2984 VSS.n2983 2.6005
R3723 VSS.n2668 VSS.n2667 2.6005
R3724 VSS.n2960 VSS.n2959 2.6005
R3725 VSS.n2852 VSS.n2851 2.6005
R3726 VSS.n2850 VSS.n2849 2.6005
R3727 VSS.n2848 VSS.n2847 2.6005
R3728 VSS.n2846 VSS.n2845 2.6005
R3729 VSS.n2844 VSS.n2843 2.6005
R3730 VSS.n2842 VSS.n2841 2.6005
R3731 VSS.n2840 VSS.n2839 2.6005
R3732 VSS.n2837 VSS.n2836 2.6005
R3733 VSS.n2835 VSS.n2834 2.6005
R3734 VSS.n2833 VSS.n2832 2.6005
R3735 VSS.n2830 VSS.n2829 2.6005
R3736 VSS.n2828 VSS.n2827 2.6005
R3737 VSS.n2826 VSS.n2825 2.6005
R3738 VSS.n2824 VSS.n2823 2.6005
R3739 VSS.n2822 VSS.n2821 2.6005
R3740 VSS.n2820 VSS.n2819 2.6005
R3741 VSS.n2818 VSS.n2817 2.6005
R3742 VSS.n2816 VSS.n2815 2.6005
R3743 VSS.n2814 VSS.n2813 2.6005
R3744 VSS.n2812 VSS.n2811 2.6005
R3745 VSS.n2810 VSS.n2809 2.6005
R3746 VSS.n2807 VSS.n2806 2.6005
R3747 VSS.n2805 VSS.n2804 2.6005
R3748 VSS.n2803 VSS.n2802 2.6005
R3749 VSS.n2801 VSS.n2800 2.6005
R3750 VSS.n2799 VSS.n2798 2.6005
R3751 VSS.n2797 VSS.n2796 2.6005
R3752 VSS.n2794 VSS.n2793 2.6005
R3753 VSS.n2792 VSS.n2791 2.6005
R3754 VSS.n2790 VSS.n2789 2.6005
R3755 VSS.n2788 VSS.n2787 2.6005
R3756 VSS.n2786 VSS.n2785 2.6005
R3757 VSS.n2784 VSS.n2783 2.6005
R3758 VSS.n2782 VSS.n2781 2.6005
R3759 VSS.n2780 VSS.n2779 2.6005
R3760 VSS.n2777 VSS.n2776 2.6005
R3761 VSS.n2775 VSS.n2774 2.6005
R3762 VSS.n2773 VSS.n2772 2.6005
R3763 VSS.n2771 VSS.n2770 2.6005
R3764 VSS.n2769 VSS.n2768 2.6005
R3765 VSS.n2767 VSS.n2766 2.6005
R3766 VSS.n2765 VSS.n2764 2.6005
R3767 VSS.n2762 VSS.n2761 2.6005
R3768 VSS.n2760 VSS.n2759 2.6005
R3769 VSS.n2758 VSS.n2757 2.6005
R3770 VSS.n2756 VSS.n2755 2.6005
R3771 VSS.n2754 VSS.n2753 2.6005
R3772 VSS.n2752 VSS.n2751 2.6005
R3773 VSS.n2749 VSS.n2748 2.6005
R3774 VSS.n2747 VSS.n2746 2.6005
R3775 VSS.n2745 VSS.n2744 2.6005
R3776 VSS.n2742 VSS.n2741 2.6005
R3777 VSS.n2740 VSS.n2739 2.6005
R3778 VSS.n2585 VSS.n2584 2.6005
R3779 VSS.n2582 VSS.n2581 2.6005
R3780 VSS.n2580 VSS.n2579 2.6005
R3781 VSS.n2577 VSS.n2576 2.6005
R3782 VSS.n2575 VSS.n2574 2.6005
R3783 VSS.n2572 VSS.n2571 2.6005
R3784 VSS.n2570 VSS.n2569 2.6005
R3785 VSS.n2857 VSS.n2856 2.6005
R3786 VSS.n2859 VSS.n2858 2.6005
R3787 VSS.n2861 VSS.n2860 2.6005
R3788 VSS.n3970 VSS.n3969 2.6005
R3789 VSS.n4044 VSS.n4043 2.6005
R3790 VSS.n4042 VSS.n4041 2.6005
R3791 VSS.n4039 VSS.n4038 2.6005
R3792 VSS.n4037 VSS.n4036 2.6005
R3793 VSS.n4034 VSS.n4033 2.6005
R3794 VSS.n4032 VSS.n4031 2.6005
R3795 VSS.n4029 VSS.n4028 2.6005
R3796 VSS.n4027 VSS.n4026 2.6005
R3797 VSS.n4024 VSS.n4023 2.6005
R3798 VSS.n4022 VSS.n4021 2.6005
R3799 VSS.n4019 VSS.n4018 2.6005
R3800 VSS.n4017 VSS.n4016 2.6005
R3801 VSS.n4014 VSS.n4013 2.6005
R3802 VSS.n4012 VSS.n4011 2.6005
R3803 VSS.n4009 VSS.n4008 2.6005
R3804 VSS.n4007 VSS.n4006 2.6005
R3805 VSS.n4004 VSS.n4003 2.6005
R3806 VSS.n4002 VSS.n4001 2.6005
R3807 VSS.n4000 VSS.n3999 2.6005
R3808 VSS.n3998 VSS.n3997 2.6005
R3809 VSS.n3996 VSS.n3995 2.6005
R3810 VSS.n3994 VSS.n3993 2.6005
R3811 VSS.n3992 VSS.n3991 2.6005
R3812 VSS.n3990 VSS.n3989 2.6005
R3813 VSS.n3988 VSS.n3987 2.6005
R3814 VSS.n3986 VSS.n3985 2.6005
R3815 VSS.n3984 VSS.n3983 2.6005
R3816 VSS.n3982 VSS.n3981 2.6005
R3817 VSS.n3980 VSS.n3979 2.6005
R3818 VSS.n3978 VSS.n3977 2.6005
R3819 VSS.n3976 VSS.n3975 2.6005
R3820 VSS.n3974 VSS.n3973 2.6005
R3821 VSS.n3972 VSS.n3971 2.6005
R3822 VSS.n3968 VSS.n3837 2.6005
R3823 VSS.n3931 VSS.n3930 2.6005
R3824 VSS.n3934 VSS.n3933 2.6005
R3825 VSS.n3933 VSS.n3932 2.6005
R3826 VSS.n3937 VSS.n3936 2.6005
R3827 VSS.n3936 VSS.n3935 2.6005
R3828 VSS.n3941 VSS.n3940 2.6005
R3829 VSS.n3940 VSS.n3939 2.6005
R3830 VSS.n3944 VSS.n3943 2.6005
R3831 VSS.n3943 VSS.n3942 2.6005
R3832 VSS.n3952 VSS.n3951 2.6005
R3833 VSS.n3951 VSS.n3950 2.6005
R3834 VSS.n3955 VSS.n3954 2.6005
R3835 VSS.n3954 VSS.n3953 2.6005
R3836 VSS.n3958 VSS.n3957 2.6005
R3837 VSS.n3957 VSS.n3956 2.6005
R3838 VSS.n3961 VSS.n3960 2.6005
R3839 VSS.n3960 VSS.n3959 2.6005
R3840 VSS.n3964 VSS.n3963 2.6005
R3841 VSS.n3963 VSS.n3962 2.6005
R3842 VSS.n3967 VSS.n3966 2.6005
R3843 VSS.n3966 VSS.n3965 2.6005
R3844 VSS.n2957 VSS.n2956 2.6005
R3845 VSS.n2955 VSS.n2954 2.6005
R3846 VSS.n2952 VSS.n2951 2.6005
R3847 VSS.n2950 VSS.n2949 2.6005
R3848 VSS.n2945 VSS.n2944 2.6005
R3849 VSS.n2943 VSS.n2942 2.6005
R3850 VSS.n2940 VSS.n2939 2.6005
R3851 VSS.n2937 VSS.n2936 2.6005
R3852 VSS.n2935 VSS.n2934 2.6005
R3853 VSS.n2932 VSS.n2931 2.6005
R3854 VSS.n2930 VSS.n2929 2.6005
R3855 VSS.n2927 VSS.n2926 2.6005
R3856 VSS.n2924 VSS.n2923 2.6005
R3857 VSS.n2922 VSS.n2921 2.6005
R3858 VSS.n2920 VSS.n2919 2.6005
R3859 VSS.n2918 VSS.n2917 2.6005
R3860 VSS.n2916 VSS.n2915 2.6005
R3861 VSS.n2914 VSS.n2913 2.6005
R3862 VSS.n2912 VSS.n2911 2.6005
R3863 VSS.n2910 VSS.n2909 2.6005
R3864 VSS.n2908 VSS.n2907 2.6005
R3865 VSS.n2906 VSS.n2905 2.6005
R3866 VSS.n2904 VSS.n2903 2.6005
R3867 VSS.n2902 VSS.n2901 2.6005
R3868 VSS.n2900 VSS.n2899 2.6005
R3869 VSS.n2898 VSS.n2897 2.6005
R3870 VSS.n2896 VSS.n2895 2.6005
R3871 VSS.n2894 VSS.n2893 2.6005
R3872 VSS.n2891 VSS.n2890 2.6005
R3873 VSS.n2889 VSS.n2888 2.6005
R3874 VSS.n2887 VSS.n2886 2.6005
R3875 VSS.n2885 VSS.n2884 2.6005
R3876 VSS.n2883 VSS.n2882 2.6005
R3877 VSS.n2880 VSS.n2879 2.6005
R3878 VSS.n2878 VSS.n2877 2.6005
R3879 VSS.n2876 VSS.n2875 2.6005
R3880 VSS.n3849 VSS.n3848 2.6005
R3881 VSS.n3852 VSS.n3851 2.6005
R3882 VSS.n3854 VSS.n3853 2.6005
R3883 VSS.n3856 VSS.n3855 2.6005
R3884 VSS.n3858 VSS.n3857 2.6005
R3885 VSS.n3860 VSS.n3859 2.6005
R3886 VSS.n3863 VSS.n3862 2.6005
R3887 VSS.n3865 VSS.n3864 2.6005
R3888 VSS.n3867 VSS.n3866 2.6005
R3889 VSS.n3869 VSS.n3868 2.6005
R3890 VSS.n3872 VSS.n3871 2.6005
R3891 VSS.n3874 VSS.n3873 2.6005
R3892 VSS.n3876 VSS.n3875 2.6005
R3893 VSS.n3878 VSS.n3877 2.6005
R3894 VSS.n3881 VSS.n3880 2.6005
R3895 VSS.n3883 VSS.n3882 2.6005
R3896 VSS.n3886 VSS.n3885 2.6005
R3897 VSS.n3888 VSS.n3887 2.6005
R3898 VSS.n3890 VSS.n3889 2.6005
R3899 VSS.n2629 VSS.n2628 2.6005
R3900 VSS.n2594 VSS.n2593 2.6005
R3901 VSS.n2597 VSS.n2596 2.6005
R3902 VSS.n2596 VSS.n2595 2.6005
R3903 VSS.n2600 VSS.n2599 2.6005
R3904 VSS.n2599 VSS.n2598 2.6005
R3905 VSS.n2604 VSS.n2603 2.6005
R3906 VSS.n2603 VSS.n2602 2.6005
R3907 VSS.n2607 VSS.n2606 2.6005
R3908 VSS.n2606 VSS.n2605 2.6005
R3909 VSS.n2611 VSS.n2610 2.6005
R3910 VSS.n2610 VSS.n2609 2.6005
R3911 VSS.n2614 VSS.n2613 2.6005
R3912 VSS.n2613 VSS.n2612 2.6005
R3913 VSS.n2617 VSS.n2616 2.6005
R3914 VSS.n2616 VSS.n2615 2.6005
R3915 VSS.n2620 VSS.n2619 2.6005
R3916 VSS.n2619 VSS.n2618 2.6005
R3917 VSS.n2623 VSS.n2622 2.6005
R3918 VSS.n2622 VSS.n2621 2.6005
R3919 VSS.n2626 VSS.n2625 2.6005
R3920 VSS.n2625 VSS.n2624 2.6005
R3921 VSS.n3370 VSS.n3369 2.6005
R3922 VSS.n3368 VSS.n3367 2.6005
R3923 VSS.n3365 VSS.n3364 2.6005
R3924 VSS.n3363 VSS.n3362 2.6005
R3925 VSS.n3360 VSS.n3359 2.6005
R3926 VSS.n3358 VSS.n3357 2.6005
R3927 VSS.n3355 VSS.n3354 2.6005
R3928 VSS.n3353 VSS.n3352 2.6005
R3929 VSS.n3350 VSS.n3349 2.6005
R3930 VSS.n3348 VSS.n3347 2.6005
R3931 VSS.n3345 VSS.n3344 2.6005
R3932 VSS.n3343 VSS.n3342 2.6005
R3933 VSS.n3340 VSS.n3339 2.6005
R3934 VSS.n3338 VSS.n3337 2.6005
R3935 VSS.n3335 VSS.n3334 2.6005
R3936 VSS.n3333 VSS.n3332 2.6005
R3937 VSS.n3331 VSS.n3330 2.6005
R3938 VSS.n2631 VSS.n2630 2.6005
R3939 VSS.n2633 VSS.n2632 2.6005
R3940 VSS.n2635 VSS.n2634 2.6005
R3941 VSS.n2637 VSS.n2636 2.6005
R3942 VSS.n2642 VSS.n2641 2.6005
R3943 VSS.n2645 VSS.n2644 2.6005
R3944 VSS.n2647 VSS.n2646 2.6005
R3945 VSS.n2649 VSS.n2648 2.6005
R3946 VSS.n2651 VSS.n2650 2.6005
R3947 VSS.n2653 VSS.n2652 2.6005
R3948 VSS.n2656 VSS.n2655 2.6005
R3949 VSS.n2659 VSS.n2658 2.6005
R3950 VSS.n2662 VSS.n2661 2.6005
R3951 VSS.n3380 VSS.n3379 2.6005
R3952 VSS.n2530 VSS.n2529 2.6005
R3953 VSS.n2529 VSS.n2528 2.6005
R3954 VSS.n2527 VSS.n2526 2.6005
R3955 VSS.n2526 VSS.n2525 2.6005
R3956 VSS.n2524 VSS.n2523 2.6005
R3957 VSS.n2523 VSS.n2522 2.6005
R3958 VSS.n2521 VSS.n2520 2.6005
R3959 VSS.n2520 VSS.n2519 2.6005
R3960 VSS.n2517 VSS.n2516 2.6005
R3961 VSS.n2516 VSS.n2515 2.6005
R3962 VSS.n2514 VSS.n2513 2.6005
R3963 VSS.n2513 VSS.n2512 2.6005
R3964 VSS.n2510 VSS.n2509 2.6005
R3965 VSS.n2509 VSS.n2508 2.6005
R3966 VSS.n2507 VSS.n2506 2.6005
R3967 VSS.n2506 VSS.n2505 2.6005
R3968 VSS.n2504 VSS.n2503 2.6005
R3969 VSS.n2503 VSS.n2502 2.6005
R3970 VSS.n2501 VSS.n2500 2.6005
R3971 VSS.n2500 VSS.n2499 2.6005
R3972 VSS.n2498 VSS.n2497 2.6005
R3973 VSS.n2497 VSS.n2496 2.6005
R3974 VSS.n2495 VSS.n2494 2.6005
R3975 VSS.n2494 VSS.n2493 2.6005
R3976 VSS.n2492 VSS.n2491 2.6005
R3977 VSS.n2491 VSS.n2490 2.6005
R3978 VSS.n2489 VSS.n2488 2.6005
R3979 VSS.n2488 VSS.n2487 2.6005
R3980 VSS.n2485 VSS.n2484 2.6005
R3981 VSS.n2484 VSS.n2483 2.6005
R3982 VSS.n2482 VSS.n2481 2.6005
R3983 VSS.n2481 VSS.n2480 2.6005
R3984 VSS.n3789 VSS.n3788 2.6005
R3985 VSS.n3788 VSS.n3787 2.6005
R3986 VSS.n3792 VSS.n3791 2.6005
R3987 VSS.n3791 VSS.n3790 2.6005
R3988 VSS.n3795 VSS.n3794 2.6005
R3989 VSS.n3794 VSS.n3793 2.6005
R3990 VSS.n3798 VSS.n3797 2.6005
R3991 VSS.n3797 VSS.n3796 2.6005
R3992 VSS.n3801 VSS.n3800 2.6005
R3993 VSS.n3800 VSS.n3799 2.6005
R3994 VSS.n3804 VSS.n3803 2.6005
R3995 VSS.n3803 VSS.n3802 2.6005
R3996 VSS.n3807 VSS.n3806 2.6005
R3997 VSS.n3806 VSS.n3805 2.6005
R3998 VSS.n3810 VSS.n3809 2.6005
R3999 VSS.n3809 VSS.n3808 2.6005
R4000 VSS.n3813 VSS.n3812 2.6005
R4001 VSS.n3812 VSS.n3811 2.6005
R4002 VSS.n3816 VSS.n3815 2.6005
R4003 VSS.n3815 VSS.n3814 2.6005
R4004 VSS.n3820 VSS.n3819 2.6005
R4005 VSS.n3819 VSS.n3818 2.6005
R4006 VSS.n3823 VSS.n3822 2.6005
R4007 VSS.n3822 VSS.n3821 2.6005
R4008 VSS.n3827 VSS.n3826 2.6005
R4009 VSS.n3826 VSS.n3825 2.6005
R4010 VSS.n3830 VSS.n3829 2.6005
R4011 VSS.n3829 VSS.n3828 2.6005
R4012 VSS.n3833 VSS.n3832 2.6005
R4013 VSS.n3832 VSS.n3831 2.6005
R4014 VSS.n3836 VSS.n3835 2.6005
R4015 VSS.n3835 VSS.n3834 2.6005
R4016 VSS.n4057 VSS.n4056 2.6005
R4017 VSS.n357 VSS.n356 2.6005
R4018 VSS.n355 VSS.n354 2.6005
R4019 VSS.n352 VSS.n351 2.6005
R4020 VSS.n349 VSS.n348 2.6005
R4021 VSS.n347 VSS.n346 2.6005
R4022 VSS.n345 VSS.n344 2.6005
R4023 VSS.n342 VSS.n341 2.6005
R4024 VSS.n340 VSS.n339 2.6005
R4025 VSS.n338 VSS.n337 2.6005
R4026 VSS.n336 VSS.n335 2.6005
R4027 VSS.n333 VSS.n332 2.6005
R4028 VSS.n331 VSS.n330 2.6005
R4029 VSS.n329 VSS.n328 2.6005
R4030 VSS.n326 VSS.n325 2.6005
R4031 VSS.n324 VSS.n323 2.6005
R4032 VSS.n322 VSS.n321 2.6005
R4033 VSS.n320 VSS.n319 2.6005
R4034 VSS.n317 VSS.n316 2.6005
R4035 VSS.n315 VSS.n314 2.6005
R4036 VSS.n313 VSS.n312 2.6005
R4037 VSS.n307 VSS.n306 2.6005
R4038 VSS.n304 VSS.n303 2.6005
R4039 VSS.n302 VSS.n301 2.6005
R4040 VSS.n3732 VSS.n3731 2.6005
R4041 VSS.n4063 VSS.n4062 2.6005
R4042 VSS.n4062 VSS.n4061 2.6005
R4043 VSS.n3772 VSS.n3771 2.6005
R4044 VSS.n3771 VSS.n3770 2.6005
R4045 VSS.n3752 VSS.n3751 2.6005
R4046 VSS.n3751 VSS.n3750 2.6005
R4047 VSS.n3749 VSS.n3748 2.6005
R4048 VSS.n3748 VSS.n3747 2.6005
R4049 VSS.n3746 VSS.n3745 2.6005
R4050 VSS.n3745 VSS.n3744 2.6005
R4051 VSS.n3742 VSS.n3741 2.6005
R4052 VSS.n3741 VSS.n3740 2.6005
R4053 VSS.n3738 VSS.n3737 2.6005
R4054 VSS.n3737 VSS.n3736 2.6005
R4055 VSS.n3735 VSS.n3734 2.6005
R4056 VSS.n3734 VSS.n3733 2.6005
R4057 VSS.n2214 VSS.n2213 2.6005
R4058 VSS.n2218 VSS.n2217 2.6005
R4059 VSS.n2220 VSS.n2219 2.6005
R4060 VSS.n2222 VSS.n2221 2.6005
R4061 VSS.n2224 VSS.n2223 2.6005
R4062 VSS.n2226 VSS.n2225 2.6005
R4063 VSS.n2228 VSS.n2227 2.6005
R4064 VSS.n2230 VSS.n2229 2.6005
R4065 VSS.n2232 VSS.n2231 2.6005
R4066 VSS.n2234 VSS.n2233 2.6005
R4067 VSS.n2236 VSS.n2235 2.6005
R4068 VSS.n2238 VSS.n2237 2.6005
R4069 VSS.n2240 VSS.n2239 2.6005
R4070 VSS.n2242 VSS.n2241 2.6005
R4071 VSS.n2244 VSS.n2243 2.6005
R4072 VSS.n2246 VSS.n2245 2.6005
R4073 VSS.n2248 VSS.n2247 2.6005
R4074 VSS.n2250 VSS.n2249 2.6005
R4075 VSS.n2252 VSS.n2251 2.6005
R4076 VSS.n2254 VSS.n2253 2.6005
R4077 VSS.n2256 VSS.n2255 2.6005
R4078 VSS.n2258 VSS.n2257 2.6005
R4079 VSS.n2260 VSS.n2259 2.6005
R4080 VSS.n2262 VSS.n2261 2.6005
R4081 VSS.n2264 VSS.n2263 2.6005
R4082 VSS.n2266 VSS.n2265 2.6005
R4083 VSS.n2268 VSS.n2267 2.6005
R4084 VSS.n2270 VSS.n2269 2.6005
R4085 VSS.n2272 VSS.n2271 2.6005
R4086 VSS.n2275 VSS.n2274 2.6005
R4087 VSS.n2277 VSS.n2276 2.6005
R4088 VSS.n2280 VSS.n2279 2.6005
R4089 VSS.n2282 VSS.n2281 2.6005
R4090 VSS.n2285 VSS.n2284 2.6005
R4091 VSS.n2287 VSS.n2286 2.6005
R4092 VSS.n2290 VSS.n2289 2.6005
R4093 VSS.n2292 VSS.n2291 2.6005
R4094 VSS.n2295 VSS.n2294 2.6005
R4095 VSS.n2216 VSS.n2215 2.6005
R4096 VSS.n2297 VSS.n2296 2.6005
R4097 VSS VSS.n3472 2.6005
R4098 VSS.n3386 VSS.n3385 2.6005
R4099 VSS.n3385 VSS.n3384 2.6005
R4100 VSS.n3389 VSS.n3388 2.6005
R4101 VSS.n3388 VSS.n3387 2.6005
R4102 VSS.n3392 VSS.n3391 2.6005
R4103 VSS.n3391 VSS.n3390 2.6005
R4104 VSS.n3395 VSS.n3394 2.6005
R4105 VSS.n3394 VSS.n3393 2.6005
R4106 VSS.n3398 VSS.n3397 2.6005
R4107 VSS.n3397 VSS.n3396 2.6005
R4108 VSS.n3401 VSS.n3400 2.6005
R4109 VSS.n3400 VSS.n3399 2.6005
R4110 VSS.n3404 VSS.n3403 2.6005
R4111 VSS.n3403 VSS.n3402 2.6005
R4112 VSS.n3407 VSS.n3406 2.6005
R4113 VSS.n3406 VSS.n3405 2.6005
R4114 VSS.n3410 VSS.n3409 2.6005
R4115 VSS.n3409 VSS.n3408 2.6005
R4116 VSS.n3413 VSS.n3412 2.6005
R4117 VSS.n3412 VSS.n3411 2.6005
R4118 VSS.n3416 VSS.n3415 2.6005
R4119 VSS.n3415 VSS.n3414 2.6005
R4120 VSS.n3419 VSS.n3418 2.6005
R4121 VSS.n3418 VSS.n3417 2.6005
R4122 VSS.n3423 VSS.n3422 2.6005
R4123 VSS.n3422 VSS.n3421 2.6005
R4124 VSS.n3426 VSS.n3425 2.6005
R4125 VSS.n3425 VSS.n3424 2.6005
R4126 VSS.n3430 VSS.n3429 2.6005
R4127 VSS.n3429 VSS.n3428 2.6005
R4128 VSS.n4113 VSS.n4112 2.6005
R4129 VSS.n4112 VSS.n4111 2.6005
R4130 VSS.n4110 VSS.n4109 2.6005
R4131 VSS.n4109 VSS.n4108 2.6005
R4132 VSS.n4106 VSS.n4105 2.6005
R4133 VSS.n4105 VSS.n4104 2.6005
R4134 VSS.n4102 VSS.n4101 2.6005
R4135 VSS.n4101 VSS.n4100 2.6005
R4136 VSS.n4099 VSS.n4098 2.6005
R4137 VSS.n4098 VSS.n4097 2.6005
R4138 VSS.n4096 VSS.n4095 2.6005
R4139 VSS.n4095 VSS.n4094 2.6005
R4140 VSS.n4092 VSS.n4091 2.6005
R4141 VSS.n4091 VSS.n4090 2.6005
R4142 VSS.n4089 VSS.n4088 2.6005
R4143 VSS.n4088 VSS.n4087 2.6005
R4144 VSS.n4086 VSS.n4085 2.6005
R4145 VSS.n4085 VSS.n4084 2.6005
R4146 VSS.n4083 VSS.n4082 2.6005
R4147 VSS.n4082 VSS.n4081 2.6005
R4148 VSS.n4079 VSS.n4078 2.6005
R4149 VSS.n4078 VSS.n4077 2.6005
R4150 VSS.n4076 VSS.n4075 2.6005
R4151 VSS.n4075 VSS.n4074 2.6005
R4152 VSS.n4073 VSS.n4072 2.6005
R4153 VSS.n4072 VSS.n4071 2.6005
R4154 VSS.n4069 VSS.n4068 2.6005
R4155 VSS.n4068 VSS.n4067 2.6005
R4156 VSS.n4066 VSS.n4065 2.6005
R4157 VSS.n4065 VSS.n4064 2.6005
R4158 VSS.n2461 VSS.n2460 2.6005
R4159 VSS.n2460 VSS.n2459 2.6005
R4160 VSS.n2465 VSS.n2464 2.6005
R4161 VSS.n2464 VSS.n2463 2.6005
R4162 VSS.n2420 VSS.n2419 2.6005
R4163 VSS.n2419 VSS.n2418 2.6005
R4164 VSS.n2424 VSS.n2423 2.6005
R4165 VSS.n2423 VSS.n2422 2.6005
R4166 VSS.n2427 VSS.n2426 2.6005
R4167 VSS.n2426 VSS.n2425 2.6005
R4168 VSS.n2437 VSS.n2436 2.6005
R4169 VSS.n2436 VSS.n2435 2.6005
R4170 VSS.n2440 VSS.n2439 2.6005
R4171 VSS.n2439 VSS.n2438 2.6005
R4172 VSS.n2443 VSS.n2442 2.6005
R4173 VSS.n2442 VSS.n2441 2.6005
R4174 VSS.n2446 VSS.n2445 2.6005
R4175 VSS.n2445 VSS.n2444 2.6005
R4176 VSS.n2449 VSS.n2448 2.6005
R4177 VSS.n2448 VSS.n2447 2.6005
R4178 VSS.n2452 VSS.n2451 2.6005
R4179 VSS.n2451 VSS.n2450 2.6005
R4180 VSS.n2455 VSS.n2454 2.6005
R4181 VSS.n2454 VSS.n2453 2.6005
R4182 VSS.n2458 VSS.n2457 2.6005
R4183 VSS.n2457 VSS.n2456 2.6005
R4184 VSS.n2417 VSS.n2416 2.6005
R4185 VSS.n2212 VSS.n2211 2.6005
R4186 VSS.n2313 VSS.n2312 2.6005
R4187 VSS.n5 VSS.n4 2.6005
R4188 VSS.n8 VSS.n7 2.6005
R4189 VSS.n10 VSS.n9 2.6005
R4190 VSS.n13 VSS.n12 2.6005
R4191 VSS.n15 VSS.n14 2.6005
R4192 VSS.n18 VSS.n17 2.6005
R4193 VSS.n20 VSS.n19 2.6005
R4194 VSS.n22 VSS.n21 2.6005
R4195 VSS.n24 VSS.n23 2.6005
R4196 VSS.n26 VSS.n25 2.6005
R4197 VSS.n28 VSS.n27 2.6005
R4198 VSS.n30 VSS.n29 2.6005
R4199 VSS.n32 VSS.n31 2.6005
R4200 VSS.n34 VSS.n33 2.6005
R4201 VSS.n37 VSS.n36 2.6005
R4202 VSS.n39 VSS.n38 2.6005
R4203 VSS.n41 VSS.n40 2.6005
R4204 VSS.n43 VSS.n42 2.6005
R4205 VSS.n45 VSS.n44 2.6005
R4206 VSS.n47 VSS.n46 2.6005
R4207 VSS.n49 VSS.n48 2.6005
R4208 VSS.n52 VSS.n51 2.6005
R4209 VSS.n54 VSS.n53 2.6005
R4210 VSS.n56 VSS.n55 2.6005
R4211 VSS.n58 VSS.n57 2.6005
R4212 VSS.n61 VSS.n60 2.6005
R4213 VSS.n63 VSS.n62 2.6005
R4214 VSS.n66 VSS.n65 2.6005
R4215 VSS.n237 VSS.n236 2.6005
R4216 VSS.n68 VSS.n67 2.6005
R4217 VSS.n226 VSS.n225 2.6005
R4218 VSS.n224 VSS.n223 2.6005
R4219 VSS.n222 VSS.n221 2.6005
R4220 VSS.n228 VSS.n227 2.6005
R4221 VSS.n2209 VSS.n2208 2.6005
R4222 VSS.n2181 VSS.n2180 2.6005
R4223 VSS.n2183 VSS.n2182 2.6005
R4224 VSS.n2185 VSS.n2184 2.6005
R4225 VSS.n2187 VSS.n2186 2.6005
R4226 VSS.n2189 VSS.n2188 2.6005
R4227 VSS.n2191 VSS.n2190 2.6005
R4228 VSS.n2193 VSS.n2192 2.6005
R4229 VSS.n2195 VSS.n2194 2.6005
R4230 VSS.n2197 VSS.n2196 2.6005
R4231 VSS.n2199 VSS.n2198 2.6005
R4232 VSS.n2201 VSS.n2200 2.6005
R4233 VSS.n2203 VSS.n2202 2.6005
R4234 VSS.n2205 VSS.n2204 2.6005
R4235 VSS.n2207 VSS.n2206 2.6005
R4236 VSS.n2179 VSS.n2178 2.6005
R4237 VSS.n2169 VSS.n2168 2.6005
R4238 VSS.n2176 VSS.n2173 2.6005
R4239 VSS.n2176 VSS.n2175 2.6005
R4240 VSS.n2023 VSS.n1412 2.6005
R4241 VSS.n2142 VSS.n2141 2.6005
R4242 VSS.n2139 VSS.n2138 2.6005
R4243 VSS.n2137 VSS.n2136 2.6005
R4244 VSS.n2134 VSS.n2133 2.6005
R4245 VSS.n2132 VSS.n2131 2.6005
R4246 VSS.n2129 VSS.n2128 2.6005
R4247 VSS.n2127 VSS.n2126 2.6005
R4248 VSS.n2124 VSS.n2123 2.6005
R4249 VSS.n2122 VSS.n2121 2.6005
R4250 VSS.n2119 VSS.n2118 2.6005
R4251 VSS.n2117 VSS.n2116 2.6005
R4252 VSS.n2114 VSS.n2113 2.6005
R4253 VSS.n2112 VSS.n2111 2.6005
R4254 VSS.n2109 VSS.n2108 2.6005
R4255 VSS.n2107 VSS.n2106 2.6005
R4256 VSS.n2104 VSS.n2103 2.6005
R4257 VSS.n2102 VSS.n2101 2.6005
R4258 VSS.n2099 VSS.n2098 2.6005
R4259 VSS.n2097 VSS.n2096 2.6005
R4260 VSS.n2095 VSS.n2094 2.6005
R4261 VSS.n2093 VSS.n2092 2.6005
R4262 VSS.n2091 VSS.n2090 2.6005
R4263 VSS.n2089 VSS.n2088 2.6005
R4264 VSS.n2087 VSS.n2086 2.6005
R4265 VSS.n2085 VSS.n2084 2.6005
R4266 VSS.n2083 VSS.n2082 2.6005
R4267 VSS.n2081 VSS.n2080 2.6005
R4268 VSS.n2079 VSS.n2078 2.6005
R4269 VSS.n2077 VSS.n2076 2.6005
R4270 VSS.n2075 VSS.n2074 2.6005
R4271 VSS.n2073 VSS.n2072 2.6005
R4272 VSS.n2071 VSS.n2070 2.6005
R4273 VSS.n2069 VSS.n2068 2.6005
R4274 VSS.n2067 VSS.n2066 2.6005
R4275 VSS.n2065 VSS.n2064 2.6005
R4276 VSS.n2063 VSS.n2062 2.6005
R4277 VSS.n2061 VSS.n2060 2.6005
R4278 VSS.n2059 VSS.n2058 2.6005
R4279 VSS.n2057 VSS.n2056 2.6005
R4280 VSS.n2055 VSS.n2054 2.6005
R4281 VSS.n2053 VSS.n2052 2.6005
R4282 VSS.n2051 VSS.n2050 2.6005
R4283 VSS.n2049 VSS.n2048 2.6005
R4284 VSS.n2047 VSS.n2046 2.6005
R4285 VSS.n2045 VSS.n2044 2.6005
R4286 VSS.n2043 VSS.n2042 2.6005
R4287 VSS.n2041 VSS.n2040 2.6005
R4288 VSS.n2039 VSS.n2038 2.6005
R4289 VSS.n2037 VSS.n2036 2.6005
R4290 VSS.n2035 VSS.n2034 2.6005
R4291 VSS.n2033 VSS.n2032 2.6005
R4292 VSS.n2031 VSS.n2030 2.6005
R4293 VSS.n2029 VSS.n2028 2.6005
R4294 VSS.n2027 VSS.n2026 2.6005
R4295 VSS.n2025 VSS.n2024 2.6005
R4296 VSS.n1950 VSS.n1949 2.6005
R4297 VSS.n1954 VSS.n1953 2.6005
R4298 VSS.n1956 VSS.n1955 2.6005
R4299 VSS.n1958 VSS.n1957 2.6005
R4300 VSS.n1960 VSS.n1959 2.6005
R4301 VSS.n1962 VSS.n1961 2.6005
R4302 VSS.n1964 VSS.n1963 2.6005
R4303 VSS.n1967 VSS.n1966 2.6005
R4304 VSS.n1970 VSS.n1969 2.6005
R4305 VSS.n1972 VSS.n1971 2.6005
R4306 VSS.n1974 VSS.n1973 2.6005
R4307 VSS.n1977 VSS.n1976 2.6005
R4308 VSS.n1979 VSS.n1978 2.6005
R4309 VSS.n1981 VSS.n1980 2.6005
R4310 VSS.n1983 VSS.n1982 2.6005
R4311 VSS.n1985 VSS.n1984 2.6005
R4312 VSS.n1987 VSS.n1986 2.6005
R4313 VSS.n1989 VSS.n1988 2.6005
R4314 VSS.n1991 VSS.n1990 2.6005
R4315 VSS.n1993 VSS.n1992 2.6005
R4316 VSS.n1995 VSS.n1994 2.6005
R4317 VSS.n1997 VSS.n1996 2.6005
R4318 VSS.n1999 VSS.n1998 2.6005
R4319 VSS.n2001 VSS.n2000 2.6005
R4320 VSS.n2003 VSS.n2002 2.6005
R4321 VSS.n2006 VSS.n2005 2.6005
R4322 VSS.n2009 VSS.n2008 2.6005
R4323 VSS.n2011 VSS.n2010 2.6005
R4324 VSS.n2013 VSS.n2012 2.6005
R4325 VSS.n2015 VSS.n2014 2.6005
R4326 VSS.n2017 VSS.n2016 2.6005
R4327 VSS.n2019 VSS.n2018 2.6005
R4328 VSS.n1950 VSS.n1948 2.6005
R4329 VSS.n1872 VSS.n1871 2.6005
R4330 VSS.n1876 VSS.n1875 2.6005
R4331 VSS.n1878 VSS.n1877 2.6005
R4332 VSS.n1880 VSS.n1879 2.6005
R4333 VSS.n1882 VSS.n1881 2.6005
R4334 VSS.n1884 VSS.n1883 2.6005
R4335 VSS.n1886 VSS.n1885 2.6005
R4336 VSS.n1889 VSS.n1888 2.6005
R4337 VSS.n1892 VSS.n1891 2.6005
R4338 VSS.n1894 VSS.n1893 2.6005
R4339 VSS.n1896 VSS.n1895 2.6005
R4340 VSS.n1898 VSS.n1897 2.6005
R4341 VSS.n1900 VSS.n1899 2.6005
R4342 VSS.n1902 VSS.n1901 2.6005
R4343 VSS.n1904 VSS.n1903 2.6005
R4344 VSS.n1906 VSS.n1905 2.6005
R4345 VSS.n1908 VSS.n1907 2.6005
R4346 VSS.n1910 VSS.n1909 2.6005
R4347 VSS.n1912 VSS.n1911 2.6005
R4348 VSS.n1914 VSS.n1913 2.6005
R4349 VSS.n1916 VSS.n1915 2.6005
R4350 VSS.n1918 VSS.n1917 2.6005
R4351 VSS.n1921 VSS.n1920 2.6005
R4352 VSS.n1923 VSS.n1922 2.6005
R4353 VSS.n1925 VSS.n1924 2.6005
R4354 VSS.n1928 VSS.n1927 2.6005
R4355 VSS.n1931 VSS.n1930 2.6005
R4356 VSS.n1933 VSS.n1932 2.6005
R4357 VSS.n1935 VSS.n1934 2.6005
R4358 VSS.n1937 VSS.n1936 2.6005
R4359 VSS.n1939 VSS.n1938 2.6005
R4360 VSS.n1941 VSS.n1940 2.6005
R4361 VSS.n1872 VSS.n1870 2.6005
R4362 VSS.n1791 VSS.n1790 2.6005
R4363 VSS.n1794 VSS.n1793 2.6005
R4364 VSS.n1796 VSS.n1795 2.6005
R4365 VSS.n1798 VSS.n1797 2.6005
R4366 VSS.n1800 VSS.n1799 2.6005
R4367 VSS.n1802 VSS.n1801 2.6005
R4368 VSS.n1804 VSS.n1803 2.6005
R4369 VSS.n1811 VSS.n1810 2.6005
R4370 VSS.n1814 VSS.n1813 2.6005
R4371 VSS.n1816 VSS.n1815 2.6005
R4372 VSS.n1818 VSS.n1817 2.6005
R4373 VSS.n1821 VSS.n1820 2.6005
R4374 VSS.n1823 VSS.n1822 2.6005
R4375 VSS.n1825 VSS.n1824 2.6005
R4376 VSS.n1827 VSS.n1826 2.6005
R4377 VSS.n1829 VSS.n1828 2.6005
R4378 VSS.n1831 VSS.n1830 2.6005
R4379 VSS.n1833 VSS.n1832 2.6005
R4380 VSS.n1835 VSS.n1834 2.6005
R4381 VSS.n1837 VSS.n1836 2.6005
R4382 VSS.n1839 VSS.n1838 2.6005
R4383 VSS.n1841 VSS.n1840 2.6005
R4384 VSS.n1843 VSS.n1842 2.6005
R4385 VSS.n1845 VSS.n1844 2.6005
R4386 VSS.n1847 VSS.n1846 2.6005
R4387 VSS.n1850 VSS.n1849 2.6005
R4388 VSS.n1853 VSS.n1852 2.6005
R4389 VSS.n1855 VSS.n1854 2.6005
R4390 VSS.n1857 VSS.n1856 2.6005
R4391 VSS.n1859 VSS.n1858 2.6005
R4392 VSS.n1861 VSS.n1860 2.6005
R4393 VSS.n1863 VSS.n1862 2.6005
R4394 VSS.n1791 VSS.n1789 2.6005
R4395 VSS.n1294 VSS.n1293 2.6005
R4396 VSS.n1111 VSS.n1110 2.6005
R4397 VSS.n928 VSS.n927 2.6005
R4398 VSS.n234 VSS.n233 2.6005
R4399 VSS.n1298 VSS.n1297 2.6005
R4400 VSS.n1297 VSS.n1296 2.6005
R4401 VSS.n1301 VSS.n1300 2.6005
R4402 VSS.n1300 VSS.n1299 2.6005
R4403 VSS.n1304 VSS.n1303 2.6005
R4404 VSS.n1303 VSS.n1302 2.6005
R4405 VSS.n1307 VSS.n1306 2.6005
R4406 VSS.n1306 VSS.n1305 2.6005
R4407 VSS.n1310 VSS.n1309 2.6005
R4408 VSS.n1309 VSS.n1308 2.6005
R4409 VSS.n1313 VSS.n1312 2.6005
R4410 VSS.n1312 VSS.n1311 2.6005
R4411 VSS.n1317 VSS.n1316 2.6005
R4412 VSS.n1316 VSS.n1315 2.6005
R4413 VSS.n1321 VSS.n1320 2.6005
R4414 VSS.n1320 VSS.n1319 2.6005
R4415 VSS.n1324 VSS.n1323 2.6005
R4416 VSS.n1323 VSS.n1322 2.6005
R4417 VSS.n1327 VSS.n1326 2.6005
R4418 VSS.n1326 VSS.n1325 2.6005
R4419 VSS.n1330 VSS.n1329 2.6005
R4420 VSS.n1329 VSS.n1328 2.6005
R4421 VSS.n1333 VSS.n1332 2.6005
R4422 VSS.n1332 VSS.n1331 2.6005
R4423 VSS.n1336 VSS.n1335 2.6005
R4424 VSS.n1335 VSS.n1334 2.6005
R4425 VSS.n1339 VSS.n1338 2.6005
R4426 VSS.n1338 VSS.n1337 2.6005
R4427 VSS.n1342 VSS.n1341 2.6005
R4428 VSS.n1341 VSS.n1340 2.6005
R4429 VSS.n1345 VSS.n1344 2.6005
R4430 VSS.n1344 VSS.n1343 2.6005
R4431 VSS.n1348 VSS.n1347 2.6005
R4432 VSS.n1347 VSS.n1346 2.6005
R4433 VSS.n1351 VSS.n1350 2.6005
R4434 VSS.n1350 VSS.n1349 2.6005
R4435 VSS.n1354 VSS.n1353 2.6005
R4436 VSS.n1353 VSS.n1352 2.6005
R4437 VSS.n1357 VSS.n1356 2.6005
R4438 VSS.n1356 VSS.n1355 2.6005
R4439 VSS.n1360 VSS.n1359 2.6005
R4440 VSS.n1359 VSS.n1358 2.6005
R4441 VSS.n1363 VSS.n1362 2.6005
R4442 VSS.n1362 VSS.n1361 2.6005
R4443 VSS.n1366 VSS.n1365 2.6005
R4444 VSS.n1365 VSS.n1364 2.6005
R4445 VSS.n1369 VSS.n1368 2.6005
R4446 VSS.n1368 VSS.n1367 2.6005
R4447 VSS.n1373 VSS.n1372 2.6005
R4448 VSS.n1372 VSS.n1371 2.6005
R4449 VSS.n1377 VSS.n1376 2.6005
R4450 VSS.n1376 VSS.n1375 2.6005
R4451 VSS.n1380 VSS.n1379 2.6005
R4452 VSS.n1379 VSS.n1378 2.6005
R4453 VSS.n1383 VSS.n1382 2.6005
R4454 VSS.n1382 VSS.n1381 2.6005
R4455 VSS.n1386 VSS.n1385 2.6005
R4456 VSS.n1385 VSS.n1384 2.6005
R4457 VSS.n1389 VSS.n1388 2.6005
R4458 VSS.n1388 VSS.n1387 2.6005
R4459 VSS.n1392 VSS.n1391 2.6005
R4460 VSS.n1391 VSS.n1390 2.6005
R4461 VSS.n1397 VSS.n1396 2.6005
R4462 VSS.n1115 VSS.n1114 2.6005
R4463 VSS.n1114 VSS.n1113 2.6005
R4464 VSS.n1118 VSS.n1117 2.6005
R4465 VSS.n1117 VSS.n1116 2.6005
R4466 VSS.n1121 VSS.n1120 2.6005
R4467 VSS.n1120 VSS.n1119 2.6005
R4468 VSS.n1124 VSS.n1123 2.6005
R4469 VSS.n1123 VSS.n1122 2.6005
R4470 VSS.n1127 VSS.n1126 2.6005
R4471 VSS.n1126 VSS.n1125 2.6005
R4472 VSS.n1130 VSS.n1129 2.6005
R4473 VSS.n1129 VSS.n1128 2.6005
R4474 VSS.n1134 VSS.n1133 2.6005
R4475 VSS.n1133 VSS.n1132 2.6005
R4476 VSS.n1138 VSS.n1137 2.6005
R4477 VSS.n1137 VSS.n1136 2.6005
R4478 VSS.n1141 VSS.n1140 2.6005
R4479 VSS.n1140 VSS.n1139 2.6005
R4480 VSS.n1144 VSS.n1143 2.6005
R4481 VSS.n1143 VSS.n1142 2.6005
R4482 VSS.n1147 VSS.n1146 2.6005
R4483 VSS.n1146 VSS.n1145 2.6005
R4484 VSS.n1150 VSS.n1149 2.6005
R4485 VSS.n1149 VSS.n1148 2.6005
R4486 VSS.n1153 VSS.n1152 2.6005
R4487 VSS.n1152 VSS.n1151 2.6005
R4488 VSS.n1156 VSS.n1155 2.6005
R4489 VSS.n1155 VSS.n1154 2.6005
R4490 VSS.n1159 VSS.n1158 2.6005
R4491 VSS.n1158 VSS.n1157 2.6005
R4492 VSS.n1162 VSS.n1161 2.6005
R4493 VSS.n1161 VSS.n1160 2.6005
R4494 VSS.n1165 VSS.n1164 2.6005
R4495 VSS.n1164 VSS.n1163 2.6005
R4496 VSS.n1168 VSS.n1167 2.6005
R4497 VSS.n1167 VSS.n1166 2.6005
R4498 VSS.n1171 VSS.n1170 2.6005
R4499 VSS.n1170 VSS.n1169 2.6005
R4500 VSS.n1174 VSS.n1173 2.6005
R4501 VSS.n1173 VSS.n1172 2.6005
R4502 VSS.n1177 VSS.n1176 2.6005
R4503 VSS.n1176 VSS.n1175 2.6005
R4504 VSS.n1180 VSS.n1179 2.6005
R4505 VSS.n1179 VSS.n1178 2.6005
R4506 VSS.n1183 VSS.n1182 2.6005
R4507 VSS.n1182 VSS.n1181 2.6005
R4508 VSS.n1186 VSS.n1185 2.6005
R4509 VSS.n1185 VSS.n1184 2.6005
R4510 VSS.n1190 VSS.n1189 2.6005
R4511 VSS.n1189 VSS.n1188 2.6005
R4512 VSS.n1194 VSS.n1193 2.6005
R4513 VSS.n1193 VSS.n1192 2.6005
R4514 VSS.n1197 VSS.n1196 2.6005
R4515 VSS.n1196 VSS.n1195 2.6005
R4516 VSS.n1200 VSS.n1199 2.6005
R4517 VSS.n1199 VSS.n1198 2.6005
R4518 VSS.n1203 VSS.n1202 2.6005
R4519 VSS.n1202 VSS.n1201 2.6005
R4520 VSS.n1206 VSS.n1205 2.6005
R4521 VSS.n1205 VSS.n1204 2.6005
R4522 VSS.n1209 VSS.n1208 2.6005
R4523 VSS.n1208 VSS.n1207 2.6005
R4524 VSS.n1242 VSS.n1241 2.6005
R4525 VSS.n932 VSS.n931 2.6005
R4526 VSS.n931 VSS.n930 2.6005
R4527 VSS.n935 VSS.n934 2.6005
R4528 VSS.n934 VSS.n933 2.6005
R4529 VSS.n938 VSS.n937 2.6005
R4530 VSS.n937 VSS.n936 2.6005
R4531 VSS.n941 VSS.n940 2.6005
R4532 VSS.n940 VSS.n939 2.6005
R4533 VSS.n944 VSS.n943 2.6005
R4534 VSS.n943 VSS.n942 2.6005
R4535 VSS.n947 VSS.n946 2.6005
R4536 VSS.n946 VSS.n945 2.6005
R4537 VSS.n951 VSS.n950 2.6005
R4538 VSS.n950 VSS.n949 2.6005
R4539 VSS.n955 VSS.n954 2.6005
R4540 VSS.n954 VSS.n953 2.6005
R4541 VSS.n958 VSS.n957 2.6005
R4542 VSS.n957 VSS.n956 2.6005
R4543 VSS.n961 VSS.n960 2.6005
R4544 VSS.n960 VSS.n959 2.6005
R4545 VSS.n964 VSS.n963 2.6005
R4546 VSS.n963 VSS.n962 2.6005
R4547 VSS.n967 VSS.n966 2.6005
R4548 VSS.n966 VSS.n965 2.6005
R4549 VSS.n970 VSS.n969 2.6005
R4550 VSS.n969 VSS.n968 2.6005
R4551 VSS.n973 VSS.n972 2.6005
R4552 VSS.n972 VSS.n971 2.6005
R4553 VSS.n976 VSS.n975 2.6005
R4554 VSS.n975 VSS.n974 2.6005
R4555 VSS.n979 VSS.n978 2.6005
R4556 VSS.n978 VSS.n977 2.6005
R4557 VSS.n982 VSS.n981 2.6005
R4558 VSS.n981 VSS.n980 2.6005
R4559 VSS.n985 VSS.n984 2.6005
R4560 VSS.n984 VSS.n983 2.6005
R4561 VSS.n988 VSS.n987 2.6005
R4562 VSS.n987 VSS.n986 2.6005
R4563 VSS.n991 VSS.n990 2.6005
R4564 VSS.n990 VSS.n989 2.6005
R4565 VSS.n994 VSS.n993 2.6005
R4566 VSS.n993 VSS.n992 2.6005
R4567 VSS.n997 VSS.n996 2.6005
R4568 VSS.n996 VSS.n995 2.6005
R4569 VSS.n1000 VSS.n999 2.6005
R4570 VSS.n999 VSS.n998 2.6005
R4571 VSS.n1003 VSS.n1002 2.6005
R4572 VSS.n1002 VSS.n1001 2.6005
R4573 VSS.n1007 VSS.n1006 2.6005
R4574 VSS.n1006 VSS.n1005 2.6005
R4575 VSS.n1011 VSS.n1010 2.6005
R4576 VSS.n1010 VSS.n1009 2.6005
R4577 VSS.n1014 VSS.n1013 2.6005
R4578 VSS.n1013 VSS.n1012 2.6005
R4579 VSS.n1017 VSS.n1016 2.6005
R4580 VSS.n1016 VSS.n1015 2.6005
R4581 VSS.n1020 VSS.n1019 2.6005
R4582 VSS.n1019 VSS.n1018 2.6005
R4583 VSS.n1023 VSS.n1022 2.6005
R4584 VSS.n1022 VSS.n1021 2.6005
R4585 VSS.n1026 VSS.n1025 2.6005
R4586 VSS.n1025 VSS.n1024 2.6005
R4587 VSS.n1059 VSS.n1058 2.6005
R4588 VSS.n3793 VSS.t279 2.55687
R4589 VSS.n2734 VSS.n2733 2.43319
R4590 VSS.n219 VSS.n218 2.43319
R4591 VSS.n216 VSS.n215 2.43319
R4592 VSS.n213 VSS.n212 2.43319
R4593 VSS.n210 VSS.n209 2.43319
R4594 VSS.n207 VSS.n206 2.43319
R4595 VSS.n204 VSS.n203 2.43319
R4596 VSS.n201 VSS.n200 2.43319
R4597 VSS.n198 VSS.n197 2.43319
R4598 VSS.n195 VSS.n194 2.43319
R4599 VSS.n192 VSS.n191 2.43319
R4600 VSS.n189 VSS.n188 2.43319
R4601 VSS.n186 VSS.n185 2.43319
R4602 VSS.n183 VSS.n182 2.43319
R4603 VSS.n180 VSS.n179 2.43319
R4604 VSS.n177 VSS.n176 2.43319
R4605 VSS.n174 VSS.n173 2.43319
R4606 VSS.n171 VSS.n170 2.43319
R4607 VSS.n168 VSS.n167 2.43319
R4608 VSS.n634 VSS.n633 2.43319
R4609 VSS.n631 VSS.n630 2.43319
R4610 VSS.n628 VSS.n627 2.43319
R4611 VSS.n625 VSS.n624 2.43319
R4612 VSS.n622 VSS.n621 2.43319
R4613 VSS.n619 VSS.n618 2.43319
R4614 VSS.n616 VSS.n615 2.43319
R4615 VSS.n613 VSS.n612 2.43319
R4616 VSS.n610 VSS.n609 2.43319
R4617 VSS.n607 VSS.n606 2.43319
R4618 VSS.n604 VSS.n603 2.43319
R4619 VSS.n601 VSS.n600 2.43319
R4620 VSS.n598 VSS.n597 2.43319
R4621 VSS.n595 VSS.n594 2.43319
R4622 VSS.n592 VSS.n591 2.43319
R4623 VSS.n589 VSS.n588 2.43319
R4624 VSS.n586 VSS.n585 2.43319
R4625 VSS.n583 VSS.n582 2.43319
R4626 VSS.n2658 VSS.n2657 2.43319
R4627 VSS.n2655 VSS.n2654 2.43319
R4628 VSS.n1747 VSS.n1744 2.29321
R4629 VSS.n1617 VSS.n1614 2.29321
R4630 VSS.n1487 VSS.n1484 2.29321
R4631 VSS.n2714 VSS.n2711 2.18289
R4632 VSS.n2512 VSS.t23 2.13081
R4633 VSS.n2496 VSS.t26 2.13081
R4634 VSS.n3799 VSS.t253 2.13081
R4635 VSS.n3821 VSS.t519 2.13081
R4636 VSS.n2170 VSS.n2169 2.08372
R4637 VSS.n2700 VSS.n2696 2.07475
R4638 VSS.n2680 VSS.n2676 2.07475
R4639 VSS.n1748 VSS.n1747 1.9805
R4640 VSS.n1618 VSS.n1617 1.9805
R4641 VSS.n1488 VSS.n1487 1.9805
R4642 VSS.n1702 VSS.n1699 1.96158
R4643 VSS.n1722 VSS.n1719 1.96158
R4644 VSS.n1572 VSS.n1569 1.96158
R4645 VSS.n1592 VSS.n1589 1.96158
R4646 VSS.n1442 VSS.n1439 1.96158
R4647 VSS.n1462 VSS.n1459 1.96158
R4648 VSS.n1727 VSS.n1726 1.95148
R4649 VSS.n1597 VSS.n1596 1.95148
R4650 VSS.n1467 VSS.n1466 1.95148
R4651 VSS.n1758 VSS.n1757 1.91002
R4652 VSS.n1734 VSS.n1733 1.91002
R4653 VSS.n1628 VSS.n1627 1.91002
R4654 VSS.n1604 VSS.n1603 1.91002
R4655 VSS.n1498 VSS.n1497 1.91002
R4656 VSS.n1474 VSS.n1473 1.91002
R4657 VSS.n1763 VSS.n1760 1.90218
R4658 VSS.n1633 VSS.n1630 1.90218
R4659 VSS.n1503 VSS.n1500 1.90218
R4660 VSS.n1728 VSS.n1727 1.89955
R4661 VSS.n1598 VSS.n1597 1.89955
R4662 VSS.n1468 VSS.n1467 1.89955
R4663 VSS.n758 VSS.n757 1.8318
R4664 VSS.n1674 VSS.n1673 1.8318
R4665 VSS.n764 VSS.n763 1.8318
R4666 VSS.n1680 VSS.n1679 1.8318
R4667 VSS.n495 VSS.n494 1.8318
R4668 VSS.n1640 VSS.n1639 1.8318
R4669 VSS.n501 VSS.n500 1.8318
R4670 VSS.n1646 VSS.n1645 1.8318
R4671 VSS.n485 VSS.n484 1.8318
R4672 VSS.n1544 VSS.n1543 1.8318
R4673 VSS.n491 VSS.n490 1.8318
R4674 VSS.n1550 VSS.n1549 1.8318
R4675 VSS.n80 VSS.n79 1.8318
R4676 VSS.n1510 VSS.n1509 1.8318
R4677 VSS.n86 VSS.n85 1.8318
R4678 VSS.n1516 VSS.n1515 1.8318
R4679 VSS.n70 VSS.n69 1.8318
R4680 VSS.n1414 VSS.n1413 1.8318
R4681 VSS.n76 VSS.n75 1.8318
R4682 VSS.n1420 VSS.n1419 1.8318
R4683 VSS.n774 VSS.n773 1.8318
R4684 VSS.n1806 VSS.n1805 1.8318
R4685 VSS.n768 VSS.n767 1.8318
R4686 VSS.n1772 VSS.n1771 1.8318
R4687 VSS.n1766 VSS.n1765 1.76495
R4688 VSS.n1636 VSS.n1635 1.76495
R4689 VSS.n1506 VSS.n1505 1.76495
R4690 VSS.n2486 VSS.t497 1.70475
R4691 VSS.n2487 VSS.t262 1.70475
R4692 VSS.t255 VSS.t44 1.70475
R4693 VSS.n2299 VSS.n2298 1.68702
R4694 VSS.n2305 VSS.n2304 1.68702
R4695 VSS.n289 VSS.n288 1.68702
R4696 VSS.n288 VSS.n287 1.68702
R4697 VSS.n3541 VSS.n3540 1.68702
R4698 VSS.n3542 VSS.n3541 1.68702
R4699 VSS.n3543 VSS.n3542 1.68702
R4700 VSS.n286 VSS.n285 1.68702
R4701 VSS.n285 VSS.n284 1.68702
R4702 VSS.n3759 VSS.n3756 1.68702
R4703 VSS.n3762 VSS.n3759 1.68702
R4704 VSS.n3765 VSS.n3762 1.68702
R4705 VSS.n3768 VSS.n3765 1.68702
R4706 VSS.n277 VSS.n276 1.68702
R4707 VSS.n276 VSS.n275 1.68702
R4708 VSS.n3522 VSS.n3519 1.68702
R4709 VSS.n3525 VSS.n3522 1.68702
R4710 VSS.n3528 VSS.n3525 1.68702
R4711 VSS.n3531 VSS.n3528 1.68702
R4712 VSS.n268 VSS.n267 1.68702
R4713 VSS.n267 VSS.n266 1.68702
R4714 VSS.n3507 VSS.n3504 1.68702
R4715 VSS.n3510 VSS.n3507 1.68702
R4716 VSS.n3513 VSS.n3510 1.68702
R4717 VSS.n3516 VSS.n3513 1.68702
R4718 VSS.n259 VSS.n258 1.68702
R4719 VSS.n258 VSS.n257 1.68702
R4720 VSS.n3492 VSS.n3489 1.68702
R4721 VSS.n3495 VSS.n3492 1.68702
R4722 VSS.n3498 VSS.n3495 1.68702
R4723 VSS.n3501 VSS.n3498 1.68702
R4724 VSS.n250 VSS.n249 1.68702
R4725 VSS.n249 VSS.n248 1.68702
R4726 VSS.n3482 VSS.n3481 1.68702
R4727 VSS.n3483 VSS.n3482 1.68702
R4728 VSS.n3484 VSS.n3483 1.68702
R4729 VSS.n247 VSS.n246 1.68702
R4730 VSS.n246 VSS.n245 1.68702
R4731 VSS.n3476 VSS.n3475 1.68702
R4732 VSS.n3477 VSS.n3476 1.68702
R4733 VSS.n3478 VSS.n3477 1.68702
R4734 VSS.n310 VSS.n309 1.68702
R4735 VSS.n309 VSS.n308 1.68702
R4736 VSS.n3533 VSS.n3532 1.68702
R4737 VSS.n3534 VSS.n3533 1.68702
R4738 VSS.n3535 VSS.n3534 1.68702
R4739 VSS.n2429 VSS.n2428 1.68702
R4740 VSS.n2309 VSS.n2308 1.68702
R4741 VSS.n477 VSS.n476 1.65879
R4742 VSS.n472 VSS.n471 1.65879
R4743 VSS.n467 VSS.n466 1.65879
R4744 VSS.n462 VSS.n461 1.65879
R4745 VSS.n457 VSS.n456 1.65879
R4746 VSS.n750 VSS.n749 1.65879
R4747 VSS.n745 VSS.n744 1.65879
R4748 VSS.n740 VSS.n739 1.65879
R4749 VSS.n735 VSS.n734 1.65879
R4750 VSS.n730 VSS.n729 1.65879
R4751 VSS.n893 VSS.n892 1.65879
R4752 VSS.n888 VSS.n887 1.65879
R4753 VSS.n883 VSS.n882 1.65879
R4754 VSS.n878 VSS.n877 1.65879
R4755 VSS.n873 VSS.n872 1.65879
R4756 VSS.n868 VSS.n867 1.65879
R4757 VSS.n3143 VSS.n3142 1.65879
R4758 VSS.n3723 VSS.n3721 1.65879
R4759 VSS.n3720 VSS.n3718 1.65879
R4760 VSS.n3717 VSS.n3715 1.65879
R4761 VSS.n3714 VSS.n3712 1.65879
R4762 VSS.n3711 VSS.n3709 1.65879
R4763 VSS.n3708 VSS.n3706 1.65879
R4764 VSS.n3705 VSS.n3703 1.65879
R4765 VSS.n3702 VSS.n3700 1.65879
R4766 VSS.n3699 VSS.n3697 1.65879
R4767 VSS.n3696 VSS.n3695 1.65879
R4768 VSS.n3924 VSS.n3923 1.65879
R4769 VSS.n3919 VSS.n3918 1.65879
R4770 VSS.n3914 VSS.n3913 1.65879
R4771 VSS.n3909 VSS.n3908 1.65879
R4772 VSS.n3904 VSS.n3903 1.65879
R4773 VSS.n3899 VSS.n3898 1.65879
R4774 VSS.n2584 VSS.n2583 1.65879
R4775 VSS.n2579 VSS.n2578 1.65879
R4776 VSS.n2574 VSS.n2573 1.65879
R4777 VSS.n3367 VSS.n3366 1.65879
R4778 VSS.n3362 VSS.n3361 1.65879
R4779 VSS.n3357 VSS.n3356 1.65879
R4780 VSS.n3352 VSS.n3351 1.65879
R4781 VSS.n3347 VSS.n3346 1.65879
R4782 VSS.n3342 VSS.n3341 1.65879
R4783 VSS.n3337 VSS.n3336 1.65879
R4784 VSS.n2167 VSS.n2144 1.65879
R4785 VSS.n2141 VSS.n2140 1.65879
R4786 VSS.n2136 VSS.n2135 1.65879
R4787 VSS.n2131 VSS.n2130 1.65879
R4788 VSS.n2126 VSS.n2125 1.65879
R4789 VSS.n2121 VSS.n2120 1.65879
R4790 VSS.n2116 VSS.n2115 1.65879
R4791 VSS.n2111 VSS.n2110 1.65879
R4792 VSS.n2106 VSS.n2105 1.65879
R4793 VSS.n2101 VSS.n2100 1.65879
R4794 VSS.n3138 VSS.n3137 1.65822
R4795 VSS.n2375 VSS.n2374 1.65822
R4796 VSS.n2380 VSS.n2379 1.65822
R4797 VSS.n2385 VSS.n2384 1.65822
R4798 VSS.n2390 VSS.n2389 1.65822
R4799 VSS.n2395 VSS.n2394 1.65822
R4800 VSS.n3729 VSS.n3728 1.65822
R4801 VSS.n3670 VSS.n3669 1.65822
R4802 VSS.n3665 VSS.n3664 1.65822
R4803 VSS.n3660 VSS.n3659 1.65822
R4804 VSS.n3655 VSS.n3654 1.65822
R4805 VSS.n3650 VSS.n3649 1.65822
R4806 VSS.n3645 VSS.n3644 1.65822
R4807 VSS.n3699 VSS.n3698 1.65822
R4808 VSS.n3702 VSS.n3701 1.65822
R4809 VSS.n3705 VSS.n3704 1.65822
R4810 VSS.n3708 VSS.n3707 1.65822
R4811 VSS.n3711 VSS.n3710 1.65822
R4812 VSS.n3714 VSS.n3713 1.65822
R4813 VSS.n3717 VSS.n3716 1.65822
R4814 VSS.n3720 VSS.n3719 1.65822
R4815 VSS.n3723 VSS.n3722 1.65822
R4816 VSS.n3894 VSS.n3893 1.65822
R4817 VSS.n2994 VSS.n2993 1.65811
R4818 VSS.n2999 VSS.n2998 1.65811
R4819 VSS.n3004 VSS.n3003 1.65811
R4820 VSS.n2988 VSS.n2987 1.65811
R4821 VSS.n4041 VSS.n4040 1.65811
R4822 VSS.n4036 VSS.n4035 1.65811
R4823 VSS.n4031 VSS.n4030 1.65811
R4824 VSS.n4026 VSS.n4025 1.65811
R4825 VSS.n4021 VSS.n4020 1.65811
R4826 VSS.n4016 VSS.n4015 1.65811
R4827 VSS.n4011 VSS.n4010 1.65811
R4828 VSS.n4006 VSS.n4005 1.65811
R4829 VSS.n2274 VSS.n2273 1.65811
R4830 VSS.n2279 VSS.n2278 1.65811
R4831 VSS.n2284 VSS.n2283 1.65811
R4832 VSS.n2289 VSS.n2288 1.65811
R4833 VSS.n2294 VSS.n2293 1.65811
R4834 VSS.n244 VSS.n243 1.65811
R4835 VSS.n3467 VSS.n3465 1.65811
R4836 VSS.n3464 VSS.n3462 1.65811
R4837 VSS.n3464 VSS.n3463 1.65811
R4838 VSS.n3461 VSS.n3460 1.65811
R4839 VSS.n3467 VSS.n3466 1.65811
R4840 VSS.n2946 VSS.t391 1.6385
R4841 VSS.n2867 VSS.t382 1.6385
R4842 VSS.n2868 VSS.t297 1.6385
R4843 VSS.n2869 VSS.t455 1.6385
R4844 VSS.n2870 VSS.t474 1.6385
R4845 VSS.n2872 VSS.t288 1.6385
R4846 VSS.n2872 VSS.n2871 1.6385
R4847 VSS.n2874 VSS.t254 1.6385
R4848 VSS.n2874 VSS.n2873 1.6385
R4849 VSS.n3847 VSS.t518 1.6385
R4850 VSS.n3847 VSS.n3846 1.6385
R4851 VSS.n3845 VSS.t628 1.6385
R4852 VSS.n3845 VSS.n3844 1.6385
R4853 VSS.n3843 VSS.t626 1.6385
R4854 VSS.n3843 VSS.n3842 1.6385
R4855 VSS.n2532 VSS.t366 1.6385
R4856 VSS.n2532 VSS.n2531 1.6385
R4857 VSS.n2534 VSS.t36 1.6385
R4858 VSS.n2534 VSS.n2533 1.6385
R4859 VSS.n2536 VSS.t38 1.6385
R4860 VSS.n2536 VSS.n2535 1.6385
R4861 VSS.n2538 VSS.t40 1.6385
R4862 VSS.n2538 VSS.n2537 1.6385
R4863 VSS.n2540 VSS.t568 1.6385
R4864 VSS.n2540 VSS.n2539 1.6385
R4865 VSS.n2542 VSS.t45 1.6385
R4866 VSS.n2542 VSS.n2541 1.6385
R4867 VSS.n2544 VSS.t225 1.6385
R4868 VSS.n2544 VSS.n2543 1.6385
R4869 VSS.n2546 VSS.t501 1.6385
R4870 VSS.n2546 VSS.n2545 1.6385
R4871 VSS.n2548 VSS.t259 1.6385
R4872 VSS.n2548 VSS.n2547 1.6385
R4873 VSS.n363 VSS 1.59665
R4874 VSS VSS.n362 1.59578
R4875 VSS.n4094 VSS.t56 1.53406
R4876 VSS.n3750 VSS.t5 1.53406
R4877 VSS.n1699 VSS.n1698 1.48796
R4878 VSS.n1687 VSS.n1686 1.48796
R4879 VSS.n1719 VSS.n1718 1.48796
R4880 VSS.n1707 VSS.n1706 1.48796
R4881 VSS.n1569 VSS.n1568 1.48796
R4882 VSS.n1557 VSS.n1556 1.48796
R4883 VSS.n1589 VSS.n1588 1.48796
R4884 VSS.n1577 VSS.n1576 1.48796
R4885 VSS.n1439 VSS.n1438 1.48796
R4886 VSS.n1427 VSS.n1426 1.48796
R4887 VSS.n1459 VSS.n1458 1.48796
R4888 VSS.n1447 VSS.n1446 1.48796
R4889 VSS.n1691 VSS.n1690 1.47979
R4890 VSS.n1711 VSS.n1710 1.47979
R4891 VSS.n1731 VSS.n1730 1.47979
R4892 VSS.n1740 VSS.n1739 1.47979
R4893 VSS.n1755 VSS.n1754 1.47979
R4894 VSS.n1561 VSS.n1560 1.47979
R4895 VSS.n1601 VSS.n1600 1.47979
R4896 VSS.n1610 VSS.n1609 1.47979
R4897 VSS.n1625 VSS.n1624 1.47979
R4898 VSS.n1581 VSS.n1580 1.47979
R4899 VSS.n1431 VSS.n1430 1.47979
R4900 VSS.n1451 VSS.n1450 1.47979
R4901 VSS.n1471 VSS.n1470 1.47979
R4902 VSS.n1480 VSS.n1479 1.47979
R4903 VSS.n1495 VSS.n1494 1.47979
R4904 VSS.n2709 VSS.n2708 1.40389
R4905 VSS.n2729 VSS.n2728 1.40389
R4906 VSS.n2661 VSS.n2660 1.40389
R4907 VSS.n2737 VSS.n2736 1.40375
R4908 VSS.n1402 VSS.n1401 1.40375
R4909 VSS.n1405 VSS.n1404 1.40375
R4910 VSS.n1410 VSS.n1409 1.40375
R4911 VSS.n480 VSS.n479 1.40375
R4912 VSS.n753 VSS.n752 1.40375
R4913 VSS.n2644 VSS.n2643 1.40375
R4914 VSS.n1290 VSS.n1248 1.38491
R4915 VSS.n1290 VSS.n1249 1.38491
R4916 VSS.n1290 VSS.n1250 1.38491
R4917 VSS.n1290 VSS.n1251 1.38491
R4918 VSS.n1290 VSS.n1252 1.38491
R4919 VSS.n1290 VSS.n1253 1.38491
R4920 VSS.n1290 VSS.n1254 1.38491
R4921 VSS.n1290 VSS.n1255 1.38491
R4922 VSS.n1290 VSS.n1256 1.38491
R4923 VSS.n1290 VSS.n1257 1.38491
R4924 VSS.n1290 VSS.n1258 1.38491
R4925 VSS.n1290 VSS.n1259 1.38491
R4926 VSS.n1290 VSS.n1260 1.38491
R4927 VSS.n1290 VSS.n1261 1.38491
R4928 VSS.n1290 VSS.n1262 1.38491
R4929 VSS.n1290 VSS.n1263 1.38491
R4930 VSS.n1290 VSS.n1264 1.38491
R4931 VSS.n1290 VSS.n1265 1.38491
R4932 VSS.n1290 VSS.n1266 1.38491
R4933 VSS.n1290 VSS.n1267 1.38491
R4934 VSS.n1290 VSS.n1268 1.38491
R4935 VSS.n1290 VSS.n1269 1.38491
R4936 VSS.n1290 VSS.n1270 1.38491
R4937 VSS.n1290 VSS.n1271 1.38491
R4938 VSS.n1290 VSS.n1272 1.38491
R4939 VSS.n1290 VSS.n1273 1.38491
R4940 VSS.n1290 VSS.n1274 1.38491
R4941 VSS.n1290 VSS.n1275 1.38491
R4942 VSS.n1290 VSS.n1276 1.38491
R4943 VSS.n1290 VSS.n1277 1.38491
R4944 VSS.n1290 VSS.n1278 1.38491
R4945 VSS.n1290 VSS.n1279 1.38491
R4946 VSS.n1290 VSS.n1280 1.38491
R4947 VSS.n1290 VSS.n1281 1.38491
R4948 VSS.n1290 VSS.n1282 1.38491
R4949 VSS.n1290 VSS.n1283 1.38491
R4950 VSS.n1290 VSS.n1284 1.38491
R4951 VSS.n1290 VSS.n1285 1.38491
R4952 VSS.n1290 VSS.n1286 1.38491
R4953 VSS.n1290 VSS.n1287 1.38491
R4954 VSS.n1290 VSS.n1288 1.38491
R4955 VSS.n1290 VSS.n1289 1.38491
R4956 VSS.n1107 VSS.n1065 1.38491
R4957 VSS.n1107 VSS.n1066 1.38491
R4958 VSS.n1107 VSS.n1067 1.38491
R4959 VSS.n1107 VSS.n1068 1.38491
R4960 VSS.n1107 VSS.n1069 1.38491
R4961 VSS.n1107 VSS.n1070 1.38491
R4962 VSS.n1107 VSS.n1071 1.38491
R4963 VSS.n1107 VSS.n1072 1.38491
R4964 VSS.n1107 VSS.n1073 1.38491
R4965 VSS.n1107 VSS.n1074 1.38491
R4966 VSS.n1107 VSS.n1075 1.38491
R4967 VSS.n1107 VSS.n1076 1.38491
R4968 VSS.n1107 VSS.n1077 1.38491
R4969 VSS.n1107 VSS.n1078 1.38491
R4970 VSS.n1107 VSS.n1079 1.38491
R4971 VSS.n1107 VSS.n1080 1.38491
R4972 VSS.n1107 VSS.n1081 1.38491
R4973 VSS.n1107 VSS.n1082 1.38491
R4974 VSS.n1107 VSS.n1083 1.38491
R4975 VSS.n1107 VSS.n1084 1.38491
R4976 VSS.n1107 VSS.n1085 1.38491
R4977 VSS.n1107 VSS.n1086 1.38491
R4978 VSS.n1107 VSS.n1087 1.38491
R4979 VSS.n1107 VSS.n1088 1.38491
R4980 VSS.n1107 VSS.n1089 1.38491
R4981 VSS.n1107 VSS.n1090 1.38491
R4982 VSS.n1107 VSS.n1091 1.38491
R4983 VSS.n1107 VSS.n1092 1.38491
R4984 VSS.n1107 VSS.n1093 1.38491
R4985 VSS.n1107 VSS.n1094 1.38491
R4986 VSS.n1107 VSS.n1095 1.38491
R4987 VSS.n1107 VSS.n1096 1.38491
R4988 VSS.n1107 VSS.n1097 1.38491
R4989 VSS.n1107 VSS.n1098 1.38491
R4990 VSS.n1107 VSS.n1099 1.38491
R4991 VSS.n1107 VSS.n1100 1.38491
R4992 VSS.n1107 VSS.n1101 1.38491
R4993 VSS.n1107 VSS.n1102 1.38491
R4994 VSS.n1107 VSS.n1103 1.38491
R4995 VSS.n1107 VSS.n1104 1.38491
R4996 VSS.n1107 VSS.n1105 1.38491
R4997 VSS.n1107 VSS.n1106 1.38491
R4998 VSS.n3377 VSS.n3371 1.38491
R4999 VSS.n3377 VSS.n3372 1.38491
R5000 VSS.n3377 VSS.n3373 1.38491
R5001 VSS.n3377 VSS.n3374 1.38491
R5002 VSS.n3377 VSS.n3375 1.38491
R5003 VSS.n3377 VSS.n3376 1.38491
R5004 VSS.n1688 VSS.n1687 1.3649
R5005 VSS.n1708 VSS.n1707 1.3649
R5006 VSS.n1558 VSS.n1557 1.3649
R5007 VSS.n1578 VSS.n1577 1.3649
R5008 VSS.n1428 VSS.n1427 1.3649
R5009 VSS.n1448 VSS.n1447 1.3649
R5010 VSS.n3128 VSS.n3125 1.3543
R5011 VSS.n3726 VSS.n3724 1.3543
R5012 VSS.n2022 VSS.n2020 1.3543
R5013 VSS.n1946 VSS.n1944 1.3543
R5014 VSS.n1868 VSS.n1866 1.3543
R5015 VSS.n3726 VSS.n3725 1.35379
R5016 VSS.n3324 VSS.n3317 1.35379
R5017 VSS.n3930 VSS.n3929 1.35379
R5018 VSS.n3379 VSS.n3378 1.35379
R5019 VSS.n2416 VSS.n2415 1.35379
R5020 VSS.n2022 VSS.n2021 1.35379
R5021 VSS.n1946 VSS.n1945 1.35379
R5022 VSS.n1868 VSS.n1867 1.35379
R5023 VSS.n3469 VSS.n3468 1.35364
R5024 VSS.n4056 VSS.n4055 1.35364
R5025 VSS.n3472 VSS.n3471 1.35364
R5026 VSS.n959 VSS.t98 1.3127
R5027 VSS.n995 VSS.t75 1.3127
R5028 VSS.n1142 VSS.t70 1.3127
R5029 VSS.n1178 VSS.t84 1.3127
R5030 VSS.n1325 VSS.t80 1.3127
R5031 VSS.n1361 VSS.t67 1.3127
R5032 VSS.n1812 VSS.n1774 1.30746
R5033 VSS.n1004 VSS.n766 1.30746
R5034 VSS.n1008 VSS.n762 1.30746
R5035 VSS.n1848 VSS.n1682 1.30746
R5036 VSS.n1851 VSS.n1678 1.30746
R5037 VSS.n1131 VSS.n503 1.30746
R5038 VSS.n1135 VSS.n499 1.30746
R5039 VSS.n1887 VSS.n1648 1.30746
R5040 VSS.n1890 VSS.n1644 1.30746
R5041 VSS.n1187 VSS.n493 1.30746
R5042 VSS.n1191 VSS.n489 1.30746
R5043 VSS.n1926 VSS.n1552 1.30746
R5044 VSS.n1929 VSS.n1548 1.30746
R5045 VSS.n1314 VSS.n88 1.30746
R5046 VSS.n1318 VSS.n84 1.30746
R5047 VSS.n1965 VSS.n1518 1.30746
R5048 VSS.n1968 VSS.n1514 1.30746
R5049 VSS.n1370 VSS.n78 1.30746
R5050 VSS.n1374 VSS.n74 1.30746
R5051 VSS.n2004 VSS.n1422 1.30746
R5052 VSS.n2007 VSS.n1418 1.30746
R5053 VSS.n3280 VSS.n3012 1.30746
R5054 VSS.n3269 VSS.n3018 1.30746
R5055 VSS.n3203 VSS.n3035 1.30746
R5056 VSS.n3181 VSS.n3040 1.30746
R5057 VSS.n3162 VSS.n3046 1.30746
R5058 VSS.n3152 VSS.n3048 1.30746
R5059 VSS.n2743 VSS.n2706 1.30746
R5060 VSS.n2750 VSS.n2704 1.30746
R5061 VSS.n3228 VSS.n3030 1.30746
R5062 VSS.n2795 VSS.n2690 1.30746
R5063 VSS.n3247 VSS.n3024 1.30746
R5064 VSS.n2808 VSS.n2687 1.30746
R5065 VSS.n3294 VSS.n3009 1.30746
R5066 VSS.n3284 VSS.n3011 1.30746
R5067 VSS.n2831 VSS.n2684 1.30746
R5068 VSS.n2838 VSS.n2682 1.30746
R5069 VSS.n1809 VSS.n1808 1.30746
R5070 VSS.n952 VSS.n772 1.30746
R5071 VSS.n948 VSS.n776 1.30746
R5072 VSS.n1737 VSS.n1736 1.3055
R5073 VSS.n1607 VSS.n1606 1.3055
R5074 VSS.n1477 VSS.n1476 1.3055
R5075 VSS.n1749 VSS.n1748 1.29992
R5076 VSS.n1619 VSS.n1618 1.29992
R5077 VSS.n1489 VSS.n1488 1.29992
R5078 VSS.n3166 VSS.t16 1.27869
R5079 VSS.n3241 VSS.t527 1.27869
R5080 VSS.n2612 VSS.t221 1.27869
R5081 VSS.n3965 VSS.t59 1.27869
R5082 VSS.n4059 VSS.n4058 1.2071
R5083 VSS.n3382 VSS.n3381 1.20692
R5084 VSS.n2565 VSS.n2556 1.19007
R5085 VSS.n2556 VSS.n2555 1.19007
R5086 VSS.n4060 VSS.n4059 1.12625
R5087 VSS.n3383 VSS.n3382 1.12625
R5088 VSS.n1696 VSS.n1695 1.1255
R5089 VSS.n1716 VSS.n1715 1.1255
R5090 VSS.n1736 VSS.n1735 1.1255
R5091 VSS.n1751 VSS.n1750 1.1255
R5092 VSS.n1760 VSS.n1759 1.1255
R5093 VSS.n1566 VSS.n1565 1.1255
R5094 VSS.n1606 VSS.n1605 1.1255
R5095 VSS.n1621 VSS.n1620 1.1255
R5096 VSS.n1630 VSS.n1629 1.1255
R5097 VSS.n1586 VSS.n1585 1.1255
R5098 VSS.n1436 VSS.n1435 1.1255
R5099 VSS.n1456 VSS.n1455 1.1255
R5100 VSS.n1476 VSS.n1475 1.1255
R5101 VSS.n1491 VSS.n1490 1.1255
R5102 VSS.n1500 VSS.n1499 1.1255
R5103 VSS.n305 VSS.n289 1.12354
R5104 VSS.n318 VSS.n286 1.12354
R5105 VSS.n327 VSS.n277 1.12354
R5106 VSS.n334 VSS.n268 1.12354
R5107 VSS.n343 VSS.n259 1.12354
R5108 VSS.n350 VSS.n250 1.12354
R5109 VSS.n353 VSS.n247 1.12354
R5110 VSS.n311 VSS.n310 1.12354
R5111 VSS.n4070 VSS.n3531 1.12159
R5112 VSS.n4080 VSS.n3516 1.12159
R5113 VSS.n4093 VSS.n3501 1.12159
R5114 VSS.n4107 VSS.n3480 1.12159
R5115 VSS.n4103 VSS.n3486 1.12159
R5116 VSS.n3743 VSS.n3539 1.12159
R5117 VSS.n3739 VSS.n3545 1.12159
R5118 VSS.n3769 VSS.n3768 1.10202
R5119 VSS.n2628 VSS.n2627 1.09195
R5120 VSS.n1789 VSS.n1788 1.09195
R5121 VSS.n64 VSS.n0 1.08441
R5122 VSS.n59 VSS.n1 1.08441
R5123 VSS.n3420 VSS.n2307 1.08441
R5124 VSS.n3427 VSS.n2303 1.08441
R5125 VSS.n2421 VSS.n2311 1.08441
R5126 VSS.n11 VSS.n2 1.08441
R5127 VSS.n2434 VSS.n2433 1.08441
R5128 VSS.n6 VSS.n3 1.08441
R5129 VSS.n3018 VSS.n3017 1.0492
R5130 VSS.n3046 VSS.n3045 1.0492
R5131 VSS.n3048 VSS.n3047 1.0492
R5132 VSS.n3030 VSS.n3029 1.0492
R5133 VSS.n3024 VSS.n3023 1.0492
R5134 VSS.n3009 VSS.n3008 1.0492
R5135 VSS.n3011 VSS.n3010 1.0492
R5136 VSS.n3780 VSS.n3779 1.0492
R5137 VSS.n3779 VSS.n3778 1.0492
R5138 VSS.n3778 VSS.n3777 1.0492
R5139 VSS.n3786 VSS.n3785 1.0492
R5140 VSS.n3785 VSS.n3784 1.0492
R5141 VSS.n3784 VSS.n3783 1.0492
R5142 VSS.n2479 VSS.n2478 1.0492
R5143 VSS.n2478 VSS.n2477 1.0492
R5144 VSS.n2477 VSS.n2476 1.0492
R5145 VSS.n2473 VSS.n2472 1.0492
R5146 VSS.n2472 VSS.n2471 1.0492
R5147 VSS.n2471 VSS.n2470 1.0492
R5148 VSS.n2715 VSS.n2714 1.00704
R5149 VSS.n1727 VSS.n1724 0.95333
R5150 VSS.n1597 VSS.n1594 0.95333
R5151 VSS.n1467 VSS.n1464 0.95333
R5152 VSS.n1702 VSS.n1701 0.949983
R5153 VSS.n1722 VSS.n1721 0.949983
R5154 VSS.n1763 VSS.n1762 0.949983
R5155 VSS.n1572 VSS.n1571 0.949983
R5156 VSS.n1633 VSS.n1632 0.949983
R5157 VSS.n1592 VSS.n1591 0.949983
R5158 VSS.n1442 VSS.n1441 0.949983
R5159 VSS.n1462 VSS.n1461 0.949983
R5160 VSS.n1503 VSS.n1502 0.949983
R5161 VSS.n2696 VSS.n2695 0.890378
R5162 VSS.n2676 VSS.n2675 0.890378
R5163 VSS.n1774 VSS.n1773 0.871152
R5164 VSS.n766 VSS.n765 0.871152
R5165 VSS.n762 VSS.n761 0.871152
R5166 VSS.n761 VSS.n758 0.871152
R5167 VSS.n1677 VSS.n1674 0.871152
R5168 VSS.n765 VSS.n764 0.871152
R5169 VSS.n1681 VSS.n1680 0.871152
R5170 VSS.n1682 VSS.n1681 0.871152
R5171 VSS.n1678 VSS.n1677 0.871152
R5172 VSS.n503 VSS.n502 0.871152
R5173 VSS.n499 VSS.n498 0.871152
R5174 VSS.n498 VSS.n495 0.871152
R5175 VSS.n1643 VSS.n1640 0.871152
R5176 VSS.n502 VSS.n501 0.871152
R5177 VSS.n1647 VSS.n1646 0.871152
R5178 VSS.n1648 VSS.n1647 0.871152
R5179 VSS.n1644 VSS.n1643 0.871152
R5180 VSS.n493 VSS.n492 0.871152
R5181 VSS.n489 VSS.n488 0.871152
R5182 VSS.n488 VSS.n485 0.871152
R5183 VSS.n1547 VSS.n1544 0.871152
R5184 VSS.n492 VSS.n491 0.871152
R5185 VSS.n1551 VSS.n1550 0.871152
R5186 VSS.n1552 VSS.n1551 0.871152
R5187 VSS.n1548 VSS.n1547 0.871152
R5188 VSS.n88 VSS.n87 0.871152
R5189 VSS.n84 VSS.n83 0.871152
R5190 VSS.n83 VSS.n80 0.871152
R5191 VSS.n1513 VSS.n1510 0.871152
R5192 VSS.n87 VSS.n86 0.871152
R5193 VSS.n1517 VSS.n1516 0.871152
R5194 VSS.n1518 VSS.n1517 0.871152
R5195 VSS.n1514 VSS.n1513 0.871152
R5196 VSS.n78 VSS.n77 0.871152
R5197 VSS.n74 VSS.n73 0.871152
R5198 VSS.n73 VSS.n70 0.871152
R5199 VSS.n1417 VSS.n1414 0.871152
R5200 VSS.n77 VSS.n76 0.871152
R5201 VSS.n1421 VSS.n1420 0.871152
R5202 VSS.n1422 VSS.n1421 0.871152
R5203 VSS.n1418 VSS.n1417 0.871152
R5204 VSS.n775 VSS.n774 0.871152
R5205 VSS.n1807 VSS.n1806 0.871152
R5206 VSS.n1808 VSS.n1807 0.871152
R5207 VSS.n772 VSS.n771 0.871152
R5208 VSS.n771 VSS.n768 0.871152
R5209 VSS.n1773 VSS.n1772 0.871152
R5210 VSS.n776 VSS.n775 0.871152
R5211 VSS.n3013 VSS.t547 0.8195
R5212 VSS.n3014 VSS.t546 0.8195
R5213 VSS.n3016 VSS.t564 0.8195
R5214 VSS.n3016 VSS.n3015 0.8195
R5215 VSS.n3032 VSS.t559 0.8195
R5216 VSS.n3032 VSS.n3031 0.8195
R5217 VSS.n3034 VSS.t20 0.8195
R5218 VSS.n3034 VSS.n3033 0.8195
R5219 VSS.n3037 VSS.t617 0.8195
R5220 VSS.n3037 VSS.n3036 0.8195
R5221 VSS.n3039 VSS.t15 0.8195
R5222 VSS.n3039 VSS.n3038 0.8195
R5223 VSS.n2703 VSS.t344 0.8195
R5224 VSS.n2703 VSS.n2702 0.8195
R5225 VSS.n3044 VSS.t368 0.8195
R5226 VSS.n3044 VSS.n3043 0.8195
R5227 VSS.n3042 VSS.t379 0.8195
R5228 VSS.n3042 VSS.n3041 0.8195
R5229 VSS.n2694 VSS.t616 0.8195
R5230 VSS.n2694 VSS.n2693 0.8195
R5231 VSS.n2692 VSS.t29 0.8195
R5232 VSS.n2692 VSS.n2691 0.8195
R5233 VSS.n2689 VSS.t246 0.8195
R5234 VSS.n2689 VSS.n2688 0.8195
R5235 VSS.n3028 VSS.t533 0.8195
R5236 VSS.n3028 VSS.n3027 0.8195
R5237 VSS.n3026 VSS.t534 0.8195
R5238 VSS.n3026 VSS.n3025 0.8195
R5239 VSS.n2686 VSS.t528 0.8195
R5240 VSS.n2686 VSS.n2685 0.8195
R5241 VSS.n3022 VSS.t531 0.8195
R5242 VSS.n3022 VSS.n3021 0.8195
R5243 VSS.n3020 VSS.t532 0.8195
R5244 VSS.n3020 VSS.n3019 0.8195
R5245 VSS.n2715 VSS.n2709 0.799363
R5246 VSS.n1290 VSS.n1247 0.799163
R5247 VSS.n1107 VSS.n1064 0.799163
R5248 VSS.n924 VSS.n898 0.799163
R5249 VSS.n2302 VSS.n2299 0.798761
R5250 VSS.n2306 VSS.n2305 0.798761
R5251 VSS.n2307 VSS.n2306 0.798761
R5252 VSS.n2303 VSS.n2302 0.798761
R5253 VSS.n3544 VSS.n3543 0.798761
R5254 VSS.n3480 VSS.n3479 0.798761
R5255 VSS.n3485 VSS.n3484 0.798761
R5256 VSS.n3486 VSS.n3485 0.798761
R5257 VSS.n3479 VSS.n3478 0.798761
R5258 VSS.n3538 VSS.n3535 0.798761
R5259 VSS.n3539 VSS.n3538 0.798761
R5260 VSS.n3545 VSS.n3544 0.798761
R5261 VSS.n2311 VSS.n2310 0.798761
R5262 VSS.n2432 VSS.n2429 0.798761
R5263 VSS.n2433 VSS.n2432 0.798761
R5264 VSS.n2310 VSS.n2309 0.798761
R5265 VSS.n3938 VSS.n3839 0.775283
R5266 VSS.n3949 VSS.n3948 0.775283
R5267 VSS.n2608 VSS.n2566 0.775283
R5268 VSS.n2601 VSS.n2568 0.775283
R5269 VSS.n4104 VSS.t340 0.767281
R5270 VSS.n3740 VSS.t314 0.767281
R5271 VSS.n3824 VSS.n3780 0.738109
R5272 VSS.n3817 VSS.n3786 0.738109
R5273 VSS.n2511 VSS.n2479 0.738109
R5274 VSS.n2518 VSS.n2473 0.738109
R5275 VSS.n2706 VSS.n2705 0.68137
R5276 VSS.n2704 VSS.n2701 0.68137
R5277 VSS.n2684 VSS.n2683 0.68137
R5278 VSS.n2682 VSS.n2681 0.68137
R5279 VSS.n949 VSS.t320 0.656602
R5280 VSS.n1005 VSS.t290 0.656602
R5281 VSS.n1132 VSS.t293 0.656602
R5282 VSS.n1188 VSS.t305 0.656602
R5283 VSS.n1315 VSS.t299 0.656602
R5284 VSS.n1371 VSS.t302 0.656602
R5285 VSS.n2023 VSS.n2022 0.640666
R5286 VSS.n1768 VSS.n1767 0.626587
R5287 VSS.n1767 VSS.n1766 0.626587
R5288 VSS.n1637 VSS.n1636 0.626587
R5289 VSS.n1638 VSS.n1637 0.626587
R5290 VSS.n1508 VSS.n1507 0.626587
R5291 VSS.n1507 VSS.n1506 0.626587
R5292 VSS.n2554 VSS.n2553 0.626587
R5293 VSS.n2553 VSS.n2552 0.626587
R5294 VSS.n2552 VSS.n2551 0.626587
R5295 VSS.n2551 VSS.n2550 0.626587
R5296 VSS.n2550 VSS.n2549 0.626587
R5297 VSS.n3131 VSS.n3128 0.624916
R5298 VSS.n3727 VSS.n3726 0.624916
R5299 VSS.n3326 VSS.n3324 0.624916
R5300 VSS.n2590 VSS.n2589 0.624916
R5301 VSS.n3929 VSS.n3928 0.624916
R5302 VSS.n3378 VSS.n3377 0.624916
R5303 VSS.n2415 VSS.n2414 0.624916
R5304 VSS.n2414 VSS.n2413 0.624916
R5305 VSS.n1290 VSS.n1245 0.624916
R5306 VSS.n1947 VSS.n1946 0.624916
R5307 VSS.n1107 VSS.n1062 0.624916
R5308 VSS.n1869 VSS.n1868 0.624916
R5309 VSS.n1291 VSS.n1290 0.624916
R5310 VSS.n1108 VSS.n1107 0.624916
R5311 VSS.n925 VSS.n924 0.624916
R5312 VSS.n1238 VSS.n1237 0.624916
R5313 VSS.n1055 VSS.n1054 0.624916
R5314 VSS.n4054 VSS.n4053 0.62468
R5315 VSS.n4055 VSS.n4054 0.62468
R5316 VSS.n3470 VSS.n3445 0.62468
R5317 VSS.n3471 VSS.n3470 0.62468
R5318 VSS.n3470 VSS.n3469 0.62468
R5319 VSS.n2953 VSS.n2866 0.608978
R5320 VSS.n3879 VSS.n3841 0.608978
R5321 VSS.n3884 VSS.n3840 0.608978
R5322 VSS.n2948 VSS.n2947 0.608978
R5323 VSS.n1950 VSS.n1947 0.6035
R5324 VSS.n3839 VSS.n3838 0.57963
R5325 VSS.n3948 VSS.n3947 0.57963
R5326 VSS.n2568 VSS.n2567 0.57963
R5327 VSS.n3767 VSS.t268 0.56925
R5328 VSS.n3767 VSS.n3766 0.56925
R5329 VSS.n3764 VSS.t215 0.56925
R5330 VSS.n3764 VSS.n3763 0.56925
R5331 VSS.n3761 VSS.t505 0.56925
R5332 VSS.n3761 VSS.n3760 0.56925
R5333 VSS.n3758 VSS.t492 0.56925
R5334 VSS.n3758 VSS.n3757 0.56925
R5335 VSS.n3755 VSS.t205 0.56925
R5336 VSS.n3755 VSS.n3754 0.56925
R5337 VSS.n283 VSS.t239 0.56925
R5338 VSS.n283 VSS.n282 0.56925
R5339 VSS.n281 VSS.t270 0.56925
R5340 VSS.n281 VSS.n280 0.56925
R5341 VSS.n279 VSS.t208 0.56925
R5342 VSS.n279 VSS.n278 0.56925
R5343 VSS.n3530 VSS.t237 0.56925
R5344 VSS.n3530 VSS.n3529 0.56925
R5345 VSS.n3527 VSS.t513 0.56925
R5346 VSS.n3527 VSS.n3526 0.56925
R5347 VSS.n3524 VSS.t610 0.56925
R5348 VSS.n3524 VSS.n3523 0.56925
R5349 VSS.n3521 VSS.t236 0.56925
R5350 VSS.n3521 VSS.n3520 0.56925
R5351 VSS.n3518 VSS.t510 0.56925
R5352 VSS.n3518 VSS.n3517 0.56925
R5353 VSS.n274 VSS.t496 0.56925
R5354 VSS.n274 VSS.n273 0.56925
R5355 VSS.n272 VSS.t207 0.56925
R5356 VSS.n272 VSS.n271 0.56925
R5357 VSS.n270 VSS.t550 0.56925
R5358 VSS.n270 VSS.n269 0.56925
R5359 VSS.n3515 VSS.t200 0.56925
R5360 VSS.n3515 VSS.n3514 0.56925
R5361 VSS.n3512 VSS.t11 0.56925
R5362 VSS.n3512 VSS.n3511 0.56925
R5363 VSS.n3509 VSS.t46 0.56925
R5364 VSS.n3509 VSS.n3508 0.56925
R5365 VSS.n3506 VSS.t556 0.56925
R5366 VSS.n3506 VSS.n3505 0.56925
R5367 VSS.n3503 VSS.t214 0.56925
R5368 VSS.n3503 VSS.n3502 0.56925
R5369 VSS.n265 VSS.t4 0.56925
R5370 VSS.n265 VSS.n264 0.56925
R5371 VSS.n263 VSS.t613 0.56925
R5372 VSS.n263 VSS.n262 0.56925
R5373 VSS.n261 VSS.t216 0.56925
R5374 VSS.n261 VSS.n260 0.56925
R5375 VSS.n3500 VSS.t229 0.56925
R5376 VSS.n3500 VSS.n3499 0.56925
R5377 VSS.n3497 VSS.t493 0.56925
R5378 VSS.n3497 VSS.n3496 0.56925
R5379 VSS.n3494 VSS.t269 0.56925
R5380 VSS.n3494 VSS.n3493 0.56925
R5381 VSS.n3491 VSS.t491 0.56925
R5382 VSS.n3491 VSS.n3490 0.56925
R5383 VSS.n3488 VSS.t57 0.56925
R5384 VSS.n3488 VSS.n3487 0.56925
R5385 VSS.n256 VSS.t238 0.56925
R5386 VSS.n256 VSS.n255 0.56925
R5387 VSS.n254 VSS.t551 0.56925
R5388 VSS.n254 VSS.n253 0.56925
R5389 VSS.n252 VSS.t201 0.56925
R5390 VSS.n252 VSS.n251 0.56925
R5391 VSS.n2555 VSS.n2554 0.563978
R5392 VSS.n3331 VSS.n3326 0.556813
R5393 VSS.n1698 VSS.t635 0.5465
R5394 VSS.n1698 VSS.n1697 0.5465
R5395 VSS.n1690 VSS.t119 0.5465
R5396 VSS.n1690 VSS.n1689 0.5465
R5397 VSS.n1693 VSS.t187 0.5465
R5398 VSS.n1693 VSS.n1692 0.5465
R5399 VSS.n1686 VSS.t598 0.5465
R5400 VSS.n1686 VSS.n1685 0.5465
R5401 VSS.n1684 VSS.t107 0.5465
R5402 VSS.n1684 VSS.n1683 0.5465
R5403 VSS.n1701 VSS.t99 0.5465
R5404 VSS.n1701 VSS.n1700 0.5465
R5405 VSS.n1718 VSS.t112 0.5465
R5406 VSS.n1718 VSS.n1717 0.5465
R5407 VSS.n1710 VSS.t589 0.5465
R5408 VSS.n1710 VSS.n1709 0.5465
R5409 VSS.n1713 VSS.t604 0.5465
R5410 VSS.n1713 VSS.n1712 0.5465
R5411 VSS.n1706 VSS.t88 0.5465
R5412 VSS.n1706 VSS.n1705 0.5465
R5413 VSS.n1704 VSS.t593 0.5465
R5414 VSS.n1704 VSS.n1703 0.5465
R5415 VSS.n1721 VSS.t573 0.5465
R5416 VSS.n1721 VSS.n1720 0.5465
R5417 VSS.n1754 VSS.t576 0.5465
R5418 VSS.n1754 VSS.n1753 0.5465
R5419 VSS.n1757 VSS.t162 0.5465
R5420 VSS.n1757 VSS.n1756 0.5465
R5421 VSS.n1739 VSS.t79 0.5465
R5422 VSS.n1739 VSS.n1738 0.5465
R5423 VSS.n1742 VSS.t111 0.5465
R5424 VSS.n1742 VSS.n1741 0.5465
R5425 VSS.n1746 VSS.t581 0.5465
R5426 VSS.n1746 VSS.n1745 0.5465
R5427 VSS.n1744 VSS.t668 0.5465
R5428 VSS.n1744 VSS.n1743 0.5465
R5429 VSS.n1730 VSS.t655 0.5465
R5430 VSS.n1730 VSS.n1729 0.5465
R5431 VSS.n1733 VSS.t150 0.5465
R5432 VSS.n1733 VSS.n1732 0.5465
R5433 VSS.n1724 VSS.t195 0.5465
R5434 VSS.n1724 VSS.n1723 0.5465
R5435 VSS.n1726 VSS.t676 0.5465
R5436 VSS.n1726 VSS.n1725 0.5465
R5437 VSS.n1762 VSS.t166 0.5465
R5438 VSS.n1762 VSS.n1761 0.5465
R5439 VSS.n1765 VSS.t662 0.5465
R5440 VSS.n1765 VSS.n1764 0.5465
R5441 VSS.n1568 VSS.t130 0.5465
R5442 VSS.n1568 VSS.n1567 0.5465
R5443 VSS.n1560 VSS.t675 0.5465
R5444 VSS.n1560 VSS.n1559 0.5465
R5445 VSS.n1563 VSS.t592 0.5465
R5446 VSS.n1563 VSS.n1562 0.5465
R5447 VSS.n1556 VSS.t143 0.5465
R5448 VSS.n1556 VSS.n1555 0.5465
R5449 VSS.n1554 VSS.t680 0.5465
R5450 VSS.n1554 VSS.n1553 0.5465
R5451 VSS.n1571 VSS.t683 0.5465
R5452 VSS.n1571 VSS.n1570 0.5465
R5453 VSS.n1635 VSS.t71 0.5465
R5454 VSS.n1635 VSS.n1634 0.5465
R5455 VSS.n1624 VSS.t196 0.5465
R5456 VSS.n1624 VSS.n1623 0.5465
R5457 VSS.n1627 VSS.t663 0.5465
R5458 VSS.n1627 VSS.n1626 0.5465
R5459 VSS.n1609 VSS.t636 0.5465
R5460 VSS.n1609 VSS.n1608 0.5465
R5461 VSS.n1612 VSS.t666 0.5465
R5462 VSS.n1612 VSS.n1611 0.5465
R5463 VSS.n1616 VSS.t161 0.5465
R5464 VSS.n1616 VSS.n1615 0.5465
R5465 VSS.n1614 VSS.t110 0.5465
R5466 VSS.n1614 VSS.n1613 0.5465
R5467 VSS.n1600 VSS.t186 0.5465
R5468 VSS.n1600 VSS.n1599 0.5465
R5469 VSS.n1603 VSS.t605 0.5465
R5470 VSS.n1603 VSS.n1602 0.5465
R5471 VSS.n1594 VSS.t641 0.5465
R5472 VSS.n1594 VSS.n1593 0.5465
R5473 VSS.n1596 VSS.t97 0.5465
R5474 VSS.n1596 VSS.n1595 0.5465
R5475 VSS.n1632 VSS.t597 0.5465
R5476 VSS.n1632 VSS.n1631 0.5465
R5477 VSS.n1588 VSS.t699 0.5465
R5478 VSS.n1588 VSS.n1587 0.5465
R5479 VSS.n1580 VSS.t163 0.5465
R5480 VSS.n1580 VSS.n1579 0.5465
R5481 VSS.n1583 VSS.t114 0.5465
R5482 VSS.n1583 VSS.n1582 0.5465
R5483 VSS.n1576 VSS.t579 0.5465
R5484 VSS.n1576 VSS.n1575 0.5465
R5485 VSS.n1574 VSS.t148 0.5465
R5486 VSS.n1574 VSS.n1573 0.5465
R5487 VSS.n1591 VSS.t172 0.5465
R5488 VSS.n1591 VSS.n1590 0.5465
R5489 VSS.n1438 VSS.t652 0.5465
R5490 VSS.n1438 VSS.n1437 0.5465
R5491 VSS.n1430 VSS.t153 0.5465
R5492 VSS.n1430 VSS.n1429 0.5465
R5493 VSS.n1433 VSS.t171 0.5465
R5494 VSS.n1433 VSS.n1432 0.5465
R5495 VSS.n1426 VSS.t588 0.5465
R5496 VSS.n1426 VSS.n1425 0.5465
R5497 VSS.n1424 VSS.t139 0.5465
R5498 VSS.n1424 VSS.n1423 0.5465
R5499 VSS.n1441 VSS.t81 0.5465
R5500 VSS.n1441 VSS.n1440 0.5465
R5501 VSS.n1458 VSS.t109 0.5465
R5502 VSS.n1458 VSS.n1457 0.5465
R5503 VSS.n1450 VSS.t679 0.5465
R5504 VSS.n1450 VSS.n1449 0.5465
R5505 VSS.n1453 VSS.t629 0.5465
R5506 VSS.n1453 VSS.n1452 0.5465
R5507 VSS.n1446 VSS.t135 0.5465
R5508 VSS.n1446 VSS.n1445 0.5465
R5509 VSS.n1444 VSS.t686 0.5465
R5510 VSS.n1444 VSS.n1443 0.5465
R5511 VSS.n1461 VSS.t580 0.5465
R5512 VSS.n1461 VSS.n1460 0.5465
R5513 VSS.n1494 VSS.t582 0.5465
R5514 VSS.n1494 VSS.n1493 0.5465
R5515 VSS.n1497 VSS.t157 0.5465
R5516 VSS.n1497 VSS.n1496 0.5465
R5517 VSS.n1479 VSS.t128 0.5465
R5518 VSS.n1479 VSS.n1478 0.5465
R5519 VSS.n1482 VSS.t104 0.5465
R5520 VSS.n1482 VSS.n1481 0.5465
R5521 VSS.n1486 VSS.t585 0.5465
R5522 VSS.n1486 VSS.n1485 0.5465
R5523 VSS.n1484 VSS.t601 0.5465
R5524 VSS.n1484 VSS.n1483 0.5465
R5525 VSS.n1470 VSS.t596 0.5465
R5526 VSS.n1470 VSS.n1469 0.5465
R5527 VSS.n1473 VSS.t194 0.5465
R5528 VSS.n1473 VSS.n1472 0.5465
R5529 VSS.n1464 VSS.t115 0.5465
R5530 VSS.n1464 VSS.n1463 0.5465
R5531 VSS.n1466 VSS.t632 0.5465
R5532 VSS.n1466 VSS.n1465 0.5465
R5533 VSS.n1502 VSS.t158 0.5465
R5534 VSS.n1502 VSS.n1501 0.5465
R5535 VSS.n1505 VSS.t667 0.5465
R5536 VSS.n1505 VSS.n1504 0.5465
R5537 VSS.n1819 VSS.n1768 0.5405
R5538 VSS.n1919 VSS.n1638 0.5405
R5539 VSS.n1975 VSS.n1508 0.5405
R5540 VSS.n3782 VSS.n3781 0.479848
R5541 VSS.n3777 VSS.n3776 0.479848
R5542 VSS.n3776 VSS.n3773 0.479848
R5543 VSS.n3783 VSS.n3782 0.479848
R5544 VSS.n2469 VSS.n2466 0.479848
R5545 VSS.n2476 VSS.n2475 0.479848
R5546 VSS.n2475 VSS.n2474 0.479848
R5547 VSS.n2470 VSS.n2469 0.479848
R5548 VSS.n1290 VSS.n1246 0.472687
R5549 VSS.n1237 VSS.n1236 0.472687
R5550 VSS.n1237 VSS.n1235 0.472687
R5551 VSS.n1237 VSS.n1234 0.472687
R5552 VSS.n1237 VSS.n1233 0.472687
R5553 VSS.n1237 VSS.n1232 0.472687
R5554 VSS.n1237 VSS.n1231 0.472687
R5555 VSS.n1237 VSS.n1230 0.472687
R5556 VSS.n1237 VSS.n1229 0.472687
R5557 VSS.n1237 VSS.n1228 0.472687
R5558 VSS.n1237 VSS.n1227 0.472687
R5559 VSS.n1237 VSS.n1226 0.472687
R5560 VSS.n1237 VSS.n1225 0.472687
R5561 VSS.n1237 VSS.n1224 0.472687
R5562 VSS.n1237 VSS.n1223 0.472687
R5563 VSS.n1237 VSS.n1222 0.472687
R5564 VSS.n1237 VSS.n1221 0.472687
R5565 VSS.n1237 VSS.n1220 0.472687
R5566 VSS.n1237 VSS.n1219 0.472687
R5567 VSS.n1237 VSS.n1218 0.472687
R5568 VSS.n1237 VSS.n1217 0.472687
R5569 VSS.n1237 VSS.n1216 0.472687
R5570 VSS.n1237 VSS.n1215 0.472687
R5571 VSS.n1237 VSS.n1214 0.472687
R5572 VSS.n1237 VSS.n1213 0.472687
R5573 VSS.n1237 VSS.n1212 0.472687
R5574 VSS.n1237 VSS.n1211 0.472687
R5575 VSS.n1107 VSS.n1063 0.472687
R5576 VSS.n1054 VSS.n1053 0.472687
R5577 VSS.n1054 VSS.n1052 0.472687
R5578 VSS.n1054 VSS.n1051 0.472687
R5579 VSS.n1054 VSS.n1050 0.472687
R5580 VSS.n1054 VSS.n1049 0.472687
R5581 VSS.n1054 VSS.n1048 0.472687
R5582 VSS.n1054 VSS.n1047 0.472687
R5583 VSS.n1054 VSS.n1046 0.472687
R5584 VSS.n1054 VSS.n1045 0.472687
R5585 VSS.n1054 VSS.n1044 0.472687
R5586 VSS.n1054 VSS.n1043 0.472687
R5587 VSS.n1054 VSS.n1042 0.472687
R5588 VSS.n1054 VSS.n1041 0.472687
R5589 VSS.n1054 VSS.n1040 0.472687
R5590 VSS.n1054 VSS.n1039 0.472687
R5591 VSS.n1054 VSS.n1038 0.472687
R5592 VSS.n1054 VSS.n1037 0.472687
R5593 VSS.n1054 VSS.n1036 0.472687
R5594 VSS.n1054 VSS.n1035 0.472687
R5595 VSS.n1054 VSS.n1034 0.472687
R5596 VSS.n1054 VSS.n1033 0.472687
R5597 VSS.n1054 VSS.n1032 0.472687
R5598 VSS.n1054 VSS.n1031 0.472687
R5599 VSS.n1054 VSS.n1030 0.472687
R5600 VSS.n1054 VSS.n1029 0.472687
R5601 VSS.n1054 VSS.n1028 0.472687
R5602 VSS.n924 VSS.n923 0.472687
R5603 VSS.n924 VSS.n922 0.472687
R5604 VSS.n924 VSS.n921 0.472687
R5605 VSS.n924 VSS.n920 0.472687
R5606 VSS.n924 VSS.n919 0.472687
R5607 VSS.n924 VSS.n918 0.472687
R5608 VSS.n924 VSS.n917 0.472687
R5609 VSS.n924 VSS.n916 0.472687
R5610 VSS.n924 VSS.n915 0.472687
R5611 VSS.n924 VSS.n914 0.472687
R5612 VSS.n924 VSS.n913 0.472687
R5613 VSS.n924 VSS.n912 0.472687
R5614 VSS.n924 VSS.n911 0.472687
R5615 VSS.n924 VSS.n910 0.472687
R5616 VSS.n924 VSS.n909 0.472687
R5617 VSS.n924 VSS.n908 0.472687
R5618 VSS.n924 VSS.n907 0.472687
R5619 VSS.n924 VSS.n906 0.472687
R5620 VSS.n924 VSS.n905 0.472687
R5621 VSS.n924 VSS.n904 0.472687
R5622 VSS.n924 VSS.n903 0.472687
R5623 VSS.n924 VSS.n902 0.472687
R5624 VSS.n924 VSS.n901 0.472687
R5625 VSS.n924 VSS.n900 0.472687
R5626 VSS.n924 VSS.n899 0.472687
R5627 VSS.n2713 VSS.n2712 0.472687
R5628 VSS.n3127 VSS.n3126 0.472687
R5629 VSS.n3727 VSS.n3720 0.472687
R5630 VSS.n3727 VSS.n3717 0.472687
R5631 VSS.n3727 VSS.n3714 0.472687
R5632 VSS.n3727 VSS.n3711 0.472687
R5633 VSS.n3727 VSS.n3708 0.472687
R5634 VSS.n3727 VSS.n3705 0.472687
R5635 VSS.n3727 VSS.n3702 0.472687
R5636 VSS.n3727 VSS.n3699 0.472687
R5637 VSS.n3727 VSS.n3696 0.472687
R5638 VSS.n3727 VSS.n3693 0.472687
R5639 VSS.n3727 VSS.n3692 0.472687
R5640 VSS.n3727 VSS.n3691 0.472687
R5641 VSS.n3727 VSS.n3690 0.472687
R5642 VSS.n3727 VSS.n3689 0.472687
R5643 VSS.n3727 VSS.n3688 0.472687
R5644 VSS.n3727 VSS.n3687 0.472687
R5645 VSS.n3727 VSS.n3686 0.472687
R5646 VSS.n3727 VSS.n3685 0.472687
R5647 VSS.n3727 VSS.n3684 0.472687
R5648 VSS.n3727 VSS.n3683 0.472687
R5649 VSS.n3727 VSS.n3682 0.472687
R5650 VSS.n3727 VSS.n3681 0.472687
R5651 VSS.n3727 VSS.n3680 0.472687
R5652 VSS.n3727 VSS.n3679 0.472687
R5653 VSS.n3727 VSS.n3678 0.472687
R5654 VSS.n3727 VSS.n3677 0.472687
R5655 VSS.n3727 VSS.n3676 0.472687
R5656 VSS.n3727 VSS.n3675 0.472687
R5657 VSS.n3727 VSS.n3674 0.472687
R5658 VSS.n3728 VSS.n3727 0.472687
R5659 VSS.n2414 VSS.n2412 0.472687
R5660 VSS.n2414 VSS.n2411 0.472687
R5661 VSS.n2414 VSS.n2410 0.472687
R5662 VSS.n2414 VSS.n2409 0.472687
R5663 VSS.n2414 VSS.n2408 0.472687
R5664 VSS.n2414 VSS.n2407 0.472687
R5665 VSS.n2414 VSS.n2406 0.472687
R5666 VSS.n2414 VSS.n2405 0.472687
R5667 VSS.n2414 VSS.n2404 0.472687
R5668 VSS.n2414 VSS.n2403 0.472687
R5669 VSS.n2414 VSS.n2402 0.472687
R5670 VSS.n2414 VSS.n2401 0.472687
R5671 VSS.n2414 VSS.n2400 0.472687
R5672 VSS.n2414 VSS.n2399 0.472687
R5673 VSS.n3727 VSS.n3723 0.472687
R5674 VSS.n3323 VSS.n3322 0.472687
R5675 VSS.n2594 VSS.n2592 0.472687
R5676 VSS.n2674 VSS.n2670 0.472687
R5677 VSS.n3322 VSS.n3321 0.472687
R5678 VSS.n3322 VSS.n3320 0.472687
R5679 VSS.n3322 VSS.n3319 0.472687
R5680 VSS.n3322 VSS.n3318 0.472687
R5681 VSS.n2960 VSS.n2855 0.472687
R5682 VSS.n2668 VSS.n2665 0.472687
R5683 VSS.n2674 VSS.n2673 0.472687
R5684 VSS.n2589 VSS.n2588 0.472687
R5685 VSS.n2958 VSS.n2864 0.472687
R5686 VSS.n3331 VSS.n3329 0.472687
R5687 VSS.n2642 VSS.n2640 0.472687
R5688 VSS.n2169 VSS.n2167 0.472687
R5689 VSS.n2166 VSS.n2165 0.472687
R5690 VSS.n2176 VSS.n2174 0.472687
R5691 VSS.n2165 VSS.n2164 0.472687
R5692 VSS.n2165 VSS.n2163 0.472687
R5693 VSS.n2165 VSS.n2162 0.472687
R5694 VSS.n2165 VSS.n2161 0.472687
R5695 VSS.n2165 VSS.n2160 0.472687
R5696 VSS.n2165 VSS.n2159 0.472687
R5697 VSS.n2165 VSS.n2158 0.472687
R5698 VSS.n2165 VSS.n2157 0.472687
R5699 VSS.n2165 VSS.n2156 0.472687
R5700 VSS.n2165 VSS.n2155 0.472687
R5701 VSS.n2165 VSS.n2154 0.472687
R5702 VSS.n2165 VSS.n2153 0.472687
R5703 VSS.n2165 VSS.n2152 0.472687
R5704 VSS.n2165 VSS.n2151 0.472687
R5705 VSS.n2165 VSS.n2150 0.472687
R5706 VSS.n2165 VSS.n2149 0.472687
R5707 VSS.n2165 VSS.n2148 0.472687
R5708 VSS.n2165 VSS.n2147 0.472687
R5709 VSS.n2165 VSS.n2146 0.472687
R5710 VSS.n234 VSS.n232 0.472687
R5711 VSS.n1397 VSS.n1395 0.472687
R5712 VSS.n1294 VSS.n1292 0.472687
R5713 VSS.n1242 VSS.n1240 0.472687
R5714 VSS.n1111 VSS.n1109 0.472687
R5715 VSS.n1059 VSS.n1057 0.472687
R5716 VSS.n928 VSS.n926 0.472687
R5717 VSS.n4054 VSS.n4052 0.472445
R5718 VSS.n4054 VSS.n4051 0.472445
R5719 VSS.n4054 VSS.n4050 0.472445
R5720 VSS.n4054 VSS.n4049 0.472445
R5721 VSS.n4054 VSS.n4048 0.472445
R5722 VSS.n4054 VSS.n4047 0.472445
R5723 VSS.n4054 VSS.n4046 0.472445
R5724 VSS.n4054 VSS.n4045 0.472445
R5725 VSS.n3470 VSS.n3444 0.472445
R5726 VSS.n3470 VSS.n3443 0.472445
R5727 VSS.n3470 VSS.n3442 0.472445
R5728 VSS.n3470 VSS.n3441 0.472445
R5729 VSS.n3470 VSS.n3440 0.472445
R5730 VSS.n3470 VSS.n3439 0.472445
R5731 VSS.n3470 VSS.n3438 0.472445
R5732 VSS.n3470 VSS.n3437 0.472445
R5733 VSS.n3470 VSS.n3436 0.472445
R5734 VSS.n3470 VSS.n3435 0.472445
R5735 VSS.n3470 VSS.n3434 0.472445
R5736 VSS.n3470 VSS.n3433 0.472445
R5737 VSS.n3470 VSS.n3432 0.472445
R5738 VSS.n3470 VSS.n3431 0.472445
R5739 VSS.n358 VSS.n244 0.472445
R5740 VSS.n3470 VSS.n3461 0.472445
R5741 VSS.n3470 VSS.n3467 0.472445
R5742 VSS.n3470 VSS.n3464 0.472445
R5743 VSS.n3470 VSS.n3457 0.472445
R5744 VSS.n3470 VSS.n3456 0.472445
R5745 VSS.n3470 VSS.n3458 0.472445
R5746 VSS.n3470 VSS.n3446 0.472445
R5747 VSS.n3470 VSS.n3453 0.472445
R5748 VSS.n3470 VSS.n3451 0.472445
R5749 VSS.n3470 VSS.n3450 0.472445
R5750 VSS.n3470 VSS.n3449 0.472445
R5751 VSS.n3470 VSS.n3448 0.472445
R5752 VSS.n3470 VSS.n3447 0.472445
R5753 VSS.n3470 VSS.n3454 0.472445
R5754 VSS.n3470 VSS.n3455 0.472445
R5755 VSS.n3470 VSS.n3459 0.472445
R5756 VSS.n3470 VSS.n3452 0.459997
R5757 VSS.n3727 VSS.n3694 0.457229
R5758 VSS.n2528 VSS.t473 0.426562
R5759 VSS.n3787 VSS.t242 0.426562
R5760 VSS.t265 VSS.t311 0.426562
R5761 VSS.n1243 VSS.n1242 0.320562
R5762 VSS.n1294 VSS.n1243 0.283437
R5763 VSS.n2566 VSS.n2565 0.282239
R5764 VSS.n1872 VSS.n1869 0.270781
R5765 VSS.n2960 VSS.n2958 0.266
R5766 VSS.n362 VSS.n361 0.229438
R5767 VSS.n2171 VSS.n2170 0.229438
R5768 VSS.n230 VSS.n229 0.229438
R5769 VSS.n2565 VSS.n2564 0.207891
R5770 VSS.n361 VSS.n360 0.198781
R5771 VSS.n2172 VSS.n2171 0.198781
R5772 VSS.n231 VSS.n230 0.198781
R5773 VSS.n1768 VSS.n1702 0.190381
R5774 VSS.n1767 VSS.n1722 0.190381
R5775 VSS.n1766 VSS.n1763 0.190381
R5776 VSS.n1638 VSS.n1572 0.190381
R5777 VSS.n1636 VSS.n1633 0.190381
R5778 VSS.n1637 VSS.n1592 0.190381
R5779 VSS.n1508 VSS.n1442 0.190381
R5780 VSS.n1507 VSS.n1462 0.190381
R5781 VSS.n1506 VSS.n1503 0.190381
R5782 VSS.n360 VSS.n359 0.188375
R5783 VSS.n2177 VSS.n2172 0.188375
R5784 VSS.n235 VSS.n231 0.188375
R5785 VSS.n761 VSS.n760 0.157022
R5786 VSS.n1677 VSS.n1676 0.157022
R5787 VSS.n498 VSS.n497 0.157022
R5788 VSS.n1643 VSS.n1642 0.157022
R5789 VSS.n488 VSS.n487 0.157022
R5790 VSS.n1547 VSS.n1546 0.157022
R5791 VSS.n83 VSS.n82 0.157022
R5792 VSS.n1513 VSS.n1512 0.157022
R5793 VSS.n73 VSS.n72 0.157022
R5794 VSS.n1417 VSS.n1416 0.157022
R5795 VSS.n2302 VSS.n2301 0.157022
R5796 VSS.n3947 VSS.n3946 0.157022
R5797 VSS.n2564 VSS.n2563 0.157022
R5798 VSS.n3776 VSS.n3775 0.157022
R5799 VSS.n2469 VSS.n2468 0.157022
R5800 VSS.n3479 VSS.n3474 0.157022
R5801 VSS.n3538 VSS.n3537 0.157022
R5802 VSS.n2432 VSS.n2431 0.157022
R5803 VSS.n1773 VSS.n1770 0.157022
R5804 VSS.n771 VSS.n770 0.157022
R5805 VSS.n1060 VSS.n636 0.148156
R5806 VSS.n1243 VSS.n363 0.148156
R5807 VSS.n1111 VSS.n1060 0.138594
R5808 VSS.n1060 VSS.n1059 0.132688
R5809 VSS.n1696 VSS.n1688 0.123658
R5810 VSS.n1716 VSS.n1708 0.123658
R5811 VSS.n1736 VSS.n1728 0.123658
R5812 VSS.n1751 VSS.n1737 0.123658
R5813 VSS.n1760 VSS.n1752 0.123658
R5814 VSS.n1566 VSS.n1558 0.123658
R5815 VSS.n1606 VSS.n1598 0.123658
R5816 VSS.n1621 VSS.n1607 0.123658
R5817 VSS.n1630 VSS.n1622 0.123658
R5818 VSS.n1586 VSS.n1578 0.123658
R5819 VSS.n1436 VSS.n1428 0.123658
R5820 VSS.n1456 VSS.n1448 0.123658
R5821 VSS.n1476 VSS.n1468 0.123658
R5822 VSS.n1491 VSS.n1477 0.123658
R5823 VSS.n1500 VSS.n1492 0.123658
R5824 VSS.n1695 VSS.n1691 0.109963
R5825 VSS.n1715 VSS.n1711 0.109963
R5826 VSS.n1759 VSS.n1755 0.109963
R5827 VSS.n1750 VSS.n1740 0.109963
R5828 VSS.n1735 VSS.n1731 0.109963
R5829 VSS.n1565 VSS.n1561 0.109963
R5830 VSS.n1629 VSS.n1625 0.109963
R5831 VSS.n1620 VSS.n1610 0.109963
R5832 VSS.n1605 VSS.n1601 0.109963
R5833 VSS.n1585 VSS.n1581 0.109963
R5834 VSS.n1435 VSS.n1431 0.109963
R5835 VSS.n1455 VSS.n1451 0.109963
R5836 VSS.n1499 VSS.n1495 0.109963
R5837 VSS.n1490 VSS.n1480 0.109963
R5838 VSS.n1475 VSS.n1471 0.109963
R5839 VSS.n3561 VSS.n3559 0.0800536
R5840 VSS.n3563 VSS.n3561 0.07925
R5841 VSS.n2317 VSS.n2315 0.0760357
R5842 VSS.n2319 VSS.n2317 0.0760357
R5843 VSS.n2321 VSS.n2319 0.0760357
R5844 VSS.n2323 VSS.n2321 0.0760357
R5845 VSS.n2325 VSS.n2323 0.0760357
R5846 VSS.n2327 VSS.n2325 0.0760357
R5847 VSS.n2329 VSS.n2327 0.0760357
R5848 VSS.n2331 VSS.n2329 0.0760357
R5849 VSS.n2333 VSS.n2331 0.0760357
R5850 VSS.n2335 VSS.n2333 0.0760357
R5851 VSS.n2337 VSS.n2335 0.0760357
R5852 VSS.n2339 VSS.n2337 0.0760357
R5853 VSS.n2341 VSS.n2339 0.0760357
R5854 VSS.n2343 VSS.n2341 0.0760357
R5855 VSS.n2345 VSS.n2343 0.0760357
R5856 VSS.n2347 VSS.n2345 0.0760357
R5857 VSS.n2349 VSS.n2347 0.0760357
R5858 VSS.n2351 VSS.n2349 0.0760357
R5859 VSS.n2353 VSS.n2351 0.0760357
R5860 VSS.n2355 VSS.n2353 0.0760357
R5861 VSS.n2357 VSS.n2355 0.0760357
R5862 VSS.n2359 VSS.n2357 0.0760357
R5863 VSS.n2361 VSS.n2359 0.0760357
R5864 VSS.n2363 VSS.n2361 0.0760357
R5865 VSS.n2365 VSS.n2363 0.0760357
R5866 VSS.n2367 VSS.n2365 0.0760357
R5867 VSS.n2369 VSS.n2367 0.0760357
R5868 VSS.n2371 VSS.n2369 0.0760357
R5869 VSS.n2373 VSS.n2371 0.0760357
R5870 VSS.n2376 VSS.n2373 0.0760357
R5871 VSS.n2378 VSS.n2376 0.0760357
R5872 VSS.n2381 VSS.n2378 0.0760357
R5873 VSS.n2383 VSS.n2381 0.0760357
R5874 VSS.n2386 VSS.n2383 0.0760357
R5875 VSS.n2388 VSS.n2386 0.0760357
R5876 VSS.n2391 VSS.n2388 0.0760357
R5877 VSS.n2393 VSS.n2391 0.0760357
R5878 VSS.n2396 VSS.n2393 0.0760357
R5879 VSS.n2398 VSS.n2396 0.0760357
R5880 VSS.n299 VSS.n298 0.0760357
R5881 VSS.n298 VSS.n297 0.0760357
R5882 VSS.n297 VSS.n296 0.0760357
R5883 VSS.n296 VSS.n295 0.0760357
R5884 VSS.n295 VSS.n294 0.0760357
R5885 VSS.n294 VSS.n293 0.0760357
R5886 VSS.n293 VSS.n292 0.0760357
R5887 VSS.n292 VSS.n291 0.0760357
R5888 VSS.n291 VSS.n290 0.0760357
R5889 VSS.n3547 VSS.n3546 0.0760357
R5890 VSS.n3548 VSS.n3547 0.0760357
R5891 VSS.n3549 VSS.n3548 0.0760357
R5892 VSS.n3550 VSS.n3549 0.0760357
R5893 VSS.n3551 VSS.n3550 0.0760357
R5894 VSS.n3552 VSS.n3551 0.0760357
R5895 VSS.n3553 VSS.n3552 0.0760357
R5896 VSS.n3554 VSS.n3553 0.0760357
R5897 VSS.n3555 VSS.n3554 0.0760357
R5898 VSS.n3557 VSS.n3555 0.0760357
R5899 VSS.n3559 VSS.n3557 0.0760357
R5900 VSS.n3565 VSS.n3563 0.0760357
R5901 VSS.n3567 VSS.n3565 0.0760357
R5902 VSS.n3569 VSS.n3567 0.0760357
R5903 VSS.n3571 VSS.n3569 0.0760357
R5904 VSS.n3573 VSS.n3571 0.0760357
R5905 VSS.n3575 VSS.n3573 0.0760357
R5906 VSS.n3577 VSS.n3575 0.0760357
R5907 VSS.n3579 VSS.n3577 0.0760357
R5908 VSS.n3581 VSS.n3579 0.0760357
R5909 VSS.n3583 VSS.n3581 0.0760357
R5910 VSS.n3585 VSS.n3583 0.0760357
R5911 VSS.n3587 VSS.n3585 0.0760357
R5912 VSS.n3589 VSS.n3587 0.0760357
R5913 VSS.n3591 VSS.n3589 0.0760357
R5914 VSS.n3593 VSS.n3591 0.0760357
R5915 VSS.n3595 VSS.n3593 0.0760357
R5916 VSS.n3597 VSS.n3595 0.0760357
R5917 VSS.n3599 VSS.n3597 0.0760357
R5918 VSS.n3601 VSS.n3599 0.0760357
R5919 VSS.n3603 VSS.n3601 0.0760357
R5920 VSS.n3605 VSS.n3603 0.0760357
R5921 VSS.n3607 VSS.n3605 0.0760357
R5922 VSS.n3609 VSS.n3607 0.0760357
R5923 VSS.n3611 VSS.n3609 0.0760357
R5924 VSS.n3613 VSS.n3611 0.0760357
R5925 VSS.n3615 VSS.n3613 0.0760357
R5926 VSS.n3617 VSS.n3615 0.0760357
R5927 VSS.n3619 VSS.n3617 0.0760357
R5928 VSS.n3621 VSS.n3619 0.0760357
R5929 VSS.n3623 VSS.n3621 0.0760357
R5930 VSS.n3625 VSS.n3623 0.0760357
R5931 VSS.n3627 VSS.n3625 0.0760357
R5932 VSS.n3629 VSS.n3627 0.0760357
R5933 VSS.n3631 VSS.n3629 0.0760357
R5934 VSS.n3633 VSS.n3631 0.0760357
R5935 VSS.n3635 VSS.n3633 0.0760357
R5936 VSS.n3637 VSS.n3635 0.0760357
R5937 VSS.n3639 VSS.n3637 0.0760357
R5938 VSS.n3641 VSS.n3639 0.0760357
R5939 VSS.n3643 VSS.n3641 0.0760357
R5940 VSS.n3646 VSS.n3643 0.0760357
R5941 VSS.n3648 VSS.n3646 0.0760357
R5942 VSS.n3651 VSS.n3648 0.0760357
R5943 VSS.n3653 VSS.n3651 0.0760357
R5944 VSS.n3656 VSS.n3653 0.0760357
R5945 VSS.n3658 VSS.n3656 0.0760357
R5946 VSS.n3661 VSS.n3658 0.0760357
R5947 VSS.n3663 VSS.n3661 0.0760357
R5948 VSS.n3666 VSS.n3663 0.0760357
R5949 VSS.n3668 VSS.n3666 0.0760357
R5950 VSS.n3671 VSS.n3668 0.0760357
R5951 VSS.n3673 VSS.n3671 0.0760357
R5952 VSS.n3730 VSS.n3673 0.0760357
R5953 VSS.n2216 VSS.n2214 0.0760357
R5954 VSS.n2218 VSS.n2216 0.0760357
R5955 VSS.n2220 VSS.n2218 0.0760357
R5956 VSS.n2222 VSS.n2220 0.0760357
R5957 VSS.n2224 VSS.n2222 0.0760357
R5958 VSS.n2226 VSS.n2224 0.0760357
R5959 VSS.n2228 VSS.n2226 0.0760357
R5960 VSS.n2230 VSS.n2228 0.0760357
R5961 VSS.n2232 VSS.n2230 0.0760357
R5962 VSS.n2234 VSS.n2232 0.0760357
R5963 VSS.n2236 VSS.n2234 0.0760357
R5964 VSS.n2238 VSS.n2236 0.0760357
R5965 VSS.n2240 VSS.n2238 0.0760357
R5966 VSS.n2242 VSS.n2240 0.0760357
R5967 VSS.n2244 VSS.n2242 0.0760357
R5968 VSS.n2246 VSS.n2244 0.0760357
R5969 VSS.n2248 VSS.n2246 0.0760357
R5970 VSS.n2250 VSS.n2248 0.0760357
R5971 VSS.n2252 VSS.n2250 0.0760357
R5972 VSS.n2254 VSS.n2252 0.0760357
R5973 VSS.n2256 VSS.n2254 0.0760357
R5974 VSS.n2258 VSS.n2256 0.0760357
R5975 VSS.n2260 VSS.n2258 0.0760357
R5976 VSS.n2262 VSS.n2260 0.0760357
R5977 VSS.n2264 VSS.n2262 0.0760357
R5978 VSS.n2266 VSS.n2264 0.0760357
R5979 VSS.n2268 VSS.n2266 0.0760357
R5980 VSS.n2270 VSS.n2268 0.0760357
R5981 VSS.n2272 VSS.n2270 0.0760357
R5982 VSS.n2275 VSS.n2272 0.0760357
R5983 VSS.n2277 VSS.n2275 0.0760357
R5984 VSS.n2280 VSS.n2277 0.0760357
R5985 VSS.n2282 VSS.n2280 0.0760357
R5986 VSS.n2285 VSS.n2282 0.0760357
R5987 VSS.n2287 VSS.n2285 0.0760357
R5988 VSS.n2290 VSS.n2287 0.0760357
R5989 VSS.n2292 VSS.n2290 0.0760357
R5990 VSS.n2295 VSS.n2292 0.0760357
R5991 VSS.n2297 VSS.n2295 0.0760357
R5992 VSS.n2701 VSS.n2700 0.068
R5993 VSS.n2681 VSS.n2680 0.068
R5994 VSS.n2183 VSS.n2181 0.0561875
R5995 VSS.n2185 VSS.n2183 0.055625
R5996 VSS.n2662 VSS.n2659 0.053375
R5997 VSS.n2659 VSS.n2656 0.053375
R5998 VSS.n2656 VSS.n2653 0.053375
R5999 VSS.n2653 VSS.n2651 0.053375
R6000 VSS.n2651 VSS.n2649 0.053375
R6001 VSS.n2649 VSS.n2647 0.053375
R6002 VSS.n2647 VSS.n2645 0.053375
R6003 VSS.n3370 VSS.n3368 0.053375
R6004 VSS.n3368 VSS.n3365 0.053375
R6005 VSS.n3365 VSS.n3363 0.053375
R6006 VSS.n3363 VSS.n3360 0.053375
R6007 VSS.n3360 VSS.n3358 0.053375
R6008 VSS.n3358 VSS.n3355 0.053375
R6009 VSS.n3355 VSS.n3353 0.053375
R6010 VSS.n3353 VSS.n3350 0.053375
R6011 VSS.n3350 VSS.n3348 0.053375
R6012 VSS.n3348 VSS.n3345 0.053375
R6013 VSS.n3345 VSS.n3343 0.053375
R6014 VSS.n3343 VSS.n3340 0.053375
R6015 VSS.n3340 VSS.n3338 0.053375
R6016 VSS.n3338 VSS.n3335 0.053375
R6017 VSS.n3335 VSS.n3333 0.053375
R6018 VSS.n2637 VSS.n2635 0.053375
R6019 VSS.n2635 VSS.n2633 0.053375
R6020 VSS.n2633 VSS.n2631 0.053375
R6021 VSS.n2587 VSS.n2585 0.053375
R6022 VSS.n2585 VSS.n2582 0.053375
R6023 VSS.n2582 VSS.n2580 0.053375
R6024 VSS.n2580 VSS.n2577 0.053375
R6025 VSS.n2577 VSS.n2575 0.053375
R6026 VSS.n2575 VSS.n2572 0.053375
R6027 VSS.n2572 VSS.n2570 0.053375
R6028 VSS.n2859 VSS.n2857 0.053375
R6029 VSS.n2861 VSS.n2859 0.053375
R6030 VSS.n3927 VSS.n3925 0.053375
R6031 VSS.n3925 VSS.n3922 0.053375
R6032 VSS.n3922 VSS.n3920 0.053375
R6033 VSS.n3920 VSS.n3917 0.053375
R6034 VSS.n3917 VSS.n3915 0.053375
R6035 VSS.n3915 VSS.n3912 0.053375
R6036 VSS.n3912 VSS.n3910 0.053375
R6037 VSS.n3910 VSS.n3907 0.053375
R6038 VSS.n3907 VSS.n3905 0.053375
R6039 VSS.n3905 VSS.n3902 0.053375
R6040 VSS.n3902 VSS.n3900 0.053375
R6041 VSS.n3900 VSS.n3897 0.053375
R6042 VSS.n3897 VSS.n3895 0.053375
R6043 VSS.n3895 VSS.n3892 0.053375
R6044 VSS.n242 VSS.n241 0.053375
R6045 VSS.n241 VSS.n240 0.053375
R6046 VSS.n240 VSS.n239 0.053375
R6047 VSS.n239 VSS.n238 0.053375
R6048 VSS.n238 VSS.n237 0.053375
R6049 VSS.n4044 VSS.n4042 0.053375
R6050 VSS.n4042 VSS.n4039 0.053375
R6051 VSS.n4039 VSS.n4037 0.053375
R6052 VSS.n4037 VSS.n4034 0.053375
R6053 VSS.n4034 VSS.n4032 0.053375
R6054 VSS.n4032 VSS.n4029 0.053375
R6055 VSS.n4029 VSS.n4027 0.053375
R6056 VSS.n4027 VSS.n4024 0.053375
R6057 VSS.n4024 VSS.n4022 0.053375
R6058 VSS.n4022 VSS.n4019 0.053375
R6059 VSS.n4019 VSS.n4017 0.053375
R6060 VSS.n4017 VSS.n4014 0.053375
R6061 VSS.n4014 VSS.n4012 0.053375
R6062 VSS.n4012 VSS.n4009 0.053375
R6063 VSS.n4009 VSS.n4007 0.053375
R6064 VSS.n4007 VSS.n4004 0.053375
R6065 VSS.n4004 VSS.n4002 0.053375
R6066 VSS.n4002 VSS.n4000 0.053375
R6067 VSS.n4000 VSS.n3998 0.053375
R6068 VSS.n3998 VSS.n3996 0.053375
R6069 VSS.n3996 VSS.n3994 0.053375
R6070 VSS.n3994 VSS.n3992 0.053375
R6071 VSS.n3992 VSS.n3990 0.053375
R6072 VSS.n3990 VSS.n3988 0.053375
R6073 VSS.n3988 VSS.n3986 0.053375
R6074 VSS.n3986 VSS.n3984 0.053375
R6075 VSS.n3984 VSS.n3982 0.053375
R6076 VSS.n3982 VSS.n3980 0.053375
R6077 VSS.n3980 VSS.n3978 0.053375
R6078 VSS.n3978 VSS.n3976 0.053375
R6079 VSS.n3976 VSS.n3974 0.053375
R6080 VSS.n3974 VSS.n3972 0.053375
R6081 VSS.n3972 VSS.n3970 0.053375
R6082 VSS.n3968 VSS.n3967 0.053375
R6083 VSS.n3967 VSS.n3964 0.053375
R6084 VSS.n3964 VSS.n3961 0.053375
R6085 VSS.n3961 VSS.n3958 0.053375
R6086 VSS.n3958 VSS.n3955 0.053375
R6087 VSS.n3955 VSS.n3952 0.053375
R6088 VSS.n3944 VSS.n3941 0.053375
R6089 VSS.n3937 VSS.n3934 0.053375
R6090 VSS.n3934 VSS.n3931 0.053375
R6091 VSS.n2957 VSS.n2955 0.053375
R6092 VSS.n2952 VSS.n2950 0.053375
R6093 VSS.n2945 VSS.n2943 0.053375
R6094 VSS.n2937 VSS.n2935 0.053375
R6095 VSS.n2932 VSS.n2930 0.053375
R6096 VSS.n2924 VSS.n2922 0.053375
R6097 VSS.n2922 VSS.n2920 0.053375
R6098 VSS.n2920 VSS.n2918 0.053375
R6099 VSS.n2918 VSS.n2916 0.053375
R6100 VSS.n2916 VSS.n2914 0.053375
R6101 VSS.n2914 VSS.n2912 0.053375
R6102 VSS.n2912 VSS.n2910 0.053375
R6103 VSS.n2910 VSS.n2908 0.053375
R6104 VSS.n2908 VSS.n2906 0.053375
R6105 VSS.n2906 VSS.n2904 0.053375
R6106 VSS.n2904 VSS.n2902 0.053375
R6107 VSS.n2902 VSS.n2900 0.053375
R6108 VSS.n2900 VSS.n2898 0.053375
R6109 VSS.n2898 VSS.n2896 0.053375
R6110 VSS.n2896 VSS.n2894 0.053375
R6111 VSS.n2891 VSS.n2889 0.053375
R6112 VSS.n2889 VSS.n2887 0.053375
R6113 VSS.n2887 VSS.n2885 0.053375
R6114 VSS.n2885 VSS.n2883 0.053375
R6115 VSS.n2880 VSS.n2878 0.053375
R6116 VSS.n2878 VSS.n2876 0.053375
R6117 VSS.n3854 VSS.n3852 0.053375
R6118 VSS.n3856 VSS.n3854 0.053375
R6119 VSS.n3858 VSS.n3856 0.053375
R6120 VSS.n3860 VSS.n3858 0.053375
R6121 VSS.n3865 VSS.n3863 0.053375
R6122 VSS.n3867 VSS.n3865 0.053375
R6123 VSS.n3869 VSS.n3867 0.053375
R6124 VSS.n3874 VSS.n3872 0.053375
R6125 VSS.n3876 VSS.n3874 0.053375
R6126 VSS.n3878 VSS.n3876 0.053375
R6127 VSS.n3883 VSS.n3881 0.053375
R6128 VSS.n3888 VSS.n3886 0.053375
R6129 VSS.n3890 VSS.n3888 0.053375
R6130 VSS.n2600 VSS.n2597 0.053375
R6131 VSS.n2607 VSS.n2604 0.053375
R6132 VSS.n2614 VSS.n2611 0.053375
R6133 VSS.n2617 VSS.n2614 0.053375
R6134 VSS.n2620 VSS.n2617 0.053375
R6135 VSS.n2623 VSS.n2620 0.053375
R6136 VSS.n2626 VSS.n2623 0.053375
R6137 VSS.n2629 VSS.n2626 0.053375
R6138 VSS.n2530 VSS.n2527 0.053375
R6139 VSS.n2527 VSS.n2524 0.053375
R6140 VSS.n2524 VSS.n2521 0.053375
R6141 VSS.n2517 VSS.n2514 0.053375
R6142 VSS.n2510 VSS.n2507 0.053375
R6143 VSS.n2507 VSS.n2504 0.053375
R6144 VSS.n2504 VSS.n2501 0.053375
R6145 VSS.n2501 VSS.n2498 0.053375
R6146 VSS.n2498 VSS.n2495 0.053375
R6147 VSS.n2495 VSS.n2492 0.053375
R6148 VSS.n2492 VSS.n2489 0.053375
R6149 VSS.n2489 VSS.n2485 0.053375
R6150 VSS.n2485 VSS.n2482 0.053375
R6151 VSS.n3792 VSS.n3789 0.053375
R6152 VSS.n3795 VSS.n3792 0.053375
R6153 VSS.n3798 VSS.n3795 0.053375
R6154 VSS.n3801 VSS.n3798 0.053375
R6155 VSS.n3804 VSS.n3801 0.053375
R6156 VSS.n3807 VSS.n3804 0.053375
R6157 VSS.n3810 VSS.n3807 0.053375
R6158 VSS.n3813 VSS.n3810 0.053375
R6159 VSS.n3816 VSS.n3813 0.053375
R6160 VSS.n3823 VSS.n3820 0.053375
R6161 VSS.n3830 VSS.n3827 0.053375
R6162 VSS.n3833 VSS.n3830 0.053375
R6163 VSS.n3836 VSS.n3833 0.053375
R6164 VSS.n357 VSS.n355 0.053375
R6165 VSS.n349 VSS.n347 0.053375
R6166 VSS.n347 VSS.n345 0.053375
R6167 VSS.n342 VSS.n340 0.053375
R6168 VSS.n340 VSS.n338 0.053375
R6169 VSS.n338 VSS.n336 0.053375
R6170 VSS.n333 VSS.n331 0.053375
R6171 VSS.n331 VSS.n329 0.053375
R6172 VSS.n326 VSS.n324 0.053375
R6173 VSS.n324 VSS.n322 0.053375
R6174 VSS.n322 VSS.n320 0.053375
R6175 VSS.n317 VSS.n315 0.053375
R6176 VSS.n315 VSS.n313 0.053375
R6177 VSS.n304 VSS.n302 0.053375
R6178 VSS.n302 VSS.n300 0.053375
R6179 VSS.n3752 VSS.n3749 0.053375
R6180 VSS.n3749 VSS.n3746 0.053375
R6181 VSS.n3738 VSS.n3735 0.053375
R6182 VSS.n3735 VSS.n3732 0.053375
R6183 VSS.n3389 VSS.n3386 0.053375
R6184 VSS.n3392 VSS.n3389 0.053375
R6185 VSS.n3395 VSS.n3392 0.053375
R6186 VSS.n3398 VSS.n3395 0.053375
R6187 VSS.n3401 VSS.n3398 0.053375
R6188 VSS.n3404 VSS.n3401 0.053375
R6189 VSS.n3407 VSS.n3404 0.053375
R6190 VSS.n3410 VSS.n3407 0.053375
R6191 VSS.n3413 VSS.n3410 0.053375
R6192 VSS.n3416 VSS.n3413 0.053375
R6193 VSS.n3419 VSS.n3416 0.053375
R6194 VSS.n3426 VSS.n3423 0.053375
R6195 VSS VSS.n3430 0.053375
R6196 VSS VSS.n4113 0.053375
R6197 VSS.n4113 VSS.n4110 0.053375
R6198 VSS.n4102 VSS.n4099 0.053375
R6199 VSS.n4099 VSS.n4096 0.053375
R6200 VSS.n4092 VSS.n4089 0.053375
R6201 VSS.n4089 VSS.n4086 0.053375
R6202 VSS.n4086 VSS.n4083 0.053375
R6203 VSS.n4079 VSS.n4076 0.053375
R6204 VSS.n4076 VSS.n4073 0.053375
R6205 VSS.n4069 VSS.n4066 0.053375
R6206 VSS.n2420 VSS.n2417 0.053375
R6207 VSS.n2427 VSS.n2424 0.053375
R6208 VSS.n2440 VSS.n2437 0.053375
R6209 VSS.n2443 VSS.n2440 0.053375
R6210 VSS.n2446 VSS.n2443 0.053375
R6211 VSS.n2449 VSS.n2446 0.053375
R6212 VSS.n2452 VSS.n2449 0.053375
R6213 VSS.n2455 VSS.n2452 0.053375
R6214 VSS.n2458 VSS.n2455 0.053375
R6215 VSS.n10 VSS.n8 0.053375
R6216 VSS.n15 VSS.n13 0.053375
R6217 VSS.n20 VSS.n18 0.053375
R6218 VSS.n22 VSS.n20 0.053375
R6219 VSS.n24 VSS.n22 0.053375
R6220 VSS.n26 VSS.n24 0.053375
R6221 VSS.n28 VSS.n26 0.053375
R6222 VSS.n30 VSS.n28 0.053375
R6223 VSS.n32 VSS.n30 0.053375
R6224 VSS.n34 VSS.n32 0.053375
R6225 VSS.n39 VSS.n37 0.053375
R6226 VSS.n41 VSS.n39 0.053375
R6227 VSS.n43 VSS.n41 0.053375
R6228 VSS.n45 VSS.n43 0.053375
R6229 VSS.n47 VSS.n45 0.053375
R6230 VSS.n49 VSS.n47 0.053375
R6231 VSS.n54 VSS.n52 0.053375
R6232 VSS.n56 VSS.n54 0.053375
R6233 VSS.n58 VSS.n56 0.053375
R6234 VSS.n63 VSS.n61 0.053375
R6235 VSS.n228 VSS.n226 0.053375
R6236 VSS.n226 VSS.n224 0.053375
R6237 VSS.n224 VSS.n222 0.053375
R6238 VSS.n222 VSS.n68 0.053375
R6239 VSS.n2181 VSS.n2179 0.053375
R6240 VSS.n2187 VSS.n2185 0.053375
R6241 VSS.n2189 VSS.n2187 0.053375
R6242 VSS.n2191 VSS.n2189 0.053375
R6243 VSS.n2193 VSS.n2191 0.053375
R6244 VSS.n2195 VSS.n2193 0.053375
R6245 VSS.n2197 VSS.n2195 0.053375
R6246 VSS.n2199 VSS.n2197 0.053375
R6247 VSS.n2201 VSS.n2199 0.053375
R6248 VSS.n2203 VSS.n2201 0.053375
R6249 VSS.n2205 VSS.n2203 0.053375
R6250 VSS.n2207 VSS.n2205 0.053375
R6251 VSS.n2209 VSS.n2207 0.053375
R6252 VSS.n4066 VSS.n4063 0.0530441
R6253 VSS.n3870 VSS.n3869 0.0528125
R6254 VSS.n2461 VSS.n2458 0.05275
R6255 VSS.n2941 VSS.n2940 0.0505625
R6256 VSS.n2179 VSS.n2177 0.0505625
R6257 VSS.n2521 VSS.n2518 0.05
R6258 VSS.n3827 VSS.n3824 0.048875
R6259 VSS.n3430 VSS.n3427 0.0483125
R6260 VSS.n2421 VSS.n2420 0.0483125
R6261 VSS.n6 VSS.n5 0.0483125
R6262 VSS.n66 VSS.n64 0.0483125
R6263 VSS.n345 VSS.n343 0.04775
R6264 VSS.n318 VSS.n317 0.04775
R6265 VSS.n4096 VSS.n4093 0.04775
R6266 VSS.n353 VSS.n352 0.046625
R6267 VSS.n307 VSS.n305 0.046625
R6268 VSS.n3742 VSS.n3739 0.046625
R6269 VSS.n4107 VSS.n4106 0.046625
R6270 VSS.n2927 VSS.n2925 0.0460625
R6271 VSS.n37 VSS.n35 0.0460625
R6272 VSS.n2928 VSS.n2927 0.0449375
R6273 VSS.n352 VSS.n350 0.044375
R6274 VSS.n311 VSS.n307 0.044375
R6275 VSS.n3743 VSS.n3742 0.044375
R6276 VSS.n4106 VSS.n4103 0.044375
R6277 VSS.n2881 VSS.n2880 0.0426875
R6278 VSS.n3850 VSS.n3849 0.0426875
R6279 VSS.n2700 VSS.n2699 0.0410839
R6280 VSS.n2680 VSS.n2679 0.0410839
R6281 VSS.n2940 VSS.n2938 0.0404375
R6282 VSS.n2210 VSS.n66 0.039875
R6283 VSS.n358 VSS.n357 0.037625
R6284 VSS.n334 VSS.n333 0.037625
R6285 VSS.n329 VSS.n327 0.037625
R6286 VSS.n4080 VSS.n4079 0.037625
R6287 VSS.n4073 VSS.n4070 0.037625
R6288 VSS.n4060 VSS.n3772 0.0354412
R6289 VSS.n4058 VSS.n3836 0.0349634
R6290 VSS.n3381 VSS.n2530 0.0349492
R6291 VSS.n3952 VSS.n3949 0.0348125
R6292 VSS.n3938 VSS.n3937 0.0348125
R6293 VSS.n2955 VSS.n2953 0.0348125
R6294 VSS.n2948 VSS.n2945 0.0348125
R6295 VSS.n3879 VSS.n3878 0.0348125
R6296 VSS.n3886 VSS.n3884 0.0348125
R6297 VSS.n2601 VSS.n2600 0.0348125
R6298 VSS.n2611 VSS.n2608 0.0348125
R6299 VSS.n2177 VSS.n68 0.0348125
R6300 VSS.n2514 VSS.n2511 0.03425
R6301 VSS.n50 VSS.n49 0.03425
R6302 VSS.n2465 VSS.n2462 0.0335
R6303 VSS.n3820 VSS.n3817 0.033125
R6304 VSS.n2894 VSS.n2892 0.0325625
R6305 VSS.n3863 VSS.n3861 0.0325625
R6306 VSS.n3423 VSS.n3420 0.0325625
R6307 VSS.n2434 VSS.n2427 0.0325625
R6308 VSS.n11 VSS.n10 0.0325625
R6309 VSS.n61 VSS.n59 0.0325625
R6310 VSS.n2597 VSS.n2594 0.030875
R6311 VSS.n2958 VSS.n2957 0.030875
R6312 VSS.n3753 VSS.n3752 0.0307426
R6313 VSS.n3386 VSS.n3383 0.029625
R6314 VSS.n2933 VSS.n2932 0.0291875
R6315 VSS.n18 VSS.n16 0.0280625
R6316 VSS.n3007 VSS.n3005 0.0269375
R6317 VSS.n3005 VSS.n3002 0.0269375
R6318 VSS.n3002 VSS.n3000 0.0269375
R6319 VSS.n3000 VSS.n2997 0.0269375
R6320 VSS.n2997 VSS.n2995 0.0269375
R6321 VSS.n2995 VSS.n2992 0.0269375
R6322 VSS.n2989 VSS.n2986 0.0269375
R6323 VSS.n2986 VSS.n2984 0.0269375
R6324 VSS.n2981 VSS.n2979 0.0269375
R6325 VSS.n2979 VSS.n2977 0.0269375
R6326 VSS.n2977 VSS.n2975 0.0269375
R6327 VSS.n2975 VSS.n2973 0.0269375
R6328 VSS.n2973 VSS.n2971 0.0269375
R6329 VSS.n2971 VSS.n2969 0.0269375
R6330 VSS.n2969 VSS.n2967 0.0269375
R6331 VSS.n2967 VSS.n2965 0.0269375
R6332 VSS.n2965 VSS.n2963 0.0269375
R6333 VSS.n2730 VSS.n2727 0.0269375
R6334 VSS.n2732 VSS.n2730 0.0269375
R6335 VSS.n2735 VSS.n2732 0.0269375
R6336 VSS.n2738 VSS.n2735 0.0269375
R6337 VSS.n2740 VSS.n2738 0.0269375
R6338 VSS.n2742 VSS.n2740 0.0269375
R6339 VSS.n2747 VSS.n2745 0.0269375
R6340 VSS.n2749 VSS.n2747 0.0269375
R6341 VSS.n2754 VSS.n2752 0.0269375
R6342 VSS.n2756 VSS.n2754 0.0269375
R6343 VSS.n2758 VSS.n2756 0.0269375
R6344 VSS.n2760 VSS.n2758 0.0269375
R6345 VSS.n2762 VSS.n2760 0.0269375
R6346 VSS.n2767 VSS.n2765 0.0269375
R6347 VSS.n2769 VSS.n2767 0.0269375
R6348 VSS.n2771 VSS.n2769 0.0269375
R6349 VSS.n2773 VSS.n2771 0.0269375
R6350 VSS.n2775 VSS.n2773 0.0269375
R6351 VSS.n2777 VSS.n2775 0.0269375
R6352 VSS.n2782 VSS.n2780 0.0269375
R6353 VSS.n2784 VSS.n2782 0.0269375
R6354 VSS.n2786 VSS.n2784 0.0269375
R6355 VSS.n2788 VSS.n2786 0.0269375
R6356 VSS.n2790 VSS.n2788 0.0269375
R6357 VSS.n2792 VSS.n2790 0.0269375
R6358 VSS.n2794 VSS.n2792 0.0269375
R6359 VSS.n2799 VSS.n2797 0.0269375
R6360 VSS.n2801 VSS.n2799 0.0269375
R6361 VSS.n2803 VSS.n2801 0.0269375
R6362 VSS.n2805 VSS.n2803 0.0269375
R6363 VSS.n2807 VSS.n2805 0.0269375
R6364 VSS.n2812 VSS.n2810 0.0269375
R6365 VSS.n2814 VSS.n2812 0.0269375
R6366 VSS.n2816 VSS.n2814 0.0269375
R6367 VSS.n2818 VSS.n2816 0.0269375
R6368 VSS.n2820 VSS.n2818 0.0269375
R6369 VSS.n2822 VSS.n2820 0.0269375
R6370 VSS.n2824 VSS.n2822 0.0269375
R6371 VSS.n2826 VSS.n2824 0.0269375
R6372 VSS.n2828 VSS.n2826 0.0269375
R6373 VSS.n2830 VSS.n2828 0.0269375
R6374 VSS.n2835 VSS.n2833 0.0269375
R6375 VSS.n2837 VSS.n2835 0.0269375
R6376 VSS.n2842 VSS.n2840 0.0269375
R6377 VSS.n2844 VSS.n2842 0.0269375
R6378 VSS.n2846 VSS.n2844 0.0269375
R6379 VSS.n2848 VSS.n2846 0.0269375
R6380 VSS.n2850 VSS.n2848 0.0269375
R6381 VSS.n2852 VSS.n2850 0.0269375
R6382 VSS.n3123 VSS.n3120 0.0269375
R6383 VSS.n3120 VSS.n3117 0.0269375
R6384 VSS.n3117 VSS.n3114 0.0269375
R6385 VSS.n3114 VSS.n3111 0.0269375
R6386 VSS.n3111 VSS.n3108 0.0269375
R6387 VSS.n3108 VSS.n3105 0.0269375
R6388 VSS.n3105 VSS.n3102 0.0269375
R6389 VSS.n3102 VSS.n3099 0.0269375
R6390 VSS.n3099 VSS.n3096 0.0269375
R6391 VSS.n3096 VSS.n3093 0.0269375
R6392 VSS.n3093 VSS.n3090 0.0269375
R6393 VSS.n3090 VSS.n3087 0.0269375
R6394 VSS.n3087 VSS.n3084 0.0269375
R6395 VSS.n3084 VSS.n3081 0.0269375
R6396 VSS.n3081 VSS.n3078 0.0269375
R6397 VSS.n3078 VSS.n3075 0.0269375
R6398 VSS.n3075 VSS.n3072 0.0269375
R6399 VSS.n3072 VSS.n3069 0.0269375
R6400 VSS.n3069 VSS.n3066 0.0269375
R6401 VSS.n3066 VSS.n3063 0.0269375
R6402 VSS.n3063 VSS.n3060 0.0269375
R6403 VSS.n3060 VSS.n3057 0.0269375
R6404 VSS.n3057 VSS.n3054 0.0269375
R6405 VSS.n3054 VSS.n3051 0.0269375
R6406 VSS.n2721 VSS.n2718 0.0269375
R6407 VSS.n2724 VSS.n2721 0.0269375
R6408 VSS.n3136 VSS.n3134 0.0269375
R6409 VSS.n3139 VSS.n3136 0.0269375
R6410 VSS.n3141 VSS.n3139 0.0269375
R6411 VSS.n3144 VSS.n3141 0.0269375
R6412 VSS.n3148 VSS.n3144 0.0269375
R6413 VSS.n3151 VSS.n3148 0.0269375
R6414 VSS.n3158 VSS.n3155 0.0269375
R6415 VSS.n3161 VSS.n3158 0.0269375
R6416 VSS.n3168 VSS.n3165 0.0269375
R6417 VSS.n3171 VSS.n3168 0.0269375
R6418 VSS.n3174 VSS.n3171 0.0269375
R6419 VSS.n3177 VSS.n3174 0.0269375
R6420 VSS.n3180 VSS.n3177 0.0269375
R6421 VSS.n3187 VSS.n3184 0.0269375
R6422 VSS.n3190 VSS.n3187 0.0269375
R6423 VSS.n3193 VSS.n3190 0.0269375
R6424 VSS.n3196 VSS.n3193 0.0269375
R6425 VSS.n3199 VSS.n3196 0.0269375
R6426 VSS.n3202 VSS.n3199 0.0269375
R6427 VSS.n3209 VSS.n3206 0.0269375
R6428 VSS.n3212 VSS.n3209 0.0269375
R6429 VSS.n3215 VSS.n3212 0.0269375
R6430 VSS.n3218 VSS.n3215 0.0269375
R6431 VSS.n3221 VSS.n3218 0.0269375
R6432 VSS.n3224 VSS.n3221 0.0269375
R6433 VSS.n3227 VSS.n3224 0.0269375
R6434 VSS.n3234 VSS.n3231 0.0269375
R6435 VSS.n3237 VSS.n3234 0.0269375
R6436 VSS.n3240 VSS.n3237 0.0269375
R6437 VSS.n3243 VSS.n3240 0.0269375
R6438 VSS.n3246 VSS.n3243 0.0269375
R6439 VSS.n3253 VSS.n3250 0.0269375
R6440 VSS.n3256 VSS.n3253 0.0269375
R6441 VSS.n3259 VSS.n3256 0.0269375
R6442 VSS.n3262 VSS.n3259 0.0269375
R6443 VSS.n3265 VSS.n3262 0.0269375
R6444 VSS.n3268 VSS.n3265 0.0269375
R6445 VSS.n3279 VSS.n3276 0.0269375
R6446 VSS.n3290 VSS.n3287 0.0269375
R6447 VSS.n3293 VSS.n3290 0.0269375
R6448 VSS.n3300 VSS.n3297 0.0269375
R6449 VSS.n3303 VSS.n3300 0.0269375
R6450 VSS.n3306 VSS.n3303 0.0269375
R6451 VSS.n3309 VSS.n3306 0.0269375
R6452 VSS.n3312 VSS.n3309 0.0269375
R6453 VSS.n3315 VSS.n3312 0.0269375
R6454 VSS.n1400 VSS.n1398 0.0269375
R6455 VSS.n1403 VSS.n1400 0.0269375
R6456 VSS.n1406 VSS.n1403 0.0269375
R6457 VSS.n1408 VSS.n1406 0.0269375
R6458 VSS.n1411 VSS.n1408 0.0269375
R6459 VSS.n1295 VSS.n220 0.0269375
R6460 VSS.n220 VSS.n217 0.0269375
R6461 VSS.n217 VSS.n214 0.0269375
R6462 VSS.n214 VSS.n211 0.0269375
R6463 VSS.n211 VSS.n208 0.0269375
R6464 VSS.n208 VSS.n205 0.0269375
R6465 VSS.n205 VSS.n202 0.0269375
R6466 VSS.n202 VSS.n199 0.0269375
R6467 VSS.n199 VSS.n196 0.0269375
R6468 VSS.n196 VSS.n193 0.0269375
R6469 VSS.n193 VSS.n190 0.0269375
R6470 VSS.n190 VSS.n187 0.0269375
R6471 VSS.n187 VSS.n184 0.0269375
R6472 VSS.n184 VSS.n181 0.0269375
R6473 VSS.n181 VSS.n178 0.0269375
R6474 VSS.n178 VSS.n175 0.0269375
R6475 VSS.n175 VSS.n172 0.0269375
R6476 VSS.n172 VSS.n169 0.0269375
R6477 VSS.n169 VSS.n166 0.0269375
R6478 VSS.n166 VSS.n164 0.0269375
R6479 VSS.n164 VSS.n162 0.0269375
R6480 VSS.n162 VSS.n160 0.0269375
R6481 VSS.n160 VSS.n158 0.0269375
R6482 VSS.n158 VSS.n156 0.0269375
R6483 VSS.n156 VSS.n154 0.0269375
R6484 VSS.n154 VSS.n152 0.0269375
R6485 VSS.n152 VSS.n150 0.0269375
R6486 VSS.n150 VSS.n148 0.0269375
R6487 VSS.n148 VSS.n146 0.0269375
R6488 VSS.n146 VSS.n144 0.0269375
R6489 VSS.n144 VSS.n142 0.0269375
R6490 VSS.n142 VSS.n140 0.0269375
R6491 VSS.n140 VSS.n138 0.0269375
R6492 VSS.n138 VSS.n136 0.0269375
R6493 VSS.n136 VSS.n134 0.0269375
R6494 VSS.n134 VSS.n132 0.0269375
R6495 VSS.n132 VSS.n130 0.0269375
R6496 VSS.n130 VSS.n128 0.0269375
R6497 VSS.n128 VSS.n126 0.0269375
R6498 VSS.n126 VSS.n124 0.0269375
R6499 VSS.n124 VSS.n122 0.0269375
R6500 VSS.n122 VSS.n120 0.0269375
R6501 VSS.n120 VSS.n118 0.0269375
R6502 VSS.n118 VSS.n116 0.0269375
R6503 VSS.n116 VSS.n114 0.0269375
R6504 VSS.n114 VSS.n112 0.0269375
R6505 VSS.n112 VSS.n110 0.0269375
R6506 VSS.n110 VSS.n108 0.0269375
R6507 VSS.n108 VSS.n106 0.0269375
R6508 VSS.n106 VSS.n104 0.0269375
R6509 VSS.n104 VSS.n102 0.0269375
R6510 VSS.n102 VSS.n100 0.0269375
R6511 VSS.n100 VSS.n98 0.0269375
R6512 VSS.n98 VSS.n96 0.0269375
R6513 VSS.n96 VSS.n94 0.0269375
R6514 VSS.n94 VSS.n92 0.0269375
R6515 VSS.n92 VSS.n90 0.0269375
R6516 VSS.n1522 VSS.n1520 0.0269375
R6517 VSS.n1524 VSS.n1522 0.0269375
R6518 VSS.n1526 VSS.n1524 0.0269375
R6519 VSS.n1528 VSS.n1526 0.0269375
R6520 VSS.n1530 VSS.n1528 0.0269375
R6521 VSS.n1952 VSS.n1530 0.0269375
R6522 VSS.n1210 VSS.n483 0.0269375
R6523 VSS.n483 VSS.n481 0.0269375
R6524 VSS.n481 VSS.n478 0.0269375
R6525 VSS.n478 VSS.n475 0.0269375
R6526 VSS.n475 VSS.n473 0.0269375
R6527 VSS.n473 VSS.n470 0.0269375
R6528 VSS.n470 VSS.n468 0.0269375
R6529 VSS.n468 VSS.n465 0.0269375
R6530 VSS.n465 VSS.n463 0.0269375
R6531 VSS.n463 VSS.n460 0.0269375
R6532 VSS.n460 VSS.n458 0.0269375
R6533 VSS.n458 VSS.n455 0.0269375
R6534 VSS.n455 VSS.n453 0.0269375
R6535 VSS.n453 VSS.n451 0.0269375
R6536 VSS.n451 VSS.n449 0.0269375
R6537 VSS.n449 VSS.n447 0.0269375
R6538 VSS.n447 VSS.n445 0.0269375
R6539 VSS.n445 VSS.n443 0.0269375
R6540 VSS.n443 VSS.n441 0.0269375
R6541 VSS.n441 VSS.n439 0.0269375
R6542 VSS.n439 VSS.n437 0.0269375
R6543 VSS.n437 VSS.n435 0.0269375
R6544 VSS.n435 VSS.n433 0.0269375
R6545 VSS.n433 VSS.n431 0.0269375
R6546 VSS.n431 VSS.n429 0.0269375
R6547 VSS.n429 VSS.n427 0.0269375
R6548 VSS.n427 VSS.n425 0.0269375
R6549 VSS.n425 VSS.n423 0.0269375
R6550 VSS.n423 VSS.n421 0.0269375
R6551 VSS.n421 VSS.n419 0.0269375
R6552 VSS.n419 VSS.n417 0.0269375
R6553 VSS.n417 VSS.n415 0.0269375
R6554 VSS.n415 VSS.n413 0.0269375
R6555 VSS.n413 VSS.n411 0.0269375
R6556 VSS.n411 VSS.n409 0.0269375
R6557 VSS.n409 VSS.n407 0.0269375
R6558 VSS.n407 VSS.n405 0.0269375
R6559 VSS.n405 VSS.n403 0.0269375
R6560 VSS.n403 VSS.n401 0.0269375
R6561 VSS.n401 VSS.n399 0.0269375
R6562 VSS.n399 VSS.n397 0.0269375
R6563 VSS.n397 VSS.n395 0.0269375
R6564 VSS.n395 VSS.n393 0.0269375
R6565 VSS.n393 VSS.n391 0.0269375
R6566 VSS.n391 VSS.n389 0.0269375
R6567 VSS.n389 VSS.n387 0.0269375
R6568 VSS.n387 VSS.n385 0.0269375
R6569 VSS.n385 VSS.n383 0.0269375
R6570 VSS.n383 VSS.n381 0.0269375
R6571 VSS.n381 VSS.n379 0.0269375
R6572 VSS.n379 VSS.n377 0.0269375
R6573 VSS.n377 VSS.n375 0.0269375
R6574 VSS.n375 VSS.n373 0.0269375
R6575 VSS.n373 VSS.n371 0.0269375
R6576 VSS.n371 VSS.n369 0.0269375
R6577 VSS.n369 VSS.n367 0.0269375
R6578 VSS.n367 VSS.n365 0.0269375
R6579 VSS.n1534 VSS.n1532 0.0269375
R6580 VSS.n1536 VSS.n1534 0.0269375
R6581 VSS.n1538 VSS.n1536 0.0269375
R6582 VSS.n1540 VSS.n1538 0.0269375
R6583 VSS.n1542 VSS.n1540 0.0269375
R6584 VSS.n1943 VSS.n1542 0.0269375
R6585 VSS.n1112 VSS.n635 0.0269375
R6586 VSS.n635 VSS.n632 0.0269375
R6587 VSS.n632 VSS.n629 0.0269375
R6588 VSS.n629 VSS.n626 0.0269375
R6589 VSS.n626 VSS.n623 0.0269375
R6590 VSS.n623 VSS.n620 0.0269375
R6591 VSS.n620 VSS.n617 0.0269375
R6592 VSS.n617 VSS.n614 0.0269375
R6593 VSS.n614 VSS.n611 0.0269375
R6594 VSS.n611 VSS.n608 0.0269375
R6595 VSS.n608 VSS.n605 0.0269375
R6596 VSS.n605 VSS.n602 0.0269375
R6597 VSS.n602 VSS.n599 0.0269375
R6598 VSS.n599 VSS.n596 0.0269375
R6599 VSS.n596 VSS.n593 0.0269375
R6600 VSS.n593 VSS.n590 0.0269375
R6601 VSS.n590 VSS.n587 0.0269375
R6602 VSS.n587 VSS.n584 0.0269375
R6603 VSS.n584 VSS.n581 0.0269375
R6604 VSS.n581 VSS.n579 0.0269375
R6605 VSS.n579 VSS.n577 0.0269375
R6606 VSS.n577 VSS.n575 0.0269375
R6607 VSS.n575 VSS.n573 0.0269375
R6608 VSS.n573 VSS.n571 0.0269375
R6609 VSS.n571 VSS.n569 0.0269375
R6610 VSS.n569 VSS.n567 0.0269375
R6611 VSS.n567 VSS.n565 0.0269375
R6612 VSS.n565 VSS.n563 0.0269375
R6613 VSS.n563 VSS.n561 0.0269375
R6614 VSS.n561 VSS.n559 0.0269375
R6615 VSS.n559 VSS.n557 0.0269375
R6616 VSS.n557 VSS.n555 0.0269375
R6617 VSS.n555 VSS.n553 0.0269375
R6618 VSS.n553 VSS.n551 0.0269375
R6619 VSS.n551 VSS.n549 0.0269375
R6620 VSS.n549 VSS.n547 0.0269375
R6621 VSS.n547 VSS.n545 0.0269375
R6622 VSS.n545 VSS.n543 0.0269375
R6623 VSS.n543 VSS.n541 0.0269375
R6624 VSS.n541 VSS.n539 0.0269375
R6625 VSS.n539 VSS.n537 0.0269375
R6626 VSS.n537 VSS.n535 0.0269375
R6627 VSS.n535 VSS.n533 0.0269375
R6628 VSS.n533 VSS.n531 0.0269375
R6629 VSS.n531 VSS.n529 0.0269375
R6630 VSS.n529 VSS.n527 0.0269375
R6631 VSS.n527 VSS.n525 0.0269375
R6632 VSS.n525 VSS.n523 0.0269375
R6633 VSS.n523 VSS.n521 0.0269375
R6634 VSS.n521 VSS.n519 0.0269375
R6635 VSS.n519 VSS.n517 0.0269375
R6636 VSS.n517 VSS.n515 0.0269375
R6637 VSS.n515 VSS.n513 0.0269375
R6638 VSS.n513 VSS.n511 0.0269375
R6639 VSS.n511 VSS.n509 0.0269375
R6640 VSS.n509 VSS.n507 0.0269375
R6641 VSS.n507 VSS.n505 0.0269375
R6642 VSS.n1652 VSS.n1650 0.0269375
R6643 VSS.n1654 VSS.n1652 0.0269375
R6644 VSS.n1656 VSS.n1654 0.0269375
R6645 VSS.n1658 VSS.n1656 0.0269375
R6646 VSS.n1660 VSS.n1658 0.0269375
R6647 VSS.n1874 VSS.n1660 0.0269375
R6648 VSS.n1027 VSS.n756 0.0269375
R6649 VSS.n756 VSS.n754 0.0269375
R6650 VSS.n754 VSS.n751 0.0269375
R6651 VSS.n751 VSS.n748 0.0269375
R6652 VSS.n748 VSS.n746 0.0269375
R6653 VSS.n746 VSS.n743 0.0269375
R6654 VSS.n743 VSS.n741 0.0269375
R6655 VSS.n741 VSS.n738 0.0269375
R6656 VSS.n738 VSS.n736 0.0269375
R6657 VSS.n736 VSS.n733 0.0269375
R6658 VSS.n733 VSS.n731 0.0269375
R6659 VSS.n731 VSS.n728 0.0269375
R6660 VSS.n728 VSS.n726 0.0269375
R6661 VSS.n726 VSS.n724 0.0269375
R6662 VSS.n724 VSS.n722 0.0269375
R6663 VSS.n722 VSS.n720 0.0269375
R6664 VSS.n720 VSS.n718 0.0269375
R6665 VSS.n718 VSS.n716 0.0269375
R6666 VSS.n716 VSS.n714 0.0269375
R6667 VSS.n714 VSS.n712 0.0269375
R6668 VSS.n712 VSS.n710 0.0269375
R6669 VSS.n710 VSS.n708 0.0269375
R6670 VSS.n708 VSS.n706 0.0269375
R6671 VSS.n706 VSS.n704 0.0269375
R6672 VSS.n704 VSS.n702 0.0269375
R6673 VSS.n702 VSS.n700 0.0269375
R6674 VSS.n700 VSS.n698 0.0269375
R6675 VSS.n698 VSS.n696 0.0269375
R6676 VSS.n696 VSS.n694 0.0269375
R6677 VSS.n694 VSS.n692 0.0269375
R6678 VSS.n692 VSS.n690 0.0269375
R6679 VSS.n690 VSS.n688 0.0269375
R6680 VSS.n688 VSS.n686 0.0269375
R6681 VSS.n686 VSS.n684 0.0269375
R6682 VSS.n684 VSS.n682 0.0269375
R6683 VSS.n682 VSS.n680 0.0269375
R6684 VSS.n680 VSS.n678 0.0269375
R6685 VSS.n678 VSS.n676 0.0269375
R6686 VSS.n676 VSS.n674 0.0269375
R6687 VSS.n674 VSS.n672 0.0269375
R6688 VSS.n672 VSS.n670 0.0269375
R6689 VSS.n670 VSS.n668 0.0269375
R6690 VSS.n668 VSS.n666 0.0269375
R6691 VSS.n666 VSS.n664 0.0269375
R6692 VSS.n664 VSS.n662 0.0269375
R6693 VSS.n662 VSS.n660 0.0269375
R6694 VSS.n660 VSS.n658 0.0269375
R6695 VSS.n658 VSS.n656 0.0269375
R6696 VSS.n656 VSS.n654 0.0269375
R6697 VSS.n654 VSS.n652 0.0269375
R6698 VSS.n652 VSS.n650 0.0269375
R6699 VSS.n650 VSS.n648 0.0269375
R6700 VSS.n648 VSS.n646 0.0269375
R6701 VSS.n646 VSS.n644 0.0269375
R6702 VSS.n644 VSS.n642 0.0269375
R6703 VSS.n642 VSS.n640 0.0269375
R6704 VSS.n640 VSS.n638 0.0269375
R6705 VSS.n1664 VSS.n1662 0.0269375
R6706 VSS.n1666 VSS.n1664 0.0269375
R6707 VSS.n1668 VSS.n1666 0.0269375
R6708 VSS.n1670 VSS.n1668 0.0269375
R6709 VSS.n1672 VSS.n1670 0.0269375
R6710 VSS.n1865 VSS.n1672 0.0269375
R6711 VSS.n929 VSS.n896 0.0269375
R6712 VSS.n896 VSS.n894 0.0269375
R6713 VSS.n894 VSS.n891 0.0269375
R6714 VSS.n891 VSS.n889 0.0269375
R6715 VSS.n889 VSS.n886 0.0269375
R6716 VSS.n886 VSS.n884 0.0269375
R6717 VSS.n884 VSS.n881 0.0269375
R6718 VSS.n881 VSS.n879 0.0269375
R6719 VSS.n879 VSS.n876 0.0269375
R6720 VSS.n876 VSS.n874 0.0269375
R6721 VSS.n874 VSS.n871 0.0269375
R6722 VSS.n871 VSS.n869 0.0269375
R6723 VSS.n869 VSS.n866 0.0269375
R6724 VSS.n866 VSS.n864 0.0269375
R6725 VSS.n864 VSS.n862 0.0269375
R6726 VSS.n862 VSS.n860 0.0269375
R6727 VSS.n860 VSS.n858 0.0269375
R6728 VSS.n858 VSS.n856 0.0269375
R6729 VSS.n856 VSS.n854 0.0269375
R6730 VSS.n854 VSS.n852 0.0269375
R6731 VSS.n852 VSS.n850 0.0269375
R6732 VSS.n850 VSS.n848 0.0269375
R6733 VSS.n848 VSS.n846 0.0269375
R6734 VSS.n846 VSS.n844 0.0269375
R6735 VSS.n844 VSS.n842 0.0269375
R6736 VSS.n842 VSS.n840 0.0269375
R6737 VSS.n840 VSS.n838 0.0269375
R6738 VSS.n838 VSS.n836 0.0269375
R6739 VSS.n836 VSS.n834 0.0269375
R6740 VSS.n834 VSS.n832 0.0269375
R6741 VSS.n832 VSS.n830 0.0269375
R6742 VSS.n830 VSS.n828 0.0269375
R6743 VSS.n828 VSS.n826 0.0269375
R6744 VSS.n826 VSS.n824 0.0269375
R6745 VSS.n824 VSS.n822 0.0269375
R6746 VSS.n822 VSS.n820 0.0269375
R6747 VSS.n820 VSS.n818 0.0269375
R6748 VSS.n818 VSS.n816 0.0269375
R6749 VSS.n816 VSS.n814 0.0269375
R6750 VSS.n814 VSS.n812 0.0269375
R6751 VSS.n812 VSS.n810 0.0269375
R6752 VSS.n810 VSS.n808 0.0269375
R6753 VSS.n808 VSS.n806 0.0269375
R6754 VSS.n806 VSS.n804 0.0269375
R6755 VSS.n804 VSS.n802 0.0269375
R6756 VSS.n802 VSS.n800 0.0269375
R6757 VSS.n800 VSS.n798 0.0269375
R6758 VSS.n798 VSS.n796 0.0269375
R6759 VSS.n796 VSS.n794 0.0269375
R6760 VSS.n794 VSS.n792 0.0269375
R6761 VSS.n792 VSS.n790 0.0269375
R6762 VSS.n790 VSS.n788 0.0269375
R6763 VSS.n788 VSS.n786 0.0269375
R6764 VSS.n786 VSS.n784 0.0269375
R6765 VSS.n784 VSS.n782 0.0269375
R6766 VSS.n782 VSS.n780 0.0269375
R6767 VSS.n780 VSS.n778 0.0269375
R6768 VSS.n1778 VSS.n1776 0.0269375
R6769 VSS.n1780 VSS.n1778 0.0269375
R6770 VSS.n1782 VSS.n1780 0.0269375
R6771 VSS.n1784 VSS.n1782 0.0269375
R6772 VSS.n1786 VSS.n1784 0.0269375
R6773 VSS.n1792 VSS.n1786 0.0269375
R6774 VSS.n2142 VSS.n2139 0.0269375
R6775 VSS.n2139 VSS.n2137 0.0269375
R6776 VSS.n2137 VSS.n2134 0.0269375
R6777 VSS.n2134 VSS.n2132 0.0269375
R6778 VSS.n2132 VSS.n2129 0.0269375
R6779 VSS.n2129 VSS.n2127 0.0269375
R6780 VSS.n2127 VSS.n2124 0.0269375
R6781 VSS.n2124 VSS.n2122 0.0269375
R6782 VSS.n2122 VSS.n2119 0.0269375
R6783 VSS.n2119 VSS.n2117 0.0269375
R6784 VSS.n2117 VSS.n2114 0.0269375
R6785 VSS.n2114 VSS.n2112 0.0269375
R6786 VSS.n2112 VSS.n2109 0.0269375
R6787 VSS.n2109 VSS.n2107 0.0269375
R6788 VSS.n2107 VSS.n2104 0.0269375
R6789 VSS.n2104 VSS.n2102 0.0269375
R6790 VSS.n2102 VSS.n2099 0.0269375
R6791 VSS.n2099 VSS.n2097 0.0269375
R6792 VSS.n2097 VSS.n2095 0.0269375
R6793 VSS.n2095 VSS.n2093 0.0269375
R6794 VSS.n2093 VSS.n2091 0.0269375
R6795 VSS.n2091 VSS.n2089 0.0269375
R6796 VSS.n2089 VSS.n2087 0.0269375
R6797 VSS.n2087 VSS.n2085 0.0269375
R6798 VSS.n2085 VSS.n2083 0.0269375
R6799 VSS.n2083 VSS.n2081 0.0269375
R6800 VSS.n2081 VSS.n2079 0.0269375
R6801 VSS.n2079 VSS.n2077 0.0269375
R6802 VSS.n2077 VSS.n2075 0.0269375
R6803 VSS.n2075 VSS.n2073 0.0269375
R6804 VSS.n2073 VSS.n2071 0.0269375
R6805 VSS.n2071 VSS.n2069 0.0269375
R6806 VSS.n2069 VSS.n2067 0.0269375
R6807 VSS.n2067 VSS.n2065 0.0269375
R6808 VSS.n2065 VSS.n2063 0.0269375
R6809 VSS.n2063 VSS.n2061 0.0269375
R6810 VSS.n2061 VSS.n2059 0.0269375
R6811 VSS.n2059 VSS.n2057 0.0269375
R6812 VSS.n2057 VSS.n2055 0.0269375
R6813 VSS.n2055 VSS.n2053 0.0269375
R6814 VSS.n2053 VSS.n2051 0.0269375
R6815 VSS.n2051 VSS.n2049 0.0269375
R6816 VSS.n2049 VSS.n2047 0.0269375
R6817 VSS.n2047 VSS.n2045 0.0269375
R6818 VSS.n2045 VSS.n2043 0.0269375
R6819 VSS.n2043 VSS.n2041 0.0269375
R6820 VSS.n2041 VSS.n2039 0.0269375
R6821 VSS.n2039 VSS.n2037 0.0269375
R6822 VSS.n2037 VSS.n2035 0.0269375
R6823 VSS.n2035 VSS.n2033 0.0269375
R6824 VSS.n2033 VSS.n2031 0.0269375
R6825 VSS.n2031 VSS.n2029 0.0269375
R6826 VSS.n2029 VSS.n2027 0.0269375
R6827 VSS.n2027 VSS.n2025 0.0269375
R6828 VSS.n2025 VSS.n2023 0.0269375
R6829 VSS.n1796 VSS.n1794 0.0269375
R6830 VSS.n1798 VSS.n1796 0.0269375
R6831 VSS.n1800 VSS.n1798 0.0269375
R6832 VSS.n1802 VSS.n1800 0.0269375
R6833 VSS.n1804 VSS.n1802 0.0269375
R6834 VSS.n1816 VSS.n1814 0.0269375
R6835 VSS.n1818 VSS.n1816 0.0269375
R6836 VSS.n1823 VSS.n1821 0.0269375
R6837 VSS.n1825 VSS.n1823 0.0269375
R6838 VSS.n1827 VSS.n1825 0.0269375
R6839 VSS.n1829 VSS.n1827 0.0269375
R6840 VSS.n1831 VSS.n1829 0.0269375
R6841 VSS.n1833 VSS.n1831 0.0269375
R6842 VSS.n1835 VSS.n1833 0.0269375
R6843 VSS.n1837 VSS.n1835 0.0269375
R6844 VSS.n1839 VSS.n1837 0.0269375
R6845 VSS.n1841 VSS.n1839 0.0269375
R6846 VSS.n1843 VSS.n1841 0.0269375
R6847 VSS.n1845 VSS.n1843 0.0269375
R6848 VSS.n1847 VSS.n1845 0.0269375
R6849 VSS.n1855 VSS.n1853 0.0269375
R6850 VSS.n1857 VSS.n1855 0.0269375
R6851 VSS.n1859 VSS.n1857 0.0269375
R6852 VSS.n1861 VSS.n1859 0.0269375
R6853 VSS.n1863 VSS.n1861 0.0269375
R6854 VSS.n1878 VSS.n1876 0.0269375
R6855 VSS.n1880 VSS.n1878 0.0269375
R6856 VSS.n1882 VSS.n1880 0.0269375
R6857 VSS.n1884 VSS.n1882 0.0269375
R6858 VSS.n1886 VSS.n1884 0.0269375
R6859 VSS.n1894 VSS.n1892 0.0269375
R6860 VSS.n1896 VSS.n1894 0.0269375
R6861 VSS.n1898 VSS.n1896 0.0269375
R6862 VSS.n1900 VSS.n1898 0.0269375
R6863 VSS.n1902 VSS.n1900 0.0269375
R6864 VSS.n1904 VSS.n1902 0.0269375
R6865 VSS.n1906 VSS.n1904 0.0269375
R6866 VSS.n1908 VSS.n1906 0.0269375
R6867 VSS.n1910 VSS.n1908 0.0269375
R6868 VSS.n1912 VSS.n1910 0.0269375
R6869 VSS.n1914 VSS.n1912 0.0269375
R6870 VSS.n1916 VSS.n1914 0.0269375
R6871 VSS.n1918 VSS.n1916 0.0269375
R6872 VSS.n1923 VSS.n1921 0.0269375
R6873 VSS.n1925 VSS.n1923 0.0269375
R6874 VSS.n1933 VSS.n1931 0.0269375
R6875 VSS.n1935 VSS.n1933 0.0269375
R6876 VSS.n1937 VSS.n1935 0.0269375
R6877 VSS.n1939 VSS.n1937 0.0269375
R6878 VSS.n1941 VSS.n1939 0.0269375
R6879 VSS.n1956 VSS.n1954 0.0269375
R6880 VSS.n1958 VSS.n1956 0.0269375
R6881 VSS.n1960 VSS.n1958 0.0269375
R6882 VSS.n1962 VSS.n1960 0.0269375
R6883 VSS.n1964 VSS.n1962 0.0269375
R6884 VSS.n1972 VSS.n1970 0.0269375
R6885 VSS.n1974 VSS.n1972 0.0269375
R6886 VSS.n1979 VSS.n1977 0.0269375
R6887 VSS.n1981 VSS.n1979 0.0269375
R6888 VSS.n1983 VSS.n1981 0.0269375
R6889 VSS.n1985 VSS.n1983 0.0269375
R6890 VSS.n1987 VSS.n1985 0.0269375
R6891 VSS.n1989 VSS.n1987 0.0269375
R6892 VSS.n1991 VSS.n1989 0.0269375
R6893 VSS.n1993 VSS.n1991 0.0269375
R6894 VSS.n1995 VSS.n1993 0.0269375
R6895 VSS.n1997 VSS.n1995 0.0269375
R6896 VSS.n1999 VSS.n1997 0.0269375
R6897 VSS.n2001 VSS.n1999 0.0269375
R6898 VSS.n2003 VSS.n2001 0.0269375
R6899 VSS.n2011 VSS.n2009 0.0269375
R6900 VSS.n2013 VSS.n2011 0.0269375
R6901 VSS.n2015 VSS.n2013 0.0269375
R6902 VSS.n2017 VSS.n2015 0.0269375
R6903 VSS.n2019 VSS.n2017 0.0269375
R6904 VSS.n935 VSS.n932 0.0269375
R6905 VSS.n938 VSS.n935 0.0269375
R6906 VSS.n941 VSS.n938 0.0269375
R6907 VSS.n944 VSS.n941 0.0269375
R6908 VSS.n947 VSS.n944 0.0269375
R6909 VSS.n958 VSS.n955 0.0269375
R6910 VSS.n961 VSS.n958 0.0269375
R6911 VSS.n964 VSS.n961 0.0269375
R6912 VSS.n967 VSS.n964 0.0269375
R6913 VSS.n970 VSS.n967 0.0269375
R6914 VSS.n973 VSS.n970 0.0269375
R6915 VSS.n976 VSS.n973 0.0269375
R6916 VSS.n979 VSS.n976 0.0269375
R6917 VSS.n982 VSS.n979 0.0269375
R6918 VSS.n985 VSS.n982 0.0269375
R6919 VSS.n988 VSS.n985 0.0269375
R6920 VSS.n991 VSS.n988 0.0269375
R6921 VSS.n994 VSS.n991 0.0269375
R6922 VSS.n997 VSS.n994 0.0269375
R6923 VSS.n1000 VSS.n997 0.0269375
R6924 VSS.n1003 VSS.n1000 0.0269375
R6925 VSS.n1014 VSS.n1011 0.0269375
R6926 VSS.n1017 VSS.n1014 0.0269375
R6927 VSS.n1020 VSS.n1017 0.0269375
R6928 VSS.n1023 VSS.n1020 0.0269375
R6929 VSS.n1026 VSS.n1023 0.0269375
R6930 VSS.n1118 VSS.n1115 0.0269375
R6931 VSS.n1121 VSS.n1118 0.0269375
R6932 VSS.n1124 VSS.n1121 0.0269375
R6933 VSS.n1127 VSS.n1124 0.0269375
R6934 VSS.n1130 VSS.n1127 0.0269375
R6935 VSS.n1141 VSS.n1138 0.0269375
R6936 VSS.n1144 VSS.n1141 0.0269375
R6937 VSS.n1147 VSS.n1144 0.0269375
R6938 VSS.n1150 VSS.n1147 0.0269375
R6939 VSS.n1153 VSS.n1150 0.0269375
R6940 VSS.n1156 VSS.n1153 0.0269375
R6941 VSS.n1159 VSS.n1156 0.0269375
R6942 VSS.n1162 VSS.n1159 0.0269375
R6943 VSS.n1165 VSS.n1162 0.0269375
R6944 VSS.n1168 VSS.n1165 0.0269375
R6945 VSS.n1171 VSS.n1168 0.0269375
R6946 VSS.n1174 VSS.n1171 0.0269375
R6947 VSS.n1177 VSS.n1174 0.0269375
R6948 VSS.n1180 VSS.n1177 0.0269375
R6949 VSS.n1183 VSS.n1180 0.0269375
R6950 VSS.n1186 VSS.n1183 0.0269375
R6951 VSS.n1197 VSS.n1194 0.0269375
R6952 VSS.n1200 VSS.n1197 0.0269375
R6953 VSS.n1203 VSS.n1200 0.0269375
R6954 VSS.n1206 VSS.n1203 0.0269375
R6955 VSS.n1209 VSS.n1206 0.0269375
R6956 VSS.n1301 VSS.n1298 0.0269375
R6957 VSS.n1304 VSS.n1301 0.0269375
R6958 VSS.n1307 VSS.n1304 0.0269375
R6959 VSS.n1310 VSS.n1307 0.0269375
R6960 VSS.n1313 VSS.n1310 0.0269375
R6961 VSS.n1324 VSS.n1321 0.0269375
R6962 VSS.n1327 VSS.n1324 0.0269375
R6963 VSS.n1330 VSS.n1327 0.0269375
R6964 VSS.n1333 VSS.n1330 0.0269375
R6965 VSS.n1336 VSS.n1333 0.0269375
R6966 VSS.n1339 VSS.n1336 0.0269375
R6967 VSS.n1342 VSS.n1339 0.0269375
R6968 VSS.n1345 VSS.n1342 0.0269375
R6969 VSS.n1348 VSS.n1345 0.0269375
R6970 VSS.n1351 VSS.n1348 0.0269375
R6971 VSS.n1354 VSS.n1351 0.0269375
R6972 VSS.n1357 VSS.n1354 0.0269375
R6973 VSS.n1360 VSS.n1357 0.0269375
R6974 VSS.n1363 VSS.n1360 0.0269375
R6975 VSS.n1366 VSS.n1363 0.0269375
R6976 VSS.n1369 VSS.n1366 0.0269375
R6977 VSS.n1380 VSS.n1377 0.0269375
R6978 VSS.n1383 VSS.n1380 0.0269375
R6979 VSS.n1386 VSS.n1383 0.0269375
R6980 VSS.n1389 VSS.n1386 0.0269375
R6981 VSS.n1392 VSS.n1389 0.0269375
R6982 VSS.n2982 VSS.n2981 0.0266563
R6983 VSS.n2990 VSS.n2989 0.0260938
R6984 VSS.n16 VSS.n15 0.0258125
R6985 VSS.n3272 VSS.n3269 0.0255312
R6986 VSS.n2935 VSS.n2933 0.0246875
R6987 VSS.n235 VSS.n228 0.0246875
R6988 VSS.n3316 VSS.n3007 0.0244062
R6989 VSS.n2963 VSS.n2961 0.0244062
R6990 VSS.n3132 VSS.n3123 0.0244062
R6991 VSS.n2725 VSS.n2724 0.0244062
R6992 VSS.n2594 VSS.n2587 0.024125
R6993 VSS.n2958 VSS.n2861 0.024125
R6994 VSS.n359 VSS.n242 0.024125
R6995 VSS.n1819 VSS.n1818 0.024125
R6996 VSS.n1921 VSS.n1919 0.024125
R6997 VSS.n1975 VSS.n1974 0.024125
R6998 VSS.n2745 VSS.n2743 0.0238437
R6999 VSS.n2797 VSS.n2795 0.0238437
R7000 VSS.n2838 VSS.n2837 0.0238437
R7001 VSS.n3155 VSS.n3152 0.0238437
R7002 VSS.n3231 VSS.n3228 0.0238437
R7003 VSS.n3294 VSS.n3293 0.0238437
R7004 VSS.n1811 VSS.n1809 0.0235625
R7005 VSS.n1851 VSS.n1850 0.0235625
R7006 VSS.n1889 VSS.n1887 0.0235625
R7007 VSS.n1929 VSS.n1928 0.0235625
R7008 VSS.n1967 VSS.n1965 0.0235625
R7009 VSS.n2007 VSS.n2006 0.0235625
R7010 VSS.n951 VSS.n948 0.0235625
R7011 VSS.n1008 VSS.n1007 0.0235625
R7012 VSS.n1134 VSS.n1131 0.0235625
R7013 VSS.n1191 VSS.n1190 0.0235625
R7014 VSS.n1317 VSS.n1314 0.0235625
R7015 VSS.n1374 VSS.n1373 0.0235625
R7016 VSS.n2642 VSS.n2637 0.023
R7017 VSS.n1812 VSS.n1811 0.0224375
R7018 VSS.n1850 VSS.n1848 0.0224375
R7019 VSS.n1890 VSS.n1889 0.0224375
R7020 VSS.n1928 VSS.n1926 0.0224375
R7021 VSS.n1968 VSS.n1967 0.0224375
R7022 VSS.n2006 VSS.n2004 0.0224375
R7023 VSS.n952 VSS.n951 0.0224375
R7024 VSS.n1007 VSS.n1004 0.0224375
R7025 VSS.n1135 VSS.n1134 0.0224375
R7026 VSS.n1190 VSS.n1187 0.0224375
R7027 VSS.n1318 VSS.n1317 0.0224375
R7028 VSS.n1373 VSS.n1370 0.0224375
R7029 VSS.n2763 VSS.n2762 0.0221563
R7030 VSS.n3181 VSS.n3180 0.0221563
R7031 VSS.n2892 VSS.n2891 0.0213125
R7032 VSS.n3861 VSS.n3860 0.0213125
R7033 VSS.n3420 VSS.n3419 0.0213125
R7034 VSS.n2437 VSS.n2434 0.0213125
R7035 VSS.n13 VSS.n11 0.0213125
R7036 VSS.n59 VSS.n58 0.0213125
R7037 VSS.n2699 VSS.n2698 0.0210419
R7038 VSS.n2679 VSS.n2678 0.0210419
R7039 VSS.n3817 VSS.n3816 0.02075
R7040 VSS.n3331 VSS.n2662 0.019625
R7041 VSS.n2511 VSS.n2510 0.019625
R7042 VSS.n52 VSS.n50 0.019625
R7043 VSS.n3383 VSS.n2465 0.0195
R7044 VSS.n2780 VSS.n2778 0.0193437
R7045 VSS.n3206 VSS.n3203 0.0193437
R7046 VSS.n3283 VSS.n3280 0.0193437
R7047 VSS.n3949 VSS.n3944 0.0190625
R7048 VSS.n3941 VSS.n3938 0.0190625
R7049 VSS.n2953 VSS.n2952 0.0190625
R7050 VSS.n2950 VSS.n2948 0.0190625
R7051 VSS.n3881 VSS.n3879 0.0190625
R7052 VSS.n3884 VSS.n3883 0.0190625
R7053 VSS.n2604 VSS.n2601 0.0190625
R7054 VSS.n2608 VSS.n2607 0.0190625
R7055 VSS.n3273 VSS.n3272 0.0182187
R7056 VSS.n2752 VSS.n2750 0.0176563
R7057 VSS.n2831 VSS.n2830 0.0176563
R7058 VSS.n3165 VSS.n3162 0.0176563
R7059 VSS.n3284 VSS.n3283 0.0176563
R7060 VSS.n2992 VSS.n2990 0.0170938
R7061 VSS.n1695 VSS.n1694 0.0167343
R7062 VSS.n1715 VSS.n1714 0.0167343
R7063 VSS.n1759 VSS.n1758 0.0167343
R7064 VSS.n1750 VSS.n1749 0.0167343
R7065 VSS.n1735 VSS.n1734 0.0167343
R7066 VSS.n1565 VSS.n1564 0.0167343
R7067 VSS.n1629 VSS.n1628 0.0167343
R7068 VSS.n1620 VSS.n1619 0.0167343
R7069 VSS.n1605 VSS.n1604 0.0167343
R7070 VSS.n1585 VSS.n1584 0.0167343
R7071 VSS.n1435 VSS.n1434 0.0167343
R7072 VSS.n1455 VSS.n1454 0.0167343
R7073 VSS.n1499 VSS.n1498 0.0167343
R7074 VSS.n1490 VSS.n1489 0.0167343
R7075 VSS.n1475 VSS.n1474 0.0167343
R7076 VSS.n2984 VSS.n2982 0.0165313
R7077 VSS.n336 VSS.n334 0.01625
R7078 VSS.n327 VSS.n326 0.01625
R7079 VSS.n4083 VSS.n4080 0.01625
R7080 VSS.n4070 VSS.n4069 0.01625
R7081 VSS.n2169 VSS.n2143 0.01625
R7082 VSS.n1792 VSS.n1791 0.01625
R7083 VSS.n1869 VSS.n1865 0.01625
R7084 VSS.n1874 VSS.n1872 0.01625
R7085 VSS.n1947 VSS.n1943 0.01625
R7086 VSS.n1952 VSS.n1950 0.01625
R7087 VSS.n929 VSS.n928 0.01625
R7088 VSS.n1059 VSS.n1027 0.01625
R7089 VSS.n1112 VSS.n1111 0.01625
R7090 VSS.n1242 VSS.n1210 0.01625
R7091 VSS.n1295 VSS.n1294 0.01625
R7092 VSS.n1398 VSS.n1397 0.01625
R7093 VSS.n2808 VSS.n2807 0.0159688
R7094 VSS.n3247 VSS.n3246 0.0159688
R7095 VSS.n4063 VSS.n4060 0.0153235
R7096 VSS.n3769 VSS.n3753 0.0153235
R7097 VSS.n2462 VSS.n2461 0.0145
R7098 VSS.n2990 VSS.n2668 0.0142813
R7099 VSS.n2982 VSS.n2674 0.0142813
R7100 VSS.n2725 VSS.n2715 0.0142813
R7101 VSS.n2961 VSS.n2960 0.0142813
R7102 VSS.n3132 VSS.n3131 0.0142813
R7103 VSS.n3326 VSS.n3316 0.0142813
R7104 VSS.n3381 VSS.n3380 0.0140074
R7105 VSS.n2212 VSS.n2210 0.014
R7106 VSS.n4058 VSS.n4057 0.0139933
R7107 VSS.n2938 VSS.n2937 0.0134375
R7108 VSS.n2143 VSS.n2142 0.0134375
R7109 VSS.n2727 VSS.n2725 0.0131563
R7110 VSS.n2961 VSS.n2852 0.0131563
R7111 VSS.n3134 VSS.n3132 0.0131563
R7112 VSS.n3316 VSS.n3315 0.0131563
R7113 VSS.n3333 VSS.n3331 0.012875
R7114 VSS.n2315 VSS.n2313 0.01175
R7115 VSS.n2417 VSS.n2398 0.01175
R7116 VSS.n300 VSS.n299 0.01175
R7117 VSS.n3732 VSS.n3730 0.01175
R7118 VSS.n2214 VSS.n2212 0.01175
R7119 VSS VSS.n2297 0.01175
R7120 VSS.n2810 VSS.n2808 0.0114688
R7121 VSS.n3250 VSS.n3247 0.0114688
R7122 VSS.n2883 VSS.n2881 0.0111875
R7123 VSS.n3852 VSS.n3850 0.0111875
R7124 VSS.n1794 VSS.n1792 0.0111875
R7125 VSS.n1865 VSS.n1863 0.0111875
R7126 VSS.n1876 VSS.n1874 0.0111875
R7127 VSS.n1943 VSS.n1941 0.0111875
R7128 VSS.n1954 VSS.n1952 0.0111875
R7129 VSS.n2023 VSS.n2019 0.0111875
R7130 VSS.n932 VSS.n929 0.0111875
R7131 VSS.n1027 VSS.n1026 0.0111875
R7132 VSS.n1115 VSS.n1112 0.0111875
R7133 VSS.n1210 VSS.n1209 0.0111875
R7134 VSS.n1298 VSS.n1295 0.0111875
R7135 VSS.n1398 VSS.n1392 0.0111875
R7136 VSS.n2750 VSS.n2749 0.00978125
R7137 VSS.n2833 VSS.n2831 0.00978125
R7138 VSS.n3162 VSS.n3161 0.00978125
R7139 VSS.n3287 VSS.n3284 0.00978125
R7140 VSS.n2645 VSS.n2642 0.0095
R7141 VSS.n350 VSS.n349 0.0095
R7142 VSS.n313 VSS.n311 0.0095
R7143 VSS.n3746 VSS.n3743 0.0095
R7144 VSS.n4103 VSS.n4102 0.0095
R7145 VSS.n3276 VSS.n3273 0.00921875
R7146 VSS.n2930 VSS.n2928 0.0089375
R7147 VSS.n2631 VSS.n2629 0.008375
R7148 VSS.n3931 VSS.n3927 0.008375
R7149 VSS.n3892 VSS.n3890 0.008375
R7150 VSS.n3970 VSS.n3968 0.008375
R7151 VSS.n2210 VSS.n2209 0.008375
R7152 VSS.n2778 VSS.n2777 0.00809375
R7153 VSS.n3203 VSS.n3202 0.00809375
R7154 VSS.n3280 VSS.n3279 0.00809375
R7155 VSS.n237 VSS.n235 0.0078125
R7156 VSS.n2925 VSS.n2924 0.0078125
R7157 VSS.n35 VSS.n34 0.0078125
R7158 VSS.n359 VSS.n358 0.00725
R7159 VSS.n355 VSS.n353 0.00725
R7160 VSS.n305 VSS.n304 0.00725
R7161 VSS.n3739 VSS.n3738 0.00725
R7162 VSS.n4110 VSS.n4107 0.00725
R7163 VSS.n2177 VSS.n2176 0.00725
R7164 VSS.n235 VSS.n234 0.00725
R7165 VSS.n343 VSS.n342 0.006125
R7166 VSS.n320 VSS.n318 0.006125
R7167 VSS.n4093 VSS.n4092 0.006125
R7168 VSS.n3772 VSS.n3769 0.00579412
R7169 VSS.n3427 VSS.n3426 0.0055625
R7170 VSS.n2424 VSS.n2421 0.0055625
R7171 VSS.n8 VSS.n6 0.0055625
R7172 VSS.n64 VSS.n63 0.0055625
R7173 VSS.n2765 VSS.n2763 0.00528125
R7174 VSS.n3184 VSS.n3181 0.00528125
R7175 VSS.n3824 VSS.n3823 0.005
R7176 VSS.n1814 VSS.n1812 0.005
R7177 VSS.n1848 VSS.n1847 0.005
R7178 VSS.n1892 VSS.n1890 0.005
R7179 VSS.n1926 VSS.n1925 0.005
R7180 VSS.n1970 VSS.n1968 0.005
R7181 VSS.n2004 VSS.n2003 0.005
R7182 VSS.n955 VSS.n952 0.005
R7183 VSS.n1004 VSS.n1003 0.005
R7184 VSS.n1138 VSS.n1135 0.005
R7185 VSS.n1187 VSS.n1186 0.005
R7186 VSS.n1321 VSS.n1318 0.005
R7187 VSS.n1370 VSS.n1369 0.005
R7188 VSS.n2518 VSS.n2517 0.003875
R7189 VSS.n1809 VSS.n1804 0.003875
R7190 VSS.n1853 VSS.n1851 0.003875
R7191 VSS.n1887 VSS.n1886 0.003875
R7192 VSS.n1931 VSS.n1929 0.003875
R7193 VSS.n1965 VSS.n1964 0.003875
R7194 VSS.n2009 VSS.n2007 0.003875
R7195 VSS.n948 VSS.n947 0.003875
R7196 VSS.n1011 VSS.n1008 0.003875
R7197 VSS.n1131 VSS.n1130 0.003875
R7198 VSS.n1194 VSS.n1191 0.003875
R7199 VSS.n1314 VSS.n1313 0.003875
R7200 VSS.n1377 VSS.n1374 0.003875
R7201 VSS.n2743 VSS.n2742 0.00359375
R7202 VSS.n2795 VSS.n2794 0.00359375
R7203 VSS.n2840 VSS.n2838 0.00359375
R7204 VSS.n3152 VSS.n3151 0.00359375
R7205 VSS.n3228 VSS.n3227 0.00359375
R7206 VSS.n3297 VSS.n3294 0.00359375
R7207 VSS.n2143 VSS.n1411 0.0033125
R7208 VSS.n2943 VSS.n2941 0.0033125
R7209 VSS.n1821 VSS.n1819 0.0033125
R7210 VSS.n1919 VSS.n1918 0.0033125
R7211 VSS.n1977 VSS.n1975 0.0033125
R7212 VSS.n3380 VSS.n3370 0.00275
R7213 VSS.n4057 VSS.n4044 0.00275
R7214 VSS.n3269 VSS.n3268 0.00190625
R7215 VSS.n3872 VSS.n3870 0.0010625
R7216 VDD.t237 VDD.t329 147.304
R7217 VDD.t164 VDD.t237 147.304
R7218 VDD.t207 VDD.t164 147.304
R7219 VDD.t395 VDD.t207 147.304
R7220 VDD.t343 VDD.t389 147.304
R7221 VDD.t267 VDD.t343 147.304
R7222 VDD.t387 VDD.t267 147.304
R7223 VDD.t339 VDD.t387 147.304
R7224 VDD.t375 VDD.t371 135.05
R7225 VDD.t393 VDD.t375 135.05
R7226 VDD.t222 VDD.t337 135.05
R7227 VDD.t279 VDD.t222 135.05
R7228 VDD.t345 VDD.t313 135.05
R7229 VDD.t373 VDD.t345 135.05
R7230 VDD.t181 VDD.t175 135.05
R7231 VDD.t210 VDD.t181 135.05
R7232 VDD.t251 VDD.t155 118.626
R7233 VDD.t391 VDD.t326 118.626
R7234 VDD.n7971 VDD.t185 103.504
R7235 VDD.n6625 VDD.t393 74.5648
R7236 VDD.n547 VDD.t279 74.5648
R7237 VDD.n555 VDD.t373 74.5648
R7238 VDD.n1028 VDD.t210 74.5648
R7239 VDD.n305 VDD.t395 72.6094
R7240 VDD.n305 VDD.t349 72.6094
R7241 VDD.n6860 VDD.t339 72.6094
R7242 VDD.n6860 VDD.t264 72.6094
R7243 VDD.n5623 VDD.t288 68.0469
R7244 VDD.n5623 VDD.t320 68.0469
R7245 VDD.n4238 VDD.t316 68.0469
R7246 VDD.n4238 VDD.t335 68.0469
R7247 VDD.n5573 VDD.t230 68.0469
R7248 VDD.n4179 VDD.t363 68.0469
R7249 VDD.n4179 VDD.t333 68.0469
R7250 VDD.n5573 VDD.t284 68.0469
R7251 VDD.n5539 VDD.t361 68.0469
R7252 VDD.n3947 VDD.t277 68.0469
R7253 VDD.n3947 VDD.t225 68.0469
R7254 VDD.n5539 VDD.t379 68.0469
R7255 VDD.n5489 VDD.t331 68.0469
R7256 VDD.n3887 VDD.t309 68.0469
R7257 VDD.n3887 VDD.t253 68.0469
R7258 VDD.n5489 VDD.t353 68.0469
R7259 VDD.n2667 VDD.t244 68.0469
R7260 VDD.n2830 VDD.t324 68.0469
R7261 VDD.n2830 VDD.t291 68.0469
R7262 VDD.n2667 VDD.t299 68.0469
R7263 VDD.n6216 VDD.t233 68.0469
R7264 VDD.n2898 VDD.t247 68.0469
R7265 VDD.n2898 VDD.t212 68.0469
R7266 VDD.n6216 VDD.t286 68.0469
R7267 VDD.n6039 VDD.t256 68.0469
R7268 VDD.n3387 VDD.t385 68.0469
R7269 VDD.n3387 VDD.t367 68.0469
R7270 VDD.n6039 VDD.t311 68.0469
R7271 VDD.n5393 VDD.t239 68.0469
R7272 VDD.n5393 VDD.t293 68.0469
R7273 VDD.n3446 VDD.t318 68.0469
R7274 VDD.n3446 VDD.t341 68.0469
R7275 VDD.n5420 VDD.t140 68.0469
R7276 VDD.n5420 VDD.t187 68.0469
R7277 VDD.n3700 VDD.t242 68.0469
R7278 VDD.n3700 VDD.t295 68.0469
R7279 VDD.n5470 VDD.t249 68.0469
R7280 VDD.n5470 VDD.t305 68.0469
R7281 VDD.n3760 VDD.t146 68.0469
R7282 VDD.n3760 VDD.t189 68.0469
R7283 VDD.n6160 VDD.t149 68.0469
R7284 VDD.n6160 VDD.t191 68.0469
R7285 VDD.n2957 VDD.t220 68.0469
R7286 VDD.n2957 VDD.t259 68.0469
R7287 VDD.n5283 VDD.t322 68.0469
R7288 VDD.n5283 VDD.t347 68.0469
R7289 VDD.n3196 VDD.t167 68.0469
R7290 VDD.n3196 VDD.t197 68.0469
R7291 VDD.n5333 VDD.t158 68.0469
R7292 VDD.n5333 VDD.t193 68.0469
R7293 VDD.n3256 VDD.t355 68.0469
R7294 VDD.n3256 VDD.t377 68.0469
R7295 VDD.n2580 VDD.t173 68.0469
R7296 VDD.n2580 VDD.t199 68.0469
R7297 VDD.n2889 VDD.t381 68.0469
R7298 VDD.n2889 VDD.t143 68.0469
R7299 VDD.n391 VDD.t391 63.8344
R7300 VDD.n402 VDD.t204 63.8344
R7301 VDD.n7904 VDD.t152 62.6612
R7302 VDD.n7969 VDD.t170 62.6612
R7303 VDD.n318 VDD.t281 62.4005
R7304 VDD.n315 VDD.t261 62.4005
R7305 VDD.n7971 VDD.t251 58.6612
R7306 VDD.n6625 VDD.t161 58.4005
R7307 VDD.n547 VDD.t307 58.4005
R7308 VDD.n555 VDD.t383 58.4005
R7309 VDD.n1028 VDD.t235 58.4005
R7310 VDD.t201 VDD.t369 49.6666
R7311 VDD.t215 VDD.t201 49.6666
R7312 VDD.t359 VDD.t228 49.6666
R7313 VDD.t365 VDD.t359 49.6666
R7314 VDD.n1447 VDD.t270 46.9291
R7315 VDD.n1125 VDD.t297 46.9291
R7316 VDD.n1125 VDD.t351 46.9291
R7317 VDD.n1447 VDD.t273 46.9291
R7318 VDD.n1439 VDD.t301 46.9291
R7319 VDD.n1439 VDD.t303 46.9291
R7320 VDD.n1345 VDD.t178 46.9291
R7321 VDD.n1099 VDD.t195 46.9291
R7322 VDD.n1099 VDD.t275 46.9291
R7323 VDD.n1345 VDD.t183 46.9291
R7324 VDD.n7887 VDD.t215 24.8335
R7325 VDD.n7887 VDD.t357 24.8335
R7326 VDD.n6 VDD.t365 24.8335
R7327 VDD.n6 VDD.t217 24.8335
R7328 VDD.n374 VDD.t940 13.6237
R7329 VDD.n144 VDD.t268 12.939
R7330 VDD.n203 VDD.t165 12.939
R7331 VDD.t568 VDD.t61 12.7541
R7332 VDD.n7020 VDD.n7019 12.7307
R7333 VDD.n8328 VDD.t26 12.7307
R7334 VDD.n7913 VDD.t572 12.4643
R7335 VDD.n7948 VDD.t564 12.4643
R7336 VDD.n157 VDD.t458 12.3639
R7337 VDD.n190 VDD.t470 12.3639
R7338 VDD.n6987 VDD.t265 12.189
R7339 VDD.n7049 VDD.t208 12.189
R7340 VDD.n371 VDD.t565 11.8846
R7341 VDD.n7000 VDD.t457 11.6473
R7342 VDD.n7035 VDD.t501 11.6473
R7343 VDD.n7938 VDD.t507 11.3048
R7344 VDD.n358 VDD.t464 10.7251
R7345 VDD.n355 VDD.t91 10.7251
R7346 VDD.n7200 VDD.t4 10.5639
R7347 VDD.n8346 VDD.t23 10.0222
R7348 VDD.n1086 VDD.t176 9.91676
R7349 VDD.n785 VDD.t314 9.91676
R7350 VDD.n7929 VDD.t566 9.56572
R7351 VDD.n7932 VDD.t571 9.56572
R7352 VDD.n172 VDD.t499 9.48871
R7353 VDD.n175 VDD.t468 9.48871
R7354 VDD.n1073 VDD.t961 9.47604
R7355 VDD.n773 VDD.t970 9.47604
R7356 VDD.n2480 VDD.t75 9.23695
R7357 VDD.n7016 VDD.t459 8.93874
R7358 VDD.n7020 VDD.t498 8.93874
R7359 VDD.n2110 VDD.t411 8.82644
R7360 VDD.n2421 VDD.t135 8.82644
R7361 VDD.n828 VDD.t575 8.59459
R7362 VDD.n849 VDD.t578 8.59459
R7363 VDD.n4418 VDD.t900 8.54751
R7364 VDD.n4438 VDD.t1100 8.54751
R7365 VDD.n4889 VDD.t1053 8.54751
R7366 VDD.n4909 VDD.t1022 8.54751
R7367 VDD.n5036 VDD.t1059 8.54751
R7368 VDD.n5056 VDD.t746 8.54751
R7369 VDD.n4587 VDD.t632 8.54751
R7370 VDD.n4607 VDD.t1201 8.54751
R7371 VDD.n4734 VDD.t822 8.54751
R7372 VDD.n4754 VDD.t770 8.54751
R7373 VDD.n5191 VDD.t776 8.54751
R7374 VDD.n5211 VDD.t895 8.54751
R7375 VDD.n6513 VDD.t671 8.54751
R7376 VDD.n6533 VDD.t668 8.54751
R7377 VDD.n2101 VDD.t66 8.41594
R7378 VDD.n2441 VDD.t78 8.41594
R7379 VDD.n331 VDD.t327 8.4063
R7380 VDD.n7916 VDD.t433 8.4063
R7381 VDD.n8132 VDD.t156 8.4063
R7382 VDD.n2092 VDD.t139 8.00543
R7383 VDD.n2202 VDD.t33 8.00543
R7384 VDD.n7221 VDD.t15 7.85532
R7385 VDD.n2083 VDD.t412 7.59492
R7386 VDD.n2211 VDD.t54 7.59492
R7387 VDD.n2295 VDD.t491 7.59492
R7388 VDD.n7209 VDD.t7 7.31361
R7389 VDD.n1056 VDD.t943 7.27243
R7390 VDD.n756 VDD.t951 7.27243
R7391 VDD.n837 VDD.t574 7.27243
R7392 VDD.n840 VDD.t583 7.27243
R7393 VDD.n374 VDD.t562 7.24688
R7394 VDD.n2175 VDD.t115 7.18441
R7395 VDD.n2283 VDD.t488 7.18441
R7396 VDD.n2463 VDD.t93 7.18441
R7397 VDD.n1456 VDD.t431 7.0395
R7398 VDD.n1455 VDD.t494 7.0395
R7399 VDD.n1928 VDD.t475 7.0395
R7400 VDD.n1929 VDD.t493 7.0395
R7401 VDD.n4398 VDD.t615 6.91951
R7402 VDD.n4458 VDD.t759 6.91951
R7403 VDD.n4869 VDD.t765 6.91951
R7404 VDD.n4929 VDD.t685 6.91951
R7405 VDD.n5016 VDD.t1044 6.91951
R7406 VDD.n5076 VDD.t762 6.91951
R7407 VDD.n4567 VDD.t1098 6.91951
R7408 VDD.n4627 VDD.t882 6.91951
R7409 VDD.n4714 VDD.t1016 6.91951
R7410 VDD.n4774 VDD.t626 6.91951
R7411 VDD.n5171 VDD.t678 6.91951
R7412 VDD.n5231 VDD.t695 6.91951
R7413 VDD.n6493 VDD.t1205 6.91951
R7414 VDD.n6553 VDD.t594 6.91951
R7415 VDD.n7732 VDD.t479 6.87803
R7416 VDD.n7710 VDD.t585 6.87803
R7417 VDD.n7697 VDD.t586 6.87803
R7418 VDD.n7689 VDD.t41 6.87803
R7419 VDD.n7673 VDD.t42 6.87803
R7420 VDD.n7629 VDD.t59 6.87803
R7421 VDD.n7613 VDD.t60 6.87803
R7422 VDD.n7605 VDD.t489 6.87803
R7423 VDD.n7592 VDD.t490 6.87803
R7424 VDD.n7570 VDD.t415 6.87803
R7425 VDD.n7719 VDD.t480 6.87615
R7426 VDD.n7583 VDD.t414 6.87615
R7427 VDD.n7886 VDD.t502 6.83706
R7428 VDD.n7808 VDD.t35 6.83492
R7429 VDD.n7478 VDD.t43 6.83492
R7430 VDD.n7271 VDD.t46 6.82906
R7431 VDD.n7257 VDD.t45 6.82906
R7432 VDD.n7249 VDD.t503 6.82906
R7433 VDD.n7841 VDD.t65 6.82906
R7434 VDD.n7826 VDD.t64 6.82906
R7435 VDD.n7333 VDD.t497 6.82906
R7436 VDD.n7340 VDD.t496 6.82906
R7437 VDD.n7349 VDD.t37 6.82906
R7438 VDD.n7362 VDD.t36 6.82906
R7439 VDD.n7369 VDD.t443 6.82906
R7440 VDD.n7382 VDD.t442 6.82906
R7441 VDD.n2190 VDD.t413 6.7739
R7442 VDD.n2274 VDD.t410 6.7739
R7443 VDD.n2400 VDD.t446 6.7739
R7444 VDD.n2403 VDD.t428 6.7739
R7445 VDD.n7916 VDD.t569 6.66717
R7446 VDD.n160 VDD.t463 6.6135
R7447 VDD.n187 VDD.t469 6.6135
R7448 VDD.n4402 VDD.t1030 6.51251
R7449 VDD.n4454 VDD.t914 6.51251
R7450 VDD.n4873 VDD.t740 6.51251
R7451 VDD.n4925 VDD.t1035 6.51251
R7452 VDD.n5020 VDD.t817 6.51251
R7453 VDD.n5072 VDD.t870 6.51251
R7454 VDD.n4571 VDD.t1048 6.51251
R7455 VDD.n4623 VDD.t813 6.51251
R7456 VDD.n4718 VDD.t612 6.51251
R7457 VDD.n4770 VDD.t791 6.51251
R7458 VDD.n5175 VDD.t835 6.51251
R7459 VDD.n5227 VDD.t815 6.51251
R7460 VDD.n6497 VDD.t844 6.51251
R7461 VDD.n6549 VDD.t701 6.51251
R7462 VDD.n1795 VDD.t116 6.4095
R7463 VDD.n1794 VDD.t117 6.4095
R7464 VDD.n1793 VDD.t513 6.4095
R7465 VDD.n1544 VDD.t514 6.4095
R7466 VDD.n1456 VDD.t432 6.4095
R7467 VDD.n1455 VDD.t495 6.4095
R7468 VDD.n1792 VDD.t87 6.4095
R7469 VDD.n1791 VDD.t88 6.4095
R7470 VDD.n1790 VDD.t484 6.4095
R7471 VDD.n1454 VDD.t485 6.4095
R7472 VDD.n1928 VDD.t474 6.4095
R7473 VDD.n1929 VDD.t492 6.4095
R7474 VDD.n2459 VDD.t106 6.36339
R7475 VDD.n393 VDD.t328 6.2405
R7476 VDD.n7980 VDD.t157 6.2405
R7477 VDD.n7004 VDD.t456 6.23019
R7478 VDD.n7032 VDD.t462 6.23019
R7479 VDD.n7802 VDD.t114 6.21361
R7480 VDD.n7487 VDD.t34 6.21361
R7481 VDD.n2122 VDD.t473 5.95288
R7482 VDD.t481 VDD.t567 5.7976
R7483 VDD.n331 VDD.t282 5.50775
R7484 VDD.n387 VDD.t119 5.50775
R7485 VDD.n371 VDD.t471 5.50775
R7486 VDD.n367 VDD.t938 5.50775
R7487 VDD.n7929 VDD.t587 5.50775
R7488 VDD.n8334 VDD.t11 5.14676
R7489 VDD.n8311 VDD.t202 5.14676
R7490 VDD.n2446 VDD.t72 5.13186
R7491 VDD.n1069 VDD.t948 5.06881
R7492 VDD.n769 VDD.t963 5.06881
R7493 VDD.n803 VDD.t223 5.06881
R7494 VDD.n6637 VDD.t162 5.06881
R7495 VDD.n4415 VDD.t698 4.88451
R7496 VDD.n4441 VDD.t676 4.88451
R7497 VDD.n4886 VDD.t620 4.88451
R7498 VDD.n4912 VDD.t607 4.88451
R7499 VDD.n5033 VDD.t922 4.88451
R7500 VDD.n5059 VDD.t838 4.88451
R7501 VDD.n4584 VDD.t623 4.88451
R7502 VDD.n4610 VDD.t885 4.88451
R7503 VDD.n4731 VDD.t1012 4.88451
R7504 VDD.n4757 VDD.t693 4.88451
R7505 VDD.n5188 VDD.t929 4.88451
R7506 VDD.n5214 VDD.t666 4.88451
R7507 VDD.n6510 VDD.t778 4.88451
R7508 VDD.n6536 VDD.t710 4.88451
R7509 VDD.n2386 VDD.t519 4.72135
R7510 VDD.n2417 VDD.t398 4.72135
R7511 VDD.n7466 VDD.t0 4.66033
R7512 VDD.n1436 VDD.n1435 4.64717
R7513 VDD.n4385 VDD.t664 4.4775
R7514 VDD.n4471 VDD.t602 4.4775
R7515 VDD.n4856 VDD.t1119 4.4775
R7516 VDD.n4942 VDD.t919 4.4775
R7517 VDD.n5003 VDD.t1094 4.4775
R7518 VDD.n5089 VDD.t609 4.4775
R7519 VDD.n4554 VDD.t1005 4.4775
R7520 VDD.n4640 VDD.t673 4.4775
R7521 VDD.n4701 VDD.t831 4.4775
R7522 VDD.n4787 VDD.t800 4.4775
R7523 VDD.n5158 VDD.t1051 4.4775
R7524 VDD.n5244 VDD.t794 4.4775
R7525 VDD.n6480 VDD.t605 4.4775
R7526 VDD.n6566 VDD.t688 4.4775
R7527 VDD.n338 VDD.t580 4.34833
R7528 VDD.n342 VDD.t205 4.34833
R7529 VDD.n348 VDD.t481 4.34833
R7530 VDD.n358 VDD.t570 4.34833
R7531 VDD.n7955 VDD.t171 4.34833
R7532 VDD.n7966 VDD.n7965 4.31441
R7533 VDD.n2476 VDD.t80 4.31084
R7534 VDD.n400 VDD.n399 4.09528
R7535 VDD.n8159 VDD.n8156 4.09137
R7536 VDD.n8148 VDD.n8145 4.09137
R7537 VDD.n7897 VDD.n7894 4.09137
R7538 VDD.n1362 VDD.n1361 4.0405
R7539 VDD.n1373 VDD.n1372 4.0405
R7540 VDD.n1384 VDD.n1383 4.0405
R7541 VDD.n1395 VDD.n1394 4.0405
R7542 VDD.n1406 VDD.n1405 4.0405
R7543 VDD.n1417 VDD.n1416 4.0405
R7544 VDD.n7419 VDD.t49 4.03902
R7545 VDD.n7498 VDD.t118 4.03902
R7546 VDD.n557 VDD.t384 4.02914
R7547 VDD.n5574 VDD.n5573 4.0005
R7548 VDD.n4180 VDD.n4179 4.0005
R7549 VDD.n5540 VDD.n5539 4.0005
R7550 VDD.n3948 VDD.n3947 4.0005
R7551 VDD.n5490 VDD.n5489 4.0005
R7552 VDD.n3888 VDD.n3887 4.0005
R7553 VDD.n3447 VDD.n3446 4.0005
R7554 VDD.n5394 VDD.n5393 4.0005
R7555 VDD.n3701 VDD.n3700 4.0005
R7556 VDD.n5421 VDD.n5420 4.0005
R7557 VDD.n3761 VDD.n3760 4.0005
R7558 VDD.n5471 VDD.n5470 4.0005
R7559 VDD.n6040 VDD.n6039 4.0005
R7560 VDD.n3388 VDD.n3387 4.0005
R7561 VDD.n2958 VDD.n2957 4.0005
R7562 VDD.n6161 VDD.n6160 4.0005
R7563 VDD.n3197 VDD.n3196 4.0005
R7564 VDD.n5284 VDD.n5283 4.0005
R7565 VDD.n3257 VDD.n3256 4.0005
R7566 VDD.n5334 VDD.n5333 4.0005
R7567 VDD.n6217 VDD.n6216 4.0005
R7568 VDD.n2899 VDD.n2898 4.0005
R7569 VDD.n2890 VDD.n2889 4.0005
R7570 VDD.n2581 VDD.n2580 4.0005
R7571 VDD.n2668 VDD.n2667 4.0005
R7572 VDD.n2831 VDD.n2830 4.0005
R7573 VDD.n548 VDD.n547 4.0005
R7574 VDD.n556 VDD.n555 4.0005
R7575 VDD.n1029 VDD.n1028 4.0005
R7576 VDD.n6626 VDD.n6625 4.0005
R7577 VDD.n306 VDD.n305 4.0005
R7578 VDD.n6861 VDD.n6860 4.0005
R7579 VDD.n7 VDD.n6 4.0005
R7580 VDD.n7888 VDD.n7887 4.0005
R7581 VDD.n7972 VDD.n7971 4.0005
R7582 VDD.n1448 VDD.n1447 4.0005
R7583 VDD.n1126 VDD.n1125 4.0005
R7584 VDD.n1440 VDD.n1439 4.0005
R7585 VDD.n1346 VDD.n1345 4.0005
R7586 VDD.n1100 VDD.n1099 4.0005
R7587 VDD.n4239 VDD.n4238 4.0005
R7588 VDD.n5624 VDD.n5623 4.0005
R7589 VDD.n403 VDD.t206 3.9242
R7590 VDD.n7905 VDD.t154 3.90659
R7591 VDD.n7970 VDD.t172 3.90659
R7592 VDD.n5598 VDD.n5597 3.89963
R7593 VDD.n4202 VDD.n4201 3.89963
R7594 VDD.n4211 VDD.n4210 3.89963
R7595 VDD.n5520 VDD.n5519 3.89963
R7596 VDD.n3920 VDD.n3919 3.89963
R7597 VDD.n3929 VDD.n3928 3.89963
R7598 VDD.n3420 VDD.n3419 3.89963
R7599 VDD.n3425 VDD.n3424 3.89963
R7600 VDD.n5377 VDD.n5376 3.89963
R7601 VDD.n3724 VDD.n3723 3.89963
R7602 VDD.n3729 VDD.n3728 3.89963
R7603 VDD.n5448 VDD.n5447 3.89963
R7604 VDD.n2931 VDD.n2930 3.89963
R7605 VDD.n2936 VDD.n2935 3.89963
R7606 VDD.n6185 VDD.n6184 3.89963
R7607 VDD.n3220 VDD.n3219 3.89963
R7608 VDD.n3225 VDD.n3224 3.89963
R7609 VDD.n5311 VDD.n5310 3.89963
R7610 VDD.n2853 VDD.n2852 3.89963
R7611 VDD.n2858 VDD.n2857 3.89963
R7612 VDD.n2558 VDD.n2557 3.89963
R7613 VDD.n1441 VDD.t304 3.88217
R7614 VDD.n7941 VDD.n7907 3.88202
R7615 VDD.n7928 VDD.n7909 3.88202
R7616 VDD.n7912 VDD.n7911 3.88202
R7617 VDD.n370 VDD.n354 3.88202
R7618 VDD.n383 VDD.n352 3.88202
R7619 VDD.n4424 VDD.n4219 3.83311
R7620 VDD.n4434 VDD.n4217 3.83311
R7621 VDD.n4593 VDD.n3915 3.83311
R7622 VDD.n4603 VDD.n3913 3.83311
R7623 VDD.n6519 VDD.n2870 3.83311
R7624 VDD.n6529 VDD.n2868 3.83311
R7625 VDD.n5042 VDD.n3237 3.83311
R7626 VDD.n5052 VDD.n3235 3.83311
R7627 VDD.n5197 VDD.n2926 3.83311
R7628 VDD.n5207 VDD.n2924 3.83311
R7629 VDD.n4740 VDD.n3741 3.83311
R7630 VDD.n4750 VDD.n3739 3.83311
R7631 VDD.n4895 VDD.n3415 3.83311
R7632 VDD.n4905 VDD.n3413 3.83311
R7633 VDD.n813 VDD.t584 3.74664
R7634 VDD.n864 VDD.t576 3.74664
R7635 VDD.n407 VDD.n406 3.6405
R7636 VDD.n7234 VDD.n7233 3.56977
R7637 VDD.n7237 VDD.n7236 3.56963
R7638 VDD.n7237 VDD.n7235 3.5691
R7639 VDD.n2375 VDD.t50 3.48983
R7640 VDD.n2487 VDD.t84 3.48983
R7641 VDD.t119 VDD.t560 3.47876
R7642 VDD.n7883 VDD.n7850 3.4707
R7643 VDD.n7883 VDD.n7882 3.47018
R7644 VDD.n400 VDD.n397 3.4692
R7645 VDD.n401 VDD.n395 3.4692
R7646 VDD.n7966 VDD.n7963 3.4692
R7647 VDD.n7967 VDD.n7961 3.4692
R7648 VDD.n319 VDD.n317 3.44767
R7649 VDD.n316 VDD.n314 3.44767
R7650 VDD.n1123 VDD.n1122 3.3285
R7651 VDD.n1121 VDD.n1120 3.3285
R7652 VDD.n5598 VDD.n5595 3.27354
R7653 VDD.n4202 VDD.n4199 3.27354
R7654 VDD.n4211 VDD.n4208 3.27354
R7655 VDD.n5520 VDD.n5517 3.27354
R7656 VDD.n3920 VDD.n3917 3.27354
R7657 VDD.n3929 VDD.n3926 3.27354
R7658 VDD.n3420 VDD.n3417 3.27354
R7659 VDD.n3425 VDD.n3422 3.27354
R7660 VDD.n5377 VDD.n5374 3.27354
R7661 VDD.n3724 VDD.n3721 3.27354
R7662 VDD.n3729 VDD.n3726 3.27354
R7663 VDD.n5448 VDD.n5445 3.27354
R7664 VDD.n2931 VDD.n2928 3.27354
R7665 VDD.n2936 VDD.n2933 3.27354
R7666 VDD.n6185 VDD.n6182 3.27354
R7667 VDD.n3220 VDD.n3217 3.27354
R7668 VDD.n3225 VDD.n3222 3.27354
R7669 VDD.n5311 VDD.n5308 3.27354
R7670 VDD.n2853 VDD.n2850 3.27354
R7671 VDD.n2858 VDD.n2855 3.27354
R7672 VDD.n2558 VDD.n2555 3.27354
R7673 VDD.n4375 VDD.t289 3.2565
R7674 VDD.n4481 VDD.t231 3.2565
R7675 VDD.n4846 VDD.t240 3.2565
R7676 VDD.n4952 VDD.t257 3.2565
R7677 VDD.n4993 VDD.t159 3.2565
R7678 VDD.n5099 VDD.t168 3.2565
R7679 VDD.n4544 VDD.t226 3.2565
R7680 VDD.n4650 VDD.t254 3.2565
R7681 VDD.n4691 VDD.t147 3.2565
R7682 VDD.n4797 VDD.t141 3.2565
R7683 VDD.n5148 VDD.t150 3.2565
R7684 VDD.n5254 VDD.t213 3.2565
R7685 VDD.n6470 VDD.t144 3.2565
R7686 VDD.n6576 VDD.t245 3.2565
R7687 VDD.n4240 VDD.t317 3.20717
R7688 VDD.n5622 VDD.t321 3.20717
R7689 VDD.n4242 VDD.t336 3.20717
R7690 VDD.n4182 VDD.t364 3.20717
R7691 VDD.n4178 VDD.t334 3.20717
R7692 VDD.n5572 VDD.t285 3.20717
R7693 VDD.n5576 VDD.t232 3.20717
R7694 VDD.n3950 VDD.t278 3.20717
R7695 VDD.n3946 VDD.t227 3.20717
R7696 VDD.n5538 VDD.t380 3.20717
R7697 VDD.n5542 VDD.t362 3.20717
R7698 VDD.n3890 VDD.t310 3.20717
R7699 VDD.n3886 VDD.t255 3.20717
R7700 VDD.n5488 VDD.t354 3.20717
R7701 VDD.n5492 VDD.t332 3.20717
R7702 VDD.n2833 VDD.t325 3.20717
R7703 VDD.n2829 VDD.t292 3.20717
R7704 VDD.n2666 VDD.t300 3.20717
R7705 VDD.n2670 VDD.t246 3.20717
R7706 VDD.n2901 VDD.t248 3.20717
R7707 VDD.n2897 VDD.t214 3.20717
R7708 VDD.n6215 VDD.t287 3.20717
R7709 VDD.n6219 VDD.t234 3.20717
R7710 VDD.n3390 VDD.t386 3.20717
R7711 VDD.n3386 VDD.t368 3.20717
R7712 VDD.n6038 VDD.t312 3.20717
R7713 VDD.n6042 VDD.t258 3.20717
R7714 VDD.n3448 VDD.t319 3.20717
R7715 VDD.n5392 VDD.t294 3.20717
R7716 VDD.n3450 VDD.t342 3.20717
R7717 VDD.n5396 VDD.t241 3.20717
R7718 VDD.n3702 VDD.t243 3.20717
R7719 VDD.n5419 VDD.t188 3.20717
R7720 VDD.n3704 VDD.t296 3.20717
R7721 VDD.n5423 VDD.t142 3.20717
R7722 VDD.n3762 VDD.t148 3.20717
R7723 VDD.n5469 VDD.t306 3.20717
R7724 VDD.n3764 VDD.t190 3.20717
R7725 VDD.n5473 VDD.t250 3.20717
R7726 VDD.n2959 VDD.t221 3.20717
R7727 VDD.n6159 VDD.t192 3.20717
R7728 VDD.n2961 VDD.t260 3.20717
R7729 VDD.n6163 VDD.t151 3.20717
R7730 VDD.n3198 VDD.t169 3.20717
R7731 VDD.n5282 VDD.t348 3.20717
R7732 VDD.n3200 VDD.t198 3.20717
R7733 VDD.n5286 VDD.t323 3.20717
R7734 VDD.n3258 VDD.t356 3.20717
R7735 VDD.n5332 VDD.t194 3.20717
R7736 VDD.n3260 VDD.t378 3.20717
R7737 VDD.n5336 VDD.t160 3.20717
R7738 VDD.n2891 VDD.t382 3.20717
R7739 VDD.n2579 VDD.t200 3.20717
R7740 VDD.n2893 VDD.t145 3.20717
R7741 VDD.n2583 VDD.t174 3.20717
R7742 VDD.n1438 VDD.n1432 3.20717
R7743 VDD.n1437 VDD.n1433 3.20717
R7744 VDD.n1436 VDD.n1434 3.20717
R7745 VDD.n1128 VDD.t298 3.20717
R7746 VDD.n1446 VDD.t274 3.20717
R7747 VDD.n1124 VDD.t352 3.20717
R7748 VDD.n1450 VDD.t272 3.20717
R7749 VDD.n1442 VDD.t302 3.20717
R7750 VDD.n1102 VDD.t196 3.20717
R7751 VDD.n1344 VDD.t184 3.20717
R7752 VDD.n1098 VDD.t276 3.20717
R7753 VDD.n1348 VDD.t180 3.20717
R7754 VDD.n5626 VDD.t290 3.20717
R7755 VDD.n1459 VDD.n1457 3.1914
R7756 VDD.n5749 VDD.n5748 3.1914
R7757 VDD.n2341 VDD.n2340 3.19093
R7758 VDD.n2150 VDD.n2149 3.19093
R7759 VDD.n2047 VDD.n2046 3.19093
R7760 VDD.n5644 VDD.n5643 3.19093
R7761 VDD.n5745 VDD.n5744 3.1908
R7762 VDD.n4518 VDD.n4517 3.1908
R7763 VDD.n6154 VDD.n6153 3.1908
R7764 VDD.n2532 VDD.n2531 3.1908
R7765 VDD.n1241 VDD.n1240 3.1908
R7766 VDD.n7945 VDD.t536 3.18891
R7767 VDD.n6628 VDD.t163 3.18197
R7768 VDD.n6624 VDD.t394 3.18197
R7769 VDD.n6623 VDD.t376 3.18197
R7770 VDD.n6647 VDD.t372 3.18197
R7771 VDD.n550 VDD.t308 3.18197
R7772 VDD.n546 VDD.t280 3.18197
R7773 VDD.n545 VDD.t224 3.18197
R7774 VDD.n6648 VDD.t338 3.18197
R7775 VDD.n558 VDD.t374 3.18197
R7776 VDD.n559 VDD.t346 3.18197
R7777 VDD.n560 VDD.t315 3.18197
R7778 VDD.n872 VDD.t177 3.18197
R7779 VDD.n1030 VDD.t182 3.18197
R7780 VDD.n1031 VDD.t211 3.18197
R7781 VDD.n1033 VDD.t236 3.18197
R7782 VDD.n7890 VDD.t358 3.18197
R7783 VDD.n7057 VDD.t219 3.18197
R7784 VDD.n4350 VDD.n4349 3.1505
R7785 VDD.n5641 VDD.n5640 3.1505
R7786 VDD.n5639 VDD.n5638 3.1505
R7787 VDD.n5636 VDD.n5635 3.1505
R7788 VDD.n5634 VDD.n5633 3.1505
R7789 VDD.n5631 VDD.n5630 3.1505
R7790 VDD.n4244 VDD.n4243 3.1505
R7791 VDD.n4247 VDD.n4246 3.1505
R7792 VDD.n4249 VDD.n4248 3.1505
R7793 VDD.n4252 VDD.n4251 3.1505
R7794 VDD.n4254 VDD.n4253 3.1505
R7795 VDD.n4257 VDD.n4256 3.1505
R7796 VDD.n4259 VDD.n4258 3.1505
R7797 VDD.n4262 VDD.n4261 3.1505
R7798 VDD.n4264 VDD.n4263 3.1505
R7799 VDD.n4267 VDD.n4266 3.1505
R7800 VDD.n4269 VDD.n4268 3.1505
R7801 VDD.n4272 VDD.n4271 3.1505
R7802 VDD.n4274 VDD.n4273 3.1505
R7803 VDD.n4277 VDD.n4276 3.1505
R7804 VDD.n4279 VDD.n4278 3.1505
R7805 VDD.n4282 VDD.n4281 3.1505
R7806 VDD.n4284 VDD.n4283 3.1505
R7807 VDD.n4287 VDD.n4286 3.1505
R7808 VDD.n4289 VDD.n4288 3.1505
R7809 VDD.n4292 VDD.n4291 3.1505
R7810 VDD.n4294 VDD.n4293 3.1505
R7811 VDD.n4297 VDD.n4296 3.1505
R7812 VDD.n4299 VDD.n4298 3.1505
R7813 VDD.n4302 VDD.n4301 3.1505
R7814 VDD.n4304 VDD.n4303 3.1505
R7815 VDD.n4307 VDD.n4306 3.1505
R7816 VDD.n4309 VDD.n4308 3.1505
R7817 VDD.n4312 VDD.n4311 3.1505
R7818 VDD.n4314 VDD.n4313 3.1505
R7819 VDD.n4317 VDD.n4316 3.1505
R7820 VDD.n4319 VDD.n4318 3.1505
R7821 VDD.n4322 VDD.n4321 3.1505
R7822 VDD.n4324 VDD.n4323 3.1505
R7823 VDD.n4327 VDD.n4326 3.1505
R7824 VDD.n4329 VDD.n4328 3.1505
R7825 VDD.n4332 VDD.n4331 3.1505
R7826 VDD.n4334 VDD.n4333 3.1505
R7827 VDD.n4337 VDD.n4336 3.1505
R7828 VDD.n4339 VDD.n4338 3.1505
R7829 VDD.n4342 VDD.n4341 3.1505
R7830 VDD.n4345 VDD.n4344 3.1505
R7831 VDD.n4347 VDD.n4346 3.1505
R7832 VDD.n4177 VDD.n4176 3.1505
R7833 VDD.n5567 VDD.n5566 3.1505
R7834 VDD.n5565 VDD.n5564 3.1505
R7835 VDD.n5563 VDD.n5562 3.1505
R7836 VDD.n4084 VDD.n4083 3.1505
R7837 VDD.n4086 VDD.n4085 3.1505
R7838 VDD.n4088 VDD.n4087 3.1505
R7839 VDD.n4090 VDD.n4089 3.1505
R7840 VDD.n4092 VDD.n4091 3.1505
R7841 VDD.n4094 VDD.n4093 3.1505
R7842 VDD.n4096 VDD.n4095 3.1505
R7843 VDD.n4098 VDD.n4097 3.1505
R7844 VDD.n4100 VDD.n4099 3.1505
R7845 VDD.n4102 VDD.n4101 3.1505
R7846 VDD.n4104 VDD.n4103 3.1505
R7847 VDD.n4106 VDD.n4105 3.1505
R7848 VDD.n4108 VDD.n4107 3.1505
R7849 VDD.n4110 VDD.n4109 3.1505
R7850 VDD.n4112 VDD.n4111 3.1505
R7851 VDD.n4114 VDD.n4113 3.1505
R7852 VDD.n4116 VDD.n4115 3.1505
R7853 VDD.n4118 VDD.n4117 3.1505
R7854 VDD.n4120 VDD.n4119 3.1505
R7855 VDD.n4122 VDD.n4121 3.1505
R7856 VDD.n4124 VDD.n4123 3.1505
R7857 VDD.n4126 VDD.n4125 3.1505
R7858 VDD.n4128 VDD.n4127 3.1505
R7859 VDD.n4130 VDD.n4129 3.1505
R7860 VDD.n4132 VDD.n4131 3.1505
R7861 VDD.n4135 VDD.n4134 3.1505
R7862 VDD.n4137 VDD.n4136 3.1505
R7863 VDD.n4140 VDD.n4139 3.1505
R7864 VDD.n4142 VDD.n4141 3.1505
R7865 VDD.n4145 VDD.n4144 3.1505
R7866 VDD.n4147 VDD.n4146 3.1505
R7867 VDD.n4150 VDD.n4149 3.1505
R7868 VDD.n4152 VDD.n4151 3.1505
R7869 VDD.n4155 VDD.n4154 3.1505
R7870 VDD.n4157 VDD.n4156 3.1505
R7871 VDD.n4160 VDD.n4159 3.1505
R7872 VDD.n4162 VDD.n4161 3.1505
R7873 VDD.n4165 VDD.n4164 3.1505
R7874 VDD.n4167 VDD.n4166 3.1505
R7875 VDD.n4170 VDD.n4169 3.1505
R7876 VDD.n4172 VDD.n4171 3.1505
R7877 VDD.n4175 VDD.n4174 3.1505
R7878 VDD.n5569 VDD.n5568 3.1505
R7879 VDD.n5571 VDD.n5570 3.1505
R7880 VDD.n3385 VDD.n3384 3.1505
R7881 VDD.n3272 VDD.n3271 3.1505
R7882 VDD.n3275 VDD.n3274 3.1505
R7883 VDD.n3277 VDD.n3276 3.1505
R7884 VDD.n3280 VDD.n3279 3.1505
R7885 VDD.n3282 VDD.n3281 3.1505
R7886 VDD.n3285 VDD.n3284 3.1505
R7887 VDD.n3287 VDD.n3286 3.1505
R7888 VDD.n3290 VDD.n3289 3.1505
R7889 VDD.n3292 VDD.n3291 3.1505
R7890 VDD.n3295 VDD.n3294 3.1505
R7891 VDD.n3297 VDD.n3296 3.1505
R7892 VDD.n3300 VDD.n3299 3.1505
R7893 VDD.n3302 VDD.n3301 3.1505
R7894 VDD.n3305 VDD.n3304 3.1505
R7895 VDD.n3307 VDD.n3306 3.1505
R7896 VDD.n3310 VDD.n3309 3.1505
R7897 VDD.n3312 VDD.n3311 3.1505
R7898 VDD.n3315 VDD.n3314 3.1505
R7899 VDD.n3317 VDD.n3316 3.1505
R7900 VDD.n3320 VDD.n3319 3.1505
R7901 VDD.n3322 VDD.n3321 3.1505
R7902 VDD.n3325 VDD.n3324 3.1505
R7903 VDD.n3327 VDD.n3326 3.1505
R7904 VDD.n3330 VDD.n3329 3.1505
R7905 VDD.n3332 VDD.n3331 3.1505
R7906 VDD.n3335 VDD.n3334 3.1505
R7907 VDD.n3337 VDD.n3336 3.1505
R7908 VDD.n3340 VDD.n3339 3.1505
R7909 VDD.n3342 VDD.n3341 3.1505
R7910 VDD.n3345 VDD.n3344 3.1505
R7911 VDD.n3347 VDD.n3346 3.1505
R7912 VDD.n3350 VDD.n3349 3.1505
R7913 VDD.n3352 VDD.n3351 3.1505
R7914 VDD.n3355 VDD.n3354 3.1505
R7915 VDD.n3357 VDD.n3356 3.1505
R7916 VDD.n3360 VDD.n3359 3.1505
R7917 VDD.n3362 VDD.n3361 3.1505
R7918 VDD.n3365 VDD.n3364 3.1505
R7919 VDD.n3367 VDD.n3366 3.1505
R7920 VDD.n3370 VDD.n3369 3.1505
R7921 VDD.n3372 VDD.n3371 3.1505
R7922 VDD.n3375 VDD.n3374 3.1505
R7923 VDD.n3377 VDD.n3376 3.1505
R7924 VDD.n3380 VDD.n3379 3.1505
R7925 VDD.n3382 VDD.n3381 3.1505
R7926 VDD.n3270 VDD.n3269 3.1505
R7927 VDD.n3267 VDD.n3266 3.1505
R7928 VDD.n3265 VDD.n3264 3.1505
R7929 VDD.n5346 VDD.n5345 3.1505
R7930 VDD.n3586 VDD.n3585 3.1505
R7931 VDD.n5410 VDD.n5409 3.1505
R7932 VDD.n3581 VDD.n3580 3.1505
R7933 VDD.n3578 VDD.n3577 3.1505
R7934 VDD.n3575 VDD.n3574 3.1505
R7935 VDD.n3572 VDD.n3571 3.1505
R7936 VDD.n3569 VDD.n3568 3.1505
R7937 VDD.n3566 VDD.n3565 3.1505
R7938 VDD.n3563 VDD.n3562 3.1505
R7939 VDD.n3560 VDD.n3559 3.1505
R7940 VDD.n3557 VDD.n3556 3.1505
R7941 VDD.n3554 VDD.n3553 3.1505
R7942 VDD.n3551 VDD.n3550 3.1505
R7943 VDD.n3548 VDD.n3547 3.1505
R7944 VDD.n3545 VDD.n3544 3.1505
R7945 VDD.n3542 VDD.n3541 3.1505
R7946 VDD.n3539 VDD.n3538 3.1505
R7947 VDD.n3536 VDD.n3535 3.1505
R7948 VDD.n3533 VDD.n3532 3.1505
R7949 VDD.n3530 VDD.n3529 3.1505
R7950 VDD.n3527 VDD.n3526 3.1505
R7951 VDD.n3524 VDD.n3523 3.1505
R7952 VDD.n3521 VDD.n3520 3.1505
R7953 VDD.n3518 VDD.n3517 3.1505
R7954 VDD.n3515 VDD.n3514 3.1505
R7955 VDD.n3512 VDD.n3511 3.1505
R7956 VDD.n3509 VDD.n3508 3.1505
R7957 VDD.n3506 VDD.n3505 3.1505
R7958 VDD.n3503 VDD.n3502 3.1505
R7959 VDD.n3500 VDD.n3499 3.1505
R7960 VDD.n3497 VDD.n3496 3.1505
R7961 VDD.n3494 VDD.n3493 3.1505
R7962 VDD.n3491 VDD.n3490 3.1505
R7963 VDD.n3488 VDD.n3487 3.1505
R7964 VDD.n3485 VDD.n3484 3.1505
R7965 VDD.n3482 VDD.n3481 3.1505
R7966 VDD.n3479 VDD.n3478 3.1505
R7967 VDD.n3476 VDD.n3475 3.1505
R7968 VDD.n3473 VDD.n3472 3.1505
R7969 VDD.n3470 VDD.n3469 3.1505
R7970 VDD.n3467 VDD.n3466 3.1505
R7971 VDD.n3464 VDD.n3463 3.1505
R7972 VDD.n3461 VDD.n3460 3.1505
R7973 VDD.n3458 VDD.n3457 3.1505
R7974 VDD.n3455 VDD.n3454 3.1505
R7975 VDD.n5404 VDD.n5403 3.1505
R7976 VDD.n5407 VDD.n5406 3.1505
R7977 VDD.n3583 VDD.n3582 3.1505
R7978 VDD.n4081 VDD.n4080 3.1505
R7979 VDD.n5561 VDD.n5560 3.1505
R7980 VDD.n4076 VDD.n4075 3.1505
R7981 VDD.n4073 VDD.n4072 3.1505
R7982 VDD.n4070 VDD.n4069 3.1505
R7983 VDD.n4067 VDD.n4066 3.1505
R7984 VDD.n4064 VDD.n4063 3.1505
R7985 VDD.n4061 VDD.n4060 3.1505
R7986 VDD.n4058 VDD.n4057 3.1505
R7987 VDD.n4055 VDD.n4054 3.1505
R7988 VDD.n4052 VDD.n4051 3.1505
R7989 VDD.n4049 VDD.n4048 3.1505
R7990 VDD.n4046 VDD.n4045 3.1505
R7991 VDD.n4043 VDD.n4042 3.1505
R7992 VDD.n4040 VDD.n4039 3.1505
R7993 VDD.n4037 VDD.n4036 3.1505
R7994 VDD.n4034 VDD.n4033 3.1505
R7995 VDD.n4031 VDD.n4030 3.1505
R7996 VDD.n4028 VDD.n4027 3.1505
R7997 VDD.n4025 VDD.n4024 3.1505
R7998 VDD.n4022 VDD.n4021 3.1505
R7999 VDD.n4019 VDD.n4018 3.1505
R8000 VDD.n4016 VDD.n4015 3.1505
R8001 VDD.n4013 VDD.n4012 3.1505
R8002 VDD.n4010 VDD.n4009 3.1505
R8003 VDD.n4007 VDD.n4006 3.1505
R8004 VDD.n4004 VDD.n4003 3.1505
R8005 VDD.n4001 VDD.n4000 3.1505
R8006 VDD.n3998 VDD.n3997 3.1505
R8007 VDD.n3995 VDD.n3994 3.1505
R8008 VDD.n3992 VDD.n3991 3.1505
R8009 VDD.n3989 VDD.n3988 3.1505
R8010 VDD.n3986 VDD.n3985 3.1505
R8011 VDD.n3983 VDD.n3982 3.1505
R8012 VDD.n3980 VDD.n3979 3.1505
R8013 VDD.n3977 VDD.n3976 3.1505
R8014 VDD.n3974 VDD.n3973 3.1505
R8015 VDD.n3971 VDD.n3970 3.1505
R8016 VDD.n3968 VDD.n3967 3.1505
R8017 VDD.n3965 VDD.n3964 3.1505
R8018 VDD.n3962 VDD.n3961 3.1505
R8019 VDD.n3959 VDD.n3958 3.1505
R8020 VDD.n3956 VDD.n3955 3.1505
R8021 VDD.n5550 VDD.n5549 3.1505
R8022 VDD.n5553 VDD.n5552 3.1505
R8023 VDD.n5556 VDD.n5555 3.1505
R8024 VDD.n5559 VDD.n5558 3.1505
R8025 VDD.n4078 VDD.n4077 3.1505
R8026 VDD.n3885 VDD.n3884 3.1505
R8027 VDD.n3772 VDD.n3771 3.1505
R8028 VDD.n3775 VDD.n3774 3.1505
R8029 VDD.n3777 VDD.n3776 3.1505
R8030 VDD.n3780 VDD.n3779 3.1505
R8031 VDD.n3782 VDD.n3781 3.1505
R8032 VDD.n3785 VDD.n3784 3.1505
R8033 VDD.n3787 VDD.n3786 3.1505
R8034 VDD.n3790 VDD.n3789 3.1505
R8035 VDD.n3792 VDD.n3791 3.1505
R8036 VDD.n3795 VDD.n3794 3.1505
R8037 VDD.n3797 VDD.n3796 3.1505
R8038 VDD.n3800 VDD.n3799 3.1505
R8039 VDD.n3802 VDD.n3801 3.1505
R8040 VDD.n3805 VDD.n3804 3.1505
R8041 VDD.n3807 VDD.n3806 3.1505
R8042 VDD.n3810 VDD.n3809 3.1505
R8043 VDD.n3812 VDD.n3811 3.1505
R8044 VDD.n3815 VDD.n3814 3.1505
R8045 VDD.n3817 VDD.n3816 3.1505
R8046 VDD.n3820 VDD.n3819 3.1505
R8047 VDD.n3822 VDD.n3821 3.1505
R8048 VDD.n3825 VDD.n3824 3.1505
R8049 VDD.n3827 VDD.n3826 3.1505
R8050 VDD.n3830 VDD.n3829 3.1505
R8051 VDD.n3832 VDD.n3831 3.1505
R8052 VDD.n3835 VDD.n3834 3.1505
R8053 VDD.n3837 VDD.n3836 3.1505
R8054 VDD.n3840 VDD.n3839 3.1505
R8055 VDD.n3842 VDD.n3841 3.1505
R8056 VDD.n3845 VDD.n3844 3.1505
R8057 VDD.n3847 VDD.n3846 3.1505
R8058 VDD.n3850 VDD.n3849 3.1505
R8059 VDD.n3852 VDD.n3851 3.1505
R8060 VDD.n3855 VDD.n3854 3.1505
R8061 VDD.n3857 VDD.n3856 3.1505
R8062 VDD.n3860 VDD.n3859 3.1505
R8063 VDD.n3862 VDD.n3861 3.1505
R8064 VDD.n3865 VDD.n3864 3.1505
R8065 VDD.n3867 VDD.n3866 3.1505
R8066 VDD.n3870 VDD.n3869 3.1505
R8067 VDD.n3872 VDD.n3871 3.1505
R8068 VDD.n3875 VDD.n3874 3.1505
R8069 VDD.n3877 VDD.n3876 3.1505
R8070 VDD.n3880 VDD.n3879 3.1505
R8071 VDD.n3882 VDD.n3881 3.1505
R8072 VDD.n3770 VDD.n3769 3.1505
R8073 VDD.n5485 VDD.n5484 3.1505
R8074 VDD.n5487 VDD.n5486 3.1505
R8075 VDD.n5483 VDD.n5482 3.1505
R8076 VDD.n3699 VDD.n3698 3.1505
R8077 VDD.n5413 VDD.n5412 3.1505
R8078 VDD.n3588 VDD.n3587 3.1505
R8079 VDD.n3591 VDD.n3590 3.1505
R8080 VDD.n3593 VDD.n3592 3.1505
R8081 VDD.n3596 VDD.n3595 3.1505
R8082 VDD.n3598 VDD.n3597 3.1505
R8083 VDD.n3601 VDD.n3600 3.1505
R8084 VDD.n3603 VDD.n3602 3.1505
R8085 VDD.n3606 VDD.n3605 3.1505
R8086 VDD.n3608 VDD.n3607 3.1505
R8087 VDD.n3611 VDD.n3610 3.1505
R8088 VDD.n3613 VDD.n3612 3.1505
R8089 VDD.n3616 VDD.n3615 3.1505
R8090 VDD.n3618 VDD.n3617 3.1505
R8091 VDD.n3621 VDD.n3620 3.1505
R8092 VDD.n3623 VDD.n3622 3.1505
R8093 VDD.n3626 VDD.n3625 3.1505
R8094 VDD.n3628 VDD.n3627 3.1505
R8095 VDD.n3631 VDD.n3630 3.1505
R8096 VDD.n3633 VDD.n3632 3.1505
R8097 VDD.n3636 VDD.n3635 3.1505
R8098 VDD.n3638 VDD.n3637 3.1505
R8099 VDD.n3641 VDD.n3640 3.1505
R8100 VDD.n3643 VDD.n3642 3.1505
R8101 VDD.n3646 VDD.n3645 3.1505
R8102 VDD.n3648 VDD.n3647 3.1505
R8103 VDD.n3651 VDD.n3650 3.1505
R8104 VDD.n3653 VDD.n3652 3.1505
R8105 VDD.n3656 VDD.n3655 3.1505
R8106 VDD.n3658 VDD.n3657 3.1505
R8107 VDD.n3661 VDD.n3660 3.1505
R8108 VDD.n3663 VDD.n3662 3.1505
R8109 VDD.n3666 VDD.n3665 3.1505
R8110 VDD.n3668 VDD.n3667 3.1505
R8111 VDD.n3671 VDD.n3670 3.1505
R8112 VDD.n3673 VDD.n3672 3.1505
R8113 VDD.n3676 VDD.n3675 3.1505
R8114 VDD.n3678 VDD.n3677 3.1505
R8115 VDD.n3681 VDD.n3680 3.1505
R8116 VDD.n3683 VDD.n3682 3.1505
R8117 VDD.n3686 VDD.n3685 3.1505
R8118 VDD.n3688 VDD.n3687 3.1505
R8119 VDD.n3691 VDD.n3690 3.1505
R8120 VDD.n3694 VDD.n3693 3.1505
R8121 VDD.n3696 VDD.n3695 3.1505
R8122 VDD.n5415 VDD.n5414 3.1505
R8123 VDD.n5418 VDD.n5417 3.1505
R8124 VDD.n5947 VDD.n5946 3.1505
R8125 VDD.n5848 VDD.n5847 3.1505
R8126 VDD.n5850 VDD.n5849 3.1505
R8127 VDD.n5852 VDD.n5851 3.1505
R8128 VDD.n5854 VDD.n5853 3.1505
R8129 VDD.n5857 VDD.n5856 3.1505
R8130 VDD.n5859 VDD.n5858 3.1505
R8131 VDD.n5862 VDD.n5861 3.1505
R8132 VDD.n5864 VDD.n5863 3.1505
R8133 VDD.n5866 VDD.n5865 3.1505
R8134 VDD.n5869 VDD.n5868 3.1505
R8135 VDD.n5871 VDD.n5870 3.1505
R8136 VDD.n5873 VDD.n5872 3.1505
R8137 VDD.n5876 VDD.n5875 3.1505
R8138 VDD.n5878 VDD.n5877 3.1505
R8139 VDD.n5880 VDD.n5879 3.1505
R8140 VDD.n5883 VDD.n5882 3.1505
R8141 VDD.n5885 VDD.n5884 3.1505
R8142 VDD.n5887 VDD.n5886 3.1505
R8143 VDD.n5889 VDD.n5888 3.1505
R8144 VDD.n5891 VDD.n5890 3.1505
R8145 VDD.n5893 VDD.n5892 3.1505
R8146 VDD.n5895 VDD.n5894 3.1505
R8147 VDD.n5897 VDD.n5896 3.1505
R8148 VDD.n5899 VDD.n5898 3.1505
R8149 VDD.n5901 VDD.n5900 3.1505
R8150 VDD.n5903 VDD.n5902 3.1505
R8151 VDD.n5906 VDD.n5905 3.1505
R8152 VDD.n5908 VDD.n5907 3.1505
R8153 VDD.n5910 VDD.n5909 3.1505
R8154 VDD.n5913 VDD.n5912 3.1505
R8155 VDD.n5915 VDD.n5914 3.1505
R8156 VDD.n5917 VDD.n5916 3.1505
R8157 VDD.n5920 VDD.n5919 3.1505
R8158 VDD.n5922 VDD.n5921 3.1505
R8159 VDD.n5924 VDD.n5923 3.1505
R8160 VDD.n5927 VDD.n5926 3.1505
R8161 VDD.n5929 VDD.n5928 3.1505
R8162 VDD.n5932 VDD.n5931 3.1505
R8163 VDD.n5934 VDD.n5933 3.1505
R8164 VDD.n5936 VDD.n5935 3.1505
R8165 VDD.n5938 VDD.n5937 3.1505
R8166 VDD.n5940 VDD.n5939 3.1505
R8167 VDD.n5947 VDD.n5944 3.1505
R8168 VDD.n5951 VDD.n5950 3.1505
R8169 VDD.n5951 VDD.n5948 3.1505
R8170 VDD.n5954 VDD.n5953 3.1505
R8171 VDD.n5956 VDD.n5955 3.1505
R8172 VDD.n5958 VDD.n5957 3.1505
R8173 VDD.n5960 VDD.n5959 3.1505
R8174 VDD.n5962 VDD.n5961 3.1505
R8175 VDD.n5965 VDD.n5964 3.1505
R8176 VDD.n5967 VDD.n5966 3.1505
R8177 VDD.n5970 VDD.n5969 3.1505
R8178 VDD.n5972 VDD.n5971 3.1505
R8179 VDD.n5974 VDD.n5973 3.1505
R8180 VDD.n5977 VDD.n5976 3.1505
R8181 VDD.n5979 VDD.n5978 3.1505
R8182 VDD.n5981 VDD.n5980 3.1505
R8183 VDD.n5984 VDD.n5983 3.1505
R8184 VDD.n5986 VDD.n5985 3.1505
R8185 VDD.n5988 VDD.n5987 3.1505
R8186 VDD.n5991 VDD.n5990 3.1505
R8187 VDD.n5993 VDD.n5992 3.1505
R8188 VDD.n5995 VDD.n5994 3.1505
R8189 VDD.n5997 VDD.n5996 3.1505
R8190 VDD.n5999 VDD.n5998 3.1505
R8191 VDD.n6001 VDD.n6000 3.1505
R8192 VDD.n6003 VDD.n6002 3.1505
R8193 VDD.n6005 VDD.n6004 3.1505
R8194 VDD.n6007 VDD.n6006 3.1505
R8195 VDD.n6009 VDD.n6008 3.1505
R8196 VDD.n6011 VDD.n6010 3.1505
R8197 VDD.n6014 VDD.n6013 3.1505
R8198 VDD.n6016 VDD.n6015 3.1505
R8199 VDD.n6018 VDD.n6017 3.1505
R8200 VDD.n6021 VDD.n6020 3.1505
R8201 VDD.n6023 VDD.n6022 3.1505
R8202 VDD.n6025 VDD.n6024 3.1505
R8203 VDD.n6028 VDD.n6027 3.1505
R8204 VDD.n6030 VDD.n6029 3.1505
R8205 VDD.n6032 VDD.n6031 3.1505
R8206 VDD.n6035 VDD.n6034 3.1505
R8207 VDD.n6037 VDD.n6036 3.1505
R8208 VDD.n6045 VDD.n6044 3.1505
R8209 VDD.n6047 VDD.n6046 3.1505
R8210 VDD.n6049 VDD.n6048 3.1505
R8211 VDD.n6051 VDD.n6050 3.1505
R8212 VDD.n4673 VDD.n4669 3.1505
R8213 VDD.n4818 VDD.n4817 3.1505
R8214 VDD.n4815 VDD.n4814 3.1505
R8215 VDD.n4814 VDD.n4813 3.1505
R8216 VDD.n4812 VDD.n4811 3.1505
R8217 VDD.n4811 VDD.n4810 3.1505
R8218 VDD.n4809 VDD.n4808 3.1505
R8219 VDD.n4808 VDD.n4807 3.1505
R8220 VDD.n4806 VDD.n4805 3.1505
R8221 VDD.n4805 VDD.n4804 3.1505
R8222 VDD.n4803 VDD.n4802 3.1505
R8223 VDD.n4802 VDD.n4801 3.1505
R8224 VDD.n4799 VDD.n4798 3.1505
R8225 VDD.n4798 VDD.n4797 3.1505
R8226 VDD.n4796 VDD.n4795 3.1505
R8227 VDD.n4795 VDD.n4794 3.1505
R8228 VDD.n4792 VDD.n4791 3.1505
R8229 VDD.n4791 VDD.n4790 3.1505
R8230 VDD.n4789 VDD.n4788 3.1505
R8231 VDD.n4788 VDD.n4787 3.1505
R8232 VDD.n4786 VDD.n4785 3.1505
R8233 VDD.n4785 VDD.n4784 3.1505
R8234 VDD.n4782 VDD.n4781 3.1505
R8235 VDD.n4781 VDD.n4780 3.1505
R8236 VDD.n4779 VDD.n4778 3.1505
R8237 VDD.n4778 VDD.n4777 3.1505
R8238 VDD.n4776 VDD.n4775 3.1505
R8239 VDD.n4775 VDD.n4774 3.1505
R8240 VDD.n4772 VDD.n4771 3.1505
R8241 VDD.n4771 VDD.n4770 3.1505
R8242 VDD.n4769 VDD.n4768 3.1505
R8243 VDD.n4768 VDD.n4767 3.1505
R8244 VDD.n4766 VDD.n4765 3.1505
R8245 VDD.n4765 VDD.n4764 3.1505
R8246 VDD.n4762 VDD.n4761 3.1505
R8247 VDD.n4761 VDD.n4760 3.1505
R8248 VDD.n4759 VDD.n4758 3.1505
R8249 VDD.n4758 VDD.n4757 3.1505
R8250 VDD.n4756 VDD.n4755 3.1505
R8251 VDD.n4755 VDD.n4754 3.1505
R8252 VDD.n4753 VDD.n4752 3.1505
R8253 VDD.n4752 VDD.n4751 3.1505
R8254 VDD.n4749 VDD.n4748 3.1505
R8255 VDD.n4748 VDD.n4747 3.1505
R8256 VDD.n4746 VDD.n4745 3.1505
R8257 VDD.n4745 VDD.n4744 3.1505
R8258 VDD.n4743 VDD.n4742 3.1505
R8259 VDD.n4742 VDD.n4741 3.1505
R8260 VDD.n4739 VDD.n4738 3.1505
R8261 VDD.n4738 VDD.n4737 3.1505
R8262 VDD.n4736 VDD.n4735 3.1505
R8263 VDD.n4735 VDD.n4734 3.1505
R8264 VDD.n4733 VDD.n4732 3.1505
R8265 VDD.n4732 VDD.n4731 3.1505
R8266 VDD.n4730 VDD.n4729 3.1505
R8267 VDD.n4729 VDD.n4728 3.1505
R8268 VDD.n4726 VDD.n4725 3.1505
R8269 VDD.n4725 VDD.n4724 3.1505
R8270 VDD.n4723 VDD.n4722 3.1505
R8271 VDD.n4722 VDD.n4721 3.1505
R8272 VDD.n4720 VDD.n4719 3.1505
R8273 VDD.n4719 VDD.n4718 3.1505
R8274 VDD.n4716 VDD.n4715 3.1505
R8275 VDD.n4715 VDD.n4714 3.1505
R8276 VDD.n4713 VDD.n4712 3.1505
R8277 VDD.n4712 VDD.n4711 3.1505
R8278 VDD.n4710 VDD.n4709 3.1505
R8279 VDD.n4709 VDD.n4708 3.1505
R8280 VDD.n4706 VDD.n4705 3.1505
R8281 VDD.n4705 VDD.n4704 3.1505
R8282 VDD.n4703 VDD.n4702 3.1505
R8283 VDD.n4702 VDD.n4701 3.1505
R8284 VDD.n4700 VDD.n4699 3.1505
R8285 VDD.n4699 VDD.n4698 3.1505
R8286 VDD.n4696 VDD.n4695 3.1505
R8287 VDD.n4695 VDD.n4694 3.1505
R8288 VDD.n4693 VDD.n4692 3.1505
R8289 VDD.n4692 VDD.n4691 3.1505
R8290 VDD.n4689 VDD.n4688 3.1505
R8291 VDD.n4688 VDD.n4687 3.1505
R8292 VDD.n4686 VDD.n4685 3.1505
R8293 VDD.n4685 VDD.n4684 3.1505
R8294 VDD.n4683 VDD.n4682 3.1505
R8295 VDD.n4682 VDD.n4681 3.1505
R8296 VDD.n4680 VDD.n4679 3.1505
R8297 VDD.n4679 VDD.n4678 3.1505
R8298 VDD.n4677 VDD.n4676 3.1505
R8299 VDD.n4676 VDD.n4675 3.1505
R8300 VDD.n4673 VDD.n4672 3.1505
R8301 VDD.n4668 VDD.n4667 3.1505
R8302 VDD.n4667 VDD.n4666 3.1505
R8303 VDD.n4827 VDD.n4823 3.1505
R8304 VDD.n4827 VDD.n4826 3.1505
R8305 VDD.n4967 VDD.n4966 3.1505
R8306 VDD.n4966 VDD.n4965 3.1505
R8307 VDD.n4964 VDD.n4963 3.1505
R8308 VDD.n4963 VDD.n4962 3.1505
R8309 VDD.n4961 VDD.n4960 3.1505
R8310 VDD.n4960 VDD.n4959 3.1505
R8311 VDD.n4958 VDD.n4957 3.1505
R8312 VDD.n4957 VDD.n4956 3.1505
R8313 VDD.n4954 VDD.n4953 3.1505
R8314 VDD.n4953 VDD.n4952 3.1505
R8315 VDD.n4951 VDD.n4950 3.1505
R8316 VDD.n4950 VDD.n4949 3.1505
R8317 VDD.n4947 VDD.n4946 3.1505
R8318 VDD.n4946 VDD.n4945 3.1505
R8319 VDD.n4944 VDD.n4943 3.1505
R8320 VDD.n4943 VDD.n4942 3.1505
R8321 VDD.n4941 VDD.n4940 3.1505
R8322 VDD.n4940 VDD.n4939 3.1505
R8323 VDD.n4937 VDD.n4936 3.1505
R8324 VDD.n4936 VDD.n4935 3.1505
R8325 VDD.n4934 VDD.n4933 3.1505
R8326 VDD.n4933 VDD.n4932 3.1505
R8327 VDD.n4931 VDD.n4930 3.1505
R8328 VDD.n4930 VDD.n4929 3.1505
R8329 VDD.n4927 VDD.n4926 3.1505
R8330 VDD.n4926 VDD.n4925 3.1505
R8331 VDD.n4924 VDD.n4923 3.1505
R8332 VDD.n4923 VDD.n4922 3.1505
R8333 VDD.n4921 VDD.n4920 3.1505
R8334 VDD.n4920 VDD.n4919 3.1505
R8335 VDD.n4917 VDD.n4916 3.1505
R8336 VDD.n4916 VDD.n4915 3.1505
R8337 VDD.n4914 VDD.n4913 3.1505
R8338 VDD.n4913 VDD.n4912 3.1505
R8339 VDD.n4911 VDD.n4910 3.1505
R8340 VDD.n4910 VDD.n4909 3.1505
R8341 VDD.n4908 VDD.n4907 3.1505
R8342 VDD.n4907 VDD.n4906 3.1505
R8343 VDD.n4904 VDD.n4903 3.1505
R8344 VDD.n4903 VDD.n4902 3.1505
R8345 VDD.n4901 VDD.n4900 3.1505
R8346 VDD.n4900 VDD.n4899 3.1505
R8347 VDD.n4898 VDD.n4897 3.1505
R8348 VDD.n4897 VDD.n4896 3.1505
R8349 VDD.n4894 VDD.n4893 3.1505
R8350 VDD.n4893 VDD.n4892 3.1505
R8351 VDD.n4891 VDD.n4890 3.1505
R8352 VDD.n4890 VDD.n4889 3.1505
R8353 VDD.n4888 VDD.n4887 3.1505
R8354 VDD.n4887 VDD.n4886 3.1505
R8355 VDD.n4885 VDD.n4884 3.1505
R8356 VDD.n4884 VDD.n4883 3.1505
R8357 VDD.n4881 VDD.n4880 3.1505
R8358 VDD.n4880 VDD.n4879 3.1505
R8359 VDD.n4878 VDD.n4877 3.1505
R8360 VDD.n4877 VDD.n4876 3.1505
R8361 VDD.n4875 VDD.n4874 3.1505
R8362 VDD.n4874 VDD.n4873 3.1505
R8363 VDD.n4871 VDD.n4870 3.1505
R8364 VDD.n4870 VDD.n4869 3.1505
R8365 VDD.n4868 VDD.n4867 3.1505
R8366 VDD.n4867 VDD.n4866 3.1505
R8367 VDD.n4865 VDD.n4864 3.1505
R8368 VDD.n4864 VDD.n4863 3.1505
R8369 VDD.n4861 VDD.n4860 3.1505
R8370 VDD.n4860 VDD.n4859 3.1505
R8371 VDD.n4858 VDD.n4857 3.1505
R8372 VDD.n4857 VDD.n4856 3.1505
R8373 VDD.n4855 VDD.n4854 3.1505
R8374 VDD.n4854 VDD.n4853 3.1505
R8375 VDD.n4851 VDD.n4850 3.1505
R8376 VDD.n4850 VDD.n4849 3.1505
R8377 VDD.n4848 VDD.n4847 3.1505
R8378 VDD.n4847 VDD.n4846 3.1505
R8379 VDD.n4844 VDD.n4843 3.1505
R8380 VDD.n4843 VDD.n4842 3.1505
R8381 VDD.n4841 VDD.n4840 3.1505
R8382 VDD.n4840 VDD.n4839 3.1505
R8383 VDD.n4838 VDD.n4837 3.1505
R8384 VDD.n4837 VDD.n4836 3.1505
R8385 VDD.n4835 VDD.n4834 3.1505
R8386 VDD.n4834 VDD.n4833 3.1505
R8387 VDD.n4832 VDD.n4831 3.1505
R8388 VDD.n4831 VDD.n4830 3.1505
R8389 VDD.n3195 VDD.n3194 3.1505
R8390 VDD.n3082 VDD.n3081 3.1505
R8391 VDD.n3084 VDD.n3083 3.1505
R8392 VDD.n3087 VDD.n3086 3.1505
R8393 VDD.n3089 VDD.n3088 3.1505
R8394 VDD.n3092 VDD.n3091 3.1505
R8395 VDD.n3094 VDD.n3093 3.1505
R8396 VDD.n3097 VDD.n3096 3.1505
R8397 VDD.n3099 VDD.n3098 3.1505
R8398 VDD.n3102 VDD.n3101 3.1505
R8399 VDD.n3104 VDD.n3103 3.1505
R8400 VDD.n3107 VDD.n3106 3.1505
R8401 VDD.n3109 VDD.n3108 3.1505
R8402 VDD.n3112 VDD.n3111 3.1505
R8403 VDD.n3114 VDD.n3113 3.1505
R8404 VDD.n3117 VDD.n3116 3.1505
R8405 VDD.n3119 VDD.n3118 3.1505
R8406 VDD.n3122 VDD.n3121 3.1505
R8407 VDD.n3124 VDD.n3123 3.1505
R8408 VDD.n3127 VDD.n3126 3.1505
R8409 VDD.n3129 VDD.n3128 3.1505
R8410 VDD.n3132 VDD.n3131 3.1505
R8411 VDD.n3134 VDD.n3133 3.1505
R8412 VDD.n3137 VDD.n3136 3.1505
R8413 VDD.n3139 VDD.n3138 3.1505
R8414 VDD.n3142 VDD.n3141 3.1505
R8415 VDD.n3144 VDD.n3143 3.1505
R8416 VDD.n3147 VDD.n3146 3.1505
R8417 VDD.n3149 VDD.n3148 3.1505
R8418 VDD.n3152 VDD.n3151 3.1505
R8419 VDD.n3154 VDD.n3153 3.1505
R8420 VDD.n3157 VDD.n3156 3.1505
R8421 VDD.n3159 VDD.n3158 3.1505
R8422 VDD.n3162 VDD.n3161 3.1505
R8423 VDD.n3164 VDD.n3163 3.1505
R8424 VDD.n3167 VDD.n3166 3.1505
R8425 VDD.n3169 VDD.n3168 3.1505
R8426 VDD.n3172 VDD.n3171 3.1505
R8427 VDD.n3174 VDD.n3173 3.1505
R8428 VDD.n3177 VDD.n3176 3.1505
R8429 VDD.n3179 VDD.n3178 3.1505
R8430 VDD.n3182 VDD.n3181 3.1505
R8431 VDD.n3184 VDD.n3183 3.1505
R8432 VDD.n3187 VDD.n3186 3.1505
R8433 VDD.n3190 VDD.n3189 3.1505
R8434 VDD.n3192 VDD.n3191 3.1505
R8435 VDD.n5278 VDD.n5277 3.1505
R8436 VDD.n5281 VDD.n5280 3.1505
R8437 VDD.n3079 VDD.n3078 3.1505
R8438 VDD.n5275 VDD.n5274 3.1505
R8439 VDD.n3074 VDD.n3073 3.1505
R8440 VDD.n3072 VDD.n3071 3.1505
R8441 VDD.n3069 VDD.n3068 3.1505
R8442 VDD.n3067 VDD.n3066 3.1505
R8443 VDD.n3064 VDD.n3063 3.1505
R8444 VDD.n3062 VDD.n3061 3.1505
R8445 VDD.n3059 VDD.n3058 3.1505
R8446 VDD.n3057 VDD.n3056 3.1505
R8447 VDD.n3054 VDD.n3053 3.1505
R8448 VDD.n3052 VDD.n3051 3.1505
R8449 VDD.n3049 VDD.n3048 3.1505
R8450 VDD.n3047 VDD.n3046 3.1505
R8451 VDD.n3044 VDD.n3043 3.1505
R8452 VDD.n3042 VDD.n3041 3.1505
R8453 VDD.n3039 VDD.n3038 3.1505
R8454 VDD.n3037 VDD.n3036 3.1505
R8455 VDD.n3034 VDD.n3033 3.1505
R8456 VDD.n3032 VDD.n3031 3.1505
R8457 VDD.n3029 VDD.n3028 3.1505
R8458 VDD.n3027 VDD.n3026 3.1505
R8459 VDD.n3024 VDD.n3023 3.1505
R8460 VDD.n3022 VDD.n3021 3.1505
R8461 VDD.n3019 VDD.n3018 3.1505
R8462 VDD.n3017 VDD.n3016 3.1505
R8463 VDD.n3014 VDD.n3013 3.1505
R8464 VDD.n3012 VDD.n3011 3.1505
R8465 VDD.n3009 VDD.n3008 3.1505
R8466 VDD.n3007 VDD.n3006 3.1505
R8467 VDD.n3004 VDD.n3003 3.1505
R8468 VDD.n3002 VDD.n3001 3.1505
R8469 VDD.n2999 VDD.n2998 3.1505
R8470 VDD.n2997 VDD.n2996 3.1505
R8471 VDD.n2994 VDD.n2993 3.1505
R8472 VDD.n2992 VDD.n2991 3.1505
R8473 VDD.n2989 VDD.n2988 3.1505
R8474 VDD.n2987 VDD.n2986 3.1505
R8475 VDD.n2984 VDD.n2983 3.1505
R8476 VDD.n2982 VDD.n2981 3.1505
R8477 VDD.n2979 VDD.n2978 3.1505
R8478 VDD.n2977 VDD.n2976 3.1505
R8479 VDD.n2974 VDD.n2973 3.1505
R8480 VDD.n2972 VDD.n2971 3.1505
R8481 VDD.n2969 VDD.n2968 3.1505
R8482 VDD.n2967 VDD.n2966 3.1505
R8483 VDD.n5273 VDD.n5272 3.1505
R8484 VDD.n3077 VDD.n3076 3.1505
R8485 VDD.n6054 VDD.n6053 3.1505
R8486 VDD.n6056 VDD.n6055 3.1505
R8487 VDD.n6058 VDD.n6057 3.1505
R8488 VDD.n6060 VDD.n6059 3.1505
R8489 VDD.n6063 VDD.n6062 3.1505
R8490 VDD.n6065 VDD.n6064 3.1505
R8491 VDD.n6068 VDD.n6067 3.1505
R8492 VDD.n6070 VDD.n6069 3.1505
R8493 VDD.n6072 VDD.n6071 3.1505
R8494 VDD.n6075 VDD.n6074 3.1505
R8495 VDD.n6077 VDD.n6076 3.1505
R8496 VDD.n6079 VDD.n6078 3.1505
R8497 VDD.n6082 VDD.n6081 3.1505
R8498 VDD.n6084 VDD.n6083 3.1505
R8499 VDD.n6086 VDD.n6085 3.1505
R8500 VDD.n6089 VDD.n6088 3.1505
R8501 VDD.n6091 VDD.n6090 3.1505
R8502 VDD.n6093 VDD.n6092 3.1505
R8503 VDD.n6095 VDD.n6094 3.1505
R8504 VDD.n6097 VDD.n6096 3.1505
R8505 VDD.n6099 VDD.n6098 3.1505
R8506 VDD.n6101 VDD.n6100 3.1505
R8507 VDD.n6103 VDD.n6102 3.1505
R8508 VDD.n6105 VDD.n6104 3.1505
R8509 VDD.n6107 VDD.n6106 3.1505
R8510 VDD.n6109 VDD.n6108 3.1505
R8511 VDD.n6112 VDD.n6111 3.1505
R8512 VDD.n6114 VDD.n6113 3.1505
R8513 VDD.n6116 VDD.n6115 3.1505
R8514 VDD.n6119 VDD.n6118 3.1505
R8515 VDD.n6121 VDD.n6120 3.1505
R8516 VDD.n6123 VDD.n6122 3.1505
R8517 VDD.n6126 VDD.n6125 3.1505
R8518 VDD.n6128 VDD.n6127 3.1505
R8519 VDD.n6130 VDD.n6129 3.1505
R8520 VDD.n6133 VDD.n6132 3.1505
R8521 VDD.n6135 VDD.n6134 3.1505
R8522 VDD.n6138 VDD.n6137 3.1505
R8523 VDD.n6140 VDD.n6139 3.1505
R8524 VDD.n6142 VDD.n6141 3.1505
R8525 VDD.n6144 VDD.n6143 3.1505
R8526 VDD.n6146 VDD.n6145 3.1505
R8527 VDD.n6305 VDD.n6304 3.1505
R8528 VDD.n6303 VDD.n6302 3.1505
R8529 VDD.n6301 VDD.n6300 3.1505
R8530 VDD.n6299 VDD.n6298 3.1505
R8531 VDD.n6297 VDD.n6296 3.1505
R8532 VDD.n6294 VDD.n6293 3.1505
R8533 VDD.n6292 VDD.n6291 3.1505
R8534 VDD.n6289 VDD.n6288 3.1505
R8535 VDD.n6287 VDD.n6286 3.1505
R8536 VDD.n6285 VDD.n6284 3.1505
R8537 VDD.n6282 VDD.n6281 3.1505
R8538 VDD.n6280 VDD.n6279 3.1505
R8539 VDD.n6278 VDD.n6277 3.1505
R8540 VDD.n6275 VDD.n6274 3.1505
R8541 VDD.n6273 VDD.n6272 3.1505
R8542 VDD.n6271 VDD.n6270 3.1505
R8543 VDD.n6268 VDD.n6267 3.1505
R8544 VDD.n6266 VDD.n6265 3.1505
R8545 VDD.n6264 VDD.n6263 3.1505
R8546 VDD.n6262 VDD.n6261 3.1505
R8547 VDD.n6260 VDD.n6259 3.1505
R8548 VDD.n6258 VDD.n6257 3.1505
R8549 VDD.n6256 VDD.n6255 3.1505
R8550 VDD.n6254 VDD.n6253 3.1505
R8551 VDD.n6252 VDD.n6251 3.1505
R8552 VDD.n6250 VDD.n6249 3.1505
R8553 VDD.n6248 VDD.n6247 3.1505
R8554 VDD.n6245 VDD.n6244 3.1505
R8555 VDD.n6243 VDD.n6242 3.1505
R8556 VDD.n6241 VDD.n6240 3.1505
R8557 VDD.n6238 VDD.n6237 3.1505
R8558 VDD.n6236 VDD.n6235 3.1505
R8559 VDD.n6234 VDD.n6233 3.1505
R8560 VDD.n6231 VDD.n6230 3.1505
R8561 VDD.n6229 VDD.n6228 3.1505
R8562 VDD.n6227 VDD.n6226 3.1505
R8563 VDD.n6224 VDD.n6223 3.1505
R8564 VDD.n6222 VDD.n6221 3.1505
R8565 VDD.n6214 VDD.n6213 3.1505
R8566 VDD.n6212 VDD.n6211 3.1505
R8567 VDD.n6210 VDD.n6209 3.1505
R8568 VDD.n5271 VDD.n5270 3.1505
R8569 VDD.n5123 VDD.n5122 3.1505
R8570 VDD.n4975 VDD.n4971 3.1505
R8571 VDD.n5123 VDD.n5119 3.1505
R8572 VDD.n5117 VDD.n5116 3.1505
R8573 VDD.n5116 VDD.n5115 3.1505
R8574 VDD.n5114 VDD.n5113 3.1505
R8575 VDD.n5113 VDD.n5112 3.1505
R8576 VDD.n5111 VDD.n5110 3.1505
R8577 VDD.n5110 VDD.n5109 3.1505
R8578 VDD.n5108 VDD.n5107 3.1505
R8579 VDD.n5107 VDD.n5106 3.1505
R8580 VDD.n5105 VDD.n5104 3.1505
R8581 VDD.n5104 VDD.n5103 3.1505
R8582 VDD.n5101 VDD.n5100 3.1505
R8583 VDD.n5100 VDD.n5099 3.1505
R8584 VDD.n5098 VDD.n5097 3.1505
R8585 VDD.n5097 VDD.n5096 3.1505
R8586 VDD.n5094 VDD.n5093 3.1505
R8587 VDD.n5093 VDD.n5092 3.1505
R8588 VDD.n5091 VDD.n5090 3.1505
R8589 VDD.n5090 VDD.n5089 3.1505
R8590 VDD.n5088 VDD.n5087 3.1505
R8591 VDD.n5087 VDD.n5086 3.1505
R8592 VDD.n5084 VDD.n5083 3.1505
R8593 VDD.n5083 VDD.n5082 3.1505
R8594 VDD.n5081 VDD.n5080 3.1505
R8595 VDD.n5080 VDD.n5079 3.1505
R8596 VDD.n5078 VDD.n5077 3.1505
R8597 VDD.n5077 VDD.n5076 3.1505
R8598 VDD.n5074 VDD.n5073 3.1505
R8599 VDD.n5073 VDD.n5072 3.1505
R8600 VDD.n5071 VDD.n5070 3.1505
R8601 VDD.n5070 VDD.n5069 3.1505
R8602 VDD.n5068 VDD.n5067 3.1505
R8603 VDD.n5067 VDD.n5066 3.1505
R8604 VDD.n5064 VDD.n5063 3.1505
R8605 VDD.n5063 VDD.n5062 3.1505
R8606 VDD.n5061 VDD.n5060 3.1505
R8607 VDD.n5060 VDD.n5059 3.1505
R8608 VDD.n5058 VDD.n5057 3.1505
R8609 VDD.n5057 VDD.n5056 3.1505
R8610 VDD.n5055 VDD.n5054 3.1505
R8611 VDD.n5054 VDD.n5053 3.1505
R8612 VDD.n5051 VDD.n5050 3.1505
R8613 VDD.n5050 VDD.n5049 3.1505
R8614 VDD.n5048 VDD.n5047 3.1505
R8615 VDD.n5047 VDD.n5046 3.1505
R8616 VDD.n5045 VDD.n5044 3.1505
R8617 VDD.n5044 VDD.n5043 3.1505
R8618 VDD.n5041 VDD.n5040 3.1505
R8619 VDD.n5040 VDD.n5039 3.1505
R8620 VDD.n5038 VDD.n5037 3.1505
R8621 VDD.n5037 VDD.n5036 3.1505
R8622 VDD.n5035 VDD.n5034 3.1505
R8623 VDD.n5034 VDD.n5033 3.1505
R8624 VDD.n5032 VDD.n5031 3.1505
R8625 VDD.n5031 VDD.n5030 3.1505
R8626 VDD.n5028 VDD.n5027 3.1505
R8627 VDD.n5027 VDD.n5026 3.1505
R8628 VDD.n5025 VDD.n5024 3.1505
R8629 VDD.n5024 VDD.n5023 3.1505
R8630 VDD.n5022 VDD.n5021 3.1505
R8631 VDD.n5021 VDD.n5020 3.1505
R8632 VDD.n5018 VDD.n5017 3.1505
R8633 VDD.n5017 VDD.n5016 3.1505
R8634 VDD.n5015 VDD.n5014 3.1505
R8635 VDD.n5014 VDD.n5013 3.1505
R8636 VDD.n5012 VDD.n5011 3.1505
R8637 VDD.n5011 VDD.n5010 3.1505
R8638 VDD.n5008 VDD.n5007 3.1505
R8639 VDD.n5007 VDD.n5006 3.1505
R8640 VDD.n5005 VDD.n5004 3.1505
R8641 VDD.n5004 VDD.n5003 3.1505
R8642 VDD.n5002 VDD.n5001 3.1505
R8643 VDD.n5001 VDD.n5000 3.1505
R8644 VDD.n4998 VDD.n4997 3.1505
R8645 VDD.n4997 VDD.n4996 3.1505
R8646 VDD.n4995 VDD.n4994 3.1505
R8647 VDD.n4994 VDD.n4993 3.1505
R8648 VDD.n4991 VDD.n4990 3.1505
R8649 VDD.n4990 VDD.n4989 3.1505
R8650 VDD.n4988 VDD.n4987 3.1505
R8651 VDD.n4987 VDD.n4986 3.1505
R8652 VDD.n4985 VDD.n4984 3.1505
R8653 VDD.n4984 VDD.n4983 3.1505
R8654 VDD.n4982 VDD.n4981 3.1505
R8655 VDD.n4981 VDD.n4980 3.1505
R8656 VDD.n4979 VDD.n4978 3.1505
R8657 VDD.n4978 VDD.n4977 3.1505
R8658 VDD.n4975 VDD.n4974 3.1505
R8659 VDD.n4970 VDD.n4969 3.1505
R8660 VDD.n4969 VDD.n4968 3.1505
R8661 VDD.n5129 VDD.n5127 3.1505
R8662 VDD.n5129 VDD.n5128 3.1505
R8663 VDD.n5269 VDD.n5268 3.1505
R8664 VDD.n5268 VDD.n5267 3.1505
R8665 VDD.n5266 VDD.n5265 3.1505
R8666 VDD.n5265 VDD.n5264 3.1505
R8667 VDD.n5263 VDD.n5262 3.1505
R8668 VDD.n5262 VDD.n5261 3.1505
R8669 VDD.n5260 VDD.n5259 3.1505
R8670 VDD.n5259 VDD.n5258 3.1505
R8671 VDD.n5256 VDD.n5255 3.1505
R8672 VDD.n5255 VDD.n5254 3.1505
R8673 VDD.n5253 VDD.n5252 3.1505
R8674 VDD.n5252 VDD.n5251 3.1505
R8675 VDD.n5249 VDD.n5248 3.1505
R8676 VDD.n5248 VDD.n5247 3.1505
R8677 VDD.n5246 VDD.n5245 3.1505
R8678 VDD.n5245 VDD.n5244 3.1505
R8679 VDD.n5243 VDD.n5242 3.1505
R8680 VDD.n5242 VDD.n5241 3.1505
R8681 VDD.n5239 VDD.n5238 3.1505
R8682 VDD.n5238 VDD.n5237 3.1505
R8683 VDD.n5236 VDD.n5235 3.1505
R8684 VDD.n5235 VDD.n5234 3.1505
R8685 VDD.n5233 VDD.n5232 3.1505
R8686 VDD.n5232 VDD.n5231 3.1505
R8687 VDD.n5229 VDD.n5228 3.1505
R8688 VDD.n5228 VDD.n5227 3.1505
R8689 VDD.n5226 VDD.n5225 3.1505
R8690 VDD.n5225 VDD.n5224 3.1505
R8691 VDD.n5223 VDD.n5222 3.1505
R8692 VDD.n5222 VDD.n5221 3.1505
R8693 VDD.n5219 VDD.n5218 3.1505
R8694 VDD.n5218 VDD.n5217 3.1505
R8695 VDD.n5216 VDD.n5215 3.1505
R8696 VDD.n5215 VDD.n5214 3.1505
R8697 VDD.n5213 VDD.n5212 3.1505
R8698 VDD.n5212 VDD.n5211 3.1505
R8699 VDD.n5210 VDD.n5209 3.1505
R8700 VDD.n5209 VDD.n5208 3.1505
R8701 VDD.n5206 VDD.n5205 3.1505
R8702 VDD.n5205 VDD.n5204 3.1505
R8703 VDD.n5203 VDD.n5202 3.1505
R8704 VDD.n5202 VDD.n5201 3.1505
R8705 VDD.n5200 VDD.n5199 3.1505
R8706 VDD.n5199 VDD.n5198 3.1505
R8707 VDD.n5196 VDD.n5195 3.1505
R8708 VDD.n5195 VDD.n5194 3.1505
R8709 VDD.n5193 VDD.n5192 3.1505
R8710 VDD.n5192 VDD.n5191 3.1505
R8711 VDD.n5190 VDD.n5189 3.1505
R8712 VDD.n5189 VDD.n5188 3.1505
R8713 VDD.n5187 VDD.n5186 3.1505
R8714 VDD.n5186 VDD.n5185 3.1505
R8715 VDD.n5183 VDD.n5182 3.1505
R8716 VDD.n5182 VDD.n5181 3.1505
R8717 VDD.n5180 VDD.n5179 3.1505
R8718 VDD.n5179 VDD.n5178 3.1505
R8719 VDD.n5177 VDD.n5176 3.1505
R8720 VDD.n5176 VDD.n5175 3.1505
R8721 VDD.n5173 VDD.n5172 3.1505
R8722 VDD.n5172 VDD.n5171 3.1505
R8723 VDD.n5170 VDD.n5169 3.1505
R8724 VDD.n5169 VDD.n5168 3.1505
R8725 VDD.n5167 VDD.n5166 3.1505
R8726 VDD.n5166 VDD.n5165 3.1505
R8727 VDD.n5163 VDD.n5162 3.1505
R8728 VDD.n5162 VDD.n5161 3.1505
R8729 VDD.n5160 VDD.n5159 3.1505
R8730 VDD.n5159 VDD.n5158 3.1505
R8731 VDD.n5157 VDD.n5156 3.1505
R8732 VDD.n5156 VDD.n5155 3.1505
R8733 VDD.n5153 VDD.n5152 3.1505
R8734 VDD.n5152 VDD.n5151 3.1505
R8735 VDD.n5150 VDD.n5149 3.1505
R8736 VDD.n5149 VDD.n5148 3.1505
R8737 VDD.n5146 VDD.n5145 3.1505
R8738 VDD.n5145 VDD.n5144 3.1505
R8739 VDD.n5143 VDD.n5142 3.1505
R8740 VDD.n5142 VDD.n5141 3.1505
R8741 VDD.n5140 VDD.n5139 3.1505
R8742 VDD.n5139 VDD.n5138 3.1505
R8743 VDD.n5137 VDD.n5136 3.1505
R8744 VDD.n5136 VDD.n5135 3.1505
R8745 VDD.n5134 VDD.n5133 3.1505
R8746 VDD.n5133 VDD.n5132 3.1505
R8747 VDD.n6450 VDD.n6449 3.1505
R8748 VDD.n6447 VDD.n6446 3.1505
R8749 VDD.n6444 VDD.n6443 3.1505
R8750 VDD.n6330 VDD.n6329 3.1505
R8751 VDD.n6332 VDD.n6331 3.1505
R8752 VDD.n6335 VDD.n6334 3.1505
R8753 VDD.n6337 VDD.n6336 3.1505
R8754 VDD.n6340 VDD.n6339 3.1505
R8755 VDD.n6342 VDD.n6341 3.1505
R8756 VDD.n6345 VDD.n6344 3.1505
R8757 VDD.n6347 VDD.n6346 3.1505
R8758 VDD.n6350 VDD.n6349 3.1505
R8759 VDD.n6352 VDD.n6351 3.1505
R8760 VDD.n6355 VDD.n6354 3.1505
R8761 VDD.n6357 VDD.n6356 3.1505
R8762 VDD.n6360 VDD.n6359 3.1505
R8763 VDD.n6362 VDD.n6361 3.1505
R8764 VDD.n6365 VDD.n6364 3.1505
R8765 VDD.n6367 VDD.n6366 3.1505
R8766 VDD.n6370 VDD.n6369 3.1505
R8767 VDD.n6372 VDD.n6371 3.1505
R8768 VDD.n6375 VDD.n6374 3.1505
R8769 VDD.n6377 VDD.n6376 3.1505
R8770 VDD.n6380 VDD.n6379 3.1505
R8771 VDD.n6382 VDD.n6381 3.1505
R8772 VDD.n6385 VDD.n6384 3.1505
R8773 VDD.n6387 VDD.n6386 3.1505
R8774 VDD.n6390 VDD.n6389 3.1505
R8775 VDD.n6392 VDD.n6391 3.1505
R8776 VDD.n6395 VDD.n6394 3.1505
R8777 VDD.n6397 VDD.n6396 3.1505
R8778 VDD.n6400 VDD.n6399 3.1505
R8779 VDD.n6402 VDD.n6401 3.1505
R8780 VDD.n6405 VDD.n6404 3.1505
R8781 VDD.n6407 VDD.n6406 3.1505
R8782 VDD.n6410 VDD.n6409 3.1505
R8783 VDD.n6412 VDD.n6411 3.1505
R8784 VDD.n6415 VDD.n6414 3.1505
R8785 VDD.n6417 VDD.n6416 3.1505
R8786 VDD.n6420 VDD.n6419 3.1505
R8787 VDD.n6422 VDD.n6421 3.1505
R8788 VDD.n6425 VDD.n6424 3.1505
R8789 VDD.n6427 VDD.n6426 3.1505
R8790 VDD.n6430 VDD.n6429 3.1505
R8791 VDD.n6432 VDD.n6431 3.1505
R8792 VDD.n6436 VDD.n6435 3.1505
R8793 VDD.n6439 VDD.n6438 3.1505
R8794 VDD.n6441 VDD.n6440 3.1505
R8795 VDD.n6327 VDD.n6326 3.1505
R8796 VDD.n6324 VDD.n6323 3.1505
R8797 VDD.n6321 VDD.n6320 3.1505
R8798 VDD.n6453 VDD.n6452 3.1505
R8799 VDD.n6314 VDD.n6313 3.1505
R8800 VDD.n2828 VDD.n2827 3.1505
R8801 VDD.n2825 VDD.n2824 3.1505
R8802 VDD.n2822 VDD.n2821 3.1505
R8803 VDD.n2819 VDD.n2818 3.1505
R8804 VDD.n2816 VDD.n2815 3.1505
R8805 VDD.n2813 VDD.n2812 3.1505
R8806 VDD.n2810 VDD.n2809 3.1505
R8807 VDD.n2807 VDD.n2806 3.1505
R8808 VDD.n2804 VDD.n2803 3.1505
R8809 VDD.n2801 VDD.n2800 3.1505
R8810 VDD.n2798 VDD.n2797 3.1505
R8811 VDD.n2795 VDD.n2794 3.1505
R8812 VDD.n2792 VDD.n2791 3.1505
R8813 VDD.n2789 VDD.n2788 3.1505
R8814 VDD.n2786 VDD.n2785 3.1505
R8815 VDD.n2783 VDD.n2782 3.1505
R8816 VDD.n2780 VDD.n2779 3.1505
R8817 VDD.n2777 VDD.n2776 3.1505
R8818 VDD.n2774 VDD.n2773 3.1505
R8819 VDD.n2771 VDD.n2770 3.1505
R8820 VDD.n2768 VDD.n2767 3.1505
R8821 VDD.n2765 VDD.n2764 3.1505
R8822 VDD.n2762 VDD.n2761 3.1505
R8823 VDD.n2759 VDD.n2758 3.1505
R8824 VDD.n2756 VDD.n2755 3.1505
R8825 VDD.n2753 VDD.n2752 3.1505
R8826 VDD.n2750 VDD.n2749 3.1505
R8827 VDD.n2747 VDD.n2746 3.1505
R8828 VDD.n2744 VDD.n2743 3.1505
R8829 VDD.n2741 VDD.n2740 3.1505
R8830 VDD.n2738 VDD.n2737 3.1505
R8831 VDD.n2735 VDD.n2734 3.1505
R8832 VDD.n2732 VDD.n2731 3.1505
R8833 VDD.n2729 VDD.n2728 3.1505
R8834 VDD.n2726 VDD.n2725 3.1505
R8835 VDD.n2723 VDD.n2722 3.1505
R8836 VDD.n2720 VDD.n2719 3.1505
R8837 VDD.n2717 VDD.n2716 3.1505
R8838 VDD.n2714 VDD.n2713 3.1505
R8839 VDD.n2711 VDD.n2710 3.1505
R8840 VDD.n2708 VDD.n2707 3.1505
R8841 VDD.n2705 VDD.n2704 3.1505
R8842 VDD.n2702 VDD.n2701 3.1505
R8843 VDD.n2699 VDD.n2698 3.1505
R8844 VDD.n2696 VDD.n2695 3.1505
R8845 VDD.n2693 VDD.n2692 3.1505
R8846 VDD.n2690 VDD.n2689 3.1505
R8847 VDD.n2687 VDD.n2686 3.1505
R8848 VDD.n6318 VDD.n6317 3.1505
R8849 VDD.n6316 VDD.n6315 3.1505
R8850 VDD.n2588 VDD.n2587 3.1505
R8851 VDD.n2590 VDD.n2589 3.1505
R8852 VDD.n2593 VDD.n2592 3.1505
R8853 VDD.n2595 VDD.n2594 3.1505
R8854 VDD.n2598 VDD.n2597 3.1505
R8855 VDD.n2600 VDD.n2599 3.1505
R8856 VDD.n2602 VDD.n2601 3.1505
R8857 VDD.n2605 VDD.n2604 3.1505
R8858 VDD.n2607 VDD.n2606 3.1505
R8859 VDD.n2609 VDD.n2608 3.1505
R8860 VDD.n2612 VDD.n2611 3.1505
R8861 VDD.n2614 VDD.n2613 3.1505
R8862 VDD.n2616 VDD.n2615 3.1505
R8863 VDD.n2619 VDD.n2618 3.1505
R8864 VDD.n2621 VDD.n2620 3.1505
R8865 VDD.n2623 VDD.n2622 3.1505
R8866 VDD.n2625 VDD.n2624 3.1505
R8867 VDD.n2627 VDD.n2626 3.1505
R8868 VDD.n2629 VDD.n2628 3.1505
R8869 VDD.n2631 VDD.n2630 3.1505
R8870 VDD.n2633 VDD.n2632 3.1505
R8871 VDD.n2635 VDD.n2634 3.1505
R8872 VDD.n2637 VDD.n2636 3.1505
R8873 VDD.n2639 VDD.n2638 3.1505
R8874 VDD.n2642 VDD.n2641 3.1505
R8875 VDD.n2644 VDD.n2643 3.1505
R8876 VDD.n2646 VDD.n2645 3.1505
R8877 VDD.n2649 VDD.n2648 3.1505
R8878 VDD.n2651 VDD.n2650 3.1505
R8879 VDD.n2653 VDD.n2652 3.1505
R8880 VDD.n2656 VDD.n2655 3.1505
R8881 VDD.n2658 VDD.n2657 3.1505
R8882 VDD.n2660 VDD.n2659 3.1505
R8883 VDD.n2663 VDD.n2662 3.1505
R8884 VDD.n2665 VDD.n2664 3.1505
R8885 VDD.n2673 VDD.n2672 3.1505
R8886 VDD.n2675 VDD.n2674 3.1505
R8887 VDD.n2677 VDD.n2676 3.1505
R8888 VDD.n2679 VDD.n2678 3.1505
R8889 VDD.n2681 VDD.n2680 3.1505
R8890 VDD.n6599 VDD.n6595 3.1505
R8891 VDD.n6599 VDD.n6598 3.1505
R8892 VDD.n6594 VDD.n6593 3.1505
R8893 VDD.n6593 VDD.n6592 3.1505
R8894 VDD.n6591 VDD.n6590 3.1505
R8895 VDD.n6590 VDD.n6589 3.1505
R8896 VDD.n6588 VDD.n6587 3.1505
R8897 VDD.n6587 VDD.n6586 3.1505
R8898 VDD.n6585 VDD.n6584 3.1505
R8899 VDD.n6584 VDD.n6583 3.1505
R8900 VDD.n6582 VDD.n6581 3.1505
R8901 VDD.n6581 VDD.n6580 3.1505
R8902 VDD.n6578 VDD.n6577 3.1505
R8903 VDD.n6577 VDD.n6576 3.1505
R8904 VDD.n6575 VDD.n6574 3.1505
R8905 VDD.n6574 VDD.n6573 3.1505
R8906 VDD.n6571 VDD.n6570 3.1505
R8907 VDD.n6570 VDD.n6569 3.1505
R8908 VDD.n6568 VDD.n6567 3.1505
R8909 VDD.n6567 VDD.n6566 3.1505
R8910 VDD.n6565 VDD.n6564 3.1505
R8911 VDD.n6564 VDD.n6563 3.1505
R8912 VDD.n6561 VDD.n6560 3.1505
R8913 VDD.n6560 VDD.n6559 3.1505
R8914 VDD.n6558 VDD.n6557 3.1505
R8915 VDD.n6557 VDD.n6556 3.1505
R8916 VDD.n6555 VDD.n6554 3.1505
R8917 VDD.n6554 VDD.n6553 3.1505
R8918 VDD.n6551 VDD.n6550 3.1505
R8919 VDD.n6550 VDD.n6549 3.1505
R8920 VDD.n6548 VDD.n6547 3.1505
R8921 VDD.n6547 VDD.n6546 3.1505
R8922 VDD.n6545 VDD.n6544 3.1505
R8923 VDD.n6544 VDD.n6543 3.1505
R8924 VDD.n6541 VDD.n6540 3.1505
R8925 VDD.n6540 VDD.n6539 3.1505
R8926 VDD.n6538 VDD.n6537 3.1505
R8927 VDD.n6537 VDD.n6536 3.1505
R8928 VDD.n6535 VDD.n6534 3.1505
R8929 VDD.n6534 VDD.n6533 3.1505
R8930 VDD.n6532 VDD.n6531 3.1505
R8931 VDD.n6531 VDD.n6530 3.1505
R8932 VDD.n6528 VDD.n6527 3.1505
R8933 VDD.n6527 VDD.n6526 3.1505
R8934 VDD.n6525 VDD.n6524 3.1505
R8935 VDD.n6524 VDD.n6523 3.1505
R8936 VDD.n6522 VDD.n6521 3.1505
R8937 VDD.n6521 VDD.n6520 3.1505
R8938 VDD.n6518 VDD.n6517 3.1505
R8939 VDD.n6517 VDD.n6516 3.1505
R8940 VDD.n6515 VDD.n6514 3.1505
R8941 VDD.n6514 VDD.n6513 3.1505
R8942 VDD.n6512 VDD.n6511 3.1505
R8943 VDD.n6511 VDD.n6510 3.1505
R8944 VDD.n6509 VDD.n6508 3.1505
R8945 VDD.n6508 VDD.n6507 3.1505
R8946 VDD.n6505 VDD.n6504 3.1505
R8947 VDD.n6504 VDD.n6503 3.1505
R8948 VDD.n6502 VDD.n6501 3.1505
R8949 VDD.n6501 VDD.n6500 3.1505
R8950 VDD.n6499 VDD.n6498 3.1505
R8951 VDD.n6498 VDD.n6497 3.1505
R8952 VDD.n6495 VDD.n6494 3.1505
R8953 VDD.n6494 VDD.n6493 3.1505
R8954 VDD.n6492 VDD.n6491 3.1505
R8955 VDD.n6491 VDD.n6490 3.1505
R8956 VDD.n6489 VDD.n6488 3.1505
R8957 VDD.n6488 VDD.n6487 3.1505
R8958 VDD.n6485 VDD.n6484 3.1505
R8959 VDD.n6484 VDD.n6483 3.1505
R8960 VDD.n6482 VDD.n6481 3.1505
R8961 VDD.n6481 VDD.n6480 3.1505
R8962 VDD.n6479 VDD.n6478 3.1505
R8963 VDD.n6478 VDD.n6477 3.1505
R8964 VDD.n6475 VDD.n6474 3.1505
R8965 VDD.n6474 VDD.n6473 3.1505
R8966 VDD.n6472 VDD.n6471 3.1505
R8967 VDD.n6471 VDD.n6470 3.1505
R8968 VDD.n6468 VDD.n6467 3.1505
R8969 VDD.n6467 VDD.n6466 3.1505
R8970 VDD.n6465 VDD.n6464 3.1505
R8971 VDD.n6464 VDD.n6463 3.1505
R8972 VDD.n6462 VDD.n6461 3.1505
R8973 VDD.n6461 VDD.n6460 3.1505
R8974 VDD.n6459 VDD.n6458 3.1505
R8975 VDD.n6458 VDD.n6457 3.1505
R8976 VDD.n737 VDD.n736 3.1505
R8977 VDD.n6851 VDD.n6850 3.1505
R8978 VDD.n6828 VDD.n6827 3.1505
R8979 VDD.n6825 VDD.n6824 3.1505
R8980 VDD.n6822 VDD.n6821 3.1505
R8981 VDD.n6819 VDD.n6818 3.1505
R8982 VDD.n6816 VDD.n6815 3.1505
R8983 VDD.n6813 VDD.n6812 3.1505
R8984 VDD.n6810 VDD.n6809 3.1505
R8985 VDD.n6807 VDD.n6806 3.1505
R8986 VDD.n6804 VDD.n6803 3.1505
R8987 VDD.n6801 VDD.n6800 3.1505
R8988 VDD.n6798 VDD.n6797 3.1505
R8989 VDD.n6795 VDD.n6794 3.1505
R8990 VDD.n6792 VDD.n6791 3.1505
R8991 VDD.n6789 VDD.n6788 3.1505
R8992 VDD.n6786 VDD.n6785 3.1505
R8993 VDD.n6783 VDD.n6782 3.1505
R8994 VDD.n6780 VDD.n6779 3.1505
R8995 VDD.n6777 VDD.n6776 3.1505
R8996 VDD.n6774 VDD.n6773 3.1505
R8997 VDD.n6771 VDD.n6770 3.1505
R8998 VDD.n6768 VDD.n6767 3.1505
R8999 VDD.n6765 VDD.n6764 3.1505
R9000 VDD.n6762 VDD.n6761 3.1505
R9001 VDD.n6759 VDD.n6758 3.1505
R9002 VDD.n6756 VDD.n6755 3.1505
R9003 VDD.n6753 VDD.n6752 3.1505
R9004 VDD.n6750 VDD.n6749 3.1505
R9005 VDD.n6748 VDD.n6747 3.1505
R9006 VDD.n6746 VDD.n6745 3.1505
R9007 VDD.n6744 VDD.n6743 3.1505
R9008 VDD.n6742 VDD.n6741 3.1505
R9009 VDD.n6740 VDD.n6739 3.1505
R9010 VDD.n6738 VDD.n6737 3.1505
R9011 VDD.n6736 VDD.n6735 3.1505
R9012 VDD.n6734 VDD.n6733 3.1505
R9013 VDD.n6732 VDD.n6731 3.1505
R9014 VDD.n6730 VDD.n6729 3.1505
R9015 VDD.n6728 VDD.n6727 3.1505
R9016 VDD.n6726 VDD.n6725 3.1505
R9017 VDD.n6724 VDD.n6723 3.1505
R9018 VDD.n6722 VDD.n6721 3.1505
R9019 VDD.n6720 VDD.n6719 3.1505
R9020 VDD.n6718 VDD.n6717 3.1505
R9021 VDD.n6716 VDD.n6715 3.1505
R9022 VDD.n6714 VDD.n6713 3.1505
R9023 VDD.n602 VDD.n601 3.1505
R9024 VDD.n712 VDD.n711 3.1505
R9025 VDD.n709 VDD.n708 3.1505
R9026 VDD.n706 VDD.n705 3.1505
R9027 VDD.n703 VDD.n702 3.1505
R9028 VDD.n700 VDD.n699 3.1505
R9029 VDD.n697 VDD.n696 3.1505
R9030 VDD.n694 VDD.n693 3.1505
R9031 VDD.n691 VDD.n690 3.1505
R9032 VDD.n688 VDD.n687 3.1505
R9033 VDD.n685 VDD.n684 3.1505
R9034 VDD.n682 VDD.n681 3.1505
R9035 VDD.n679 VDD.n678 3.1505
R9036 VDD.n676 VDD.n675 3.1505
R9037 VDD.n673 VDD.n672 3.1505
R9038 VDD.n670 VDD.n669 3.1505
R9039 VDD.n667 VDD.n666 3.1505
R9040 VDD.n664 VDD.n663 3.1505
R9041 VDD.n661 VDD.n660 3.1505
R9042 VDD.n658 VDD.n657 3.1505
R9043 VDD.n655 VDD.n654 3.1505
R9044 VDD.n652 VDD.n651 3.1505
R9045 VDD.n649 VDD.n648 3.1505
R9046 VDD.n646 VDD.n645 3.1505
R9047 VDD.n643 VDD.n642 3.1505
R9048 VDD.n640 VDD.n639 3.1505
R9049 VDD.n638 VDD.n637 3.1505
R9050 VDD.n636 VDD.n635 3.1505
R9051 VDD.n634 VDD.n633 3.1505
R9052 VDD.n632 VDD.n631 3.1505
R9053 VDD.n630 VDD.n629 3.1505
R9054 VDD.n628 VDD.n627 3.1505
R9055 VDD.n626 VDD.n625 3.1505
R9056 VDD.n624 VDD.n623 3.1505
R9057 VDD.n622 VDD.n621 3.1505
R9058 VDD.n620 VDD.n619 3.1505
R9059 VDD.n618 VDD.n617 3.1505
R9060 VDD.n616 VDD.n615 3.1505
R9061 VDD.n614 VDD.n613 3.1505
R9062 VDD.n612 VDD.n611 3.1505
R9063 VDD.n610 VDD.n609 3.1505
R9064 VDD.n608 VDD.n607 3.1505
R9065 VDD.n606 VDD.n605 3.1505
R9066 VDD.n604 VDD.n603 3.1505
R9067 VDD.n714 VDD.n713 3.1505
R9068 VDD.n1008 VDD.n1007 3.1505
R9069 VDD.n910 VDD.n909 3.1505
R9070 VDD.n912 VDD.n911 3.1505
R9071 VDD.n914 VDD.n913 3.1505
R9072 VDD.n916 VDD.n915 3.1505
R9073 VDD.n918 VDD.n917 3.1505
R9074 VDD.n920 VDD.n919 3.1505
R9075 VDD.n922 VDD.n921 3.1505
R9076 VDD.n924 VDD.n923 3.1505
R9077 VDD.n926 VDD.n925 3.1505
R9078 VDD.n928 VDD.n927 3.1505
R9079 VDD.n930 VDD.n929 3.1505
R9080 VDD.n932 VDD.n931 3.1505
R9081 VDD.n934 VDD.n933 3.1505
R9082 VDD.n936 VDD.n935 3.1505
R9083 VDD.n938 VDD.n937 3.1505
R9084 VDD.n940 VDD.n939 3.1505
R9085 VDD.n942 VDD.n941 3.1505
R9086 VDD.n944 VDD.n943 3.1505
R9087 VDD.n946 VDD.n945 3.1505
R9088 VDD.n948 VDD.n947 3.1505
R9089 VDD.n950 VDD.n949 3.1505
R9090 VDD.n952 VDD.n951 3.1505
R9091 VDD.n954 VDD.n953 3.1505
R9092 VDD.n956 VDD.n955 3.1505
R9093 VDD.n958 VDD.n957 3.1505
R9094 VDD.n960 VDD.n959 3.1505
R9095 VDD.n962 VDD.n961 3.1505
R9096 VDD.n964 VDD.n963 3.1505
R9097 VDD.n966 VDD.n965 3.1505
R9098 VDD.n968 VDD.n967 3.1505
R9099 VDD.n971 VDD.n970 3.1505
R9100 VDD.n973 VDD.n972 3.1505
R9101 VDD.n976 VDD.n975 3.1505
R9102 VDD.n978 VDD.n977 3.1505
R9103 VDD.n981 VDD.n980 3.1505
R9104 VDD.n983 VDD.n982 3.1505
R9105 VDD.n986 VDD.n985 3.1505
R9106 VDD.n988 VDD.n987 3.1505
R9107 VDD.n991 VDD.n990 3.1505
R9108 VDD.n993 VDD.n992 3.1505
R9109 VDD.n996 VDD.n995 3.1505
R9110 VDD.n998 VDD.n997 3.1505
R9111 VDD.n1001 VDD.n1000 3.1505
R9112 VDD.n1003 VDD.n1002 3.1505
R9113 VDD.n1006 VDD.n1005 3.1505
R9114 VDD.n908 VDD.n871 3.1505
R9115 VDD.n907 VDD.n906 3.1505
R9116 VDD.n905 VDD.n904 3.1505
R9117 VDD.n902 VDD.n901 3.1505
R9118 VDD.n900 VDD.n899 3.1505
R9119 VDD.n897 VDD.n896 3.1505
R9120 VDD.n895 VDD.n894 3.1505
R9121 VDD.n893 VDD.n892 3.1505
R9122 VDD.n890 VDD.n889 3.1505
R9123 VDD.n888 VDD.n887 3.1505
R9124 VDD.n886 VDD.n885 3.1505
R9125 VDD.n883 VDD.n882 3.1505
R9126 VDD.n881 VDD.n880 3.1505
R9127 VDD.n572 VDD.n571 3.1505
R9128 VDD.n574 VDD.n573 3.1505
R9129 VDD.n577 VDD.n576 3.1505
R9130 VDD.n579 VDD.n578 3.1505
R9131 VDD.n581 VDD.n580 3.1505
R9132 VDD.n584 VDD.n583 3.1505
R9133 VDD.n586 VDD.n585 3.1505
R9134 VDD.n588 VDD.n587 3.1505
R9135 VDD.n591 VDD.n590 3.1505
R9136 VDD.n593 VDD.n592 3.1505
R9137 VDD.n596 VDD.n595 3.1505
R9138 VDD.n598 VDD.n597 3.1505
R9139 VDD.n600 VDD.n599 3.1505
R9140 VDD.n6651 VDD.n6650 3.1505
R9141 VDD.n6654 VDD.n6653 3.1505
R9142 VDD.n6656 VDD.n6655 3.1505
R9143 VDD.n6659 VDD.n6658 3.1505
R9144 VDD.n6661 VDD.n6660 3.1505
R9145 VDD.n6663 VDD.n6662 3.1505
R9146 VDD.n6665 VDD.n6664 3.1505
R9147 VDD.n6667 VDD.n6666 3.1505
R9148 VDD.n6669 VDD.n6668 3.1505
R9149 VDD.n6671 VDD.n6670 3.1505
R9150 VDD.n6673 VDD.n6672 3.1505
R9151 VDD.n6675 VDD.n6674 3.1505
R9152 VDD.n6677 VDD.n6676 3.1505
R9153 VDD.n6679 VDD.n6678 3.1505
R9154 VDD.n6681 VDD.n6680 3.1505
R9155 VDD.n6683 VDD.n6682 3.1505
R9156 VDD.n6685 VDD.n6684 3.1505
R9157 VDD.n6687 VDD.n6686 3.1505
R9158 VDD.n6689 VDD.n6688 3.1505
R9159 VDD.n6691 VDD.n6690 3.1505
R9160 VDD.n6693 VDD.n6692 3.1505
R9161 VDD.n6695 VDD.n6694 3.1505
R9162 VDD.n6697 VDD.n6696 3.1505
R9163 VDD.n6699 VDD.n6698 3.1505
R9164 VDD.n6701 VDD.n6700 3.1505
R9165 VDD.n6705 VDD.n6704 3.1505
R9166 VDD.n6707 VDD.n6706 3.1505
R9167 VDD.n6710 VDD.n6709 3.1505
R9168 VDD.n6712 VDD.n6711 3.1505
R9169 VDD.n7640 VDD.n7639 3.1505
R9170 VDD.n7388 VDD.n7387 3.1505
R9171 VDD.n7565 VDD.n7564 3.1505
R9172 VDD.n7635 VDD.n7634 3.1505
R9173 VDD.n7632 VDD.n7631 3.1505
R9174 VDD.n7628 VDD.n7627 3.1505
R9175 VDD.n7626 VDD.n7625 3.1505
R9176 VDD.n7623 VDD.n7622 3.1505
R9177 VDD.n7621 VDD.n7620 3.1505
R9178 VDD.n7618 VDD.n7617 3.1505
R9179 VDD.n7616 VDD.n7615 3.1505
R9180 VDD.n7612 VDD.n7611 3.1505
R9181 VDD.n7610 VDD.n7609 3.1505
R9182 VDD.n7607 VDD.n7606 3.1505
R9183 VDD.n7604 VDD.n7603 3.1505
R9184 VDD.n7602 VDD.n7601 3.1505
R9185 VDD.n7600 VDD.n7599 3.1505
R9186 VDD.n7598 VDD.n7597 3.1505
R9187 VDD.n7596 VDD.n7595 3.1505
R9188 VDD.n7594 VDD.n7593 3.1505
R9189 VDD.n7591 VDD.n7590 3.1505
R9190 VDD.n7589 VDD.n7588 3.1505
R9191 VDD.n7587 VDD.n7586 3.1505
R9192 VDD.n7585 VDD.n7584 3.1505
R9193 VDD.n7582 VDD.n7581 3.1505
R9194 VDD.n7580 VDD.n7579 3.1505
R9195 VDD.n7578 VDD.n7577 3.1505
R9196 VDD.n7576 VDD.n7575 3.1505
R9197 VDD.n7574 VDD.n7573 3.1505
R9198 VDD.n7572 VDD.n7571 3.1505
R9199 VDD.n7569 VDD.n7568 3.1505
R9200 VDD.n7567 VDD.n7566 3.1505
R9201 VDD.n7637 VDD.n7636 3.1505
R9202 VDD.n7390 VDD.n7389 3.1505
R9203 VDD.n7394 VDD.n7392 3.1505
R9204 VDD.n7397 VDD.n7395 3.1505
R9205 VDD.n7400 VDD.n7398 3.1505
R9206 VDD.n7403 VDD.n7401 3.1505
R9207 VDD.n7406 VDD.n7404 3.1505
R9208 VDD.n7409 VDD.n7407 3.1505
R9209 VDD.n7413 VDD.n7410 3.1505
R9210 VDD.n7417 VDD.n7414 3.1505
R9211 VDD.n7421 VDD.n7418 3.1505
R9212 VDD.n7425 VDD.n7423 3.1505
R9213 VDD.n7423 VDD.n7422 3.1505
R9214 VDD.n7429 VDD.n7427 3.1505
R9215 VDD.n7427 VDD.n7426 3.1505
R9216 VDD.n7433 VDD.n7430 3.1505
R9217 VDD.n7437 VDD.n7435 3.1505
R9218 VDD.n7435 VDD.n7434 3.1505
R9219 VDD.n7441 VDD.n7439 3.1505
R9220 VDD.n7439 VDD.n7438 3.1505
R9221 VDD.n7445 VDD.n7443 3.1505
R9222 VDD.n7443 VDD.n7442 3.1505
R9223 VDD.n7449 VDD.n7447 3.1505
R9224 VDD.n7447 VDD.n7446 3.1505
R9225 VDD.n7453 VDD.n7450 3.1505
R9226 VDD.n7457 VDD.n7455 3.1505
R9227 VDD.n7455 VDD.n7454 3.1505
R9228 VDD.n7461 VDD.n7459 3.1505
R9229 VDD.n7459 VDD.n7458 3.1505
R9230 VDD.n7465 VDD.n7462 3.1505
R9231 VDD.n7469 VDD.n7467 3.1505
R9232 VDD.n7467 VDD.n7466 3.1505
R9233 VDD.n7473 VDD.n7471 3.1505
R9234 VDD.n7471 VDD.n7470 3.1505
R9235 VDD.n7477 VDD.n7475 3.1505
R9236 VDD.n7475 VDD.n7474 3.1505
R9237 VDD.n7481 VDD.n7479 3.1505
R9238 VDD.n7479 VDD.n7478 3.1505
R9239 VDD.n7485 VDD.n7482 3.1505
R9240 VDD.n7489 VDD.n7486 3.1505
R9241 VDD.n7493 VDD.n7491 3.1505
R9242 VDD.n7491 VDD.n7490 3.1505
R9243 VDD.n7497 VDD.n7495 3.1505
R9244 VDD.n7495 VDD.n7494 3.1505
R9245 VDD.n7501 VDD.n7499 3.1505
R9246 VDD.n7499 VDD.n7498 3.1505
R9247 VDD.n7505 VDD.n7503 3.1505
R9248 VDD.n7503 VDD.n7502 3.1505
R9249 VDD.n7509 VDD.n7506 3.1505
R9250 VDD.n7513 VDD.n7511 3.1505
R9251 VDD.n7511 VDD.n7510 3.1505
R9252 VDD.n7517 VDD.n7514 3.1505
R9253 VDD.n7521 VDD.n7518 3.1505
R9254 VDD.n7525 VDD.n7522 3.1505
R9255 VDD.n7529 VDD.n7526 3.1505
R9256 VDD.n7533 VDD.n7530 3.1505
R9257 VDD.n7537 VDD.n7535 3.1505
R9258 VDD.n7535 VDD.n7534 3.1505
R9259 VDD.n7386 VDD.n7385 3.1505
R9260 VDD.n7384 VDD.n7383 3.1505
R9261 VDD.n7381 VDD.n7380 3.1505
R9262 VDD.n7379 VDD.n7378 3.1505
R9263 VDD.n7377 VDD.n7376 3.1505
R9264 VDD.n7375 VDD.n7374 3.1505
R9265 VDD.n7373 VDD.n7372 3.1505
R9266 VDD.n7371 VDD.n7370 3.1505
R9267 VDD.n7368 VDD.n7367 3.1505
R9268 VDD.n7366 VDD.n7365 3.1505
R9269 VDD.n7364 VDD.n7363 3.1505
R9270 VDD.n7361 VDD.n7360 3.1505
R9271 VDD.n7359 VDD.n7358 3.1505
R9272 VDD.n7357 VDD.n7356 3.1505
R9273 VDD.n7355 VDD.n7354 3.1505
R9274 VDD.n7353 VDD.n7352 3.1505
R9275 VDD.n7351 VDD.n7350 3.1505
R9276 VDD.n7348 VDD.n7347 3.1505
R9277 VDD.n7346 VDD.n7345 3.1505
R9278 VDD.n7344 VDD.n7343 3.1505
R9279 VDD.n7342 VDD.n7341 3.1505
R9280 VDD.n7329 VDD.n7328 3.1505
R9281 VDD.n7327 VDD.n7326 3.1505
R9282 VDD.n7325 VDD.n7324 3.1505
R9283 VDD.n7323 VDD.n7322 3.1505
R9284 VDD.n7321 VDD.n7320 3.1505
R9285 VDD.n7319 VDD.n7318 3.1505
R9286 VDD.n7317 VDD.n7316 3.1505
R9287 VDD.n7315 VDD.n7314 3.1505
R9288 VDD.n7313 VDD.n7312 3.1505
R9289 VDD.n7311 VDD.n7310 3.1505
R9290 VDD.n7309 VDD.n7308 3.1505
R9291 VDD.n7307 VDD.n7306 3.1505
R9292 VDD.n7305 VDD.n7304 3.1505
R9293 VDD.n7303 VDD.n7302 3.1505
R9294 VDD.n7301 VDD.n7300 3.1505
R9295 VDD.n7299 VDD.n7298 3.1505
R9296 VDD.n7297 VDD.n7296 3.1505
R9297 VDD.n7295 VDD.n7294 3.1505
R9298 VDD.n7293 VDD.n7292 3.1505
R9299 VDD.n7291 VDD.n7290 3.1505
R9300 VDD.n7289 VDD.n7288 3.1505
R9301 VDD.n7287 VDD.n7286 3.1505
R9302 VDD.n7285 VDD.n7284 3.1505
R9303 VDD.n7283 VDD.n7282 3.1505
R9304 VDD.n7281 VDD.n7280 3.1505
R9305 VDD.n7539 VDD.n7538 3.1505
R9306 VDD.n7541 VDD.n7540 3.1505
R9307 VDD.n7543 VDD.n7542 3.1505
R9308 VDD.n7545 VDD.n7544 3.1505
R9309 VDD.n7547 VDD.n7546 3.1505
R9310 VDD.n7549 VDD.n7548 3.1505
R9311 VDD.n7551 VDD.n7550 3.1505
R9312 VDD.n7553 VDD.n7552 3.1505
R9313 VDD.n7555 VDD.n7554 3.1505
R9314 VDD.n7557 VDD.n7556 3.1505
R9315 VDD.n7559 VDD.n7558 3.1505
R9316 VDD.n7561 VDD.n7560 3.1505
R9317 VDD.n7563 VDD.n7562 3.1505
R9318 VDD.n7820 VDD.n7242 3.1505
R9319 VDD.n7819 VDD.n7818 3.1505
R9320 VDD.n7818 VDD.n7817 3.1505
R9321 VDD.n7816 VDD.n7815 3.1505
R9322 VDD.n7815 VDD.n7814 3.1505
R9323 VDD.n7813 VDD.n7812 3.1505
R9324 VDD.n7812 VDD.n7811 3.1505
R9325 VDD.n7810 VDD.n7809 3.1505
R9326 VDD.n7809 VDD.n7808 3.1505
R9327 VDD.n7807 VDD.n7806 3.1505
R9328 VDD.n7806 VDD.n7805 3.1505
R9329 VDD.n7804 VDD.n7803 3.1505
R9330 VDD.n7803 VDD.n7802 3.1505
R9331 VDD.n7801 VDD.n7800 3.1505
R9332 VDD.n7799 VDD.n7798 3.1505
R9333 VDD.n7797 VDD.n7796 3.1505
R9334 VDD.n7795 VDD.n7794 3.1505
R9335 VDD.n7793 VDD.n7792 3.1505
R9336 VDD.n7791 VDD.n7790 3.1505
R9337 VDD.n7789 VDD.n7788 3.1505
R9338 VDD.n7787 VDD.n7786 3.1505
R9339 VDD.n7785 VDD.n7784 3.1505
R9340 VDD.n7783 VDD.n7782 3.1505
R9341 VDD.n7781 VDD.n7780 3.1505
R9342 VDD.n7779 VDD.n7778 3.1505
R9343 VDD.n7777 VDD.n7776 3.1505
R9344 VDD.n7775 VDD.n7774 3.1505
R9345 VDD.n7773 VDD.n7772 3.1505
R9346 VDD.n7771 VDD.n7770 3.1505
R9347 VDD.n7769 VDD.n7768 3.1505
R9348 VDD.n7767 VDD.n7766 3.1505
R9349 VDD.n7765 VDD.n7764 3.1505
R9350 VDD.n7763 VDD.n7762 3.1505
R9351 VDD.n7761 VDD.n7760 3.1505
R9352 VDD.n7759 VDD.n7758 3.1505
R9353 VDD.n7757 VDD.n7756 3.1505
R9354 VDD.n7755 VDD.n7754 3.1505
R9355 VDD.n7753 VDD.n7752 3.1505
R9356 VDD.n7751 VDD.n7750 3.1505
R9357 VDD.n7749 VDD.n7748 3.1505
R9358 VDD.n7747 VDD.n7746 3.1505
R9359 VDD.n7745 VDD.n7744 3.1505
R9360 VDD.n7743 VDD.n7742 3.1505
R9361 VDD.n7741 VDD.n7740 3.1505
R9362 VDD.n7739 VDD.n7738 3.1505
R9363 VDD.n7737 VDD.n7243 3.1505
R9364 VDD.n7736 VDD.n7735 3.1505
R9365 VDD.n7734 VDD.n7733 3.1505
R9366 VDD.n7731 VDD.n7730 3.1505
R9367 VDD.n7729 VDD.n7728 3.1505
R9368 VDD.n7727 VDD.n7726 3.1505
R9369 VDD.n7725 VDD.n7724 3.1505
R9370 VDD.n7723 VDD.n7722 3.1505
R9371 VDD.n7721 VDD.n7720 3.1505
R9372 VDD.n7718 VDD.n7717 3.1505
R9373 VDD.n7716 VDD.n7715 3.1505
R9374 VDD.n7714 VDD.n7713 3.1505
R9375 VDD.n7712 VDD.n7711 3.1505
R9376 VDD.n7709 VDD.n7708 3.1505
R9377 VDD.n7707 VDD.n7706 3.1505
R9378 VDD.n7705 VDD.n7704 3.1505
R9379 VDD.n7703 VDD.n7702 3.1505
R9380 VDD.n7701 VDD.n7700 3.1505
R9381 VDD.n7699 VDD.n7698 3.1505
R9382 VDD.n7696 VDD.n7695 3.1505
R9383 VDD.n7694 VDD.n7693 3.1505
R9384 VDD.n7692 VDD.n7691 3.1505
R9385 VDD.n7688 VDD.n7687 3.1505
R9386 VDD.n7686 VDD.n7685 3.1505
R9387 VDD.n7683 VDD.n7682 3.1505
R9388 VDD.n7681 VDD.n7680 3.1505
R9389 VDD.n7678 VDD.n7677 3.1505
R9390 VDD.n7676 VDD.n7675 3.1505
R9391 VDD.n7672 VDD.n7671 3.1505
R9392 VDD.n7670 VDD.n7669 3.1505
R9393 VDD.n7667 VDD.n7666 3.1505
R9394 VDD.n7665 VDD.n7664 3.1505
R9395 VDD.n7394 VDD.n7393 3.1505
R9396 VDD.n7397 VDD.n7396 3.1505
R9397 VDD.n7400 VDD.n7399 3.1505
R9398 VDD.n7403 VDD.n7402 3.1505
R9399 VDD.n7406 VDD.n7405 3.1505
R9400 VDD.n7409 VDD.n7408 3.1505
R9401 VDD.n7413 VDD.n7412 3.1505
R9402 VDD.n7412 VDD.n7411 3.1505
R9403 VDD.n7417 VDD.n7416 3.1505
R9404 VDD.n7416 VDD.n7415 3.1505
R9405 VDD.n7421 VDD.n7420 3.1505
R9406 VDD.n7420 VDD.n7419 3.1505
R9407 VDD.n7425 VDD.n7424 3.1505
R9408 VDD.n7429 VDD.n7428 3.1505
R9409 VDD.n7433 VDD.n7432 3.1505
R9410 VDD.n7432 VDD.n7431 3.1505
R9411 VDD.n7437 VDD.n7436 3.1505
R9412 VDD.n7441 VDD.n7440 3.1505
R9413 VDD.n7445 VDD.n7444 3.1505
R9414 VDD.n7449 VDD.n7448 3.1505
R9415 VDD.n7453 VDD.n7452 3.1505
R9416 VDD.n7452 VDD.n7451 3.1505
R9417 VDD.n7457 VDD.n7456 3.1505
R9418 VDD.n7461 VDD.n7460 3.1505
R9419 VDD.n7465 VDD.n7464 3.1505
R9420 VDD.n7464 VDD.n7463 3.1505
R9421 VDD.n7469 VDD.n7468 3.1505
R9422 VDD.n7473 VDD.n7472 3.1505
R9423 VDD.n7477 VDD.n7476 3.1505
R9424 VDD.n7481 VDD.n7480 3.1505
R9425 VDD.n7485 VDD.n7484 3.1505
R9426 VDD.n7484 VDD.n7483 3.1505
R9427 VDD.n7489 VDD.n7488 3.1505
R9428 VDD.n7488 VDD.n7487 3.1505
R9429 VDD.n7493 VDD.n7492 3.1505
R9430 VDD.n7497 VDD.n7496 3.1505
R9431 VDD.n7501 VDD.n7500 3.1505
R9432 VDD.n7505 VDD.n7504 3.1505
R9433 VDD.n7509 VDD.n7508 3.1505
R9434 VDD.n7508 VDD.n7507 3.1505
R9435 VDD.n7513 VDD.n7512 3.1505
R9436 VDD.n7517 VDD.n7516 3.1505
R9437 VDD.n7516 VDD.n7515 3.1505
R9438 VDD.n7521 VDD.n7520 3.1505
R9439 VDD.n7520 VDD.n7519 3.1505
R9440 VDD.n7525 VDD.n7524 3.1505
R9441 VDD.n7524 VDD.n7523 3.1505
R9442 VDD.n7529 VDD.n7528 3.1505
R9443 VDD.n7528 VDD.n7527 3.1505
R9444 VDD.n7533 VDD.n7532 3.1505
R9445 VDD.n7532 VDD.n7531 3.1505
R9446 VDD.n7537 VDD.n7536 3.1505
R9447 VDD.n7279 VDD.n7278 3.1505
R9448 VDD.n7844 VDD.n7843 3.1505
R9449 VDD.n7840 VDD.n7839 3.1505
R9450 VDD.n7838 VDD.n7837 3.1505
R9451 VDD.n7835 VDD.n7834 3.1505
R9452 VDD.n7833 VDD.n7832 3.1505
R9453 VDD.n7830 VDD.n7829 3.1505
R9454 VDD.n7828 VDD.n7827 3.1505
R9455 VDD.n7825 VDD.n7824 3.1505
R9456 VDD.n7823 VDD.n7822 3.1505
R9457 VDD.n7846 VDD.n7845 3.1505
R9458 VDD.n7849 VDD.n7848 3.1505
R9459 VDD.n7241 VDD.n7240 3.1505
R9460 VDD.n7245 VDD.n7244 3.1505
R9461 VDD.n7248 VDD.n7247 3.1505
R9462 VDD.n7251 VDD.n7250 3.1505
R9463 VDD.n7254 VDD.n7253 3.1505
R9464 VDD.n7256 VDD.n7255 3.1505
R9465 VDD.n7260 VDD.n7259 3.1505
R9466 VDD.n7262 VDD.n7261 3.1505
R9467 VDD.n7264 VDD.n7263 3.1505
R9468 VDD.n7266 VDD.n7265 3.1505
R9469 VDD.n7268 VDD.n7267 3.1505
R9470 VDD.n7270 VDD.n7269 3.1505
R9471 VDD.n7273 VDD.n7272 3.1505
R9472 VDD.n7275 VDD.n7274 3.1505
R9473 VDD.n7277 VDD.n7276 3.1505
R9474 VDD.n7886 VDD.n7884 3.1505
R9475 VDD.n7886 VDD.n7885 3.1505
R9476 VDD.n138 VDD.n137 3.1505
R9477 VDD.n46 VDD.n45 3.1505
R9478 VDD.n48 VDD.n47 3.1505
R9479 VDD.n50 VDD.n49 3.1505
R9480 VDD.n52 VDD.n51 3.1505
R9481 VDD.n54 VDD.n53 3.1505
R9482 VDD.n56 VDD.n55 3.1505
R9483 VDD.n58 VDD.n57 3.1505
R9484 VDD.n60 VDD.n59 3.1505
R9485 VDD.n62 VDD.n61 3.1505
R9486 VDD.n64 VDD.n63 3.1505
R9487 VDD.n66 VDD.n65 3.1505
R9488 VDD.n68 VDD.n67 3.1505
R9489 VDD.n70 VDD.n69 3.1505
R9490 VDD.n73 VDD.n72 3.1505
R9491 VDD.n76 VDD.n75 3.1505
R9492 VDD.n79 VDD.n78 3.1505
R9493 VDD.n82 VDD.n81 3.1505
R9494 VDD.n85 VDD.n84 3.1505
R9495 VDD.n88 VDD.n87 3.1505
R9496 VDD.n91 VDD.n90 3.1505
R9497 VDD.n94 VDD.n93 3.1505
R9498 VDD.n97 VDD.n96 3.1505
R9499 VDD.n100 VDD.n99 3.1505
R9500 VDD.n103 VDD.n102 3.1505
R9501 VDD.n106 VDD.n105 3.1505
R9502 VDD.n109 VDD.n108 3.1505
R9503 VDD.n112 VDD.n111 3.1505
R9504 VDD.n115 VDD.n114 3.1505
R9505 VDD.n118 VDD.n117 3.1505
R9506 VDD.n121 VDD.n120 3.1505
R9507 VDD.n124 VDD.n123 3.1505
R9508 VDD.n127 VDD.n126 3.1505
R9509 VDD.n130 VDD.n129 3.1505
R9510 VDD.n133 VDD.n132 3.1505
R9511 VDD.n136 VDD.n135 3.1505
R9512 VDD.n139 VDD.n42 3.1505
R9513 VDD.n142 VDD.n141 3.1505
R9514 VDD.n141 VDD.n140 3.1505
R9515 VDD.n146 VDD.n145 3.1505
R9516 VDD.n145 VDD.n144 3.1505
R9517 VDD.n149 VDD.n148 3.1505
R9518 VDD.n148 VDD.n147 3.1505
R9519 VDD.n153 VDD.n152 3.1505
R9520 VDD.n152 VDD.n151 3.1505
R9521 VDD.n156 VDD.n155 3.1505
R9522 VDD.n155 VDD.n154 3.1505
R9523 VDD.n159 VDD.n158 3.1505
R9524 VDD.n158 VDD.n157 3.1505
R9525 VDD.n162 VDD.n161 3.1505
R9526 VDD.n161 VDD.n160 3.1505
R9527 VDD.n165 VDD.n164 3.1505
R9528 VDD.n164 VDD.n163 3.1505
R9529 VDD.n168 VDD.n167 3.1505
R9530 VDD.n167 VDD.n166 3.1505
R9531 VDD.n171 VDD.n170 3.1505
R9532 VDD.n170 VDD.n169 3.1505
R9533 VDD.n174 VDD.n173 3.1505
R9534 VDD.n173 VDD.n172 3.1505
R9535 VDD.n177 VDD.n176 3.1505
R9536 VDD.n176 VDD.n175 3.1505
R9537 VDD.n180 VDD.n179 3.1505
R9538 VDD.n179 VDD.n178 3.1505
R9539 VDD.n183 VDD.n182 3.1505
R9540 VDD.n182 VDD.n181 3.1505
R9541 VDD.n186 VDD.n185 3.1505
R9542 VDD.n185 VDD.n184 3.1505
R9543 VDD.n189 VDD.n188 3.1505
R9544 VDD.n188 VDD.n187 3.1505
R9545 VDD.n192 VDD.n191 3.1505
R9546 VDD.n191 VDD.n190 3.1505
R9547 VDD.n195 VDD.n194 3.1505
R9548 VDD.n194 VDD.n193 3.1505
R9549 VDD.n198 VDD.n197 3.1505
R9550 VDD.n197 VDD.n196 3.1505
R9551 VDD.n202 VDD.n201 3.1505
R9552 VDD.n201 VDD.n200 3.1505
R9553 VDD.n205 VDD.n204 3.1505
R9554 VDD.n204 VDD.n203 3.1505
R9555 VDD.n209 VDD.n208 3.1505
R9556 VDD.n208 VDD.n207 3.1505
R9557 VDD.n211 VDD.n210 3.1505
R9558 VDD.n8215 VDD.n8214 3.1505
R9559 VDD.n6979 VDD.n6978 3.1505
R9560 VDD.n6965 VDD.n6964 3.1505
R9561 VDD.n6962 VDD.n6961 3.1505
R9562 VDD.n6959 VDD.n6958 3.1505
R9563 VDD.n6956 VDD.n6955 3.1505
R9564 VDD.n6953 VDD.n6952 3.1505
R9565 VDD.n6950 VDD.n6949 3.1505
R9566 VDD.n6947 VDD.n6946 3.1505
R9567 VDD.n6944 VDD.n6943 3.1505
R9568 VDD.n6941 VDD.n6940 3.1505
R9569 VDD.n6938 VDD.n6937 3.1505
R9570 VDD.n6935 VDD.n6934 3.1505
R9571 VDD.n6932 VDD.n6931 3.1505
R9572 VDD.n6929 VDD.n6928 3.1505
R9573 VDD.n6926 VDD.n6925 3.1505
R9574 VDD.n6923 VDD.n6922 3.1505
R9575 VDD.n6920 VDD.n6919 3.1505
R9576 VDD.n6917 VDD.n6916 3.1505
R9577 VDD.n6914 VDD.n6913 3.1505
R9578 VDD.n6911 VDD.n6910 3.1505
R9579 VDD.n6908 VDD.n6907 3.1505
R9580 VDD.n6905 VDD.n6904 3.1505
R9581 VDD.n6902 VDD.n6901 3.1505
R9582 VDD.n6899 VDD.n6898 3.1505
R9583 VDD.n6896 VDD.n6895 3.1505
R9584 VDD.n6893 VDD.n6892 3.1505
R9585 VDD.n6890 VDD.n6889 3.1505
R9586 VDD.n6887 VDD.n6886 3.1505
R9587 VDD.n6885 VDD.n6884 3.1505
R9588 VDD.n6883 VDD.n6882 3.1505
R9589 VDD.n6881 VDD.n6880 3.1505
R9590 VDD.n6879 VDD.n6878 3.1505
R9591 VDD.n6877 VDD.n6876 3.1505
R9592 VDD.n6875 VDD.n6874 3.1505
R9593 VDD.n6873 VDD.n6872 3.1505
R9594 VDD.n6871 VDD.n6870 3.1505
R9595 VDD.n6869 VDD.n6868 3.1505
R9596 VDD.n44 VDD.n43 3.1505
R9597 VDD.n8251 VDD.n7238 3.1505
R9598 VDD.n8285 VDD.n8284 3.1505
R9599 VDD.n8283 VDD.n8282 3.1505
R9600 VDD.n8280 VDD.n8279 3.1505
R9601 VDD.n8278 VDD.n8277 3.1505
R9602 VDD.n8275 VDD.n8274 3.1505
R9603 VDD.n8273 VDD.n8272 3.1505
R9604 VDD.n8270 VDD.n8269 3.1505
R9605 VDD.n8268 VDD.n8267 3.1505
R9606 VDD.n8265 VDD.n8264 3.1505
R9607 VDD.n8263 VDD.n8262 3.1505
R9608 VDD.n8260 VDD.n8259 3.1505
R9609 VDD.n8258 VDD.n8257 3.1505
R9610 VDD.n8255 VDD.n8254 3.1505
R9611 VDD.n8253 VDD.n8252 3.1505
R9612 VDD.n8250 VDD.n8249 3.1505
R9613 VDD.n8247 VDD.n8246 3.1505
R9614 VDD.n8245 VDD.n8244 3.1505
R9615 VDD.n8243 VDD.n8242 3.1505
R9616 VDD.n8241 VDD.n8240 3.1505
R9617 VDD.n8239 VDD.n8238 3.1505
R9618 VDD.n8237 VDD.n8236 3.1505
R9619 VDD.n8235 VDD.n8234 3.1505
R9620 VDD.n8233 VDD.n8232 3.1505
R9621 VDD.n8231 VDD.n8230 3.1505
R9622 VDD.n8229 VDD.n8228 3.1505
R9623 VDD.n8227 VDD.n8226 3.1505
R9624 VDD.n8225 VDD.n8224 3.1505
R9625 VDD.n8223 VDD.n8222 3.1505
R9626 VDD.n8221 VDD.n8220 3.1505
R9627 VDD.n8219 VDD.n8218 3.1505
R9628 VDD.n8217 VDD.n8216 3.1505
R9629 VDD.n7085 VDD.n7084 3.1505
R9630 VDD.n7089 VDD.n7088 3.1505
R9631 VDD.n7091 VDD.n7090 3.1505
R9632 VDD.n7093 VDD.n7092 3.1505
R9633 VDD.n7095 VDD.n7094 3.1505
R9634 VDD.n7097 VDD.n7096 3.1505
R9635 VDD.n7099 VDD.n7098 3.1505
R9636 VDD.n7101 VDD.n7100 3.1505
R9637 VDD.n7103 VDD.n7102 3.1505
R9638 VDD.n7105 VDD.n7104 3.1505
R9639 VDD.n7107 VDD.n7106 3.1505
R9640 VDD.n7109 VDD.n7108 3.1505
R9641 VDD.n7111 VDD.n7110 3.1505
R9642 VDD.n7113 VDD.n7112 3.1505
R9643 VDD.n7115 VDD.n7114 3.1505
R9644 VDD.n7117 VDD.n7116 3.1505
R9645 VDD.n7119 VDD.n7118 3.1505
R9646 VDD.n7121 VDD.n7120 3.1505
R9647 VDD.n7123 VDD.n7122 3.1505
R9648 VDD.n7125 VDD.n7124 3.1505
R9649 VDD.n7128 VDD.n7127 3.1505
R9650 VDD.n7130 VDD.n7129 3.1505
R9651 VDD.n7133 VDD.n7132 3.1505
R9652 VDD.n7135 VDD.n7134 3.1505
R9653 VDD.n7138 VDD.n7137 3.1505
R9654 VDD.n7140 VDD.n7139 3.1505
R9655 VDD.n7143 VDD.n7142 3.1505
R9656 VDD.n7145 VDD.n7144 3.1505
R9657 VDD.n7148 VDD.n7147 3.1505
R9658 VDD.n7150 VDD.n7149 3.1505
R9659 VDD.n7153 VDD.n7152 3.1505
R9660 VDD.n7155 VDD.n7154 3.1505
R9661 VDD.n7158 VDD.n7157 3.1505
R9662 VDD.n7160 VDD.n7159 3.1505
R9663 VDD.n7163 VDD.n7162 3.1505
R9664 VDD.n7165 VDD.n7164 3.1505
R9665 VDD.n7087 VDD.n7086 3.1505
R9666 VDD.n215 VDD.n214 3.1505
R9667 VDD.n217 VDD.n216 3.1505
R9668 VDD.n219 VDD.n218 3.1505
R9669 VDD.n221 VDD.n220 3.1505
R9670 VDD.n223 VDD.n222 3.1505
R9671 VDD.n225 VDD.n224 3.1505
R9672 VDD.n227 VDD.n226 3.1505
R9673 VDD.n229 VDD.n228 3.1505
R9674 VDD.n231 VDD.n230 3.1505
R9675 VDD.n233 VDD.n232 3.1505
R9676 VDD.n235 VDD.n234 3.1505
R9677 VDD.n237 VDD.n236 3.1505
R9678 VDD.n239 VDD.n238 3.1505
R9679 VDD.n241 VDD.n240 3.1505
R9680 VDD.n243 VDD.n242 3.1505
R9681 VDD.n245 VDD.n244 3.1505
R9682 VDD.n248 VDD.n247 3.1505
R9683 VDD.n250 VDD.n249 3.1505
R9684 VDD.n253 VDD.n252 3.1505
R9685 VDD.n255 VDD.n254 3.1505
R9686 VDD.n258 VDD.n257 3.1505
R9687 VDD.n260 VDD.n259 3.1505
R9688 VDD.n263 VDD.n262 3.1505
R9689 VDD.n265 VDD.n264 3.1505
R9690 VDD.n268 VDD.n267 3.1505
R9691 VDD.n270 VDD.n269 3.1505
R9692 VDD.n273 VDD.n272 3.1505
R9693 VDD.n275 VDD.n274 3.1505
R9694 VDD.n278 VDD.n277 3.1505
R9695 VDD.n280 VDD.n279 3.1505
R9696 VDD.n283 VDD.n282 3.1505
R9697 VDD.n285 VDD.n284 3.1505
R9698 VDD.n288 VDD.n287 3.1505
R9699 VDD.n290 VDD.n289 3.1505
R9700 VDD.n302 VDD.n301 3.1505
R9701 VDD.n213 VDD.n212 3.1505
R9702 VDD.n7179 VDD.n7178 3.1505
R9703 VDD.n7182 VDD.n7181 3.1505
R9704 VDD.n7181 VDD.n7180 3.1505
R9705 VDD.n7185 VDD.n7184 3.1505
R9706 VDD.n7184 VDD.n7183 3.1505
R9707 VDD.n7188 VDD.n7187 3.1505
R9708 VDD.n7187 VDD.n7186 3.1505
R9709 VDD.n7192 VDD.n7191 3.1505
R9710 VDD.n7191 VDD.n7190 3.1505
R9711 VDD.n7195 VDD.n7194 3.1505
R9712 VDD.n7194 VDD.n7193 3.1505
R9713 VDD.n7198 VDD.n7197 3.1505
R9714 VDD.n7197 VDD.n7196 3.1505
R9715 VDD.n7202 VDD.n7201 3.1505
R9716 VDD.n7201 VDD.n7200 3.1505
R9717 VDD.n7205 VDD.n7204 3.1505
R9718 VDD.n7204 VDD.n7203 3.1505
R9719 VDD.n7208 VDD.n7207 3.1505
R9720 VDD.n7207 VDD.n7206 3.1505
R9721 VDD.n7211 VDD.n7210 3.1505
R9722 VDD.n7210 VDD.n7209 3.1505
R9723 VDD.n7214 VDD.n7213 3.1505
R9724 VDD.n7213 VDD.n7212 3.1505
R9725 VDD.n7217 VDD.n7216 3.1505
R9726 VDD.n7216 VDD.n7215 3.1505
R9727 VDD.n7220 VDD.n7219 3.1505
R9728 VDD.n7219 VDD.n7218 3.1505
R9729 VDD.n7223 VDD.n7222 3.1505
R9730 VDD.n7222 VDD.n7221 3.1505
R9731 VDD.n7226 VDD.n7225 3.1505
R9732 VDD.n7225 VDD.n7224 3.1505
R9733 VDD.n7229 VDD.n7228 3.1505
R9734 VDD.n7228 VDD.n7227 3.1505
R9735 VDD VDD.n8347 3.1505
R9736 VDD.n8347 VDD.n8346 3.1505
R9737 VDD.n8345 VDD.n8344 3.1505
R9738 VDD.n8344 VDD.n8343 3.1505
R9739 VDD.n8342 VDD.n8341 3.1505
R9740 VDD.n8341 VDD.n8340 3.1505
R9741 VDD.n8339 VDD.n8338 3.1505
R9742 VDD.n8338 VDD.n8337 3.1505
R9743 VDD.n8336 VDD.n8335 3.1505
R9744 VDD.n8335 VDD.n8334 3.1505
R9745 VDD.n8333 VDD.n8332 3.1505
R9746 VDD.n8332 VDD.n8331 3.1505
R9747 VDD.n8330 VDD.n8329 3.1505
R9748 VDD.n8329 VDD.n8328 3.1505
R9749 VDD.n8327 VDD.n8326 3.1505
R9750 VDD.n8326 VDD.n8325 3.1505
R9751 VDD.n8316 VDD.n8315 3.1505
R9752 VDD.n8315 VDD.n8314 3.1505
R9753 VDD.n8313 VDD.n8312 3.1505
R9754 VDD.n8312 VDD.n8311 3.1505
R9755 VDD.n8309 VDD.n8308 3.1505
R9756 VDD.n8308 VDD.n8307 3.1505
R9757 VDD.n8306 VDD.n8305 3.1505
R9758 VDD.n8305 VDD.n8304 3.1505
R9759 VDD.n8303 VDD.n8302 3.1505
R9760 VDD.n8302 VDD.n8301 3.1505
R9761 VDD.n8300 VDD.n8299 3.1505
R9762 VDD.n8299 VDD.n8298 3.1505
R9763 VDD.n8297 VDD.n8296 3.1505
R9764 VDD.n532 VDD.n531 3.1505
R9765 VDD.n530 VDD.n529 3.1505
R9766 VDD.n527 VDD.n526 3.1505
R9767 VDD.n525 VDD.n524 3.1505
R9768 VDD.n522 VDD.n521 3.1505
R9769 VDD.n520 VDD.n519 3.1505
R9770 VDD.n517 VDD.n516 3.1505
R9771 VDD.n515 VDD.n514 3.1505
R9772 VDD.n512 VDD.n511 3.1505
R9773 VDD.n510 VDD.n509 3.1505
R9774 VDD.n507 VDD.n506 3.1505
R9775 VDD.n505 VDD.n504 3.1505
R9776 VDD.n502 VDD.n501 3.1505
R9777 VDD.n500 VDD.n499 3.1505
R9778 VDD.n497 VDD.n496 3.1505
R9779 VDD.n495 VDD.n494 3.1505
R9780 VDD.n492 VDD.n491 3.1505
R9781 VDD.n490 VDD.n489 3.1505
R9782 VDD.n487 VDD.n486 3.1505
R9783 VDD.n485 VDD.n484 3.1505
R9784 VDD.n482 VDD.n481 3.1505
R9785 VDD.n480 VDD.n479 3.1505
R9786 VDD.n477 VDD.n476 3.1505
R9787 VDD.n475 VDD.n474 3.1505
R9788 VDD.n473 VDD.n472 3.1505
R9789 VDD.n471 VDD.n470 3.1505
R9790 VDD.n469 VDD.n468 3.1505
R9791 VDD.n467 VDD.n466 3.1505
R9792 VDD.n465 VDD.n464 3.1505
R9793 VDD.n463 VDD.n462 3.1505
R9794 VDD.n461 VDD.n460 3.1505
R9795 VDD.n459 VDD.n458 3.1505
R9796 VDD.n457 VDD.n456 3.1505
R9797 VDD.n455 VDD.n454 3.1505
R9798 VDD.n8109 VDD.n8108 3.1505
R9799 VDD.n8032 VDD.n8031 3.1505
R9800 VDD.n8104 VDD.n8103 3.1505
R9801 VDD.n8102 VDD.n8101 3.1505
R9802 VDD.n8099 VDD.n8098 3.1505
R9803 VDD.n8097 VDD.n8096 3.1505
R9804 VDD.n8094 VDD.n8093 3.1505
R9805 VDD.n8092 VDD.n8091 3.1505
R9806 VDD.n8089 VDD.n8088 3.1505
R9807 VDD.n8087 VDD.n8086 3.1505
R9808 VDD.n8084 VDD.n8083 3.1505
R9809 VDD.n8082 VDD.n8081 3.1505
R9810 VDD.n8079 VDD.n8078 3.1505
R9811 VDD.n8077 VDD.n8076 3.1505
R9812 VDD.n8074 VDD.n8073 3.1505
R9813 VDD.n8072 VDD.n8071 3.1505
R9814 VDD.n8069 VDD.n8068 3.1505
R9815 VDD.n8067 VDD.n8066 3.1505
R9816 VDD.n8064 VDD.n8063 3.1505
R9817 VDD.n8062 VDD.n8061 3.1505
R9818 VDD.n8059 VDD.n8058 3.1505
R9819 VDD.n8057 VDD.n8056 3.1505
R9820 VDD.n8054 VDD.n8053 3.1505
R9821 VDD.n8052 VDD.n8051 3.1505
R9822 VDD.n8050 VDD.n8049 3.1505
R9823 VDD.n8048 VDD.n8047 3.1505
R9824 VDD.n8046 VDD.n8045 3.1505
R9825 VDD.n8044 VDD.n8043 3.1505
R9826 VDD.n8042 VDD.n8041 3.1505
R9827 VDD.n8040 VDD.n8039 3.1505
R9828 VDD.n8038 VDD.n8037 3.1505
R9829 VDD.n8036 VDD.n8035 3.1505
R9830 VDD.n8034 VDD.n8033 3.1505
R9831 VDD.n8107 VDD.n8106 3.1505
R9832 VDD.n8029 VDD.n8028 3.1505
R9833 VDD.n450 VDD.n449 3.1505
R9834 VDD.n448 VDD.n447 3.1505
R9835 VDD.n446 VDD.n445 3.1505
R9836 VDD.n443 VDD.n442 3.1505
R9837 VDD.n441 VDD.n440 3.1505
R9838 VDD.n438 VDD.n437 3.1505
R9839 VDD.n436 VDD.n435 3.1505
R9840 VDD.n434 VDD.n433 3.1505
R9841 VDD.n432 VDD.n431 3.1505
R9842 VDD.n430 VDD.n429 3.1505
R9843 VDD.n428 VDD.n427 3.1505
R9844 VDD.n426 VDD.n425 3.1505
R9845 VDD.n424 VDD.n423 3.1505
R9846 VDD.n422 VDD.n421 3.1505
R9847 VDD.n420 VDD.n419 3.1505
R9848 VDD.n418 VDD.n417 3.1505
R9849 VDD.n416 VDD.n415 3.1505
R9850 VDD.n414 VDD.n413 3.1505
R9851 VDD.n412 VDD.n411 3.1505
R9852 VDD.n410 VDD.n409 3.1505
R9853 VDD.n7982 VDD.n7981 3.1505
R9854 VDD.n7984 VDD.n7983 3.1505
R9855 VDD.n7986 VDD.n7985 3.1505
R9856 VDD.n7988 VDD.n7987 3.1505
R9857 VDD.n7990 VDD.n7989 3.1505
R9858 VDD.n7992 VDD.n7991 3.1505
R9859 VDD.n7994 VDD.n7993 3.1505
R9860 VDD.n7996 VDD.n7995 3.1505
R9861 VDD.n7998 VDD.n7997 3.1505
R9862 VDD.n8000 VDD.n7999 3.1505
R9863 VDD.n8002 VDD.n8001 3.1505
R9864 VDD.n8004 VDD.n8003 3.1505
R9865 VDD.n8006 VDD.n8005 3.1505
R9866 VDD.n8008 VDD.n8007 3.1505
R9867 VDD.n8010 VDD.n8009 3.1505
R9868 VDD.n8012 VDD.n8011 3.1505
R9869 VDD.n8014 VDD.n8013 3.1505
R9870 VDD.n8018 VDD.n8017 3.1505
R9871 VDD.n8020 VDD.n8019 3.1505
R9872 VDD.n8023 VDD.n8022 3.1505
R9873 VDD.n8025 VDD.n8024 3.1505
R9874 VDD.n8027 VDD.n8026 3.1505
R9875 VDD.n452 VDD.n451 3.1505
R9876 VDD.n8118 VDD.n8117 3.1505
R9877 VDD.n544 VDD.n540 3.1505
R9878 VDD.n543 VDD.n542 3.1505
R9879 VDD.n542 VDD.n541 3.1505
R9880 VDD.n323 VDD.n322 3.1505
R9881 VDD.n322 VDD.n321 3.1505
R9882 VDD.n326 VDD.n325 3.1505
R9883 VDD.n325 VDD.n324 3.1505
R9884 VDD.n329 VDD.n328 3.1505
R9885 VDD.n328 VDD.n327 3.1505
R9886 VDD.n333 VDD.n332 3.1505
R9887 VDD.n332 VDD.n331 3.1505
R9888 VDD.n336 VDD.n335 3.1505
R9889 VDD.n335 VDD.n334 3.1505
R9890 VDD.n340 VDD.n339 3.1505
R9891 VDD.n339 VDD.n338 3.1505
R9892 VDD.n344 VDD.n343 3.1505
R9893 VDD.n343 VDD.n342 3.1505
R9894 VDD.n347 VDD.n346 3.1505
R9895 VDD.n346 VDD.n345 3.1505
R9896 VDD.n350 VDD.n349 3.1505
R9897 VDD.n349 VDD.n348 3.1505
R9898 VDD.n389 VDD.n388 3.1505
R9899 VDD.n388 VDD.n387 3.1505
R9900 VDD.n386 VDD.n385 3.1505
R9901 VDD.n385 VDD.n384 3.1505
R9902 VDD.n382 VDD.n381 3.1505
R9903 VDD.n381 VDD.n380 3.1505
R9904 VDD.n379 VDD.n378 3.1505
R9905 VDD.n378 VDD.n377 3.1505
R9906 VDD.n376 VDD.n375 3.1505
R9907 VDD.n375 VDD.n374 3.1505
R9908 VDD.n373 VDD.n372 3.1505
R9909 VDD.n372 VDD.n371 3.1505
R9910 VDD.n369 VDD.n368 3.1505
R9911 VDD.n368 VDD.n367 3.1505
R9912 VDD.n366 VDD.n365 3.1505
R9913 VDD.n365 VDD.n364 3.1505
R9914 VDD.n363 VDD.n362 3.1505
R9915 VDD.n362 VDD.n361 3.1505
R9916 VDD.n360 VDD.n359 3.1505
R9917 VDD.n359 VDD.n358 3.1505
R9918 VDD.n357 VDD.n356 3.1505
R9919 VDD.n356 VDD.n355 3.1505
R9920 VDD.n7915 VDD.n7914 3.1505
R9921 VDD.n7914 VDD.n7913 3.1505
R9922 VDD.n7918 VDD.n7917 3.1505
R9923 VDD.n7917 VDD.n7916 3.1505
R9924 VDD.n7921 VDD.n7920 3.1505
R9925 VDD.n7920 VDD.n7919 3.1505
R9926 VDD.n7924 VDD.n7923 3.1505
R9927 VDD.n7923 VDD.n7922 3.1505
R9928 VDD.n7927 VDD.n7926 3.1505
R9929 VDD.n7926 VDD.n7925 3.1505
R9930 VDD.n7931 VDD.n7930 3.1505
R9931 VDD.n7930 VDD.n7929 3.1505
R9932 VDD.n7934 VDD.n7933 3.1505
R9933 VDD.n7933 VDD.n7932 3.1505
R9934 VDD.n7937 VDD.n7936 3.1505
R9935 VDD.n7936 VDD.n7935 3.1505
R9936 VDD.n7940 VDD.n7939 3.1505
R9937 VDD.n7939 VDD.n7938 3.1505
R9938 VDD.n7944 VDD.n7943 3.1505
R9939 VDD.n7943 VDD.n7942 3.1505
R9940 VDD.n7947 VDD.n7946 3.1505
R9941 VDD.n7946 VDD.n7945 3.1505
R9942 VDD.n7950 VDD.n7949 3.1505
R9943 VDD.n7949 VDD.n7948 3.1505
R9944 VDD.n7953 VDD.n7952 3.1505
R9945 VDD.n7952 VDD.n7951 3.1505
R9946 VDD.n7957 VDD.n7956 3.1505
R9947 VDD.n7956 VDD.n7955 3.1505
R9948 VDD.n8142 VDD.n8141 3.1505
R9949 VDD.n8141 VDD.n8140 3.1505
R9950 VDD.n8138 VDD.n8137 3.1505
R9951 VDD.n8137 VDD.n8136 3.1505
R9952 VDD.n8134 VDD.n8133 3.1505
R9953 VDD.n8133 VDD.n8132 3.1505
R9954 VDD.n8131 VDD.n8130 3.1505
R9955 VDD.n8130 VDD.n8129 3.1505
R9956 VDD.n8127 VDD.n8126 3.1505
R9957 VDD.n8126 VDD.n8125 3.1505
R9958 VDD.n8124 VDD.n8123 3.1505
R9959 VDD.n8123 VDD.n8122 3.1505
R9960 VDD.n8121 VDD.n8120 3.1505
R9961 VDD.n8120 VDD.n8119 3.1505
R9962 VDD.n7083 VDD.n7056 3.1505
R9963 VDD.n6985 VDD.n6984 3.1505
R9964 VDD.n6984 VDD.n6983 3.1505
R9965 VDD.n6989 VDD.n6988 3.1505
R9966 VDD.n6988 VDD.n6987 3.1505
R9967 VDD.n6992 VDD.n6991 3.1505
R9968 VDD.n6991 VDD.n6990 3.1505
R9969 VDD.n6996 VDD.n6995 3.1505
R9970 VDD.n6995 VDD.n6994 3.1505
R9971 VDD.n6999 VDD.n6998 3.1505
R9972 VDD.n6998 VDD.n6997 3.1505
R9973 VDD.n7002 VDD.n7001 3.1505
R9974 VDD.n7001 VDD.n7000 3.1505
R9975 VDD.n7006 VDD.n7005 3.1505
R9976 VDD.n7005 VDD.n7004 3.1505
R9977 VDD.n7009 VDD.n7008 3.1505
R9978 VDD.n7008 VDD.n7007 3.1505
R9979 VDD.n7012 VDD.n7011 3.1505
R9980 VDD.n7011 VDD.n7010 3.1505
R9981 VDD.n7015 VDD.n7014 3.1505
R9982 VDD.n7014 VDD.n7013 3.1505
R9983 VDD.n7018 VDD.n7017 3.1505
R9984 VDD.n7017 VDD.n7016 3.1505
R9985 VDD.n7022 VDD.n7021 3.1505
R9986 VDD.n7021 VDD.n7020 3.1505
R9987 VDD.n7025 VDD.n7024 3.1505
R9988 VDD.n7024 VDD.n7023 3.1505
R9989 VDD.n7028 VDD.n7027 3.1505
R9990 VDD.n7027 VDD.n7026 3.1505
R9991 VDD.n7031 VDD.n7030 3.1505
R9992 VDD.n7030 VDD.n7029 3.1505
R9993 VDD.n7034 VDD.n7033 3.1505
R9994 VDD.n7033 VDD.n7032 3.1505
R9995 VDD.n7037 VDD.n7036 3.1505
R9996 VDD.n7036 VDD.n7035 3.1505
R9997 VDD.n7041 VDD.n7040 3.1505
R9998 VDD.n7040 VDD.n7039 3.1505
R9999 VDD.n7044 VDD.n7043 3.1505
R10000 VDD.n7043 VDD.n7042 3.1505
R10001 VDD.n7048 VDD.n7047 3.1505
R10002 VDD.n7047 VDD.n7046 3.1505
R10003 VDD.n7051 VDD.n7050 3.1505
R10004 VDD.n7050 VDD.n7049 3.1505
R10005 VDD.n7055 VDD.n7054 3.1505
R10006 VDD.n7054 VDD.n7053 3.1505
R10007 VDD.n7082 VDD.n7081 3.1505
R10008 VDD.n7080 VDD.n7079 3.1505
R10009 VDD.n7078 VDD.n7077 3.1505
R10010 VDD.n7075 VDD.n7074 3.1505
R10011 VDD.n7073 VDD.n7072 3.1505
R10012 VDD.n7071 VDD.n7070 3.1505
R10013 VDD.n7068 VDD.n7067 3.1505
R10014 VDD.n7066 VDD.n7065 3.1505
R10015 VDD.n7064 VDD.n7063 3.1505
R10016 VDD.n7062 VDD.n7061 3.1505
R10017 VDD.n8168 VDD.n8167 3.1505
R10018 VDD.n8170 VDD.n8169 3.1505
R10019 VDD.n8172 VDD.n8171 3.1505
R10020 VDD.n8174 VDD.n8173 3.1505
R10021 VDD.n8176 VDD.n8175 3.1505
R10022 VDD.n8179 VDD.n8178 3.1505
R10023 VDD.n8181 VDD.n8180 3.1505
R10024 VDD.n8183 VDD.n8182 3.1505
R10025 VDD.n8186 VDD.n8185 3.1505
R10026 VDD.n8188 VDD.n8187 3.1505
R10027 VDD.n8191 VDD.n8190 3.1505
R10028 VDD.n8193 VDD.n8192 3.1505
R10029 VDD.n8195 VDD.n8194 3.1505
R10030 VDD.n8197 VDD.n8196 3.1505
R10031 VDD.n8200 VDD.n8199 3.1505
R10032 VDD.n8202 VDD.n8201 3.1505
R10033 VDD.n8205 VDD.n8204 3.1505
R10034 VDD.n8207 VDD.n8206 3.1505
R10035 VDD.n8209 VDD.n8208 3.1505
R10036 VDD.n8211 VDD.n8210 3.1505
R10037 VDD.n8213 VDD.n8212 3.1505
R10038 VDD.n6981 VDD.n6980 3.1505
R10039 VDD.n1027 VDD.n1026 3.1505
R10040 VDD.n6853 VDD.n6852 3.1505
R10041 VDD.n6646 VDD.n6645 3.1505
R10042 VDD.n6645 VDD.n6644 3.1505
R10043 VDD.n6642 VDD.n6641 3.1505
R10044 VDD.n6641 VDD.n6640 3.1505
R10045 VDD.n6639 VDD.n6638 3.1505
R10046 VDD.n6638 VDD.n6637 3.1505
R10047 VDD.n6635 VDD.n6634 3.1505
R10048 VDD.n6634 VDD.n6633 3.1505
R10049 VDD.n869 VDD.n868 3.1505
R10050 VDD.n868 VDD.n867 3.1505
R10051 VDD.n866 VDD.n865 3.1505
R10052 VDD.n865 VDD.n864 3.1505
R10053 VDD.n863 VDD.n862 3.1505
R10054 VDD.n862 VDD.n861 3.1505
R10055 VDD.n860 VDD.n859 3.1505
R10056 VDD.n859 VDD.n858 3.1505
R10057 VDD.n857 VDD.n856 3.1505
R10058 VDD.n856 VDD.n855 3.1505
R10059 VDD.n854 VDD.n853 3.1505
R10060 VDD.n853 VDD.n852 3.1505
R10061 VDD.n851 VDD.n850 3.1505
R10062 VDD.n850 VDD.n849 3.1505
R10063 VDD.n848 VDD.n847 3.1505
R10064 VDD.n847 VDD.n846 3.1505
R10065 VDD.n845 VDD.n844 3.1505
R10066 VDD.n844 VDD.n843 3.1505
R10067 VDD.n842 VDD.n841 3.1505
R10068 VDD.n841 VDD.n840 3.1505
R10069 VDD.n839 VDD.n838 3.1505
R10070 VDD.n838 VDD.n837 3.1505
R10071 VDD.n836 VDD.n835 3.1505
R10072 VDD.n835 VDD.n834 3.1505
R10073 VDD.n833 VDD.n832 3.1505
R10074 VDD.n832 VDD.n831 3.1505
R10075 VDD.n830 VDD.n829 3.1505
R10076 VDD.n829 VDD.n828 3.1505
R10077 VDD.n827 VDD.n826 3.1505
R10078 VDD.n826 VDD.n825 3.1505
R10079 VDD.n824 VDD.n823 3.1505
R10080 VDD.n823 VDD.n822 3.1505
R10081 VDD.n821 VDD.n820 3.1505
R10082 VDD.n820 VDD.n819 3.1505
R10083 VDD.n818 VDD.n817 3.1505
R10084 VDD.n817 VDD.n816 3.1505
R10085 VDD.n815 VDD.n814 3.1505
R10086 VDD.n814 VDD.n813 3.1505
R10087 VDD.n812 VDD.n811 3.1505
R10088 VDD.n811 VDD.n810 3.1505
R10089 VDD.n809 VDD.n808 3.1505
R10090 VDD.n808 VDD.n807 3.1505
R10091 VDD.n805 VDD.n804 3.1505
R10092 VDD.n804 VDD.n803 3.1505
R10093 VDD.n802 VDD.n801 3.1505
R10094 VDD.n801 VDD.n800 3.1505
R10095 VDD.n798 VDD.n797 3.1505
R10096 VDD.n797 VDD.n796 3.1505
R10097 VDD.n795 VDD.n794 3.1505
R10098 VDD.n793 VDD.n792 3.1505
R10099 VDD.n792 VDD.n791 3.1505
R10100 VDD.n790 VDD.n789 3.1505
R10101 VDD.n789 VDD.n788 3.1505
R10102 VDD.n787 VDD.n786 3.1505
R10103 VDD.n786 VDD.n785 3.1505
R10104 VDD.n784 VDD.n783 3.1505
R10105 VDD.n783 VDD.n782 3.1505
R10106 VDD.n781 VDD.n780 3.1505
R10107 VDD.n780 VDD.n779 3.1505
R10108 VDD.n778 VDD.n777 3.1505
R10109 VDD.n777 VDD.n776 3.1505
R10110 VDD.n775 VDD.n774 3.1505
R10111 VDD.n774 VDD.n773 3.1505
R10112 VDD.n771 VDD.n770 3.1505
R10113 VDD.n770 VDD.n769 3.1505
R10114 VDD.n768 VDD.n767 3.1505
R10115 VDD.n767 VDD.n766 3.1505
R10116 VDD.n765 VDD.n764 3.1505
R10117 VDD.n764 VDD.n763 3.1505
R10118 VDD.n761 VDD.n760 3.1505
R10119 VDD.n760 VDD.n759 3.1505
R10120 VDD.n758 VDD.n757 3.1505
R10121 VDD.n757 VDD.n756 3.1505
R10122 VDD.n1058 VDD.n1057 3.1505
R10123 VDD.n1057 VDD.n1056 3.1505
R10124 VDD.n1061 VDD.n1060 3.1505
R10125 VDD.n1060 VDD.n1059 3.1505
R10126 VDD.n1065 VDD.n1064 3.1505
R10127 VDD.n1064 VDD.n1063 3.1505
R10128 VDD.n1068 VDD.n1067 3.1505
R10129 VDD.n1067 VDD.n1066 3.1505
R10130 VDD.n1071 VDD.n1070 3.1505
R10131 VDD.n1070 VDD.n1069 3.1505
R10132 VDD.n1075 VDD.n1074 3.1505
R10133 VDD.n1074 VDD.n1073 3.1505
R10134 VDD.n1078 VDD.n1077 3.1505
R10135 VDD.n1077 VDD.n1076 3.1505
R10136 VDD.n1081 VDD.n1080 3.1505
R10137 VDD.n1080 VDD.n1079 3.1505
R10138 VDD.n1085 VDD.n1084 3.1505
R10139 VDD.n1084 VDD.n1083 3.1505
R10140 VDD.n1088 VDD.n1087 3.1505
R10141 VDD.n1087 VDD.n1086 3.1505
R10142 VDD.n1092 VDD.n1091 3.1505
R10143 VDD.n1091 VDD.n1090 3.1505
R10144 VDD.n1095 VDD.n1094 3.1505
R10145 VDD.n1094 VDD.n1093 3.1505
R10146 VDD.n1789 VDD.n1788 3.1505
R10147 VDD.n1927 VDD.n1926 3.1505
R10148 VDD.n2031 VDD.n2030 3.1505
R10149 VDD.n1664 VDD.n1663 3.1505
R10150 VDD.n1666 VDD.n1665 3.1505
R10151 VDD.n1668 VDD.n1667 3.1505
R10152 VDD.n1670 VDD.n1669 3.1505
R10153 VDD.n1673 VDD.n1672 3.1505
R10154 VDD.n1676 VDD.n1675 3.1505
R10155 VDD.n1679 VDD.n1678 3.1505
R10156 VDD.n1682 VDD.n1681 3.1505
R10157 VDD.n1685 VDD.n1684 3.1505
R10158 VDD.n1688 VDD.n1687 3.1505
R10159 VDD.n1691 VDD.n1690 3.1505
R10160 VDD.n1694 VDD.n1693 3.1505
R10161 VDD.n1697 VDD.n1696 3.1505
R10162 VDD.n1700 VDD.n1699 3.1505
R10163 VDD.n1703 VDD.n1702 3.1505
R10164 VDD.n1706 VDD.n1705 3.1505
R10165 VDD.n1709 VDD.n1708 3.1505
R10166 VDD.n1712 VDD.n1711 3.1505
R10167 VDD.n1715 VDD.n1714 3.1505
R10168 VDD.n1718 VDD.n1717 3.1505
R10169 VDD.n1721 VDD.n1720 3.1505
R10170 VDD.n1724 VDD.n1723 3.1505
R10171 VDD.n1727 VDD.n1726 3.1505
R10172 VDD.n1730 VDD.n1729 3.1505
R10173 VDD.n1733 VDD.n1732 3.1505
R10174 VDD.n1736 VDD.n1735 3.1505
R10175 VDD.n1739 VDD.n1738 3.1505
R10176 VDD.n1742 VDD.n1741 3.1505
R10177 VDD.n1745 VDD.n1744 3.1505
R10178 VDD.n1748 VDD.n1747 3.1505
R10179 VDD.n1751 VDD.n1750 3.1505
R10180 VDD.n1754 VDD.n1753 3.1505
R10181 VDD.n1757 VDD.n1756 3.1505
R10182 VDD.n1760 VDD.n1759 3.1505
R10183 VDD.n1763 VDD.n1762 3.1505
R10184 VDD.n1766 VDD.n1765 3.1505
R10185 VDD.n1769 VDD.n1768 3.1505
R10186 VDD.n1772 VDD.n1771 3.1505
R10187 VDD.n1775 VDD.n1774 3.1505
R10188 VDD.n1778 VDD.n1777 3.1505
R10189 VDD.n1781 VDD.n1780 3.1505
R10190 VDD.n1784 VDD.n1783 3.1505
R10191 VDD.n1787 VDD.n1786 3.1505
R10192 VDD.n1661 VDD.n1660 3.1505
R10193 VDD.n1659 VDD.n1658 3.1505
R10194 VDD.n1802 VDD.n1801 3.1505
R10195 VDD.n1804 VDD.n1803 3.1505
R10196 VDD.n1806 VDD.n1805 3.1505
R10197 VDD.n1808 VDD.n1807 3.1505
R10198 VDD.n1811 VDD.n1810 3.1505
R10199 VDD.n1814 VDD.n1813 3.1505
R10200 VDD.n1817 VDD.n1816 3.1505
R10201 VDD.n1820 VDD.n1819 3.1505
R10202 VDD.n1823 VDD.n1822 3.1505
R10203 VDD.n1826 VDD.n1825 3.1505
R10204 VDD.n1829 VDD.n1828 3.1505
R10205 VDD.n1832 VDD.n1831 3.1505
R10206 VDD.n1835 VDD.n1834 3.1505
R10207 VDD.n1838 VDD.n1837 3.1505
R10208 VDD.n1841 VDD.n1840 3.1505
R10209 VDD.n1844 VDD.n1843 3.1505
R10210 VDD.n1847 VDD.n1846 3.1505
R10211 VDD.n1850 VDD.n1849 3.1505
R10212 VDD.n1853 VDD.n1852 3.1505
R10213 VDD.n1856 VDD.n1855 3.1505
R10214 VDD.n1859 VDD.n1858 3.1505
R10215 VDD.n1862 VDD.n1861 3.1505
R10216 VDD.n1865 VDD.n1864 3.1505
R10217 VDD.n1868 VDD.n1867 3.1505
R10218 VDD.n1871 VDD.n1870 3.1505
R10219 VDD.n1874 VDD.n1873 3.1505
R10220 VDD.n1877 VDD.n1876 3.1505
R10221 VDD.n1880 VDD.n1879 3.1505
R10222 VDD.n1883 VDD.n1882 3.1505
R10223 VDD.n1886 VDD.n1885 3.1505
R10224 VDD.n1889 VDD.n1888 3.1505
R10225 VDD.n1892 VDD.n1891 3.1505
R10226 VDD.n1895 VDD.n1894 3.1505
R10227 VDD.n1898 VDD.n1897 3.1505
R10228 VDD.n1901 VDD.n1900 3.1505
R10229 VDD.n1904 VDD.n1903 3.1505
R10230 VDD.n1907 VDD.n1906 3.1505
R10231 VDD.n1910 VDD.n1909 3.1505
R10232 VDD.n1913 VDD.n1912 3.1505
R10233 VDD.n1916 VDD.n1915 3.1505
R10234 VDD.n1919 VDD.n1918 3.1505
R10235 VDD.n1922 VDD.n1921 3.1505
R10236 VDD.n1925 VDD.n1924 3.1505
R10237 VDD.n1799 VDD.n1798 3.1505
R10238 VDD.n1797 VDD.n1796 3.1505
R10239 VDD.n2029 VDD.n2028 3.1505
R10240 VDD.n2026 VDD.n2025 3.1505
R10241 VDD.n2024 VDD.n2023 3.1505
R10242 VDD.n2021 VDD.n2020 3.1505
R10243 VDD.n2019 VDD.n2018 3.1505
R10244 VDD.n2016 VDD.n2015 3.1505
R10245 VDD.n2014 VDD.n2013 3.1505
R10246 VDD.n2011 VDD.n2010 3.1505
R10247 VDD.n2009 VDD.n2008 3.1505
R10248 VDD.n2006 VDD.n2005 3.1505
R10249 VDD.n2004 VDD.n2003 3.1505
R10250 VDD.n2001 VDD.n2000 3.1505
R10251 VDD.n1999 VDD.n1998 3.1505
R10252 VDD.n1996 VDD.n1995 3.1505
R10253 VDD.n1994 VDD.n1993 3.1505
R10254 VDD.n1991 VDD.n1990 3.1505
R10255 VDD.n1989 VDD.n1988 3.1505
R10256 VDD.n1986 VDD.n1985 3.1505
R10257 VDD.n1984 VDD.n1983 3.1505
R10258 VDD.n1981 VDD.n1980 3.1505
R10259 VDD.n1979 VDD.n1978 3.1505
R10260 VDD.n1977 VDD.n1976 3.1505
R10261 VDD.n1975 VDD.n1974 3.1505
R10262 VDD.n1973 VDD.n1972 3.1505
R10263 VDD.n1971 VDD.n1970 3.1505
R10264 VDD.n1969 VDD.n1968 3.1505
R10265 VDD.n1967 VDD.n1966 3.1505
R10266 VDD.n1965 VDD.n1964 3.1505
R10267 VDD.n1963 VDD.n1962 3.1505
R10268 VDD.n1961 VDD.n1960 3.1505
R10269 VDD.n1959 VDD.n1958 3.1505
R10270 VDD.n1957 VDD.n1956 3.1505
R10271 VDD.n1955 VDD.n1954 3.1505
R10272 VDD.n1953 VDD.n1952 3.1505
R10273 VDD.n1951 VDD.n1950 3.1505
R10274 VDD.n1949 VDD.n1948 3.1505
R10275 VDD.n1947 VDD.n1946 3.1505
R10276 VDD.n1945 VDD.n1944 3.1505
R10277 VDD.n1943 VDD.n1942 3.1505
R10278 VDD.n1941 VDD.n1940 3.1505
R10279 VDD.n1939 VDD.n1938 3.1505
R10280 VDD.n1937 VDD.n1936 3.1505
R10281 VDD.n1935 VDD.n1934 3.1505
R10282 VDD.n1933 VDD.n1932 3.1505
R10283 VDD.n1931 VDD.n1930 3.1505
R10284 VDD.n1343 VDD.n1097 3.1505
R10285 VDD.n1244 VDD.n1243 3.1505
R10286 VDD.n1339 VDD.n1338 3.1505
R10287 VDD.n1337 VDD.n1336 3.1505
R10288 VDD.n1334 VDD.n1333 3.1505
R10289 VDD.n1332 VDD.n1331 3.1505
R10290 VDD.n1329 VDD.n1328 3.1505
R10291 VDD.n1327 VDD.n1326 3.1505
R10292 VDD.n1324 VDD.n1323 3.1505
R10293 VDD.n1322 VDD.n1321 3.1505
R10294 VDD.n1319 VDD.n1318 3.1505
R10295 VDD.n1317 VDD.n1316 3.1505
R10296 VDD.n1314 VDD.n1313 3.1505
R10297 VDD.n1312 VDD.n1311 3.1505
R10298 VDD.n1309 VDD.n1308 3.1505
R10299 VDD.n1307 VDD.n1306 3.1505
R10300 VDD.n1304 VDD.n1303 3.1505
R10301 VDD.n1302 VDD.n1301 3.1505
R10302 VDD.n1299 VDD.n1298 3.1505
R10303 VDD.n1297 VDD.n1296 3.1505
R10304 VDD.n1294 VDD.n1293 3.1505
R10305 VDD.n1292 VDD.n1291 3.1505
R10306 VDD.n1290 VDD.n1289 3.1505
R10307 VDD.n1288 VDD.n1287 3.1505
R10308 VDD.n1286 VDD.n1285 3.1505
R10309 VDD.n1284 VDD.n1283 3.1505
R10310 VDD.n1282 VDD.n1281 3.1505
R10311 VDD.n1280 VDD.n1279 3.1505
R10312 VDD.n1278 VDD.n1277 3.1505
R10313 VDD.n1276 VDD.n1275 3.1505
R10314 VDD.n1274 VDD.n1273 3.1505
R10315 VDD.n1272 VDD.n1271 3.1505
R10316 VDD.n1270 VDD.n1269 3.1505
R10317 VDD.n1268 VDD.n1267 3.1505
R10318 VDD.n1266 VDD.n1265 3.1505
R10319 VDD.n1264 VDD.n1263 3.1505
R10320 VDD.n1262 VDD.n1261 3.1505
R10321 VDD.n1260 VDD.n1259 3.1505
R10322 VDD.n1258 VDD.n1257 3.1505
R10323 VDD.n1256 VDD.n1255 3.1505
R10324 VDD.n1254 VDD.n1253 3.1505
R10325 VDD.n1252 VDD.n1251 3.1505
R10326 VDD.n1250 VDD.n1249 3.1505
R10327 VDD.n1248 VDD.n1247 3.1505
R10328 VDD.n1246 VDD.n1245 3.1505
R10329 VDD.n1342 VDD.n1341 3.1505
R10330 VDD.n1462 VDD.n1461 3.1505
R10331 VDD.n1464 VDD.n1463 3.1505
R10332 VDD.n1466 VDD.n1465 3.1505
R10333 VDD.n1468 VDD.n1467 3.1505
R10334 VDD.n1470 VDD.n1469 3.1505
R10335 VDD.n1472 VDD.n1471 3.1505
R10336 VDD.n1475 VDD.n1474 3.1505
R10337 VDD.n1477 VDD.n1476 3.1505
R10338 VDD.n1479 VDD.n1478 3.1505
R10339 VDD.n1481 VDD.n1480 3.1505
R10340 VDD.n1483 VDD.n1482 3.1505
R10341 VDD.n1485 VDD.n1484 3.1505
R10342 VDD.n1487 VDD.n1486 3.1505
R10343 VDD.n1489 VDD.n1488 3.1505
R10344 VDD.n1491 VDD.n1490 3.1505
R10345 VDD.n1493 VDD.n1492 3.1505
R10346 VDD.n1495 VDD.n1494 3.1505
R10347 VDD.n1497 VDD.n1496 3.1505
R10348 VDD.n1499 VDD.n1498 3.1505
R10349 VDD.n1501 VDD.n1500 3.1505
R10350 VDD.n1503 VDD.n1502 3.1505
R10351 VDD.n1505 VDD.n1504 3.1505
R10352 VDD.n1507 VDD.n1506 3.1505
R10353 VDD.n1509 VDD.n1508 3.1505
R10354 VDD.n1511 VDD.n1510 3.1505
R10355 VDD.n1514 VDD.n1513 3.1505
R10356 VDD.n1516 VDD.n1515 3.1505
R10357 VDD.n1518 VDD.n1517 3.1505
R10358 VDD.n1520 VDD.n1519 3.1505
R10359 VDD.n1522 VDD.n1521 3.1505
R10360 VDD.n1524 VDD.n1523 3.1505
R10361 VDD.n1531 VDD.n1530 3.1505
R10362 VDD.n1533 VDD.n1532 3.1505
R10363 VDD.n1535 VDD.n1534 3.1505
R10364 VDD.n1537 VDD.n1536 3.1505
R10365 VDD.n1539 VDD.n1538 3.1505
R10366 VDD.n1541 VDD.n1540 3.1505
R10367 VDD.n1543 VDD.n1542 3.1505
R10368 VDD.n1547 VDD.n1546 3.1505
R10369 VDD.n1549 VDD.n1548 3.1505
R10370 VDD.n1551 VDD.n1550 3.1505
R10371 VDD.n1553 VDD.n1552 3.1505
R10372 VDD.n1555 VDD.n1554 3.1505
R10373 VDD.n1557 VDD.n1556 3.1505
R10374 VDD.n1559 VDD.n1558 3.1505
R10375 VDD.n1561 VDD.n1560 3.1505
R10376 VDD.n1563 VDD.n1562 3.1505
R10377 VDD.n1565 VDD.n1564 3.1505
R10378 VDD.n1567 VDD.n1566 3.1505
R10379 VDD.n1569 VDD.n1568 3.1505
R10380 VDD.n1571 VDD.n1570 3.1505
R10381 VDD.n1573 VDD.n1572 3.1505
R10382 VDD.n1575 VDD.n1574 3.1505
R10383 VDD.n1577 VDD.n1576 3.1505
R10384 VDD.n1579 VDD.n1578 3.1505
R10385 VDD.n1581 VDD.n1580 3.1505
R10386 VDD.n1583 VDD.n1582 3.1505
R10387 VDD.n1585 VDD.n1584 3.1505
R10388 VDD.n1587 VDD.n1586 3.1505
R10389 VDD.n1589 VDD.n1588 3.1505
R10390 VDD.n1591 VDD.n1590 3.1505
R10391 VDD.n1593 VDD.n1592 3.1505
R10392 VDD.n1595 VDD.n1594 3.1505
R10393 VDD.n1597 VDD.n1596 3.1505
R10394 VDD.n1599 VDD.n1598 3.1505
R10395 VDD.n1601 VDD.n1600 3.1505
R10396 VDD.n1603 VDD.n1602 3.1505
R10397 VDD.n1605 VDD.n1604 3.1505
R10398 VDD.n1607 VDD.n1606 3.1505
R10399 VDD.n1609 VDD.n1608 3.1505
R10400 VDD.n1611 VDD.n1610 3.1505
R10401 VDD.n1613 VDD.n1612 3.1505
R10402 VDD.n1615 VDD.n1614 3.1505
R10403 VDD.n1617 VDD.n1616 3.1505
R10404 VDD.n1619 VDD.n1618 3.1505
R10405 VDD.n1621 VDD.n1620 3.1505
R10406 VDD.n1623 VDD.n1622 3.1505
R10407 VDD.n1625 VDD.n1624 3.1505
R10408 VDD.n1627 VDD.n1626 3.1505
R10409 VDD.n1629 VDD.n1628 3.1505
R10410 VDD.n1631 VDD.n1630 3.1505
R10411 VDD.n1633 VDD.n1632 3.1505
R10412 VDD.n1635 VDD.n1634 3.1505
R10413 VDD.n1637 VDD.n1636 3.1505
R10414 VDD.n1640 VDD.n1639 3.1505
R10415 VDD.n1642 VDD.n1641 3.1505
R10416 VDD.n1644 VDD.n1643 3.1505
R10417 VDD.n1646 VDD.n1645 3.1505
R10418 VDD.n1648 VDD.n1647 3.1505
R10419 VDD.n1650 VDD.n1649 3.1505
R10420 VDD.n1652 VDD.n1651 3.1505
R10421 VDD.n1133 VDD.n1132 3.1505
R10422 VDD.n1135 VDD.n1134 3.1505
R10423 VDD.n1137 VDD.n1136 3.1505
R10424 VDD.n1139 VDD.n1138 3.1505
R10425 VDD.n1141 VDD.n1140 3.1505
R10426 VDD.n1143 VDD.n1142 3.1505
R10427 VDD.n1146 VDD.n1145 3.1505
R10428 VDD.n1149 VDD.n1148 3.1505
R10429 VDD.n1151 VDD.n1150 3.1505
R10430 VDD.n1154 VDD.n1153 3.1505
R10431 VDD.n1156 VDD.n1155 3.1505
R10432 VDD.n1158 VDD.n1157 3.1505
R10433 VDD.n1160 VDD.n1159 3.1505
R10434 VDD.n1162 VDD.n1161 3.1505
R10435 VDD.n1164 VDD.n1163 3.1505
R10436 VDD.n1167 VDD.n1166 3.1505
R10437 VDD.n1169 VDD.n1168 3.1505
R10438 VDD.n1171 VDD.n1170 3.1505
R10439 VDD.n1173 VDD.n1172 3.1505
R10440 VDD.n1176 VDD.n1175 3.1505
R10441 VDD.n1178 VDD.n1177 3.1505
R10442 VDD.n1180 VDD.n1179 3.1505
R10443 VDD.n1182 VDD.n1181 3.1505
R10444 VDD.n1184 VDD.n1183 3.1505
R10445 VDD.n1186 VDD.n1185 3.1505
R10446 VDD.n1188 VDD.n1187 3.1505
R10447 VDD.n1190 VDD.n1189 3.1505
R10448 VDD.n1192 VDD.n1191 3.1505
R10449 VDD.n1194 VDD.n1193 3.1505
R10450 VDD.n1196 VDD.n1195 3.1505
R10451 VDD.n1198 VDD.n1197 3.1505
R10452 VDD.n1200 VDD.n1199 3.1505
R10453 VDD.n1202 VDD.n1201 3.1505
R10454 VDD.n1204 VDD.n1203 3.1505
R10455 VDD.n1206 VDD.n1205 3.1505
R10456 VDD.n1208 VDD.n1207 3.1505
R10457 VDD.n1210 VDD.n1209 3.1505
R10458 VDD.n1212 VDD.n1211 3.1505
R10459 VDD.n1214 VDD.n1213 3.1505
R10460 VDD.n1216 VDD.n1215 3.1505
R10461 VDD.n1218 VDD.n1217 3.1505
R10462 VDD.n1220 VDD.n1219 3.1505
R10463 VDD.n1222 VDD.n1221 3.1505
R10464 VDD.n1225 VDD.n1224 3.1505
R10465 VDD.n1228 VDD.n1227 3.1505
R10466 VDD.n1230 VDD.n1229 3.1505
R10467 VDD.n1232 VDD.n1231 3.1505
R10468 VDD.n1234 VDD.n1233 3.1505
R10469 VDD.n1236 VDD.n1235 3.1505
R10470 VDD.n1238 VDD.n1237 3.1505
R10471 VDD.n2051 VDD.n2050 3.1505
R10472 VDD.n2050 VDD.n2049 3.1505
R10473 VDD.n2054 VDD.n2053 3.1505
R10474 VDD.n2053 VDD.n2052 3.1505
R10475 VDD.n2057 VDD.n2056 3.1505
R10476 VDD.n2056 VDD.n2055 3.1505
R10477 VDD.n2060 VDD.n2059 3.1505
R10478 VDD.n2059 VDD.n2058 3.1505
R10479 VDD.n2063 VDD.n2062 3.1505
R10480 VDD.n2062 VDD.n2061 3.1505
R10481 VDD.n2066 VDD.n2065 3.1505
R10482 VDD.n2065 VDD.n2064 3.1505
R10483 VDD.n2070 VDD.n2069 3.1505
R10484 VDD.n2069 VDD.n2068 3.1505
R10485 VDD.n2073 VDD.n2072 3.1505
R10486 VDD.n2072 VDD.n2071 3.1505
R10487 VDD.n2076 VDD.n2075 3.1505
R10488 VDD.n2075 VDD.n2074 3.1505
R10489 VDD.n2079 VDD.n2078 3.1505
R10490 VDD.n2078 VDD.n2077 3.1505
R10491 VDD.n2082 VDD.n2081 3.1505
R10492 VDD.n2081 VDD.n2080 3.1505
R10493 VDD.n2085 VDD.n2084 3.1505
R10494 VDD.n2084 VDD.n2083 3.1505
R10495 VDD.n2088 VDD.n2087 3.1505
R10496 VDD.n2087 VDD.n2086 3.1505
R10497 VDD.n2091 VDD.n2090 3.1505
R10498 VDD.n2090 VDD.n2089 3.1505
R10499 VDD.n2094 VDD.n2093 3.1505
R10500 VDD.n2093 VDD.n2092 3.1505
R10501 VDD.n2097 VDD.n2096 3.1505
R10502 VDD.n2096 VDD.n2095 3.1505
R10503 VDD.n2100 VDD.n2099 3.1505
R10504 VDD.n2099 VDD.n2098 3.1505
R10505 VDD.n2103 VDD.n2102 3.1505
R10506 VDD.n2102 VDD.n2101 3.1505
R10507 VDD.n2106 VDD.n2105 3.1505
R10508 VDD.n2105 VDD.n2104 3.1505
R10509 VDD.n2109 VDD.n2108 3.1505
R10510 VDD.n2108 VDD.n2107 3.1505
R10511 VDD.n2112 VDD.n2111 3.1505
R10512 VDD.n2111 VDD.n2110 3.1505
R10513 VDD.n2115 VDD.n2114 3.1505
R10514 VDD.n2114 VDD.n2113 3.1505
R10515 VDD.n2118 VDD.n2117 3.1505
R10516 VDD.n2117 VDD.n2116 3.1505
R10517 VDD.n2121 VDD.n2120 3.1505
R10518 VDD.n2120 VDD.n2119 3.1505
R10519 VDD.n2124 VDD.n2123 3.1505
R10520 VDD.n2123 VDD.n2122 3.1505
R10521 VDD.n2128 VDD.n2127 3.1505
R10522 VDD.n2127 VDD.n2126 3.1505
R10523 VDD.n2131 VDD.n2130 3.1505
R10524 VDD.n2130 VDD.n2129 3.1505
R10525 VDD.n2134 VDD.n2133 3.1505
R10526 VDD.n2133 VDD.n2132 3.1505
R10527 VDD.n2137 VDD.n2136 3.1505
R10528 VDD.n2136 VDD.n2135 3.1505
R10529 VDD.n2140 VDD.n2139 3.1505
R10530 VDD.n2139 VDD.n2138 3.1505
R10531 VDD.n2143 VDD.n2142 3.1505
R10532 VDD.n2142 VDD.n2141 3.1505
R10533 VDD.n2155 VDD.n2154 3.1505
R10534 VDD.n2154 VDD.n2153 3.1505
R10535 VDD.n2158 VDD.n2157 3.1505
R10536 VDD.n2157 VDD.n2156 3.1505
R10537 VDD.n2161 VDD.n2160 3.1505
R10538 VDD.n2160 VDD.n2159 3.1505
R10539 VDD.n2164 VDD.n2163 3.1505
R10540 VDD.n2163 VDD.n2162 3.1505
R10541 VDD.n2167 VDD.n2166 3.1505
R10542 VDD.n2166 VDD.n2165 3.1505
R10543 VDD.n2170 VDD.n2169 3.1505
R10544 VDD.n2169 VDD.n2168 3.1505
R10545 VDD.n2173 VDD.n2172 3.1505
R10546 VDD.n2172 VDD.n2171 3.1505
R10547 VDD.n2177 VDD.n2176 3.1505
R10548 VDD.n2176 VDD.n2175 3.1505
R10549 VDD.n2180 VDD.n2179 3.1505
R10550 VDD.n2179 VDD.n2178 3.1505
R10551 VDD.n2183 VDD.n2182 3.1505
R10552 VDD.n2182 VDD.n2181 3.1505
R10553 VDD.n2186 VDD.n2185 3.1505
R10554 VDD.n2185 VDD.n2184 3.1505
R10555 VDD.n2189 VDD.n2188 3.1505
R10556 VDD.n2188 VDD.n2187 3.1505
R10557 VDD.n2192 VDD.n2191 3.1505
R10558 VDD.n2191 VDD.n2190 3.1505
R10559 VDD.n2195 VDD.n2194 3.1505
R10560 VDD.n2194 VDD.n2193 3.1505
R10561 VDD.n2198 VDD.n2197 3.1505
R10562 VDD.n2197 VDD.n2196 3.1505
R10563 VDD.n2201 VDD.n2200 3.1505
R10564 VDD.n2200 VDD.n2199 3.1505
R10565 VDD.n2204 VDD.n2203 3.1505
R10566 VDD.n2203 VDD.n2202 3.1505
R10567 VDD.n2207 VDD.n2206 3.1505
R10568 VDD.n2206 VDD.n2205 3.1505
R10569 VDD.n2210 VDD.n2209 3.1505
R10570 VDD.n2209 VDD.n2208 3.1505
R10571 VDD.n2213 VDD.n2212 3.1505
R10572 VDD.n2212 VDD.n2211 3.1505
R10573 VDD.n2216 VDD.n2215 3.1505
R10574 VDD.n2215 VDD.n2214 3.1505
R10575 VDD.n2219 VDD.n2218 3.1505
R10576 VDD.n2218 VDD.n2217 3.1505
R10577 VDD.n2222 VDD.n2221 3.1505
R10578 VDD.n2221 VDD.n2220 3.1505
R10579 VDD.n2225 VDD.n2224 3.1505
R10580 VDD.n2224 VDD.n2223 3.1505
R10581 VDD.n2228 VDD.n2227 3.1505
R10582 VDD.n2227 VDD.n2226 3.1505
R10583 VDD.n2231 VDD.n2230 3.1505
R10584 VDD.n2230 VDD.n2229 3.1505
R10585 VDD.n2234 VDD.n2233 3.1505
R10586 VDD.n2233 VDD.n2232 3.1505
R10587 VDD.n2237 VDD.n2236 3.1505
R10588 VDD.n2236 VDD.n2235 3.1505
R10589 VDD.n2240 VDD.n2239 3.1505
R10590 VDD.n2239 VDD.n2238 3.1505
R10591 VDD.n2243 VDD.n2242 3.1505
R10592 VDD.n2242 VDD.n2241 3.1505
R10593 VDD.n2246 VDD.n2245 3.1505
R10594 VDD.n2245 VDD.n2244 3.1505
R10595 VDD.n2249 VDD.n2248 3.1505
R10596 VDD.n2248 VDD.n2247 3.1505
R10597 VDD.n2252 VDD.n2251 3.1505
R10598 VDD.n2251 VDD.n2250 3.1505
R10599 VDD.n2255 VDD.n2254 3.1505
R10600 VDD.n2254 VDD.n2253 3.1505
R10601 VDD.n2258 VDD.n2257 3.1505
R10602 VDD.n2257 VDD.n2256 3.1505
R10603 VDD.n2261 VDD.n2260 3.1505
R10604 VDD.n2260 VDD.n2259 3.1505
R10605 VDD.n2264 VDD.n2263 3.1505
R10606 VDD.n2263 VDD.n2262 3.1505
R10607 VDD.n2267 VDD.n2266 3.1505
R10608 VDD.n2266 VDD.n2265 3.1505
R10609 VDD.n2270 VDD.n2269 3.1505
R10610 VDD.n2269 VDD.n2268 3.1505
R10611 VDD.n2273 VDD.n2272 3.1505
R10612 VDD.n2272 VDD.n2271 3.1505
R10613 VDD.n2276 VDD.n2275 3.1505
R10614 VDD.n2275 VDD.n2274 3.1505
R10615 VDD.n2279 VDD.n2278 3.1505
R10616 VDD.n2278 VDD.n2277 3.1505
R10617 VDD.n2282 VDD.n2281 3.1505
R10618 VDD.n2281 VDD.n2280 3.1505
R10619 VDD.n2285 VDD.n2284 3.1505
R10620 VDD.n2284 VDD.n2283 3.1505
R10621 VDD.n2288 VDD.n2287 3.1505
R10622 VDD.n2287 VDD.n2286 3.1505
R10623 VDD.n2291 VDD.n2290 3.1505
R10624 VDD.n2290 VDD.n2289 3.1505
R10625 VDD.n2294 VDD.n2293 3.1505
R10626 VDD.n2293 VDD.n2292 3.1505
R10627 VDD.n2297 VDD.n2296 3.1505
R10628 VDD.n2296 VDD.n2295 3.1505
R10629 VDD.n2300 VDD.n2299 3.1505
R10630 VDD.n2299 VDD.n2298 3.1505
R10631 VDD.n2303 VDD.n2302 3.1505
R10632 VDD.n2302 VDD.n2301 3.1505
R10633 VDD.n2306 VDD.n2305 3.1505
R10634 VDD.n2305 VDD.n2304 3.1505
R10635 VDD.n2309 VDD.n2308 3.1505
R10636 VDD.n2308 VDD.n2307 3.1505
R10637 VDD.n2312 VDD.n2311 3.1505
R10638 VDD.n2311 VDD.n2310 3.1505
R10639 VDD.n2316 VDD.n2315 3.1505
R10640 VDD.n2315 VDD.n2314 3.1505
R10641 VDD.n2319 VDD.n2318 3.1505
R10642 VDD.n2318 VDD.n2317 3.1505
R10643 VDD.n2322 VDD.n2321 3.1505
R10644 VDD.n2321 VDD.n2320 3.1505
R10645 VDD.n2325 VDD.n2324 3.1505
R10646 VDD.n2324 VDD.n2323 3.1505
R10647 VDD.n2328 VDD.n2327 3.1505
R10648 VDD.n2327 VDD.n2326 3.1505
R10649 VDD.n2331 VDD.n2330 3.1505
R10650 VDD.n2330 VDD.n2329 3.1505
R10651 VDD.n2334 VDD.n2333 3.1505
R10652 VDD.n2333 VDD.n2332 3.1505
R10653 VDD.n2346 VDD.n2345 3.1505
R10654 VDD.n2345 VDD.n2344 3.1505
R10655 VDD.n2349 VDD.n2348 3.1505
R10656 VDD.n2348 VDD.n2347 3.1505
R10657 VDD.n2352 VDD.n2351 3.1505
R10658 VDD.n2351 VDD.n2350 3.1505
R10659 VDD.n2355 VDD.n2354 3.1505
R10660 VDD.n2354 VDD.n2353 3.1505
R10661 VDD.n2358 VDD.n2357 3.1505
R10662 VDD.n2357 VDD.n2356 3.1505
R10663 VDD.n2361 VDD.n2360 3.1505
R10664 VDD.n2360 VDD.n2359 3.1505
R10665 VDD.n2365 VDD.n2364 3.1505
R10666 VDD.n2364 VDD.n2363 3.1505
R10667 VDD.n2369 VDD.n2368 3.1505
R10668 VDD.n2368 VDD.n2367 3.1505
R10669 VDD.n2373 VDD.n2372 3.1505
R10670 VDD.n2372 VDD.n2371 3.1505
R10671 VDD.n2377 VDD.n2376 3.1505
R10672 VDD.n2376 VDD.n2375 3.1505
R10673 VDD.n2380 VDD.n2379 3.1505
R10674 VDD.n2379 VDD.n2378 3.1505
R10675 VDD.n2384 VDD.n2383 3.1505
R10676 VDD.n2383 VDD.n2382 3.1505
R10677 VDD.n2388 VDD.n2387 3.1505
R10678 VDD.n2387 VDD.n2386 3.1505
R10679 VDD.n2392 VDD.n2391 3.1505
R10680 VDD.n2391 VDD.n2390 3.1505
R10681 VDD.n2395 VDD.n2394 3.1505
R10682 VDD.n2394 VDD.n2393 3.1505
R10683 VDD.n2399 VDD.n2398 3.1505
R10684 VDD.n2398 VDD.n2397 3.1505
R10685 VDD.n2402 VDD.n2401 3.1505
R10686 VDD.n2401 VDD.n2400 3.1505
R10687 VDD.n2405 VDD.n2404 3.1505
R10688 VDD.n2404 VDD.n2403 3.1505
R10689 VDD.n2408 VDD.n2407 3.1505
R10690 VDD.n2407 VDD.n2406 3.1505
R10691 VDD.n2413 VDD.n2412 3.1505
R10692 VDD.n2412 VDD.n2411 3.1505
R10693 VDD.n2416 VDD.n2415 3.1505
R10694 VDD.n2415 VDD.n2414 3.1505
R10695 VDD.n2419 VDD.n2418 3.1505
R10696 VDD.n2418 VDD.n2417 3.1505
R10697 VDD.n2423 VDD.n2422 3.1505
R10698 VDD.n2422 VDD.n2421 3.1505
R10699 VDD.n2426 VDD.n2425 3.1505
R10700 VDD.n2425 VDD.n2424 3.1505
R10701 VDD.n2430 VDD.n2429 3.1505
R10702 VDD.n2429 VDD.n2428 3.1505
R10703 VDD.n2433 VDD.n2432 3.1505
R10704 VDD.n2432 VDD.n2431 3.1505
R10705 VDD.n2437 VDD.n2436 3.1505
R10706 VDD.n2436 VDD.n2435 3.1505
R10707 VDD.n2440 VDD.n2439 3.1505
R10708 VDD.n2439 VDD.n2438 3.1505
R10709 VDD.n2443 VDD.n2442 3.1505
R10710 VDD.n2442 VDD.n2441 3.1505
R10711 VDD.n2448 VDD.n2447 3.1505
R10712 VDD.n2447 VDD.n2446 3.1505
R10713 VDD.n2451 VDD.n2450 3.1505
R10714 VDD.n2450 VDD.n2449 3.1505
R10715 VDD.n2454 VDD.n2453 3.1505
R10716 VDD.n2453 VDD.n2452 3.1505
R10717 VDD.n2458 VDD.n2457 3.1505
R10718 VDD.n2457 VDD.n2456 3.1505
R10719 VDD.n2461 VDD.n2460 3.1505
R10720 VDD.n2460 VDD.n2459 3.1505
R10721 VDD.n2465 VDD.n2464 3.1505
R10722 VDD.n2464 VDD.n2463 3.1505
R10723 VDD.n2468 VDD.n2467 3.1505
R10724 VDD.n2467 VDD.n2466 3.1505
R10725 VDD.n2472 VDD.n2471 3.1505
R10726 VDD.n2471 VDD.n2470 3.1505
R10727 VDD.n2475 VDD.n2474 3.1505
R10728 VDD.n2474 VDD.n2473 3.1505
R10729 VDD.n2478 VDD.n2477 3.1505
R10730 VDD.n2477 VDD.n2476 3.1505
R10731 VDD.n2482 VDD.n2481 3.1505
R10732 VDD.n2481 VDD.n2480 3.1505
R10733 VDD.n2486 VDD.n2485 3.1505
R10734 VDD.n2485 VDD.n2484 3.1505
R10735 VDD.n2489 VDD.n2488 3.1505
R10736 VDD.n2488 VDD.n2487 3.1505
R10737 VDD.n2492 VDD.n2491 3.1505
R10738 VDD.n2491 VDD.n2490 3.1505
R10739 VDD.n2496 VDD.n2495 3.1505
R10740 VDD.n2495 VDD.n2494 3.1505
R10741 VDD.n2500 VDD.n2499 3.1505
R10742 VDD.n2499 VDD.n2498 3.1505
R10743 VDD.n2504 VDD.n2503 3.1505
R10744 VDD.n2503 VDD.n2502 3.1505
R10745 VDD.n2507 VDD.n2506 3.1505
R10746 VDD.n2506 VDD.n2505 3.1505
R10747 VDD.n2510 VDD.n2509 3.1505
R10748 VDD.n2509 VDD.n2508 3.1505
R10749 VDD.n2513 VDD.n2512 3.1505
R10750 VDD.n2512 VDD.n2511 3.1505
R10751 VDD.n2516 VDD.n2515 3.1505
R10752 VDD.n2515 VDD.n2514 3.1505
R10753 VDD.n4665 VDD.n4664 3.1505
R10754 VDD.n4664 VDD.n4663 3.1505
R10755 VDD.n4662 VDD.n4661 3.1505
R10756 VDD.n4661 VDD.n4660 3.1505
R10757 VDD.n4659 VDD.n4658 3.1505
R10758 VDD.n4658 VDD.n4657 3.1505
R10759 VDD.n4656 VDD.n4655 3.1505
R10760 VDD.n4655 VDD.n4654 3.1505
R10761 VDD.n4652 VDD.n4651 3.1505
R10762 VDD.n4651 VDD.n4650 3.1505
R10763 VDD.n4649 VDD.n4648 3.1505
R10764 VDD.n4648 VDD.n4647 3.1505
R10765 VDD.n4645 VDD.n4644 3.1505
R10766 VDD.n4644 VDD.n4643 3.1505
R10767 VDD.n4642 VDD.n4641 3.1505
R10768 VDD.n4641 VDD.n4640 3.1505
R10769 VDD.n4639 VDD.n4638 3.1505
R10770 VDD.n4638 VDD.n4637 3.1505
R10771 VDD.n4635 VDD.n4634 3.1505
R10772 VDD.n4634 VDD.n4633 3.1505
R10773 VDD.n4632 VDD.n4631 3.1505
R10774 VDD.n4631 VDD.n4630 3.1505
R10775 VDD.n4629 VDD.n4628 3.1505
R10776 VDD.n4628 VDD.n4627 3.1505
R10777 VDD.n4625 VDD.n4624 3.1505
R10778 VDD.n4624 VDD.n4623 3.1505
R10779 VDD.n4622 VDD.n4621 3.1505
R10780 VDD.n4621 VDD.n4620 3.1505
R10781 VDD.n4619 VDD.n4618 3.1505
R10782 VDD.n4618 VDD.n4617 3.1505
R10783 VDD.n4615 VDD.n4614 3.1505
R10784 VDD.n4614 VDD.n4613 3.1505
R10785 VDD.n4612 VDD.n4611 3.1505
R10786 VDD.n4611 VDD.n4610 3.1505
R10787 VDD.n4609 VDD.n4608 3.1505
R10788 VDD.n4608 VDD.n4607 3.1505
R10789 VDD.n4606 VDD.n4605 3.1505
R10790 VDD.n4605 VDD.n4604 3.1505
R10791 VDD.n4602 VDD.n4601 3.1505
R10792 VDD.n4601 VDD.n4600 3.1505
R10793 VDD.n4599 VDD.n4598 3.1505
R10794 VDD.n4598 VDD.n4597 3.1505
R10795 VDD.n4596 VDD.n4595 3.1505
R10796 VDD.n4595 VDD.n4594 3.1505
R10797 VDD.n4592 VDD.n4591 3.1505
R10798 VDD.n4591 VDD.n4590 3.1505
R10799 VDD.n4589 VDD.n4588 3.1505
R10800 VDD.n4588 VDD.n4587 3.1505
R10801 VDD.n4586 VDD.n4585 3.1505
R10802 VDD.n4585 VDD.n4584 3.1505
R10803 VDD.n4583 VDD.n4582 3.1505
R10804 VDD.n4582 VDD.n4581 3.1505
R10805 VDD.n4579 VDD.n4578 3.1505
R10806 VDD.n4578 VDD.n4577 3.1505
R10807 VDD.n4576 VDD.n4575 3.1505
R10808 VDD.n4575 VDD.n4574 3.1505
R10809 VDD.n4573 VDD.n4572 3.1505
R10810 VDD.n4572 VDD.n4571 3.1505
R10811 VDD.n4569 VDD.n4568 3.1505
R10812 VDD.n4568 VDD.n4567 3.1505
R10813 VDD.n4566 VDD.n4565 3.1505
R10814 VDD.n4565 VDD.n4564 3.1505
R10815 VDD.n4563 VDD.n4562 3.1505
R10816 VDD.n4562 VDD.n4561 3.1505
R10817 VDD.n4559 VDD.n4558 3.1505
R10818 VDD.n4558 VDD.n4557 3.1505
R10819 VDD.n4556 VDD.n4555 3.1505
R10820 VDD.n4555 VDD.n4554 3.1505
R10821 VDD.n4553 VDD.n4552 3.1505
R10822 VDD.n4552 VDD.n4551 3.1505
R10823 VDD.n4549 VDD.n4548 3.1505
R10824 VDD.n4548 VDD.n4547 3.1505
R10825 VDD.n4546 VDD.n4545 3.1505
R10826 VDD.n4545 VDD.n4544 3.1505
R10827 VDD.n4542 VDD.n4541 3.1505
R10828 VDD.n4541 VDD.n4540 3.1505
R10829 VDD.n4539 VDD.n4538 3.1505
R10830 VDD.n4538 VDD.n4537 3.1505
R10831 VDD.n4536 VDD.n4535 3.1505
R10832 VDD.n4535 VDD.n4534 3.1505
R10833 VDD.n4533 VDD.n4532 3.1505
R10834 VDD.n4532 VDD.n4531 3.1505
R10835 VDD.n4529 VDD.n4528 3.1505
R10836 VDD.n4528 VDD.n4527 3.1505
R10837 VDD.n4523 VDD.n4522 3.1505
R10838 VDD.n4499 VDD.n4498 3.1505
R10839 VDD.n4498 VDD.n4497 3.1505
R10840 VDD.n4496 VDD.n4495 3.1505
R10841 VDD.n4495 VDD.n4494 3.1505
R10842 VDD.n4493 VDD.n4492 3.1505
R10843 VDD.n4492 VDD.n4491 3.1505
R10844 VDD.n4490 VDD.n4489 3.1505
R10845 VDD.n4489 VDD.n4488 3.1505
R10846 VDD.n4487 VDD.n4486 3.1505
R10847 VDD.n4486 VDD.n4485 3.1505
R10848 VDD.n4483 VDD.n4482 3.1505
R10849 VDD.n4482 VDD.n4481 3.1505
R10850 VDD.n4480 VDD.n4479 3.1505
R10851 VDD.n4479 VDD.n4478 3.1505
R10852 VDD.n4476 VDD.n4475 3.1505
R10853 VDD.n4475 VDD.n4474 3.1505
R10854 VDD.n4473 VDD.n4472 3.1505
R10855 VDD.n4472 VDD.n4471 3.1505
R10856 VDD.n4470 VDD.n4469 3.1505
R10857 VDD.n4469 VDD.n4468 3.1505
R10858 VDD.n4466 VDD.n4465 3.1505
R10859 VDD.n4465 VDD.n4464 3.1505
R10860 VDD.n4463 VDD.n4462 3.1505
R10861 VDD.n4462 VDD.n4461 3.1505
R10862 VDD.n4460 VDD.n4459 3.1505
R10863 VDD.n4459 VDD.n4458 3.1505
R10864 VDD.n4456 VDD.n4455 3.1505
R10865 VDD.n4455 VDD.n4454 3.1505
R10866 VDD.n4453 VDD.n4452 3.1505
R10867 VDD.n4452 VDD.n4451 3.1505
R10868 VDD.n4450 VDD.n4449 3.1505
R10869 VDD.n4449 VDD.n4448 3.1505
R10870 VDD.n4446 VDD.n4445 3.1505
R10871 VDD.n4445 VDD.n4444 3.1505
R10872 VDD.n4443 VDD.n4442 3.1505
R10873 VDD.n4442 VDD.n4441 3.1505
R10874 VDD.n4440 VDD.n4439 3.1505
R10875 VDD.n4439 VDD.n4438 3.1505
R10876 VDD.n4437 VDD.n4436 3.1505
R10877 VDD.n4436 VDD.n4435 3.1505
R10878 VDD.n4433 VDD.n4432 3.1505
R10879 VDD.n4432 VDD.n4431 3.1505
R10880 VDD.n4430 VDD.n4429 3.1505
R10881 VDD.n4429 VDD.n4428 3.1505
R10882 VDD.n4427 VDD.n4426 3.1505
R10883 VDD.n4426 VDD.n4425 3.1505
R10884 VDD.n4423 VDD.n4422 3.1505
R10885 VDD.n4422 VDD.n4421 3.1505
R10886 VDD.n4420 VDD.n4419 3.1505
R10887 VDD.n4419 VDD.n4418 3.1505
R10888 VDD.n4417 VDD.n4416 3.1505
R10889 VDD.n4416 VDD.n4415 3.1505
R10890 VDD.n4414 VDD.n4413 3.1505
R10891 VDD.n4413 VDD.n4412 3.1505
R10892 VDD.n4410 VDD.n4409 3.1505
R10893 VDD.n4409 VDD.n4408 3.1505
R10894 VDD.n4407 VDD.n4406 3.1505
R10895 VDD.n4406 VDD.n4405 3.1505
R10896 VDD.n4404 VDD.n4403 3.1505
R10897 VDD.n4403 VDD.n4402 3.1505
R10898 VDD.n4400 VDD.n4399 3.1505
R10899 VDD.n4399 VDD.n4398 3.1505
R10900 VDD.n4397 VDD.n4396 3.1505
R10901 VDD.n4396 VDD.n4395 3.1505
R10902 VDD.n4394 VDD.n4393 3.1505
R10903 VDD.n4393 VDD.n4392 3.1505
R10904 VDD.n4390 VDD.n4389 3.1505
R10905 VDD.n4389 VDD.n4388 3.1505
R10906 VDD.n4387 VDD.n4386 3.1505
R10907 VDD.n4386 VDD.n4385 3.1505
R10908 VDD.n4384 VDD.n4383 3.1505
R10909 VDD.n4383 VDD.n4382 3.1505
R10910 VDD.n4380 VDD.n4379 3.1505
R10911 VDD.n4379 VDD.n4378 3.1505
R10912 VDD.n4377 VDD.n4376 3.1505
R10913 VDD.n4376 VDD.n4375 3.1505
R10914 VDD.n4370 VDD.n4369 3.1505
R10915 VDD.n4369 VDD.n4368 3.1505
R10916 VDD.n4367 VDD.n4366 3.1505
R10917 VDD.n4366 VDD.n4365 3.1505
R10918 VDD.n4364 VDD.n4363 3.1505
R10919 VDD.n4363 VDD.n4362 3.1505
R10920 VDD.n4361 VDD.n4360 3.1505
R10921 VDD.n4360 VDD.n4359 3.1505
R10922 VDD.n4358 VDD.n4357 3.1505
R10923 VDD.n4357 VDD.n4356 3.1505
R10924 VDD.n4353 VDD.n4352 3.1505
R10925 VDD.n5753 VDD.n5752 3.1505
R10926 VDD.n5755 VDD.n5754 3.1505
R10927 VDD.n5757 VDD.n5756 3.1505
R10928 VDD.n5759 VDD.n5758 3.1505
R10929 VDD.n5761 VDD.n5760 3.1505
R10930 VDD.n5764 VDD.n5763 3.1505
R10931 VDD.n5766 VDD.n5765 3.1505
R10932 VDD.n5769 VDD.n5768 3.1505
R10933 VDD.n5771 VDD.n5770 3.1505
R10934 VDD.n5773 VDD.n5772 3.1505
R10935 VDD.n5776 VDD.n5775 3.1505
R10936 VDD.n5778 VDD.n5777 3.1505
R10937 VDD.n5780 VDD.n5779 3.1505
R10938 VDD.n5783 VDD.n5782 3.1505
R10939 VDD.n5785 VDD.n5784 3.1505
R10940 VDD.n5787 VDD.n5786 3.1505
R10941 VDD.n5790 VDD.n5789 3.1505
R10942 VDD.n5792 VDD.n5791 3.1505
R10943 VDD.n5794 VDD.n5793 3.1505
R10944 VDD.n5796 VDD.n5795 3.1505
R10945 VDD.n5798 VDD.n5797 3.1505
R10946 VDD.n5800 VDD.n5799 3.1505
R10947 VDD.n5802 VDD.n5801 3.1505
R10948 VDD.n5804 VDD.n5803 3.1505
R10949 VDD.n5806 VDD.n5805 3.1505
R10950 VDD.n5808 VDD.n5807 3.1505
R10951 VDD.n5810 VDD.n5809 3.1505
R10952 VDD.n5813 VDD.n5812 3.1505
R10953 VDD.n5815 VDD.n5814 3.1505
R10954 VDD.n5817 VDD.n5816 3.1505
R10955 VDD.n5820 VDD.n5819 3.1505
R10956 VDD.n5822 VDD.n5821 3.1505
R10957 VDD.n5824 VDD.n5823 3.1505
R10958 VDD.n5827 VDD.n5826 3.1505
R10959 VDD.n5829 VDD.n5828 3.1505
R10960 VDD.n5831 VDD.n5830 3.1505
R10961 VDD.n5834 VDD.n5833 3.1505
R10962 VDD.n5836 VDD.n5835 3.1505
R10963 VDD.n5839 VDD.n5838 3.1505
R10964 VDD.n5841 VDD.n5840 3.1505
R10965 VDD.n5843 VDD.n5842 3.1505
R10966 VDD.n5845 VDD.n5844 3.1505
R10967 VDD.n5647 VDD.n5646 3.1505
R10968 VDD.n5649 VDD.n5648 3.1505
R10969 VDD.n5651 VDD.n5650 3.1505
R10970 VDD.n5653 VDD.n5652 3.1505
R10971 VDD.n5655 VDD.n5654 3.1505
R10972 VDD.n5658 VDD.n5657 3.1505
R10973 VDD.n5660 VDD.n5659 3.1505
R10974 VDD.n5663 VDD.n5662 3.1505
R10975 VDD.n5665 VDD.n5664 3.1505
R10976 VDD.n5667 VDD.n5666 3.1505
R10977 VDD.n5670 VDD.n5669 3.1505
R10978 VDD.n5672 VDD.n5671 3.1505
R10979 VDD.n5674 VDD.n5673 3.1505
R10980 VDD.n5677 VDD.n5676 3.1505
R10981 VDD.n5679 VDD.n5678 3.1505
R10982 VDD.n5681 VDD.n5680 3.1505
R10983 VDD.n5684 VDD.n5683 3.1505
R10984 VDD.n5686 VDD.n5685 3.1505
R10985 VDD.n5688 VDD.n5687 3.1505
R10986 VDD.n5690 VDD.n5689 3.1505
R10987 VDD.n5692 VDD.n5691 3.1505
R10988 VDD.n5694 VDD.n5693 3.1505
R10989 VDD.n5696 VDD.n5695 3.1505
R10990 VDD.n5698 VDD.n5697 3.1505
R10991 VDD.n5700 VDD.n5699 3.1505
R10992 VDD.n5702 VDD.n5701 3.1505
R10993 VDD.n5704 VDD.n5703 3.1505
R10994 VDD.n5707 VDD.n5706 3.1505
R10995 VDD.n5709 VDD.n5708 3.1505
R10996 VDD.n5711 VDD.n5710 3.1505
R10997 VDD.n5714 VDD.n5713 3.1505
R10998 VDD.n5716 VDD.n5715 3.1505
R10999 VDD.n5718 VDD.n5717 3.1505
R11000 VDD.n5721 VDD.n5720 3.1505
R11001 VDD.n5723 VDD.n5722 3.1505
R11002 VDD.n5725 VDD.n5724 3.1505
R11003 VDD.n5728 VDD.n5727 3.1505
R11004 VDD.n5730 VDD.n5729 3.1505
R11005 VDD.n5733 VDD.n5732 3.1505
R11006 VDD.n5735 VDD.n5734 3.1505
R11007 VDD.n5737 VDD.n5736 3.1505
R11008 VDD.n5739 VDD.n5738 3.1505
R11009 VDD.n5741 VDD.n5740 3.1505
R11010 VDD.n308 VDD.t350 3.08583
R11011 VDD.n304 VDD.t396 3.08583
R11012 VDD.n303 VDD.t209 3.08583
R11013 VDD.n16 VDD.t166 3.08583
R11014 VDD.n17 VDD.t238 3.08583
R11015 VDD.n18 VDD.t330 3.08583
R11016 VDD.n6863 VDD.t266 3.08583
R11017 VDD.n6859 VDD.t340 3.08583
R11018 VDD.n6858 VDD.t388 3.08583
R11019 VDD.n22 VDD.t269 3.08583
R11020 VDD.n23 VDD.t344 3.08583
R11021 VDD.n24 VDD.t390 3.08583
R11022 VDD.n2068 VDD.t430 3.07932
R11023 VDD.n2226 VDD.t32 3.07932
R11024 VDD.n2310 VDD.t86 3.07932
R11025 VDD.n2428 VDD.t403 3.07932
R11026 VDD.n7959 VDD.t252 3.0555
R11027 VDD.n392 VDD.t392 3.0555
R11028 VDD.n7974 VDD.t186 3.0555
R11029 VDD.n7193 VDD.t218 2.97991
R11030 VDD.n6451 VDD.n6448 2.93268
R11031 VDD.n6150 VDD.n6149 2.87353
R11032 VDD.n2684 VDD.n2683 2.87353
R11033 VDD.n4425 VDD.t726 2.8495
R11034 VDD.n4431 VDD.t712 2.8495
R11035 VDD.n4896 VDD.t721 2.8495
R11036 VDD.n4902 VDD.t650 2.8495
R11037 VDD.n5043 VDD.t714 2.8495
R11038 VDD.n5049 VDD.t729 2.8495
R11039 VDD.n4594 VDD.t636 2.8495
R11040 VDD.n4600 VDD.t719 2.8495
R11041 VDD.n4741 VDD.t641 2.8495
R11042 VDD.n4747 VDD.t657 2.8495
R11043 VDD.n5198 VDD.t661 2.8495
R11044 VDD.n5204 VDD.t644 2.8495
R11045 VDD.n6520 VDD.t646 2.8495
R11046 VDD.n6526 VDD.t639 2.8495
R11047 VDD.n2235 VDD.t478 2.66881
R11048 VDD.n2435 VDD.t67 2.66881
R11049 VDD.n338 VDD.t262 2.6092
R11050 VDD.n345 VDD.t504 2.6092
R11051 VDD.n364 VDD.t436 2.6092
R11052 VDD.n361 VDD.t56 2.6092
R11053 VDD.n4237 VDD.n4236 2.6005
R11054 VDD.n4234 VDD.n4233 2.6005
R11055 VDD.n5620 VDD.n5619 2.6005
R11056 VDD.n5621 VDD.n5617 2.6005
R11057 VDD.n4231 VDD.n4230 2.6005
R11058 VDD.n4228 VDD.n4227 2.6005
R11059 VDD.n5614 VDD.n5613 2.6005
R11060 VDD.n5615 VDD.n5611 2.6005
R11061 VDD.n4225 VDD.n4224 2.6005
R11062 VDD.n4222 VDD.n4221 2.6005
R11063 VDD.n5608 VDD.n5607 2.6005
R11064 VDD.n5609 VDD.n5605 2.6005
R11065 VDD.n5603 VDD.n5593 2.6005
R11066 VDD.n5601 VDD.n5600 2.6005
R11067 VDD.n4206 VDD.n4205 2.6005
R11068 VDD.n4215 VDD.n4214 2.6005
R11069 VDD.n4197 VDD.n4196 2.6005
R11070 VDD.n4194 VDD.n4193 2.6005
R11071 VDD.n5590 VDD.n5589 2.6005
R11072 VDD.n5591 VDD.n5587 2.6005
R11073 VDD.n4191 VDD.n4190 2.6005
R11074 VDD.n4188 VDD.n4187 2.6005
R11075 VDD.n5584 VDD.n5583 2.6005
R11076 VDD.n5585 VDD.n5581 2.6005
R11077 VDD.n3945 VDD.n3944 2.6005
R11078 VDD.n3942 VDD.n3941 2.6005
R11079 VDD.n5536 VDD.n5535 2.6005
R11080 VDD.n5537 VDD.n5533 2.6005
R11081 VDD.n3939 VDD.n3938 2.6005
R11082 VDD.n3936 VDD.n3935 2.6005
R11083 VDD.n5530 VDD.n5529 2.6005
R11084 VDD.n5531 VDD.n5527 2.6005
R11085 VDD.n5525 VDD.n5515 2.6005
R11086 VDD.n5523 VDD.n5522 2.6005
R11087 VDD.n3924 VDD.n3923 2.6005
R11088 VDD.n3933 VDD.n3932 2.6005
R11089 VDD.n3911 VDD.n3910 2.6005
R11090 VDD.n3908 VDD.n3907 2.6005
R11091 VDD.n5512 VDD.n5511 2.6005
R11092 VDD.n5513 VDD.n5509 2.6005
R11093 VDD.n3905 VDD.n3904 2.6005
R11094 VDD.n3902 VDD.n3901 2.6005
R11095 VDD.n5506 VDD.n5505 2.6005
R11096 VDD.n5507 VDD.n5503 2.6005
R11097 VDD.n3899 VDD.n3898 2.6005
R11098 VDD.n3896 VDD.n3895 2.6005
R11099 VDD.n5500 VDD.n5499 2.6005
R11100 VDD.n5501 VDD.n5497 2.6005
R11101 VDD.n3399 VDD.n3398 2.6005
R11102 VDD.n3396 VDD.n3395 2.6005
R11103 VDD.n5354 VDD.n5353 2.6005
R11104 VDD.n5355 VDD.n5351 2.6005
R11105 VDD.n3405 VDD.n3404 2.6005
R11106 VDD.n3402 VDD.n3401 2.6005
R11107 VDD.n5360 VDD.n5359 2.6005
R11108 VDD.n5361 VDD.n5357 2.6005
R11109 VDD.n3411 VDD.n3410 2.6005
R11110 VDD.n3408 VDD.n3407 2.6005
R11111 VDD.n5366 VDD.n5365 2.6005
R11112 VDD.n5367 VDD.n5363 2.6005
R11113 VDD.n3433 VDD.n3432 2.6005
R11114 VDD.n3429 VDD.n3428 2.6005
R11115 VDD.n5372 VDD.n5371 2.6005
R11116 VDD.n5379 VDD.n5369 2.6005
R11117 VDD.n3439 VDD.n3438 2.6005
R11118 VDD.n3436 VDD.n3435 2.6005
R11119 VDD.n5384 VDD.n5383 2.6005
R11120 VDD.n5385 VDD.n5381 2.6005
R11121 VDD.n3445 VDD.n3444 2.6005
R11122 VDD.n3442 VDD.n3441 2.6005
R11123 VDD.n5390 VDD.n5389 2.6005
R11124 VDD.n5391 VDD.n5387 2.6005
R11125 VDD.n3713 VDD.n3712 2.6005
R11126 VDD.n3710 VDD.n3709 2.6005
R11127 VDD.n5431 VDD.n5430 2.6005
R11128 VDD.n5432 VDD.n5428 2.6005
R11129 VDD.n3719 VDD.n3718 2.6005
R11130 VDD.n3716 VDD.n3715 2.6005
R11131 VDD.n5437 VDD.n5436 2.6005
R11132 VDD.n5438 VDD.n5434 2.6005
R11133 VDD.n3737 VDD.n3736 2.6005
R11134 VDD.n3733 VDD.n3732 2.6005
R11135 VDD.n5443 VDD.n5442 2.6005
R11136 VDD.n5450 VDD.n5440 2.6005
R11137 VDD.n3747 VDD.n3746 2.6005
R11138 VDD.n3744 VDD.n3743 2.6005
R11139 VDD.n5455 VDD.n5454 2.6005
R11140 VDD.n5456 VDD.n5452 2.6005
R11141 VDD.n3753 VDD.n3752 2.6005
R11142 VDD.n3750 VDD.n3749 2.6005
R11143 VDD.n5461 VDD.n5460 2.6005
R11144 VDD.n5462 VDD.n5458 2.6005
R11145 VDD.n3759 VDD.n3758 2.6005
R11146 VDD.n3756 VDD.n3755 2.6005
R11147 VDD.n5467 VDD.n5466 2.6005
R11148 VDD.n5468 VDD.n5464 2.6005
R11149 VDD.n2910 VDD.n2909 2.6005
R11150 VDD.n2907 VDD.n2906 2.6005
R11151 VDD.n6204 VDD.n6203 2.6005
R11152 VDD.n6205 VDD.n6201 2.6005
R11153 VDD.n2916 VDD.n2915 2.6005
R11154 VDD.n2913 VDD.n2912 2.6005
R11155 VDD.n6198 VDD.n6197 2.6005
R11156 VDD.n6199 VDD.n6195 2.6005
R11157 VDD.n2922 VDD.n2921 2.6005
R11158 VDD.n2919 VDD.n2918 2.6005
R11159 VDD.n6192 VDD.n6191 2.6005
R11160 VDD.n6193 VDD.n6189 2.6005
R11161 VDD.n2944 VDD.n2943 2.6005
R11162 VDD.n2940 VDD.n2939 2.6005
R11163 VDD.n6180 VDD.n6179 2.6005
R11164 VDD.n6187 VDD.n6177 2.6005
R11165 VDD.n2950 VDD.n2949 2.6005
R11166 VDD.n2947 VDD.n2946 2.6005
R11167 VDD.n6174 VDD.n6173 2.6005
R11168 VDD.n6175 VDD.n6171 2.6005
R11169 VDD.n2956 VDD.n2955 2.6005
R11170 VDD.n2953 VDD.n2952 2.6005
R11171 VDD.n6168 VDD.n6167 2.6005
R11172 VDD.n6169 VDD.n6165 2.6005
R11173 VDD.n3209 VDD.n3208 2.6005
R11174 VDD.n3206 VDD.n3205 2.6005
R11175 VDD.n5294 VDD.n5293 2.6005
R11176 VDD.n5295 VDD.n5291 2.6005
R11177 VDD.n3215 VDD.n3214 2.6005
R11178 VDD.n3212 VDD.n3211 2.6005
R11179 VDD.n5300 VDD.n5299 2.6005
R11180 VDD.n5301 VDD.n5297 2.6005
R11181 VDD.n3233 VDD.n3232 2.6005
R11182 VDD.n3229 VDD.n3228 2.6005
R11183 VDD.n5306 VDD.n5305 2.6005
R11184 VDD.n5313 VDD.n5303 2.6005
R11185 VDD.n3243 VDD.n3242 2.6005
R11186 VDD.n3240 VDD.n3239 2.6005
R11187 VDD.n5318 VDD.n5317 2.6005
R11188 VDD.n5319 VDD.n5315 2.6005
R11189 VDD.n3249 VDD.n3248 2.6005
R11190 VDD.n3246 VDD.n3245 2.6005
R11191 VDD.n5324 VDD.n5323 2.6005
R11192 VDD.n5325 VDD.n5321 2.6005
R11193 VDD.n3255 VDD.n3254 2.6005
R11194 VDD.n3252 VDD.n3251 2.6005
R11195 VDD.n5330 VDD.n5329 2.6005
R11196 VDD.n5331 VDD.n5327 2.6005
R11197 VDD.n2842 VDD.n2841 2.6005
R11198 VDD.n2839 VDD.n2838 2.6005
R11199 VDD.n2541 VDD.n2540 2.6005
R11200 VDD.n2542 VDD.n2538 2.6005
R11201 VDD.n2848 VDD.n2847 2.6005
R11202 VDD.n2845 VDD.n2844 2.6005
R11203 VDD.n2547 VDD.n2546 2.6005
R11204 VDD.n2548 VDD.n2544 2.6005
R11205 VDD.n2866 VDD.n2865 2.6005
R11206 VDD.n2862 VDD.n2861 2.6005
R11207 VDD.n2553 VDD.n2552 2.6005
R11208 VDD.n2560 VDD.n2550 2.6005
R11209 VDD.n2876 VDD.n2875 2.6005
R11210 VDD.n2873 VDD.n2872 2.6005
R11211 VDD.n2565 VDD.n2564 2.6005
R11212 VDD.n2566 VDD.n2562 2.6005
R11213 VDD.n2882 VDD.n2881 2.6005
R11214 VDD.n2879 VDD.n2878 2.6005
R11215 VDD.n2571 VDD.n2570 2.6005
R11216 VDD.n2572 VDD.n2568 2.6005
R11217 VDD.n2888 VDD.n2887 2.6005
R11218 VDD.n2885 VDD.n2884 2.6005
R11219 VDD.n2577 VDD.n2576 2.6005
R11220 VDD.n2578 VDD.n2574 2.6005
R11221 VDD.n746 VDD.n745 2.6005
R11222 VDD.n743 VDD.n742 2.6005
R11223 VDD.n740 VDD.n739 2.6005
R11224 VDD.n567 VDD.n566 2.6005
R11225 VDD.n755 VDD.n754 2.6005
R11226 VDD.n752 VDD.n751 2.6005
R11227 VDD.n749 VDD.n748 2.6005
R11228 VDD.n570 VDD.n569 2.6005
R11229 VDD.n1055 VDD.n1054 2.6005
R11230 VDD.n1052 VDD.n1051 2.6005
R11231 VDD.n1049 VDD.n1048 2.6005
R11232 VDD.n879 VDD.n878 2.6005
R11233 VDD.n1046 VDD.n1045 2.6005
R11234 VDD.n1043 VDD.n1042 2.6005
R11235 VDD.n1040 VDD.n1039 2.6005
R11236 VDD.n876 VDD.n875 2.6005
R11237 VDD.n8159 VDD.n8158 2.6005
R11238 VDD.n8162 VDD.n8161 2.6005
R11239 VDD.n8165 VDD.n8164 2.6005
R11240 VDD.n8148 VDD.n8147 2.6005
R11241 VDD.n8151 VDD.n8150 2.6005
R11242 VDD.n8154 VDD.n8153 2.6005
R11243 VDD.n7897 VDD.n7896 2.6005
R11244 VDD.n7900 VDD.n7899 2.6005
R11245 VDD.n7903 VDD.n7902 2.6005
R11246 VDD.n11 VDD.n1 2.6005
R11247 VDD.n10 VDD.n3 2.6005
R11248 VDD.n9 VDD.n5 2.6005
R11249 VDD.n7060 VDD.n7059 2.6005
R11250 VDD.n8321 VDD.n8319 2.6005
R11251 VDD.n8322 VDD.n8318 2.6005
R11252 VDD.n8323 VDD.n8317 2.6005
R11253 VDD.n7892 VDD.n7891 2.6005
R11254 VDD.n408 VDD.n407 2.6005
R11255 VDD.n1362 VDD.n1359 2.6005
R11256 VDD.n1363 VDD.n1357 2.6005
R11257 VDD.n1364 VDD.n1355 2.6005
R11258 VDD.n1373 VDD.n1370 2.6005
R11259 VDD.n1374 VDD.n1368 2.6005
R11260 VDD.n1375 VDD.n1366 2.6005
R11261 VDD.n1384 VDD.n1381 2.6005
R11262 VDD.n1385 VDD.n1379 2.6005
R11263 VDD.n1386 VDD.n1377 2.6005
R11264 VDD.n1395 VDD.n1392 2.6005
R11265 VDD.n1396 VDD.n1390 2.6005
R11266 VDD.n1397 VDD.n1388 2.6005
R11267 VDD.n1406 VDD.n1403 2.6005
R11268 VDD.n1407 VDD.n1401 2.6005
R11269 VDD.n1408 VDD.n1399 2.6005
R11270 VDD.n1417 VDD.n1414 2.6005
R11271 VDD.n1418 VDD.n1412 2.6005
R11272 VDD.n1419 VDD.n1410 2.6005
R11273 VDD.n1431 VDD.n1427 2.6005
R11274 VDD.n1430 VDD.n1429 2.6005
R11275 VDD.n1116 VDD.n1115 2.6005
R11276 VDD.n1119 VDD.n1118 2.6005
R11277 VDD.n1425 VDD.n1421 2.6005
R11278 VDD.n1424 VDD.n1423 2.6005
R11279 VDD.n1110 VDD.n1109 2.6005
R11280 VDD.n1113 VDD.n1112 2.6005
R11281 VDD.n1353 VDD.n1349 2.6005
R11282 VDD.n1104 VDD.n1103 2.6005
R11283 VDD.n1351 VDD.n1350 2.6005
R11284 VDD.n1107 VDD.n1106 2.6005
R11285 VDD.n2689 VDD.n2688 2.48924
R11286 VDD.n2692 VDD.n2691 2.48924
R11287 VDD.n2695 VDD.n2694 2.48924
R11288 VDD.n2698 VDD.n2697 2.48924
R11289 VDD.n2701 VDD.n2700 2.48924
R11290 VDD.n2704 VDD.n2703 2.48924
R11291 VDD.n2707 VDD.n2706 2.48924
R11292 VDD.n2710 VDD.n2709 2.48924
R11293 VDD.n2713 VDD.n2712 2.48924
R11294 VDD.n2716 VDD.n2715 2.48924
R11295 VDD.n2719 VDD.n2718 2.48924
R11296 VDD.n2722 VDD.n2721 2.48924
R11297 VDD.n2725 VDD.n2724 2.48924
R11298 VDD.n2728 VDD.n2727 2.48924
R11299 VDD.n2731 VDD.n2730 2.48924
R11300 VDD.n2734 VDD.n2733 2.48924
R11301 VDD.n2737 VDD.n2736 2.48924
R11302 VDD.n2740 VDD.n2739 2.48924
R11303 VDD.n2743 VDD.n2742 2.48924
R11304 VDD.n2746 VDD.n2745 2.48924
R11305 VDD.n2749 VDD.n2748 2.48924
R11306 VDD.n2752 VDD.n2751 2.48924
R11307 VDD.n2755 VDD.n2754 2.48924
R11308 VDD.n2758 VDD.n2757 2.48924
R11309 VDD.n2761 VDD.n2760 2.48924
R11310 VDD.n2764 VDD.n2763 2.48924
R11311 VDD.n2767 VDD.n2766 2.48924
R11312 VDD.n2770 VDD.n2769 2.48924
R11313 VDD.n2773 VDD.n2772 2.48924
R11314 VDD.n2776 VDD.n2775 2.48924
R11315 VDD.n2779 VDD.n2778 2.48924
R11316 VDD.n2782 VDD.n2781 2.48924
R11317 VDD.n2785 VDD.n2784 2.48924
R11318 VDD.n2788 VDD.n2787 2.48924
R11319 VDD.n2791 VDD.n2790 2.48924
R11320 VDD.n2794 VDD.n2793 2.48924
R11321 VDD.n2797 VDD.n2796 2.48924
R11322 VDD.n2800 VDD.n2799 2.48924
R11323 VDD.n2803 VDD.n2802 2.48924
R11324 VDD.n2806 VDD.n2805 2.48924
R11325 VDD.n2809 VDD.n2808 2.48924
R11326 VDD.n2812 VDD.n2811 2.48924
R11327 VDD.n2815 VDD.n2814 2.48924
R11328 VDD.n2818 VDD.n2817 2.48924
R11329 VDD.n2821 VDD.n2820 2.48924
R11330 VDD.n2824 VDD.n2823 2.48924
R11331 VDD.n6323 VDD.n6322 2.48924
R11332 VDD.n6326 VDD.n6325 2.48924
R11333 VDD.n6443 VDD.n6442 2.48924
R11334 VDD.n3457 VDD.n3456 2.48924
R11335 VDD.n3460 VDD.n3459 2.48924
R11336 VDD.n3463 VDD.n3462 2.48924
R11337 VDD.n3466 VDD.n3465 2.48924
R11338 VDD.n3469 VDD.n3468 2.48924
R11339 VDD.n3472 VDD.n3471 2.48924
R11340 VDD.n3475 VDD.n3474 2.48924
R11341 VDD.n3478 VDD.n3477 2.48924
R11342 VDD.n3481 VDD.n3480 2.48924
R11343 VDD.n3484 VDD.n3483 2.48924
R11344 VDD.n3487 VDD.n3486 2.48924
R11345 VDD.n3490 VDD.n3489 2.48924
R11346 VDD.n3493 VDD.n3492 2.48924
R11347 VDD.n3496 VDD.n3495 2.48924
R11348 VDD.n3499 VDD.n3498 2.48924
R11349 VDD.n3502 VDD.n3501 2.48924
R11350 VDD.n3505 VDD.n3504 2.48924
R11351 VDD.n3508 VDD.n3507 2.48924
R11352 VDD.n3511 VDD.n3510 2.48924
R11353 VDD.n3514 VDD.n3513 2.48924
R11354 VDD.n3517 VDD.n3516 2.48924
R11355 VDD.n3520 VDD.n3519 2.48924
R11356 VDD.n3523 VDD.n3522 2.48924
R11357 VDD.n3526 VDD.n3525 2.48924
R11358 VDD.n3529 VDD.n3528 2.48924
R11359 VDD.n3532 VDD.n3531 2.48924
R11360 VDD.n3535 VDD.n3534 2.48924
R11361 VDD.n3538 VDD.n3537 2.48924
R11362 VDD.n3541 VDD.n3540 2.48924
R11363 VDD.n3544 VDD.n3543 2.48924
R11364 VDD.n3547 VDD.n3546 2.48924
R11365 VDD.n3550 VDD.n3549 2.48924
R11366 VDD.n3553 VDD.n3552 2.48924
R11367 VDD.n3556 VDD.n3555 2.48924
R11368 VDD.n3559 VDD.n3558 2.48924
R11369 VDD.n3562 VDD.n3561 2.48924
R11370 VDD.n3565 VDD.n3564 2.48924
R11371 VDD.n3568 VDD.n3567 2.48924
R11372 VDD.n3571 VDD.n3570 2.48924
R11373 VDD.n3574 VDD.n3573 2.48924
R11374 VDD.n3577 VDD.n3576 2.48924
R11375 VDD.n5403 VDD.n5402 2.48924
R11376 VDD.n3958 VDD.n3957 2.48924
R11377 VDD.n3961 VDD.n3960 2.48924
R11378 VDD.n3964 VDD.n3963 2.48924
R11379 VDD.n3967 VDD.n3966 2.48924
R11380 VDD.n3970 VDD.n3969 2.48924
R11381 VDD.n3973 VDD.n3972 2.48924
R11382 VDD.n3976 VDD.n3975 2.48924
R11383 VDD.n3979 VDD.n3978 2.48924
R11384 VDD.n3982 VDD.n3981 2.48924
R11385 VDD.n3985 VDD.n3984 2.48924
R11386 VDD.n3988 VDD.n3987 2.48924
R11387 VDD.n3991 VDD.n3990 2.48924
R11388 VDD.n3994 VDD.n3993 2.48924
R11389 VDD.n3997 VDD.n3996 2.48924
R11390 VDD.n4000 VDD.n3999 2.48924
R11391 VDD.n4003 VDD.n4002 2.48924
R11392 VDD.n4006 VDD.n4005 2.48924
R11393 VDD.n4009 VDD.n4008 2.48924
R11394 VDD.n4012 VDD.n4011 2.48924
R11395 VDD.n4015 VDD.n4014 2.48924
R11396 VDD.n4018 VDD.n4017 2.48924
R11397 VDD.n4021 VDD.n4020 2.48924
R11398 VDD.n4024 VDD.n4023 2.48924
R11399 VDD.n4027 VDD.n4026 2.48924
R11400 VDD.n4030 VDD.n4029 2.48924
R11401 VDD.n4033 VDD.n4032 2.48924
R11402 VDD.n4036 VDD.n4035 2.48924
R11403 VDD.n4039 VDD.n4038 2.48924
R11404 VDD.n4042 VDD.n4041 2.48924
R11405 VDD.n4045 VDD.n4044 2.48924
R11406 VDD.n4048 VDD.n4047 2.48924
R11407 VDD.n4051 VDD.n4050 2.48924
R11408 VDD.n4054 VDD.n4053 2.48924
R11409 VDD.n4057 VDD.n4056 2.48924
R11410 VDD.n4060 VDD.n4059 2.48924
R11411 VDD.n4063 VDD.n4062 2.48924
R11412 VDD.n4066 VDD.n4065 2.48924
R11413 VDD.n4069 VDD.n4068 2.48924
R11414 VDD.n4072 VDD.n4071 2.48924
R11415 VDD.n5555 VDD.n5554 2.48924
R11416 VDD.n5552 VDD.n5551 2.48924
R11417 VDD.n5549 VDD.n5548 2.48924
R11418 VDD.n5417 VDD.n5416 2.48924
R11419 VDD.n5946 VDD.n5945 2.48924
R11420 VDD.n5280 VDD.n5279 2.48924
R11421 VDD.n6752 VDD.n6751 2.48924
R11422 VDD.n6755 VDD.n6754 2.48924
R11423 VDD.n6758 VDD.n6757 2.48924
R11424 VDD.n6761 VDD.n6760 2.48924
R11425 VDD.n6764 VDD.n6763 2.48924
R11426 VDD.n6767 VDD.n6766 2.48924
R11427 VDD.n6770 VDD.n6769 2.48924
R11428 VDD.n6773 VDD.n6772 2.48924
R11429 VDD.n6776 VDD.n6775 2.48924
R11430 VDD.n6779 VDD.n6778 2.48924
R11431 VDD.n6782 VDD.n6781 2.48924
R11432 VDD.n6785 VDD.n6784 2.48924
R11433 VDD.n6788 VDD.n6787 2.48924
R11434 VDD.n6791 VDD.n6790 2.48924
R11435 VDD.n6794 VDD.n6793 2.48924
R11436 VDD.n6797 VDD.n6796 2.48924
R11437 VDD.n6800 VDD.n6799 2.48924
R11438 VDD.n6803 VDD.n6802 2.48924
R11439 VDD.n6806 VDD.n6805 2.48924
R11440 VDD.n6809 VDD.n6808 2.48924
R11441 VDD.n6812 VDD.n6811 2.48924
R11442 VDD.n6815 VDD.n6814 2.48924
R11443 VDD.n6818 VDD.n6817 2.48924
R11444 VDD.n6821 VDD.n6820 2.48924
R11445 VDD.n6824 VDD.n6823 2.48924
R11446 VDD.n6827 VDD.n6826 2.48924
R11447 VDD.n642 VDD.n641 2.48924
R11448 VDD.n645 VDD.n644 2.48924
R11449 VDD.n648 VDD.n647 2.48924
R11450 VDD.n651 VDD.n650 2.48924
R11451 VDD.n654 VDD.n653 2.48924
R11452 VDD.n657 VDD.n656 2.48924
R11453 VDD.n660 VDD.n659 2.48924
R11454 VDD.n663 VDD.n662 2.48924
R11455 VDD.n666 VDD.n665 2.48924
R11456 VDD.n669 VDD.n668 2.48924
R11457 VDD.n672 VDD.n671 2.48924
R11458 VDD.n675 VDD.n674 2.48924
R11459 VDD.n678 VDD.n677 2.48924
R11460 VDD.n681 VDD.n680 2.48924
R11461 VDD.n684 VDD.n683 2.48924
R11462 VDD.n687 VDD.n686 2.48924
R11463 VDD.n690 VDD.n689 2.48924
R11464 VDD.n693 VDD.n692 2.48924
R11465 VDD.n696 VDD.n695 2.48924
R11466 VDD.n699 VDD.n698 2.48924
R11467 VDD.n702 VDD.n701 2.48924
R11468 VDD.n705 VDD.n704 2.48924
R11469 VDD.n708 VDD.n707 2.48924
R11470 VDD.n6889 VDD.n6888 2.48924
R11471 VDD.n6892 VDD.n6891 2.48924
R11472 VDD.n6895 VDD.n6894 2.48924
R11473 VDD.n6898 VDD.n6897 2.48924
R11474 VDD.n6901 VDD.n6900 2.48924
R11475 VDD.n6904 VDD.n6903 2.48924
R11476 VDD.n6907 VDD.n6906 2.48924
R11477 VDD.n6910 VDD.n6909 2.48924
R11478 VDD.n6913 VDD.n6912 2.48924
R11479 VDD.n6916 VDD.n6915 2.48924
R11480 VDD.n6919 VDD.n6918 2.48924
R11481 VDD.n6922 VDD.n6921 2.48924
R11482 VDD.n6925 VDD.n6924 2.48924
R11483 VDD.n6928 VDD.n6927 2.48924
R11484 VDD.n6931 VDD.n6930 2.48924
R11485 VDD.n6934 VDD.n6933 2.48924
R11486 VDD.n6937 VDD.n6936 2.48924
R11487 VDD.n6940 VDD.n6939 2.48924
R11488 VDD.n6943 VDD.n6942 2.48924
R11489 VDD.n6946 VDD.n6945 2.48924
R11490 VDD.n6949 VDD.n6948 2.48924
R11491 VDD.n6952 VDD.n6951 2.48924
R11492 VDD.n6955 VDD.n6954 2.48924
R11493 VDD.n6958 VDD.n6957 2.48924
R11494 VDD.n6961 VDD.n6960 2.48924
R11495 VDD.n6964 VDD.n6963 2.48924
R11496 VDD.n132 VDD.n131 2.48924
R11497 VDD.n129 VDD.n128 2.48924
R11498 VDD.n126 VDD.n125 2.48924
R11499 VDD.n123 VDD.n122 2.48924
R11500 VDD.n120 VDD.n119 2.48924
R11501 VDD.n117 VDD.n116 2.48924
R11502 VDD.n114 VDD.n113 2.48924
R11503 VDD.n111 VDD.n110 2.48924
R11504 VDD.n108 VDD.n107 2.48924
R11505 VDD.n105 VDD.n104 2.48924
R11506 VDD.n102 VDD.n101 2.48924
R11507 VDD.n99 VDD.n98 2.48924
R11508 VDD.n96 VDD.n95 2.48924
R11509 VDD.n93 VDD.n92 2.48924
R11510 VDD.n90 VDD.n89 2.48924
R11511 VDD.n87 VDD.n86 2.48924
R11512 VDD.n84 VDD.n83 2.48924
R11513 VDD.n81 VDD.n80 2.48924
R11514 VDD.n78 VDD.n77 2.48924
R11515 VDD.n75 VDD.n74 2.48924
R11516 VDD.n72 VDD.n71 2.48924
R11517 VDD.n1783 VDD.n1782 2.48924
R11518 VDD.n1780 VDD.n1779 2.48924
R11519 VDD.n1777 VDD.n1776 2.48924
R11520 VDD.n1774 VDD.n1773 2.48924
R11521 VDD.n1771 VDD.n1770 2.48924
R11522 VDD.n1768 VDD.n1767 2.48924
R11523 VDD.n1765 VDD.n1764 2.48924
R11524 VDD.n1762 VDD.n1761 2.48924
R11525 VDD.n1759 VDD.n1758 2.48924
R11526 VDD.n1756 VDD.n1755 2.48924
R11527 VDD.n1753 VDD.n1752 2.48924
R11528 VDD.n1750 VDD.n1749 2.48924
R11529 VDD.n1747 VDD.n1746 2.48924
R11530 VDD.n1744 VDD.n1743 2.48924
R11531 VDD.n1741 VDD.n1740 2.48924
R11532 VDD.n1738 VDD.n1737 2.48924
R11533 VDD.n1735 VDD.n1734 2.48924
R11534 VDD.n1732 VDD.n1731 2.48924
R11535 VDD.n1729 VDD.n1728 2.48924
R11536 VDD.n1726 VDD.n1725 2.48924
R11537 VDD.n1723 VDD.n1722 2.48924
R11538 VDD.n1720 VDD.n1719 2.48924
R11539 VDD.n1717 VDD.n1716 2.48924
R11540 VDD.n1714 VDD.n1713 2.48924
R11541 VDD.n1711 VDD.n1710 2.48924
R11542 VDD.n1708 VDD.n1707 2.48924
R11543 VDD.n1705 VDD.n1704 2.48924
R11544 VDD.n1702 VDD.n1701 2.48924
R11545 VDD.n1699 VDD.n1698 2.48924
R11546 VDD.n1696 VDD.n1695 2.48924
R11547 VDD.n1693 VDD.n1692 2.48924
R11548 VDD.n1690 VDD.n1689 2.48924
R11549 VDD.n1687 VDD.n1686 2.48924
R11550 VDD.n1684 VDD.n1683 2.48924
R11551 VDD.n1681 VDD.n1680 2.48924
R11552 VDD.n1678 VDD.n1677 2.48924
R11553 VDD.n1675 VDD.n1674 2.48924
R11554 VDD.n1672 VDD.n1671 2.48924
R11555 VDD.n1921 VDD.n1920 2.48924
R11556 VDD.n1918 VDD.n1917 2.48924
R11557 VDD.n1915 VDD.n1914 2.48924
R11558 VDD.n1912 VDD.n1911 2.48924
R11559 VDD.n1909 VDD.n1908 2.48924
R11560 VDD.n1906 VDD.n1905 2.48924
R11561 VDD.n1903 VDD.n1902 2.48924
R11562 VDD.n1900 VDD.n1899 2.48924
R11563 VDD.n1897 VDD.n1896 2.48924
R11564 VDD.n1894 VDD.n1893 2.48924
R11565 VDD.n1891 VDD.n1890 2.48924
R11566 VDD.n1888 VDD.n1887 2.48924
R11567 VDD.n1885 VDD.n1884 2.48924
R11568 VDD.n1882 VDD.n1881 2.48924
R11569 VDD.n1879 VDD.n1878 2.48924
R11570 VDD.n1876 VDD.n1875 2.48924
R11571 VDD.n1873 VDD.n1872 2.48924
R11572 VDD.n1870 VDD.n1869 2.48924
R11573 VDD.n1867 VDD.n1866 2.48924
R11574 VDD.n1864 VDD.n1863 2.48924
R11575 VDD.n1861 VDD.n1860 2.48924
R11576 VDD.n1858 VDD.n1857 2.48924
R11577 VDD.n1855 VDD.n1854 2.48924
R11578 VDD.n1852 VDD.n1851 2.48924
R11579 VDD.n1849 VDD.n1848 2.48924
R11580 VDD.n1846 VDD.n1845 2.48924
R11581 VDD.n1843 VDD.n1842 2.48924
R11582 VDD.n1840 VDD.n1839 2.48924
R11583 VDD.n1837 VDD.n1836 2.48924
R11584 VDD.n1834 VDD.n1833 2.48924
R11585 VDD.n1831 VDD.n1830 2.48924
R11586 VDD.n1828 VDD.n1827 2.48924
R11587 VDD.n1825 VDD.n1824 2.48924
R11588 VDD.n1822 VDD.n1821 2.48924
R11589 VDD.n1819 VDD.n1818 2.48924
R11590 VDD.n1816 VDD.n1815 2.48924
R11591 VDD.n1813 VDD.n1812 2.48924
R11592 VDD.n1810 VDD.n1809 2.48924
R11593 VDD.n7454 VDD.t44 2.48574
R11594 VDD.n8340 VDD.t9 2.4382
R11595 VDD.n822 VDD.t577 2.42448
R11596 VDD.n855 VDD.t579 2.42448
R11597 VDD.t433 VDD.t1 2.31934
R11598 VDD.t587 VDD.t439 2.31934
R11599 VDD.t507 VDD.t38 2.31934
R11600 VDD.t536 VDD.t862 2.31934
R11601 VDD.t171 VDD.t153 2.31934
R11602 VDD.n2259 VDD.t48 2.2583
R11603 VDD.n2363 VDD.t271 2.2583
R11604 VDD.n2494 VDD.t179 2.2583
R11605 VDD.n18 VDD.n17 2.21137
R11606 VDD.n17 VDD.n16 2.21137
R11607 VDD.n304 VDD.n303 2.21137
R11608 VDD.n21 VDD.n20 2.21137
R11609 VDD.n20 VDD.n19 2.21137
R11610 VDD.n310 VDD.n309 2.21137
R11611 VDD.n24 VDD.n23 2.21137
R11612 VDD.n23 VDD.n22 2.21137
R11613 VDD.n6859 VDD.n6858 2.21137
R11614 VDD.n27 VDD.n26 2.21137
R11615 VDD.n26 VDD.n25 2.21137
R11616 VDD.n6865 VDD.n6864 2.21137
R11617 VDD.n5621 VDD.n5620 2.07441
R11618 VDD.n4237 VDD.n4234 2.07441
R11619 VDD.n5615 VDD.n5614 2.07441
R11620 VDD.n4231 VDD.n4228 2.07441
R11621 VDD.n5609 VDD.n5608 2.07441
R11622 VDD.n4225 VDD.n4222 2.07441
R11623 VDD.n5591 VDD.n5590 2.07441
R11624 VDD.n4197 VDD.n4194 2.07441
R11625 VDD.n5585 VDD.n5584 2.07441
R11626 VDD.n4191 VDD.n4188 2.07441
R11627 VDD.n5537 VDD.n5536 2.07441
R11628 VDD.n3945 VDD.n3942 2.07441
R11629 VDD.n5531 VDD.n5530 2.07441
R11630 VDD.n3939 VDD.n3936 2.07441
R11631 VDD.n5513 VDD.n5512 2.07441
R11632 VDD.n3911 VDD.n3908 2.07441
R11633 VDD.n5507 VDD.n5506 2.07441
R11634 VDD.n3905 VDD.n3902 2.07441
R11635 VDD.n5501 VDD.n5500 2.07441
R11636 VDD.n3899 VDD.n3896 2.07441
R11637 VDD.n5355 VDD.n5354 2.07441
R11638 VDD.n3399 VDD.n3396 2.07441
R11639 VDD.n5361 VDD.n5360 2.07441
R11640 VDD.n3405 VDD.n3402 2.07441
R11641 VDD.n5367 VDD.n5366 2.07441
R11642 VDD.n3411 VDD.n3408 2.07441
R11643 VDD.n5385 VDD.n5384 2.07441
R11644 VDD.n3439 VDD.n3436 2.07441
R11645 VDD.n5391 VDD.n5390 2.07441
R11646 VDD.n3445 VDD.n3442 2.07441
R11647 VDD.n5432 VDD.n5431 2.07441
R11648 VDD.n3713 VDD.n3710 2.07441
R11649 VDD.n5438 VDD.n5437 2.07441
R11650 VDD.n3719 VDD.n3716 2.07441
R11651 VDD.n5456 VDD.n5455 2.07441
R11652 VDD.n3747 VDD.n3744 2.07441
R11653 VDD.n5462 VDD.n5461 2.07441
R11654 VDD.n3753 VDD.n3750 2.07441
R11655 VDD.n5468 VDD.n5467 2.07441
R11656 VDD.n3759 VDD.n3756 2.07441
R11657 VDD.n6205 VDD.n6204 2.07441
R11658 VDD.n2910 VDD.n2907 2.07441
R11659 VDD.n6199 VDD.n6198 2.07441
R11660 VDD.n2916 VDD.n2913 2.07441
R11661 VDD.n6193 VDD.n6192 2.07441
R11662 VDD.n2922 VDD.n2919 2.07441
R11663 VDD.n6175 VDD.n6174 2.07441
R11664 VDD.n2950 VDD.n2947 2.07441
R11665 VDD.n6169 VDD.n6168 2.07441
R11666 VDD.n2956 VDD.n2953 2.07441
R11667 VDD.n5295 VDD.n5294 2.07441
R11668 VDD.n3209 VDD.n3206 2.07441
R11669 VDD.n5301 VDD.n5300 2.07441
R11670 VDD.n3215 VDD.n3212 2.07441
R11671 VDD.n5319 VDD.n5318 2.07441
R11672 VDD.n3243 VDD.n3240 2.07441
R11673 VDD.n5325 VDD.n5324 2.07441
R11674 VDD.n3249 VDD.n3246 2.07441
R11675 VDD.n5331 VDD.n5330 2.07441
R11676 VDD.n3255 VDD.n3252 2.07441
R11677 VDD.n2542 VDD.n2541 2.07441
R11678 VDD.n2842 VDD.n2839 2.07441
R11679 VDD.n2548 VDD.n2547 2.07441
R11680 VDD.n2848 VDD.n2845 2.07441
R11681 VDD.n2566 VDD.n2565 2.07441
R11682 VDD.n2876 VDD.n2873 2.07441
R11683 VDD.n2572 VDD.n2571 2.07441
R11684 VDD.n2882 VDD.n2879 2.07441
R11685 VDD.n2578 VDD.n2577 2.07441
R11686 VDD.n2888 VDD.n2885 2.07441
R11687 VDD.n6624 VDD.n6623 2.02746
R11688 VDD.n546 VDD.n545 2.02746
R11689 VDD.n552 VDD.n551 2.02746
R11690 VDD.n560 VDD.n559 2.02746
R11691 VDD.n559 VDD.n558 2.02746
R11692 VDD.n564 VDD.n563 2.02746
R11693 VDD.n563 VDD.n562 2.02746
R11694 VDD.n743 VDD.n740 2.02746
R11695 VDD.n746 VDD.n743 2.02746
R11696 VDD.n752 VDD.n749 2.02746
R11697 VDD.n755 VDD.n752 2.02746
R11698 VDD.n1052 VDD.n1049 2.02746
R11699 VDD.n1055 VDD.n1052 2.02746
R11700 VDD.n1043 VDD.n1040 2.02746
R11701 VDD.n1046 VDD.n1043 2.02746
R11702 VDD.n1035 VDD.n1034 2.02746
R11703 VDD.n1031 VDD.n1030 2.02746
R11704 VDD.n6630 VDD.n6629 2.02746
R11705 VDD.n2479 VDD.n1364 1.9805
R11706 VDD.n2469 VDD.n1375 1.9805
R11707 VDD.n2455 VDD.n1386 1.9805
R11708 VDD.n2444 VDD.n1397 1.9805
R11709 VDD.n2434 VDD.n1408 1.9805
R11710 VDD.n2420 VDD.n1419 1.9805
R11711 VDD.n2385 VDD.n1438 1.9805
R11712 VDD.n2362 VDD.n1453 1.9805
R11713 VDD.n2366 VDD.n1450 1.9805
R11714 VDD.n1144 VDD.n1131 1.9805
R11715 VDD.n1147 VDD.n1128 1.9805
R11716 VDD.n2374 VDD.n1445 1.9805
R11717 VDD.n2381 VDD.n1442 1.9805
R11718 VDD.n2396 VDD.n1431 1.9805
R11719 VDD.n1165 VDD.n1119 1.9805
R11720 VDD.n2410 VDD.n1425 1.9805
R11721 VDD.n1174 VDD.n1113 1.9805
R11722 VDD.n2493 VDD.n1353 1.9805
R11723 VDD.n2497 VDD.n1348 1.9805
R11724 VDD.n1223 VDD.n1107 1.9805
R11725 VDD.n1226 VDD.n1102 1.9805
R11726 VDD.n6848 VDD.n6829 1.90688
R11727 VDD.n6848 VDD.n6830 1.90688
R11728 VDD.n6848 VDD.n6831 1.90688
R11729 VDD.n6848 VDD.n6832 1.90688
R11730 VDD.n6848 VDD.n6833 1.90688
R11731 VDD.n6848 VDD.n6834 1.90688
R11732 VDD.n6848 VDD.n6835 1.90688
R11733 VDD.n6848 VDD.n6836 1.90688
R11734 VDD.n6848 VDD.n6837 1.90688
R11735 VDD.n6848 VDD.n6838 1.90688
R11736 VDD.n6848 VDD.n6839 1.90688
R11737 VDD.n6848 VDD.n6840 1.90688
R11738 VDD.n6848 VDD.n6841 1.90688
R11739 VDD.n6848 VDD.n6842 1.90688
R11740 VDD.n6848 VDD.n6843 1.90688
R11741 VDD.n6848 VDD.n6844 1.90688
R11742 VDD.n6848 VDD.n6845 1.90688
R11743 VDD.n6848 VDD.n6846 1.90688
R11744 VDD.n734 VDD.n715 1.90688
R11745 VDD.n734 VDD.n716 1.90688
R11746 VDD.n734 VDD.n717 1.90688
R11747 VDD.n734 VDD.n718 1.90688
R11748 VDD.n734 VDD.n719 1.90688
R11749 VDD.n734 VDD.n720 1.90688
R11750 VDD.n734 VDD.n721 1.90688
R11751 VDD.n734 VDD.n722 1.90688
R11752 VDD.n734 VDD.n723 1.90688
R11753 VDD.n734 VDD.n724 1.90688
R11754 VDD.n734 VDD.n725 1.90688
R11755 VDD.n734 VDD.n726 1.90688
R11756 VDD.n734 VDD.n727 1.90688
R11757 VDD.n734 VDD.n728 1.90688
R11758 VDD.n734 VDD.n729 1.90688
R11759 VDD.n734 VDD.n730 1.90688
R11760 VDD.n734 VDD.n731 1.90688
R11761 VDD.n40 VDD.n29 1.90688
R11762 VDD.n40 VDD.n30 1.90688
R11763 VDD.n40 VDD.n31 1.90688
R11764 VDD.n40 VDD.n32 1.90688
R11765 VDD.n40 VDD.n33 1.90688
R11766 VDD.n40 VDD.n34 1.90688
R11767 VDD.n40 VDD.n35 1.90688
R11768 VDD.n40 VDD.n36 1.90688
R11769 VDD.n40 VDD.n37 1.90688
R11770 VDD.n40 VDD.n38 1.90688
R11771 VDD.n40 VDD.n39 1.90688
R11772 VDD.n6976 VDD.n6966 1.90688
R11773 VDD.n6976 VDD.n6967 1.90688
R11774 VDD.n6976 VDD.n6968 1.90688
R11775 VDD.n6976 VDD.n6969 1.90688
R11776 VDD.n6976 VDD.n6970 1.90688
R11777 VDD.n6976 VDD.n6971 1.90688
R11778 VDD.n6976 VDD.n6972 1.90688
R11779 VDD.n6976 VDD.n6973 1.90688
R11780 VDD.n6976 VDD.n6974 1.90688
R11781 VDD.n2339 VDD.n2337 1.90688
R11782 VDD.n2339 VDD.n2338 1.90688
R11783 VDD.n2148 VDD.n2146 1.90688
R11784 VDD.n2148 VDD.n2147 1.90688
R11785 VDD.n1152 VDD.n1123 1.88267
R11786 VDD.n7431 VDD.t55 1.86443
R11787 VDD.n7510 VDD.t90 1.86443
R11788 VDD.n2250 VDD.t53 1.84779
R11789 VDD.n5638 VDD.n5637 1.7854
R11790 VDD.n5633 VDD.n5632 1.7854
R11791 VDD.n3585 VDD.n3584 1.7854
R11792 VDD.n4080 VDD.n4079 1.7854
R11793 VDD.n6312 VDD.n6309 1.7854
R11794 VDD.n736 VDD.n735 1.7854
R11795 VDD.n8282 VDD.n8281 1.7854
R11796 VDD.n8277 VDD.n8276 1.7854
R11797 VDD.n8272 VDD.n8271 1.7854
R11798 VDD.n8267 VDD.n8266 1.7854
R11799 VDD.n8262 VDD.n8261 1.7854
R11800 VDD.n8257 VDD.n8256 1.7854
R11801 VDD.n8249 VDD.n8248 1.7854
R11802 VDD.n529 VDD.n528 1.7854
R11803 VDD.n524 VDD.n523 1.7854
R11804 VDD.n519 VDD.n518 1.7854
R11805 VDD.n514 VDD.n513 1.7854
R11806 VDD.n509 VDD.n508 1.7854
R11807 VDD.n504 VDD.n503 1.7854
R11808 VDD.n499 VDD.n498 1.7854
R11809 VDD.n494 VDD.n493 1.7854
R11810 VDD.n489 VDD.n488 1.7854
R11811 VDD.n484 VDD.n483 1.7854
R11812 VDD.n479 VDD.n478 1.7854
R11813 VDD.n2028 VDD.n2027 1.7854
R11814 VDD.n2023 VDD.n2022 1.7854
R11815 VDD.n2018 VDD.n2017 1.7854
R11816 VDD.n2013 VDD.n2012 1.7854
R11817 VDD.n2008 VDD.n2007 1.7854
R11818 VDD.n2003 VDD.n2002 1.7854
R11819 VDD.n1998 VDD.n1997 1.7854
R11820 VDD.n1993 VDD.n1992 1.7854
R11821 VDD.n1988 VDD.n1987 1.7854
R11822 VDD.n1983 VDD.n1982 1.7854
R11823 VDD.n4246 VDD.n4245 1.78487
R11824 VDD.n4251 VDD.n4250 1.78487
R11825 VDD.n4256 VDD.n4255 1.78487
R11826 VDD.n4261 VDD.n4260 1.78487
R11827 VDD.n4266 VDD.n4265 1.78487
R11828 VDD.n4271 VDD.n4270 1.78487
R11829 VDD.n4276 VDD.n4275 1.78487
R11830 VDD.n4281 VDD.n4280 1.78487
R11831 VDD.n4286 VDD.n4285 1.78487
R11832 VDD.n4291 VDD.n4290 1.78487
R11833 VDD.n4296 VDD.n4295 1.78487
R11834 VDD.n4301 VDD.n4300 1.78487
R11835 VDD.n4306 VDD.n4305 1.78487
R11836 VDD.n4311 VDD.n4310 1.78487
R11837 VDD.n4316 VDD.n4315 1.78487
R11838 VDD.n4321 VDD.n4320 1.78487
R11839 VDD.n4326 VDD.n4325 1.78487
R11840 VDD.n4331 VDD.n4330 1.78487
R11841 VDD.n4336 VDD.n4335 1.78487
R11842 VDD.n4341 VDD.n4340 1.78487
R11843 VDD.n3690 VDD.n3689 1.78487
R11844 VDD.n3685 VDD.n3684 1.78487
R11845 VDD.n3680 VDD.n3679 1.78487
R11846 VDD.n3675 VDD.n3674 1.78487
R11847 VDD.n3670 VDD.n3669 1.78487
R11848 VDD.n3665 VDD.n3664 1.78487
R11849 VDD.n3660 VDD.n3659 1.78487
R11850 VDD.n3655 VDD.n3654 1.78487
R11851 VDD.n3650 VDD.n3649 1.78487
R11852 VDD.n3645 VDD.n3644 1.78487
R11853 VDD.n3640 VDD.n3639 1.78487
R11854 VDD.n3635 VDD.n3634 1.78487
R11855 VDD.n3630 VDD.n3629 1.78487
R11856 VDD.n3625 VDD.n3624 1.78487
R11857 VDD.n3620 VDD.n3619 1.78487
R11858 VDD.n3615 VDD.n3614 1.78487
R11859 VDD.n3610 VDD.n3609 1.78487
R11860 VDD.n3605 VDD.n3604 1.78487
R11861 VDD.n3600 VDD.n3599 1.78487
R11862 VDD.n3595 VDD.n3594 1.78487
R11863 VDD.n3590 VDD.n3589 1.78487
R11864 VDD.n3186 VDD.n3185 1.78487
R11865 VDD.n3181 VDD.n3180 1.78487
R11866 VDD.n3176 VDD.n3175 1.78487
R11867 VDD.n3171 VDD.n3170 1.78487
R11868 VDD.n3166 VDD.n3165 1.78487
R11869 VDD.n3161 VDD.n3160 1.78487
R11870 VDD.n3156 VDD.n3155 1.78487
R11871 VDD.n3151 VDD.n3150 1.78487
R11872 VDD.n3146 VDD.n3145 1.78487
R11873 VDD.n3141 VDD.n3140 1.78487
R11874 VDD.n3136 VDD.n3135 1.78487
R11875 VDD.n3131 VDD.n3130 1.78487
R11876 VDD.n3126 VDD.n3125 1.78487
R11877 VDD.n3121 VDD.n3120 1.78487
R11878 VDD.n3116 VDD.n3115 1.78487
R11879 VDD.n3111 VDD.n3110 1.78487
R11880 VDD.n3106 VDD.n3105 1.78487
R11881 VDD.n3101 VDD.n3100 1.78487
R11882 VDD.n3096 VDD.n3095 1.78487
R11883 VDD.n3091 VDD.n3090 1.78487
R11884 VDD.n3086 VDD.n3085 1.78487
R11885 VDD.n6312 VDD.n6311 1.78487
R11886 VDD.n6435 VDD.n6434 1.78487
R11887 VDD.n6429 VDD.n6428 1.78487
R11888 VDD.n6424 VDD.n6423 1.78487
R11889 VDD.n6419 VDD.n6418 1.78487
R11890 VDD.n6414 VDD.n6413 1.78487
R11891 VDD.n6409 VDD.n6408 1.78487
R11892 VDD.n6404 VDD.n6403 1.78487
R11893 VDD.n6399 VDD.n6398 1.78487
R11894 VDD.n6394 VDD.n6393 1.78487
R11895 VDD.n6389 VDD.n6388 1.78487
R11896 VDD.n6384 VDD.n6383 1.78487
R11897 VDD.n6379 VDD.n6378 1.78487
R11898 VDD.n6374 VDD.n6373 1.78487
R11899 VDD.n6369 VDD.n6368 1.78487
R11900 VDD.n6364 VDD.n6363 1.78487
R11901 VDD.n6359 VDD.n6358 1.78487
R11902 VDD.n6354 VDD.n6353 1.78487
R11903 VDD.n6349 VDD.n6348 1.78487
R11904 VDD.n6344 VDD.n6343 1.78487
R11905 VDD.n6339 VDD.n6338 1.78487
R11906 VDD.n6334 VDD.n6333 1.78487
R11907 VDD.n4174 VDD.n4173 1.78473
R11908 VDD.n4169 VDD.n4168 1.78473
R11909 VDD.n4164 VDD.n4163 1.78473
R11910 VDD.n4159 VDD.n4158 1.78473
R11911 VDD.n4154 VDD.n4153 1.78473
R11912 VDD.n4149 VDD.n4148 1.78473
R11913 VDD.n4144 VDD.n4143 1.78473
R11914 VDD.n4139 VDD.n4138 1.78473
R11915 VDD.n4134 VDD.n4133 1.78473
R11916 VDD.n3384 VDD.n3383 1.78473
R11917 VDD.n3379 VDD.n3378 1.78473
R11918 VDD.n3374 VDD.n3373 1.78473
R11919 VDD.n3369 VDD.n3368 1.78473
R11920 VDD.n3364 VDD.n3363 1.78473
R11921 VDD.n3359 VDD.n3358 1.78473
R11922 VDD.n3354 VDD.n3353 1.78473
R11923 VDD.n3349 VDD.n3348 1.78473
R11924 VDD.n3344 VDD.n3343 1.78473
R11925 VDD.n3339 VDD.n3338 1.78473
R11926 VDD.n3334 VDD.n3333 1.78473
R11927 VDD.n3329 VDD.n3328 1.78473
R11928 VDD.n3324 VDD.n3323 1.78473
R11929 VDD.n3319 VDD.n3318 1.78473
R11930 VDD.n3314 VDD.n3313 1.78473
R11931 VDD.n3309 VDD.n3308 1.78473
R11932 VDD.n3304 VDD.n3303 1.78473
R11933 VDD.n3299 VDD.n3298 1.78473
R11934 VDD.n3294 VDD.n3293 1.78473
R11935 VDD.n3289 VDD.n3288 1.78473
R11936 VDD.n3284 VDD.n3283 1.78473
R11937 VDD.n3279 VDD.n3278 1.78473
R11938 VDD.n3274 VDD.n3273 1.78473
R11939 VDD.n3269 VDD.n3268 1.78473
R11940 VDD.n5344 VDD.n5341 1.78473
R11941 VDD.n5344 VDD.n5343 1.78473
R11942 VDD.n3884 VDD.n3883 1.78473
R11943 VDD.n3879 VDD.n3878 1.78473
R11944 VDD.n3874 VDD.n3873 1.78473
R11945 VDD.n3869 VDD.n3868 1.78473
R11946 VDD.n3864 VDD.n3863 1.78473
R11947 VDD.n3859 VDD.n3858 1.78473
R11948 VDD.n3854 VDD.n3853 1.78473
R11949 VDD.n3849 VDD.n3848 1.78473
R11950 VDD.n3844 VDD.n3843 1.78473
R11951 VDD.n3839 VDD.n3838 1.78473
R11952 VDD.n3834 VDD.n3833 1.78473
R11953 VDD.n3829 VDD.n3828 1.78473
R11954 VDD.n3824 VDD.n3823 1.78473
R11955 VDD.n3819 VDD.n3818 1.78473
R11956 VDD.n3814 VDD.n3813 1.78473
R11957 VDD.n3809 VDD.n3808 1.78473
R11958 VDD.n3804 VDD.n3803 1.78473
R11959 VDD.n3799 VDD.n3798 1.78473
R11960 VDD.n3794 VDD.n3793 1.78473
R11961 VDD.n3789 VDD.n3788 1.78473
R11962 VDD.n3784 VDD.n3783 1.78473
R11963 VDD.n3779 VDD.n3778 1.78473
R11964 VDD.n3774 VDD.n3773 1.78473
R11965 VDD.n3769 VDD.n3768 1.78473
R11966 VDD.n5481 VDD.n5478 1.78473
R11967 VDD.n5481 VDD.n5480 1.78473
R11968 VDD.n2966 VDD.n2965 1.78473
R11969 VDD.n2971 VDD.n2970 1.78473
R11970 VDD.n2976 VDD.n2975 1.78473
R11971 VDD.n2981 VDD.n2980 1.78473
R11972 VDD.n2986 VDD.n2985 1.78473
R11973 VDD.n2991 VDD.n2990 1.78473
R11974 VDD.n2996 VDD.n2995 1.78473
R11975 VDD.n3001 VDD.n3000 1.78473
R11976 VDD.n3006 VDD.n3005 1.78473
R11977 VDD.n3011 VDD.n3010 1.78473
R11978 VDD.n3016 VDD.n3015 1.78473
R11979 VDD.n3021 VDD.n3020 1.78473
R11980 VDD.n3026 VDD.n3025 1.78473
R11981 VDD.n3031 VDD.n3030 1.78473
R11982 VDD.n3036 VDD.n3035 1.78473
R11983 VDD.n3041 VDD.n3040 1.78473
R11984 VDD.n3046 VDD.n3045 1.78473
R11985 VDD.n3051 VDD.n3050 1.78473
R11986 VDD.n3056 VDD.n3055 1.78473
R11987 VDD.n3061 VDD.n3060 1.78473
R11988 VDD.n3066 VDD.n3065 1.78473
R11989 VDD.n3071 VDD.n3070 1.78473
R11990 VDD.n3076 VDD.n3075 1.78473
R11991 VDD.n970 VDD.n969 1.78473
R11992 VDD.n975 VDD.n974 1.78473
R11993 VDD.n980 VDD.n979 1.78473
R11994 VDD.n985 VDD.n984 1.78473
R11995 VDD.n990 VDD.n989 1.78473
R11996 VDD.n995 VDD.n994 1.78473
R11997 VDD.n1000 VDD.n999 1.78473
R11998 VDD.n1005 VDD.n1004 1.78473
R11999 VDD.n7162 VDD.n7161 1.78473
R12000 VDD.n7157 VDD.n7156 1.78473
R12001 VDD.n7152 VDD.n7151 1.78473
R12002 VDD.n7147 VDD.n7146 1.78473
R12003 VDD.n7142 VDD.n7141 1.78473
R12004 VDD.n7137 VDD.n7136 1.78473
R12005 VDD.n7132 VDD.n7131 1.78473
R12006 VDD.n7127 VDD.n7126 1.78473
R12007 VDD.n247 VDD.n246 1.78473
R12008 VDD.n252 VDD.n251 1.78473
R12009 VDD.n257 VDD.n256 1.78473
R12010 VDD.n262 VDD.n261 1.78473
R12011 VDD.n267 VDD.n266 1.78473
R12012 VDD.n272 VDD.n271 1.78473
R12013 VDD.n277 VDD.n276 1.78473
R12014 VDD.n282 VDD.n281 1.78473
R12015 VDD.n287 VDD.n286 1.78473
R12016 VDD.n301 VDD.n300 1.78473
R12017 VDD.n8056 VDD.n8055 1.78473
R12018 VDD.n8061 VDD.n8060 1.78473
R12019 VDD.n8066 VDD.n8065 1.78473
R12020 VDD.n8071 VDD.n8070 1.78473
R12021 VDD.n8076 VDD.n8075 1.78473
R12022 VDD.n8081 VDD.n8080 1.78473
R12023 VDD.n8086 VDD.n8085 1.78473
R12024 VDD.n8091 VDD.n8090 1.78473
R12025 VDD.n8096 VDD.n8095 1.78473
R12026 VDD.n8101 VDD.n8100 1.78473
R12027 VDD.n8106 VDD.n8105 1.78473
R12028 VDD.n1296 VDD.n1295 1.78473
R12029 VDD.n1301 VDD.n1300 1.78473
R12030 VDD.n1306 VDD.n1305 1.78473
R12031 VDD.n1311 VDD.n1310 1.78473
R12032 VDD.n1316 VDD.n1315 1.78473
R12033 VDD.n1321 VDD.n1320 1.78473
R12034 VDD.n1326 VDD.n1325 1.78473
R12035 VDD.n1331 VDD.n1330 1.78473
R12036 VDD.n1336 VDD.n1335 1.78473
R12037 VDD.n1341 VDD.n1340 1.78473
R12038 VDD.n393 VDD.n392 1.78093
R12039 VDD.n408 VDD.n405 1.78093
R12040 VDD.n7631 VDD.n7630 1.73593
R12041 VDD.n7625 VDD.n7624 1.73593
R12042 VDD.n7620 VDD.n7619 1.73593
R12043 VDD.n7615 VDD.n7614 1.73593
R12044 VDD.n7609 VDD.n7608 1.73593
R12045 VDD.n7866 VDD.n7864 1.73593
R12046 VDD.n7869 VDD.n7867 1.73593
R12047 VDD.n7872 VDD.n7870 1.73593
R12048 VDD.n7863 VDD.n7862 1.73541
R12049 VDD.n7866 VDD.n7865 1.73541
R12050 VDD.n7869 VDD.n7868 1.73541
R12051 VDD.n7872 VDD.n7871 1.73541
R12052 VDD.n7691 VDD.n7690 1.73527
R12053 VDD.n7685 VDD.n7684 1.73527
R12054 VDD.n7680 VDD.n7679 1.73527
R12055 VDD.n7675 VDD.n7674 1.73527
R12056 VDD.n7669 VDD.n7668 1.73527
R12057 VDD.n7832 VDD.n7831 1.73527
R12058 VDD.n7837 VDD.n7836 1.73527
R12059 VDD.n7843 VDD.n7842 1.73527
R12060 VDD.n7848 VDD.n7847 1.73527
R12061 VDD.n7240 VDD.n7239 1.73527
R12062 VDD.n7247 VDD.n7246 1.73527
R12063 VDD.n7253 VDD.n7252 1.73527
R12064 VDD.n7259 VDD.n7258 1.73527
R12065 VDD.n6611 VDD.n6610 1.61319
R12066 VDD.n7968 VDD.n7967 1.54224
R12067 VDD.n7974 VDD.n7973 1.52463
R12068 VDD.n7978 VDD.n7977 1.52463
R12069 VDD.n8162 VDD.n8159 1.49137
R12070 VDD.n8165 VDD.n8162 1.49137
R12071 VDD.n8151 VDD.n8148 1.49137
R12072 VDD.n8154 VDD.n8151 1.49137
R12073 VDD.n7900 VDD.n7897 1.49137
R12074 VDD.n7903 VDD.n7900 1.49137
R12075 VDD.n7232 VDD.n7231 1.49137
R12076 VDD.n7231 VDD.n7230 1.49137
R12077 VDD.n11 VDD.n10 1.49137
R12078 VDD.n10 VDD.n9 1.49137
R12079 VDD.n15 VDD.n14 1.49137
R12080 VDD.n14 VDD.n13 1.49137
R12081 VDD.n8323 VDD.n8322 1.49137
R12082 VDD.n8322 VDD.n8321 1.49137
R12083 VDD.n5406 VDD.n5405 1.467
R12084 VDD.n5558 VDD.n5557 1.467
R12085 VDD.n135 VDD.n134 1.467
R12086 VDD.n1786 VDD.n1785 1.467
R12087 VDD.n1924 VDD.n1923 1.467
R12088 VDD.n4344 VDD.n4343 1.46684
R12089 VDD.n4349 VDD.n4348 1.46684
R12090 VDD.n2827 VDD.n2826 1.46684
R12091 VDD.n6329 VDD.n6328 1.46684
R12092 VDD.n6438 VDD.n6437 1.46684
R12093 VDD.n6446 VDD.n6445 1.46684
R12094 VDD.n5409 VDD.n5408 1.46684
R12095 VDD.n3580 VDD.n3579 1.46684
R12096 VDD.n4075 VDD.n4074 1.46684
R12097 VDD.n5412 VDD.n5411 1.46684
R12098 VDD.n3693 VDD.n3692 1.46684
R12099 VDD.n3698 VDD.n3697 1.46684
R12100 VDD.n3081 VDD.n3080 1.46684
R12101 VDD.n3189 VDD.n3188 1.46684
R12102 VDD.n3194 VDD.n3193 1.46684
R12103 VDD.n6451 VDD.n6450 1.46684
R12104 VDD.n6454 VDD.n6453 1.46684
R12105 VDD.n6850 VDD.n6849 1.46684
R12106 VDD.n711 VDD.n710 1.46684
R12107 VDD.n6978 VDD.n6977 1.46684
R12108 VDD.n1801 VDD.n1800 1.46684
R12109 VDD.n1663 VDD.n1662 1.46684
R12110 VDD.n7938 VDD.t563 1.44978
R12111 VDD.n7875 VDD.n7873 1.44895
R12112 VDD.n7875 VDD.n7874 1.44847
R12113 VDD.n7822 VDD.n7821 1.4483
R12114 VDD.n1364 VDD.n1363 1.4405
R12115 VDD.n1363 VDD.n1362 1.4405
R12116 VDD.n1375 VDD.n1374 1.4405
R12117 VDD.n1374 VDD.n1373 1.4405
R12118 VDD.n1386 VDD.n1385 1.4405
R12119 VDD.n1385 VDD.n1384 1.4405
R12120 VDD.n1397 VDD.n1396 1.4405
R12121 VDD.n1396 VDD.n1395 1.4405
R12122 VDD.n1408 VDD.n1407 1.4405
R12123 VDD.n1407 VDD.n1406 1.4405
R12124 VDD.n1419 VDD.n1418 1.4405
R12125 VDD.n1418 VDD.n1417 1.4405
R12126 VDD.n1438 VDD.n1437 1.4405
R12127 VDD.n1437 VDD.n1436 1.4405
R12128 VDD.n1123 VDD.n1121 1.4405
R12129 VDD.n1431 VDD.n1430 1.4405
R12130 VDD.n1119 VDD.n1116 1.4405
R12131 VDD.n1425 VDD.n1424 1.4405
R12132 VDD.n1113 VDD.n1110 1.4405
R12133 VDD.n166 VDD.t467 1.43811
R12134 VDD.n181 VDD.t500 1.43811
R12135 VDD.n2470 VDD.t97 1.43728
R12136 VDD.n7634 VDD.n7633 1.41705
R12137 VDD.n4518 VDD.n4501 1.40703
R12138 VDD.n4820 VDD.n4818 1.40703
R12139 VDD.n5122 VDD.n5121 1.40703
R12140 VDD.n6154 VDD.n6152 1.40703
R12141 VDD.n42 VDD.n41 1.40703
R12142 VDD.n454 VDD.n453 1.40703
R12143 VDD.n1241 VDD.n1239 1.40703
R12144 VDD.n1655 VDD.n1653 1.40703
R12145 VDD.n1527 VDD.n1525 1.40703
R12146 VDD.n2341 VDD.n2335 1.40703
R12147 VDD.n2150 VDD.n2144 1.40703
R12148 VDD.n2047 VDD.n2032 1.40703
R12149 VDD.n2532 VDD.n2517 1.40703
R12150 VDD.n4354 VDD.n4351 1.40703
R12151 VDD.n4524 VDD.n4521 1.40703
R12152 VDD.n5644 VDD.n5642 1.40703
R12153 VDD.n5745 VDD.n5743 1.40703
R12154 VDD.n4820 VDD.n4819 1.40656
R12155 VDD.n6150 VDD.n6148 1.40656
R12156 VDD.n2684 VDD.n2682 1.40656
R12157 VDD.n8296 VDD.n8295 1.40656
R12158 VDD.n540 VDD.n539 1.40656
R12159 VDD.n1527 VDD.n1526 1.40656
R12160 VDD.n1655 VDD.n1654 1.40656
R12161 VDD.n1459 VDD.n1458 1.40656
R12162 VDD.n4524 VDD.n4523 1.40656
R12163 VDD.n4354 VDD.n4353 1.40656
R12164 VDD.n5749 VDD.n5747 1.40656
R12165 VDD.n6598 VDD.n6597 1.40638
R12166 VDD.n5343 VDD.n5342 1.40638
R12167 VDD.n4974 VDD.n4973 1.40638
R12168 VDD.n4826 VDD.n4825 1.40638
R12169 VDD.n5480 VDD.n5479 1.40638
R12170 VDD.n4672 VDD.n4671 1.40638
R12171 VDD.n5127 VDD.n5126 1.40638
R12172 VDD.n1026 VDD.n1025 1.40638
R12173 VDD.n7178 VDD.n7177 1.40638
R12174 VDD.n8117 VDD.n8116 1.40638
R12175 VDD.n8031 VDD.n8030 1.40638
R12176 VDD.n6848 VDD.n6847 1.36744
R12177 VDD.n7010 VDD.t460 1.35478
R12178 VDD.n7026 VDD.t461 1.35478
R12179 VDD.n7662 VDD.n7642 1.34143
R12180 VDD.n7038 VDD.n390 1.33475
R12181 VDD.n8184 VDD.n8143 1.33475
R12182 VDD.n7664 VDD.n7663 1.32491
R12183 VDD.n5602 VDD.n5601 1.31137
R12184 VDD.n4206 VDD.n4203 1.31137
R12185 VDD.n4215 VDD.n4212 1.31137
R12186 VDD.n5524 VDD.n5523 1.31137
R12187 VDD.n3924 VDD.n3921 1.31137
R12188 VDD.n3933 VDD.n3930 1.31137
R12189 VDD.n3433 VDD.n3430 1.31137
R12190 VDD.n3429 VDD.n3426 1.31137
R12191 VDD.n5378 VDD.n5372 1.31137
R12192 VDD.n3737 VDD.n3734 1.31137
R12193 VDD.n3733 VDD.n3730 1.31137
R12194 VDD.n5449 VDD.n5443 1.31137
R12195 VDD.n2944 VDD.n2941 1.31137
R12196 VDD.n2940 VDD.n2937 1.31137
R12197 VDD.n6186 VDD.n6180 1.31137
R12198 VDD.n3233 VDD.n3230 1.31137
R12199 VDD.n3229 VDD.n3226 1.31137
R12200 VDD.n5312 VDD.n5306 1.31137
R12201 VDD.n2866 VDD.n2863 1.31137
R12202 VDD.n2862 VDD.n2859 1.31137
R12203 VDD.n2559 VDD.n2553 1.31137
R12204 VDD.n6622 VDD.n6621 1.30325
R12205 VDD.n4381 VDD.n4242 1.23311
R12206 VDD.n5668 VDD.n5621 1.23311
R12207 VDD.n4391 VDD.n4237 1.23311
R12208 VDD.n5675 VDD.n5615 1.23311
R12209 VDD.n4401 VDD.n4231 1.23311
R12210 VDD.n5682 VDD.n5609 1.23311
R12211 VDD.n4411 VDD.n4225 1.23311
R12212 VDD.n5705 VDD.n5603 1.23311
R12213 VDD.n4447 VDD.n4215 1.23311
R12214 VDD.n5712 VDD.n5591 1.23311
R12215 VDD.n4457 VDD.n4197 1.23311
R12216 VDD.n5719 VDD.n5585 1.23311
R12217 VDD.n4467 VDD.n4191 1.23311
R12218 VDD.n5726 VDD.n5579 1.23311
R12219 VDD.n5731 VDD.n5576 1.23311
R12220 VDD.n4477 VDD.n4185 1.23311
R12221 VDD.n4484 VDD.n4182 1.23311
R12222 VDD.n5762 VDD.n5545 1.23311
R12223 VDD.n5767 VDD.n5542 1.23311
R12224 VDD.n4543 VDD.n3953 1.23311
R12225 VDD.n4550 VDD.n3950 1.23311
R12226 VDD.n5774 VDD.n5537 1.23311
R12227 VDD.n4560 VDD.n3945 1.23311
R12228 VDD.n5781 VDD.n5531 1.23311
R12229 VDD.n4570 VDD.n3939 1.23311
R12230 VDD.n5788 VDD.n5525 1.23311
R12231 VDD.n4580 VDD.n3933 1.23311
R12232 VDD.n5811 VDD.n5513 1.23311
R12233 VDD.n4616 VDD.n3911 1.23311
R12234 VDD.n5818 VDD.n5507 1.23311
R12235 VDD.n4626 VDD.n3905 1.23311
R12236 VDD.n5825 VDD.n5501 1.23311
R12237 VDD.n4636 VDD.n3899 1.23311
R12238 VDD.n5832 VDD.n5495 1.23311
R12239 VDD.n5837 VDD.n5492 1.23311
R12240 VDD.n4646 VDD.n3893 1.23311
R12241 VDD.n4653 VDD.n3890 1.23311
R12242 VDD.n6033 VDD.n5349 1.23311
R12243 VDD.n6026 VDD.n5355 1.23311
R12244 VDD.n4938 VDD.n3399 1.23311
R12245 VDD.n6019 VDD.n5361 1.23311
R12246 VDD.n4928 VDD.n3405 1.23311
R12247 VDD.n6012 VDD.n5367 1.23311
R12248 VDD.n4918 VDD.n3411 1.23311
R12249 VDD.n4882 VDD.n3433 1.23311
R12250 VDD.n5989 VDD.n5379 1.23311
R12251 VDD.n5982 VDD.n5385 1.23311
R12252 VDD.n4872 VDD.n3439 1.23311
R12253 VDD.n5975 VDD.n5391 1.23311
R12254 VDD.n4862 VDD.n3445 1.23311
R12255 VDD.n4852 VDD.n3450 1.23311
R12256 VDD.n4845 VDD.n3453 1.23311
R12257 VDD.n5968 VDD.n5396 1.23311
R12258 VDD.n5963 VDD.n5399 1.23311
R12259 VDD.n4800 VDD.n3704 1.23311
R12260 VDD.n4793 VDD.n3707 1.23311
R12261 VDD.n5930 VDD.n5423 1.23311
R12262 VDD.n5925 VDD.n5426 1.23311
R12263 VDD.n5918 VDD.n5432 1.23311
R12264 VDD.n4783 VDD.n3713 1.23311
R12265 VDD.n5911 VDD.n5438 1.23311
R12266 VDD.n4773 VDD.n3719 1.23311
R12267 VDD.n4763 VDD.n3737 1.23311
R12268 VDD.n5904 VDD.n5450 1.23311
R12269 VDD.n5881 VDD.n5456 1.23311
R12270 VDD.n4727 VDD.n3747 1.23311
R12271 VDD.n5874 VDD.n5462 1.23311
R12272 VDD.n4717 VDD.n3753 1.23311
R12273 VDD.n5867 VDD.n5468 1.23311
R12274 VDD.n4707 VDD.n3759 1.23311
R12275 VDD.n4697 VDD.n3764 1.23311
R12276 VDD.n4690 VDD.n3767 1.23311
R12277 VDD.n5860 VDD.n5473 1.23311
R12278 VDD.n5855 VDD.n5476 1.23311
R12279 VDD.n6043 VDD.n6042 1.23311
R12280 VDD.n4948 VDD.n3393 1.23311
R12281 VDD.n4955 VDD.n3390 1.23311
R12282 VDD.n6225 VDD.n6208 1.23311
R12283 VDD.n6232 VDD.n6205 1.23311
R12284 VDD.n5240 VDD.n2910 1.23311
R12285 VDD.n6239 VDD.n6199 1.23311
R12286 VDD.n5230 VDD.n2916 1.23311
R12287 VDD.n6246 VDD.n6193 1.23311
R12288 VDD.n5220 VDD.n2922 1.23311
R12289 VDD.n5184 VDD.n2944 1.23311
R12290 VDD.n6269 VDD.n6187 1.23311
R12291 VDD.n6276 VDD.n6175 1.23311
R12292 VDD.n5174 VDD.n2950 1.23311
R12293 VDD.n6283 VDD.n6169 1.23311
R12294 VDD.n5164 VDD.n2956 1.23311
R12295 VDD.n5154 VDD.n2961 1.23311
R12296 VDD.n5147 VDD.n2964 1.23311
R12297 VDD.n6290 VDD.n6163 1.23311
R12298 VDD.n6295 VDD.n6158 1.23311
R12299 VDD.n5102 VDD.n3200 1.23311
R12300 VDD.n5095 VDD.n3203 1.23311
R12301 VDD.n6136 VDD.n5286 1.23311
R12302 VDD.n6131 VDD.n5289 1.23311
R12303 VDD.n6124 VDD.n5295 1.23311
R12304 VDD.n5085 VDD.n3209 1.23311
R12305 VDD.n6117 VDD.n5301 1.23311
R12306 VDD.n5075 VDD.n3215 1.23311
R12307 VDD.n5065 VDD.n3233 1.23311
R12308 VDD.n6110 VDD.n5313 1.23311
R12309 VDD.n6087 VDD.n5319 1.23311
R12310 VDD.n5029 VDD.n3243 1.23311
R12311 VDD.n6080 VDD.n5325 1.23311
R12312 VDD.n5019 VDD.n3249 1.23311
R12313 VDD.n6073 VDD.n5331 1.23311
R12314 VDD.n5009 VDD.n3255 1.23311
R12315 VDD.n4999 VDD.n3260 1.23311
R12316 VDD.n4992 VDD.n3263 1.23311
R12317 VDD.n6066 VDD.n5336 1.23311
R12318 VDD.n6061 VDD.n5339 1.23311
R12319 VDD.n6220 VDD.n6219 1.23311
R12320 VDD.n5250 VDD.n2904 1.23311
R12321 VDD.n5257 VDD.n2901 1.23311
R12322 VDD.n2661 VDD.n2536 1.23311
R12323 VDD.n2654 VDD.n2542 1.23311
R12324 VDD.n6562 VDD.n2842 1.23311
R12325 VDD.n2647 VDD.n2548 1.23311
R12326 VDD.n6552 VDD.n2848 1.23311
R12327 VDD.n6542 VDD.n2866 1.23311
R12328 VDD.n2640 VDD.n2560 1.23311
R12329 VDD.n2617 VDD.n2566 1.23311
R12330 VDD.n6506 VDD.n2876 1.23311
R12331 VDD.n2610 VDD.n2572 1.23311
R12332 VDD.n6496 VDD.n2882 1.23311
R12333 VDD.n2603 VDD.n2578 1.23311
R12334 VDD.n6486 VDD.n2888 1.23311
R12335 VDD.n6476 VDD.n2893 1.23311
R12336 VDD.n6469 VDD.n2896 1.23311
R12337 VDD.n2596 VDD.n2583 1.23311
R12338 VDD.n2591 VDD.n2586 1.23311
R12339 VDD.n2671 VDD.n2670 1.23311
R12340 VDD.n6572 VDD.n2836 1.23311
R12341 VDD.n6579 VDD.n2833 1.23311
R12342 VDD.n206 VDD.n18 1.23311
R12343 VDD.n199 VDD.n21 1.23311
R12344 VDD.n150 VDD.n24 1.23311
R12345 VDD.n143 VDD.n27 1.23311
R12346 VDD.n4374 VDD.n4373 1.23311
R12347 VDD.n5661 VDD.n5626 1.23311
R12348 VDD.n5656 VDD.n5629 1.23311
R12349 VDD.n4392 VDD.t1152 1.2215
R12350 VDD.n4464 VDD.t910 1.2215
R12351 VDD.n4863 VDD.t682 1.2215
R12352 VDD.n4935 VDD.t1041 1.2215
R12353 VDD.n5010 VDD.t828 1.2215
R12354 VDD.n5082 VDD.t806 1.2215
R12355 VDD.n4561 VDD.t773 1.2215
R12356 VDD.n4633 VDD.t898 1.2215
R12357 VDD.n4708 VDD.t617 1.2215
R12358 VDD.n4780 VDD.t705 1.2215
R12359 VDD.n5165 VDD.t866 1.2215
R12360 VDD.n5237 VDD.t783 1.2215
R12361 VDD.n6487 VDD.t755 1.2215
R12362 VDD.n6559 VDD.t781 1.2215
R12363 VDD.n7045 VDD.n312 1.21354
R12364 VDD.n7052 VDD.n308 1.21354
R12365 VDD.n6986 VDD.n6867 1.21354
R12366 VDD.n6993 VDD.n6863 1.21354
R12367 VDD.t436 VDD.t561 1.15992
R12368 VDD.t573 VDD.t530 1.15992
R12369 VDD.t476 VDD.t573 1.15992
R12370 VDD.t862 VDD.t559 1.15992
R12371 VDD.n7662 VDD.n7643 1.15696
R12372 VDD.n6602 VDD.n6601 1.15363
R12373 VDD.n6604 VDD.n6603 1.15363
R12374 VDD.n6605 VDD.n6604 1.15363
R12375 VDD.n6607 VDD.n6606 1.15363
R12376 VDD.n6608 VDD.n6607 1.15363
R12377 VDD.n6856 VDD.n6855 1.14664
R12378 VDD.n8166 VDD.n8165 1.13137
R12379 VDD.n8177 VDD.n8154 1.13137
R12380 VDD.n8189 VDD.n7903 1.13137
R12381 VDD.n7076 VDD.n7057 1.13137
R12382 VDD.n7069 VDD.n7060 1.13137
R12383 VDD.n8198 VDD.n7892 1.13137
R12384 VDD.n8203 VDD.n7890 1.13137
R12385 VDD.n6708 VDD.n6647 1.1255
R12386 VDD.n799 VDD.n554 1.1255
R12387 VDD.n6657 VDD.n6648 1.1255
R12388 VDD.n806 VDD.n550 1.1255
R12389 VDD.n6652 VDD.n6649 1.1255
R12390 VDD.n594 VDD.n560 1.1255
R12391 VDD.n589 VDD.n564 1.1255
R12392 VDD.n582 VDD.n567 1.1255
R12393 VDD.n772 VDD.n746 1.1255
R12394 VDD.n575 VDD.n570 1.1255
R12395 VDD.n762 VDD.n755 1.1255
R12396 VDD.n884 VDD.n879 1.1255
R12397 VDD.n1062 VDD.n1055 1.1255
R12398 VDD.n891 VDD.n876 1.1255
R12399 VDD.n1072 VDD.n1046 1.1255
R12400 VDD.n1089 VDD.n1033 1.1255
R12401 VDD.n898 VDD.n873 1.1255
R12402 VDD.n1082 VDD.n1037 1.1255
R12403 VDD.n903 VDD.n872 1.1255
R12404 VDD.n6703 VDD.n6702 1.1255
R12405 VDD.n6636 VDD.n6632 1.1255
R12406 VDD.n6643 VDD.n6628 1.1255
R12407 VDD.n734 VDD.n732 1.12396
R12408 VDD.n6976 VDD.n6975 1.12396
R12409 VDD.n6455 VDD.n6451 1.12377
R12410 VDD.n6455 VDD.n6454 1.12377
R12411 VDD.n6849 VDD.n6848 1.12377
R12412 VDD.n40 VDD.n28 1.12377
R12413 VDD.n6977 VDD.n6976 1.12377
R12414 VDD.n1063 VDD.t946 1.10231
R12415 VDD.n763 VDD.t954 1.10231
R12416 VDD.n6311 VDD.n6310 1.1018
R12417 VDD.n5944 VDD.n5943 1.1016
R12418 VDD.n5950 VDD.n5949 1.1016
R12419 VDD.n401 VDD.n400 1.09615
R12420 VDD.n6627 VDD.n6624 1.09028
R12421 VDD.n549 VDD.n546 1.09028
R12422 VDD.n553 VDD.n552 1.09028
R12423 VDD.n558 VDD.n557 1.09028
R12424 VDD.n562 VDD.n561 1.09028
R12425 VDD.n1036 VDD.n1035 1.09028
R12426 VDD.n1032 VDD.n1031 1.09028
R12427 VDD.n6631 VDD.n6630 1.09028
R12428 VDD.n8310 VDD.n7232 1.07267
R12429 VDD.n7199 VDD.n11 1.07267
R12430 VDD.n7189 VDD.n15 1.07267
R12431 VDD.n8324 VDD.n8323 1.07267
R12432 VDD.n312 VDD.n311 1.06093
R12433 VDD.n307 VDD.n304 1.06093
R12434 VDD.n308 VDD.n307 1.06093
R12435 VDD.n311 VDD.n310 1.06093
R12436 VDD.n6867 VDD.n6866 1.06093
R12437 VDD.n6862 VDD.n6859 1.06093
R12438 VDD.n6863 VDD.n6862 1.06093
R12439 VDD.n6866 VDD.n6865 1.06093
R12440 VDD.n7639 VDD.n7638 1.0274
R12441 VDD.n2393 VDD.t524 1.02677
R12442 VDD.n2411 VDD.t109 1.02677
R12443 VDD.n392 VDD.n391 1.02572
R12444 VDD.n7969 VDD.n7968 1.00811
R12445 VDD.n4242 VDD.n4241 0.992457
R12446 VDD.n5579 VDD.n5578 0.992457
R12447 VDD.n5576 VDD.n5575 0.992457
R12448 VDD.n5575 VDD.n5572 0.992457
R12449 VDD.n4181 VDD.n4178 0.992457
R12450 VDD.n5578 VDD.n5577 0.992457
R12451 VDD.n4184 VDD.n4183 0.992457
R12452 VDD.n4185 VDD.n4184 0.992457
R12453 VDD.n4182 VDD.n4181 0.992457
R12454 VDD.n5545 VDD.n5544 0.992457
R12455 VDD.n5542 VDD.n5541 0.992457
R12456 VDD.n5541 VDD.n5538 0.992457
R12457 VDD.n3949 VDD.n3946 0.992457
R12458 VDD.n5544 VDD.n5543 0.992457
R12459 VDD.n3952 VDD.n3951 0.992457
R12460 VDD.n3953 VDD.n3952 0.992457
R12461 VDD.n3950 VDD.n3949 0.992457
R12462 VDD.n5495 VDD.n5494 0.992457
R12463 VDD.n5492 VDD.n5491 0.992457
R12464 VDD.n5491 VDD.n5488 0.992457
R12465 VDD.n3889 VDD.n3886 0.992457
R12466 VDD.n5494 VDD.n5493 0.992457
R12467 VDD.n3892 VDD.n3891 0.992457
R12468 VDD.n3893 VDD.n3892 0.992457
R12469 VDD.n3890 VDD.n3889 0.992457
R12470 VDD.n5349 VDD.n5348 0.992457
R12471 VDD.n3450 VDD.n3449 0.992457
R12472 VDD.n5398 VDD.n5397 0.992457
R12473 VDD.n3452 VDD.n3451 0.992457
R12474 VDD.n3453 VDD.n3452 0.992457
R12475 VDD.n5396 VDD.n5395 0.992457
R12476 VDD.n5395 VDD.n5392 0.992457
R12477 VDD.n3449 VDD.n3448 0.992457
R12478 VDD.n5399 VDD.n5398 0.992457
R12479 VDD.n3704 VDD.n3703 0.992457
R12480 VDD.n5425 VDD.n5424 0.992457
R12481 VDD.n3706 VDD.n3705 0.992457
R12482 VDD.n3707 VDD.n3706 0.992457
R12483 VDD.n5423 VDD.n5422 0.992457
R12484 VDD.n5422 VDD.n5419 0.992457
R12485 VDD.n3703 VDD.n3702 0.992457
R12486 VDD.n5426 VDD.n5425 0.992457
R12487 VDD.n3764 VDD.n3763 0.992457
R12488 VDD.n5475 VDD.n5474 0.992457
R12489 VDD.n3766 VDD.n3765 0.992457
R12490 VDD.n3767 VDD.n3766 0.992457
R12491 VDD.n5473 VDD.n5472 0.992457
R12492 VDD.n5472 VDD.n5469 0.992457
R12493 VDD.n3763 VDD.n3762 0.992457
R12494 VDD.n5476 VDD.n5475 0.992457
R12495 VDD.n6042 VDD.n6041 0.992457
R12496 VDD.n6041 VDD.n6038 0.992457
R12497 VDD.n3389 VDD.n3386 0.992457
R12498 VDD.n5348 VDD.n5347 0.992457
R12499 VDD.n3392 VDD.n3391 0.992457
R12500 VDD.n3393 VDD.n3392 0.992457
R12501 VDD.n3390 VDD.n3389 0.992457
R12502 VDD.n6208 VDD.n6207 0.992457
R12503 VDD.n2961 VDD.n2960 0.992457
R12504 VDD.n6157 VDD.n6156 0.992457
R12505 VDD.n2963 VDD.n2962 0.992457
R12506 VDD.n2964 VDD.n2963 0.992457
R12507 VDD.n6163 VDD.n6162 0.992457
R12508 VDD.n6162 VDD.n6159 0.992457
R12509 VDD.n2960 VDD.n2959 0.992457
R12510 VDD.n6158 VDD.n6157 0.992457
R12511 VDD.n3200 VDD.n3199 0.992457
R12512 VDD.n5288 VDD.n5287 0.992457
R12513 VDD.n3202 VDD.n3201 0.992457
R12514 VDD.n3203 VDD.n3202 0.992457
R12515 VDD.n5286 VDD.n5285 0.992457
R12516 VDD.n5285 VDD.n5282 0.992457
R12517 VDD.n3199 VDD.n3198 0.992457
R12518 VDD.n5289 VDD.n5288 0.992457
R12519 VDD.n3260 VDD.n3259 0.992457
R12520 VDD.n5338 VDD.n5337 0.992457
R12521 VDD.n3262 VDD.n3261 0.992457
R12522 VDD.n3263 VDD.n3262 0.992457
R12523 VDD.n5336 VDD.n5335 0.992457
R12524 VDD.n5335 VDD.n5332 0.992457
R12525 VDD.n3259 VDD.n3258 0.992457
R12526 VDD.n5339 VDD.n5338 0.992457
R12527 VDD.n6219 VDD.n6218 0.992457
R12528 VDD.n6218 VDD.n6215 0.992457
R12529 VDD.n2900 VDD.n2897 0.992457
R12530 VDD.n6207 VDD.n6206 0.992457
R12531 VDD.n2903 VDD.n2902 0.992457
R12532 VDD.n2904 VDD.n2903 0.992457
R12533 VDD.n2901 VDD.n2900 0.992457
R12534 VDD.n2536 VDD.n2535 0.992457
R12535 VDD.n2893 VDD.n2892 0.992457
R12536 VDD.n2585 VDD.n2584 0.992457
R12537 VDD.n2895 VDD.n2894 0.992457
R12538 VDD.n2896 VDD.n2895 0.992457
R12539 VDD.n2583 VDD.n2582 0.992457
R12540 VDD.n2582 VDD.n2579 0.992457
R12541 VDD.n2892 VDD.n2891 0.992457
R12542 VDD.n2586 VDD.n2585 0.992457
R12543 VDD.n2670 VDD.n2669 0.992457
R12544 VDD.n2669 VDD.n2666 0.992457
R12545 VDD.n2832 VDD.n2829 0.992457
R12546 VDD.n2535 VDD.n2534 0.992457
R12547 VDD.n2835 VDD.n2834 0.992457
R12548 VDD.n2836 VDD.n2835 0.992457
R12549 VDD.n2833 VDD.n2832 0.992457
R12550 VDD.n5628 VDD.n5627 0.992457
R12551 VDD.n4372 VDD.n4371 0.992457
R12552 VDD.n4373 VDD.n4372 0.992457
R12553 VDD.n5626 VDD.n5625 0.992457
R12554 VDD.n5625 VDD.n5622 0.992457
R12555 VDD.n4241 VDD.n4240 0.992457
R12556 VDD.n5629 VDD.n5628 0.992457
R12557 VDD.n6857 VDD.n544 0.932563
R12558 VDD.n7881 VDD.n7851 0.914272
R12559 VDD.n7663 VDD.n7662 0.914044
R12560 VDD.n7881 VDD.n7876 0.914044
R12561 VDD.n8251 VDD.n7886 0.8809
R12562 VDD.n2685 VDD.n2684 0.878601
R12563 VDD.n4355 VDD.n4354 0.878601
R12564 VDD.n5645 VDD.n5644 0.878601
R12565 VDD.n1460 VDD.n1459 0.875507
R12566 VDD.n1242 VDD.n1241 0.875507
R12567 VDD.n2533 VDD.n2532 0.875507
R12568 VDD.n2048 VDD.n2047 0.875507
R12569 VDD.n4821 VDD.n4820 0.873539
R12570 VDD.n6155 VDD.n6154 0.873539
R12571 VDD.n6151 VDD.n6150 0.873539
R12572 VDD.n5121 VDD.n5120 0.873539
R12573 VDD.n734 VDD.n733 0.873539
R12574 VDD.n41 VDD.n40 0.873539
R12575 VDD.n8295 VDD.n8294 0.873539
R12576 VDD.n539 VDD.n538 0.873539
R12577 VDD.n1656 VDD.n1655 0.873539
R12578 VDD.n1528 VDD.n1527 0.873539
R12579 VDD.n2151 VDD.n2150 0.873539
R12580 VDD.n2342 VDD.n2341 0.873539
R12581 VDD.n4519 VDD.n4518 0.873539
R12582 VDD.n4525 VDD.n4524 0.873539
R12583 VDD.n5746 VDD.n5745 0.873539
R12584 VDD.n5750 VDD.n5749 0.873539
R12585 VDD.n4671 VDD.n4670 0.873308
R12586 VDD.n4825 VDD.n4824 0.873308
R12587 VDD.n4973 VDD.n4972 0.873308
R12588 VDD.n5126 VDD.n5125 0.873308
R12589 VDD.n6597 VDD.n6596 0.873308
R12590 VDD.n1024 VDD.n1009 0.873308
R12591 VDD.n7177 VDD.n7176 0.873308
R12592 VDD.n8116 VDD.n8115 0.873308
R12593 VDD.n1025 VDD.n1024 0.873308
R12594 VDD.n380 VDD.t568 0.870065
R12595 VDD.n405 VDD.n404 0.869196
R12596 VDD.n7881 VDD.n7875 0.852583
R12597 VDD.n7662 VDD.n7661 0.852583
R12598 VDD.n7977 VDD.n7976 0.851587
R12599 VDD.n7975 VDD.n7974 0.851587
R12600 VDD.n7973 VDD.n7959 0.851587
R12601 VDD.n7979 VDD.n7978 0.851587
R12602 VDD.n554 VDD.n553 0.847674
R12603 VDD.n550 VDD.n549 0.847674
R12604 VDD.n1033 VDD.n1032 0.847674
R12605 VDD.n1037 VDD.n1036 0.847674
R12606 VDD.n6632 VDD.n6631 0.847674
R12607 VDD.n6628 VDD.n6627 0.847674
R12608 VDD.n6610 VDD.n6609 0.8465
R12609 VDD.n7967 VDD.n7966 0.845717
R12610 VDD.n4408 VDD.t847 0.814501
R12611 VDD.n4448 VDD.t849 0.814501
R12612 VDD.n4879 VDD.t826 0.814501
R12613 VDD.n4919 VDD.t767 0.814501
R12614 VDD.n5026 VDD.t634 0.814501
R12615 VDD.n5066 VDD.t629 0.814501
R12616 VDD.n4577 VDD.t592 0.814501
R12617 VDD.n4617 VDD.t599 0.814501
R12618 VDD.n4724 VDD.t925 0.814501
R12619 VDD.n4764 VDD.t907 0.814501
R12620 VDD.n5181 VDD.t597 0.814501
R12621 VDD.n5221 VDD.t707 0.814501
R12622 VDD.n6503 VDD.t680 0.814501
R12623 VDD.n6543 VDD.t797 0.814501
R12624 VDD.n7662 VDD.n7651 0.709103
R12625 VDD.n7662 VDD.n7650 0.709103
R12626 VDD.n7662 VDD.n7649 0.709103
R12627 VDD.n7662 VDD.n7648 0.709103
R12628 VDD.n7662 VDD.n7647 0.709103
R12629 VDD.n7662 VDD.n7646 0.709103
R12630 VDD.n7662 VDD.n7645 0.709103
R12631 VDD.n7662 VDD.n7644 0.709103
R12632 VDD.n7881 VDD.n7852 0.709103
R12633 VDD.n7881 VDD.n7853 0.709103
R12634 VDD.n7881 VDD.n7854 0.709103
R12635 VDD.n7881 VDD.n7855 0.709103
R12636 VDD.n7881 VDD.n7856 0.709103
R12637 VDD.n7881 VDD.n7857 0.709103
R12638 VDD.n7881 VDD.n7858 0.709103
R12639 VDD.n7881 VDD.n7859 0.709103
R12640 VDD.n7881 VDD.n7860 0.709103
R12641 VDD.n7881 VDD.n7861 0.709103
R12642 VDD.n7881 VDD.n7863 0.709103
R12643 VDD.n7881 VDD.n7866 0.709103
R12644 VDD.n7881 VDD.n7869 0.709103
R12645 VDD.n7881 VDD.n7872 0.709103
R12646 VDD.n7886 VDD.n7883 0.709103
R12647 VDD.n7662 VDD.n7660 0.708865
R12648 VDD.n7662 VDD.n7659 0.708865
R12649 VDD.n7662 VDD.n7658 0.708865
R12650 VDD.n7662 VDD.n7657 0.708865
R12651 VDD.n7662 VDD.n7656 0.708865
R12652 VDD.n7662 VDD.n7655 0.708865
R12653 VDD.n7662 VDD.n7654 0.708865
R12654 VDD.n7662 VDD.n7653 0.708865
R12655 VDD.n7662 VDD.n7652 0.708865
R12656 VDD.n7881 VDD.n7879 0.708865
R12657 VDD.n7881 VDD.n7878 0.708865
R12658 VDD.n7881 VDD.n7877 0.708865
R12659 VDD.n7881 VDD.n7880 0.708865
R12660 VDD.n7882 VDD.n7881 0.708865
R12661 VDD.n9 VDD.n8 0.700935
R12662 VDD.n13 VDD.n12 0.700935
R12663 VDD.n8321 VDD.n8320 0.700935
R12664 VDD.n7890 VDD.n7889 0.700935
R12665 VDD.n8251 VDD.n7234 0.684371
R12666 VDD.n2340 VDD.n2339 0.684371
R12667 VDD.n2149 VDD.n2148 0.684371
R12668 VDD.n2046 VDD.n2045 0.684371
R12669 VDD.n6434 VDD.n6433 0.684371
R12670 VDD.n6314 VDD.n6312 0.684371
R12671 VDD.n735 VDD.n734 0.684371
R12672 VDD.n8294 VDD.n8293 0.684371
R12673 VDD.n8294 VDD.n8292 0.684371
R12674 VDD.n8294 VDD.n8291 0.684371
R12675 VDD.n8294 VDD.n8290 0.684371
R12676 VDD.n8294 VDD.n8289 0.684371
R12677 VDD.n8294 VDD.n8288 0.684371
R12678 VDD.n8294 VDD.n8287 0.684371
R12679 VDD.n8294 VDD.n8286 0.684371
R12680 VDD.n538 VDD.n537 0.684371
R12681 VDD.n538 VDD.n536 0.684371
R12682 VDD.n538 VDD.n535 0.684371
R12683 VDD.n538 VDD.n534 0.684371
R12684 VDD.n538 VDD.n533 0.684371
R12685 VDD.n2339 VDD.n2336 0.684371
R12686 VDD.n2148 VDD.n2145 0.684371
R12687 VDD.n2045 VDD.n2044 0.684371
R12688 VDD.n2045 VDD.n2043 0.684371
R12689 VDD.n2045 VDD.n2042 0.684371
R12690 VDD.n2045 VDD.n2041 0.684371
R12691 VDD.n2045 VDD.n2040 0.684371
R12692 VDD.n2045 VDD.n2039 0.684371
R12693 VDD.n2045 VDD.n2038 0.684371
R12694 VDD.n2045 VDD.n2037 0.684371
R12695 VDD.n2045 VDD.n2036 0.684371
R12696 VDD.n2045 VDD.n2035 0.684371
R12697 VDD.n2045 VDD.n2034 0.684371
R12698 VDD.n2045 VDD.n2033 0.684371
R12699 VDD.n4516 VDD.n4515 0.684132
R12700 VDD.n4516 VDD.n4514 0.684132
R12701 VDD.n4516 VDD.n4513 0.684132
R12702 VDD.n4516 VDD.n4512 0.684132
R12703 VDD.n4516 VDD.n4511 0.684132
R12704 VDD.n4516 VDD.n4510 0.684132
R12705 VDD.n4516 VDD.n4509 0.684132
R12706 VDD.n4516 VDD.n4508 0.684132
R12707 VDD.n4516 VDD.n4507 0.684132
R12708 VDD.n4516 VDD.n4506 0.684132
R12709 VDD.n4516 VDD.n4505 0.684132
R12710 VDD.n4516 VDD.n4504 0.684132
R12711 VDD.n4516 VDD.n4503 0.684132
R12712 VDD.n4516 VDD.n4502 0.684132
R12713 VDD.n5346 VDD.n5344 0.684132
R12714 VDD.n5483 VDD.n5481 0.684132
R12715 VDD.n1024 VDD.n1010 0.684132
R12716 VDD.n1024 VDD.n1011 0.684132
R12717 VDD.n1024 VDD.n1012 0.684132
R12718 VDD.n1024 VDD.n1013 0.684132
R12719 VDD.n1024 VDD.n1014 0.684132
R12720 VDD.n1024 VDD.n1015 0.684132
R12721 VDD.n1024 VDD.n1016 0.684132
R12722 VDD.n1024 VDD.n1017 0.684132
R12723 VDD.n1024 VDD.n1018 0.684132
R12724 VDD.n1024 VDD.n1019 0.684132
R12725 VDD.n1024 VDD.n1020 0.684132
R12726 VDD.n1024 VDD.n1021 0.684132
R12727 VDD.n1024 VDD.n1022 0.684132
R12728 VDD.n1024 VDD.n1023 0.684132
R12729 VDD.n8251 VDD.n7237 0.684132
R12730 VDD.n7176 VDD.n7166 0.684132
R12731 VDD.n7176 VDD.n7167 0.684132
R12732 VDD.n7176 VDD.n7168 0.684132
R12733 VDD.n7176 VDD.n7169 0.684132
R12734 VDD.n7176 VDD.n7170 0.684132
R12735 VDD.n7176 VDD.n7171 0.684132
R12736 VDD.n7176 VDD.n7172 0.684132
R12737 VDD.n7176 VDD.n7173 0.684132
R12738 VDD.n7176 VDD.n7174 0.684132
R12739 VDD.n7176 VDD.n7175 0.684132
R12740 VDD.n299 VDD.n298 0.684132
R12741 VDD.n299 VDD.n297 0.684132
R12742 VDD.n299 VDD.n296 0.684132
R12743 VDD.n299 VDD.n295 0.684132
R12744 VDD.n299 VDD.n294 0.684132
R12745 VDD.n299 VDD.n293 0.684132
R12746 VDD.n299 VDD.n292 0.684132
R12747 VDD.n299 VDD.n291 0.684132
R12748 VDD.n300 VDD.n299 0.684132
R12749 VDD.n8115 VDD.n8110 0.684132
R12750 VDD.n8115 VDD.n8111 0.684132
R12751 VDD.n8115 VDD.n8112 0.684132
R12752 VDD.n8115 VDD.n8113 0.684132
R12753 VDD.n8115 VDD.n8114 0.684132
R12754 VDD.n2530 VDD.n2518 0.684132
R12755 VDD.n2530 VDD.n2519 0.684132
R12756 VDD.n2530 VDD.n2520 0.684132
R12757 VDD.n2530 VDD.n2521 0.684132
R12758 VDD.n2530 VDD.n2522 0.684132
R12759 VDD.n2530 VDD.n2523 0.684132
R12760 VDD.n2530 VDD.n2524 0.684132
R12761 VDD.n2530 VDD.n2525 0.684132
R12762 VDD.n2530 VDD.n2526 0.684132
R12763 VDD.n2530 VDD.n2527 0.684132
R12764 VDD.n2530 VDD.n2528 0.684132
R12765 VDD.n2530 VDD.n2529 0.684132
R12766 VDD.n2531 VDD.n2530 0.684132
R12767 VDD.n4517 VDD.n4516 0.684132
R12768 VDD.n1453 VDD.n1452 0.6755
R12769 VDD.n1450 VDD.n1449 0.6755
R12770 VDD.n1449 VDD.n1446 0.6755
R12771 VDD.n1127 VDD.n1124 0.6755
R12772 VDD.n1452 VDD.n1451 0.6755
R12773 VDD.n1130 VDD.n1129 0.6755
R12774 VDD.n1131 VDD.n1130 0.6755
R12775 VDD.n1128 VDD.n1127 0.6755
R12776 VDD.n1445 VDD.n1444 0.6755
R12777 VDD.n1442 VDD.n1441 0.6755
R12778 VDD.n1444 VDD.n1443 0.6755
R12779 VDD.n1353 VDD.n1352 0.6755
R12780 VDD.n1348 VDD.n1347 0.6755
R12781 VDD.n1347 VDD.n1344 0.6755
R12782 VDD.n1101 VDD.n1098 0.6755
R12783 VDD.n1352 VDD.n1351 0.6755
R12784 VDD.n1105 VDD.n1104 0.6755
R12785 VDD.n1107 VDD.n1105 0.6755
R12786 VDD.n1102 VDD.n1101 0.6755
R12787 VDD.n5603 VDD.n5602 0.673543
R12788 VDD.n4212 VDD.n4206 0.673543
R12789 VDD.n5525 VDD.n5524 0.673543
R12790 VDD.n3930 VDD.n3924 0.673543
R12791 VDD.n3430 VDD.n3429 0.673543
R12792 VDD.n5379 VDD.n5378 0.673543
R12793 VDD.n3734 VDD.n3733 0.673543
R12794 VDD.n5450 VDD.n5449 0.673543
R12795 VDD.n2941 VDD.n2940 0.673543
R12796 VDD.n6187 VDD.n6186 0.673543
R12797 VDD.n3230 VDD.n3229 0.673543
R12798 VDD.n5313 VDD.n5312 0.673543
R12799 VDD.n2863 VDD.n2862 0.673543
R12800 VDD.n2560 VDD.n2559 0.673543
R12801 VDD VDD.n6307 0.666861
R12802 VDD.n5602 VDD.n5598 0.626587
R12803 VDD.n4203 VDD.n4202 0.626587
R12804 VDD.n4212 VDD.n4211 0.626587
R12805 VDD.n5524 VDD.n5520 0.626587
R12806 VDD.n3921 VDD.n3920 0.626587
R12807 VDD.n3930 VDD.n3929 0.626587
R12808 VDD.n3430 VDD.n3420 0.626587
R12809 VDD.n3426 VDD.n3425 0.626587
R12810 VDD.n5378 VDD.n5377 0.626587
R12811 VDD.n3734 VDD.n3724 0.626587
R12812 VDD.n3730 VDD.n3729 0.626587
R12813 VDD.n5449 VDD.n5448 0.626587
R12814 VDD.n2941 VDD.n2931 0.626587
R12815 VDD.n2937 VDD.n2936 0.626587
R12816 VDD.n6186 VDD.n6185 0.626587
R12817 VDD.n3230 VDD.n3220 0.626587
R12818 VDD.n3226 VDD.n3225 0.626587
R12819 VDD.n5312 VDD.n5311 0.626587
R12820 VDD.n2863 VDD.n2853 0.626587
R12821 VDD.n2859 VDD.n2858 0.626587
R12822 VDD.n2559 VDD.n2558 0.626587
R12823 VDD.n2452 VDD.t121 0.616264
R12824 VDD.n5617 VDD.t665 0.607167
R12825 VDD.n5617 VDD.n5616 0.607167
R12826 VDD.n5619 VDD.t1376 0.607167
R12827 VDD.n5619 VDD.n5618 0.607167
R12828 VDD.n4233 VDD.t1436 0.607167
R12829 VDD.n4233 VDD.n4232 0.607167
R12830 VDD.n4236 VDD.t1093 0.607167
R12831 VDD.n4236 VDD.n4235 0.607167
R12832 VDD.n5611 VDD.t872 0.607167
R12833 VDD.n5611 VDD.n5610 0.607167
R12834 VDD.n5613 VDD.t616 0.607167
R12835 VDD.n5613 VDD.n5612 0.607167
R12836 VDD.n4227 VDD.t1082 0.607167
R12837 VDD.n4227 VDD.n4226 0.607167
R12838 VDD.n4230 VDD.t1043 0.607167
R12839 VDD.n4230 VDD.n4229 0.607167
R12840 VDD.n5605 VDD.t1335 0.607167
R12841 VDD.n5605 VDD.n5604 0.607167
R12842 VDD.n5607 VDD.t928 0.607167
R12843 VDD.n5607 VDD.n5606 0.607167
R12844 VDD.n4221 VDD.t848 0.607167
R12845 VDD.n4221 VDD.n4220 0.607167
R12846 VDD.n4224 VDD.t1068 0.607167
R12847 VDD.n4224 VDD.n4223 0.607167
R12848 VDD.n4219 VDD.t904 0.607167
R12849 VDD.n4219 VDD.n4218 0.607167
R12850 VDD.n4217 VDD.t1311 0.607167
R12851 VDD.n4217 VDD.n4216 0.607167
R12852 VDD.n4214 VDD.t1382 0.607167
R12853 VDD.n4214 VDD.n4213 0.607167
R12854 VDD.n4205 VDD.t677 0.607167
R12855 VDD.n4205 VDD.n4204 0.607167
R12856 VDD.n5600 VDD.t1427 0.607167
R12857 VDD.n5600 VDD.n5599 0.607167
R12858 VDD.n5593 VDD.t810 0.607167
R12859 VDD.n5593 VDD.n5592 0.607167
R12860 VDD.n5597 VDD.t1214 0.607167
R12861 VDD.n5597 VDD.n5596 0.607167
R12862 VDD.n5595 VDD.t713 0.607167
R12863 VDD.n5595 VDD.n5594 0.607167
R12864 VDD.n4201 VDD.t901 0.607167
R12865 VDD.n4201 VDD.n4200 0.607167
R12866 VDD.n4199 VDD.t1253 0.607167
R12867 VDD.n4199 VDD.n4198 0.607167
R12868 VDD.n4210 VDD.t1412 0.607167
R12869 VDD.n4210 VDD.n4209 0.607167
R12870 VDD.n4208 VDD.t1220 0.607167
R12871 VDD.n4208 VDD.n4207 0.607167
R12872 VDD.n5587 VDD.t915 0.607167
R12873 VDD.n5587 VDD.n5586 0.607167
R12874 VDD.n5589 VDD.t1298 0.607167
R12875 VDD.n5589 VDD.n5588 0.607167
R12876 VDD.n4193 VDD.t1088 0.607167
R12877 VDD.n4193 VDD.n4192 0.607167
R12878 VDD.n4196 VDD.t1303 0.607167
R12879 VDD.n4196 VDD.n4195 0.607167
R12880 VDD.n5581 VDD.t1319 0.607167
R12881 VDD.n5581 VDD.n5580 0.607167
R12882 VDD.n5583 VDD.t1362 0.607167
R12883 VDD.n5583 VDD.n5582 0.607167
R12884 VDD.n4187 VDD.t911 0.607167
R12885 VDD.n4187 VDD.n4186 0.607167
R12886 VDD.n4190 VDD.t1320 0.607167
R12887 VDD.n4190 VDD.n4189 0.607167
R12888 VDD.n5533 VDD.t1190 0.607167
R12889 VDD.n5533 VDD.n5532 0.607167
R12890 VDD.n5535 VDD.t1264 0.607167
R12891 VDD.n5535 VDD.n5534 0.607167
R12892 VDD.n3941 VDD.t1006 0.607167
R12893 VDD.n3941 VDD.n3940 0.607167
R12894 VDD.n3944 VDD.t1271 0.607167
R12895 VDD.n3944 VDD.n3943 0.607167
R12896 VDD.n5527 VDD.t1099 0.607167
R12897 VDD.n5527 VDD.n5526 0.607167
R12898 VDD.n5529 VDD.t1420 0.607167
R12899 VDD.n5529 VDD.n5528 0.607167
R12900 VDD.n3935 VDD.t1238 0.607167
R12901 VDD.n3935 VDD.n3934 0.607167
R12902 VDD.n3938 VDD.t1424 0.607167
R12903 VDD.n3938 VDD.n3937 0.607167
R12904 VDD.n3932 VDD.t593 0.607167
R12905 VDD.n3932 VDD.n3931 0.607167
R12906 VDD.n3923 VDD.t1196 0.607167
R12907 VDD.n3923 VDD.n3922 0.607167
R12908 VDD.n5522 VDD.t879 0.607167
R12909 VDD.n5522 VDD.n5521 0.607167
R12910 VDD.n5515 VDD.t1384 0.607167
R12911 VDD.n5515 VDD.n5514 0.607167
R12912 VDD.n5517 VDD.t633 0.607167
R12913 VDD.n5517 VDD.n5516 0.607167
R12914 VDD.n5519 VDD.t1221 0.607167
R12915 VDD.n5519 VDD.n5518 0.607167
R12916 VDD.n3917 VDD.t1162 0.607167
R12917 VDD.n3917 VDD.n3916 0.607167
R12918 VDD.n3919 VDD.t1312 0.607167
R12919 VDD.n3919 VDD.n3918 0.607167
R12920 VDD.n3926 VDD.t1283 0.607167
R12921 VDD.n3926 VDD.n3925 0.607167
R12922 VDD.n3928 VDD.t734 0.607167
R12923 VDD.n3928 VDD.n3927 0.607167
R12924 VDD.n3915 VDD.t1127 0.607167
R12925 VDD.n3915 VDD.n3914 0.607167
R12926 VDD.n3913 VDD.t720 0.607167
R12927 VDD.n3913 VDD.n3912 0.607167
R12928 VDD.n5509 VDD.t1215 0.607167
R12929 VDD.n5509 VDD.n5508 0.607167
R12930 VDD.n5511 VDD.t902 0.607167
R12931 VDD.n5511 VDD.n5510 0.607167
R12932 VDD.n3907 VDD.t1204 0.607167
R12933 VDD.n3907 VDD.n3906 0.607167
R12934 VDD.n3910 VDD.t886 0.607167
R12935 VDD.n3910 VDD.n3909 0.607167
R12936 VDD.n5503 VDD.t1004 0.607167
R12937 VDD.n5503 VDD.n5502 0.607167
R12938 VDD.n5505 VDD.t1272 0.607167
R12939 VDD.n5505 VDD.n5504 0.607167
R12940 VDD.n3901 VDD.t814 0.607167
R12941 VDD.n3901 VDD.n3900 0.607167
R12942 VDD.n3904 VDD.t1430 0.607167
R12943 VDD.n3904 VDD.n3903 0.607167
R12944 VDD.n5497 VDD.t1435 0.607167
R12945 VDD.n5497 VDD.n5496 0.607167
R12946 VDD.n5499 VDD.t1087 0.607167
R12947 VDD.n5499 VDD.n5498 0.607167
R12948 VDD.n3895 VDD.t899 0.607167
R12949 VDD.n3895 VDD.n3894 0.607167
R12950 VDD.n3898 VDD.t1001 0.607167
R12951 VDD.n3898 VDD.n3897 0.607167
R12952 VDD.n2870 VDD.t927 0.607167
R12953 VDD.n2870 VDD.n2869 0.607167
R12954 VDD.n2868 VDD.t1291 0.607167
R12955 VDD.n2868 VDD.n2867 0.607167
R12956 VDD.n3237 VDD.t1141 0.607167
R12957 VDD.n3237 VDD.n3236 0.607167
R12958 VDD.n3235 VDD.t789 0.607167
R12959 VDD.n3235 VDD.n3234 0.607167
R12960 VDD.n2926 VDD.t777 0.607167
R12961 VDD.n2926 VDD.n2925 0.607167
R12962 VDD.n2924 VDD.t1297 0.607167
R12963 VDD.n2924 VDD.n2923 0.607167
R12964 VDD.n3741 VDD.t823 0.607167
R12965 VDD.n3741 VDD.n3740 0.607167
R12966 VDD.n3739 VDD.t658 0.607167
R12967 VDD.n3739 VDD.n3738 0.607167
R12968 VDD.n3415 VDD.t1363 0.607167
R12969 VDD.n3415 VDD.n3414 0.607167
R12970 VDD.n3413 VDD.t1396 0.607167
R12971 VDD.n3413 VDD.n3412 0.607167
R12972 VDD.n5351 VDD.t1081 0.607167
R12973 VDD.n5351 VDD.n5350 0.607167
R12974 VDD.n5353 VDD.t1042 0.607167
R12975 VDD.n5353 VDD.n5352 0.607167
R12976 VDD.n3395 VDD.t1114 0.607167
R12977 VDD.n3395 VDD.n3394 0.607167
R12978 VDD.n3398 VDD.t1223 0.607167
R12979 VDD.n3398 VDD.n3397 0.607167
R12980 VDD.n5357 VDD.t1235 0.607167
R12981 VDD.n5357 VDD.n5356 0.607167
R12982 VDD.n5359 VDD.t1423 0.607167
R12983 VDD.n5359 VDD.n5358 0.607167
R12984 VDD.n3401 VDD.t1036 0.607167
R12985 VDD.n3401 VDD.n3400 0.607167
R12986 VDD.n3404 VDD.t1447 0.607167
R12987 VDD.n3404 VDD.n3403 0.607167
R12988 VDD.n5363 VDD.t608 0.607167
R12989 VDD.n5363 VDD.n5362 0.607167
R12990 VDD.n5365 VDD.t1241 0.607167
R12991 VDD.n5365 VDD.n5364 0.607167
R12992 VDD.n3407 VDD.t1139 0.607167
R12993 VDD.n3407 VDD.n3406 0.607167
R12994 VDD.n3410 VDD.t1349 0.607167
R12995 VDD.n3410 VDD.n3409 0.607167
R12996 VDD.n5369 VDD.t840 0.607167
R12997 VDD.n5369 VDD.n5368 0.607167
R12998 VDD.n5371 VDD.t1057 0.607167
R12999 VDD.n5371 VDD.n5370 0.607167
R13000 VDD.n3428 VDD.t1304 0.607167
R13001 VDD.n3428 VDD.n3427 0.607167
R13002 VDD.n3432 VDD.t827 0.607167
R13003 VDD.n3432 VDD.n3431 0.607167
R13004 VDD.n3417 VDD.t1321 0.607167
R13005 VDD.n3417 VDD.n3416 0.607167
R13006 VDD.n3419 VDD.t731 0.607167
R13007 VDD.n3419 VDD.n3418 0.607167
R13008 VDD.n3422 VDD.t1134 0.607167
R13009 VDD.n3422 VDD.n3421 0.607167
R13010 VDD.n3424 VDD.t725 0.607167
R13011 VDD.n3424 VDD.n3423 0.607167
R13012 VDD.n5374 VDD.t1054 0.607167
R13013 VDD.n5374 VDD.n5373 0.607167
R13014 VDD.n5376 VDD.t651 0.607167
R13015 VDD.n5376 VDD.n5375 0.607167
R13016 VDD.n5381 VDD.t766 0.607167
R13017 VDD.n5381 VDD.n5380 0.607167
R13018 VDD.n5383 VDD.t1157 0.607167
R13019 VDD.n5383 VDD.n5382 0.607167
R13020 VDD.n3435 VDD.t808 0.607167
R13021 VDD.n3435 VDD.n3434 0.607167
R13022 VDD.n3438 VDD.t1330 0.607167
R13023 VDD.n3438 VDD.n3437 0.607167
R13024 VDD.n5387 VDD.t1279 0.607167
R13025 VDD.n5387 VDD.n5386 0.607167
R13026 VDD.n5389 VDD.t1120 0.607167
R13027 VDD.n5389 VDD.n5388 0.607167
R13028 VDD.n3441 VDD.t1225 0.607167
R13029 VDD.n3441 VDD.n3440 0.607167
R13030 VDD.n3444 VDD.t1385 0.607167
R13031 VDD.n3444 VDD.n3443 0.607167
R13032 VDD.n5428 VDD.t1107 0.607167
R13033 VDD.n5428 VDD.n5427 0.607167
R13034 VDD.n5430 VDD.t706 0.607167
R13035 VDD.n5430 VDD.n5429 0.607167
R13036 VDD.n3709 VDD.t1284 0.607167
R13037 VDD.n3709 VDD.n3708 0.607167
R13038 VDD.n3712 VDD.t1129 0.607167
R13039 VDD.n3712 VDD.n3711 0.607167
R13040 VDD.n5434 VDD.t1038 0.607167
R13041 VDD.n5434 VDD.n5433 0.607167
R13042 VDD.n5436 VDD.t1166 0.607167
R13043 VDD.n5436 VDD.n5435 0.607167
R13044 VDD.n3715 VDD.t792 0.607167
R13045 VDD.n3715 VDD.n3714 0.607167
R13046 VDD.n3718 VDD.t1268 0.607167
R13047 VDD.n3718 VDD.n3717 0.607167
R13048 VDD.n5440 VDD.t743 0.607167
R13049 VDD.n5440 VDD.n5439 0.607167
R13050 VDD.n5442 VDD.t1073 0.607167
R13051 VDD.n5442 VDD.n5441 0.607167
R13052 VDD.n3732 VDD.t694 0.607167
R13053 VDD.n3732 VDD.n3731 0.607167
R13054 VDD.n3736 VDD.t903 0.607167
R13055 VDD.n3736 VDD.n3735 0.607167
R13056 VDD.n3723 VDD.t1444 0.607167
R13057 VDD.n3723 VDD.n3722 0.607167
R13058 VDD.n3721 VDD.t1252 0.607167
R13059 VDD.n3721 VDD.n3720 0.607167
R13060 VDD.n3728 VDD.t1267 0.607167
R13061 VDD.n3728 VDD.n3727 0.607167
R13062 VDD.n3726 VDD.t735 0.607167
R13063 VDD.n3726 VDD.n3725 0.607167
R13064 VDD.n5447 VDD.t1195 0.607167
R13065 VDD.n5447 VDD.n5446 0.607167
R13066 VDD.n5445 VDD.t1309 0.607167
R13067 VDD.n5445 VDD.n5444 0.607167
R13068 VDD.n5452 VDD.t1037 0.607167
R13069 VDD.n5452 VDD.n5451 0.607167
R13070 VDD.n5454 VDD.t1448 0.607167
R13071 VDD.n5454 VDD.n5453 0.607167
R13072 VDD.n3743 VDD.t926 0.607167
R13073 VDD.n3743 VDD.n3742 0.607167
R13074 VDD.n3746 VDD.t1211 0.607167
R13075 VDD.n3746 VDD.n3745 0.607167
R13076 VDD.n5458 VDD.t1369 0.607167
R13077 VDD.n5458 VDD.n5457 0.607167
R13078 VDD.n5460 VDD.t1181 0.607167
R13079 VDD.n5460 VDD.n5459 0.607167
R13080 VDD.n3749 VDD.t1017 0.607167
R13081 VDD.n3749 VDD.n3748 0.607167
R13082 VDD.n3752 VDD.t1172 0.607167
R13083 VDD.n3752 VDD.n3751 0.607167
R13084 VDD.n5464 VDD.t1305 0.607167
R13085 VDD.n5464 VDD.n5463 0.607167
R13086 VDD.n5466 VDD.t832 0.607167
R13087 VDD.n5466 VDD.n5465 0.607167
R13088 VDD.n3755 VDD.t1358 0.607167
R13089 VDD.n3755 VDD.n3754 0.607167
R13090 VDD.n3758 VDD.t1178 0.607167
R13091 VDD.n3758 VDD.n3757 0.607167
R13092 VDD.n6201 VDD.t843 0.607167
R13093 VDD.n6201 VDD.n6200 0.607167
R13094 VDD.n6203 VDD.t1063 0.607167
R13095 VDD.n6203 VDD.n6202 0.607167
R13096 VDD.n2906 VDD.t784 0.607167
R13097 VDD.n2906 VDD.n2905 0.607167
R13098 VDD.n2909 VDD.t809 0.607167
R13099 VDD.n2909 VDD.n2908 0.607167
R13100 VDD.n6195 VDD.t816 0.607167
R13101 VDD.n6195 VDD.n6194 0.607167
R13102 VDD.n6197 VDD.t1431 0.607167
R13103 VDD.n6197 VDD.n6196 0.607167
R13104 VDD.n2912 VDD.t1434 0.607167
R13105 VDD.n2912 VDD.n2911 0.607167
R13106 VDD.n2915 VDD.t918 0.607167
R13107 VDD.n2915 VDD.n2914 0.607167
R13108 VDD.n6189 VDD.t1025 0.607167
R13109 VDD.n6189 VDD.n6188 0.607167
R13110 VDD.n6191 VDD.t1439 0.607167
R13111 VDD.n6191 VDD.n6190 0.607167
R13112 VDD.n2918 VDD.t887 0.607167
R13113 VDD.n2918 VDD.n2917 0.607167
R13114 VDD.n2921 VDD.t667 0.607167
R13115 VDD.n2921 VDD.n2920 0.607167
R13116 VDD.n6177 VDD.t1406 0.607167
R13117 VDD.n6177 VDD.n6176 0.607167
R13118 VDD.n6179 VDD.t1224 0.607167
R13119 VDD.n6179 VDD.n6178 0.607167
R13120 VDD.n2939 VDD.t598 0.607167
R13121 VDD.n2939 VDD.n2938 0.607167
R13122 VDD.n2943 VDD.t1234 0.607167
R13123 VDD.n2943 VDD.n2942 0.607167
R13124 VDD.n2928 VDD.t1128 0.607167
R13125 VDD.n2928 VDD.n2927 0.607167
R13126 VDD.n2930 VDD.t645 0.607167
R13127 VDD.n2930 VDD.n2929 0.607167
R13128 VDD.n2933 VDD.t1355 0.607167
R13129 VDD.n2933 VDD.n2932 0.607167
R13130 VDD.n2935 VDD.t656 0.607167
R13131 VDD.n2935 VDD.n2934 0.607167
R13132 VDD.n6182 VDD.t1388 0.607167
R13133 VDD.n6182 VDD.n6181 0.607167
R13134 VDD.n6184 VDD.t1251 0.607167
R13135 VDD.n6184 VDD.n6183 0.607167
R13136 VDD.n6171 VDD.t679 0.607167
R13137 VDD.n6171 VDD.n6170 0.607167
R13138 VDD.n6173 VDD.t1383 0.607167
R13139 VDD.n6173 VDD.n6172 0.607167
R13140 VDD.n2946 VDD.t758 0.607167
R13141 VDD.n2946 VDD.n2945 0.607167
R13142 VDD.n2949 VDD.t1080 0.607167
R13143 VDD.n2949 VDD.n2948 0.607167
R13144 VDD.n6165 VDD.t1160 0.607167
R13145 VDD.n6165 VDD.n6164 0.607167
R13146 VDD.n6167 VDD.t1409 0.607167
R13147 VDD.n6167 VDD.n6166 0.607167
R13148 VDD.n2952 VDD.t1121 0.607167
R13149 VDD.n2952 VDD.n2951 0.607167
R13150 VDD.n2955 VDD.t1052 0.607167
R13151 VDD.n2955 VDD.n2954 0.607167
R13152 VDD.n5291 VDD.t1352 0.607167
R13153 VDD.n5291 VDD.n5290 0.607167
R13154 VDD.n5293 VDD.t807 0.607167
R13155 VDD.n5293 VDD.n5292 0.607167
R13156 VDD.n3205 VDD.t1324 0.607167
R13157 VDD.n3205 VDD.n3204 0.607167
R13158 VDD.n3208 VDD.t1364 0.607167
R13159 VDD.n3208 VDD.n3207 0.607167
R13160 VDD.n5297 VDD.t1058 0.607167
R13161 VDD.n5297 VDD.n5296 0.607167
R13162 VDD.n5299 VDD.t1140 0.607167
R13163 VDD.n5299 VDD.n5298 0.607167
R13164 VDD.n3211 VDD.t1375 0.607167
R13165 VDD.n3211 VDD.n3210 0.607167
R13166 VDD.n3214 VDD.t871 0.607167
R13167 VDD.n3214 VDD.n3213 0.607167
R13168 VDD.n5303 VDD.t1417 0.607167
R13169 VDD.n5303 VDD.n5302 0.607167
R13170 VDD.n5305 VDD.t839 0.607167
R13171 VDD.n5305 VDD.n5304 0.607167
R13172 VDD.n3228 VDD.t1149 0.607167
R13173 VDD.n3228 VDD.n3227 0.607167
R13174 VDD.n3232 VDD.t1403 0.607167
R13175 VDD.n3232 VDD.n3231 0.607167
R13176 VDD.n3219 VDD.t1060 0.607167
R13177 VDD.n3219 VDD.n3218 0.607167
R13178 VDD.n3217 VDD.t1310 0.607167
R13179 VDD.n3217 VDD.n3216 0.607167
R13180 VDD.n3224 VDD.t1124 0.607167
R13181 VDD.n3224 VDD.n3223 0.607167
R13182 VDD.n3222 VDD.t730 0.607167
R13183 VDD.n3222 VDD.n3221 0.607167
R13184 VDD.n5310 VDD.t1280 0.607167
R13185 VDD.n5310 VDD.n5309 0.607167
R13186 VDD.n5308 VDD.t1294 0.607167
R13187 VDD.n5308 VDD.n5307 0.607167
R13188 VDD.n5315 VDD.t1287 0.607167
R13189 VDD.n5315 VDD.n5314 0.607167
R13190 VDD.n5317 VDD.t1011 0.607167
R13191 VDD.n5317 VDD.n5316 0.607167
R13192 VDD.n3239 VDD.t635 0.607167
R13193 VDD.n3239 VDD.n3238 0.607167
R13194 VDD.n3242 VDD.t1165 0.607167
R13195 VDD.n3242 VDD.n3241 0.607167
R13196 VDD.n5321 VDD.t1222 0.607167
R13197 VDD.n5321 VDD.n5320 0.607167
R13198 VDD.n5323 VDD.t1288 0.607167
R13199 VDD.n5323 VDD.n5322 0.607167
R13200 VDD.n3245 VDD.t1045 0.607167
R13201 VDD.n3245 VDD.n3244 0.607167
R13202 VDD.n3248 VDD.t1148 0.607167
R13203 VDD.n3248 VDD.n3247 0.607167
R13204 VDD.n5327 VDD.t1171 0.607167
R13205 VDD.n5327 VDD.n5326 0.607167
R13206 VDD.n5329 VDD.t1113 0.607167
R13207 VDD.n5329 VDD.n5328 0.607167
R13208 VDD.n3251 VDD.t1095 0.607167
R13209 VDD.n3251 VDD.n3250 0.607167
R13210 VDD.n3254 VDD.t1306 0.607167
R13211 VDD.n3254 VDD.n3253 0.607167
R13212 VDD.n2538 VDD.t1019 0.607167
R13213 VDD.n2538 VDD.n2537 0.607167
R13214 VDD.n2540 VDD.t782 0.607167
R13215 VDD.n2540 VDD.n2539 0.607167
R13216 VDD.n2838 VDD.t1348 0.607167
R13217 VDD.n2838 VDD.n2837 0.607167
R13218 VDD.n2841 VDD.t793 0.607167
R13219 VDD.n2841 VDD.n2840 0.607167
R13220 VDD.n2544 VDD.t1015 0.607167
R13221 VDD.n2544 VDD.n2543 0.607167
R13222 VDD.n2546 VDD.t1173 0.607167
R13223 VDD.n2546 VDD.n2545 0.607167
R13224 VDD.n2844 VDD.t937 0.607167
R13225 VDD.n2844 VDD.n2843 0.607167
R13226 VDD.n2847 VDD.t702 0.607167
R13227 VDD.n2847 VDD.n2846 0.607167
R13228 VDD.n2550 VDD.t790 0.607167
R13229 VDD.n2550 VDD.n2549 0.607167
R13230 VDD.n2552 VDD.t1018 0.607167
R13231 VDD.n2552 VDD.n2551 0.607167
R13232 VDD.n2861 VDD.t1112 0.607167
R13233 VDD.n2861 VDD.n2860 0.607167
R13234 VDD.n2865 VDD.t711 0.607167
R13235 VDD.n2865 VDD.n2864 0.607167
R13236 VDD.n2852 VDD.t1329 0.607167
R13237 VDD.n2852 VDD.n2851 0.607167
R13238 VDD.n2850 VDD.t640 0.607167
R13239 VDD.n2850 VDD.n2849 0.607167
R13240 VDD.n2857 VDD.t1377 0.607167
R13241 VDD.n2857 VDD.n2856 0.607167
R13242 VDD.n2855 VDD.t724 0.607167
R13243 VDD.n2855 VDD.n2854 0.607167
R13244 VDD.n2557 VDD.t672 0.607167
R13245 VDD.n2557 VDD.n2556 0.607167
R13246 VDD.n2555 VDD.t649 0.607167
R13247 VDD.n2555 VDD.n2554 0.607167
R13248 VDD.n2562 VDD.t894 0.607167
R13249 VDD.n2562 VDD.n2561 0.607167
R13250 VDD.n2564 VDD.t681 0.607167
R13251 VDD.n2564 VDD.n2563 0.607167
R13252 VDD.n2872 VDD.t1161 0.607167
R13253 VDD.n2872 VDD.n2871 0.607167
R13254 VDD.n2875 VDD.t932 0.607167
R13255 VDD.n2875 VDD.n2874 0.607167
R13256 VDD.n2568 VDD.t1244 0.607167
R13257 VDD.n2568 VDD.n2567 0.607167
R13258 VDD.n2570 VDD.t1206 0.607167
R13259 VDD.n2570 VDD.n2569 0.607167
R13260 VDD.n2878 VDD.t1395 0.607167
R13261 VDD.n2878 VDD.n2877 0.607167
R13262 VDD.n2881 VDD.t1359 0.607167
R13263 VDD.n2881 VDD.n2880 0.607167
R13264 VDD.n2574 VDD.t805 0.607167
R13265 VDD.n2574 VDD.n2573 0.607167
R13266 VDD.n2576 VDD.t606 0.607167
R13267 VDD.n2576 VDD.n2575 0.607167
R13268 VDD.n2884 VDD.t1374 0.607167
R13269 VDD.n2884 VDD.n2883 0.607167
R13270 VDD.n2887 VDD.t869 0.607167
R13271 VDD.n2887 VDD.n2886 0.607167
R13272 VDD.n1355 VDD.t83 0.607167
R13273 VDD.n1355 VDD.n1354 0.607167
R13274 VDD.n1357 VDD.t81 0.607167
R13275 VDD.n1357 VDD.n1356 0.607167
R13276 VDD.n1359 VDD.t96 0.607167
R13277 VDD.n1359 VDD.n1358 0.607167
R13278 VDD.n1361 VDD.t105 0.607167
R13279 VDD.n1361 VDD.n1360 0.607167
R13280 VDD.n1366 VDD.t94 0.607167
R13281 VDD.n1366 VDD.n1365 0.607167
R13282 VDD.n1368 VDD.t552 0.607167
R13283 VDD.n1368 VDD.n1367 0.607167
R13284 VDD.n1370 VDD.t405 0.607167
R13285 VDD.n1370 VDD.n1369 0.607167
R13286 VDD.n1372 VDD.t542 0.607167
R13287 VDD.n1372 VDD.n1371 0.607167
R13288 VDD.n1377 VDD.t402 0.607167
R13289 VDD.n1377 VDD.n1376 0.607167
R13290 VDD.n1379 VDD.t400 0.607167
R13291 VDD.n1379 VDD.n1378 0.607167
R13292 VDD.n1381 VDD.t417 0.607167
R13293 VDD.n1381 VDD.n1380 0.607167
R13294 VDD.n1383 VDD.t122 0.607167
R13295 VDD.n1383 VDD.n1382 0.607167
R13296 VDD.n1388 VDD.t82 0.607167
R13297 VDD.n1388 VDD.n1387 0.607167
R13298 VDD.n1390 VDD.t79 0.607167
R13299 VDD.n1390 VDD.n1389 0.607167
R13300 VDD.n1392 VDD.t95 0.607167
R13301 VDD.n1392 VDD.n1391 0.607167
R13302 VDD.n1394 VDD.t104 0.607167
R13303 VDD.n1394 VDD.n1393 0.607167
R13304 VDD.n1399 VDD.t553 0.607167
R13305 VDD.n1399 VDD.n1398 0.607167
R13306 VDD.n1401 VDD.t551 0.607167
R13307 VDD.n1401 VDD.n1400 0.607167
R13308 VDD.n1403 VDD.t404 0.607167
R13309 VDD.n1403 VDD.n1402 0.607167
R13310 VDD.n1405 VDD.t541 0.607167
R13311 VDD.n1405 VDD.n1404 0.607167
R13312 VDD.n1410 VDD.t401 0.607167
R13313 VDD.n1410 VDD.n1409 0.607167
R13314 VDD.n1412 VDD.t399 0.607167
R13315 VDD.n1412 VDD.n1411 0.607167
R13316 VDD.n1414 VDD.t416 0.607167
R13317 VDD.n1414 VDD.n1413 0.607167
R13318 VDD.n1416 VDD.t427 0.607167
R13319 VDD.n1416 VDD.n1415 0.607167
R13320 VDD.n1118 VDD.t859 0.607167
R13321 VDD.n1118 VDD.n1117 0.607167
R13322 VDD.n1115 VDD.t525 0.607167
R13323 VDD.n1115 VDD.n1114 0.607167
R13324 VDD.n1429 VDD.t860 0.607167
R13325 VDD.n1429 VDD.n1428 0.607167
R13326 VDD.n1427 VDD.t861 0.607167
R13327 VDD.n1427 VDD.n1426 0.607167
R13328 VDD.n1112 VDD.t445 0.607167
R13329 VDD.n1112 VDD.n1111 0.607167
R13330 VDD.n1109 VDD.t451 0.607167
R13331 VDD.n1109 VDD.n1108 0.607167
R13332 VDD.n1423 VDD.t444 0.607167
R13333 VDD.n1423 VDD.n1422 0.607167
R13334 VDD.n1421 VDD.t429 0.607167
R13335 VDD.n1421 VDD.n1420 0.607167
R13336 VDD.n1106 VDD.t426 0.607167
R13337 VDD.n1350 VDD.t138 0.607167
R13338 VDD.n1103 VDD.t85 0.607167
R13339 VDD.n1349 VDD.t397 0.607167
R13340 VDD.n444 VDD.n393 0.597239
R13341 VDD.n439 VDD.n408 0.597239
R13342 VDD.n8021 VDD.n7980 0.597239
R13343 VDD.n8016 VDD.n8015 0.597239
R13344 VDD.n566 VDD.t964 0.58197
R13345 VDD.n566 VDD.n565 0.58197
R13346 VDD.n739 VDD.t980 0.58197
R13347 VDD.n739 VDD.n738 0.58197
R13348 VDD.n742 VDD.t975 0.58197
R13349 VDD.n742 VDD.n741 0.58197
R13350 VDD.n745 VDD.t969 0.58197
R13351 VDD.n745 VDD.n744 0.58197
R13352 VDD.n569 VDD.t996 0.58197
R13353 VDD.n569 VDD.n568 0.58197
R13354 VDD.n748 VDD.t952 0.58197
R13355 VDD.n748 VDD.n747 0.58197
R13356 VDD.n751 VDD.t997 0.58197
R13357 VDD.n751 VDD.n750 0.58197
R13358 VDD.n754 VDD.t988 0.58197
R13359 VDD.n754 VDD.n753 0.58197
R13360 VDD.n878 VDD.t947 0.58197
R13361 VDD.n878 VDD.n877 0.58197
R13362 VDD.n1048 VDD.t953 0.58197
R13363 VDD.n1048 VDD.n1047 0.58197
R13364 VDD.n1051 VDD.t998 0.58197
R13365 VDD.n1051 VDD.n1050 0.58197
R13366 VDD.n1054 VDD.t989 0.58197
R13367 VDD.n1054 VDD.n1053 0.58197
R13368 VDD.n875 VDD.t962 0.58197
R13369 VDD.n875 VDD.n874 0.58197
R13370 VDD.n1039 VDD.t983 0.58197
R13371 VDD.n1039 VDD.n1038 0.58197
R13372 VDD.n1042 VDD.t979 0.58197
R13373 VDD.n1042 VDD.n1041 0.58197
R13374 VDD.n1045 VDD.t976 0.58197
R13375 VDD.n1045 VDD.n1044 0.58197
R13376 VDD.n8164 VDD.t14 0.58197
R13377 VDD.n8164 VDD.n8163 0.58197
R13378 VDD.n8161 VDD.t466 0.58197
R13379 VDD.n8161 VDD.n8160 0.58197
R13380 VDD.n8158 VDD.t865 0.58197
R13381 VDD.n8158 VDD.n8157 0.58197
R13382 VDD.n8156 VDD.t8 0.58197
R13383 VDD.n8156 VDD.n8155 0.58197
R13384 VDD.n8153 VDD.t16 0.58197
R13385 VDD.n8153 VDD.n8152 0.58197
R13386 VDD.n8150 VDD.t527 0.58197
R13387 VDD.n8150 VDD.n8149 0.58197
R13388 VDD.n8147 VDD.t21 0.58197
R13389 VDD.n8147 VDD.n8146 0.58197
R13390 VDD.n8145 VDD.t852 0.58197
R13391 VDD.n8145 VDD.n8144 0.58197
R13392 VDD.n7902 VDD.t47 0.58197
R13393 VDD.n7902 VDD.n7901 0.58197
R13394 VDD.n7899 VDD.t20 0.58197
R13395 VDD.n7899 VDD.n7898 0.58197
R13396 VDD.n7896 VDD.t22 0.58197
R13397 VDD.n7896 VDD.n7895 0.58197
R13398 VDD.n7894 VDD.t10 0.58197
R13399 VDD.n7894 VDD.n7893 0.58197
R13400 VDD.n7891 VDD.t558 0.58197
R13401 VDD.n8317 VDD.t509 0.58197
R13402 VDD.n8317 VDD.t370 0.58197
R13403 VDD.n8318 VDD.t526 0.58197
R13404 VDD.n8318 VDD.t203 0.58197
R13405 VDD.n8319 VDD.t27 0.58197
R13406 VDD.n8319 VDD.t216 0.58197
R13407 VDD.n7059 VDD.n7058 0.58197
R13408 VDD.n5 VDD.t366 0.58197
R13409 VDD.n5 VDD.n4 0.58197
R13410 VDD.n3 VDD.t360 0.58197
R13411 VDD.n3 VDD.n2 0.58197
R13412 VDD.n1 VDD.t229 0.58197
R13413 VDD.n1 VDD.n0 0.58197
R13414 VDD.n1792 VDD.n1791 0.520296
R13415 VDD.n1795 VDD.n1794 0.520296
R13416 VDD.n5346 VDD.n5340 0.480464
R13417 VDD.n5483 VDD.n5477 0.480464
R13418 VDD.n6314 VDD.n6308 0.480464
R13419 VDD.n6308 VDD 0.473954
R13420 VDD.n399 VDD.t939 0.4555
R13421 VDD.n399 VDD.n398 0.4555
R13422 VDD.n397 VDD.t510 0.4555
R13423 VDD.n397 VDD.n396 0.4555
R13424 VDD.n395 VDD.n394 0.4555
R13425 VDD.n7965 VDD.t92 0.4555
R13426 VDD.n7965 VDD.n7964 0.4555
R13427 VDD.n7963 VDD.t531 0.4555
R13428 VDD.n7963 VDD.n7962 0.4555
R13429 VDD.n7961 VDD.t39 0.4555
R13430 VDD.n7961 VDD.n7960 0.4555
R13431 VDD.n7907 VDD.t508 0.4555
R13432 VDD.n7907 VDD.n7906 0.4555
R13433 VDD.n7909 VDD.t477 0.4555
R13434 VDD.n7909 VDD.n7908 0.4555
R13435 VDD.n7911 VDD.t465 0.4555
R13436 VDD.n7911 VDD.n7910 0.4555
R13437 VDD.n354 VDD.t472 0.4555
R13438 VDD.n354 VDD.n353 0.4555
R13439 VDD.n352 VDD.t120 0.4555
R13440 VDD.n352 VDD.n351 0.4555
R13441 VDD.n317 VDD.t283 0.4555
R13442 VDD.n314 VDD.t263 0.4555
R13443 VDD.n314 VDD.n313 0.4555
R13444 VDD.n5751 VDD.n5547 0.444312
R13445 VDD.n5952 VDD.n5401 0.444312
R13446 VDD.n6147 VDD.n5276 0.444312
R13447 VDD.n6307 VDD.n6306 0.444312
R13448 VDD.n5401 VDD.n5400 0.42125
R13449 VDD.n6603 VDD.n6602 0.411125
R13450 VDD.n6606 VDD.n6605 0.411125
R13451 VDD.n5547 VDD.n5546 0.411125
R13452 VDD.n5951 VDD.n5947 0.401
R13453 VDD.n6155 VDD.n6151 0.401
R13454 VDD.n5750 VDD.n5746 0.401
R13455 VDD.n5129 VDD.n5124 0.395938
R13456 VDD.n1791 VDD.n1790 0.386214
R13457 VDD.n1794 VDD.n1793 0.386214
R13458 VDD.n4827 VDD.n4822 0.385812
R13459 VDD.n4525 VDD.n4520 0.375687
R13460 VDD.n6621 VDD.n6620 0.354031
R13461 VDD.n337 VDD.n319 0.344848
R13462 VDD.n341 VDD.n316 0.344848
R13463 VDD.n330 VDD.n320 0.344848
R13464 VDD.n8139 VDD.n7958 0.340935
R13465 VDD.n8135 VDD.n7975 0.340935
R13466 VDD.n8128 VDD.n7979 0.340935
R13467 VDD.n7954 VDD.n7905 0.340935
R13468 VDD.n7442 VDD.t89 0.311155
R13469 VDD.n7523 VDD.t40 0.311155
R13470 VDD.n7922 VDD.t476 0.290355
R13471 VDD.n2313 VDD.n1792 0.279684
R13472 VDD.n2174 VDD.n1795 0.279684
R13473 VDD.n7215 VDD.t17 0.271356
R13474 VDD.n404 VDD.n403 0.266587
R13475 VDD.n7973 VDD.n7970 0.266587
R13476 VDD.n6609 VDD.n6608 0.257
R13477 VDD.n1638 VDD.n1454 0.239276
R13478 VDD.n1545 VDD.n1544 0.239276
R13479 VDD.n6621 VDD.n1096 0.222688
R13480 VDD.n6622 VDD.n870 0.222688
R13481 VDD.n6612 VDD.n6611 0.219875
R13482 VDD.n7003 VDD.n6857 0.203563
R13483 VDD.n6620 VDD.n2533 0.195969
R13484 VDD.n1473 VDD.n1456 0.195194
R13485 VDD.n1512 VDD.n1455 0.195194
R13486 VDD.n2125 VDD.n1928 0.195194
R13487 VDD.n2067 VDD.n1929 0.195194
R13488 VDD.n8 VDD.n7 0.190283
R13489 VDD.n7889 VDD.n7888 0.190283
R13490 VDD.n5575 VDD.n5574 0.157022
R13491 VDD.n4181 VDD.n4180 0.157022
R13492 VDD.n5541 VDD.n5540 0.157022
R13493 VDD.n3949 VDD.n3948 0.157022
R13494 VDD.n5491 VDD.n5490 0.157022
R13495 VDD.n3889 VDD.n3888 0.157022
R13496 VDD.n3449 VDD.n3447 0.157022
R13497 VDD.n5395 VDD.n5394 0.157022
R13498 VDD.n3703 VDD.n3701 0.157022
R13499 VDD.n5422 VDD.n5421 0.157022
R13500 VDD.n3763 VDD.n3761 0.157022
R13501 VDD.n5472 VDD.n5471 0.157022
R13502 VDD.n6041 VDD.n6040 0.157022
R13503 VDD.n3389 VDD.n3388 0.157022
R13504 VDD.n2960 VDD.n2958 0.157022
R13505 VDD.n6162 VDD.n6161 0.157022
R13506 VDD.n3199 VDD.n3197 0.157022
R13507 VDD.n5285 VDD.n5284 0.157022
R13508 VDD.n3259 VDD.n3257 0.157022
R13509 VDD.n5335 VDD.n5334 0.157022
R13510 VDD.n6218 VDD.n6217 0.157022
R13511 VDD.n2900 VDD.n2899 0.157022
R13512 VDD.n2892 VDD.n2890 0.157022
R13513 VDD.n2582 VDD.n2581 0.157022
R13514 VDD.n2669 VDD.n2668 0.157022
R13515 VDD.n2832 VDD.n2831 0.157022
R13516 VDD.n549 VDD.n548 0.157022
R13517 VDD.n557 VDD.n556 0.157022
R13518 VDD.n1032 VDD.n1029 0.157022
R13519 VDD.n6627 VDD.n6626 0.157022
R13520 VDD.n307 VDD.n306 0.157022
R13521 VDD.n6862 VDD.n6861 0.157022
R13522 VDD.n403 VDD.n402 0.157022
R13523 VDD.n402 VDD.n401 0.157022
R13524 VDD.n7970 VDD.n7969 0.157022
R13525 VDD.n7973 VDD.n7972 0.157022
R13526 VDD.n7905 VDD.n7904 0.157022
R13527 VDD.n319 VDD.n318 0.157022
R13528 VDD.n316 VDD.n315 0.157022
R13529 VDD.n1449 VDD.n1448 0.157022
R13530 VDD.n1127 VDD.n1126 0.157022
R13531 VDD.n1441 VDD.n1440 0.157022
R13532 VDD.n1347 VDD.n1346 0.157022
R13533 VDD.n1101 VDD.n1100 0.157022
R13534 VDD.n4241 VDD.n4239 0.157022
R13535 VDD.n5625 VDD.n5624 0.157022
R13536 VDD.n6857 VDD.n6856 0.149958
R13537 VDD.n6613 VDD.n6612 0.141125
R13538 VDD.n6614 VDD.n6613 0.141125
R13539 VDD.n6615 VDD.n6614 0.141125
R13540 VDD.n6616 VDD.n6615 0.141125
R13541 VDD.n6617 VDD.n6616 0.141125
R13542 VDD.n6618 VDD.n6617 0.141125
R13543 VDD.n6619 VDD.n6618 0.141125
R13544 VDD.n6620 VDD.n6619 0.141125
R13545 VDD.n6855 VDD.n6854 0.122562
R13546 VDD.n4530 VDD.n3954 0.122281
R13547 VDD.n6608 VDD.n6600 0.122281
R13548 VDD.n4520 VDD.n4082 0.122281
R13549 VDD.n7567 VDD.n7565 0.122
R13550 VDD.n7330 VDD.n7329 0.120875
R13551 VDD.n7820 VDD.n7819 0.120875
R13552 VDD.n7245 VDD.n7241 0.11075
R13553 VDD.n7248 VDD.n7245 0.11075
R13554 VDD.n7254 VDD.n7251 0.11075
R13555 VDD.n7256 VDD.n7254 0.11075
R13556 VDD.n7262 VDD.n7260 0.11075
R13557 VDD.n7264 VDD.n7262 0.11075
R13558 VDD.n7266 VDD.n7264 0.11075
R13559 VDD.n7268 VDD.n7266 0.11075
R13560 VDD.n7270 VDD.n7268 0.11075
R13561 VDD.n7275 VDD.n7273 0.11075
R13562 VDD.n7277 VDD.n7275 0.11075
R13563 VDD.n7825 VDD.n7823 0.11075
R13564 VDD.n7830 VDD.n7828 0.11075
R13565 VDD.n7833 VDD.n7830 0.11075
R13566 VDD.n7835 VDD.n7833 0.11075
R13567 VDD.n7838 VDD.n7835 0.11075
R13568 VDD.n7840 VDD.n7838 0.11075
R13569 VDD.n7846 VDD.n7844 0.11075
R13570 VDD.n7849 VDD.n7846 0.11075
R13571 VDD.n7329 VDD.n7327 0.11075
R13572 VDD.n7327 VDD.n7325 0.11075
R13573 VDD.n7325 VDD.n7323 0.11075
R13574 VDD.n7323 VDD.n7321 0.11075
R13575 VDD.n7321 VDD.n7319 0.11075
R13576 VDD.n7319 VDD.n7317 0.11075
R13577 VDD.n7317 VDD.n7315 0.11075
R13578 VDD.n7315 VDD.n7313 0.11075
R13579 VDD.n7313 VDD.n7311 0.11075
R13580 VDD.n7311 VDD.n7309 0.11075
R13581 VDD.n7309 VDD.n7307 0.11075
R13582 VDD.n7307 VDD.n7305 0.11075
R13583 VDD.n7305 VDD.n7303 0.11075
R13584 VDD.n7303 VDD.n7301 0.11075
R13585 VDD.n7301 VDD.n7299 0.11075
R13586 VDD.n7299 VDD.n7297 0.11075
R13587 VDD.n7297 VDD.n7295 0.11075
R13588 VDD.n7295 VDD.n7293 0.11075
R13589 VDD.n7293 VDD.n7291 0.11075
R13590 VDD.n7291 VDD.n7289 0.11075
R13591 VDD.n7289 VDD.n7287 0.11075
R13592 VDD.n7287 VDD.n7285 0.11075
R13593 VDD.n7285 VDD.n7283 0.11075
R13594 VDD.n7283 VDD.n7281 0.11075
R13595 VDD.n7541 VDD.n7539 0.11075
R13596 VDD.n7543 VDD.n7541 0.11075
R13597 VDD.n7545 VDD.n7543 0.11075
R13598 VDD.n7547 VDD.n7545 0.11075
R13599 VDD.n7549 VDD.n7547 0.11075
R13600 VDD.n7551 VDD.n7549 0.11075
R13601 VDD.n7553 VDD.n7551 0.11075
R13602 VDD.n7555 VDD.n7553 0.11075
R13603 VDD.n7557 VDD.n7555 0.11075
R13604 VDD.n7559 VDD.n7557 0.11075
R13605 VDD.n7561 VDD.n7559 0.11075
R13606 VDD.n7563 VDD.n7561 0.11075
R13607 VDD.n7388 VDD.n7386 0.11075
R13608 VDD.n7386 VDD.n7384 0.11075
R13609 VDD.n7381 VDD.n7379 0.11075
R13610 VDD.n7379 VDD.n7377 0.11075
R13611 VDD.n7377 VDD.n7375 0.11075
R13612 VDD.n7375 VDD.n7373 0.11075
R13613 VDD.n7373 VDD.n7371 0.11075
R13614 VDD.n7368 VDD.n7366 0.11075
R13615 VDD.n7366 VDD.n7364 0.11075
R13616 VDD.n7361 VDD.n7359 0.11075
R13617 VDD.n7359 VDD.n7357 0.11075
R13618 VDD.n7357 VDD.n7355 0.11075
R13619 VDD.n7355 VDD.n7353 0.11075
R13620 VDD.n7353 VDD.n7351 0.11075
R13621 VDD.n7348 VDD.n7346 0.11075
R13622 VDD.n7346 VDD.n7344 0.11075
R13623 VDD.n7344 VDD.n7342 0.11075
R13624 VDD.n7339 VDD.n7338 0.11075
R13625 VDD.n7338 VDD.n7337 0.11075
R13626 VDD.n7337 VDD.n7336 0.11075
R13627 VDD.n7336 VDD.n7335 0.11075
R13628 VDD.n7335 VDD.n7334 0.11075
R13629 VDD.n7332 VDD.n7331 0.11075
R13630 VDD.n7637 VDD.n7635 0.11075
R13631 VDD.n7635 VDD.n7632 0.11075
R13632 VDD.n7628 VDD.n7626 0.11075
R13633 VDD.n7626 VDD.n7623 0.11075
R13634 VDD.n7623 VDD.n7621 0.11075
R13635 VDD.n7621 VDD.n7618 0.11075
R13636 VDD.n7618 VDD.n7616 0.11075
R13637 VDD.n7612 VDD.n7610 0.11075
R13638 VDD.n7610 VDD.n7607 0.11075
R13639 VDD.n7604 VDD.n7602 0.11075
R13640 VDD.n7602 VDD.n7600 0.11075
R13641 VDD.n7600 VDD.n7598 0.11075
R13642 VDD.n7598 VDD.n7596 0.11075
R13643 VDD.n7596 VDD.n7594 0.11075
R13644 VDD.n7591 VDD.n7589 0.11075
R13645 VDD.n7589 VDD.n7587 0.11075
R13646 VDD.n7587 VDD.n7585 0.11075
R13647 VDD.n7582 VDD.n7580 0.11075
R13648 VDD.n7580 VDD.n7578 0.11075
R13649 VDD.n7578 VDD.n7576 0.11075
R13650 VDD.n7576 VDD.n7574 0.11075
R13651 VDD.n7574 VDD.n7572 0.11075
R13652 VDD.n7569 VDD.n7567 0.11075
R13653 VDD.n7819 VDD.n7816 0.11075
R13654 VDD.n7816 VDD.n7813 0.11075
R13655 VDD.n7813 VDD.n7810 0.11075
R13656 VDD.n7810 VDD.n7807 0.11075
R13657 VDD.n7807 VDD.n7804 0.11075
R13658 VDD.n7804 VDD.n7801 0.11075
R13659 VDD.n7801 VDD.n7799 0.11075
R13660 VDD.n7799 VDD.n7797 0.11075
R13661 VDD.n7797 VDD.n7795 0.11075
R13662 VDD.n7795 VDD.n7793 0.11075
R13663 VDD.n7793 VDD.n7791 0.11075
R13664 VDD.n7791 VDD.n7789 0.11075
R13665 VDD.n7789 VDD.n7787 0.11075
R13666 VDD.n7787 VDD.n7785 0.11075
R13667 VDD.n7785 VDD.n7783 0.11075
R13668 VDD.n7783 VDD.n7781 0.11075
R13669 VDD.n7781 VDD.n7779 0.11075
R13670 VDD.n7779 VDD.n7777 0.11075
R13671 VDD.n7775 VDD.n7773 0.11075
R13672 VDD.n7773 VDD.n7771 0.11075
R13673 VDD.n7771 VDD.n7769 0.11075
R13674 VDD.n7769 VDD.n7767 0.11075
R13675 VDD.n7767 VDD.n7765 0.11075
R13676 VDD.n7765 VDD.n7763 0.11075
R13677 VDD.n7763 VDD.n7761 0.11075
R13678 VDD.n7761 VDD.n7759 0.11075
R13679 VDD.n7759 VDD.n7757 0.11075
R13680 VDD.n7757 VDD.n7755 0.11075
R13681 VDD.n7755 VDD.n7753 0.11075
R13682 VDD.n7753 VDD.n7751 0.11075
R13683 VDD.n7751 VDD.n7749 0.11075
R13684 VDD.n7749 VDD.n7747 0.11075
R13685 VDD.n7747 VDD.n7745 0.11075
R13686 VDD.n7745 VDD.n7743 0.11075
R13687 VDD.n7743 VDD.n7741 0.11075
R13688 VDD.n7741 VDD.n7739 0.11075
R13689 VDD.n7739 VDD.n7737 0.11075
R13690 VDD.n7736 VDD.n7734 0.11075
R13691 VDD.n7731 VDD.n7729 0.11075
R13692 VDD.n7729 VDD.n7727 0.11075
R13693 VDD.n7727 VDD.n7725 0.11075
R13694 VDD.n7725 VDD.n7723 0.11075
R13695 VDD.n7723 VDD.n7721 0.11075
R13696 VDD.n7718 VDD.n7716 0.11075
R13697 VDD.n7716 VDD.n7714 0.11075
R13698 VDD.n7714 VDD.n7712 0.11075
R13699 VDD.n7709 VDD.n7707 0.11075
R13700 VDD.n7707 VDD.n7705 0.11075
R13701 VDD.n7705 VDD.n7703 0.11075
R13702 VDD.n7703 VDD.n7701 0.11075
R13703 VDD.n7701 VDD.n7699 0.11075
R13704 VDD.n7696 VDD.n7694 0.11075
R13705 VDD.n7694 VDD.n7692 0.11075
R13706 VDD.n7688 VDD.n7686 0.11075
R13707 VDD.n7686 VDD.n7683 0.11075
R13708 VDD.n7683 VDD.n7681 0.11075
R13709 VDD.n7681 VDD.n7678 0.11075
R13710 VDD.n7678 VDD.n7676 0.11075
R13711 VDD.n7672 VDD.n7670 0.11075
R13712 VDD.n7670 VDD.n7667 0.11075
R13713 VDD.n7667 VDD.n7665 0.11075
R13714 VDD.n6855 VDD.n6622 0.104958
R13715 VDD.n7826 VDD.n7825 0.10175
R13716 VDD.n7333 VDD.n7332 0.10175
R13717 VDD.n7570 VDD.n7569 0.10175
R13718 VDD.n7734 VDD.n7732 0.10175
R13719 VDD.n7841 VDD.n7840 0.100625
R13720 VDD.n7340 VDD.n7339 0.100625
R13721 VDD.n7607 VDD.n7605 0.09275
R13722 VDD.n7697 VDD.n7696 0.09275
R13723 VDD.n7583 VDD.n7582 0.08825
R13724 VDD.n7721 VDD.n7719 0.08825
R13725 VDD.n7251 VDD.n7249 0.082625
R13726 VDD.n7364 VDD.n7362 0.082625
R13727 VDD.n7351 VDD.n7349 0.07925
R13728 VDD.n7823 VDD.n7820 0.077
R13729 VDD.n7331 VDD.n7330 0.077
R13730 VDD.n7641 VDD.n7640 0.077
R13731 VDD.n7737 VDD.n7736 0.077
R13732 VDD.n6716 VDD.n6714 0.0760357
R13733 VDD.n6718 VDD.n6716 0.0760357
R13734 VDD.n6720 VDD.n6718 0.0760357
R13735 VDD.n6722 VDD.n6720 0.0760357
R13736 VDD.n6724 VDD.n6722 0.0760357
R13737 VDD.n6726 VDD.n6724 0.0760357
R13738 VDD.n6728 VDD.n6726 0.0760357
R13739 VDD.n6730 VDD.n6728 0.0760357
R13740 VDD.n6732 VDD.n6730 0.0760357
R13741 VDD.n6734 VDD.n6732 0.0760357
R13742 VDD.n6736 VDD.n6734 0.0760357
R13743 VDD.n6738 VDD.n6736 0.0760357
R13744 VDD.n6740 VDD.n6738 0.0760357
R13745 VDD.n6742 VDD.n6740 0.0760357
R13746 VDD.n6744 VDD.n6742 0.0760357
R13747 VDD.n6746 VDD.n6744 0.0760357
R13748 VDD.n6748 VDD.n6746 0.0760357
R13749 VDD.n6750 VDD.n6748 0.0760357
R13750 VDD.n6753 VDD.n6750 0.0760357
R13751 VDD.n6756 VDD.n6753 0.0760357
R13752 VDD.n6759 VDD.n6756 0.0760357
R13753 VDD.n6762 VDD.n6759 0.0760357
R13754 VDD.n6765 VDD.n6762 0.0760357
R13755 VDD.n6768 VDD.n6765 0.0760357
R13756 VDD.n6771 VDD.n6768 0.0760357
R13757 VDD.n6774 VDD.n6771 0.0760357
R13758 VDD.n6777 VDD.n6774 0.0760357
R13759 VDD.n6780 VDD.n6777 0.0760357
R13760 VDD.n6783 VDD.n6780 0.0760357
R13761 VDD.n6786 VDD.n6783 0.0760357
R13762 VDD.n6789 VDD.n6786 0.0760357
R13763 VDD.n6792 VDD.n6789 0.0760357
R13764 VDD.n6795 VDD.n6792 0.0760357
R13765 VDD.n6798 VDD.n6795 0.0760357
R13766 VDD.n6801 VDD.n6798 0.0760357
R13767 VDD.n6804 VDD.n6801 0.0760357
R13768 VDD.n6807 VDD.n6804 0.0760357
R13769 VDD.n6810 VDD.n6807 0.0760357
R13770 VDD.n6813 VDD.n6810 0.0760357
R13771 VDD.n6816 VDD.n6813 0.0760357
R13772 VDD.n6819 VDD.n6816 0.0760357
R13773 VDD.n6822 VDD.n6819 0.0760357
R13774 VDD.n6825 VDD.n6822 0.0760357
R13775 VDD.n6828 VDD.n6825 0.0760357
R13776 VDD.n6851 VDD.n6828 0.0760357
R13777 VDD.n604 VDD.n602 0.0760357
R13778 VDD.n606 VDD.n604 0.0760357
R13779 VDD.n608 VDD.n606 0.0760357
R13780 VDD.n610 VDD.n608 0.0760357
R13781 VDD.n612 VDD.n610 0.0760357
R13782 VDD.n614 VDD.n612 0.0760357
R13783 VDD.n616 VDD.n614 0.0760357
R13784 VDD.n618 VDD.n616 0.0760357
R13785 VDD.n620 VDD.n618 0.0760357
R13786 VDD.n622 VDD.n620 0.0760357
R13787 VDD.n624 VDD.n622 0.0760357
R13788 VDD.n626 VDD.n624 0.0760357
R13789 VDD.n628 VDD.n626 0.0760357
R13790 VDD.n630 VDD.n628 0.0760357
R13791 VDD.n632 VDD.n630 0.0760357
R13792 VDD.n634 VDD.n632 0.0760357
R13793 VDD.n636 VDD.n634 0.0760357
R13794 VDD.n638 VDD.n636 0.0760357
R13795 VDD.n640 VDD.n638 0.0760357
R13796 VDD.n643 VDD.n640 0.0760357
R13797 VDD.n646 VDD.n643 0.0760357
R13798 VDD.n649 VDD.n646 0.0760357
R13799 VDD.n652 VDD.n649 0.0760357
R13800 VDD.n655 VDD.n652 0.0760357
R13801 VDD.n658 VDD.n655 0.0760357
R13802 VDD.n661 VDD.n658 0.0760357
R13803 VDD.n664 VDD.n661 0.0760357
R13804 VDD.n667 VDD.n664 0.0760357
R13805 VDD.n670 VDD.n667 0.0760357
R13806 VDD.n673 VDD.n670 0.0760357
R13807 VDD.n676 VDD.n673 0.0760357
R13808 VDD.n679 VDD.n676 0.0760357
R13809 VDD.n682 VDD.n679 0.0760357
R13810 VDD.n685 VDD.n682 0.0760357
R13811 VDD.n688 VDD.n685 0.0760357
R13812 VDD.n691 VDD.n688 0.0760357
R13813 VDD.n694 VDD.n691 0.0760357
R13814 VDD.n697 VDD.n694 0.0760357
R13815 VDD.n700 VDD.n697 0.0760357
R13816 VDD.n703 VDD.n700 0.0760357
R13817 VDD.n706 VDD.n703 0.0760357
R13818 VDD.n709 VDD.n706 0.0760357
R13819 VDD.n712 VDD.n709 0.0760357
R13820 VDD.n714 VDD.n712 0.0760357
R13821 VDD.n737 VDD.n714 0.0760357
R13822 VDD.n912 VDD.n910 0.0760357
R13823 VDD.n914 VDD.n912 0.0760357
R13824 VDD.n916 VDD.n914 0.0760357
R13825 VDD.n918 VDD.n916 0.0760357
R13826 VDD.n920 VDD.n918 0.0760357
R13827 VDD.n922 VDD.n920 0.0760357
R13828 VDD.n924 VDD.n922 0.0760357
R13829 VDD.n926 VDD.n924 0.0760357
R13830 VDD.n928 VDD.n926 0.0760357
R13831 VDD.n930 VDD.n928 0.0760357
R13832 VDD.n932 VDD.n930 0.0760357
R13833 VDD.n934 VDD.n932 0.0760357
R13834 VDD.n936 VDD.n934 0.0760357
R13835 VDD.n938 VDD.n936 0.0760357
R13836 VDD.n940 VDD.n938 0.0760357
R13837 VDD.n942 VDD.n940 0.0760357
R13838 VDD.n944 VDD.n942 0.0760357
R13839 VDD.n946 VDD.n944 0.0760357
R13840 VDD.n948 VDD.n946 0.0760357
R13841 VDD.n950 VDD.n948 0.0760357
R13842 VDD.n952 VDD.n950 0.0760357
R13843 VDD.n954 VDD.n952 0.0760357
R13844 VDD.n956 VDD.n954 0.0760357
R13845 VDD.n958 VDD.n956 0.0760357
R13846 VDD.n960 VDD.n958 0.0760357
R13847 VDD.n962 VDD.n960 0.0760357
R13848 VDD.n964 VDD.n962 0.0760357
R13849 VDD.n966 VDD.n964 0.0760357
R13850 VDD.n968 VDD.n966 0.0760357
R13851 VDD.n971 VDD.n968 0.0760357
R13852 VDD.n973 VDD.n971 0.0760357
R13853 VDD.n976 VDD.n973 0.0760357
R13854 VDD.n978 VDD.n976 0.0760357
R13855 VDD.n981 VDD.n978 0.0760357
R13856 VDD.n983 VDD.n981 0.0760357
R13857 VDD.n986 VDD.n983 0.0760357
R13858 VDD.n988 VDD.n986 0.0760357
R13859 VDD.n991 VDD.n988 0.0760357
R13860 VDD.n993 VDD.n991 0.0760357
R13861 VDD.n996 VDD.n993 0.0760357
R13862 VDD.n998 VDD.n996 0.0760357
R13863 VDD.n1001 VDD.n998 0.0760357
R13864 VDD.n1003 VDD.n1001 0.0760357
R13865 VDD.n8285 VDD.n8283 0.0760357
R13866 VDD.n8283 VDD.n8280 0.0760357
R13867 VDD.n8280 VDD.n8278 0.0760357
R13868 VDD.n8278 VDD.n8275 0.0760357
R13869 VDD.n8275 VDD.n8273 0.0760357
R13870 VDD.n8273 VDD.n8270 0.0760357
R13871 VDD.n8270 VDD.n8268 0.0760357
R13872 VDD.n8268 VDD.n8265 0.0760357
R13873 VDD.n8265 VDD.n8263 0.0760357
R13874 VDD.n8263 VDD.n8260 0.0760357
R13875 VDD.n8260 VDD.n8258 0.0760357
R13876 VDD.n8258 VDD.n8255 0.0760357
R13877 VDD.n8255 VDD.n8253 0.0760357
R13878 VDD.n8250 VDD.n8247 0.0760357
R13879 VDD.n8247 VDD.n8245 0.0760357
R13880 VDD.n8245 VDD.n8243 0.0760357
R13881 VDD.n8243 VDD.n8241 0.0760357
R13882 VDD.n8241 VDD.n8239 0.0760357
R13883 VDD.n8239 VDD.n8237 0.0760357
R13884 VDD.n8237 VDD.n8235 0.0760357
R13885 VDD.n8235 VDD.n8233 0.0760357
R13886 VDD.n8233 VDD.n8231 0.0760357
R13887 VDD.n8231 VDD.n8229 0.0760357
R13888 VDD.n8229 VDD.n8227 0.0760357
R13889 VDD.n8227 VDD.n8225 0.0760357
R13890 VDD.n8225 VDD.n8223 0.0760357
R13891 VDD.n8223 VDD.n8221 0.0760357
R13892 VDD.n8221 VDD.n8219 0.0760357
R13893 VDD.n8219 VDD.n8217 0.0760357
R13894 VDD.n8217 VDD.n8215 0.0760357
R13895 VDD.n215 VDD.n213 0.0760357
R13896 VDD.n217 VDD.n215 0.0760357
R13897 VDD.n219 VDD.n217 0.0760357
R13898 VDD.n221 VDD.n219 0.0760357
R13899 VDD.n223 VDD.n221 0.0760357
R13900 VDD.n225 VDD.n223 0.0760357
R13901 VDD.n227 VDD.n225 0.0760357
R13902 VDD.n229 VDD.n227 0.0760357
R13903 VDD.n231 VDD.n229 0.0760357
R13904 VDD.n233 VDD.n231 0.0760357
R13905 VDD.n235 VDD.n233 0.0760357
R13906 VDD.n237 VDD.n235 0.0760357
R13907 VDD.n239 VDD.n237 0.0760357
R13908 VDD.n241 VDD.n239 0.0760357
R13909 VDD.n243 VDD.n241 0.0760357
R13910 VDD.n245 VDD.n243 0.0760357
R13911 VDD.n248 VDD.n245 0.0760357
R13912 VDD.n250 VDD.n248 0.0760357
R13913 VDD.n253 VDD.n250 0.0760357
R13914 VDD.n255 VDD.n253 0.0760357
R13915 VDD.n258 VDD.n255 0.0760357
R13916 VDD.n260 VDD.n258 0.0760357
R13917 VDD.n263 VDD.n260 0.0760357
R13918 VDD.n265 VDD.n263 0.0760357
R13919 VDD.n268 VDD.n265 0.0760357
R13920 VDD.n270 VDD.n268 0.0760357
R13921 VDD.n273 VDD.n270 0.0760357
R13922 VDD.n275 VDD.n273 0.0760357
R13923 VDD.n278 VDD.n275 0.0760357
R13924 VDD.n280 VDD.n278 0.0760357
R13925 VDD.n283 VDD.n280 0.0760357
R13926 VDD.n285 VDD.n283 0.0760357
R13927 VDD.n288 VDD.n285 0.0760357
R13928 VDD.n290 VDD.n288 0.0760357
R13929 VDD.n302 VDD.n290 0.0760357
R13930 VDD.n138 VDD.n136 0.0760357
R13931 VDD.n136 VDD.n133 0.0760357
R13932 VDD.n133 VDD.n130 0.0760357
R13933 VDD.n130 VDD.n127 0.0760357
R13934 VDD.n127 VDD.n124 0.0760357
R13935 VDD.n124 VDD.n121 0.0760357
R13936 VDD.n121 VDD.n118 0.0760357
R13937 VDD.n118 VDD.n115 0.0760357
R13938 VDD.n115 VDD.n112 0.0760357
R13939 VDD.n112 VDD.n109 0.0760357
R13940 VDD.n109 VDD.n106 0.0760357
R13941 VDD.n106 VDD.n103 0.0760357
R13942 VDD.n103 VDD.n100 0.0760357
R13943 VDD.n100 VDD.n97 0.0760357
R13944 VDD.n97 VDD.n94 0.0760357
R13945 VDD.n94 VDD.n91 0.0760357
R13946 VDD.n91 VDD.n88 0.0760357
R13947 VDD.n88 VDD.n85 0.0760357
R13948 VDD.n85 VDD.n82 0.0760357
R13949 VDD.n82 VDD.n79 0.0760357
R13950 VDD.n79 VDD.n76 0.0760357
R13951 VDD.n76 VDD.n73 0.0760357
R13952 VDD.n73 VDD.n70 0.0760357
R13953 VDD.n70 VDD.n68 0.0760357
R13954 VDD.n68 VDD.n66 0.0760357
R13955 VDD.n66 VDD.n64 0.0760357
R13956 VDD.n64 VDD.n62 0.0760357
R13957 VDD.n62 VDD.n60 0.0760357
R13958 VDD.n60 VDD.n58 0.0760357
R13959 VDD.n58 VDD.n56 0.0760357
R13960 VDD.n56 VDD.n54 0.0760357
R13961 VDD.n54 VDD.n52 0.0760357
R13962 VDD.n52 VDD.n50 0.0760357
R13963 VDD.n50 VDD.n48 0.0760357
R13964 VDD.n48 VDD.n46 0.0760357
R13965 VDD.n46 VDD.n44 0.0760357
R13966 VDD.n6871 VDD.n6869 0.0760357
R13967 VDD.n6873 VDD.n6871 0.0760357
R13968 VDD.n6875 VDD.n6873 0.0760357
R13969 VDD.n6877 VDD.n6875 0.0760357
R13970 VDD.n6879 VDD.n6877 0.0760357
R13971 VDD.n6881 VDD.n6879 0.0760357
R13972 VDD.n6883 VDD.n6881 0.0760357
R13973 VDD.n6885 VDD.n6883 0.0760357
R13974 VDD.n6887 VDD.n6885 0.0760357
R13975 VDD.n6890 VDD.n6887 0.0760357
R13976 VDD.n6893 VDD.n6890 0.0760357
R13977 VDD.n6896 VDD.n6893 0.0760357
R13978 VDD.n6899 VDD.n6896 0.0760357
R13979 VDD.n6902 VDD.n6899 0.0760357
R13980 VDD.n6905 VDD.n6902 0.0760357
R13981 VDD.n6908 VDD.n6905 0.0760357
R13982 VDD.n6911 VDD.n6908 0.0760357
R13983 VDD.n6914 VDD.n6911 0.0760357
R13984 VDD.n6917 VDD.n6914 0.0760357
R13985 VDD.n6920 VDD.n6917 0.0760357
R13986 VDD.n6923 VDD.n6920 0.0760357
R13987 VDD.n6926 VDD.n6923 0.0760357
R13988 VDD.n6929 VDD.n6926 0.0760357
R13989 VDD.n6932 VDD.n6929 0.0760357
R13990 VDD.n6935 VDD.n6932 0.0760357
R13991 VDD.n6938 VDD.n6935 0.0760357
R13992 VDD.n6941 VDD.n6938 0.0760357
R13993 VDD.n6944 VDD.n6941 0.0760357
R13994 VDD.n6947 VDD.n6944 0.0760357
R13995 VDD.n6950 VDD.n6947 0.0760357
R13996 VDD.n6953 VDD.n6950 0.0760357
R13997 VDD.n6956 VDD.n6953 0.0760357
R13998 VDD.n6959 VDD.n6956 0.0760357
R13999 VDD.n6962 VDD.n6959 0.0760357
R14000 VDD.n6965 VDD.n6962 0.0760357
R14001 VDD.n6979 VDD.n6965 0.0760357
R14002 VDD.n7165 VDD.n7163 0.0760357
R14003 VDD.n7163 VDD.n7160 0.0760357
R14004 VDD.n7160 VDD.n7158 0.0760357
R14005 VDD.n7158 VDD.n7155 0.0760357
R14006 VDD.n7155 VDD.n7153 0.0760357
R14007 VDD.n7153 VDD.n7150 0.0760357
R14008 VDD.n7150 VDD.n7148 0.0760357
R14009 VDD.n7148 VDD.n7145 0.0760357
R14010 VDD.n7145 VDD.n7143 0.0760357
R14011 VDD.n7143 VDD.n7140 0.0760357
R14012 VDD.n7140 VDD.n7138 0.0760357
R14013 VDD.n7138 VDD.n7135 0.0760357
R14014 VDD.n7135 VDD.n7133 0.0760357
R14015 VDD.n7133 VDD.n7130 0.0760357
R14016 VDD.n7130 VDD.n7128 0.0760357
R14017 VDD.n7128 VDD.n7125 0.0760357
R14018 VDD.n7125 VDD.n7123 0.0760357
R14019 VDD.n7123 VDD.n7121 0.0760357
R14020 VDD.n7121 VDD.n7119 0.0760357
R14021 VDD.n7119 VDD.n7117 0.0760357
R14022 VDD.n7117 VDD.n7115 0.0760357
R14023 VDD.n7115 VDD.n7113 0.0760357
R14024 VDD.n7113 VDD.n7111 0.0760357
R14025 VDD.n7111 VDD.n7109 0.0760357
R14026 VDD.n7109 VDD.n7107 0.0760357
R14027 VDD.n7107 VDD.n7105 0.0760357
R14028 VDD.n7105 VDD.n7103 0.0760357
R14029 VDD.n7103 VDD.n7101 0.0760357
R14030 VDD.n7101 VDD.n7099 0.0760357
R14031 VDD.n7099 VDD.n7097 0.0760357
R14032 VDD.n7097 VDD.n7095 0.0760357
R14033 VDD.n7095 VDD.n7093 0.0760357
R14034 VDD.n7093 VDD.n7091 0.0760357
R14035 VDD.n7091 VDD.n7089 0.0760357
R14036 VDD.n7089 VDD.n7087 0.0760357
R14037 VDD.n7087 VDD.n7085 0.0760357
R14038 VDD.n7613 VDD.n7612 0.075875
R14039 VDD.n7692 VDD.n7689 0.075875
R14040 VDD.n1006 VDD.n1003 0.0745948
R14041 VDD.n1008 VDD.n1006 0.073431
R14042 VDD.n7594 VDD.n7592 0.0725
R14043 VDD.n7710 VDD.n7709 0.0725
R14044 VDD.n7271 VDD.n7270 0.071375
R14045 VDD.n7382 VDD.n7381 0.071375
R14046 VDD.n7629 VDD.n7628 0.071375
R14047 VDD.n7676 VDD.n7673 0.071375
R14048 VDD.n7257 VDD.n7256 0.07025
R14049 VDD.n7369 VDD.n7368 0.07025
R14050 VDD.n8251 VDD.n8250 0.0696071
R14051 VDD.n7391 VDD.n7279 0.068
R14052 VDD.n7391 VDD.n7390 0.068
R14053 VDD.n7279 VDD.n7277 0.06575
R14054 VDD.n7565 VDD.n7563 0.06575
R14055 VDD.n7390 VDD.n7388 0.06575
R14056 VDD.n7640 VDD.n7637 0.06575
R14057 VDD.n7777 VDD 0.062375
R14058 VDD.n908 VDD.n907 0.053375
R14059 VDD.n907 VDD.n905 0.053375
R14060 VDD.n902 VDD.n900 0.053375
R14061 VDD.n897 VDD.n895 0.053375
R14062 VDD.n895 VDD.n893 0.053375
R14063 VDD.n890 VDD.n888 0.053375
R14064 VDD.n888 VDD.n886 0.053375
R14065 VDD.n883 VDD.n881 0.053375
R14066 VDD.n574 VDD.n572 0.053375
R14067 VDD.n579 VDD.n577 0.053375
R14068 VDD.n581 VDD.n579 0.053375
R14069 VDD.n586 VDD.n584 0.053375
R14070 VDD.n588 VDD.n586 0.053375
R14071 VDD.n593 VDD.n591 0.053375
R14072 VDD.n598 VDD.n596 0.053375
R14073 VDD.n600 VDD.n598 0.053375
R14074 VDD.n6656 VDD.n6654 0.053375
R14075 VDD.n6661 VDD.n6659 0.053375
R14076 VDD.n6663 VDD.n6661 0.053375
R14077 VDD.n6665 VDD.n6663 0.053375
R14078 VDD.n6667 VDD.n6665 0.053375
R14079 VDD.n6669 VDD.n6667 0.053375
R14080 VDD.n6671 VDD.n6669 0.053375
R14081 VDD.n6673 VDD.n6671 0.053375
R14082 VDD.n6675 VDD.n6673 0.053375
R14083 VDD.n6677 VDD.n6675 0.053375
R14084 VDD.n6679 VDD.n6677 0.053375
R14085 VDD.n6681 VDD.n6679 0.053375
R14086 VDD.n6683 VDD.n6681 0.053375
R14087 VDD.n6685 VDD.n6683 0.053375
R14088 VDD.n6687 VDD.n6685 0.053375
R14089 VDD.n6689 VDD.n6687 0.053375
R14090 VDD.n6691 VDD.n6689 0.053375
R14091 VDD.n6693 VDD.n6691 0.053375
R14092 VDD.n6695 VDD.n6693 0.053375
R14093 VDD.n6697 VDD.n6695 0.053375
R14094 VDD.n6699 VDD.n6697 0.053375
R14095 VDD.n6701 VDD.n6699 0.053375
R14096 VDD.n6707 VDD.n6705 0.053375
R14097 VDD.n6712 VDD.n6710 0.053375
R14098 VDD.n142 VDD.n139 0.053375
R14099 VDD.n149 VDD.n146 0.053375
R14100 VDD.n156 VDD.n153 0.053375
R14101 VDD.n159 VDD.n156 0.053375
R14102 VDD.n162 VDD.n159 0.053375
R14103 VDD.n165 VDD.n162 0.053375
R14104 VDD.n168 VDD.n165 0.053375
R14105 VDD.n171 VDD.n168 0.053375
R14106 VDD.n174 VDD.n171 0.053375
R14107 VDD.n177 VDD.n174 0.053375
R14108 VDD.n180 VDD.n177 0.053375
R14109 VDD.n183 VDD.n180 0.053375
R14110 VDD.n186 VDD.n183 0.053375
R14111 VDD.n189 VDD.n186 0.053375
R14112 VDD.n192 VDD.n189 0.053375
R14113 VDD.n195 VDD.n192 0.053375
R14114 VDD.n198 VDD.n195 0.053375
R14115 VDD.n205 VDD.n202 0.053375
R14116 VDD.n211 VDD.n209 0.053375
R14117 VDD.n7182 VDD.n7179 0.053375
R14118 VDD.n7185 VDD.n7182 0.053375
R14119 VDD.n7188 VDD.n7185 0.053375
R14120 VDD.n7195 VDD.n7192 0.053375
R14121 VDD.n7198 VDD.n7195 0.053375
R14122 VDD.n7205 VDD.n7202 0.053375
R14123 VDD.n7208 VDD.n7205 0.053375
R14124 VDD.n7211 VDD.n7208 0.053375
R14125 VDD.n7214 VDD.n7211 0.053375
R14126 VDD.n7217 VDD.n7214 0.053375
R14127 VDD.n7220 VDD.n7217 0.053375
R14128 VDD.n7223 VDD.n7220 0.053375
R14129 VDD.n7226 VDD.n7223 0.053375
R14130 VDD.n7229 VDD.n7226 0.053375
R14131 VDD VDD.n7229 0.053375
R14132 VDD VDD.n8345 0.053375
R14133 VDD.n8345 VDD.n8342 0.053375
R14134 VDD.n8342 VDD.n8339 0.053375
R14135 VDD.n8339 VDD.n8336 0.053375
R14136 VDD.n8336 VDD.n8333 0.053375
R14137 VDD.n8333 VDD.n8330 0.053375
R14138 VDD.n8330 VDD.n8327 0.053375
R14139 VDD.n8316 VDD.n8313 0.053375
R14140 VDD.n8309 VDD.n8306 0.053375
R14141 VDD.n8306 VDD.n8303 0.053375
R14142 VDD.n8303 VDD.n8300 0.053375
R14143 VDD.n8300 VDD.n8297 0.053375
R14144 VDD.n532 VDD.n530 0.053375
R14145 VDD.n530 VDD.n527 0.053375
R14146 VDD.n527 VDD.n525 0.053375
R14147 VDD.n525 VDD.n522 0.053375
R14148 VDD.n522 VDD.n520 0.053375
R14149 VDD.n520 VDD.n517 0.053375
R14150 VDD.n517 VDD.n515 0.053375
R14151 VDD.n515 VDD.n512 0.053375
R14152 VDD.n512 VDD.n510 0.053375
R14153 VDD.n510 VDD.n507 0.053375
R14154 VDD.n507 VDD.n505 0.053375
R14155 VDD.n505 VDD.n502 0.053375
R14156 VDD.n502 VDD.n500 0.053375
R14157 VDD.n500 VDD.n497 0.053375
R14158 VDD.n497 VDD.n495 0.053375
R14159 VDD.n495 VDD.n492 0.053375
R14160 VDD.n492 VDD.n490 0.053375
R14161 VDD.n490 VDD.n487 0.053375
R14162 VDD.n487 VDD.n485 0.053375
R14163 VDD.n485 VDD.n482 0.053375
R14164 VDD.n482 VDD.n480 0.053375
R14165 VDD.n480 VDD.n477 0.053375
R14166 VDD.n477 VDD.n475 0.053375
R14167 VDD.n475 VDD.n473 0.053375
R14168 VDD.n473 VDD.n471 0.053375
R14169 VDD.n471 VDD.n469 0.053375
R14170 VDD.n469 VDD.n467 0.053375
R14171 VDD.n467 VDD.n465 0.053375
R14172 VDD.n465 VDD.n463 0.053375
R14173 VDD.n463 VDD.n461 0.053375
R14174 VDD.n461 VDD.n459 0.053375
R14175 VDD.n459 VDD.n457 0.053375
R14176 VDD.n457 VDD.n455 0.053375
R14177 VDD.n8109 VDD.n8107 0.053375
R14178 VDD.n8107 VDD.n8104 0.053375
R14179 VDD.n8104 VDD.n8102 0.053375
R14180 VDD.n8102 VDD.n8099 0.053375
R14181 VDD.n8099 VDD.n8097 0.053375
R14182 VDD.n8097 VDD.n8094 0.053375
R14183 VDD.n8094 VDD.n8092 0.053375
R14184 VDD.n8092 VDD.n8089 0.053375
R14185 VDD.n8089 VDD.n8087 0.053375
R14186 VDD.n8087 VDD.n8084 0.053375
R14187 VDD.n8084 VDD.n8082 0.053375
R14188 VDD.n8082 VDD.n8079 0.053375
R14189 VDD.n8079 VDD.n8077 0.053375
R14190 VDD.n8077 VDD.n8074 0.053375
R14191 VDD.n8074 VDD.n8072 0.053375
R14192 VDD.n8072 VDD.n8069 0.053375
R14193 VDD.n8069 VDD.n8067 0.053375
R14194 VDD.n8067 VDD.n8064 0.053375
R14195 VDD.n8064 VDD.n8062 0.053375
R14196 VDD.n8062 VDD.n8059 0.053375
R14197 VDD.n8059 VDD.n8057 0.053375
R14198 VDD.n8057 VDD.n8054 0.053375
R14199 VDD.n8054 VDD.n8052 0.053375
R14200 VDD.n8052 VDD.n8050 0.053375
R14201 VDD.n8050 VDD.n8048 0.053375
R14202 VDD.n8048 VDD.n8046 0.053375
R14203 VDD.n8046 VDD.n8044 0.053375
R14204 VDD.n8044 VDD.n8042 0.053375
R14205 VDD.n8042 VDD.n8040 0.053375
R14206 VDD.n8040 VDD.n8038 0.053375
R14207 VDD.n8038 VDD.n8036 0.053375
R14208 VDD.n8036 VDD.n8034 0.053375
R14209 VDD.n8034 VDD.n8032 0.053375
R14210 VDD.n452 VDD.n450 0.053375
R14211 VDD.n450 VDD.n448 0.053375
R14212 VDD.n448 VDD.n446 0.053375
R14213 VDD.n443 VDD.n441 0.053375
R14214 VDD.n438 VDD.n436 0.053375
R14215 VDD.n436 VDD.n434 0.053375
R14216 VDD.n434 VDD.n432 0.053375
R14217 VDD.n432 VDD.n430 0.053375
R14218 VDD.n430 VDD.n428 0.053375
R14219 VDD.n428 VDD.n426 0.053375
R14220 VDD.n426 VDD.n424 0.053375
R14221 VDD.n424 VDD.n422 0.053375
R14222 VDD.n422 VDD.n420 0.053375
R14223 VDD.n420 VDD.n418 0.053375
R14224 VDD.n418 VDD.n416 0.053375
R14225 VDD.n416 VDD.n414 0.053375
R14226 VDD.n414 VDD.n412 0.053375
R14227 VDD.n412 VDD.n410 0.053375
R14228 VDD.n7984 VDD.n7982 0.053375
R14229 VDD.n7986 VDD.n7984 0.053375
R14230 VDD.n7988 VDD.n7986 0.053375
R14231 VDD.n7990 VDD.n7988 0.053375
R14232 VDD.n7992 VDD.n7990 0.053375
R14233 VDD.n7994 VDD.n7992 0.053375
R14234 VDD.n7996 VDD.n7994 0.053375
R14235 VDD.n7998 VDD.n7996 0.053375
R14236 VDD.n8000 VDD.n7998 0.053375
R14237 VDD.n8002 VDD.n8000 0.053375
R14238 VDD.n8004 VDD.n8002 0.053375
R14239 VDD.n8006 VDD.n8004 0.053375
R14240 VDD.n8008 VDD.n8006 0.053375
R14241 VDD.n8010 VDD.n8008 0.053375
R14242 VDD.n8012 VDD.n8010 0.053375
R14243 VDD.n8014 VDD.n8012 0.053375
R14244 VDD.n8020 VDD.n8018 0.053375
R14245 VDD.n8025 VDD.n8023 0.053375
R14246 VDD.n8027 VDD.n8025 0.053375
R14247 VDD.n8029 VDD.n8027 0.053375
R14248 VDD.n544 VDD.n543 0.053375
R14249 VDD.n326 VDD.n323 0.053375
R14250 VDD.n329 VDD.n326 0.053375
R14251 VDD.n336 VDD.n333 0.053375
R14252 VDD.n347 VDD.n344 0.053375
R14253 VDD.n350 VDD.n347 0.053375
R14254 VDD.n389 VDD.n386 0.053375
R14255 VDD.n382 VDD.n379 0.053375
R14256 VDD.n379 VDD.n376 0.053375
R14257 VDD.n376 VDD.n373 0.053375
R14258 VDD.n369 VDD.n366 0.053375
R14259 VDD.n366 VDD.n363 0.053375
R14260 VDD.n363 VDD.n360 0.053375
R14261 VDD.n360 VDD.n357 0.053375
R14262 VDD.n7918 VDD.n7915 0.053375
R14263 VDD.n7921 VDD.n7918 0.053375
R14264 VDD.n7924 VDD.n7921 0.053375
R14265 VDD.n7927 VDD.n7924 0.053375
R14266 VDD.n7934 VDD.n7931 0.053375
R14267 VDD.n7937 VDD.n7934 0.053375
R14268 VDD.n7940 VDD.n7937 0.053375
R14269 VDD.n7947 VDD.n7944 0.053375
R14270 VDD.n7950 VDD.n7947 0.053375
R14271 VDD.n7953 VDD.n7950 0.053375
R14272 VDD.n8134 VDD.n8131 0.053375
R14273 VDD.n8127 VDD.n8124 0.053375
R14274 VDD.n8124 VDD.n8121 0.053375
R14275 VDD.n8121 VDD.n8118 0.053375
R14276 VDD.n6992 VDD.n6989 0.053375
R14277 VDD.n6999 VDD.n6996 0.053375
R14278 VDD.n7002 VDD.n6999 0.053375
R14279 VDD.n7009 VDD.n7006 0.053375
R14280 VDD.n7012 VDD.n7009 0.053375
R14281 VDD.n7015 VDD.n7012 0.053375
R14282 VDD.n7018 VDD.n7015 0.053375
R14283 VDD.n7022 VDD.n7018 0.053375
R14284 VDD.n7025 VDD.n7022 0.053375
R14285 VDD.n7028 VDD.n7025 0.053375
R14286 VDD.n7031 VDD.n7028 0.053375
R14287 VDD.n7034 VDD.n7031 0.053375
R14288 VDD.n7037 VDD.n7034 0.053375
R14289 VDD.n7044 VDD.n7041 0.053375
R14290 VDD.n7051 VDD.n7048 0.053375
R14291 VDD.n7083 VDD.n7055 0.053375
R14292 VDD.n7083 VDD.n7082 0.053375
R14293 VDD.n7082 VDD.n7080 0.053375
R14294 VDD.n7080 VDD.n7078 0.053375
R14295 VDD.n7075 VDD.n7073 0.053375
R14296 VDD.n7073 VDD.n7071 0.053375
R14297 VDD.n7068 VDD.n7066 0.053375
R14298 VDD.n7066 VDD.n7064 0.053375
R14299 VDD.n7064 VDD.n7062 0.053375
R14300 VDD.n8170 VDD.n8168 0.053375
R14301 VDD.n8172 VDD.n8170 0.053375
R14302 VDD.n8174 VDD.n8172 0.053375
R14303 VDD.n8176 VDD.n8174 0.053375
R14304 VDD.n8181 VDD.n8179 0.053375
R14305 VDD.n8183 VDD.n8181 0.053375
R14306 VDD.n8188 VDD.n8186 0.053375
R14307 VDD.n8193 VDD.n8191 0.053375
R14308 VDD.n8195 VDD.n8193 0.053375
R14309 VDD.n8197 VDD.n8195 0.053375
R14310 VDD.n8202 VDD.n8200 0.053375
R14311 VDD.n8207 VDD.n8205 0.053375
R14312 VDD.n8209 VDD.n8207 0.053375
R14313 VDD.n8211 VDD.n8209 0.053375
R14314 VDD.n8213 VDD.n8211 0.053375
R14315 VDD.n1095 VDD.n1092 0.053375
R14316 VDD.n1088 VDD.n1085 0.053375
R14317 VDD.n1081 VDD.n1078 0.053375
R14318 VDD.n1078 VDD.n1075 0.053375
R14319 VDD.n1071 VDD.n1068 0.053375
R14320 VDD.n1068 VDD.n1065 0.053375
R14321 VDD.n1061 VDD.n1058 0.053375
R14322 VDD.n761 VDD.n758 0.053375
R14323 VDD.n768 VDD.n765 0.053375
R14324 VDD.n771 VDD.n768 0.053375
R14325 VDD.n778 VDD.n775 0.053375
R14326 VDD.n781 VDD.n778 0.053375
R14327 VDD.n784 VDD.n781 0.053375
R14328 VDD.n787 VDD.n784 0.053375
R14329 VDD.n790 VDD.n787 0.053375
R14330 VDD.n793 VDD.n790 0.053375
R14331 VDD.n795 VDD.n793 0.053375
R14332 VDD.n798 VDD.n795 0.053375
R14333 VDD.n805 VDD.n802 0.053375
R14334 VDD.n812 VDD.n809 0.053375
R14335 VDD.n815 VDD.n812 0.053375
R14336 VDD.n818 VDD.n815 0.053375
R14337 VDD.n821 VDD.n818 0.053375
R14338 VDD.n824 VDD.n821 0.053375
R14339 VDD.n827 VDD.n824 0.053375
R14340 VDD.n830 VDD.n827 0.053375
R14341 VDD.n833 VDD.n830 0.053375
R14342 VDD.n836 VDD.n833 0.053375
R14343 VDD.n839 VDD.n836 0.053375
R14344 VDD.n842 VDD.n839 0.053375
R14345 VDD.n845 VDD.n842 0.053375
R14346 VDD.n848 VDD.n845 0.053375
R14347 VDD.n851 VDD.n848 0.053375
R14348 VDD.n854 VDD.n851 0.053375
R14349 VDD.n857 VDD.n854 0.053375
R14350 VDD.n860 VDD.n857 0.053375
R14351 VDD.n863 VDD.n860 0.053375
R14352 VDD.n866 VDD.n863 0.053375
R14353 VDD.n869 VDD.n866 0.053375
R14354 VDD.n6642 VDD.n6639 0.053375
R14355 VDD.n8143 VDD.n8142 0.0528125
R14356 VDD.n7189 VDD.n7188 0.0516875
R14357 VDD.n7078 VDD.n7076 0.0516875
R14358 VDD.n8313 VDD.n8310 0.0505625
R14359 VDD.n340 VDD.n337 0.0505625
R14360 VDD.n373 VDD.n370 0.0505625
R14361 VDD.n8191 VDD.n8189 0.0505625
R14362 VDD.n8203 VDD.n8202 0.0505625
R14363 VDD VDD.n7775 0.048875
R14364 VDD.n6652 VDD.n6651 0.0483125
R14365 VDD.n6710 VDD.n6708 0.0483125
R14366 VDD.n8139 VDD.n8138 0.0483125
R14367 VDD.n799 VDD.n798 0.0483125
R14368 VDD.n6646 VDD.n6643 0.0483125
R14369 VDD.n7931 VDD.n7928 0.0460625
R14370 VDD.n446 VDD.n444 0.0449375
R14371 VDD.n8023 VDD.n8021 0.0449375
R14372 VDD.n8128 VDD.n8127 0.0449375
R14373 VDD.n886 VDD.n884 0.0426875
R14374 VDD.n577 VDD.n575 0.0426875
R14375 VDD.n1065 VDD.n1062 0.0426875
R14376 VDD.n765 VDD.n762 0.0426875
R14377 VDD.n1096 VDD.n1095 0.042125
R14378 VDD.n7260 VDD.n7257 0.041
R14379 VDD.n7371 VDD.n7369 0.041
R14380 VDD.n8184 VDD.n8183 0.041
R14381 VDD.n341 VDD.n340 0.0404375
R14382 VDD.n7003 VDD.n7002 0.0404375
R14383 VDD.n7273 VDD.n7271 0.039875
R14384 VDD.n7384 VDD.n7382 0.039875
R14385 VDD.n7632 VDD.n7629 0.039875
R14386 VDD.n7673 VDD.n7672 0.039875
R14387 VDD.n6985 VDD.n6982 0.039875
R14388 VDD.n6854 VDD.n6646 0.039875
R14389 VDD.n7202 VDD.n7199 0.0393125
R14390 VDD.n7941 VDD.n7940 0.0393125
R14391 VDD.n7069 VDD.n7068 0.0393125
R14392 VDD.n7592 VDD.n7591 0.03875
R14393 VDD.n7712 VDD.n7710 0.03875
R14394 VDD.n7041 VDD.n7038 0.03875
R14395 VDD.n7397 VDD.n7394 0.0369463
R14396 VDD.n7400 VDD.n7397 0.0369463
R14397 VDD.n7403 VDD.n7400 0.0369463
R14398 VDD.n7406 VDD.n7403 0.0369463
R14399 VDD.n7409 VDD.n7406 0.0369463
R14400 VDD.n7413 VDD.n7409 0.0369463
R14401 VDD.n7417 VDD.n7413 0.0369463
R14402 VDD.n7421 VDD.n7417 0.0369463
R14403 VDD.n7425 VDD.n7421 0.0369463
R14404 VDD.n7429 VDD.n7425 0.0369463
R14405 VDD.n7433 VDD.n7429 0.0369463
R14406 VDD.n7437 VDD.n7433 0.0369463
R14407 VDD.n7441 VDD.n7437 0.0369463
R14408 VDD.n7445 VDD.n7441 0.0369463
R14409 VDD.n7449 VDD.n7445 0.0369463
R14410 VDD.n7453 VDD.n7449 0.0369463
R14411 VDD.n7457 VDD.n7453 0.0369463
R14412 VDD.n7461 VDD.n7457 0.0369463
R14413 VDD.n7465 VDD.n7461 0.0369463
R14414 VDD.n7469 VDD.n7465 0.0369463
R14415 VDD.n7473 VDD.n7469 0.0369463
R14416 VDD.n7477 VDD.n7473 0.0369463
R14417 VDD.n7481 VDD.n7477 0.0369463
R14418 VDD.n7485 VDD.n7481 0.0369463
R14419 VDD.n7489 VDD.n7485 0.0369463
R14420 VDD.n7493 VDD.n7489 0.0369463
R14421 VDD.n7497 VDD.n7493 0.0369463
R14422 VDD.n7501 VDD.n7497 0.0369463
R14423 VDD.n7505 VDD.n7501 0.0369463
R14424 VDD.n7509 VDD.n7505 0.0369463
R14425 VDD.n7513 VDD.n7509 0.0369463
R14426 VDD.n7517 VDD.n7513 0.0369463
R14427 VDD.n7521 VDD.n7517 0.0369463
R14428 VDD.n7525 VDD.n7521 0.0369463
R14429 VDD.n7529 VDD.n7525 0.0369463
R14430 VDD.n7533 VDD.n7529 0.0369463
R14431 VDD.n7537 VDD.n7533 0.0369463
R14432 VDD.n7886 VDD.n7241 0.0365
R14433 VDD.n898 VDD.n897 0.0359375
R14434 VDD.n589 VDD.n588 0.0359375
R14435 VDD.n153 VDD.n150 0.0359375
R14436 VDD.n199 VDD.n198 0.0359375
R14437 VDD.n6996 VDD.n6993 0.0359375
R14438 VDD.n7045 VDD.n7044 0.0359375
R14439 VDD.n1082 VDD.n1081 0.0359375
R14440 VDD.n7616 VDD.n7613 0.035375
R14441 VDD.n7689 VDD.n7688 0.035375
R14442 VDD.n8327 VDD.n8324 0.0348125
R14443 VDD.n333 VDD.n330 0.0348125
R14444 VDD.n383 VDD.n382 0.0348125
R14445 VDD.n8198 VDD.n8197 0.0348125
R14446 VDD.n905 VDD.n903 0.0336875
R14447 VDD.n596 VDD.n594 0.0336875
R14448 VDD.n143 VDD.n142 0.0336875
R14449 VDD.n209 VDD.n206 0.0336875
R14450 VDD.n6986 VDD.n6985 0.0336875
R14451 VDD.n7055 VDD.n7052 0.0336875
R14452 VDD.n1092 VDD.n1089 0.0336875
R14453 VDD.n891 VDD.n890 0.0325625
R14454 VDD.n582 VDD.n581 0.0325625
R14455 VDD.n6657 VDD.n6656 0.0325625
R14456 VDD.n6705 VDD.n6703 0.0325625
R14457 VDD.n7957 VDD.n7954 0.0325625
R14458 VDD.n1072 VDD.n1071 0.0325625
R14459 VDD.n772 VDD.n771 0.0325625
R14460 VDD.n806 VDD.n805 0.0325625
R14461 VDD.n6639 VDD.n6636 0.0325625
R14462 VDD.n7349 VDD.n7348 0.032
R14463 VDD.n7665 VDD.n7641 0.032
R14464 VDD.n441 VDD.n439 0.0291875
R14465 VDD.n8018 VDD.n8016 0.0291875
R14466 VDD.n8135 VDD.n8134 0.0291875
R14467 VDD.n8179 VDD.n8177 0.0291875
R14468 VDD.n7249 VDD.n7248 0.028625
R14469 VDD.n7362 VDD.n7361 0.028625
R14470 VDD.n390 VDD.n350 0.0280625
R14471 VDD.n5641 VDD.n5639 0.0269375
R14472 VDD.n5639 VDD.n5636 0.0269375
R14473 VDD.n5636 VDD.n5634 0.0269375
R14474 VDD.n5634 VDD.n5631 0.0269375
R14475 VDD.n4247 VDD.n4244 0.0269375
R14476 VDD.n4249 VDD.n4247 0.0269375
R14477 VDD.n4252 VDD.n4249 0.0269375
R14478 VDD.n4254 VDD.n4252 0.0269375
R14479 VDD.n4257 VDD.n4254 0.0269375
R14480 VDD.n4259 VDD.n4257 0.0269375
R14481 VDD.n4262 VDD.n4259 0.0269375
R14482 VDD.n4264 VDD.n4262 0.0269375
R14483 VDD.n4267 VDD.n4264 0.0269375
R14484 VDD.n4269 VDD.n4267 0.0269375
R14485 VDD.n4272 VDD.n4269 0.0269375
R14486 VDD.n4274 VDD.n4272 0.0269375
R14487 VDD.n4277 VDD.n4274 0.0269375
R14488 VDD.n4279 VDD.n4277 0.0269375
R14489 VDD.n4282 VDD.n4279 0.0269375
R14490 VDD.n4284 VDD.n4282 0.0269375
R14491 VDD.n4287 VDD.n4284 0.0269375
R14492 VDD.n4289 VDD.n4287 0.0269375
R14493 VDD.n4292 VDD.n4289 0.0269375
R14494 VDD.n4294 VDD.n4292 0.0269375
R14495 VDD.n4297 VDD.n4294 0.0269375
R14496 VDD.n4299 VDD.n4297 0.0269375
R14497 VDD.n4302 VDD.n4299 0.0269375
R14498 VDD.n4304 VDD.n4302 0.0269375
R14499 VDD.n4307 VDD.n4304 0.0269375
R14500 VDD.n4309 VDD.n4307 0.0269375
R14501 VDD.n4312 VDD.n4309 0.0269375
R14502 VDD.n4314 VDD.n4312 0.0269375
R14503 VDD.n4317 VDD.n4314 0.0269375
R14504 VDD.n4319 VDD.n4317 0.0269375
R14505 VDD.n4322 VDD.n4319 0.0269375
R14506 VDD.n4324 VDD.n4322 0.0269375
R14507 VDD.n4327 VDD.n4324 0.0269375
R14508 VDD.n4329 VDD.n4327 0.0269375
R14509 VDD.n4332 VDD.n4329 0.0269375
R14510 VDD.n4334 VDD.n4332 0.0269375
R14511 VDD.n4337 VDD.n4334 0.0269375
R14512 VDD.n4339 VDD.n4337 0.0269375
R14513 VDD.n4342 VDD.n4339 0.0269375
R14514 VDD.n4345 VDD.n4342 0.0269375
R14515 VDD.n4347 VDD.n4345 0.0269375
R14516 VDD.n4350 VDD.n4347 0.0269375
R14517 VDD.n5571 VDD.n5569 0.0269375
R14518 VDD.n5569 VDD.n5567 0.0269375
R14519 VDD.n5567 VDD.n5565 0.0269375
R14520 VDD.n5565 VDD.n5563 0.0269375
R14521 VDD.n4086 VDD.n4084 0.0269375
R14522 VDD.n4088 VDD.n4086 0.0269375
R14523 VDD.n4090 VDD.n4088 0.0269375
R14524 VDD.n4092 VDD.n4090 0.0269375
R14525 VDD.n4094 VDD.n4092 0.0269375
R14526 VDD.n4096 VDD.n4094 0.0269375
R14527 VDD.n4098 VDD.n4096 0.0269375
R14528 VDD.n4100 VDD.n4098 0.0269375
R14529 VDD.n4102 VDD.n4100 0.0269375
R14530 VDD.n4104 VDD.n4102 0.0269375
R14531 VDD.n4106 VDD.n4104 0.0269375
R14532 VDD.n4108 VDD.n4106 0.0269375
R14533 VDD.n4110 VDD.n4108 0.0269375
R14534 VDD.n4112 VDD.n4110 0.0269375
R14535 VDD.n4114 VDD.n4112 0.0269375
R14536 VDD.n4116 VDD.n4114 0.0269375
R14537 VDD.n4118 VDD.n4116 0.0269375
R14538 VDD.n4120 VDD.n4118 0.0269375
R14539 VDD.n4122 VDD.n4120 0.0269375
R14540 VDD.n4124 VDD.n4122 0.0269375
R14541 VDD.n4126 VDD.n4124 0.0269375
R14542 VDD.n4128 VDD.n4126 0.0269375
R14543 VDD.n4130 VDD.n4128 0.0269375
R14544 VDD.n4132 VDD.n4130 0.0269375
R14545 VDD.n4135 VDD.n4132 0.0269375
R14546 VDD.n4137 VDD.n4135 0.0269375
R14547 VDD.n4140 VDD.n4137 0.0269375
R14548 VDD.n4142 VDD.n4140 0.0269375
R14549 VDD.n4145 VDD.n4142 0.0269375
R14550 VDD.n4147 VDD.n4145 0.0269375
R14551 VDD.n4150 VDD.n4147 0.0269375
R14552 VDD.n4152 VDD.n4150 0.0269375
R14553 VDD.n4155 VDD.n4152 0.0269375
R14554 VDD.n4157 VDD.n4155 0.0269375
R14555 VDD.n4160 VDD.n4157 0.0269375
R14556 VDD.n4162 VDD.n4160 0.0269375
R14557 VDD.n4165 VDD.n4162 0.0269375
R14558 VDD.n4167 VDD.n4165 0.0269375
R14559 VDD.n4170 VDD.n4167 0.0269375
R14560 VDD.n4172 VDD.n4170 0.0269375
R14561 VDD.n4175 VDD.n4172 0.0269375
R14562 VDD.n4177 VDD.n4175 0.0269375
R14563 VDD.n5410 VDD.n5407 0.0269375
R14564 VDD.n5407 VDD.n5404 0.0269375
R14565 VDD.n3458 VDD.n3455 0.0269375
R14566 VDD.n3461 VDD.n3458 0.0269375
R14567 VDD.n3464 VDD.n3461 0.0269375
R14568 VDD.n3467 VDD.n3464 0.0269375
R14569 VDD.n3470 VDD.n3467 0.0269375
R14570 VDD.n3473 VDD.n3470 0.0269375
R14571 VDD.n3476 VDD.n3473 0.0269375
R14572 VDD.n3479 VDD.n3476 0.0269375
R14573 VDD.n3482 VDD.n3479 0.0269375
R14574 VDD.n3485 VDD.n3482 0.0269375
R14575 VDD.n3488 VDD.n3485 0.0269375
R14576 VDD.n3491 VDD.n3488 0.0269375
R14577 VDD.n3494 VDD.n3491 0.0269375
R14578 VDD.n3497 VDD.n3494 0.0269375
R14579 VDD.n3500 VDD.n3497 0.0269375
R14580 VDD.n3503 VDD.n3500 0.0269375
R14581 VDD.n3506 VDD.n3503 0.0269375
R14582 VDD.n3509 VDD.n3506 0.0269375
R14583 VDD.n3512 VDD.n3509 0.0269375
R14584 VDD.n3515 VDD.n3512 0.0269375
R14585 VDD.n3518 VDD.n3515 0.0269375
R14586 VDD.n3521 VDD.n3518 0.0269375
R14587 VDD.n3524 VDD.n3521 0.0269375
R14588 VDD.n3527 VDD.n3524 0.0269375
R14589 VDD.n3530 VDD.n3527 0.0269375
R14590 VDD.n3533 VDD.n3530 0.0269375
R14591 VDD.n3536 VDD.n3533 0.0269375
R14592 VDD.n3539 VDD.n3536 0.0269375
R14593 VDD.n3542 VDD.n3539 0.0269375
R14594 VDD.n3545 VDD.n3542 0.0269375
R14595 VDD.n3548 VDD.n3545 0.0269375
R14596 VDD.n3551 VDD.n3548 0.0269375
R14597 VDD.n3554 VDD.n3551 0.0269375
R14598 VDD.n3557 VDD.n3554 0.0269375
R14599 VDD.n3560 VDD.n3557 0.0269375
R14600 VDD.n3563 VDD.n3560 0.0269375
R14601 VDD.n3566 VDD.n3563 0.0269375
R14602 VDD.n3569 VDD.n3566 0.0269375
R14603 VDD.n3572 VDD.n3569 0.0269375
R14604 VDD.n3575 VDD.n3572 0.0269375
R14605 VDD.n3578 VDD.n3575 0.0269375
R14606 VDD.n3581 VDD.n3578 0.0269375
R14607 VDD.n3583 VDD.n3581 0.0269375
R14608 VDD.n3586 VDD.n3583 0.0269375
R14609 VDD.n5561 VDD.n5559 0.0269375
R14610 VDD.n5559 VDD.n5556 0.0269375
R14611 VDD.n5556 VDD.n5553 0.0269375
R14612 VDD.n5553 VDD.n5550 0.0269375
R14613 VDD.n3959 VDD.n3956 0.0269375
R14614 VDD.n3962 VDD.n3959 0.0269375
R14615 VDD.n3965 VDD.n3962 0.0269375
R14616 VDD.n3968 VDD.n3965 0.0269375
R14617 VDD.n3971 VDD.n3968 0.0269375
R14618 VDD.n3974 VDD.n3971 0.0269375
R14619 VDD.n3977 VDD.n3974 0.0269375
R14620 VDD.n3980 VDD.n3977 0.0269375
R14621 VDD.n3983 VDD.n3980 0.0269375
R14622 VDD.n3986 VDD.n3983 0.0269375
R14623 VDD.n3989 VDD.n3986 0.0269375
R14624 VDD.n3992 VDD.n3989 0.0269375
R14625 VDD.n3995 VDD.n3992 0.0269375
R14626 VDD.n3998 VDD.n3995 0.0269375
R14627 VDD.n4001 VDD.n3998 0.0269375
R14628 VDD.n4004 VDD.n4001 0.0269375
R14629 VDD.n4007 VDD.n4004 0.0269375
R14630 VDD.n4010 VDD.n4007 0.0269375
R14631 VDD.n4013 VDD.n4010 0.0269375
R14632 VDD.n4016 VDD.n4013 0.0269375
R14633 VDD.n4019 VDD.n4016 0.0269375
R14634 VDD.n4022 VDD.n4019 0.0269375
R14635 VDD.n4025 VDD.n4022 0.0269375
R14636 VDD.n4028 VDD.n4025 0.0269375
R14637 VDD.n4031 VDD.n4028 0.0269375
R14638 VDD.n4034 VDD.n4031 0.0269375
R14639 VDD.n4037 VDD.n4034 0.0269375
R14640 VDD.n4040 VDD.n4037 0.0269375
R14641 VDD.n4043 VDD.n4040 0.0269375
R14642 VDD.n4046 VDD.n4043 0.0269375
R14643 VDD.n4049 VDD.n4046 0.0269375
R14644 VDD.n4052 VDD.n4049 0.0269375
R14645 VDD.n4055 VDD.n4052 0.0269375
R14646 VDD.n4058 VDD.n4055 0.0269375
R14647 VDD.n4061 VDD.n4058 0.0269375
R14648 VDD.n4064 VDD.n4061 0.0269375
R14649 VDD.n4067 VDD.n4064 0.0269375
R14650 VDD.n4070 VDD.n4067 0.0269375
R14651 VDD.n4073 VDD.n4070 0.0269375
R14652 VDD.n4076 VDD.n4073 0.0269375
R14653 VDD.n4078 VDD.n4076 0.0269375
R14654 VDD.n4081 VDD.n4078 0.0269375
R14655 VDD.n5418 VDD.n5415 0.0269375
R14656 VDD.n5415 VDD.n5413 0.0269375
R14657 VDD.n3591 VDD.n3588 0.0269375
R14658 VDD.n3593 VDD.n3591 0.0269375
R14659 VDD.n3596 VDD.n3593 0.0269375
R14660 VDD.n3598 VDD.n3596 0.0269375
R14661 VDD.n3601 VDD.n3598 0.0269375
R14662 VDD.n3603 VDD.n3601 0.0269375
R14663 VDD.n3606 VDD.n3603 0.0269375
R14664 VDD.n3608 VDD.n3606 0.0269375
R14665 VDD.n3611 VDD.n3608 0.0269375
R14666 VDD.n3613 VDD.n3611 0.0269375
R14667 VDD.n3616 VDD.n3613 0.0269375
R14668 VDD.n3618 VDD.n3616 0.0269375
R14669 VDD.n3621 VDD.n3618 0.0269375
R14670 VDD.n3623 VDD.n3621 0.0269375
R14671 VDD.n3626 VDD.n3623 0.0269375
R14672 VDD.n3628 VDD.n3626 0.0269375
R14673 VDD.n3631 VDD.n3628 0.0269375
R14674 VDD.n3633 VDD.n3631 0.0269375
R14675 VDD.n3636 VDD.n3633 0.0269375
R14676 VDD.n3638 VDD.n3636 0.0269375
R14677 VDD.n3641 VDD.n3638 0.0269375
R14678 VDD.n3643 VDD.n3641 0.0269375
R14679 VDD.n3646 VDD.n3643 0.0269375
R14680 VDD.n3648 VDD.n3646 0.0269375
R14681 VDD.n3651 VDD.n3648 0.0269375
R14682 VDD.n3653 VDD.n3651 0.0269375
R14683 VDD.n3656 VDD.n3653 0.0269375
R14684 VDD.n3658 VDD.n3656 0.0269375
R14685 VDD.n3661 VDD.n3658 0.0269375
R14686 VDD.n3663 VDD.n3661 0.0269375
R14687 VDD.n3666 VDD.n3663 0.0269375
R14688 VDD.n3668 VDD.n3666 0.0269375
R14689 VDD.n3671 VDD.n3668 0.0269375
R14690 VDD.n3673 VDD.n3671 0.0269375
R14691 VDD.n3676 VDD.n3673 0.0269375
R14692 VDD.n3678 VDD.n3676 0.0269375
R14693 VDD.n3681 VDD.n3678 0.0269375
R14694 VDD.n3683 VDD.n3681 0.0269375
R14695 VDD.n3686 VDD.n3683 0.0269375
R14696 VDD.n3688 VDD.n3686 0.0269375
R14697 VDD.n3691 VDD.n3688 0.0269375
R14698 VDD.n3694 VDD.n3691 0.0269375
R14699 VDD.n3696 VDD.n3694 0.0269375
R14700 VDD.n3699 VDD.n3696 0.0269375
R14701 VDD.n5850 VDD.n5848 0.0269375
R14702 VDD.n5852 VDD.n5850 0.0269375
R14703 VDD.n5854 VDD.n5852 0.0269375
R14704 VDD.n5859 VDD.n5857 0.0269375
R14705 VDD.n5864 VDD.n5862 0.0269375
R14706 VDD.n5866 VDD.n5864 0.0269375
R14707 VDD.n5871 VDD.n5869 0.0269375
R14708 VDD.n5873 VDD.n5871 0.0269375
R14709 VDD.n5878 VDD.n5876 0.0269375
R14710 VDD.n5880 VDD.n5878 0.0269375
R14711 VDD.n5885 VDD.n5883 0.0269375
R14712 VDD.n5887 VDD.n5885 0.0269375
R14713 VDD.n5889 VDD.n5887 0.0269375
R14714 VDD.n5891 VDD.n5889 0.0269375
R14715 VDD.n5893 VDD.n5891 0.0269375
R14716 VDD.n5895 VDD.n5893 0.0269375
R14717 VDD.n5897 VDD.n5895 0.0269375
R14718 VDD.n5899 VDD.n5897 0.0269375
R14719 VDD.n5901 VDD.n5899 0.0269375
R14720 VDD.n5903 VDD.n5901 0.0269375
R14721 VDD.n5908 VDD.n5906 0.0269375
R14722 VDD.n5910 VDD.n5908 0.0269375
R14723 VDD.n5915 VDD.n5913 0.0269375
R14724 VDD.n5917 VDD.n5915 0.0269375
R14725 VDD.n5922 VDD.n5920 0.0269375
R14726 VDD.n5924 VDD.n5922 0.0269375
R14727 VDD.n5929 VDD.n5927 0.0269375
R14728 VDD.n5934 VDD.n5932 0.0269375
R14729 VDD.n5936 VDD.n5934 0.0269375
R14730 VDD.n5938 VDD.n5936 0.0269375
R14731 VDD.n5940 VDD.n5938 0.0269375
R14732 VDD.n5956 VDD.n5954 0.0269375
R14733 VDD.n5958 VDD.n5956 0.0269375
R14734 VDD.n5960 VDD.n5958 0.0269375
R14735 VDD.n5962 VDD.n5960 0.0269375
R14736 VDD.n5967 VDD.n5965 0.0269375
R14737 VDD.n5972 VDD.n5970 0.0269375
R14738 VDD.n5974 VDD.n5972 0.0269375
R14739 VDD.n5979 VDD.n5977 0.0269375
R14740 VDD.n5981 VDD.n5979 0.0269375
R14741 VDD.n5986 VDD.n5984 0.0269375
R14742 VDD.n5988 VDD.n5986 0.0269375
R14743 VDD.n5993 VDD.n5991 0.0269375
R14744 VDD.n5995 VDD.n5993 0.0269375
R14745 VDD.n5997 VDD.n5995 0.0269375
R14746 VDD.n5999 VDD.n5997 0.0269375
R14747 VDD.n6001 VDD.n5999 0.0269375
R14748 VDD.n6003 VDD.n6001 0.0269375
R14749 VDD.n6005 VDD.n6003 0.0269375
R14750 VDD.n6007 VDD.n6005 0.0269375
R14751 VDD.n6009 VDD.n6007 0.0269375
R14752 VDD.n6011 VDD.n6009 0.0269375
R14753 VDD.n6016 VDD.n6014 0.0269375
R14754 VDD.n6018 VDD.n6016 0.0269375
R14755 VDD.n6023 VDD.n6021 0.0269375
R14756 VDD.n6025 VDD.n6023 0.0269375
R14757 VDD.n6030 VDD.n6028 0.0269375
R14758 VDD.n6032 VDD.n6030 0.0269375
R14759 VDD.n6037 VDD.n6035 0.0269375
R14760 VDD.n6047 VDD.n6045 0.0269375
R14761 VDD.n6049 VDD.n6047 0.0269375
R14762 VDD.n6051 VDD.n6049 0.0269375
R14763 VDD.n4668 VDD.n4665 0.0269375
R14764 VDD.n4673 VDD.n4668 0.0269375
R14765 VDD.n4680 VDD.n4677 0.0269375
R14766 VDD.n4683 VDD.n4680 0.0269375
R14767 VDD.n4686 VDD.n4683 0.0269375
R14768 VDD.n4689 VDD.n4686 0.0269375
R14769 VDD.n4696 VDD.n4693 0.0269375
R14770 VDD.n4703 VDD.n4700 0.0269375
R14771 VDD.n4706 VDD.n4703 0.0269375
R14772 VDD.n4713 VDD.n4710 0.0269375
R14773 VDD.n4716 VDD.n4713 0.0269375
R14774 VDD.n4723 VDD.n4720 0.0269375
R14775 VDD.n4726 VDD.n4723 0.0269375
R14776 VDD.n4733 VDD.n4730 0.0269375
R14777 VDD.n4736 VDD.n4733 0.0269375
R14778 VDD.n4739 VDD.n4736 0.0269375
R14779 VDD.n4746 VDD.n4743 0.0269375
R14780 VDD.n4749 VDD.n4746 0.0269375
R14781 VDD.n4756 VDD.n4753 0.0269375
R14782 VDD.n4759 VDD.n4756 0.0269375
R14783 VDD.n4762 VDD.n4759 0.0269375
R14784 VDD.n4769 VDD.n4766 0.0269375
R14785 VDD.n4772 VDD.n4769 0.0269375
R14786 VDD.n4779 VDD.n4776 0.0269375
R14787 VDD.n4782 VDD.n4779 0.0269375
R14788 VDD.n4789 VDD.n4786 0.0269375
R14789 VDD.n4792 VDD.n4789 0.0269375
R14790 VDD.n4799 VDD.n4796 0.0269375
R14791 VDD.n4806 VDD.n4803 0.0269375
R14792 VDD.n4809 VDD.n4806 0.0269375
R14793 VDD.n4812 VDD.n4809 0.0269375
R14794 VDD.n4815 VDD.n4812 0.0269375
R14795 VDD.n4835 VDD.n4832 0.0269375
R14796 VDD.n4838 VDD.n4835 0.0269375
R14797 VDD.n4841 VDD.n4838 0.0269375
R14798 VDD.n4844 VDD.n4841 0.0269375
R14799 VDD.n4851 VDD.n4848 0.0269375
R14800 VDD.n4858 VDD.n4855 0.0269375
R14801 VDD.n4861 VDD.n4858 0.0269375
R14802 VDD.n4868 VDD.n4865 0.0269375
R14803 VDD.n4871 VDD.n4868 0.0269375
R14804 VDD.n4878 VDD.n4875 0.0269375
R14805 VDD.n4881 VDD.n4878 0.0269375
R14806 VDD.n4888 VDD.n4885 0.0269375
R14807 VDD.n4891 VDD.n4888 0.0269375
R14808 VDD.n4894 VDD.n4891 0.0269375
R14809 VDD.n4901 VDD.n4898 0.0269375
R14810 VDD.n4904 VDD.n4901 0.0269375
R14811 VDD.n4911 VDD.n4908 0.0269375
R14812 VDD.n4914 VDD.n4911 0.0269375
R14813 VDD.n4917 VDD.n4914 0.0269375
R14814 VDD.n4924 VDD.n4921 0.0269375
R14815 VDD.n4927 VDD.n4924 0.0269375
R14816 VDD.n4934 VDD.n4931 0.0269375
R14817 VDD.n4937 VDD.n4934 0.0269375
R14818 VDD.n4944 VDD.n4941 0.0269375
R14819 VDD.n4947 VDD.n4944 0.0269375
R14820 VDD.n4954 VDD.n4951 0.0269375
R14821 VDD.n4961 VDD.n4958 0.0269375
R14822 VDD.n4964 VDD.n4961 0.0269375
R14823 VDD.n4967 VDD.n4964 0.0269375
R14824 VDD.n4970 VDD.n4967 0.0269375
R14825 VDD.n5281 VDD.n5278 0.0269375
R14826 VDD.n3084 VDD.n3082 0.0269375
R14827 VDD.n3087 VDD.n3084 0.0269375
R14828 VDD.n3089 VDD.n3087 0.0269375
R14829 VDD.n3092 VDD.n3089 0.0269375
R14830 VDD.n3094 VDD.n3092 0.0269375
R14831 VDD.n3097 VDD.n3094 0.0269375
R14832 VDD.n3099 VDD.n3097 0.0269375
R14833 VDD.n3102 VDD.n3099 0.0269375
R14834 VDD.n3104 VDD.n3102 0.0269375
R14835 VDD.n3107 VDD.n3104 0.0269375
R14836 VDD.n3109 VDD.n3107 0.0269375
R14837 VDD.n3112 VDD.n3109 0.0269375
R14838 VDD.n3114 VDD.n3112 0.0269375
R14839 VDD.n3117 VDD.n3114 0.0269375
R14840 VDD.n3119 VDD.n3117 0.0269375
R14841 VDD.n3122 VDD.n3119 0.0269375
R14842 VDD.n3124 VDD.n3122 0.0269375
R14843 VDD.n3127 VDD.n3124 0.0269375
R14844 VDD.n3129 VDD.n3127 0.0269375
R14845 VDD.n3132 VDD.n3129 0.0269375
R14846 VDD.n3134 VDD.n3132 0.0269375
R14847 VDD.n3137 VDD.n3134 0.0269375
R14848 VDD.n3139 VDD.n3137 0.0269375
R14849 VDD.n3142 VDD.n3139 0.0269375
R14850 VDD.n3144 VDD.n3142 0.0269375
R14851 VDD.n3147 VDD.n3144 0.0269375
R14852 VDD.n3149 VDD.n3147 0.0269375
R14853 VDD.n3152 VDD.n3149 0.0269375
R14854 VDD.n3154 VDD.n3152 0.0269375
R14855 VDD.n3157 VDD.n3154 0.0269375
R14856 VDD.n3159 VDD.n3157 0.0269375
R14857 VDD.n3162 VDD.n3159 0.0269375
R14858 VDD.n3164 VDD.n3162 0.0269375
R14859 VDD.n3167 VDD.n3164 0.0269375
R14860 VDD.n3169 VDD.n3167 0.0269375
R14861 VDD.n3172 VDD.n3169 0.0269375
R14862 VDD.n3174 VDD.n3172 0.0269375
R14863 VDD.n3177 VDD.n3174 0.0269375
R14864 VDD.n3179 VDD.n3177 0.0269375
R14865 VDD.n3182 VDD.n3179 0.0269375
R14866 VDD.n3184 VDD.n3182 0.0269375
R14867 VDD.n3187 VDD.n3184 0.0269375
R14868 VDD.n3190 VDD.n3187 0.0269375
R14869 VDD.n3192 VDD.n3190 0.0269375
R14870 VDD.n3195 VDD.n3192 0.0269375
R14871 VDD.n5275 VDD.n5273 0.0269375
R14872 VDD.n2969 VDD.n2967 0.0269375
R14873 VDD.n2972 VDD.n2969 0.0269375
R14874 VDD.n2974 VDD.n2972 0.0269375
R14875 VDD.n2977 VDD.n2974 0.0269375
R14876 VDD.n2979 VDD.n2977 0.0269375
R14877 VDD.n2982 VDD.n2979 0.0269375
R14878 VDD.n2984 VDD.n2982 0.0269375
R14879 VDD.n2987 VDD.n2984 0.0269375
R14880 VDD.n2989 VDD.n2987 0.0269375
R14881 VDD.n2992 VDD.n2989 0.0269375
R14882 VDD.n2994 VDD.n2992 0.0269375
R14883 VDD.n2997 VDD.n2994 0.0269375
R14884 VDD.n2999 VDD.n2997 0.0269375
R14885 VDD.n3002 VDD.n2999 0.0269375
R14886 VDD.n3004 VDD.n3002 0.0269375
R14887 VDD.n3007 VDD.n3004 0.0269375
R14888 VDD.n3009 VDD.n3007 0.0269375
R14889 VDD.n3012 VDD.n3009 0.0269375
R14890 VDD.n3014 VDD.n3012 0.0269375
R14891 VDD.n3017 VDD.n3014 0.0269375
R14892 VDD.n3019 VDD.n3017 0.0269375
R14893 VDD.n3022 VDD.n3019 0.0269375
R14894 VDD.n3024 VDD.n3022 0.0269375
R14895 VDD.n3027 VDD.n3024 0.0269375
R14896 VDD.n3029 VDD.n3027 0.0269375
R14897 VDD.n3032 VDD.n3029 0.0269375
R14898 VDD.n3034 VDD.n3032 0.0269375
R14899 VDD.n3037 VDD.n3034 0.0269375
R14900 VDD.n3039 VDD.n3037 0.0269375
R14901 VDD.n3042 VDD.n3039 0.0269375
R14902 VDD.n3044 VDD.n3042 0.0269375
R14903 VDD.n3047 VDD.n3044 0.0269375
R14904 VDD.n3049 VDD.n3047 0.0269375
R14905 VDD.n3052 VDD.n3049 0.0269375
R14906 VDD.n3054 VDD.n3052 0.0269375
R14907 VDD.n3057 VDD.n3054 0.0269375
R14908 VDD.n3059 VDD.n3057 0.0269375
R14909 VDD.n3062 VDD.n3059 0.0269375
R14910 VDD.n3064 VDD.n3062 0.0269375
R14911 VDD.n3067 VDD.n3064 0.0269375
R14912 VDD.n3069 VDD.n3067 0.0269375
R14913 VDD.n3072 VDD.n3069 0.0269375
R14914 VDD.n3074 VDD.n3072 0.0269375
R14915 VDD.n3077 VDD.n3074 0.0269375
R14916 VDD.n3079 VDD.n3077 0.0269375
R14917 VDD.n6056 VDD.n6054 0.0269375
R14918 VDD.n6058 VDD.n6056 0.0269375
R14919 VDD.n6060 VDD.n6058 0.0269375
R14920 VDD.n6065 VDD.n6063 0.0269375
R14921 VDD.n6070 VDD.n6068 0.0269375
R14922 VDD.n6072 VDD.n6070 0.0269375
R14923 VDD.n6077 VDD.n6075 0.0269375
R14924 VDD.n6079 VDD.n6077 0.0269375
R14925 VDD.n6084 VDD.n6082 0.0269375
R14926 VDD.n6086 VDD.n6084 0.0269375
R14927 VDD.n6091 VDD.n6089 0.0269375
R14928 VDD.n6093 VDD.n6091 0.0269375
R14929 VDD.n6095 VDD.n6093 0.0269375
R14930 VDD.n6097 VDD.n6095 0.0269375
R14931 VDD.n6099 VDD.n6097 0.0269375
R14932 VDD.n6101 VDD.n6099 0.0269375
R14933 VDD.n6103 VDD.n6101 0.0269375
R14934 VDD.n6105 VDD.n6103 0.0269375
R14935 VDD.n6107 VDD.n6105 0.0269375
R14936 VDD.n6109 VDD.n6107 0.0269375
R14937 VDD.n6114 VDD.n6112 0.0269375
R14938 VDD.n6116 VDD.n6114 0.0269375
R14939 VDD.n6121 VDD.n6119 0.0269375
R14940 VDD.n6123 VDD.n6121 0.0269375
R14941 VDD.n6128 VDD.n6126 0.0269375
R14942 VDD.n6130 VDD.n6128 0.0269375
R14943 VDD.n6135 VDD.n6133 0.0269375
R14944 VDD.n6140 VDD.n6138 0.0269375
R14945 VDD.n6142 VDD.n6140 0.0269375
R14946 VDD.n6144 VDD.n6142 0.0269375
R14947 VDD.n6146 VDD.n6144 0.0269375
R14948 VDD.n6305 VDD.n6303 0.0269375
R14949 VDD.n6303 VDD.n6301 0.0269375
R14950 VDD.n6301 VDD.n6299 0.0269375
R14951 VDD.n6299 VDD.n6297 0.0269375
R14952 VDD.n6294 VDD.n6292 0.0269375
R14953 VDD.n6289 VDD.n6287 0.0269375
R14954 VDD.n6287 VDD.n6285 0.0269375
R14955 VDD.n6282 VDD.n6280 0.0269375
R14956 VDD.n6280 VDD.n6278 0.0269375
R14957 VDD.n6275 VDD.n6273 0.0269375
R14958 VDD.n6273 VDD.n6271 0.0269375
R14959 VDD.n6268 VDD.n6266 0.0269375
R14960 VDD.n6266 VDD.n6264 0.0269375
R14961 VDD.n6264 VDD.n6262 0.0269375
R14962 VDD.n6262 VDD.n6260 0.0269375
R14963 VDD.n6260 VDD.n6258 0.0269375
R14964 VDD.n6258 VDD.n6256 0.0269375
R14965 VDD.n6256 VDD.n6254 0.0269375
R14966 VDD.n6254 VDD.n6252 0.0269375
R14967 VDD.n6252 VDD.n6250 0.0269375
R14968 VDD.n6250 VDD.n6248 0.0269375
R14969 VDD.n6245 VDD.n6243 0.0269375
R14970 VDD.n6243 VDD.n6241 0.0269375
R14971 VDD.n6238 VDD.n6236 0.0269375
R14972 VDD.n6236 VDD.n6234 0.0269375
R14973 VDD.n6231 VDD.n6229 0.0269375
R14974 VDD.n6229 VDD.n6227 0.0269375
R14975 VDD.n6224 VDD.n6222 0.0269375
R14976 VDD.n6214 VDD.n6212 0.0269375
R14977 VDD.n6212 VDD.n6210 0.0269375
R14978 VDD.n6210 VDD.n5271 0.0269375
R14979 VDD.n4975 VDD.n4970 0.0269375
R14980 VDD.n4982 VDD.n4979 0.0269375
R14981 VDD.n4985 VDD.n4982 0.0269375
R14982 VDD.n4988 VDD.n4985 0.0269375
R14983 VDD.n4991 VDD.n4988 0.0269375
R14984 VDD.n4998 VDD.n4995 0.0269375
R14985 VDD.n5005 VDD.n5002 0.0269375
R14986 VDD.n5008 VDD.n5005 0.0269375
R14987 VDD.n5015 VDD.n5012 0.0269375
R14988 VDD.n5018 VDD.n5015 0.0269375
R14989 VDD.n5025 VDD.n5022 0.0269375
R14990 VDD.n5028 VDD.n5025 0.0269375
R14991 VDD.n5035 VDD.n5032 0.0269375
R14992 VDD.n5038 VDD.n5035 0.0269375
R14993 VDD.n5041 VDD.n5038 0.0269375
R14994 VDD.n5048 VDD.n5045 0.0269375
R14995 VDD.n5051 VDD.n5048 0.0269375
R14996 VDD.n5058 VDD.n5055 0.0269375
R14997 VDD.n5061 VDD.n5058 0.0269375
R14998 VDD.n5064 VDD.n5061 0.0269375
R14999 VDD.n5071 VDD.n5068 0.0269375
R15000 VDD.n5074 VDD.n5071 0.0269375
R15001 VDD.n5081 VDD.n5078 0.0269375
R15002 VDD.n5084 VDD.n5081 0.0269375
R15003 VDD.n5091 VDD.n5088 0.0269375
R15004 VDD.n5094 VDD.n5091 0.0269375
R15005 VDD.n5101 VDD.n5098 0.0269375
R15006 VDD.n5108 VDD.n5105 0.0269375
R15007 VDD.n5111 VDD.n5108 0.0269375
R15008 VDD.n5114 VDD.n5111 0.0269375
R15009 VDD.n5117 VDD.n5114 0.0269375
R15010 VDD.n5137 VDD.n5134 0.0269375
R15011 VDD.n5140 VDD.n5137 0.0269375
R15012 VDD.n5143 VDD.n5140 0.0269375
R15013 VDD.n5146 VDD.n5143 0.0269375
R15014 VDD.n5153 VDD.n5150 0.0269375
R15015 VDD.n5160 VDD.n5157 0.0269375
R15016 VDD.n5163 VDD.n5160 0.0269375
R15017 VDD.n5170 VDD.n5167 0.0269375
R15018 VDD.n5173 VDD.n5170 0.0269375
R15019 VDD.n5180 VDD.n5177 0.0269375
R15020 VDD.n5183 VDD.n5180 0.0269375
R15021 VDD.n5190 VDD.n5187 0.0269375
R15022 VDD.n5193 VDD.n5190 0.0269375
R15023 VDD.n5196 VDD.n5193 0.0269375
R15024 VDD.n5203 VDD.n5200 0.0269375
R15025 VDD.n5206 VDD.n5203 0.0269375
R15026 VDD.n5213 VDD.n5210 0.0269375
R15027 VDD.n5216 VDD.n5213 0.0269375
R15028 VDD.n5219 VDD.n5216 0.0269375
R15029 VDD.n5226 VDD.n5223 0.0269375
R15030 VDD.n5229 VDD.n5226 0.0269375
R15031 VDD.n5236 VDD.n5233 0.0269375
R15032 VDD.n5239 VDD.n5236 0.0269375
R15033 VDD.n5246 VDD.n5243 0.0269375
R15034 VDD.n5249 VDD.n5246 0.0269375
R15035 VDD.n5256 VDD.n5253 0.0269375
R15036 VDD.n5263 VDD.n5260 0.0269375
R15037 VDD.n5266 VDD.n5263 0.0269375
R15038 VDD.n5269 VDD.n5266 0.0269375
R15039 VDD.n2690 VDD.n2687 0.0269375
R15040 VDD.n2693 VDD.n2690 0.0269375
R15041 VDD.n2696 VDD.n2693 0.0269375
R15042 VDD.n2699 VDD.n2696 0.0269375
R15043 VDD.n2702 VDD.n2699 0.0269375
R15044 VDD.n2705 VDD.n2702 0.0269375
R15045 VDD.n2708 VDD.n2705 0.0269375
R15046 VDD.n2711 VDD.n2708 0.0269375
R15047 VDD.n2714 VDD.n2711 0.0269375
R15048 VDD.n2717 VDD.n2714 0.0269375
R15049 VDD.n2720 VDD.n2717 0.0269375
R15050 VDD.n2723 VDD.n2720 0.0269375
R15051 VDD.n2726 VDD.n2723 0.0269375
R15052 VDD.n2729 VDD.n2726 0.0269375
R15053 VDD.n2732 VDD.n2729 0.0269375
R15054 VDD.n2735 VDD.n2732 0.0269375
R15055 VDD.n2738 VDD.n2735 0.0269375
R15056 VDD.n2741 VDD.n2738 0.0269375
R15057 VDD.n2744 VDD.n2741 0.0269375
R15058 VDD.n2747 VDD.n2744 0.0269375
R15059 VDD.n2750 VDD.n2747 0.0269375
R15060 VDD.n2753 VDD.n2750 0.0269375
R15061 VDD.n2756 VDD.n2753 0.0269375
R15062 VDD.n2759 VDD.n2756 0.0269375
R15063 VDD.n2762 VDD.n2759 0.0269375
R15064 VDD.n2765 VDD.n2762 0.0269375
R15065 VDD.n2768 VDD.n2765 0.0269375
R15066 VDD.n2771 VDD.n2768 0.0269375
R15067 VDD.n2774 VDD.n2771 0.0269375
R15068 VDD.n2777 VDD.n2774 0.0269375
R15069 VDD.n2780 VDD.n2777 0.0269375
R15070 VDD.n2783 VDD.n2780 0.0269375
R15071 VDD.n2786 VDD.n2783 0.0269375
R15072 VDD.n2789 VDD.n2786 0.0269375
R15073 VDD.n2792 VDD.n2789 0.0269375
R15074 VDD.n2795 VDD.n2792 0.0269375
R15075 VDD.n2798 VDD.n2795 0.0269375
R15076 VDD.n2801 VDD.n2798 0.0269375
R15077 VDD.n2804 VDD.n2801 0.0269375
R15078 VDD.n2807 VDD.n2804 0.0269375
R15079 VDD.n2810 VDD.n2807 0.0269375
R15080 VDD.n2813 VDD.n2810 0.0269375
R15081 VDD.n2816 VDD.n2813 0.0269375
R15082 VDD.n2819 VDD.n2816 0.0269375
R15083 VDD.n2822 VDD.n2819 0.0269375
R15084 VDD.n2825 VDD.n2822 0.0269375
R15085 VDD.n2828 VDD.n2825 0.0269375
R15086 VDD.n6318 VDD.n6316 0.0269375
R15087 VDD.n2590 VDD.n2588 0.0269375
R15088 VDD.n2595 VDD.n2593 0.0269375
R15089 VDD.n2600 VDD.n2598 0.0269375
R15090 VDD.n2602 VDD.n2600 0.0269375
R15091 VDD.n2607 VDD.n2605 0.0269375
R15092 VDD.n2609 VDD.n2607 0.0269375
R15093 VDD.n2614 VDD.n2612 0.0269375
R15094 VDD.n2616 VDD.n2614 0.0269375
R15095 VDD.n2621 VDD.n2619 0.0269375
R15096 VDD.n2623 VDD.n2621 0.0269375
R15097 VDD.n2625 VDD.n2623 0.0269375
R15098 VDD.n2627 VDD.n2625 0.0269375
R15099 VDD.n2629 VDD.n2627 0.0269375
R15100 VDD.n2631 VDD.n2629 0.0269375
R15101 VDD.n2633 VDD.n2631 0.0269375
R15102 VDD.n2635 VDD.n2633 0.0269375
R15103 VDD.n2637 VDD.n2635 0.0269375
R15104 VDD.n2639 VDD.n2637 0.0269375
R15105 VDD.n2644 VDD.n2642 0.0269375
R15106 VDD.n2646 VDD.n2644 0.0269375
R15107 VDD.n2651 VDD.n2649 0.0269375
R15108 VDD.n2653 VDD.n2651 0.0269375
R15109 VDD.n2658 VDD.n2656 0.0269375
R15110 VDD.n2660 VDD.n2658 0.0269375
R15111 VDD.n2665 VDD.n2663 0.0269375
R15112 VDD.n2675 VDD.n2673 0.0269375
R15113 VDD.n2677 VDD.n2675 0.0269375
R15114 VDD.n2679 VDD.n2677 0.0269375
R15115 VDD.n2681 VDD.n2679 0.0269375
R15116 VDD.n6462 VDD.n6459 0.0269375
R15117 VDD.n6465 VDD.n6462 0.0269375
R15118 VDD.n6468 VDD.n6465 0.0269375
R15119 VDD.n6475 VDD.n6472 0.0269375
R15120 VDD.n6482 VDD.n6479 0.0269375
R15121 VDD.n6485 VDD.n6482 0.0269375
R15122 VDD.n6492 VDD.n6489 0.0269375
R15123 VDD.n6495 VDD.n6492 0.0269375
R15124 VDD.n6502 VDD.n6499 0.0269375
R15125 VDD.n6505 VDD.n6502 0.0269375
R15126 VDD.n6512 VDD.n6509 0.0269375
R15127 VDD.n6515 VDD.n6512 0.0269375
R15128 VDD.n6518 VDD.n6515 0.0269375
R15129 VDD.n6525 VDD.n6522 0.0269375
R15130 VDD.n6528 VDD.n6525 0.0269375
R15131 VDD.n6535 VDD.n6532 0.0269375
R15132 VDD.n6538 VDD.n6535 0.0269375
R15133 VDD.n6541 VDD.n6538 0.0269375
R15134 VDD.n6548 VDD.n6545 0.0269375
R15135 VDD.n6551 VDD.n6548 0.0269375
R15136 VDD.n6558 VDD.n6555 0.0269375
R15137 VDD.n6561 VDD.n6558 0.0269375
R15138 VDD.n6568 VDD.n6565 0.0269375
R15139 VDD.n6571 VDD.n6568 0.0269375
R15140 VDD.n6578 VDD.n6575 0.0269375
R15141 VDD.n6585 VDD.n6582 0.0269375
R15142 VDD.n6588 VDD.n6585 0.0269375
R15143 VDD.n6591 VDD.n6588 0.0269375
R15144 VDD.n6594 VDD.n6591 0.0269375
R15145 VDD.n2031 VDD.n2029 0.0269375
R15146 VDD.n2029 VDD.n2026 0.0269375
R15147 VDD.n2026 VDD.n2024 0.0269375
R15148 VDD.n2024 VDD.n2021 0.0269375
R15149 VDD.n2021 VDD.n2019 0.0269375
R15150 VDD.n2019 VDD.n2016 0.0269375
R15151 VDD.n2016 VDD.n2014 0.0269375
R15152 VDD.n2014 VDD.n2011 0.0269375
R15153 VDD.n2011 VDD.n2009 0.0269375
R15154 VDD.n2009 VDD.n2006 0.0269375
R15155 VDD.n2006 VDD.n2004 0.0269375
R15156 VDD.n2004 VDD.n2001 0.0269375
R15157 VDD.n2001 VDD.n1999 0.0269375
R15158 VDD.n1999 VDD.n1996 0.0269375
R15159 VDD.n1996 VDD.n1994 0.0269375
R15160 VDD.n1994 VDD.n1991 0.0269375
R15161 VDD.n1991 VDD.n1989 0.0269375
R15162 VDD.n1989 VDD.n1986 0.0269375
R15163 VDD.n1986 VDD.n1984 0.0269375
R15164 VDD.n1984 VDD.n1981 0.0269375
R15165 VDD.n1981 VDD.n1979 0.0269375
R15166 VDD.n1979 VDD.n1977 0.0269375
R15167 VDD.n1977 VDD.n1975 0.0269375
R15168 VDD.n1975 VDD.n1973 0.0269375
R15169 VDD.n1973 VDD.n1971 0.0269375
R15170 VDD.n1971 VDD.n1969 0.0269375
R15171 VDD.n1969 VDD.n1967 0.0269375
R15172 VDD.n1967 VDD.n1965 0.0269375
R15173 VDD.n1965 VDD.n1963 0.0269375
R15174 VDD.n1963 VDD.n1961 0.0269375
R15175 VDD.n1961 VDD.n1959 0.0269375
R15176 VDD.n1959 VDD.n1957 0.0269375
R15177 VDD.n1957 VDD.n1955 0.0269375
R15178 VDD.n1955 VDD.n1953 0.0269375
R15179 VDD.n1953 VDD.n1951 0.0269375
R15180 VDD.n1951 VDD.n1949 0.0269375
R15181 VDD.n1949 VDD.n1947 0.0269375
R15182 VDD.n1947 VDD.n1945 0.0269375
R15183 VDD.n1945 VDD.n1943 0.0269375
R15184 VDD.n1943 VDD.n1941 0.0269375
R15185 VDD.n1941 VDD.n1939 0.0269375
R15186 VDD.n1939 VDD.n1937 0.0269375
R15187 VDD.n1937 VDD.n1935 0.0269375
R15188 VDD.n1935 VDD.n1933 0.0269375
R15189 VDD.n1933 VDD.n1931 0.0269375
R15190 VDD.n1927 VDD.n1925 0.0269375
R15191 VDD.n1925 VDD.n1922 0.0269375
R15192 VDD.n1922 VDD.n1919 0.0269375
R15193 VDD.n1919 VDD.n1916 0.0269375
R15194 VDD.n1916 VDD.n1913 0.0269375
R15195 VDD.n1913 VDD.n1910 0.0269375
R15196 VDD.n1910 VDD.n1907 0.0269375
R15197 VDD.n1907 VDD.n1904 0.0269375
R15198 VDD.n1904 VDD.n1901 0.0269375
R15199 VDD.n1901 VDD.n1898 0.0269375
R15200 VDD.n1898 VDD.n1895 0.0269375
R15201 VDD.n1895 VDD.n1892 0.0269375
R15202 VDD.n1892 VDD.n1889 0.0269375
R15203 VDD.n1889 VDD.n1886 0.0269375
R15204 VDD.n1886 VDD.n1883 0.0269375
R15205 VDD.n1883 VDD.n1880 0.0269375
R15206 VDD.n1880 VDD.n1877 0.0269375
R15207 VDD.n1877 VDD.n1874 0.0269375
R15208 VDD.n1874 VDD.n1871 0.0269375
R15209 VDD.n1871 VDD.n1868 0.0269375
R15210 VDD.n1868 VDD.n1865 0.0269375
R15211 VDD.n1865 VDD.n1862 0.0269375
R15212 VDD.n1862 VDD.n1859 0.0269375
R15213 VDD.n1859 VDD.n1856 0.0269375
R15214 VDD.n1856 VDD.n1853 0.0269375
R15215 VDD.n1853 VDD.n1850 0.0269375
R15216 VDD.n1850 VDD.n1847 0.0269375
R15217 VDD.n1847 VDD.n1844 0.0269375
R15218 VDD.n1844 VDD.n1841 0.0269375
R15219 VDD.n1841 VDD.n1838 0.0269375
R15220 VDD.n1838 VDD.n1835 0.0269375
R15221 VDD.n1835 VDD.n1832 0.0269375
R15222 VDD.n1832 VDD.n1829 0.0269375
R15223 VDD.n1829 VDD.n1826 0.0269375
R15224 VDD.n1826 VDD.n1823 0.0269375
R15225 VDD.n1823 VDD.n1820 0.0269375
R15226 VDD.n1820 VDD.n1817 0.0269375
R15227 VDD.n1817 VDD.n1814 0.0269375
R15228 VDD.n1814 VDD.n1811 0.0269375
R15229 VDD.n1811 VDD.n1808 0.0269375
R15230 VDD.n1808 VDD.n1806 0.0269375
R15231 VDD.n1806 VDD.n1804 0.0269375
R15232 VDD.n1804 VDD.n1802 0.0269375
R15233 VDD.n1802 VDD.n1799 0.0269375
R15234 VDD.n1799 VDD.n1797 0.0269375
R15235 VDD.n1789 VDD.n1787 0.0269375
R15236 VDD.n1787 VDD.n1784 0.0269375
R15237 VDD.n1784 VDD.n1781 0.0269375
R15238 VDD.n1781 VDD.n1778 0.0269375
R15239 VDD.n1778 VDD.n1775 0.0269375
R15240 VDD.n1775 VDD.n1772 0.0269375
R15241 VDD.n1772 VDD.n1769 0.0269375
R15242 VDD.n1769 VDD.n1766 0.0269375
R15243 VDD.n1766 VDD.n1763 0.0269375
R15244 VDD.n1763 VDD.n1760 0.0269375
R15245 VDD.n1760 VDD.n1757 0.0269375
R15246 VDD.n1757 VDD.n1754 0.0269375
R15247 VDD.n1754 VDD.n1751 0.0269375
R15248 VDD.n1751 VDD.n1748 0.0269375
R15249 VDD.n1748 VDD.n1745 0.0269375
R15250 VDD.n1745 VDD.n1742 0.0269375
R15251 VDD.n1742 VDD.n1739 0.0269375
R15252 VDD.n1739 VDD.n1736 0.0269375
R15253 VDD.n1736 VDD.n1733 0.0269375
R15254 VDD.n1733 VDD.n1730 0.0269375
R15255 VDD.n1730 VDD.n1727 0.0269375
R15256 VDD.n1727 VDD.n1724 0.0269375
R15257 VDD.n1724 VDD.n1721 0.0269375
R15258 VDD.n1721 VDD.n1718 0.0269375
R15259 VDD.n1718 VDD.n1715 0.0269375
R15260 VDD.n1715 VDD.n1712 0.0269375
R15261 VDD.n1712 VDD.n1709 0.0269375
R15262 VDD.n1709 VDD.n1706 0.0269375
R15263 VDD.n1706 VDD.n1703 0.0269375
R15264 VDD.n1703 VDD.n1700 0.0269375
R15265 VDD.n1700 VDD.n1697 0.0269375
R15266 VDD.n1697 VDD.n1694 0.0269375
R15267 VDD.n1694 VDD.n1691 0.0269375
R15268 VDD.n1691 VDD.n1688 0.0269375
R15269 VDD.n1688 VDD.n1685 0.0269375
R15270 VDD.n1685 VDD.n1682 0.0269375
R15271 VDD.n1682 VDD.n1679 0.0269375
R15272 VDD.n1679 VDD.n1676 0.0269375
R15273 VDD.n1676 VDD.n1673 0.0269375
R15274 VDD.n1673 VDD.n1670 0.0269375
R15275 VDD.n1670 VDD.n1668 0.0269375
R15276 VDD.n1668 VDD.n1666 0.0269375
R15277 VDD.n1666 VDD.n1664 0.0269375
R15278 VDD.n1664 VDD.n1661 0.0269375
R15279 VDD.n1661 VDD.n1659 0.0269375
R15280 VDD.n1343 VDD.n1342 0.0269375
R15281 VDD.n1342 VDD.n1339 0.0269375
R15282 VDD.n1339 VDD.n1337 0.0269375
R15283 VDD.n1337 VDD.n1334 0.0269375
R15284 VDD.n1334 VDD.n1332 0.0269375
R15285 VDD.n1332 VDD.n1329 0.0269375
R15286 VDD.n1329 VDD.n1327 0.0269375
R15287 VDD.n1327 VDD.n1324 0.0269375
R15288 VDD.n1324 VDD.n1322 0.0269375
R15289 VDD.n1322 VDD.n1319 0.0269375
R15290 VDD.n1319 VDD.n1317 0.0269375
R15291 VDD.n1317 VDD.n1314 0.0269375
R15292 VDD.n1314 VDD.n1312 0.0269375
R15293 VDD.n1312 VDD.n1309 0.0269375
R15294 VDD.n1309 VDD.n1307 0.0269375
R15295 VDD.n1307 VDD.n1304 0.0269375
R15296 VDD.n1304 VDD.n1302 0.0269375
R15297 VDD.n1302 VDD.n1299 0.0269375
R15298 VDD.n1299 VDD.n1297 0.0269375
R15299 VDD.n1297 VDD.n1294 0.0269375
R15300 VDD.n1294 VDD.n1292 0.0269375
R15301 VDD.n1292 VDD.n1290 0.0269375
R15302 VDD.n1290 VDD.n1288 0.0269375
R15303 VDD.n1288 VDD.n1286 0.0269375
R15304 VDD.n1286 VDD.n1284 0.0269375
R15305 VDD.n1284 VDD.n1282 0.0269375
R15306 VDD.n1282 VDD.n1280 0.0269375
R15307 VDD.n1280 VDD.n1278 0.0269375
R15308 VDD.n1278 VDD.n1276 0.0269375
R15309 VDD.n1276 VDD.n1274 0.0269375
R15310 VDD.n1274 VDD.n1272 0.0269375
R15311 VDD.n1272 VDD.n1270 0.0269375
R15312 VDD.n1270 VDD.n1268 0.0269375
R15313 VDD.n1268 VDD.n1266 0.0269375
R15314 VDD.n1266 VDD.n1264 0.0269375
R15315 VDD.n1264 VDD.n1262 0.0269375
R15316 VDD.n1262 VDD.n1260 0.0269375
R15317 VDD.n1260 VDD.n1258 0.0269375
R15318 VDD.n1258 VDD.n1256 0.0269375
R15319 VDD.n1256 VDD.n1254 0.0269375
R15320 VDD.n1254 VDD.n1252 0.0269375
R15321 VDD.n1252 VDD.n1250 0.0269375
R15322 VDD.n1250 VDD.n1248 0.0269375
R15323 VDD.n1248 VDD.n1246 0.0269375
R15324 VDD.n1246 VDD.n1244 0.0269375
R15325 VDD.n1464 VDD.n1462 0.0269375
R15326 VDD.n1466 VDD.n1464 0.0269375
R15327 VDD.n1468 VDD.n1466 0.0269375
R15328 VDD.n1470 VDD.n1468 0.0269375
R15329 VDD.n1472 VDD.n1470 0.0269375
R15330 VDD.n1477 VDD.n1475 0.0269375
R15331 VDD.n1479 VDD.n1477 0.0269375
R15332 VDD.n1481 VDD.n1479 0.0269375
R15333 VDD.n1483 VDD.n1481 0.0269375
R15334 VDD.n1485 VDD.n1483 0.0269375
R15335 VDD.n1487 VDD.n1485 0.0269375
R15336 VDD.n1489 VDD.n1487 0.0269375
R15337 VDD.n1491 VDD.n1489 0.0269375
R15338 VDD.n1493 VDD.n1491 0.0269375
R15339 VDD.n1495 VDD.n1493 0.0269375
R15340 VDD.n1497 VDD.n1495 0.0269375
R15341 VDD.n1499 VDD.n1497 0.0269375
R15342 VDD.n1501 VDD.n1499 0.0269375
R15343 VDD.n1503 VDD.n1501 0.0269375
R15344 VDD.n1505 VDD.n1503 0.0269375
R15345 VDD.n1507 VDD.n1505 0.0269375
R15346 VDD.n1509 VDD.n1507 0.0269375
R15347 VDD.n1511 VDD.n1509 0.0269375
R15348 VDD.n1516 VDD.n1514 0.0269375
R15349 VDD.n1518 VDD.n1516 0.0269375
R15350 VDD.n1520 VDD.n1518 0.0269375
R15351 VDD.n1522 VDD.n1520 0.0269375
R15352 VDD.n1524 VDD.n1522 0.0269375
R15353 VDD.n1528 VDD.n1524 0.0269375
R15354 VDD.n1533 VDD.n1531 0.0269375
R15355 VDD.n1535 VDD.n1533 0.0269375
R15356 VDD.n1537 VDD.n1535 0.0269375
R15357 VDD.n1539 VDD.n1537 0.0269375
R15358 VDD.n1541 VDD.n1539 0.0269375
R15359 VDD.n1543 VDD.n1541 0.0269375
R15360 VDD.n1549 VDD.n1547 0.0269375
R15361 VDD.n1551 VDD.n1549 0.0269375
R15362 VDD.n1553 VDD.n1551 0.0269375
R15363 VDD.n1555 VDD.n1553 0.0269375
R15364 VDD.n1557 VDD.n1555 0.0269375
R15365 VDD.n1559 VDD.n1557 0.0269375
R15366 VDD.n1561 VDD.n1559 0.0269375
R15367 VDD.n1563 VDD.n1561 0.0269375
R15368 VDD.n1565 VDD.n1563 0.0269375
R15369 VDD.n1567 VDD.n1565 0.0269375
R15370 VDD.n1569 VDD.n1567 0.0269375
R15371 VDD.n1571 VDD.n1569 0.0269375
R15372 VDD.n1573 VDD.n1571 0.0269375
R15373 VDD.n1575 VDD.n1573 0.0269375
R15374 VDD.n1577 VDD.n1575 0.0269375
R15375 VDD.n1579 VDD.n1577 0.0269375
R15376 VDD.n1581 VDD.n1579 0.0269375
R15377 VDD.n1583 VDD.n1581 0.0269375
R15378 VDD.n1585 VDD.n1583 0.0269375
R15379 VDD.n1587 VDD.n1585 0.0269375
R15380 VDD.n1589 VDD.n1587 0.0269375
R15381 VDD.n1591 VDD.n1589 0.0269375
R15382 VDD.n1593 VDD.n1591 0.0269375
R15383 VDD.n1595 VDD.n1593 0.0269375
R15384 VDD.n1597 VDD.n1595 0.0269375
R15385 VDD.n1599 VDD.n1597 0.0269375
R15386 VDD.n1601 VDD.n1599 0.0269375
R15387 VDD.n1603 VDD.n1601 0.0269375
R15388 VDD.n1605 VDD.n1603 0.0269375
R15389 VDD.n1607 VDD.n1605 0.0269375
R15390 VDD.n1609 VDD.n1607 0.0269375
R15391 VDD.n1611 VDD.n1609 0.0269375
R15392 VDD.n1613 VDD.n1611 0.0269375
R15393 VDD.n1615 VDD.n1613 0.0269375
R15394 VDD.n1617 VDD.n1615 0.0269375
R15395 VDD.n1619 VDD.n1617 0.0269375
R15396 VDD.n1621 VDD.n1619 0.0269375
R15397 VDD.n1623 VDD.n1621 0.0269375
R15398 VDD.n1625 VDD.n1623 0.0269375
R15399 VDD.n1627 VDD.n1625 0.0269375
R15400 VDD.n1629 VDD.n1627 0.0269375
R15401 VDD.n1631 VDD.n1629 0.0269375
R15402 VDD.n1633 VDD.n1631 0.0269375
R15403 VDD.n1635 VDD.n1633 0.0269375
R15404 VDD.n1637 VDD.n1635 0.0269375
R15405 VDD.n1642 VDD.n1640 0.0269375
R15406 VDD.n1644 VDD.n1642 0.0269375
R15407 VDD.n1646 VDD.n1644 0.0269375
R15408 VDD.n1648 VDD.n1646 0.0269375
R15409 VDD.n1650 VDD.n1648 0.0269375
R15410 VDD.n1652 VDD.n1650 0.0269375
R15411 VDD.n1656 VDD.n1652 0.0269375
R15412 VDD.n1135 VDD.n1133 0.0269375
R15413 VDD.n1137 VDD.n1135 0.0269375
R15414 VDD.n1139 VDD.n1137 0.0269375
R15415 VDD.n1141 VDD.n1139 0.0269375
R15416 VDD.n1143 VDD.n1141 0.0269375
R15417 VDD.n1151 VDD.n1149 0.0269375
R15418 VDD.n1156 VDD.n1154 0.0269375
R15419 VDD.n1158 VDD.n1156 0.0269375
R15420 VDD.n1160 VDD.n1158 0.0269375
R15421 VDD.n1162 VDD.n1160 0.0269375
R15422 VDD.n1164 VDD.n1162 0.0269375
R15423 VDD.n1169 VDD.n1167 0.0269375
R15424 VDD.n1171 VDD.n1169 0.0269375
R15425 VDD.n1173 VDD.n1171 0.0269375
R15426 VDD.n1178 VDD.n1176 0.0269375
R15427 VDD.n1180 VDD.n1178 0.0269375
R15428 VDD.n1182 VDD.n1180 0.0269375
R15429 VDD.n1184 VDD.n1182 0.0269375
R15430 VDD.n1186 VDD.n1184 0.0269375
R15431 VDD.n1188 VDD.n1186 0.0269375
R15432 VDD.n1190 VDD.n1188 0.0269375
R15433 VDD.n1192 VDD.n1190 0.0269375
R15434 VDD.n1194 VDD.n1192 0.0269375
R15435 VDD.n1196 VDD.n1194 0.0269375
R15436 VDD.n1198 VDD.n1196 0.0269375
R15437 VDD.n1200 VDD.n1198 0.0269375
R15438 VDD.n1202 VDD.n1200 0.0269375
R15439 VDD.n1204 VDD.n1202 0.0269375
R15440 VDD.n1206 VDD.n1204 0.0269375
R15441 VDD.n1208 VDD.n1206 0.0269375
R15442 VDD.n1210 VDD.n1208 0.0269375
R15443 VDD.n1212 VDD.n1210 0.0269375
R15444 VDD.n1214 VDD.n1212 0.0269375
R15445 VDD.n1216 VDD.n1214 0.0269375
R15446 VDD.n1218 VDD.n1216 0.0269375
R15447 VDD.n1220 VDD.n1218 0.0269375
R15448 VDD.n1222 VDD.n1220 0.0269375
R15449 VDD.n1230 VDD.n1228 0.0269375
R15450 VDD.n1232 VDD.n1230 0.0269375
R15451 VDD.n1234 VDD.n1232 0.0269375
R15452 VDD.n1236 VDD.n1234 0.0269375
R15453 VDD.n1238 VDD.n1236 0.0269375
R15454 VDD.n2054 VDD.n2051 0.0269375
R15455 VDD.n2057 VDD.n2054 0.0269375
R15456 VDD.n2060 VDD.n2057 0.0269375
R15457 VDD.n2063 VDD.n2060 0.0269375
R15458 VDD.n2066 VDD.n2063 0.0269375
R15459 VDD.n2073 VDD.n2070 0.0269375
R15460 VDD.n2076 VDD.n2073 0.0269375
R15461 VDD.n2079 VDD.n2076 0.0269375
R15462 VDD.n2082 VDD.n2079 0.0269375
R15463 VDD.n2085 VDD.n2082 0.0269375
R15464 VDD.n2088 VDD.n2085 0.0269375
R15465 VDD.n2091 VDD.n2088 0.0269375
R15466 VDD.n2094 VDD.n2091 0.0269375
R15467 VDD.n2097 VDD.n2094 0.0269375
R15468 VDD.n2100 VDD.n2097 0.0269375
R15469 VDD.n2103 VDD.n2100 0.0269375
R15470 VDD.n2106 VDD.n2103 0.0269375
R15471 VDD.n2109 VDD.n2106 0.0269375
R15472 VDD.n2112 VDD.n2109 0.0269375
R15473 VDD.n2115 VDD.n2112 0.0269375
R15474 VDD.n2118 VDD.n2115 0.0269375
R15475 VDD.n2121 VDD.n2118 0.0269375
R15476 VDD.n2124 VDD.n2121 0.0269375
R15477 VDD.n2131 VDD.n2128 0.0269375
R15478 VDD.n2134 VDD.n2131 0.0269375
R15479 VDD.n2137 VDD.n2134 0.0269375
R15480 VDD.n2140 VDD.n2137 0.0269375
R15481 VDD.n2143 VDD.n2140 0.0269375
R15482 VDD.n2151 VDD.n2143 0.0269375
R15483 VDD.n2158 VDD.n2155 0.0269375
R15484 VDD.n2161 VDD.n2158 0.0269375
R15485 VDD.n2164 VDD.n2161 0.0269375
R15486 VDD.n2167 VDD.n2164 0.0269375
R15487 VDD.n2170 VDD.n2167 0.0269375
R15488 VDD.n2173 VDD.n2170 0.0269375
R15489 VDD.n2180 VDD.n2177 0.0269375
R15490 VDD.n2183 VDD.n2180 0.0269375
R15491 VDD.n2186 VDD.n2183 0.0269375
R15492 VDD.n2189 VDD.n2186 0.0269375
R15493 VDD.n2192 VDD.n2189 0.0269375
R15494 VDD.n2195 VDD.n2192 0.0269375
R15495 VDD.n2198 VDD.n2195 0.0269375
R15496 VDD.n2201 VDD.n2198 0.0269375
R15497 VDD.n2204 VDD.n2201 0.0269375
R15498 VDD.n2207 VDD.n2204 0.0269375
R15499 VDD.n2210 VDD.n2207 0.0269375
R15500 VDD.n2213 VDD.n2210 0.0269375
R15501 VDD.n2216 VDD.n2213 0.0269375
R15502 VDD.n2219 VDD.n2216 0.0269375
R15503 VDD.n2222 VDD.n2219 0.0269375
R15504 VDD.n2225 VDD.n2222 0.0269375
R15505 VDD.n2228 VDD.n2225 0.0269375
R15506 VDD.n2231 VDD.n2228 0.0269375
R15507 VDD.n2234 VDD.n2231 0.0269375
R15508 VDD.n2237 VDD.n2234 0.0269375
R15509 VDD.n2240 VDD.n2237 0.0269375
R15510 VDD.n2243 VDD.n2240 0.0269375
R15511 VDD.n2246 VDD.n2243 0.0269375
R15512 VDD.n2249 VDD.n2246 0.0269375
R15513 VDD.n2252 VDD.n2249 0.0269375
R15514 VDD.n2255 VDD.n2252 0.0269375
R15515 VDD.n2258 VDD.n2255 0.0269375
R15516 VDD.n2261 VDD.n2258 0.0269375
R15517 VDD.n2264 VDD.n2261 0.0269375
R15518 VDD.n2267 VDD.n2264 0.0269375
R15519 VDD.n2270 VDD.n2267 0.0269375
R15520 VDD.n2273 VDD.n2270 0.0269375
R15521 VDD.n2276 VDD.n2273 0.0269375
R15522 VDD.n2279 VDD.n2276 0.0269375
R15523 VDD.n2282 VDD.n2279 0.0269375
R15524 VDD.n2285 VDD.n2282 0.0269375
R15525 VDD.n2288 VDD.n2285 0.0269375
R15526 VDD.n2291 VDD.n2288 0.0269375
R15527 VDD.n2294 VDD.n2291 0.0269375
R15528 VDD.n2297 VDD.n2294 0.0269375
R15529 VDD.n2300 VDD.n2297 0.0269375
R15530 VDD.n2303 VDD.n2300 0.0269375
R15531 VDD.n2306 VDD.n2303 0.0269375
R15532 VDD.n2309 VDD.n2306 0.0269375
R15533 VDD.n2312 VDD.n2309 0.0269375
R15534 VDD.n2319 VDD.n2316 0.0269375
R15535 VDD.n2322 VDD.n2319 0.0269375
R15536 VDD.n2325 VDD.n2322 0.0269375
R15537 VDD.n2328 VDD.n2325 0.0269375
R15538 VDD.n2331 VDD.n2328 0.0269375
R15539 VDD.n2334 VDD.n2331 0.0269375
R15540 VDD.n2342 VDD.n2334 0.0269375
R15541 VDD.n2349 VDD.n2346 0.0269375
R15542 VDD.n2352 VDD.n2349 0.0269375
R15543 VDD.n2355 VDD.n2352 0.0269375
R15544 VDD.n2358 VDD.n2355 0.0269375
R15545 VDD.n2361 VDD.n2358 0.0269375
R15546 VDD.n2380 VDD.n2377 0.0269375
R15547 VDD.n2395 VDD.n2392 0.0269375
R15548 VDD.n2402 VDD.n2399 0.0269375
R15549 VDD.n2405 VDD.n2402 0.0269375
R15550 VDD.n2408 VDD.n2405 0.0269375
R15551 VDD.n2416 VDD.n2413 0.0269375
R15552 VDD.n2419 VDD.n2416 0.0269375
R15553 VDD.n2426 VDD.n2423 0.0269375
R15554 VDD.n2433 VDD.n2430 0.0269375
R15555 VDD.n2440 VDD.n2437 0.0269375
R15556 VDD.n2443 VDD.n2440 0.0269375
R15557 VDD.n2451 VDD.n2448 0.0269375
R15558 VDD.n2454 VDD.n2451 0.0269375
R15559 VDD.n2461 VDD.n2458 0.0269375
R15560 VDD.n2468 VDD.n2465 0.0269375
R15561 VDD.n2475 VDD.n2472 0.0269375
R15562 VDD.n2478 VDD.n2475 0.0269375
R15563 VDD.n2489 VDD.n2486 0.0269375
R15564 VDD.n2492 VDD.n2489 0.0269375
R15565 VDD.n2507 VDD.n2504 0.0269375
R15566 VDD.n2510 VDD.n2507 0.0269375
R15567 VDD.n2513 VDD.n2510 0.0269375
R15568 VDD.n2516 VDD.n2513 0.0269375
R15569 VDD.n4361 VDD.n4358 0.0269375
R15570 VDD.n4364 VDD.n4361 0.0269375
R15571 VDD.n4367 VDD.n4364 0.0269375
R15572 VDD.n4370 VDD.n4367 0.0269375
R15573 VDD.n4380 VDD.n4377 0.0269375
R15574 VDD.n4387 VDD.n4384 0.0269375
R15575 VDD.n4390 VDD.n4387 0.0269375
R15576 VDD.n4397 VDD.n4394 0.0269375
R15577 VDD.n4400 VDD.n4397 0.0269375
R15578 VDD.n4407 VDD.n4404 0.0269375
R15579 VDD.n4410 VDD.n4407 0.0269375
R15580 VDD.n4417 VDD.n4414 0.0269375
R15581 VDD.n4420 VDD.n4417 0.0269375
R15582 VDD.n4423 VDD.n4420 0.0269375
R15583 VDD.n4430 VDD.n4427 0.0269375
R15584 VDD.n4433 VDD.n4430 0.0269375
R15585 VDD.n4440 VDD.n4437 0.0269375
R15586 VDD.n4443 VDD.n4440 0.0269375
R15587 VDD.n4446 VDD.n4443 0.0269375
R15588 VDD.n4453 VDD.n4450 0.0269375
R15589 VDD.n4456 VDD.n4453 0.0269375
R15590 VDD.n4463 VDD.n4460 0.0269375
R15591 VDD.n4466 VDD.n4463 0.0269375
R15592 VDD.n4473 VDD.n4470 0.0269375
R15593 VDD.n4476 VDD.n4473 0.0269375
R15594 VDD.n4483 VDD.n4480 0.0269375
R15595 VDD.n4490 VDD.n4487 0.0269375
R15596 VDD.n4493 VDD.n4490 0.0269375
R15597 VDD.n4496 VDD.n4493 0.0269375
R15598 VDD.n4499 VDD.n4496 0.0269375
R15599 VDD.n4536 VDD.n4533 0.0269375
R15600 VDD.n4539 VDD.n4536 0.0269375
R15601 VDD.n4542 VDD.n4539 0.0269375
R15602 VDD.n4549 VDD.n4546 0.0269375
R15603 VDD.n4556 VDD.n4553 0.0269375
R15604 VDD.n4559 VDD.n4556 0.0269375
R15605 VDD.n4566 VDD.n4563 0.0269375
R15606 VDD.n4569 VDD.n4566 0.0269375
R15607 VDD.n4576 VDD.n4573 0.0269375
R15608 VDD.n4579 VDD.n4576 0.0269375
R15609 VDD.n4586 VDD.n4583 0.0269375
R15610 VDD.n4589 VDD.n4586 0.0269375
R15611 VDD.n4592 VDD.n4589 0.0269375
R15612 VDD.n4599 VDD.n4596 0.0269375
R15613 VDD.n4602 VDD.n4599 0.0269375
R15614 VDD.n4609 VDD.n4606 0.0269375
R15615 VDD.n4612 VDD.n4609 0.0269375
R15616 VDD.n4615 VDD.n4612 0.0269375
R15617 VDD.n4622 VDD.n4619 0.0269375
R15618 VDD.n4625 VDD.n4622 0.0269375
R15619 VDD.n4632 VDD.n4629 0.0269375
R15620 VDD.n4635 VDD.n4632 0.0269375
R15621 VDD.n4642 VDD.n4639 0.0269375
R15622 VDD.n4645 VDD.n4642 0.0269375
R15623 VDD.n4652 VDD.n4649 0.0269375
R15624 VDD.n4659 VDD.n4656 0.0269375
R15625 VDD.n4662 VDD.n4659 0.0269375
R15626 VDD.n4665 VDD.n4662 0.0269375
R15627 VDD.n5649 VDD.n5647 0.0269375
R15628 VDD.n5651 VDD.n5649 0.0269375
R15629 VDD.n5653 VDD.n5651 0.0269375
R15630 VDD.n5655 VDD.n5653 0.0269375
R15631 VDD.n5660 VDD.n5658 0.0269375
R15632 VDD.n5665 VDD.n5663 0.0269375
R15633 VDD.n5667 VDD.n5665 0.0269375
R15634 VDD.n5672 VDD.n5670 0.0269375
R15635 VDD.n5674 VDD.n5672 0.0269375
R15636 VDD.n5679 VDD.n5677 0.0269375
R15637 VDD.n5681 VDD.n5679 0.0269375
R15638 VDD.n5686 VDD.n5684 0.0269375
R15639 VDD.n5688 VDD.n5686 0.0269375
R15640 VDD.n5690 VDD.n5688 0.0269375
R15641 VDD.n5692 VDD.n5690 0.0269375
R15642 VDD.n5694 VDD.n5692 0.0269375
R15643 VDD.n5696 VDD.n5694 0.0269375
R15644 VDD.n5698 VDD.n5696 0.0269375
R15645 VDD.n5700 VDD.n5698 0.0269375
R15646 VDD.n5702 VDD.n5700 0.0269375
R15647 VDD.n5704 VDD.n5702 0.0269375
R15648 VDD.n5709 VDD.n5707 0.0269375
R15649 VDD.n5711 VDD.n5709 0.0269375
R15650 VDD.n5716 VDD.n5714 0.0269375
R15651 VDD.n5718 VDD.n5716 0.0269375
R15652 VDD.n5723 VDD.n5721 0.0269375
R15653 VDD.n5725 VDD.n5723 0.0269375
R15654 VDD.n5730 VDD.n5728 0.0269375
R15655 VDD.n5735 VDD.n5733 0.0269375
R15656 VDD.n5737 VDD.n5735 0.0269375
R15657 VDD.n5739 VDD.n5737 0.0269375
R15658 VDD.n5741 VDD.n5739 0.0269375
R15659 VDD.n5755 VDD.n5753 0.0269375
R15660 VDD.n5757 VDD.n5755 0.0269375
R15661 VDD.n5759 VDD.n5757 0.0269375
R15662 VDD.n5761 VDD.n5759 0.0269375
R15663 VDD.n5766 VDD.n5764 0.0269375
R15664 VDD.n5771 VDD.n5769 0.0269375
R15665 VDD.n5773 VDD.n5771 0.0269375
R15666 VDD.n5778 VDD.n5776 0.0269375
R15667 VDD.n5780 VDD.n5778 0.0269375
R15668 VDD.n5785 VDD.n5783 0.0269375
R15669 VDD.n5787 VDD.n5785 0.0269375
R15670 VDD.n5792 VDD.n5790 0.0269375
R15671 VDD.n5794 VDD.n5792 0.0269375
R15672 VDD.n5796 VDD.n5794 0.0269375
R15673 VDD.n5798 VDD.n5796 0.0269375
R15674 VDD.n5800 VDD.n5798 0.0269375
R15675 VDD.n5802 VDD.n5800 0.0269375
R15676 VDD.n5804 VDD.n5802 0.0269375
R15677 VDD.n5806 VDD.n5804 0.0269375
R15678 VDD.n5808 VDD.n5806 0.0269375
R15679 VDD.n5810 VDD.n5808 0.0269375
R15680 VDD.n5815 VDD.n5813 0.0269375
R15681 VDD.n5817 VDD.n5815 0.0269375
R15682 VDD.n5822 VDD.n5820 0.0269375
R15683 VDD.n5824 VDD.n5822 0.0269375
R15684 VDD.n5829 VDD.n5827 0.0269375
R15685 VDD.n5831 VDD.n5829 0.0269375
R15686 VDD.n5836 VDD.n5834 0.0269375
R15687 VDD.n5841 VDD.n5839 0.0269375
R15688 VDD.n5843 VDD.n5841 0.0269375
R15689 VDD.n5845 VDD.n5843 0.0269375
R15690 VDD.n2437 VDD.n2434 0.0266563
R15691 VDD.n5862 VDD.n5860 0.026375
R15692 VDD.n5925 VDD.n5924 0.026375
R15693 VDD.n5970 VDD.n5968 0.026375
R15694 VDD.n6033 VDD.n6032 0.026375
R15695 VDD.n4700 VDD.n4697 0.026375
R15696 VDD.n4793 VDD.n4792 0.026375
R15697 VDD.n4855 VDD.n4852 0.026375
R15698 VDD.n4948 VDD.n4947 0.026375
R15699 VDD.n6068 VDD.n6066 0.026375
R15700 VDD.n6131 VDD.n6130 0.026375
R15701 VDD.n6290 VDD.n6289 0.026375
R15702 VDD.n6227 VDD.n6225 0.026375
R15703 VDD.n5002 VDD.n4999 0.026375
R15704 VDD.n5095 VDD.n5094 0.026375
R15705 VDD.n5157 VDD.n5154 0.026375
R15706 VDD.n5250 VDD.n5249 0.026375
R15707 VDD.n2598 VDD.n2596 0.026375
R15708 VDD.n2661 VDD.n2660 0.026375
R15709 VDD.n6479 VDD.n6476 0.026375
R15710 VDD.n6572 VDD.n6571 0.026375
R15711 VDD.n870 VDD.n869 0.026375
R15712 VDD.n4384 VDD.n4381 0.026375
R15713 VDD.n4477 VDD.n4476 0.026375
R15714 VDD.n4553 VDD.n4550 0.026375
R15715 VDD.n4646 VDD.n4645 0.026375
R15716 VDD.n5663 VDD.n5661 0.026375
R15717 VDD.n5726 VDD.n5725 0.026375
R15718 VDD.n5769 VDD.n5767 0.026375
R15719 VDD.n5832 VDD.n5831 0.026375
R15720 VDD.n1147 VDD.n1146 0.0260938
R15721 VDD.n1225 VDD.n1223 0.0260938
R15722 VDD.n2366 VDD.n2365 0.0260938
R15723 VDD.n2384 VDD.n2381 0.0260938
R15724 VDD.n2462 VDD.n2461 0.0260938
R15725 VDD.n2496 VDD.n2493 0.0260938
R15726 VDD.n4674 VDD.n4673 0.0258125
R15727 VDD.n390 VDD.n389 0.0258125
R15728 VDD.n4520 VDD.n4519 0.0258125
R15729 VDD.n1462 VDD.n1460 0.0249687
R15730 VDD.n1531 VDD.n1529 0.0249687
R15731 VDD.n1242 VDD.n1238 0.0249687
R15732 VDD.n2051 VDD.n2048 0.0249687
R15733 VDD.n2155 VDD.n2152 0.0249687
R15734 VDD.n2346 VDD.n2343 0.0249687
R15735 VDD.n2533 VDD.n2516 0.0249687
R15736 VDD.n5869 VDD.n5867 0.0246875
R15737 VDD.n5918 VDD.n5917 0.0246875
R15738 VDD.n5977 VDD.n5975 0.0246875
R15739 VDD.n6026 VDD.n6025 0.0246875
R15740 VDD.n4710 VDD.n4707 0.0246875
R15741 VDD.n4783 VDD.n4782 0.0246875
R15742 VDD.n4865 VDD.n4862 0.0246875
R15743 VDD.n4938 VDD.n4937 0.0246875
R15744 VDD.n6075 VDD.n6073 0.0246875
R15745 VDD.n6124 VDD.n6123 0.0246875
R15746 VDD.n6283 VDD.n6282 0.0246875
R15747 VDD.n6234 VDD.n6232 0.0246875
R15748 VDD.n5012 VDD.n5009 0.0246875
R15749 VDD.n5085 VDD.n5084 0.0246875
R15750 VDD.n5167 VDD.n5164 0.0246875
R15751 VDD.n5240 VDD.n5239 0.0246875
R15752 VDD.n2605 VDD.n2603 0.0246875
R15753 VDD.n2654 VDD.n2653 0.0246875
R15754 VDD.n6489 VDD.n6486 0.0246875
R15755 VDD.n6562 VDD.n6561 0.0246875
R15756 VDD.n439 VDD.n438 0.0246875
R15757 VDD.n8016 VDD.n8014 0.0246875
R15758 VDD.n7915 VDD.n7912 0.0246875
R15759 VDD.n8138 VDD.n8135 0.0246875
R15760 VDD.n8177 VDD.n8176 0.0246875
R15761 VDD.n4394 VDD.n4391 0.0246875
R15762 VDD.n4467 VDD.n4466 0.0246875
R15763 VDD.n4563 VDD.n4560 0.0246875
R15764 VDD.n4636 VDD.n4635 0.0246875
R15765 VDD.n5670 VDD.n5668 0.0246875
R15766 VDD.n5719 VDD.n5718 0.0246875
R15767 VDD.n5776 VDD.n5774 0.0246875
R15768 VDD.n5825 VDD.n5824 0.0246875
R15769 VDD.n3267 VDD.n3265 0.024264
R15770 VDD.n3270 VDD.n3267 0.024264
R15771 VDD.n3272 VDD.n3270 0.024264
R15772 VDD.n3275 VDD.n3272 0.024264
R15773 VDD.n3277 VDD.n3275 0.024264
R15774 VDD.n3280 VDD.n3277 0.024264
R15775 VDD.n3282 VDD.n3280 0.024264
R15776 VDD.n3285 VDD.n3282 0.024264
R15777 VDD.n3287 VDD.n3285 0.024264
R15778 VDD.n3290 VDD.n3287 0.024264
R15779 VDD.n3292 VDD.n3290 0.024264
R15780 VDD.n3295 VDD.n3292 0.024264
R15781 VDD.n3297 VDD.n3295 0.024264
R15782 VDD.n3300 VDD.n3297 0.024264
R15783 VDD.n3302 VDD.n3300 0.024264
R15784 VDD.n3305 VDD.n3302 0.024264
R15785 VDD.n3307 VDD.n3305 0.024264
R15786 VDD.n3310 VDD.n3307 0.024264
R15787 VDD.n3312 VDD.n3310 0.024264
R15788 VDD.n3315 VDD.n3312 0.024264
R15789 VDD.n3317 VDD.n3315 0.024264
R15790 VDD.n3320 VDD.n3317 0.024264
R15791 VDD.n3322 VDD.n3320 0.024264
R15792 VDD.n3325 VDD.n3322 0.024264
R15793 VDD.n3327 VDD.n3325 0.024264
R15794 VDD.n3330 VDD.n3327 0.024264
R15795 VDD.n3332 VDD.n3330 0.024264
R15796 VDD.n3335 VDD.n3332 0.024264
R15797 VDD.n3337 VDD.n3335 0.024264
R15798 VDD.n3340 VDD.n3337 0.024264
R15799 VDD.n3342 VDD.n3340 0.024264
R15800 VDD.n3345 VDD.n3342 0.024264
R15801 VDD.n3347 VDD.n3345 0.024264
R15802 VDD.n3350 VDD.n3347 0.024264
R15803 VDD.n3352 VDD.n3350 0.024264
R15804 VDD.n3355 VDD.n3352 0.024264
R15805 VDD.n3357 VDD.n3355 0.024264
R15806 VDD.n3360 VDD.n3357 0.024264
R15807 VDD.n3362 VDD.n3360 0.024264
R15808 VDD.n3365 VDD.n3362 0.024264
R15809 VDD.n3367 VDD.n3365 0.024264
R15810 VDD.n3370 VDD.n3367 0.024264
R15811 VDD.n3372 VDD.n3370 0.024264
R15812 VDD.n3375 VDD.n3372 0.024264
R15813 VDD.n3377 VDD.n3375 0.024264
R15814 VDD.n3380 VDD.n3377 0.024264
R15815 VDD.n3382 VDD.n3380 0.024264
R15816 VDD.n3385 VDD.n3382 0.024264
R15817 VDD.n5487 VDD.n5485 0.024264
R15818 VDD.n3772 VDD.n3770 0.024264
R15819 VDD.n3775 VDD.n3772 0.024264
R15820 VDD.n3777 VDD.n3775 0.024264
R15821 VDD.n3780 VDD.n3777 0.024264
R15822 VDD.n3782 VDD.n3780 0.024264
R15823 VDD.n3785 VDD.n3782 0.024264
R15824 VDD.n3787 VDD.n3785 0.024264
R15825 VDD.n3790 VDD.n3787 0.024264
R15826 VDD.n3792 VDD.n3790 0.024264
R15827 VDD.n3795 VDD.n3792 0.024264
R15828 VDD.n3797 VDD.n3795 0.024264
R15829 VDD.n3800 VDD.n3797 0.024264
R15830 VDD.n3802 VDD.n3800 0.024264
R15831 VDD.n3805 VDD.n3802 0.024264
R15832 VDD.n3807 VDD.n3805 0.024264
R15833 VDD.n3810 VDD.n3807 0.024264
R15834 VDD.n3812 VDD.n3810 0.024264
R15835 VDD.n3815 VDD.n3812 0.024264
R15836 VDD.n3817 VDD.n3815 0.024264
R15837 VDD.n3820 VDD.n3817 0.024264
R15838 VDD.n3822 VDD.n3820 0.024264
R15839 VDD.n3825 VDD.n3822 0.024264
R15840 VDD.n3827 VDD.n3825 0.024264
R15841 VDD.n3830 VDD.n3827 0.024264
R15842 VDD.n3832 VDD.n3830 0.024264
R15843 VDD.n3835 VDD.n3832 0.024264
R15844 VDD.n3837 VDD.n3835 0.024264
R15845 VDD.n3840 VDD.n3837 0.024264
R15846 VDD.n3842 VDD.n3840 0.024264
R15847 VDD.n3845 VDD.n3842 0.024264
R15848 VDD.n3847 VDD.n3845 0.024264
R15849 VDD.n3850 VDD.n3847 0.024264
R15850 VDD.n3852 VDD.n3850 0.024264
R15851 VDD.n3855 VDD.n3852 0.024264
R15852 VDD.n3857 VDD.n3855 0.024264
R15853 VDD.n3860 VDD.n3857 0.024264
R15854 VDD.n3862 VDD.n3860 0.024264
R15855 VDD.n3865 VDD.n3862 0.024264
R15856 VDD.n3867 VDD.n3865 0.024264
R15857 VDD.n3870 VDD.n3867 0.024264
R15858 VDD.n3872 VDD.n3870 0.024264
R15859 VDD.n3875 VDD.n3872 0.024264
R15860 VDD.n3877 VDD.n3875 0.024264
R15861 VDD.n3880 VDD.n3877 0.024264
R15862 VDD.n3882 VDD.n3880 0.024264
R15863 VDD.n3885 VDD.n3882 0.024264
R15864 VDD.n6324 VDD.n6321 0.024264
R15865 VDD.n6327 VDD.n6324 0.024264
R15866 VDD.n6330 VDD.n6327 0.024264
R15867 VDD.n6332 VDD.n6330 0.024264
R15868 VDD.n6335 VDD.n6332 0.024264
R15869 VDD.n6337 VDD.n6335 0.024264
R15870 VDD.n6340 VDD.n6337 0.024264
R15871 VDD.n6342 VDD.n6340 0.024264
R15872 VDD.n6345 VDD.n6342 0.024264
R15873 VDD.n6347 VDD.n6345 0.024264
R15874 VDD.n6350 VDD.n6347 0.024264
R15875 VDD.n6352 VDD.n6350 0.024264
R15876 VDD.n6355 VDD.n6352 0.024264
R15877 VDD.n6357 VDD.n6355 0.024264
R15878 VDD.n6360 VDD.n6357 0.024264
R15879 VDD.n6362 VDD.n6360 0.024264
R15880 VDD.n6365 VDD.n6362 0.024264
R15881 VDD.n6367 VDD.n6365 0.024264
R15882 VDD.n6370 VDD.n6367 0.024264
R15883 VDD.n6372 VDD.n6370 0.024264
R15884 VDD.n6375 VDD.n6372 0.024264
R15885 VDD.n6377 VDD.n6375 0.024264
R15886 VDD.n6380 VDD.n6377 0.024264
R15887 VDD.n6382 VDD.n6380 0.024264
R15888 VDD.n6385 VDD.n6382 0.024264
R15889 VDD.n6387 VDD.n6385 0.024264
R15890 VDD.n6390 VDD.n6387 0.024264
R15891 VDD.n6392 VDD.n6390 0.024264
R15892 VDD.n6395 VDD.n6392 0.024264
R15893 VDD.n6397 VDD.n6395 0.024264
R15894 VDD.n6400 VDD.n6397 0.024264
R15895 VDD.n6402 VDD.n6400 0.024264
R15896 VDD.n6405 VDD.n6402 0.024264
R15897 VDD.n6407 VDD.n6405 0.024264
R15898 VDD.n6410 VDD.n6407 0.024264
R15899 VDD.n6412 VDD.n6410 0.024264
R15900 VDD.n6415 VDD.n6412 0.024264
R15901 VDD.n6417 VDD.n6415 0.024264
R15902 VDD.n6420 VDD.n6417 0.024264
R15903 VDD.n6422 VDD.n6420 0.024264
R15904 VDD.n6425 VDD.n6422 0.024264
R15905 VDD.n6427 VDD.n6425 0.024264
R15906 VDD.n6430 VDD.n6427 0.024264
R15907 VDD.n6432 VDD.n6430 0.024264
R15908 VDD.n6436 VDD.n6432 0.024264
R15909 VDD.n6439 VDD.n6436 0.024264
R15910 VDD.n6441 VDD.n6439 0.024264
R15911 VDD.n6444 VDD.n6441 0.024264
R15912 VDD.n6447 VDD.n6444 0.024264
R15913 VDD.n5881 VDD.n5880 0.024125
R15914 VDD.n5906 VDD.n5904 0.024125
R15915 VDD.n5989 VDD.n5988 0.024125
R15916 VDD.n6014 VDD.n6012 0.024125
R15917 VDD.n4727 VDD.n4726 0.024125
R15918 VDD.n4766 VDD.n4763 0.024125
R15919 VDD.n4882 VDD.n4881 0.024125
R15920 VDD.n4921 VDD.n4918 0.024125
R15921 VDD.n6087 VDD.n6086 0.024125
R15922 VDD.n6112 VDD.n6110 0.024125
R15923 VDD.n6271 VDD.n6269 0.024125
R15924 VDD.n6246 VDD.n6245 0.024125
R15925 VDD.n5029 VDD.n5028 0.024125
R15926 VDD.n5068 VDD.n5065 0.024125
R15927 VDD.n5184 VDD.n5183 0.024125
R15928 VDD.n5223 VDD.n5220 0.024125
R15929 VDD.n2617 VDD.n2616 0.024125
R15930 VDD.n2642 VDD.n2640 0.024125
R15931 VDD.n6506 VDD.n6505 0.024125
R15932 VDD.n6545 VDD.n6542 0.024125
R15933 VDD.n4411 VDD.n4410 0.024125
R15934 VDD.n4450 VDD.n4447 0.024125
R15935 VDD.n4580 VDD.n4579 0.024125
R15936 VDD.n4619 VDD.n4616 0.024125
R15937 VDD.n5682 VDD.n5681 0.024125
R15938 VDD.n5707 VDD.n5705 0.024125
R15939 VDD.n5788 VDD.n5787 0.024125
R15940 VDD.n5813 VDD.n5811 0.024125
R15941 VDD.n8253 VDD.n8251 0.023
R15942 VDD.n7585 VDD.n7583 0.023
R15943 VDD.n7719 VDD.n7718 0.023
R15944 VDD.n1473 VDD.n1472 0.0227188
R15945 VDD.n1640 VDD.n1638 0.0227188
R15946 VDD.n2067 VDD.n2066 0.0227188
R15947 VDD.n2316 VDD.n2313 0.0227188
R15948 VDD.n2455 VDD.n2454 0.0221563
R15949 VDD.n5954 VDD.n5952 0.021875
R15950 VDD.n4816 VDD.n4815 0.021875
R15951 VDD.n6147 VDD.n6146 0.021875
R15952 VDD.n6306 VDD.n6305 0.021875
R15953 VDD.n5118 VDD.n5117 0.021875
R15954 VDD.n2685 VDD.n2681 0.021875
R15955 VDD.n6600 VDD.n6594 0.021875
R15956 VDD.n4358 VDD.n4355 0.021875
R15957 VDD.n4500 VDD.n4499 0.021875
R15958 VDD.n4529 VDD.n4526 0.021875
R15959 VDD.n5647 VDD.n5645 0.021875
R15960 VDD.n5742 VDD.n5741 0.021875
R15961 VDD.n5753 VDD.n5751 0.021875
R15962 VDD.n1165 VDD.n1164 0.0215938
R15963 VDD.n1176 VDD.n1174 0.0215938
R15964 VDD.n2396 VDD.n2395 0.0215938
R15965 VDD.n2413 VDD.n2410 0.0215938
R15966 VDD.n893 VDD.n891 0.0213125
R15967 VDD.n584 VDD.n582 0.0213125
R15968 VDD.n6659 VDD.n6657 0.0213125
R15969 VDD.n6703 VDD.n6701 0.0213125
R15970 VDD.n7954 VDD.n7953 0.0213125
R15971 VDD.n1075 VDD.n1072 0.0213125
R15972 VDD.n775 VDD.n772 0.0213125
R15973 VDD.n809 VDD.n806 0.0213125
R15974 VDD.n6636 VDD.n6635 0.0213125
R15975 VDD.n2472 VDD.n2469 0.0210313
R15976 VDD.n4829 VDD.n4828 0.02075
R15977 VDD.n903 VDD.n902 0.0201875
R15978 VDD.n594 VDD.n593 0.0201875
R15979 VDD.n146 VDD.n143 0.0201875
R15980 VDD.n206 VDD.n205 0.0201875
R15981 VDD.n6989 VDD.n6986 0.0201875
R15982 VDD.n7052 VDD.n7051 0.0201875
R15983 VDD.n1089 VDD.n1088 0.0201875
R15984 VDD.n5846 VDD.n5487 0.0199663
R15985 VDD.n6321 VDD.n6319 0.0199663
R15986 VDD.n6456 VDD.n6447 0.0199663
R15987 VDD.n1146 VDD.n1144 0.0199062
R15988 VDD.n1226 VDD.n1225 0.0199062
R15989 VDD.n2365 VDD.n2362 0.0199062
R15990 VDD.n2497 VDD.n2496 0.0199062
R15991 VDD.n213 VDD.n211 0.0197857
R15992 VDD.n139 VDD.n138 0.0197857
R15993 VDD.n2486 VDD.n2483 0.0193437
R15994 VDD.n4743 VDD.n4740 0.0190625
R15995 VDD.n4750 VDD.n4749 0.0190625
R15996 VDD.n4898 VDD.n4895 0.0190625
R15997 VDD.n4905 VDD.n4904 0.0190625
R15998 VDD.n5045 VDD.n5042 0.0190625
R15999 VDD.n5052 VDD.n5051 0.0190625
R16000 VDD.n5200 VDD.n5197 0.0190625
R16001 VDD.n5207 VDD.n5206 0.0190625
R16002 VDD.n6522 VDD.n6519 0.0190625
R16003 VDD.n6529 VDD.n6528 0.0190625
R16004 VDD.n8324 VDD.n8316 0.0190625
R16005 VDD.n330 VDD.n329 0.0190625
R16006 VDD.n386 VDD.n383 0.0190625
R16007 VDD.n8200 VDD.n8198 0.0190625
R16008 VDD.n4427 VDD.n4424 0.0190625
R16009 VDD.n4434 VDD.n4433 0.0190625
R16010 VDD.n4596 VDD.n4593 0.0190625
R16011 VDD.n4603 VDD.n4602 0.0190625
R16012 VDD.n1514 VDD.n1512 0.0187812
R16013 VDD.n2128 VDD.n2125 0.0187812
R16014 VDD.n2389 VDD.n2388 0.0187812
R16015 VDD.n5857 VDD.n5855 0.0185
R16016 VDD.n5930 VDD.n5929 0.0185
R16017 VDD.n5965 VDD.n5963 0.0185
R16018 VDD.n6043 VDD.n6037 0.0185
R16019 VDD.n4693 VDD.n4690 0.0185
R16020 VDD.n4800 VDD.n4799 0.0185
R16021 VDD.n4848 VDD.n4845 0.0185
R16022 VDD.n4955 VDD.n4954 0.0185
R16023 VDD.n6063 VDD.n6061 0.0185
R16024 VDD.n6136 VDD.n6135 0.0185
R16025 VDD.n6295 VDD.n6294 0.0185
R16026 VDD.n6222 VDD.n6220 0.0185
R16027 VDD.n4995 VDD.n4992 0.0185
R16028 VDD.n5102 VDD.n5101 0.0185
R16029 VDD.n5150 VDD.n5147 0.0185
R16030 VDD.n5257 VDD.n5256 0.0185
R16031 VDD.n2593 VDD.n2591 0.0185
R16032 VDD.n2671 VDD.n2665 0.0185
R16033 VDD.n6472 VDD.n6469 0.0185
R16034 VDD.n6579 VDD.n6578 0.0185
R16035 VDD.n7605 VDD.n7604 0.0185
R16036 VDD.n7699 VDD.n7697 0.0185
R16037 VDD.n4377 VDD.n4374 0.0185
R16038 VDD.n4484 VDD.n4483 0.0185
R16039 VDD.n4546 VDD.n4543 0.0185
R16040 VDD.n4653 VDD.n4652 0.0185
R16041 VDD.n5658 VDD.n5656 0.0185
R16042 VDD.n5731 VDD.n5730 0.0185
R16043 VDD.n5764 VDD.n5762 0.0185
R16044 VDD.n5837 VDD.n5836 0.0185
R16045 VDD.n1154 VDD.n1152 0.0182187
R16046 VDD.n2377 VDD.n2374 0.0182187
R16047 VDD.n2430 VDD.n2427 0.0182187
R16048 VDD.n7394 VDD.n7391 0.0179793
R16049 VDD.n900 VDD.n898 0.0179375
R16050 VDD.n591 VDD.n589 0.0179375
R16051 VDD.n150 VDD.n149 0.0179375
R16052 VDD.n202 VDD.n199 0.0179375
R16053 VDD.n6993 VDD.n6992 0.0179375
R16054 VDD.n7048 VDD.n7045 0.0179375
R16055 VDD.n1085 VDD.n1082 0.0179375
R16056 VDD.n4533 VDD.n4530 0.0179375
R16057 VDD.n1545 VDD.n1543 0.0170938
R16058 VDD.n2174 VDD.n2173 0.0170938
R16059 VDD.n2373 VDD.n2370 0.0170938
R16060 VDD.n2479 VDD.n2478 0.0170938
R16061 VDD.n2388 VDD.n2385 0.0165313
R16062 VDD.n2420 VDD.n2419 0.0165313
R16063 VDD.n2501 VDD.n2500 0.0165313
R16064 VDD.n4822 VDD.n4821 0.0156875
R16065 VDD.n4976 VDD.n4975 0.0156875
R16066 VDD.n7038 VDD.n7037 0.015125
R16067 VDD.n7199 VDD.n7198 0.0145625
R16068 VDD.n7944 VDD.n7941 0.0145625
R16069 VDD.n7071 VDD.n7069 0.0145625
R16070 VDD.n5876 VDD.n5874 0.014
R16071 VDD.n5911 VDD.n5910 0.014
R16072 VDD.n5984 VDD.n5982 0.014
R16073 VDD.n6019 VDD.n6018 0.014
R16074 VDD.n4720 VDD.n4717 0.014
R16075 VDD.n4773 VDD.n4772 0.014
R16076 VDD.n4875 VDD.n4872 0.014
R16077 VDD.n4928 VDD.n4927 0.014
R16078 VDD.n6082 VDD.n6080 0.014
R16079 VDD.n6117 VDD.n6116 0.014
R16080 VDD.n6276 VDD.n6275 0.014
R16081 VDD.n6241 VDD.n6239 0.014
R16082 VDD.n5022 VDD.n5019 0.014
R16083 VDD.n5075 VDD.n5074 0.014
R16084 VDD.n5177 VDD.n5174 0.014
R16085 VDD.n5230 VDD.n5229 0.014
R16086 VDD.n2612 VDD.n2610 0.014
R16087 VDD.n2647 VDD.n2646 0.014
R16088 VDD.n6499 VDD.n6496 0.014
R16089 VDD.n6552 VDD.n6551 0.014
R16090 VDD.n6982 VDD.n6981 0.014
R16091 VDD.n6854 VDD.n6853 0.014
R16092 VDD.n4404 VDD.n4401 0.014
R16093 VDD.n4457 VDD.n4456 0.014
R16094 VDD.n4573 VDD.n4570 0.014
R16095 VDD.n4626 VDD.n4625 0.014
R16096 VDD.n5677 VDD.n5675 0.014
R16097 VDD.n5712 VDD.n5711 0.014
R16098 VDD.n5783 VDD.n5781 0.014
R16099 VDD.n5818 VDD.n5817 0.014
R16100 VDD.n5874 VDD.n5873 0.0134375
R16101 VDD.n5913 VDD.n5911 0.0134375
R16102 VDD.n5982 VDD.n5981 0.0134375
R16103 VDD.n6021 VDD.n6019 0.0134375
R16104 VDD.n4717 VDD.n4716 0.0134375
R16105 VDD.n4776 VDD.n4773 0.0134375
R16106 VDD.n4872 VDD.n4871 0.0134375
R16107 VDD.n4931 VDD.n4928 0.0134375
R16108 VDD.n6080 VDD.n6079 0.0134375
R16109 VDD.n6119 VDD.n6117 0.0134375
R16110 VDD.n6278 VDD.n6276 0.0134375
R16111 VDD.n6239 VDD.n6238 0.0134375
R16112 VDD.n5019 VDD.n5018 0.0134375
R16113 VDD.n5078 VDD.n5075 0.0134375
R16114 VDD.n5174 VDD.n5173 0.0134375
R16115 VDD.n5233 VDD.n5230 0.0134375
R16116 VDD.n2610 VDD.n2609 0.0134375
R16117 VDD.n2649 VDD.n2647 0.0134375
R16118 VDD.n6496 VDD.n6495 0.0134375
R16119 VDD.n6555 VDD.n6552 0.0134375
R16120 VDD.n344 VDD.n341 0.0134375
R16121 VDD.n7006 VDD.n7003 0.0134375
R16122 VDD.n4401 VDD.n4400 0.0134375
R16123 VDD.n4460 VDD.n4457 0.0134375
R16124 VDD.n4570 VDD.n4569 0.0134375
R16125 VDD.n4629 VDD.n4626 0.0134375
R16126 VDD.n5675 VDD.n5674 0.0134375
R16127 VDD.n5714 VDD.n5712 0.0134375
R16128 VDD.n5781 VDD.n5780 0.0134375
R16129 VDD.n5820 VDD.n5818 0.0134375
R16130 VDD.n8186 VDD.n8184 0.012875
R16131 VDD.n1027 VDD.n1008 0.0124871
R16132 VDD.n5941 VDD.n5940 0.01175
R16133 VDD.n4979 VDD.n4976 0.01175
R16134 VDD.n5134 VDD.n5131 0.01175
R16135 VDD.n6714 VDD.n6712 0.01175
R16136 VDD.n6853 VDD.n6851 0.01175
R16137 VDD.n602 VDD.n600 0.01175
R16138 VDD.n795 VDD.n737 0.01175
R16139 VDD.n910 VDD.n908 0.01175
R16140 VDD.n8297 VDD.n8285 0.01175
R16141 VDD.n8215 VDD.n8213 0.01175
R16142 VDD.n7179 VDD.n302 0.01175
R16143 VDD.n6981 VDD.n6979 0.01175
R16144 VDD.n7179 VDD.n7165 0.01175
R16145 VDD.n7085 VDD.n7083 0.01175
R16146 VDD.n1096 VDD.n1027 0.01175
R16147 VDD.n7641 VDD.n7537 0.011657
R16148 VDD.n2444 VDD.n2443 0.0114688
R16149 VDD.n884 VDD.n883 0.0111875
R16150 VDD.n575 VDD.n574 0.0111875
R16151 VDD.n1062 VDD.n1061 0.0111875
R16152 VDD.n762 VDD.n761 0.0111875
R16153 VDD.n2385 VDD.n2384 0.0109063
R16154 VDD.n2423 VDD.n2420 0.0109063
R16155 VDD.n2504 VDD.n2501 0.0109063
R16156 VDD.n5942 VDD.n5941 0.010625
R16157 VDD.n5131 VDD.n5130 0.010625
R16158 VDD.n7844 VDD.n7841 0.010625
R16159 VDD.n7342 VDD.n7340 0.010625
R16160 VDD.n1547 VDD.n1545 0.0103438
R16161 VDD.n2177 VDD.n2174 0.0103438
R16162 VDD.n2370 VDD.n2369 0.0103438
R16163 VDD.n2482 VDD.n2479 0.0103438
R16164 VDD.n2448 VDD.n2445 0.00978125
R16165 VDD.n7828 VDD.n7826 0.0095
R16166 VDD.n7886 VDD.n7849 0.0095
R16167 VDD.n7334 VDD.n7333 0.0095
R16168 VDD.n7572 VDD.n7570 0.0095
R16169 VDD.n7732 VDD.n7731 0.0095
R16170 VDD.n4530 VDD.n4529 0.0095
R16171 VDD.n1152 VDD.n1151 0.00921875
R16172 VDD.n2374 VDD.n2373 0.00921875
R16173 VDD.n2427 VDD.n2426 0.00921875
R16174 VDD.n5855 VDD.n5854 0.0089375
R16175 VDD.n5932 VDD.n5930 0.0089375
R16176 VDD.n5963 VDD.n5962 0.0089375
R16177 VDD.n6045 VDD.n6043 0.0089375
R16178 VDD.n4690 VDD.n4689 0.0089375
R16179 VDD.n4803 VDD.n4800 0.0089375
R16180 VDD.n4845 VDD.n4844 0.0089375
R16181 VDD.n4958 VDD.n4955 0.0089375
R16182 VDD.n6061 VDD.n6060 0.0089375
R16183 VDD.n6138 VDD.n6136 0.0089375
R16184 VDD.n6297 VDD.n6295 0.0089375
R16185 VDD.n6220 VDD.n6214 0.0089375
R16186 VDD.n4992 VDD.n4991 0.0089375
R16187 VDD.n5105 VDD.n5102 0.0089375
R16188 VDD.n5147 VDD.n5146 0.0089375
R16189 VDD.n5260 VDD.n5257 0.0089375
R16190 VDD.n2591 VDD.n2590 0.0089375
R16191 VDD.n2673 VDD.n2671 0.0089375
R16192 VDD.n6469 VDD.n6468 0.0089375
R16193 VDD.n6582 VDD.n6579 0.0089375
R16194 VDD.n444 VDD.n443 0.0089375
R16195 VDD.n8021 VDD.n8020 0.0089375
R16196 VDD.n8131 VDD.n8128 0.0089375
R16197 VDD.n4374 VDD.n4370 0.0089375
R16198 VDD.n4487 VDD.n4484 0.0089375
R16199 VDD.n4543 VDD.n4542 0.0089375
R16200 VDD.n4656 VDD.n4653 0.0089375
R16201 VDD.n5656 VDD.n5655 0.0089375
R16202 VDD.n5733 VDD.n5731 0.0089375
R16203 VDD.n5762 VDD.n5761 0.0089375
R16204 VDD.n5839 VDD.n5837 0.0089375
R16205 VDD.n1512 VDD.n1511 0.00865625
R16206 VDD.n2125 VDD.n2124 0.00865625
R16207 VDD.n2392 VDD.n2389 0.00865625
R16208 VDD.n4740 VDD.n4739 0.008375
R16209 VDD.n4753 VDD.n4750 0.008375
R16210 VDD.n4895 VDD.n4894 0.008375
R16211 VDD.n4908 VDD.n4905 0.008375
R16212 VDD.n5042 VDD.n5041 0.008375
R16213 VDD.n5055 VDD.n5052 0.008375
R16214 VDD.n5197 VDD.n5196 0.008375
R16215 VDD.n5210 VDD.n5207 0.008375
R16216 VDD.n6519 VDD.n6518 0.008375
R16217 VDD.n6532 VDD.n6529 0.008375
R16218 VDD.n544 VDD.n532 0.008375
R16219 VDD.n455 VDD.n452 0.008375
R16220 VDD.n8118 VDD.n8109 0.008375
R16221 VDD.n8032 VDD.n8029 0.008375
R16222 VDD.n4424 VDD.n4423 0.008375
R16223 VDD.n4437 VDD.n4434 0.008375
R16224 VDD.n4593 VDD.n4592 0.008375
R16225 VDD.n4606 VDD.n4603 0.008375
R16226 VDD.n2483 VDD.n2482 0.00809375
R16227 VDD.n7928 VDD.n7927 0.0078125
R16228 VDD.n8168 VDD.n8166 0.0078125
R16229 VDD.n1144 VDD.n1143 0.00753125
R16230 VDD.n1228 VDD.n1226 0.00753125
R16231 VDD.n2362 VDD.n2361 0.00753125
R16232 VDD.n2500 VDD.n2497 0.00753125
R16233 VDD.n2445 VDD.n2444 0.0066875
R16234 VDD.n2469 VDD.n2468 0.00640625
R16235 VDD.n1167 VDD.n1165 0.00584375
R16236 VDD.n1174 VDD.n1173 0.00584375
R16237 VDD.n2399 VDD.n2396 0.00584375
R16238 VDD.n5947 VDD.n5942 0.0055625
R16239 VDD.n5952 VDD.n5951 0.0055625
R16240 VDD.n4821 VDD.n4816 0.0055625
R16241 VDD.n4828 VDD.n4827 0.0055625
R16242 VDD.n6151 VDD.n6147 0.0055625
R16243 VDD.n6306 VDD.n6155 0.0055625
R16244 VDD.n5123 VDD.n5118 0.0055625
R16245 VDD.n5124 VDD.n5123 0.0055625
R16246 VDD.n5130 VDD.n5129 0.0055625
R16247 VDD.n6600 VDD.n6599 0.0055625
R16248 VDD.n6654 VDD.n6652 0.0055625
R16249 VDD.n6708 VDD.n6707 0.0055625
R16250 VDD.n8142 VDD.n8139 0.0055625
R16251 VDD.n802 VDD.n799 0.0055625
R16252 VDD.n6643 VDD.n6642 0.0055625
R16253 VDD.n2410 VDD.n2409 0.0055625
R16254 VDD.n4519 VDD.n4500 0.0055625
R16255 VDD.n4526 VDD.n4525 0.0055625
R16256 VDD.n5746 VDD.n5742 0.0055625
R16257 VDD.n5751 VDD.n5750 0.0055625
R16258 VDD.n2458 VDD.n2455 0.00528125
R16259 VDD.n6052 VDD.n5346 0.00479775
R16260 VDD.n5846 VDD.n5483 0.00479775
R16261 VDD.n6319 VDD.n6314 0.00479775
R16262 VDD.n6456 VDD.n6455 0.00479775
R16263 VDD.n1475 VDD.n1473 0.00471875
R16264 VDD.n1638 VDD.n1637 0.00471875
R16265 VDD.n2070 VDD.n2067 0.00471875
R16266 VDD.n2313 VDD.n2312 0.00471875
R16267 VDD.n5645 VDD.n5641 0.00359375
R16268 VDD.n4355 VDD.n4350 0.00359375
R16269 VDD.n5742 VDD.n5571 0.00359375
R16270 VDD.n4500 VDD.n4177 0.00359375
R16271 VDD.n5952 VDD.n5410 0.00359375
R16272 VDD.n4828 VDD.n3586 0.00359375
R16273 VDD.n5751 VDD.n5561 0.00359375
R16274 VDD.n4526 VDD.n4081 0.00359375
R16275 VDD.n5942 VDD.n5418 0.00359375
R16276 VDD.n4816 VDD.n3699 0.00359375
R16277 VDD.n6147 VDD.n5281 0.00359375
R16278 VDD.n5118 VDD.n3195 0.00359375
R16279 VDD.n6306 VDD.n5275 0.00359375
R16280 VDD.n5130 VDD.n3079 0.00359375
R16281 VDD.n2687 VDD.n2685 0.00359375
R16282 VDD.n6600 VDD.n2828 0.00359375
R16283 VDD.n5848 VDD.n5846 0.0033125
R16284 VDD.n5883 VDD.n5881 0.0033125
R16285 VDD.n5904 VDD.n5903 0.0033125
R16286 VDD.n5991 VDD.n5989 0.0033125
R16287 VDD.n6012 VDD.n6011 0.0033125
R16288 VDD.n6052 VDD.n6051 0.0033125
R16289 VDD.n4730 VDD.n4727 0.0033125
R16290 VDD.n4763 VDD.n4762 0.0033125
R16291 VDD.n4885 VDD.n4882 0.0033125
R16292 VDD.n4918 VDD.n4917 0.0033125
R16293 VDD.n6054 VDD.n6052 0.0033125
R16294 VDD.n6089 VDD.n6087 0.0033125
R16295 VDD.n6110 VDD.n6109 0.0033125
R16296 VDD.n6269 VDD.n6268 0.0033125
R16297 VDD.n6248 VDD.n6246 0.0033125
R16298 VDD.n6319 VDD.n5271 0.0033125
R16299 VDD.n5032 VDD.n5029 0.0033125
R16300 VDD.n5065 VDD.n5064 0.0033125
R16301 VDD.n5187 VDD.n5184 0.0033125
R16302 VDD.n5220 VDD.n5219 0.0033125
R16303 VDD.n6456 VDD.n5269 0.0033125
R16304 VDD.n6319 VDD.n6318 0.0033125
R16305 VDD.n2619 VDD.n2617 0.0033125
R16306 VDD.n2640 VDD.n2639 0.0033125
R16307 VDD.n6459 VDD.n6456 0.0033125
R16308 VDD.n6509 VDD.n6506 0.0033125
R16309 VDD.n6542 VDD.n6541 0.0033125
R16310 VDD.n8310 VDD.n8309 0.0033125
R16311 VDD.n337 VDD.n336 0.0033125
R16312 VDD.n370 VDD.n369 0.0033125
R16313 VDD.n8189 VDD.n8188 0.0033125
R16314 VDD.n8205 VDD.n8203 0.0033125
R16315 VDD.n4414 VDD.n4411 0.0033125
R16316 VDD.n4447 VDD.n4446 0.0033125
R16317 VDD.n4583 VDD.n4580 0.0033125
R16318 VDD.n4616 VDD.n4615 0.0033125
R16319 VDD.n5684 VDD.n5682 0.0033125
R16320 VDD.n5705 VDD.n5704 0.0033125
R16321 VDD.n5790 VDD.n5788 0.0033125
R16322 VDD.n5811 VDD.n5810 0.0033125
R16323 VDD.n5846 VDD.n5845 0.0033125
R16324 VDD.n4975 VDD.n3385 0.0032809
R16325 VDD.n4673 VDD.n3885 0.0032809
R16326 VDD.n5867 VDD.n5866 0.00275
R16327 VDD.n5920 VDD.n5918 0.00275
R16328 VDD.n5975 VDD.n5974 0.00275
R16329 VDD.n6028 VDD.n6026 0.00275
R16330 VDD.n4707 VDD.n4706 0.00275
R16331 VDD.n4786 VDD.n4783 0.00275
R16332 VDD.n4862 VDD.n4861 0.00275
R16333 VDD.n4941 VDD.n4938 0.00275
R16334 VDD.n6073 VDD.n6072 0.00275
R16335 VDD.n6126 VDD.n6124 0.00275
R16336 VDD.n6285 VDD.n6283 0.00275
R16337 VDD.n6232 VDD.n6231 0.00275
R16338 VDD.n5009 VDD.n5008 0.00275
R16339 VDD.n5088 VDD.n5085 0.00275
R16340 VDD.n5164 VDD.n5163 0.00275
R16341 VDD.n5243 VDD.n5240 0.00275
R16342 VDD.n2603 VDD.n2602 0.00275
R16343 VDD.n2656 VDD.n2654 0.00275
R16344 VDD.n6486 VDD.n6485 0.00275
R16345 VDD.n6565 VDD.n6562 0.00275
R16346 VDD.n4391 VDD.n4390 0.00275
R16347 VDD.n4470 VDD.n4467 0.00275
R16348 VDD.n4560 VDD.n4559 0.00275
R16349 VDD.n4639 VDD.n4636 0.00275
R16350 VDD.n5668 VDD.n5667 0.00275
R16351 VDD.n5721 VDD.n5719 0.00275
R16352 VDD.n5774 VDD.n5773 0.00275
R16353 VDD.n5827 VDD.n5825 0.00275
R16354 VDD.n1529 VDD.n1528 0.00246875
R16355 VDD.n1657 VDD.n1656 0.00246875
R16356 VDD.n2152 VDD.n2151 0.00246875
R16357 VDD.n2343 VDD.n2342 0.00246875
R16358 VDD.n7192 VDD.n7189 0.0021875
R16359 VDD.n7076 VDD.n7075 0.0021875
R16360 VDD.n4677 VDD.n4674 0.001625
R16361 VDD.n4832 VDD.n4829 0.001625
R16362 VDD.n1149 VDD.n1147 0.00134375
R16363 VDD.n1223 VDD.n1222 0.00134375
R16364 VDD.n2369 VDD.n2366 0.00134375
R16365 VDD.n2381 VDD.n2380 0.00134375
R16366 VDD.n2465 VDD.n2462 0.00134375
R16367 VDD.n2493 VDD.n2492 0.00134375
R16368 VDD.n5860 VDD.n5859 0.0010625
R16369 VDD.n5927 VDD.n5925 0.0010625
R16370 VDD.n5968 VDD.n5967 0.0010625
R16371 VDD.n6035 VDD.n6033 0.0010625
R16372 VDD.n4697 VDD.n4696 0.0010625
R16373 VDD.n4796 VDD.n4793 0.0010625
R16374 VDD.n4852 VDD.n4851 0.0010625
R16375 VDD.n4951 VDD.n4948 0.0010625
R16376 VDD.n6066 VDD.n6065 0.0010625
R16377 VDD.n6133 VDD.n6131 0.0010625
R16378 VDD.n6292 VDD.n6290 0.0010625
R16379 VDD.n6225 VDD.n6224 0.0010625
R16380 VDD.n4999 VDD.n4998 0.0010625
R16381 VDD.n5098 VDD.n5095 0.0010625
R16382 VDD.n5154 VDD.n5153 0.0010625
R16383 VDD.n5253 VDD.n5250 0.0010625
R16384 VDD.n2596 VDD.n2595 0.0010625
R16385 VDD.n2663 VDD.n2661 0.0010625
R16386 VDD.n6476 VDD.n6475 0.0010625
R16387 VDD.n6575 VDD.n6572 0.0010625
R16388 VDD.n8143 VDD.n7957 0.0010625
R16389 VDD.n4381 VDD.n4380 0.0010625
R16390 VDD.n4480 VDD.n4477 0.0010625
R16391 VDD.n4550 VDD.n4549 0.0010625
R16392 VDD.n4649 VDD.n4646 0.0010625
R16393 VDD.n5661 VDD.n5660 0.0010625
R16394 VDD.n5728 VDD.n5726 0.0010625
R16395 VDD.n5767 VDD.n5766 0.0010625
R16396 VDD.n5834 VDD.n5832 0.0010625
R16397 VDD.n2048 VDD.n2031 0.00078125
R16398 VDD.n2152 VDD.n1927 0.00078125
R16399 VDD.n2343 VDD.n1789 0.00078125
R16400 VDD.n1659 VDD.n1657 0.00078125
R16401 VDD.n2533 VDD.n1343 0.00078125
R16402 VDD.n1244 VDD.n1242 0.00078125
R16403 VDD.n2409 VDD.n2408 0.00078125
R16404 VDD.n2434 VDD.n2433 0.00078125
R16405 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n69 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t279 81.7344
R16406 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n70 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t514 81.7344
R16407 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n71 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t173 81.7344
R16408 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n72 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t408 81.7344
R16409 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n73 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t540 81.7344
R16410 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n74 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t211 81.7344
R16411 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n75 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t447 81.7344
R16412 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n86 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t431 81.7344
R16413 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n85 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t147 81.7344
R16414 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n84 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t374 81.7344
R16415 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n83 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t466 81.7344
R16416 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n82 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t274 81.7344
R16417 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n81 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t363 81.7344
R16418 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n80 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t457 81.7344
R16419 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n312 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t287 81.7344
R16420 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n313 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t247 81.7344
R16421 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n314 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t480 81.7344
R16422 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n315 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t145 81.7344
R16423 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n316 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t232 81.7344
R16424 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n317 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t464 81.7344
R16425 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n318 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t126 81.7344
R16426 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n329 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t161 81.7344
R16427 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n328 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t400 81.7344
R16428 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n327 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t487 81.7344
R16429 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n326 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t293 81.7344
R16430 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n325 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t432 81.7344
R16431 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n324 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t521 81.7344
R16432 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n323 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t327 81.7344
R16433 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n420 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t446 81.7344
R16434 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n421 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t529 81.7344
R16435 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n422 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t335 81.7344
R16436 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n423 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t428 81.7344
R16437 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n424 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t519 81.7344
R16438 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n425 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t372 81.7344
R16439 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n426 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t463 81.7344
R16440 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n437 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t454 81.7344
R16441 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n436 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t261 81.7344
R16442 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n435 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t398 81.7344
R16443 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n434 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t203 81.7344
R16444 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n433 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t291 81.7344
R16445 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n432 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t381 81.7344
R16446 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n431 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t191 81.7344
R16447 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n523 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t143 81.7344
R16448 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n524 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t370 81.7344
R16449 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n525 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t511 81.7344
R16450 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n526 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t316 81.7344
R16451 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n527 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t407 81.7344
R16452 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n528 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t496 81.7344
R16453 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n529 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t301 81.7344
R16454 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n540 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t337 81.7344
R16455 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n539 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t429 81.7344
R16456 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n538 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t238 81.7344
R16457 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n537 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t326 81.7344
R16458 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n536 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t137 81.7344
R16459 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n535 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t224 81.7344
R16460 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n534 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t362 81.7344
R16461 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n626 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t298 81.7344
R16462 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n627 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t392 81.7344
R16463 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n628 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t199 81.7344
R16464 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n629 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t333 81.7344
R16465 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n630 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t427 81.7344
R16466 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n631 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t234 81.7344
R16467 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n632 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t324 81.7344
R16468 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n643 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t356 81.7344
R16469 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n642 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t163 81.7344
R16470 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n641 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t258 81.7344
R16471 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n640 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t490 81.7344
R16472 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n639 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t154 81.7344
R16473 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n638 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t245 81.7344
R16474 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n637 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t478 81.7344
R16475 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n729 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t474 81.7344
R16476 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n730 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t283 81.7344
R16477 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n731 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t368 81.7344
R16478 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n732 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t178 81.7344
R16479 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n733 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t268 81.7344
R16480 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n734 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t355 81.7344
R16481 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n735 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t162 81.7344
R16482 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n746 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t200 81.7344
R16483 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n745 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t290 81.7344
R16484 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n744 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t524 81.7344
R16485 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n743 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t188 81.7344
R16486 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n742 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t471 81.7344
R16487 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n741 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t132 81.7344
R16488 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n740 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t223 81.7344
R16489 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n214 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t313 81.7344
R16490 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n215 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t539 81.7344
R16491 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n216 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t209 81.7344
R16492 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n217 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t445 81.7344
R16493 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n218 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t531 81.7344
R16494 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n219 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t198 81.7344
R16495 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n220 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t477 81.7344
R16496 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n231 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t462 81.7344
R16497 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n230 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t122 81.7344
R16498 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n229 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t358 81.7344
R16499 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n228 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t497 81.7344
R16500 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n227 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t304 81.7344
R16501 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n226 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t397 81.7344
R16502 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n225 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t485 81.7344
R16503 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n10 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t59 53.5894
R16504 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n7 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t9 53.5894
R16505 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n253 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t19 53.5894
R16506 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n250 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t37 53.5894
R16507 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n361 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t51 53.5894
R16508 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n358 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t75 53.5894
R16509 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n464 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t93 53.5894
R16510 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n461 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t43 53.5894
R16511 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n567 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t83 53.5894
R16512 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n564 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t113 53.5894
R16513 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n670 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t5 53.5894
R16514 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n667 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t69 53.5894
R16515 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n114 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t49 53.5894
R16516 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n109 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t111 53.5894
R16517 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n19 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t7 47.0594
R16518 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n32 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t115 47.0594
R16519 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n59 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t95 47.0594
R16520 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n87 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t71 47.0594
R16521 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n48 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t101 47.0594
R16522 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n76 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t25 47.0594
R16523 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n69 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t228 47.0594
R16524 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n70 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t460 47.0594
R16525 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n71 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t541 47.0594
R16526 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n72 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t354 47.0594
R16527 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n73 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t495 47.0594
R16528 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n74 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t158 47.0594
R16529 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n75 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t391 47.0594
R16530 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n86 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t377 47.0594
R16531 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n85 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t518 47.0594
R16532 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n84 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t323 47.0594
R16533 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n83 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t413 47.0594
R16534 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n82 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t221 47.0594
R16535 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n26 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t508 47.0594
R16536 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n12 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t144 47.0594
R16537 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n41 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t197 47.0594
R16538 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n13 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t157 47.0594
R16539 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n42 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t210 47.0594
R16540 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n14 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t280 47.0594
R16541 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n43 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t330 47.0594
R16542 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n15 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t294 47.0594
R16543 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n44 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t348 47.0594
R16544 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n16 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t275 47.0594
R16545 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n45 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t325 47.0594
R16546 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n17 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t401 47.0594
R16547 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n46 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t455 47.0594
R16548 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n18 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t414 47.0594
R16549 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n47 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t467 47.0594
R16550 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n31 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t252 47.0594
R16551 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n58 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t300 47.0594
R16552 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n30 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t230 47.0594
R16553 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n57 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t281 47.0594
R16554 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n29 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t249 47.0594
R16555 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n56 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t295 47.0594
R16556 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n28 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t367 47.0594
R16557 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n55 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t420 47.0594
R16558 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n27 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t384 47.0594
R16559 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n54 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t438 47.0594
R16560 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n25 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t206 47.0594
R16561 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n52 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t262 47.0594
R16562 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n53 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t136 47.0594
R16563 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n81 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t314 47.0594
R16564 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n80 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t404 47.0594
R16565 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n274 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t63 47.0594
R16566 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n302 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t45 47.0594
R16567 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n330 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t31 47.0594
R16568 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n263 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t91 47.0594
R16569 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n291 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t77 47.0594
R16570 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n319 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t53 47.0594
R16571 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n312 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t235 47.0594
R16572 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n313 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t194 47.0594
R16573 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n314 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t426 47.0594
R16574 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n315 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t517 47.0594
R16575 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n316 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t176 47.0594
R16576 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n317 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t411 47.0594
R16577 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n318 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t501 47.0594
R16578 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n329 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t533 47.0594
R16579 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n328 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t346 47.0594
R16580 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n327 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t434 47.0594
R16581 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n326 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t242 47.0594
R16582 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n325 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t378 47.0594
R16583 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n268 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t289 47.0594
R16584 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n256 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t334 47.0594
R16585 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n284 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t389 47.0594
R16586 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n257 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t365 47.0594
R16587 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n285 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t416 47.0594
R16588 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n258 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t380 47.0594
R16589 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n286 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t436 47.0594
R16590 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n259 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t505 47.0594
R16591 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n287 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t131 47.0594
R16592 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n260 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t201 47.0594
R16593 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n288 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t257 47.0594
R16594 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n261 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t215 47.0594
R16595 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n289 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t269 47.0594
R16596 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n262 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t339 47.0594
R16597 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n290 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t394 47.0594
R16598 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n273 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t459 47.0594
R16599 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n301 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t512 47.0594
R16600 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n272 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t475 47.0594
R16601 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n300 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t527 47.0594
R16602 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n271 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t171 47.0594
R16603 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n299 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t226 47.0594
R16604 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n270 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t190 47.0594
R16605 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n298 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t244 47.0594
R16606 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n269 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t165 47.0594
R16607 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n297 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t217 47.0594
R16608 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n267 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t308 47.0594
R16609 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n295 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t357 47.0594
R16610 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n296 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t343 47.0594
R16611 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n324 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t469 47.0594
R16612 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n323 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t277 47.0594
R16613 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n382 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t85 47.0594
R16614 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n410 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t73 47.0594
R16615 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n438 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t67 47.0594
R16616 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n371 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t13 47.0594
R16617 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n399 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t109 47.0594
R16618 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n427 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t87 47.0594
R16619 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n420 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t388 47.0594
R16620 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n421 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t482 47.0594
R16621 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n422 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t285 47.0594
R16622 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n423 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t375 47.0594
R16623 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n424 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t465 47.0594
R16624 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n425 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t320 47.0594
R16625 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n426 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t409 47.0594
R16626 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n437 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t402 47.0594
R16627 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n436 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t207 47.0594
R16628 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n435 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t344 47.0594
R16629 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n434 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t152 47.0594
R16630 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n433 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t240 47.0594
R16631 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n376 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t174 47.0594
R16632 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n364 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t123 47.0594
R16633 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n392 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t177 47.0594
R16634 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n365 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t250 47.0594
R16635 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n393 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t297 47.0594
R16636 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n366 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t265 47.0594
R16637 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n394 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t315 47.0594
R16638 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n367 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t386 47.0594
R16639 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n395 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t443 47.0594
R16640 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n368 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t513 47.0594
R16641 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n396 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t142 47.0594
R16642 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n369 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t383 47.0594
R16643 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n397 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t439 47.0594
R16644 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n370 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t507 47.0594
R16645 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n398 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t134 47.0594
R16646 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n381 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t345 47.0594
R16647 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n409 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t399 47.0594
R16648 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n380 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t361 47.0594
R16649 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n408 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t412 47.0594
R16650 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n379 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t336 47.0594
R16651 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n407 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t390 47.0594
R16652 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n378 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t352 47.0594
R16653 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n406 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t406 47.0594
R16654 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n377 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t483 47.0594
R16655 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n405 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t530 47.0594
R16656 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n375 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t195 47.0594
R16657 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n403 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t248 47.0594
R16658 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n404 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t229 47.0594
R16659 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n432 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t328 47.0594
R16660 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n431 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t140 47.0594
R16661 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n485 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t33 47.0594
R16662 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n513 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t21 47.0594
R16663 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n541 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t107 47.0594
R16664 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n474 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t35 47.0594
R16665 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n502 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t27 47.0594
R16666 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n530 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t57 47.0594
R16667 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n523 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t515 47.0594
R16668 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n524 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t318 47.0594
R16669 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n525 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t458 47.0594
R16670 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n526 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t266 47.0594
R16671 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n527 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t353 47.0594
R16672 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n528 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t448 47.0594
R16673 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n529 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t253 47.0594
R16674 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n540 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t286 47.0594
R16675 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n539 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t376 47.0594
R16676 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n538 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t185 47.0594
R16677 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n537 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t276 47.0594
R16678 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n536 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t509 47.0594
R16679 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n479 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t395 47.0594
R16680 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n467 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t456 47.0594
R16681 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n495 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t503 47.0594
R16682 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n468 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t468 47.0594
R16683 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n496 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t520 47.0594
R16684 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n469 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t451 47.0594
R16685 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n497 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t498 47.0594
R16686 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n470 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t461 47.0594
R16687 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n498 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t516 47.0594
R16688 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n471 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t160 47.0594
R16689 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n499 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t212 47.0594
R16690 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n472 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t282 47.0594
R16691 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n500 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t331 47.0594
R16692 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n473 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t296 47.0594
R16693 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n501 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t349 47.0594
R16694 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n484 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t417 47.0594
R16695 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n512 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t470 47.0594
R16696 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n483 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t538 47.0594
R16697 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n511 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t164 47.0594
R16698 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n482 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t128 47.0594
R16699 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n510 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t182 47.0594
R16700 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n481 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t254 47.0594
R16701 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n509 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t306 47.0594
R16702 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n480 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t270 47.0594
R16703 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n508 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t322 47.0594
R16704 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n478 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t369 47.0594
R16705 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n506 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t424 47.0594
R16706 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n507 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t450 47.0594
R16707 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n535 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t170 47.0594
R16708 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n534 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t311 47.0594
R16709 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n588 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t11 47.0594
R16710 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n616 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t105 47.0594
R16711 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n644 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t99 47.0594
R16712 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n577 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t39 47.0594
R16713 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n605 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t29 47.0594
R16714 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n633 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t17 47.0594
R16715 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n626 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t251 47.0594
R16716 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n627 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t338 47.0594
R16717 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n628 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t149 47.0594
R16718 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n629 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t284 47.0594
R16719 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n630 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t373 47.0594
R16720 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n631 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t180 47.0594
R16721 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n632 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t272 47.0594
R16722 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n643 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t305 47.0594
R16723 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n642 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t537 47.0594
R16724 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n641 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t204 47.0594
R16725 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n640 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t441 47.0594
R16726 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n639 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t525 47.0594
R16727 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n582 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t488 47.0594
R16728 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n570 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t440 47.0594
R16729 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n598 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t492 47.0594
R16730 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n571 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t135 47.0594
R16731 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n599 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t187 47.0594
R16732 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n572 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t153 47.0594
R16733 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n600 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t205 47.0594
R16734 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n573 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t129 47.0594
R16735 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n601 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t181 47.0594
R16736 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n574 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t255 47.0594
R16737 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n602 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t302 47.0594
R16738 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n575 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t267 47.0594
R16739 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n603 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t321 47.0594
R16740 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n576 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t393 47.0594
R16741 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n604 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t449 47.0594
R16742 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n587 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t510 47.0594
R16743 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n615 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t139 47.0594
R16744 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n586 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t526 47.0594
R16745 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n614 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t155 47.0594
R16746 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n585 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t225 47.0594
R16747 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n613 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t278 47.0594
R16748 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n584 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t241 47.0594
R16749 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n612 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t292 47.0594
R16750 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n583 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t364 47.0594
R16751 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n611 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t415 47.0594
R16752 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n581 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t502 47.0594
R16753 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n609 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t127 47.0594
R16754 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n610 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t535 47.0594
R16755 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n638 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t192 47.0594
R16756 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n637 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t423 47.0594
R16757 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n691 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t97 47.0594
R16758 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n719 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t81 47.0594
R16759 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n747 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t23 47.0594
R16760 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n680 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t103 47.0594
R16761 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n708 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t89 47.0594
R16762 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n736 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t79 47.0594
R16763 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n729 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t421 47.0594
R16764 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n730 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t231 47.0594
R16765 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n731 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t317 47.0594
R16766 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n732 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t124 47.0594
R16767 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n733 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t214 47.0594
R16768 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n734 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t303 47.0594
R16769 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n735 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t536 47.0594
R16770 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n746 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t150 47.0594
R16771 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n745 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t239 47.0594
R16772 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n744 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t473 47.0594
R16773 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n743 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t138 47.0594
R16774 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n742 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t418 47.0594
R16775 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n685 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t133 47.0594
R16776 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n673 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t196 47.0594
R16777 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n701 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t246 47.0594
R16778 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n674 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t208 47.0594
R16779 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n702 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t263 47.0594
R16780 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n675 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t329 47.0594
R16781 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n703 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t382 47.0594
R16782 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n676 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t347 47.0594
R16783 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n704 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t403 47.0594
R16784 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n677 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t472 47.0594
R16785 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n705 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t523 47.0594
R16786 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n678 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t166 47.0594
R16787 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n706 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t218 47.0594
R16788 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n679 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t183 47.0594
R16789 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n707 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t237 47.0594
R16790 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n690 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t299 47.0594
R16791 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n718 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t351 47.0594
R16792 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n689 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t425 47.0594
R16793 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n717 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t479 47.0594
R16794 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n688 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t444 47.0594
R16795 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n716 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t494 47.0594
R16796 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n687 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t141 47.0594
R16797 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n715 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t193 47.0594
R16798 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n686 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t437 47.0594
R16799 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n714 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t489 47.0594
R16800 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n684 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t259 47.0594
R16801 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n712 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t312 47.0594
R16802 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n713 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t186 47.0594
R16803 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n741 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t506 47.0594
R16804 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n740 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t169 47.0594
R16805 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n125 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t61 47.0594
R16806 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n136 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t55 47.0594
R16807 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n194 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t47 47.0594
R16808 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n205 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t41 47.0594
R16809 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n232 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t65 47.0594
R16810 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n221 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t15 47.0594
R16811 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n214 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t260 47.0594
R16812 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n215 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t493 47.0594
R16813 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n216 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t156 47.0594
R16814 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n217 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t387 47.0594
R16815 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n218 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t481 47.0594
R16816 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n219 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t146 47.0594
R16817 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n220 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t422 47.0594
R16818 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n231 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t410 47.0594
R16819 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n230 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t500 47.0594
R16820 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n229 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t309 47.0594
R16821 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n228 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t452 47.0594
R16822 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n227 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t256 47.0594
R16823 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n130 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t307 47.0594
R16824 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n118 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t366 47.0594
R16825 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n187 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t419 47.0594
R16826 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n119 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t379 47.0594
R16827 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n188 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t435 47.0594
R16828 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n120 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t504 47.0594
R16829 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n189 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t130 47.0594
R16830 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n121 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t522 47.0594
R16831 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n190 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t148 47.0594
R16832 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n122 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t216 47.0594
R16833 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n191 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t271 47.0594
R16834 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n123 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t340 47.0594
R16835 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n192 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t396 47.0594
R16836 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n124 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t213 47.0594
R16837 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n193 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t264 47.0594
R16838 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n135 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t476 47.0594
R16839 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n204 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t528 47.0594
R16840 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n134 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t172 47.0594
R16841 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n203 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t227 47.0594
R16842 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n133 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t189 47.0594
R16843 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n202 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t243 47.0594
R16844 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n132 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t167 47.0594
R16845 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n201 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t219 47.0594
R16846 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n131 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t184 47.0594
R16847 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n200 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t236 47.0594
R16848 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n129 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t430 47.0594
R16849 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n198 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t484 47.0594
R16850 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n199 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t359 47.0594
R16851 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n226 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t342 47.0594
R16852 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n225 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t433 47.0594
R16853 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n13 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n12 16.2227
R16854 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n14 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n13 16.2227
R16855 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n15 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n14 16.2227
R16856 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n16 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n15 16.2227
R16857 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n17 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n16 16.2227
R16858 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n18 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n17 16.2227
R16859 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n19 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n18 16.2227
R16860 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n32 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n31 16.2227
R16861 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n31 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n30 16.2227
R16862 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n30 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n29 16.2227
R16863 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n29 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n28 16.2227
R16864 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n28 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n27 16.2227
R16865 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n27 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n26 16.2227
R16866 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n26 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n25 16.2227
R16867 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n42 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n41 16.2227
R16868 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n43 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n42 16.2227
R16869 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n44 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n43 16.2227
R16870 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n45 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n44 16.2227
R16871 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n46 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n45 16.2227
R16872 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n47 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n46 16.2227
R16873 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n48 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n47 16.2227
R16874 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n59 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n58 16.2227
R16875 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n58 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n57 16.2227
R16876 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n57 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n56 16.2227
R16877 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n56 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n55 16.2227
R16878 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n55 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n54 16.2227
R16879 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n54 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n53 16.2227
R16880 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n53 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n52 16.2227
R16881 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n70 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n69 16.2227
R16882 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n71 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n70 16.2227
R16883 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n72 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n71 16.2227
R16884 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n73 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n72 16.2227
R16885 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n74 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n73 16.2227
R16886 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n75 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n74 16.2227
R16887 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n76 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n75 16.2227
R16888 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n87 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n86 16.2227
R16889 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n86 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n85 16.2227
R16890 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n85 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n84 16.2227
R16891 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n84 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n83 16.2227
R16892 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n83 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n82 16.2227
R16893 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n82 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n81 16.2227
R16894 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n81 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n80 16.2227
R16895 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n257 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n256 16.2227
R16896 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n258 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n257 16.2227
R16897 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n259 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n258 16.2227
R16898 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n260 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n259 16.2227
R16899 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n261 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n260 16.2227
R16900 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n262 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n261 16.2227
R16901 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n263 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n262 16.2227
R16902 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n274 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n273 16.2227
R16903 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n273 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n272 16.2227
R16904 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n272 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n271 16.2227
R16905 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n271 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n270 16.2227
R16906 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n270 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n269 16.2227
R16907 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n269 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n268 16.2227
R16908 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n268 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n267 16.2227
R16909 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n285 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n284 16.2227
R16910 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n286 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n285 16.2227
R16911 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n287 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n286 16.2227
R16912 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n288 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n287 16.2227
R16913 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n289 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n288 16.2227
R16914 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n290 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n289 16.2227
R16915 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n291 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n290 16.2227
R16916 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n302 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n301 16.2227
R16917 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n301 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n300 16.2227
R16918 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n300 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n299 16.2227
R16919 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n299 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n298 16.2227
R16920 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n298 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n297 16.2227
R16921 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n297 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n296 16.2227
R16922 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n296 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n295 16.2227
R16923 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n313 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n312 16.2227
R16924 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n314 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n313 16.2227
R16925 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n315 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n314 16.2227
R16926 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n316 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n315 16.2227
R16927 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n317 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n316 16.2227
R16928 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n318 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n317 16.2227
R16929 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n319 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n318 16.2227
R16930 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n330 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n329 16.2227
R16931 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n329 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n328 16.2227
R16932 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n328 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n327 16.2227
R16933 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n327 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n326 16.2227
R16934 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n326 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n325 16.2227
R16935 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n325 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n324 16.2227
R16936 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n324 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n323 16.2227
R16937 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n365 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n364 16.2227
R16938 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n366 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n365 16.2227
R16939 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n367 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n366 16.2227
R16940 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n368 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n367 16.2227
R16941 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n369 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n368 16.2227
R16942 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n370 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n369 16.2227
R16943 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n371 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n370 16.2227
R16944 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n382 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n381 16.2227
R16945 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n381 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n380 16.2227
R16946 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n380 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n379 16.2227
R16947 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n379 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n378 16.2227
R16948 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n378 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n377 16.2227
R16949 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n377 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n376 16.2227
R16950 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n376 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n375 16.2227
R16951 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n393 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n392 16.2227
R16952 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n394 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n393 16.2227
R16953 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n395 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n394 16.2227
R16954 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n396 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n395 16.2227
R16955 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n397 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n396 16.2227
R16956 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n398 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n397 16.2227
R16957 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n399 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n398 16.2227
R16958 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n410 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n409 16.2227
R16959 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n409 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n408 16.2227
R16960 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n408 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n407 16.2227
R16961 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n407 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n406 16.2227
R16962 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n406 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n405 16.2227
R16963 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n405 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n404 16.2227
R16964 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n404 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n403 16.2227
R16965 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n421 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n420 16.2227
R16966 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n422 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n421 16.2227
R16967 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n423 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n422 16.2227
R16968 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n424 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n423 16.2227
R16969 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n425 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n424 16.2227
R16970 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n426 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n425 16.2227
R16971 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n427 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n426 16.2227
R16972 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n438 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n437 16.2227
R16973 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n437 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n436 16.2227
R16974 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n436 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n435 16.2227
R16975 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n435 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n434 16.2227
R16976 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n434 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n433 16.2227
R16977 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n433 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n432 16.2227
R16978 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n432 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n431 16.2227
R16979 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n468 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n467 16.2227
R16980 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n469 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n468 16.2227
R16981 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n470 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n469 16.2227
R16982 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n471 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n470 16.2227
R16983 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n472 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n471 16.2227
R16984 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n473 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n472 16.2227
R16985 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n474 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n473 16.2227
R16986 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n485 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n484 16.2227
R16987 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n484 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n483 16.2227
R16988 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n483 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n482 16.2227
R16989 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n482 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n481 16.2227
R16990 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n481 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n480 16.2227
R16991 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n480 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n479 16.2227
R16992 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n479 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n478 16.2227
R16993 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n496 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n495 16.2227
R16994 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n497 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n496 16.2227
R16995 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n498 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n497 16.2227
R16996 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n499 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n498 16.2227
R16997 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n500 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n499 16.2227
R16998 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n501 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n500 16.2227
R16999 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n502 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n501 16.2227
R17000 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n513 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n512 16.2227
R17001 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n512 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n511 16.2227
R17002 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n511 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n510 16.2227
R17003 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n510 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n509 16.2227
R17004 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n509 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n508 16.2227
R17005 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n508 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n507 16.2227
R17006 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n507 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n506 16.2227
R17007 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n524 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n523 16.2227
R17008 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n525 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n524 16.2227
R17009 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n526 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n525 16.2227
R17010 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n527 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n526 16.2227
R17011 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n528 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n527 16.2227
R17012 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n529 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n528 16.2227
R17013 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n530 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n529 16.2227
R17014 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n541 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n540 16.2227
R17015 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n540 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n539 16.2227
R17016 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n539 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n538 16.2227
R17017 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n538 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n537 16.2227
R17018 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n537 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n536 16.2227
R17019 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n536 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n535 16.2227
R17020 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n535 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n534 16.2227
R17021 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n571 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n570 16.2227
R17022 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n572 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n571 16.2227
R17023 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n573 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n572 16.2227
R17024 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n574 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n573 16.2227
R17025 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n575 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n574 16.2227
R17026 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n576 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n575 16.2227
R17027 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n577 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n576 16.2227
R17028 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n588 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n587 16.2227
R17029 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n587 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n586 16.2227
R17030 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n586 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n585 16.2227
R17031 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n585 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n584 16.2227
R17032 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n584 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n583 16.2227
R17033 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n583 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n582 16.2227
R17034 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n582 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n581 16.2227
R17035 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n599 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n598 16.2227
R17036 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n600 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n599 16.2227
R17037 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n601 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n600 16.2227
R17038 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n602 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n601 16.2227
R17039 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n603 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n602 16.2227
R17040 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n604 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n603 16.2227
R17041 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n605 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n604 16.2227
R17042 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n616 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n615 16.2227
R17043 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n615 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n614 16.2227
R17044 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n614 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n613 16.2227
R17045 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n613 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n612 16.2227
R17046 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n612 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n611 16.2227
R17047 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n611 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n610 16.2227
R17048 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n610 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n609 16.2227
R17049 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n627 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n626 16.2227
R17050 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n628 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n627 16.2227
R17051 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n629 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n628 16.2227
R17052 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n630 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n629 16.2227
R17053 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n631 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n630 16.2227
R17054 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n632 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n631 16.2227
R17055 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n633 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n632 16.2227
R17056 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n644 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n643 16.2227
R17057 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n643 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n642 16.2227
R17058 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n642 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n641 16.2227
R17059 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n641 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n640 16.2227
R17060 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n640 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n639 16.2227
R17061 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n639 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n638 16.2227
R17062 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n638 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n637 16.2227
R17063 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n674 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n673 16.2227
R17064 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n675 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n674 16.2227
R17065 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n676 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n675 16.2227
R17066 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n677 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n676 16.2227
R17067 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n678 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n677 16.2227
R17068 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n679 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n678 16.2227
R17069 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n680 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n679 16.2227
R17070 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n691 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n690 16.2227
R17071 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n690 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n689 16.2227
R17072 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n689 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n688 16.2227
R17073 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n688 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n687 16.2227
R17074 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n687 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n686 16.2227
R17075 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n686 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n685 16.2227
R17076 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n685 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n684 16.2227
R17077 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n702 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n701 16.2227
R17078 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n703 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n702 16.2227
R17079 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n704 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n703 16.2227
R17080 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n705 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n704 16.2227
R17081 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n706 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n705 16.2227
R17082 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n707 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n706 16.2227
R17083 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n708 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n707 16.2227
R17084 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n719 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n718 16.2227
R17085 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n718 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n717 16.2227
R17086 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n717 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n716 16.2227
R17087 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n716 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n715 16.2227
R17088 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n715 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n714 16.2227
R17089 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n714 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n713 16.2227
R17090 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n713 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n712 16.2227
R17091 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n730 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n729 16.2227
R17092 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n731 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n730 16.2227
R17093 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n732 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n731 16.2227
R17094 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n733 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n732 16.2227
R17095 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n734 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n733 16.2227
R17096 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n735 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n734 16.2227
R17097 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n736 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n735 16.2227
R17098 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n747 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n746 16.2227
R17099 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n746 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n745 16.2227
R17100 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n745 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n744 16.2227
R17101 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n744 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n743 16.2227
R17102 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n743 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n742 16.2227
R17103 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n742 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n741 16.2227
R17104 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n741 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n740 16.2227
R17105 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n119 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n118 16.2227
R17106 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n120 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n119 16.2227
R17107 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n121 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n120 16.2227
R17108 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n122 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n121 16.2227
R17109 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n123 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n122 16.2227
R17110 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n124 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n123 16.2227
R17111 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n125 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n124 16.2227
R17112 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n136 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n135 16.2227
R17113 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n135 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n134 16.2227
R17114 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n134 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n133 16.2227
R17115 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n133 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n132 16.2227
R17116 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n132 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n131 16.2227
R17117 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n131 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n130 16.2227
R17118 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n130 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n129 16.2227
R17119 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n188 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n187 16.2227
R17120 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n189 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n188 16.2227
R17121 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n190 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n189 16.2227
R17122 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n191 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n190 16.2227
R17123 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n192 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n191 16.2227
R17124 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n193 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n192 16.2227
R17125 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n194 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n193 16.2227
R17126 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n205 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n204 16.2227
R17127 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n204 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n203 16.2227
R17128 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n203 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n202 16.2227
R17129 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n202 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n201 16.2227
R17130 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n201 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n200 16.2227
R17131 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n200 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n199 16.2227
R17132 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n199 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n198 16.2227
R17133 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n215 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n214 16.2227
R17134 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n216 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n215 16.2227
R17135 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n217 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n216 16.2227
R17136 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n218 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n217 16.2227
R17137 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n219 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n218 16.2227
R17138 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n220 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n219 16.2227
R17139 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n221 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n220 16.2227
R17140 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n232 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n231 16.2227
R17141 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n231 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n230 16.2227
R17142 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n230 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n229 16.2227
R17143 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n229 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n228 16.2227
R17144 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n228 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n227 16.2227
R17145 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n227 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n226 16.2227
R17146 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n226 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n225 16.2227
R17147 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n180 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n179 11.6793
R17148 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n142 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t119 4.65943
R17149 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n154 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n153 3.86296
R17150 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n169 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n168 3.86296
R17151 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n90 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n79 3.30289
R17152 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n62 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n51 3.30289
R17153 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n6 3.30289
R17154 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n333 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n322 3.30289
R17155 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n305 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n294 3.30289
R17156 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n277 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n266 3.30289
R17157 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n252 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n249 3.30289
R17158 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n441 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n430 3.30289
R17159 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n413 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n402 3.30289
R17160 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n385 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n374 3.30289
R17161 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n360 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n357 3.30289
R17162 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n544 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n533 3.30289
R17163 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n516 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n505 3.30289
R17164 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n488 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n477 3.30289
R17165 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n463 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n460 3.30289
R17166 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n647 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n636 3.30289
R17167 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n619 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n608 3.30289
R17168 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n591 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n580 3.30289
R17169 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n566 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n563 3.30289
R17170 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n750 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n739 3.30289
R17171 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n722 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n711 3.30289
R17172 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n694 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n683 3.30289
R17173 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n669 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n666 3.30289
R17174 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n224 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n213 3.30289
R17175 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n197 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n186 3.30289
R17176 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n128 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n117 3.30289
R17177 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n113 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n112 3.30289
R17178 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n24 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n23 3.30289
R17179 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n33 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n32 2.8805
R17180 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n49 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n48 2.8805
R17181 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n77 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n76 2.8805
R17182 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n264 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n263 2.8805
R17183 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n292 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n291 2.8805
R17184 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n320 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n319 2.8805
R17185 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n303 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n302 2.8805
R17186 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n331 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n330 2.8805
R17187 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n275 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n274 2.8805
R17188 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n372 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n371 2.8805
R17189 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n400 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n399 2.8805
R17190 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n428 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n427 2.8805
R17191 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n411 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n410 2.8805
R17192 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n439 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n438 2.8805
R17193 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n383 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n382 2.8805
R17194 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n475 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n474 2.8805
R17195 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n503 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n502 2.8805
R17196 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n531 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n530 2.8805
R17197 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n514 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n513 2.8805
R17198 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n542 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n541 2.8805
R17199 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n486 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n485 2.8805
R17200 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n578 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n577 2.8805
R17201 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n606 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n605 2.8805
R17202 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n634 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n633 2.8805
R17203 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n617 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n616 2.8805
R17204 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n645 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n644 2.8805
R17205 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n589 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n588 2.8805
R17206 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n681 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n680 2.8805
R17207 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n709 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n708 2.8805
R17208 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n737 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n736 2.8805
R17209 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n720 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n719 2.8805
R17210 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n748 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n747 2.8805
R17211 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n692 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n691 2.8805
R17212 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n137 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n136 2.8805
R17213 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n206 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n205 2.8805
R17214 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n233 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n232 2.8805
R17215 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n222 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n221 2.8805
R17216 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n195 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n194 2.8805
R17217 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n126 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n125 2.8805
R17218 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n60 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n59 2.8805
R17219 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n88 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n87 2.8805
R17220 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n20 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n19 2.8805
R17221 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n661 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n660 1.69656
R17222 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n455 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n454 1.69656
R17223 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n347 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n346 1.69656
R17224 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n159 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n158 1.44217
R17225 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n174 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n173 1.44217
R17226 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n558 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n557 1.24529
R17227 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n352 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n351 1.24529
R17228 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n244 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n243 1.24529
R17229 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n141 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n140 1.16617
R17230 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n160 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n159 1.14036
R17231 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n175 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n174 1.14036
R17232 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n144 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n143 1.1255
R17233 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n156 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n155 1.1255
R17234 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n171 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n170 1.1255
R17235 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n335 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n334 1.1228
R17236 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n307 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n306 1.1228
R17237 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n279 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n278 1.1228
R17238 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n443 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n442 1.1228
R17239 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n415 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n414 1.1228
R17240 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n387 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n386 1.1228
R17241 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n546 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n545 1.1228
R17242 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n518 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n517 1.1228
R17243 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n490 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n489 1.1228
R17244 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n649 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n648 1.1228
R17245 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n621 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n620 1.1228
R17246 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n593 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n592 1.1228
R17247 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n752 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n751 1.1228
R17248 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n724 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n723 1.1228
R17249 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n696 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n695 1.1228
R17250 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n92 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n91 1.1228
R17251 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n64 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n63 1.1228
R17252 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n36 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n34 1.12272
R17253 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n96 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n11 1.12272
R17254 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n339 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n254 1.12272
R17255 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n447 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n362 1.12272
R17256 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n550 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n465 1.12272
R17257 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n653 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n568 1.12272
R17258 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n756 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n671 1.12272
R17259 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n235 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n234 1.12272
R17260 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n208 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n207 1.12272
R17261 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n181 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n138 1.12272
R17262 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n239 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n115 1.12272
R17263 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n239 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n110 1.12243
R17264 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n346 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n345 1.11801
R17265 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n763 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n762 1.11801
R17266 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n660 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n659 1.11801
R17267 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n557 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n556 1.11801
R17268 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n454 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n453 1.11801
R17269 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n242 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n241 1.11782
R17270 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n760 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n759 1.11782
R17271 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n657 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n656 1.11782
R17272 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n554 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n553 1.11782
R17273 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n451 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n450 1.11782
R17274 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n343 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n342 1.11782
R17275 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n351 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n102 1.11782
R17276 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n140 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n139 1.07327
R17277 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n764 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n763 0.962646
R17278 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n139 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t120 0.8195
R17279 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n158 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t4 0.8195
R17280 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n158 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n157 0.8195
R17281 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n153 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t3 0.8195
R17282 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n153 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n152 0.8195
R17283 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n173 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t1 0.8195
R17284 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n173 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n172 0.8195
R17285 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n168 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t117 0.8195
R17286 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n168 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n167 0.8195
R17287 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n768 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n767 0.767554
R17288 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n4 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n3 0.7505
R17289 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n162 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n161 0.727916
R17290 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n177 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n176 0.727916
R17291 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n147 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n145 0.616779
R17292 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n79 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t26 0.607167
R17293 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n79 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n78 0.607167
R17294 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n51 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t102 0.607167
R17295 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n51 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n50 0.607167
R17296 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n6 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t10 0.607167
R17297 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n6 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n5 0.607167
R17298 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n322 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t54 0.607167
R17299 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n322 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n321 0.607167
R17300 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n294 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t78 0.607167
R17301 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n294 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n293 0.607167
R17302 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n266 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t92 0.607167
R17303 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n266 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n265 0.607167
R17304 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n249 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t38 0.607167
R17305 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n249 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n248 0.607167
R17306 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n430 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t88 0.607167
R17307 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n430 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n429 0.607167
R17308 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n402 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t110 0.607167
R17309 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n402 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n401 0.607167
R17310 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n374 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t14 0.607167
R17311 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n374 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n373 0.607167
R17312 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n357 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t76 0.607167
R17313 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n357 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n356 0.607167
R17314 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n533 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t58 0.607167
R17315 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n533 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n532 0.607167
R17316 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n505 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t28 0.607167
R17317 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n505 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n504 0.607167
R17318 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n477 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t36 0.607167
R17319 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n477 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n476 0.607167
R17320 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n460 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t44 0.607167
R17321 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n460 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n459 0.607167
R17322 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n636 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t18 0.607167
R17323 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n636 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n635 0.607167
R17324 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n608 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t30 0.607167
R17325 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n608 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n607 0.607167
R17326 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n580 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t40 0.607167
R17327 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n580 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n579 0.607167
R17328 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n563 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t114 0.607167
R17329 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n563 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n562 0.607167
R17330 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n739 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t80 0.607167
R17331 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n739 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n738 0.607167
R17332 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n711 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t90 0.607167
R17333 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n711 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n710 0.607167
R17334 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n683 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t104 0.607167
R17335 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n683 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n682 0.607167
R17336 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n666 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t70 0.607167
R17337 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n666 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n665 0.607167
R17338 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n213 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t16 0.607167
R17339 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n213 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n212 0.607167
R17340 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n186 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t48 0.607167
R17341 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n186 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n185 0.607167
R17342 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n117 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t62 0.607167
R17343 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n117 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n116 0.607167
R17344 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n112 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t112 0.607167
R17345 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n112 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n111 0.607167
R17346 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n23 Folded_Diff_Op_Amp_Layout_0.IBIAS2.t8 0.607167
R17347 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n23 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n22 0.607167
R17348 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n338 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n337 0.386051
R17349 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n310 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n309 0.386051
R17350 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n282 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n281 0.386051
R17351 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n446 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n445 0.386051
R17352 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n418 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n417 0.386051
R17353 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n390 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n389 0.386051
R17354 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n549 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n548 0.386051
R17355 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n521 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n520 0.386051
R17356 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n493 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n492 0.386051
R17357 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n652 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n651 0.386051
R17358 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n624 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n623 0.386051
R17359 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n596 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n595 0.386051
R17360 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n755 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n754 0.386051
R17361 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n727 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n726 0.386051
R17362 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n699 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n698 0.386051
R17363 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n238 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n237 0.386051
R17364 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n211 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n210 0.386051
R17365 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n184 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n183 0.386051
R17366 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n95 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n94 0.386051
R17367 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n67 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n66 0.386051
R17368 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n39 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n38 0.386051
R17369 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n342 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n341 0.380932
R17370 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n450 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n449 0.380932
R17371 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n553 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n552 0.380932
R17372 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n656 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n655 0.380932
R17373 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n759 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n758 0.380932
R17374 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n241 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n240 0.380932
R17375 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n99 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n98 0.380932
R17376 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n165 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n164 0.2775
R17377 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n150 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n149 0.2775
R17378 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n767 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n766 0.147906
R17379 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n34 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n24 0.101374
R17380 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n11 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n9 0.101374
R17381 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n254 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n252 0.101374
R17382 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n362 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n360 0.101374
R17383 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n465 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n463 0.101374
R17384 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n568 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n566 0.101374
R17385 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n671 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n669 0.101374
R17386 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n234 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n224 0.101374
R17387 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n207 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n197 0.101374
R17388 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n138 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n128 0.101374
R17389 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n115 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n113 0.101374
R17390 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n91 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n90 0.100442
R17391 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n63 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n62 0.100442
R17392 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n334 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n333 0.100442
R17393 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n306 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n305 0.100442
R17394 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n278 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n277 0.100442
R17395 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n442 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n441 0.100442
R17396 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n414 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n413 0.100442
R17397 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n386 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n385 0.100442
R17398 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n545 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n544 0.100442
R17399 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n517 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n516 0.100442
R17400 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n489 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n488 0.100442
R17401 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n648 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n647 0.100442
R17402 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n620 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n619 0.100442
R17403 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n592 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n591 0.100442
R17404 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n751 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n750 0.100442
R17405 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n723 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n722 0.100442
R17406 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n695 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n694 0.100442
R17407 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n252 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n251 0.0986789
R17408 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n360 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n359 0.0986789
R17409 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n463 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n462 0.0986789
R17410 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n566 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n565 0.0986789
R17411 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n669 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n668 0.0986789
R17412 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n197 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n196 0.0986789
R17413 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n224 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n223 0.0986789
R17414 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n128 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n127 0.0986789
R17415 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n8 0.0986789
R17416 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n90 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n89 0.0937119
R17417 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n62 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n61 0.0937119
R17418 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n333 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n332 0.0937119
R17419 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n305 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n304 0.0937119
R17420 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n277 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n276 0.0937119
R17421 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n441 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n440 0.0937119
R17422 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n413 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n412 0.0937119
R17423 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n385 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n384 0.0937119
R17424 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n544 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n543 0.0937119
R17425 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n516 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n515 0.0937119
R17426 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n488 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n487 0.0937119
R17427 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n647 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n646 0.0937119
R17428 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n619 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n618 0.0937119
R17429 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n591 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n590 0.0937119
R17430 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n750 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n749 0.0937119
R17431 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n722 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n721 0.0937119
R17432 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n694 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n693 0.0937119
R17433 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n24 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n21 0.0930698
R17434 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n161 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n160 0.0826464
R17435 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n176 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n175 0.0826464
R17436 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n768 0.0822606
R17437 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n145 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n141 0.0712285
R17438 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n145 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n144 0.0534597
R17439 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n161 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n156 0.0423164
R17440 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n176 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n171 0.0423164
R17441 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n143 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n142 0.0383947
R17442 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n768 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n4 0.0334577
R17443 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n104 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n103 0.0235313
R17444 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n100 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n99 0.0235313
R17445 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n106 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n105 0.0228651
R17446 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n350 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n349 0.0228651
R17447 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n241 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n108 0.0179841
R17448 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n759 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n664 0.0179841
R17449 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n656 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n561 0.0179841
R17450 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n553 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n458 0.0179841
R17451 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n450 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n355 0.0179841
R17452 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n342 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n247 0.0179841
R17453 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n762 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n761 0.0179841
R17454 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n663 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n662 0.0179841
R17455 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n659 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n658 0.0179841
R17456 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n560 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n559 0.0179841
R17457 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n556 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n555 0.0179841
R17458 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n457 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n456 0.0179841
R17459 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n453 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n452 0.0179841
R17460 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n354 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n353 0.0179841
R17461 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n345 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n344 0.0179841
R17462 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n246 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n245 0.0179841
R17463 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n349 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n348 0.0179841
R17464 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n108 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n107 0.0177304
R17465 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n662 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n661 0.0177304
R17466 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n559 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n558 0.0177304
R17467 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n456 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n455 0.0177304
R17468 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n353 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n352 0.0177304
R17469 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n245 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n244 0.0177304
R17470 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n348 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n347 0.0177304
R17471 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n760 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n663 0.0173591
R17472 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n657 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n560 0.0173591
R17473 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n554 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n457 0.0173591
R17474 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n451 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n354 0.0173591
R17475 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n343 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n246 0.0173591
R17476 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n242 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n104 0.0173591
R17477 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n243 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n242 0.0173591
R17478 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n763 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n760 0.0173591
R17479 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n660 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n657 0.0173591
R17480 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n557 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n554 0.0173591
R17481 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n454 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n451 0.0173591
R17482 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n346 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n343 0.0173591
R17483 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n102 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n101 0.0173591
R17484 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n155 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n154 0.0167343
R17485 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n170 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n169 0.0167343
R17486 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n2 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n1 0.0163451
R17487 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n766 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n765 0.0163451
R17488 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n21 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n20 0.0158007
R17489 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n276 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n275 0.0151658
R17490 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n304 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n303 0.0151658
R17491 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n332 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n331 0.0151658
R17492 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n384 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n383 0.0151658
R17493 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n412 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n411 0.0151658
R17494 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n440 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n439 0.0151658
R17495 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n487 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n486 0.0151658
R17496 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n515 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n514 0.0151658
R17497 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n543 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n542 0.0151658
R17498 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n590 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n589 0.0151658
R17499 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n618 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n617 0.0151658
R17500 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n646 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n645 0.0151658
R17501 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n693 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n692 0.0151658
R17502 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n721 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n720 0.0151658
R17503 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n749 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n748 0.0151658
R17504 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n61 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n60 0.0151658
R17505 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n89 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n88 0.0151658
R17506 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n147 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n146 0.014
R17507 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n101 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n100 0.0122638
R17508 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n107 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n106 0.0119325
R17509 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n351 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n350 0.0119325
R17510 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n765 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n764 0.0112521
R17511 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n251 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n250 0.0111568
R17512 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n359 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n358 0.0111568
R17513 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n462 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n461 0.0111568
R17514 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n565 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n564 0.0111568
R17515 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n668 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n667 0.0111568
R17516 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n196 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n195 0.0111568
R17517 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n223 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n222 0.0111568
R17518 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n127 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n126 0.0111568
R17519 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n7 0.0111568
R17520 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n339 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n338 0.0100339
R17521 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n279 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n255 0.0100339
R17522 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n447 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n446 0.0100339
R17523 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n387 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n363 0.0100339
R17524 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n550 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n549 0.0100339
R17525 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n490 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n466 0.0100339
R17526 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n653 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n652 0.0100339
R17527 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n593 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n569 0.0100339
R17528 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n756 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n755 0.0100339
R17529 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n696 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n672 0.0100339
R17530 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n239 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n238 0.0100339
R17531 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n235 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n211 0.0100339
R17532 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n208 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n184 0.0100339
R17533 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n181 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n180 0.0100339
R17534 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n96 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n95 0.0100339
R17535 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n36 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n35 0.0100339
R17536 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n240 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n239 0.00965254
R17537 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n3 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n2 0.00905634
R17538 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n0 0.00905634
R17539 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n110 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n109 0.00899732
R17540 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n34 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n33 0.00845754
R17541 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n11 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n10 0.00845754
R17542 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n254 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n253 0.00845754
R17543 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n362 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n361 0.00845754
R17544 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n465 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n464 0.00845754
R17545 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n568 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n567 0.00845754
R17546 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n671 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n670 0.00845754
R17547 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n234 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n233 0.00845754
R17548 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n207 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n206 0.00845754
R17549 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n138 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n137 0.00845754
R17550 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n115 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n114 0.00845754
R17551 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n91 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n77 0.00838025
R17552 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n63 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n49 0.00838025
R17553 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n334 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n320 0.00838025
R17554 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n306 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n292 0.00838025
R17555 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n278 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n264 0.00838025
R17556 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n442 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n428 0.00838025
R17557 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n414 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n400 0.00838025
R17558 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n386 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n372 0.00838025
R17559 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n545 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n531 0.00838025
R17560 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n517 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n503 0.00838025
R17561 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n489 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n475 0.00838025
R17562 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n648 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n634 0.00838025
R17563 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n620 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n606 0.00838025
R17564 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n592 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n578 0.00838025
R17565 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n751 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n737 0.00838025
R17566 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n723 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n709 0.00838025
R17567 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n695 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n681 0.00838025
R17568 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n148 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n147 0.00776379
R17569 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n281 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n280 0.00775263
R17570 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n389 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n388 0.00775263
R17571 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n492 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n491 0.00775263
R17572 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n595 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n594 0.00775263
R17573 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n698 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n697 0.00775263
R17574 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n178 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n177 0.00773989
R17575 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n166 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n165 0.00773989
R17576 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n163 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n162 0.00773989
R17577 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n151 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n150 0.00773989
R17578 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n179 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n178 0.00773989
R17579 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n177 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n166 0.00773989
R17580 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n164 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n163 0.00773989
R17581 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n162 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n151 0.00773989
R17582 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n149 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n148 0.00771607
R17583 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n38 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n37 0.00709343
R17584 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n92 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n68 0.00577753
R17585 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n64 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n40 0.00577753
R17586 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n335 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n311 0.00577753
R17587 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n307 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n283 0.00577753
R17588 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n443 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n419 0.00577753
R17589 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n415 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n391 0.00577753
R17590 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n546 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n522 0.00577753
R17591 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n518 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n494 0.00577753
R17592 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n649 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n625 0.00577753
R17593 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n621 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n597 0.00577753
R17594 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n752 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n728 0.00577753
R17595 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n724 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n700 0.00577753
R17596 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n311 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n310 0.00574631
R17597 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n283 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n282 0.00574631
R17598 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n419 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n418 0.00574631
R17599 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n391 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n390 0.00574631
R17600 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n522 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n521 0.00574631
R17601 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n494 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n493 0.00574631
R17602 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n625 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n624 0.00574631
R17603 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n597 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n596 0.00574631
R17604 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n728 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n727 0.00574631
R17605 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n700 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n699 0.00574631
R17606 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n68 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n67 0.00574631
R17607 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n40 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n39 0.00574631
R17608 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n97 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n96 0.00558603
R17609 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n340 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n339 0.00558603
R17610 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n448 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n447 0.00558603
R17611 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n551 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n550 0.00558603
R17612 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n654 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n653 0.00558603
R17613 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n757 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n756 0.00558603
R17614 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n236 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n235 0.00558603
R17615 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n209 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n208 0.00558603
R17616 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n182 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n181 0.00558603
R17617 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n336 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n335 0.00557162
R17618 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n308 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n307 0.00557162
R17619 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n309 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n308 0.00557162
R17620 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n337 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n336 0.00557162
R17621 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n444 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n443 0.00557162
R17622 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n416 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n415 0.00557162
R17623 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n417 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n416 0.00557162
R17624 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n445 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n444 0.00557162
R17625 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n547 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n546 0.00557162
R17626 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n519 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n518 0.00557162
R17627 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n520 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n519 0.00557162
R17628 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n548 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n547 0.00557162
R17629 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n650 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n649 0.00557162
R17630 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n622 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n621 0.00557162
R17631 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n623 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n622 0.00557162
R17632 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n651 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n650 0.00557162
R17633 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n753 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n752 0.00557162
R17634 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n725 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n724 0.00557162
R17635 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n726 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n725 0.00557162
R17636 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n754 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n753 0.00557162
R17637 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n93 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n92 0.00557162
R17638 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n65 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n64 0.00557162
R17639 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n66 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n65 0.00557162
R17640 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n94 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n93 0.00557162
R17641 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n341 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n340 0.00555725
R17642 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n449 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n448 0.00555725
R17643 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n552 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n551 0.00555725
R17644 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n655 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n654 0.00555725
R17645 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n758 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n757 0.00555725
R17646 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n237 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n236 0.00555725
R17647 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n210 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n209 0.00555725
R17648 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n183 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n182 0.00555725
R17649 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n98 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n97 0.00555725
R17650 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n280 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n279 0.00438682
R17651 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n388 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n387 0.00438682
R17652 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n491 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n490 0.00438682
R17653 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n594 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n593 0.00438682
R17654 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n697 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n696 0.00438682
R17655 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n37 Folded_Diff_Op_Amp_Layout_0.IBIAS2.n36 0.00404672
R17656 VOUT_P.n1976 VOUT_P.n1975 11.6357
R17657 VOUT_P.n1103 VOUT_P.t197 6.959
R17658 VOUT_P VOUT_P.t0 4.25918
R17659 VOUT_P.n1106 VOUT_P.n1105 2.40737
R17660 VOUT_P.n1974 VOUT_P.t272 2.38651
R17661 VOUT_P.n1974 VOUT_P.t273 2.2505
R17662 VOUT_P.n1987 VOUT_P.n7 2.24934
R17663 VOUT_P.n5 VOUT_P.n3 2.24889
R17664 VOUT_P.n1984 VOUT_P.n1973 2.24753
R17665 VOUT_P.n1984 VOUT_P.n1979 2.24639
R17666 VOUT_P.n1959 VOUT_P.n1957 2.24505
R17667 VOUT_P.n1985 VOUT_P.n1984 2.2449
R17668 VOUT_P.n1975 VOUT_P.n1974 2.05827
R17669 VOUT_P.n551 VOUT_P.n548 1.84464
R17670 VOUT_P.n930 VOUT_P.n929 1.76234
R17671 VOUT_P.n945 VOUT_P.n944 1.76234
R17672 VOUT_P.n539 VOUT_P.n198 1.49643
R17673 VOUT_P.n448 VOUT_P.n201 1.49371
R17674 VOUT_P.n447 VOUT_P.n203 1.49371
R17675 VOUT_P.n540 VOUT_P.n196 1.49371
R17676 VOUT_P.n973 VOUT_P.n936 1.49371
R17677 VOUT_P.n1923 VOUT_P.n543 1.49371
R17678 VOUT_P.n960 VOUT_P.n959 1.47979
R17679 VOUT_P.n924 VOUT_P.n923 1.47979
R17680 VOUT_P.n939 VOUT_P.n938 1.47979
R17681 VOUT_P.n984 VOUT_P.n983 1.47979
R17682 VOUT_P.n916 VOUT_P.n915 1.47979
R17683 VOUT_P.n908 VOUT_P.n907 1.47979
R17684 VOUT_P.n1460 VOUT_P.n1459 1.46987
R17685 VOUT_P.n1470 VOUT_P.t244 1.46987
R17686 VOUT_P.n1475 VOUT_P.n1474 1.46987
R17687 VOUT_P.n1499 VOUT_P.t249 1.46987
R17688 VOUT_P.n1490 VOUT_P.n1489 1.46987
R17689 VOUT_P.n1485 VOUT_P.t239 1.46987
R17690 VOUT_P.n8 VOUT_P.t213 1.46987
R17691 VOUT_P.n29 VOUT_P.n28 1.46987
R17692 VOUT_P.n134 VOUT_P.t199 1.46987
R17693 VOUT_P.n155 VOUT_P.n154 1.46987
R17694 VOUT_P.n164 VOUT_P.t240 1.46987
R17695 VOUT_P.n185 VOUT_P.n184 1.46987
R17696 VOUT_P.n1707 VOUT_P.n1706 1.43193
R17697 VOUT_P.n1690 VOUT_P.t101 1.43193
R17698 VOUT_P.n1686 VOUT_P.n1685 1.43193
R17699 VOUT_P.n1669 VOUT_P.t193 1.43193
R17700 VOUT_P.n1665 VOUT_P.n1664 1.43193
R17701 VOUT_P.n1648 VOUT_P.t50 1.43193
R17702 VOUT_P.n1644 VOUT_P.n1643 1.43193
R17703 VOUT_P.n1627 VOUT_P.t136 1.43193
R17704 VOUT_P.n1623 VOUT_P.n1622 1.43193
R17705 VOUT_P.n1893 VOUT_P.t22 1.43193
R17706 VOUT_P.n1862 VOUT_P.n1861 1.43193
R17707 VOUT_P.n1852 VOUT_P.t85 1.43193
R17708 VOUT_P.n1821 VOUT_P.n1820 1.43193
R17709 VOUT_P.n1606 VOUT_P.t129 1.43193
R17710 VOUT_P.n714 VOUT_P.n713 1.43193
R17711 VOUT_P.n697 VOUT_P.t173 1.43193
R17712 VOUT_P.n693 VOUT_P.n692 1.43193
R17713 VOUT_P.n676 VOUT_P.t51 1.43193
R17714 VOUT_P.n672 VOUT_P.n671 1.43193
R17715 VOUT_P.n655 VOUT_P.t102 1.43193
R17716 VOUT_P.n651 VOUT_P.n650 1.43193
R17717 VOUT_P.n634 VOUT_P.t186 1.43193
R17718 VOUT_P.n630 VOUT_P.n629 1.43193
R17719 VOUT_P.n613 VOUT_P.t59 1.43193
R17720 VOUT_P.n609 VOUT_P.n608 1.43193
R17721 VOUT_P.n592 VOUT_P.t121 1.43193
R17722 VOUT_P.n588 VOUT_P.n587 1.43193
R17723 VOUT_P.n571 VOUT_P.t45 1.43193
R17724 VOUT_P.n931 VOUT_P.n930 1.3488
R17725 VOUT_P.n946 VOUT_P.n945 1.3488
R17726 VOUT_P.n954 VOUT_P.n953 1.28777
R17727 VOUT_P.n989 VOUT_P.n987 1.28777
R17728 VOUT_P.n563 VOUT_P.n562 1.28752
R17729 VOUT_P.n1072 VOUT_P.n1065 1.26239
R17730 VOUT_P.n957 VOUT_P.n956 1.21718
R17731 VOUT_P.n994 VOUT_P.n993 1.21718
R17732 VOUT_P.n209 VOUT_P.n206 1.19506
R17733 VOUT_P.n219 VOUT_P.n218 1.19506
R17734 VOUT_P.n230 VOUT_P.n229 1.19506
R17735 VOUT_P.n241 VOUT_P.n240 1.19506
R17736 VOUT_P.n267 VOUT_P.n266 1.19506
R17737 VOUT_P.n278 VOUT_P.n277 1.19506
R17738 VOUT_P.n289 VOUT_P.n288 1.19506
R17739 VOUT_P.n300 VOUT_P.n299 1.19506
R17740 VOUT_P.n311 VOUT_P.n310 1.19506
R17741 VOUT_P.n322 VOUT_P.n321 1.19506
R17742 VOUT_P.n333 VOUT_P.n332 1.19506
R17743 VOUT_P.n344 VOUT_P.n343 1.19506
R17744 VOUT_P.n364 VOUT_P.n363 1.19506
R17745 VOUT_P.n375 VOUT_P.n374 1.19506
R17746 VOUT_P.n386 VOUT_P.n385 1.19506
R17747 VOUT_P.n397 VOUT_P.n396 1.19506
R17748 VOUT_P.n408 VOUT_P.n407 1.19506
R17749 VOUT_P.n419 VOUT_P.n418 1.19506
R17750 VOUT_P.n430 VOUT_P.n429 1.19506
R17751 VOUT_P.n441 VOUT_P.n440 1.19506
R17752 VOUT_P.n456 VOUT_P.n455 1.19506
R17753 VOUT_P.n467 VOUT_P.n466 1.19506
R17754 VOUT_P.n478 VOUT_P.n477 1.19506
R17755 VOUT_P.n489 VOUT_P.n488 1.19506
R17756 VOUT_P.n500 VOUT_P.n499 1.19506
R17757 VOUT_P.n511 VOUT_P.n510 1.19506
R17758 VOUT_P.n522 VOUT_P.n521 1.19506
R17759 VOUT_P.n533 VOUT_P.n532 1.19506
R17760 VOUT_P.n1934 VOUT_P.n1933 1.1949
R17761 VOUT_P.n1941 VOUT_P.n1938 1.1949
R17762 VOUT_P.n1300 VOUT_P.n1299 1.1948
R17763 VOUT_P.n1288 VOUT_P.n1287 1.1948
R17764 VOUT_P.n1276 VOUT_P.n1275 1.1948
R17765 VOUT_P.n1264 VOUT_P.n1263 1.1948
R17766 VOUT_P.n1252 VOUT_P.n1251 1.1948
R17767 VOUT_P.n1240 VOUT_P.n1239 1.1948
R17768 VOUT_P.n1228 VOUT_P.n1227 1.1948
R17769 VOUT_P.n1216 VOUT_P.n1215 1.1948
R17770 VOUT_P.n1204 VOUT_P.n1203 1.1948
R17771 VOUT_P.n1192 VOUT_P.n1191 1.1948
R17772 VOUT_P.n1180 VOUT_P.n1179 1.1948
R17773 VOUT_P.n1168 VOUT_P.n1167 1.1948
R17774 VOUT_P.n1156 VOUT_P.n1155 1.1948
R17775 VOUT_P.n1144 VOUT_P.n1143 1.1948
R17776 VOUT_P.n1691 VOUT_P.n1690 1.19473
R17777 VOUT_P.n1670 VOUT_P.n1669 1.19473
R17778 VOUT_P.n1649 VOUT_P.n1648 1.19473
R17779 VOUT_P.n1628 VOUT_P.n1627 1.19473
R17780 VOUT_P.n1607 VOUT_P.n1606 1.19473
R17781 VOUT_P.n715 VOUT_P.n714 1.19473
R17782 VOUT_P.n694 VOUT_P.n693 1.19473
R17783 VOUT_P.n673 VOUT_P.n672 1.19473
R17784 VOUT_P.n652 VOUT_P.n651 1.19473
R17785 VOUT_P.n631 VOUT_P.n630 1.19473
R17786 VOUT_P.n610 VOUT_P.n609 1.19473
R17787 VOUT_P.n589 VOUT_P.n588 1.19473
R17788 VOUT_P.n1114 VOUT_P.n1113 1.19461
R17789 VOUT_P.n1555 VOUT_P.n1554 1.19461
R17790 VOUT_P.n1525 VOUT_P.n1524 1.19461
R17791 VOUT_P.n45 VOUT_P.n44 1.19461
R17792 VOUT_P.n1476 VOUT_P.n1475 1.19458
R17793 VOUT_P.n1486 VOUT_P.n1485 1.19458
R17794 VOUT_P.n9 VOUT_P.n8 1.19458
R17795 VOUT_P.n30 VOUT_P.n29 1.19458
R17796 VOUT_P.n135 VOUT_P.n134 1.19458
R17797 VOUT_P.n156 VOUT_P.n155 1.19458
R17798 VOUT_P.n165 VOUT_P.n164 1.19458
R17799 VOUT_P.n186 VOUT_P.n185 1.19458
R17800 VOUT_P.n76 VOUT_P.n75 1.19458
R17801 VOUT_P.n1703 VOUT_P.n1702 1.19445
R17802 VOUT_P.n1682 VOUT_P.n1681 1.19445
R17803 VOUT_P.n1661 VOUT_P.n1660 1.19445
R17804 VOUT_P.n1640 VOUT_P.n1639 1.19445
R17805 VOUT_P.n1619 VOUT_P.n1618 1.19445
R17806 VOUT_P.n704 VOUT_P.n703 1.19445
R17807 VOUT_P.n683 VOUT_P.n682 1.19445
R17808 VOUT_P.n662 VOUT_P.n661 1.19445
R17809 VOUT_P.n641 VOUT_P.n640 1.19445
R17810 VOUT_P.n620 VOUT_P.n619 1.19445
R17811 VOUT_P.n599 VOUT_P.n598 1.19445
R17812 VOUT_P.n578 VOUT_P.n577 1.19445
R17813 VOUT_P.n1467 VOUT_P.n1466 1.19426
R17814 VOUT_P.n1497 VOUT_P.n1496 1.19426
R17815 VOUT_P.n20 VOUT_P.n19 1.19426
R17816 VOUT_P.n146 VOUT_P.n145 1.19426
R17817 VOUT_P.n176 VOUT_P.n175 1.19426
R17818 VOUT_P.n1097 VOUT_P.n1096 1.18729
R17819 VOUT_P.n1482 VOUT_P.n1481 1.17959
R17820 VOUT_P.n1461 VOUT_P.n1460 1.1793
R17821 VOUT_P.n1471 VOUT_P.n1470 1.1793
R17822 VOUT_P.n1502 VOUT_P.n1499 1.1793
R17823 VOUT_P.n1491 VOUT_P.n1490 1.1793
R17824 VOUT_P.n1697 VOUT_P.n1696 1.1791
R17825 VOUT_P.n1676 VOUT_P.n1675 1.1791
R17826 VOUT_P.n1655 VOUT_P.n1654 1.1791
R17827 VOUT_P.n1634 VOUT_P.n1633 1.1791
R17828 VOUT_P.n1613 VOUT_P.n1612 1.1791
R17829 VOUT_P.n1885 VOUT_P.n1884 1.1791
R17830 VOUT_P.n1874 VOUT_P.n1873 1.1791
R17831 VOUT_P.n1844 VOUT_P.n1843 1.1791
R17832 VOUT_P.n1833 VOUT_P.n1832 1.1791
R17833 VOUT_P.n710 VOUT_P.n709 1.1791
R17834 VOUT_P.n689 VOUT_P.n688 1.1791
R17835 VOUT_P.n668 VOUT_P.n667 1.1791
R17836 VOUT_P.n647 VOUT_P.n646 1.1791
R17837 VOUT_P.n626 VOUT_P.n625 1.1791
R17838 VOUT_P.n605 VOUT_P.n604 1.1791
R17839 VOUT_P.n584 VOUT_P.n583 1.1791
R17840 VOUT_P.n1120 VOUT_P.n1119 1.17896
R17841 VOUT_P.n1531 VOUT_P.n1530 1.17896
R17842 VOUT_P.n1549 VOUT_P.n1548 1.17896
R17843 VOUT_P.n51 VOUT_P.n50 1.17896
R17844 VOUT_P.n69 VOUT_P.n68 1.17896
R17845 VOUT_P.n1708 VOUT_P.n1707 1.17884
R17846 VOUT_P.n1687 VOUT_P.n1686 1.17884
R17847 VOUT_P.n1666 VOUT_P.n1665 1.17884
R17848 VOUT_P.n1645 VOUT_P.n1644 1.17884
R17849 VOUT_P.n1624 VOUT_P.n1623 1.17884
R17850 VOUT_P.n1894 VOUT_P.n1893 1.17884
R17851 VOUT_P.n1863 VOUT_P.n1862 1.17884
R17852 VOUT_P.n1853 VOUT_P.n1852 1.17884
R17853 VOUT_P.n1822 VOUT_P.n1821 1.17884
R17854 VOUT_P.n698 VOUT_P.n697 1.17884
R17855 VOUT_P.n677 VOUT_P.n676 1.17884
R17856 VOUT_P.n656 VOUT_P.n655 1.17884
R17857 VOUT_P.n635 VOUT_P.n634 1.17884
R17858 VOUT_P.n614 VOUT_P.n613 1.17884
R17859 VOUT_P.n593 VOUT_P.n592 1.17884
R17860 VOUT_P.n572 VOUT_P.n571 1.17884
R17861 VOUT_P.n1294 VOUT_P.n1293 1.17849
R17862 VOUT_P.n1282 VOUT_P.n1281 1.17849
R17863 VOUT_P.n1270 VOUT_P.n1269 1.17849
R17864 VOUT_P.n1258 VOUT_P.n1257 1.17849
R17865 VOUT_P.n1246 VOUT_P.n1245 1.17849
R17866 VOUT_P.n1234 VOUT_P.n1233 1.17849
R17867 VOUT_P.n1222 VOUT_P.n1221 1.17849
R17868 VOUT_P.n1210 VOUT_P.n1209 1.17849
R17869 VOUT_P.n1198 VOUT_P.n1197 1.17849
R17870 VOUT_P.n1186 VOUT_P.n1185 1.17849
R17871 VOUT_P.n1174 VOUT_P.n1173 1.17849
R17872 VOUT_P.n1162 VOUT_P.n1161 1.17849
R17873 VOUT_P.n1150 VOUT_P.n1149 1.17849
R17874 VOUT_P.n1138 VOUT_P.n1137 1.17849
R17875 VOUT_P.n989 VOUT_P.n988 1.1742
R17876 VOUT_P.n564 VOUT_P.n563 1.17419
R17877 VOUT_P.n552 VOUT_P.n551 1.14437
R17878 VOUT_P.n925 VOUT_P.n924 1.14073
R17879 VOUT_P.n940 VOUT_P.n939 1.14073
R17880 VOUT_P.n985 VOUT_P.n984 1.14073
R17881 VOUT_P.n917 VOUT_P.n916 1.14073
R17882 VOUT_P.n909 VOUT_P.n908 1.14073
R17883 VOUT_P.n356 VOUT_P.n355 1.1353
R17884 VOUT_P.n1928 VOUT_P.n1927 1.12925
R17885 VOUT_P.n210 VOUT_P.n209 1.12829
R17886 VOUT_P.n107 VOUT_P.n106 1.12829
R17887 VOUT_P.n553 VOUT_P.n552 1.12829
R17888 VOUT_P.n1503 VOUT_P.n1502 1.12829
R17889 VOUT_P.n1942 VOUT_P.n1941 1.12795
R17890 VOUT_P.n963 VOUT_P.n962 1.12795
R17891 VOUT_P.n77 VOUT_P.n76 1.12758
R17892 VOUT_P.n962 VOUT_P.n961 1.1255
R17893 VOUT_P.n933 VOUT_P.n932 1.1255
R17894 VOUT_P.n948 VOUT_P.n947 1.1255
R17895 VOUT_P.n992 VOUT_P.n991 1.1255
R17896 VOUT_P.n996 VOUT_P.n995 1.1255
R17897 VOUT_P.n920 VOUT_P.n919 1.1255
R17898 VOUT_P.n560 VOUT_P.n559 1.1255
R17899 VOUT_P.n912 VOUT_P.n911 1.1255
R17900 VOUT_P.n1064 VOUT_P.n1063 1.12145
R17901 VOUT_P.n1064 VOUT_P.n1059 1.12145
R17902 VOUT_P.n1054 VOUT_P.n1051 1.12145
R17903 VOUT_P.n1054 VOUT_P.n1053 1.12145
R17904 VOUT_P.n1095 VOUT_P.n1094 1.12145
R17905 VOUT_P.n1088 VOUT_P.n1087 1.12145
R17906 VOUT_P.n904 VOUT_P.n903 1.11801
R17907 VOUT_P.n844 VOUT_P.n843 1.11801
R17908 VOUT_P.n847 VOUT_P.n846 1.11801
R17909 VOUT_P.n123 VOUT_P.n116 1.11801
R17910 VOUT_P.n260 VOUT_P.n259 1.11801
R17911 VOUT_P.n1327 VOUT_P.n1326 1.11801
R17912 VOUT_P.n1909 VOUT_P.n1012 1.11801
R17913 VOUT_P.n1915 VOUT_P.n569 1.11801
R17914 VOUT_P.n1953 VOUT_P.n1952 1.11801
R17915 VOUT_P.n1603 VOUT_P.n1602 1.11801
R17916 VOUT_P.n1105 VOUT_P.n1098 1.11801
R17917 VOUT_P.n793 VOUT_P.n792 1.11782
R17918 VOUT_P.n87 VOUT_P.n86 1.11782
R17919 VOUT_P.n130 VOUT_P.n129 1.11782
R17920 VOUT_P.n1567 VOUT_P.n1566 1.11782
R17921 VOUT_P.n1543 VOUT_P.n1542 1.11782
R17922 VOUT_P.n62 VOUT_P.n61 1.11782
R17923 VOUT_P.n1573 VOUT_P.n1572 1.11782
R17924 VOUT_P.n1735 VOUT_P.n1734 1.11782
R17925 VOUT_P.n1324 VOUT_P.n1323 1.11782
R17926 VOUT_P.n1453 VOUT_P.n1452 1.11782
R17927 VOUT_P.n1132 VOUT_P.n1131 1.11782
R17928 VOUT_P.n1914 VOUT_P.n1913 1.11782
R17929 VOUT_P.n1905 VOUT_P.n1904 1.11782
R17930 VOUT_P.n1104 VOUT_P.n1103 1.11782
R17931 VOUT_P.n1975 VOUT_P 1.06273
R17932 VOUT_P.n1000 VOUT_P.n999 1.03835
R17933 VOUT_P.n75 VOUT_P.n74 0.923874
R17934 VOUT_P.n1113 VOUT_P.n1112 0.923611
R17935 VOUT_P.n1554 VOUT_P.n1553 0.923611
R17936 VOUT_P.n1524 VOUT_P.n1523 0.923611
R17937 VOUT_P.n44 VOUT_P.n43 0.923611
R17938 VOUT_P.n1933 VOUT_P.n1932 0.923589
R17939 VOUT_P.n1938 VOUT_P.n1937 0.923589
R17940 VOUT_P.n1119 VOUT_P.n1118 0.923589
R17941 VOUT_P.n1530 VOUT_P.n1529 0.923589
R17942 VOUT_P.n1548 VOUT_P.n1547 0.923589
R17943 VOUT_P.n50 VOUT_P.n49 0.923589
R17944 VOUT_P.n68 VOUT_P.n67 0.923589
R17945 VOUT_P.n1466 VOUT_P.n1465 0.923538
R17946 VOUT_P.n1481 VOUT_P.n1480 0.923538
R17947 VOUT_P.n1496 VOUT_P.n1495 0.923538
R17948 VOUT_P.n19 VOUT_P.n18 0.923538
R17949 VOUT_P.n145 VOUT_P.n144 0.923538
R17950 VOUT_P.n175 VOUT_P.n174 0.923538
R17951 VOUT_P.n1948 VOUT_P.n1935 0.885703
R17952 VOUT_P.n566 VOUT_P.n565 0.885703
R17953 VOUT_P.n535 VOUT_P.n534 0.885703
R17954 VOUT_P.n524 VOUT_P.n523 0.885703
R17955 VOUT_P.n513 VOUT_P.n512 0.885703
R17956 VOUT_P.n502 VOUT_P.n501 0.885703
R17957 VOUT_P.n491 VOUT_P.n490 0.885703
R17958 VOUT_P.n480 VOUT_P.n479 0.885703
R17959 VOUT_P.n469 VOUT_P.n468 0.885703
R17960 VOUT_P.n458 VOUT_P.n457 0.885703
R17961 VOUT_P.n443 VOUT_P.n442 0.885703
R17962 VOUT_P.n432 VOUT_P.n431 0.885703
R17963 VOUT_P.n421 VOUT_P.n420 0.885703
R17964 VOUT_P.n410 VOUT_P.n409 0.885703
R17965 VOUT_P.n399 VOUT_P.n398 0.885703
R17966 VOUT_P.n388 VOUT_P.n387 0.885703
R17967 VOUT_P.n377 VOUT_P.n376 0.885703
R17968 VOUT_P.n366 VOUT_P.n365 0.885703
R17969 VOUT_P.n346 VOUT_P.n345 0.885703
R17970 VOUT_P.n335 VOUT_P.n334 0.885703
R17971 VOUT_P.n324 VOUT_P.n323 0.885703
R17972 VOUT_P.n313 VOUT_P.n312 0.885703
R17973 VOUT_P.n302 VOUT_P.n301 0.885703
R17974 VOUT_P.n291 VOUT_P.n290 0.885703
R17975 VOUT_P.n280 VOUT_P.n279 0.885703
R17976 VOUT_P.n269 VOUT_P.n268 0.885703
R17977 VOUT_P.n243 VOUT_P.n242 0.885703
R17978 VOUT_P.n232 VOUT_P.n231 0.885703
R17979 VOUT_P.n221 VOUT_P.n220 0.885703
R17980 VOUT_P.n1824 VOUT_P.n1823 0.885703
R17981 VOUT_P.n1835 VOUT_P.n1834 0.885703
R17982 VOUT_P.n1846 VOUT_P.n1845 0.885703
R17983 VOUT_P.n1855 VOUT_P.n1854 0.885703
R17984 VOUT_P.n1865 VOUT_P.n1864 0.885703
R17985 VOUT_P.n1876 VOUT_P.n1875 0.885703
R17986 VOUT_P.n1887 VOUT_P.n1886 0.885703
R17987 VOUT_P.n1896 VOUT_P.n1895 0.885703
R17988 VOUT_P.n162 VOUT_P.n161 0.835535
R17989 VOUT_P.n1588 VOUT_P.n1587 0.835535
R17990 VOUT_P.n1299 VOUT_P.n1298 0.824999
R17991 VOUT_P.n1287 VOUT_P.n1286 0.824999
R17992 VOUT_P.n1275 VOUT_P.n1274 0.824999
R17993 VOUT_P.n1263 VOUT_P.n1262 0.824999
R17994 VOUT_P.n1251 VOUT_P.n1250 0.824999
R17995 VOUT_P.n1239 VOUT_P.n1238 0.824999
R17996 VOUT_P.n1227 VOUT_P.n1226 0.824999
R17997 VOUT_P.n1215 VOUT_P.n1214 0.824999
R17998 VOUT_P.n1203 VOUT_P.n1202 0.824999
R17999 VOUT_P.n1191 VOUT_P.n1190 0.824999
R18000 VOUT_P.n1179 VOUT_P.n1178 0.824999
R18001 VOUT_P.n1167 VOUT_P.n1166 0.824999
R18002 VOUT_P.n1155 VOUT_P.n1154 0.824999
R18003 VOUT_P.n1143 VOUT_P.n1142 0.824999
R18004 VOUT_P.n1293 VOUT_P.n1292 0.824997
R18005 VOUT_P.n206 VOUT_P.n205 0.824997
R18006 VOUT_P.n218 VOUT_P.n217 0.824997
R18007 VOUT_P.n229 VOUT_P.n228 0.824997
R18008 VOUT_P.n240 VOUT_P.n239 0.824997
R18009 VOUT_P.n266 VOUT_P.n265 0.824997
R18010 VOUT_P.n277 VOUT_P.n276 0.824997
R18011 VOUT_P.n288 VOUT_P.n287 0.824997
R18012 VOUT_P.n299 VOUT_P.n298 0.824997
R18013 VOUT_P.n310 VOUT_P.n309 0.824997
R18014 VOUT_P.n321 VOUT_P.n320 0.824997
R18015 VOUT_P.n332 VOUT_P.n331 0.824997
R18016 VOUT_P.n343 VOUT_P.n342 0.824997
R18017 VOUT_P.n363 VOUT_P.n362 0.824997
R18018 VOUT_P.n374 VOUT_P.n373 0.824997
R18019 VOUT_P.n385 VOUT_P.n384 0.824997
R18020 VOUT_P.n396 VOUT_P.n395 0.824997
R18021 VOUT_P.n407 VOUT_P.n406 0.824997
R18022 VOUT_P.n418 VOUT_P.n417 0.824997
R18023 VOUT_P.n429 VOUT_P.n428 0.824997
R18024 VOUT_P.n440 VOUT_P.n439 0.824997
R18025 VOUT_P.n455 VOUT_P.n454 0.824997
R18026 VOUT_P.n466 VOUT_P.n465 0.824997
R18027 VOUT_P.n477 VOUT_P.n476 0.824997
R18028 VOUT_P.n488 VOUT_P.n487 0.824997
R18029 VOUT_P.n499 VOUT_P.n498 0.824997
R18030 VOUT_P.n510 VOUT_P.n509 0.824997
R18031 VOUT_P.n521 VOUT_P.n520 0.824997
R18032 VOUT_P.n532 VOUT_P.n531 0.824997
R18033 VOUT_P.n1281 VOUT_P.n1280 0.824997
R18034 VOUT_P.n1269 VOUT_P.n1268 0.824997
R18035 VOUT_P.n1257 VOUT_P.n1256 0.824997
R18036 VOUT_P.n1245 VOUT_P.n1244 0.824997
R18037 VOUT_P.n1233 VOUT_P.n1232 0.824997
R18038 VOUT_P.n1221 VOUT_P.n1220 0.824997
R18039 VOUT_P.n1209 VOUT_P.n1208 0.824997
R18040 VOUT_P.n1197 VOUT_P.n1196 0.824997
R18041 VOUT_P.n1185 VOUT_P.n1184 0.824997
R18042 VOUT_P.n1173 VOUT_P.n1172 0.824997
R18043 VOUT_P.n1161 VOUT_P.n1160 0.824997
R18044 VOUT_P.n1149 VOUT_P.n1148 0.824997
R18045 VOUT_P.n1137 VOUT_P.n1136 0.824997
R18046 VOUT_P.n1702 VOUT_P.n1701 0.82495
R18047 VOUT_P.n1696 VOUT_P.n1695 0.82495
R18048 VOUT_P.n1681 VOUT_P.n1680 0.82495
R18049 VOUT_P.n1675 VOUT_P.n1674 0.82495
R18050 VOUT_P.n1660 VOUT_P.n1659 0.82495
R18051 VOUT_P.n1654 VOUT_P.n1653 0.82495
R18052 VOUT_P.n1639 VOUT_P.n1638 0.82495
R18053 VOUT_P.n1633 VOUT_P.n1632 0.82495
R18054 VOUT_P.n1618 VOUT_P.n1617 0.82495
R18055 VOUT_P.n1612 VOUT_P.n1611 0.82495
R18056 VOUT_P.n1884 VOUT_P.n1883 0.82495
R18057 VOUT_P.n1873 VOUT_P.n1872 0.82495
R18058 VOUT_P.n1843 VOUT_P.n1842 0.82495
R18059 VOUT_P.n1832 VOUT_P.n1831 0.82495
R18060 VOUT_P.n709 VOUT_P.n708 0.82495
R18061 VOUT_P.n703 VOUT_P.n702 0.82495
R18062 VOUT_P.n688 VOUT_P.n687 0.82495
R18063 VOUT_P.n682 VOUT_P.n681 0.82495
R18064 VOUT_P.n667 VOUT_P.n666 0.82495
R18065 VOUT_P.n661 VOUT_P.n660 0.82495
R18066 VOUT_P.n646 VOUT_P.n645 0.82495
R18067 VOUT_P.n640 VOUT_P.n639 0.82495
R18068 VOUT_P.n625 VOUT_P.n624 0.82495
R18069 VOUT_P.n619 VOUT_P.n618 0.82495
R18070 VOUT_P.n604 VOUT_P.n603 0.82495
R18071 VOUT_P.n598 VOUT_P.n597 0.82495
R18072 VOUT_P.n583 VOUT_P.n582 0.82495
R18073 VOUT_P.n577 VOUT_P.n576 0.82495
R18074 VOUT_P.n1070 VOUT_P.n1069 0.736598
R18075 VOUT_P.n13 VOUT_P.n11 0.727916
R18076 VOUT_P.n23 VOUT_P.n22 0.727916
R18077 VOUT_P.n33 VOUT_P.n32 0.727916
R18078 VOUT_P.n138 VOUT_P.n137 0.727916
R18079 VOUT_P.n149 VOUT_P.n148 0.727916
R18080 VOUT_P.n159 VOUT_P.n158 0.727916
R18081 VOUT_P.n168 VOUT_P.n167 0.727916
R18082 VOUT_P.n179 VOUT_P.n178 0.727916
R18083 VOUT_P.n189 VOUT_P.n188 0.727916
R18084 VOUT_P.n1539 VOUT_P.n1526 0.727104
R18085 VOUT_P.n1558 VOUT_P.n1556 0.727104
R18086 VOUT_P.n977 VOUT_P.n934 0.727104
R18087 VOUT_P.n1002 VOUT_P.n921 0.727104
R18088 VOUT_P.n969 VOUT_P.n949 0.727104
R18089 VOUT_P.n722 VOUT_P.n711 0.727104
R18090 VOUT_P.n731 VOUT_P.n699 0.727104
R18091 VOUT_P.n744 VOUT_P.n690 0.727104
R18092 VOUT_P.n753 VOUT_P.n678 0.727104
R18093 VOUT_P.n762 VOUT_P.n669 0.727104
R18094 VOUT_P.n771 VOUT_P.n657 0.727104
R18095 VOUT_P.n800 VOUT_P.n648 0.727104
R18096 VOUT_P.n809 VOUT_P.n636 0.727104
R18097 VOUT_P.n818 VOUT_P.n627 0.727104
R18098 VOUT_P.n827 VOUT_P.n615 0.727104
R18099 VOUT_P.n855 VOUT_P.n606 0.727104
R18100 VOUT_P.n864 VOUT_P.n594 0.727104
R18101 VOUT_P.n873 VOUT_P.n585 0.727104
R18102 VOUT_P.n882 VOUT_P.n573 0.727104
R18103 VOUT_P.n58 VOUT_P.n46 0.727104
R18104 VOUT_P.n1512 VOUT_P.n1492 0.727104
R18105 VOUT_P.n1599 VOUT_P.n1462 0.727104
R18106 VOUT_P.n1590 VOUT_P.n1472 0.727104
R18107 VOUT_P.n1581 VOUT_P.n1483 0.727104
R18108 VOUT_P.n1711 VOUT_P.n1709 0.727104
R18109 VOUT_P.n1720 VOUT_P.n1698 0.727104
R18110 VOUT_P.n1739 VOUT_P.n1688 0.727104
R18111 VOUT_P.n1748 VOUT_P.n1677 0.727104
R18112 VOUT_P.n1757 VOUT_P.n1667 0.727104
R18113 VOUT_P.n1766 VOUT_P.n1656 0.727104
R18114 VOUT_P.n1779 VOUT_P.n1646 0.727104
R18115 VOUT_P.n1788 VOUT_P.n1635 0.727104
R18116 VOUT_P.n1797 VOUT_P.n1625 0.727104
R18117 VOUT_P.n1806 VOUT_P.n1614 0.727104
R18118 VOUT_P.n1128 VOUT_P.n1115 0.727104
R18119 VOUT_P.n1303 VOUT_P.n1301 0.727104
R18120 VOUT_P.n1312 VOUT_P.n1289 0.727104
R18121 VOUT_P.n1330 VOUT_P.n1277 0.727104
R18122 VOUT_P.n1339 VOUT_P.n1265 0.727104
R18123 VOUT_P.n1348 VOUT_P.n1253 0.727104
R18124 VOUT_P.n1357 VOUT_P.n1241 0.727104
R18125 VOUT_P.n1371 VOUT_P.n1229 0.727104
R18126 VOUT_P.n1380 VOUT_P.n1217 0.727104
R18127 VOUT_P.n1389 VOUT_P.n1205 0.727104
R18128 VOUT_P.n1398 VOUT_P.n1193 0.727104
R18129 VOUT_P.n1412 VOUT_P.n1181 0.727104
R18130 VOUT_P.n1421 VOUT_P.n1169 0.727104
R18131 VOUT_P.n1430 VOUT_P.n1157 0.727104
R18132 VOUT_P.n1439 VOUT_P.n1145 0.727104
R18133 VOUT_P.n112 VOUT_P.n103 0.726858
R18134 VOUT_P.n1007 VOUT_P.n913 0.726858
R18135 VOUT_P.n1954 VOUT_P.n1953 0.696042
R18136 VOUT_P.n305 VOUT_P.n304 0.685007
R18137 VOUT_P.n402 VOUT_P.n401 0.685007
R18138 VOUT_P.n494 VOUT_P.n493 0.685007
R18139 VOUT_P.n1346 VOUT_P.n1345 0.685007
R18140 VOUT_P.n1387 VOUT_P.n1386 0.685007
R18141 VOUT_P.n1428 VOUT_P.n1427 0.685007
R18142 VOUT_P.n1951 VOUT_P.n1950 0.673915
R18143 VOUT_P.n1565 VOUT_P.n1564 0.673915
R18144 VOUT_P.n1542 VOUT_P.n1541 0.673915
R18145 VOUT_P.n99 VOUT_P.n98 0.673915
R18146 VOUT_P.n115 VOUT_P.n114 0.673915
R18147 VOUT_P.n569 VOUT_P.n568 0.673915
R18148 VOUT_P.n1010 VOUT_P.n1009 0.673915
R18149 VOUT_P.n975 VOUT_P.n974 0.673915
R18150 VOUT_P.n972 VOUT_P.n971 0.673915
R18151 VOUT_P.n61 VOUT_P.n60 0.673915
R18152 VOUT_P.n85 VOUT_P.n84 0.673915
R18153 VOUT_P.n1131 VOUT_P.n1130 0.673915
R18154 VOUT_P.n998 VOUT_P.n997 0.617177
R18155 VOUT_P.n1308 VOUT_P.n1295 0.616779
R18156 VOUT_P.n1123 VOUT_P.n1121 0.616779
R18157 VOUT_P.n1716 VOUT_P.n1704 0.616779
R18158 VOUT_P.n1725 VOUT_P.n1692 0.616779
R18159 VOUT_P.n1744 VOUT_P.n1683 0.616779
R18160 VOUT_P.n1753 VOUT_P.n1671 0.616779
R18161 VOUT_P.n1762 VOUT_P.n1662 0.616779
R18162 VOUT_P.n1771 VOUT_P.n1650 0.616779
R18163 VOUT_P.n1784 VOUT_P.n1641 0.616779
R18164 VOUT_P.n1793 VOUT_P.n1629 0.616779
R18165 VOUT_P.n1802 VOUT_P.n1620 0.616779
R18166 VOUT_P.n1811 VOUT_P.n1608 0.616779
R18167 VOUT_P.n1594 VOUT_P.n1468 0.616779
R18168 VOUT_P.n1585 VOUT_P.n1477 0.616779
R18169 VOUT_P.n1507 VOUT_P.n1498 0.616779
R18170 VOUT_P.n1576 VOUT_P.n1487 0.616779
R18171 VOUT_P.n1534 VOUT_P.n1532 0.616779
R18172 VOUT_P.n1563 VOUT_P.n1550 0.616779
R18173 VOUT_P.n718 VOUT_P.n716 0.616779
R18174 VOUT_P.n727 VOUT_P.n705 0.616779
R18175 VOUT_P.n740 VOUT_P.n695 0.616779
R18176 VOUT_P.n749 VOUT_P.n684 0.616779
R18177 VOUT_P.n758 VOUT_P.n674 0.616779
R18178 VOUT_P.n767 VOUT_P.n663 0.616779
R18179 VOUT_P.n796 VOUT_P.n653 0.616779
R18180 VOUT_P.n805 VOUT_P.n642 0.616779
R18181 VOUT_P.n814 VOUT_P.n632 0.616779
R18182 VOUT_P.n823 VOUT_P.n621 0.616779
R18183 VOUT_P.n851 VOUT_P.n611 0.616779
R18184 VOUT_P.n860 VOUT_P.n600 0.616779
R18185 VOUT_P.n869 VOUT_P.n590 0.616779
R18186 VOUT_P.n878 VOUT_P.n579 0.616779
R18187 VOUT_P.n97 VOUT_P.n90 0.616779
R18188 VOUT_P.n54 VOUT_P.n52 0.616779
R18189 VOUT_P.n82 VOUT_P.n70 0.616779
R18190 VOUT_P.n1317 VOUT_P.n1283 0.616779
R18191 VOUT_P.n1335 VOUT_P.n1271 0.616779
R18192 VOUT_P.n1344 VOUT_P.n1259 0.616779
R18193 VOUT_P.n1353 VOUT_P.n1247 0.616779
R18194 VOUT_P.n1362 VOUT_P.n1235 0.616779
R18195 VOUT_P.n1376 VOUT_P.n1223 0.616779
R18196 VOUT_P.n1385 VOUT_P.n1211 0.616779
R18197 VOUT_P.n1394 VOUT_P.n1199 0.616779
R18198 VOUT_P.n1403 VOUT_P.n1187 0.616779
R18199 VOUT_P.n1417 VOUT_P.n1175 0.616779
R18200 VOUT_P.n1426 VOUT_P.n1163 0.616779
R18201 VOUT_P.n1435 VOUT_P.n1151 0.616779
R18202 VOUT_P.n1444 VOUT_P.n1139 0.616779
R18203 VOUT_P.n1298 VOUT_P.t156 0.607167
R18204 VOUT_P.n1298 VOUT_P.n1297 0.607167
R18205 VOUT_P.n1292 VOUT_P.t174 0.607167
R18206 VOUT_P.n1292 VOUT_P.n1291 0.607167
R18207 VOUT_P.n1286 VOUT_P.t109 0.607167
R18208 VOUT_P.n1286 VOUT_P.n1285 0.607167
R18209 VOUT_P.n1701 VOUT_P.t60 0.607167
R18210 VOUT_P.n1701 VOUT_P.n1700 0.607167
R18211 VOUT_P.n1695 VOUT_P.t19 0.607167
R18212 VOUT_P.n1695 VOUT_P.n1694 0.607167
R18213 VOUT_P.n1680 VOUT_P.t167 0.607167
R18214 VOUT_P.n1680 VOUT_P.n1679 0.607167
R18215 VOUT_P.n1674 VOUT_P.t120 0.607167
R18216 VOUT_P.n1674 VOUT_P.n1673 0.607167
R18217 VOUT_P.n1659 VOUT_P.t8 0.607167
R18218 VOUT_P.n1659 VOUT_P.n1658 0.607167
R18219 VOUT_P.n1653 VOUT_P.t166 0.607167
R18220 VOUT_P.n1653 VOUT_P.n1652 0.607167
R18221 VOUT_P.n1638 VOUT_P.t41 0.607167
R18222 VOUT_P.n1638 VOUT_P.n1637 0.607167
R18223 VOUT_P.n1632 VOUT_P.t67 0.607167
R18224 VOUT_P.n1632 VOUT_P.n1631 0.607167
R18225 VOUT_P.n1617 VOUT_P.t90 0.607167
R18226 VOUT_P.n1617 VOUT_P.n1616 0.607167
R18227 VOUT_P.n1611 VOUT_P.t111 0.607167
R18228 VOUT_P.n1611 VOUT_P.n1610 0.607167
R18229 VOUT_P.n1883 VOUT_P.t141 0.607167
R18230 VOUT_P.n1883 VOUT_P.n1882 0.607167
R18231 VOUT_P.n1872 VOUT_P.t183 0.607167
R18232 VOUT_P.n1872 VOUT_P.n1871 0.607167
R18233 VOUT_P.n1842 VOUT_P.t147 0.607167
R18234 VOUT_P.n1842 VOUT_P.n1841 0.607167
R18235 VOUT_P.n1831 VOUT_P.t192 0.607167
R18236 VOUT_P.n1831 VOUT_P.n1830 0.607167
R18237 VOUT_P.n205 VOUT_P.t117 0.607167
R18238 VOUT_P.n205 VOUT_P.n204 0.607167
R18239 VOUT_P.n217 VOUT_P.t87 0.607167
R18240 VOUT_P.n217 VOUT_P.n216 0.607167
R18241 VOUT_P.n228 VOUT_P.t158 0.607167
R18242 VOUT_P.n228 VOUT_P.n227 0.607167
R18243 VOUT_P.n239 VOUT_P.t30 0.607167
R18244 VOUT_P.n239 VOUT_P.n238 0.607167
R18245 VOUT_P.n265 VOUT_P.t66 0.607167
R18246 VOUT_P.n265 VOUT_P.n264 0.607167
R18247 VOUT_P.n276 VOUT_P.t144 0.607167
R18248 VOUT_P.n276 VOUT_P.n275 0.607167
R18249 VOUT_P.n287 VOUT_P.t86 0.607167
R18250 VOUT_P.n287 VOUT_P.n286 0.607167
R18251 VOUT_P.n298 VOUT_P.t180 0.607167
R18252 VOUT_P.n298 VOUT_P.n297 0.607167
R18253 VOUT_P.n309 VOUT_P.t79 0.607167
R18254 VOUT_P.n309 VOUT_P.n308 0.607167
R18255 VOUT_P.n320 VOUT_P.t17 0.607167
R18256 VOUT_P.n320 VOUT_P.n319 0.607167
R18257 VOUT_P.n331 VOUT_P.t95 0.607167
R18258 VOUT_P.n331 VOUT_P.n330 0.607167
R18259 VOUT_P.n342 VOUT_P.t188 0.607167
R18260 VOUT_P.n342 VOUT_P.n341 0.607167
R18261 VOUT_P.n362 VOUT_P.t3 0.607167
R18262 VOUT_P.n362 VOUT_P.n361 0.607167
R18263 VOUT_P.n373 VOUT_P.t78 0.607167
R18264 VOUT_P.n373 VOUT_P.n372 0.607167
R18265 VOUT_P.n384 VOUT_P.t37 0.607167
R18266 VOUT_P.n384 VOUT_P.n383 0.607167
R18267 VOUT_P.n395 VOUT_P.t113 0.607167
R18268 VOUT_P.n395 VOUT_P.n394 0.607167
R18269 VOUT_P.n406 VOUT_P.t10 0.607167
R18270 VOUT_P.n406 VOUT_P.n405 0.607167
R18271 VOUT_P.n417 VOUT_P.t154 0.607167
R18272 VOUT_P.n417 VOUT_P.n416 0.607167
R18273 VOUT_P.n428 VOUT_P.t47 0.607167
R18274 VOUT_P.n428 VOUT_P.n427 0.607167
R18275 VOUT_P.n439 VOUT_P.t123 0.607167
R18276 VOUT_P.n439 VOUT_P.n438 0.607167
R18277 VOUT_P.n454 VOUT_P.t137 0.607167
R18278 VOUT_P.n454 VOUT_P.n453 0.607167
R18279 VOUT_P.n465 VOUT_P.t33 0.607167
R18280 VOUT_P.n465 VOUT_P.n464 0.607167
R18281 VOUT_P.n476 VOUT_P.t178 0.607167
R18282 VOUT_P.n476 VOUT_P.n475 0.607167
R18283 VOUT_P.n487 VOUT_P.t46 0.607167
R18284 VOUT_P.n487 VOUT_P.n486 0.607167
R18285 VOUT_P.n498 VOUT_P.t1 0.607167
R18286 VOUT_P.n498 VOUT_P.n497 0.607167
R18287 VOUT_P.n509 VOUT_P.t160 0.607167
R18288 VOUT_P.n509 VOUT_P.n508 0.607167
R18289 VOUT_P.n520 VOUT_P.t35 0.607167
R18290 VOUT_P.n520 VOUT_P.n519 0.607167
R18291 VOUT_P.n531 VOUT_P.t106 0.607167
R18292 VOUT_P.n531 VOUT_P.n530 0.607167
R18293 VOUT_P.n708 VOUT_P.t195 0.607167
R18294 VOUT_P.n708 VOUT_P.n707 0.607167
R18295 VOUT_P.n702 VOUT_P.t29 0.607167
R18296 VOUT_P.n702 VOUT_P.n701 0.607167
R18297 VOUT_P.n687 VOUT_P.t116 0.607167
R18298 VOUT_P.n687 VOUT_P.n686 0.607167
R18299 VOUT_P.n681 VOUT_P.t157 0.607167
R18300 VOUT_P.n681 VOUT_P.n680 0.607167
R18301 VOUT_P.n666 VOUT_P.t127 0.607167
R18302 VOUT_P.n666 VOUT_P.n665 0.607167
R18303 VOUT_P.n660 VOUT_P.t163 0.607167
R18304 VOUT_P.n660 VOUT_P.n659 0.607167
R18305 VOUT_P.n645 VOUT_P.t76 0.607167
R18306 VOUT_P.n645 VOUT_P.n644 0.607167
R18307 VOUT_P.n639 VOUT_P.t92 0.607167
R18308 VOUT_P.n639 VOUT_P.n638 0.607167
R18309 VOUT_P.n624 VOUT_P.t88 0.607167
R18310 VOUT_P.n624 VOUT_P.n623 0.607167
R18311 VOUT_P.n618 VOUT_P.t100 0.607167
R18312 VOUT_P.n618 VOUT_P.n617 0.607167
R18313 VOUT_P.n603 VOUT_P.t7 0.607167
R18314 VOUT_P.n603 VOUT_P.n602 0.607167
R18315 VOUT_P.n597 VOUT_P.t44 0.607167
R18316 VOUT_P.n597 VOUT_P.n596 0.607167
R18317 VOUT_P.n582 VOUT_P.t70 0.607167
R18318 VOUT_P.n582 VOUT_P.n581 0.607167
R18319 VOUT_P.n576 VOUT_P.t103 0.607167
R18320 VOUT_P.n576 VOUT_P.n575 0.607167
R18321 VOUT_P.n1280 VOUT_P.t43 0.607167
R18322 VOUT_P.n1280 VOUT_P.n1279 0.607167
R18323 VOUT_P.n1274 VOUT_P.t189 0.607167
R18324 VOUT_P.n1274 VOUT_P.n1273 0.607167
R18325 VOUT_P.n1268 VOUT_P.t126 0.607167
R18326 VOUT_P.n1268 VOUT_P.n1267 0.607167
R18327 VOUT_P.n1262 VOUT_P.t12 0.607167
R18328 VOUT_P.n1262 VOUT_P.n1261 0.607167
R18329 VOUT_P.n1256 VOUT_P.t82 0.607167
R18330 VOUT_P.n1256 VOUT_P.n1255 0.607167
R18331 VOUT_P.n1250 VOUT_P.t31 0.607167
R18332 VOUT_P.n1250 VOUT_P.n1249 0.607167
R18333 VOUT_P.n1244 VOUT_P.t118 0.607167
R18334 VOUT_P.n1244 VOUT_P.n1243 0.607167
R18335 VOUT_P.n1238 VOUT_P.t55 0.607167
R18336 VOUT_P.n1238 VOUT_P.n1237 0.607167
R18337 VOUT_P.n1232 VOUT_P.t125 0.607167
R18338 VOUT_P.n1232 VOUT_P.n1231 0.607167
R18339 VOUT_P.n1226 VOUT_P.t135 0.607167
R18340 VOUT_P.n1226 VOUT_P.n1225 0.607167
R18341 VOUT_P.n1220 VOUT_P.t72 0.607167
R18342 VOUT_P.n1220 VOUT_P.n1219 0.607167
R18343 VOUT_P.n1214 VOUT_P.t91 0.607167
R18344 VOUT_P.n1214 VOUT_P.n1213 0.607167
R18345 VOUT_P.n1208 VOUT_P.t23 0.607167
R18346 VOUT_P.n1208 VOUT_P.n1207 0.607167
R18347 VOUT_P.n1202 VOUT_P.t179 0.607167
R18348 VOUT_P.n1202 VOUT_P.n1201 0.607167
R18349 VOUT_P.n1196 VOUT_P.t61 0.607167
R18350 VOUT_P.n1196 VOUT_P.n1195 0.607167
R18351 VOUT_P.n1190 VOUT_P.t133 0.607167
R18352 VOUT_P.n1190 VOUT_P.n1189 0.607167
R18353 VOUT_P.n1184 VOUT_P.t71 0.607167
R18354 VOUT_P.n1184 VOUT_P.n1183 0.607167
R18355 VOUT_P.n1178 VOUT_P.t81 0.607167
R18356 VOUT_P.n1178 VOUT_P.n1177 0.607167
R18357 VOUT_P.n1172 VOUT_P.t150 0.607167
R18358 VOUT_P.n1172 VOUT_P.n1171 0.607167
R18359 VOUT_P.n1166 VOUT_P.t36 0.607167
R18360 VOUT_P.n1166 VOUT_P.n1165 0.607167
R18361 VOUT_P.n1160 VOUT_P.t175 0.607167
R18362 VOUT_P.n1160 VOUT_P.n1159 0.607167
R18363 VOUT_P.n1154 VOUT_P.t75 0.607167
R18364 VOUT_P.n1154 VOUT_P.n1153 0.607167
R18365 VOUT_P.n1148 VOUT_P.t93 0.607167
R18366 VOUT_P.n1148 VOUT_P.n1147 0.607167
R18367 VOUT_P.n1142 VOUT_P.t27 0.607167
R18368 VOUT_P.n1142 VOUT_P.n1141 0.607167
R18369 VOUT_P.n1136 VOUT_P.t164 0.607167
R18370 VOUT_P.n1136 VOUT_P.n1135 0.607167
R18371 VOUT_P.n192 VOUT_P.n191 0.572507
R18372 VOUT_P.n132 VOUT_P.n131 0.572507
R18373 VOUT_P.n36 VOUT_P.n35 0.572507
R18374 VOUT_P.n1602 VOUT_P.n1601 0.572507
R18375 VOUT_P.n1575 VOUT_P.n1574 0.572507
R18376 VOUT_P.n1515 VOUT_P.n1514 0.572507
R18377 VOUT_P.n349 VOUT_P.n348 0.555711
R18378 VOUT_P.n1364 VOUT_P.n1363 0.555711
R18379 VOUT_P.n1446 VOUT_P.n1445 0.552542
R18380 VOUT_P.n538 VOUT_P.n537 0.548033
R18381 VOUT_P.n1932 VOUT_P.t267 0.5465
R18382 VOUT_P.n1932 VOUT_P.n1931 0.5465
R18383 VOUT_P.n1937 VOUT_P.t237 0.5465
R18384 VOUT_P.n1937 VOUT_P.n1936 0.5465
R18385 VOUT_P.n1118 VOUT_P.t222 0.5465
R18386 VOUT_P.n1118 VOUT_P.n1117 0.5465
R18387 VOUT_P.n1112 VOUT_P.t208 0.5465
R18388 VOUT_P.n1112 VOUT_P.n1111 0.5465
R18389 VOUT_P.n1465 VOUT_P.t253 0.5465
R18390 VOUT_P.n1465 VOUT_P.n1464 0.5465
R18391 VOUT_P.n1480 VOUT_P.t268 0.5465
R18392 VOUT_P.n1480 VOUT_P.n1479 0.5465
R18393 VOUT_P.n1495 VOUT_P.t255 0.5465
R18394 VOUT_P.n1495 VOUT_P.n1494 0.5465
R18395 VOUT_P.n1553 VOUT_P.t216 0.5465
R18396 VOUT_P.n1553 VOUT_P.n1552 0.5465
R18397 VOUT_P.n1529 VOUT_P.t246 0.5465
R18398 VOUT_P.n1529 VOUT_P.n1528 0.5465
R18399 VOUT_P.n1523 VOUT_P.t270 0.5465
R18400 VOUT_P.n1523 VOUT_P.n1522 0.5465
R18401 VOUT_P.n1547 VOUT_P.t238 0.5465
R18402 VOUT_P.n1547 VOUT_P.n1546 0.5465
R18403 VOUT_P.n18 VOUT_P.t210 0.5465
R18404 VOUT_P.n18 VOUT_P.n17 0.5465
R18405 VOUT_P.n144 VOUT_P.t233 0.5465
R18406 VOUT_P.n144 VOUT_P.n143 0.5465
R18407 VOUT_P.n174 VOUT_P.t228 0.5465
R18408 VOUT_P.n174 VOUT_P.n173 0.5465
R18409 VOUT_P.n987 VOUT_P.t265 0.5465
R18410 VOUT_P.n987 VOUT_P.n986 0.5465
R18411 VOUT_P.n953 VOUT_P.t258 0.5465
R18412 VOUT_P.n953 VOUT_P.n952 0.5465
R18413 VOUT_P.n959 VOUT_P.t203 0.5465
R18414 VOUT_P.n959 VOUT_P.n958 0.5465
R18415 VOUT_P.n929 VOUT_P.t236 0.5465
R18416 VOUT_P.n929 VOUT_P.n928 0.5465
R18417 VOUT_P.n923 VOUT_P.t269 0.5465
R18418 VOUT_P.n923 VOUT_P.n922 0.5465
R18419 VOUT_P.n944 VOUT_P.t266 0.5465
R18420 VOUT_P.n944 VOUT_P.n943 0.5465
R18421 VOUT_P.n938 VOUT_P.t220 0.5465
R18422 VOUT_P.n938 VOUT_P.n937 0.5465
R18423 VOUT_P.n983 VOUT_P.t245 0.5465
R18424 VOUT_P.n983 VOUT_P.n982 0.5465
R18425 VOUT_P.n562 VOUT_P.t261 0.5465
R18426 VOUT_P.n562 VOUT_P.n561 0.5465
R18427 VOUT_P.n548 VOUT_P.t234 0.5465
R18428 VOUT_P.n548 VOUT_P.n547 0.5465
R18429 VOUT_P.n915 VOUT_P.t254 0.5465
R18430 VOUT_P.n915 VOUT_P.n914 0.5465
R18431 VOUT_P.n907 VOUT_P.t230 0.5465
R18432 VOUT_P.n907 VOUT_P.n906 0.5465
R18433 VOUT_P.n49 VOUT_P.t198 0.5465
R18434 VOUT_P.n49 VOUT_P.n48 0.5465
R18435 VOUT_P.n43 VOUT_P.t242 0.5465
R18436 VOUT_P.n43 VOUT_P.n42 0.5465
R18437 VOUT_P.n67 VOUT_P.t201 0.5465
R18438 VOUT_P.n67 VOUT_P.n66 0.5465
R18439 VOUT_P.n74 VOUT_P.t263 0.5465
R18440 VOUT_P.n74 VOUT_P.n73 0.5465
R18441 VOUT_P.n261 VOUT_P.n260 0.543352
R18442 VOUT_P.n1328 VOUT_P.n1327 0.543352
R18443 VOUT_P.n446 VOUT_P.n445 0.542718
R18444 VOUT_P.n1405 VOUT_P.n1404 0.542718
R18445 VOUT_P.n450 VOUT_P.n449 0.529408
R18446 VOUT_P.n1410 VOUT_P.n1409 0.529408
R18447 VOUT_P.n246 VOUT_P.n245 0.528775
R18448 VOUT_P.n1319 VOUT_P.n1318 0.528775
R18449 VOUT_P.n358 VOUT_P.n357 0.516415
R18450 VOUT_P.n1369 VOUT_P.n1368 0.516415
R18451 VOUT_P.n756 VOUT_P.n755 0.482824
R18452 VOUT_P.n812 VOUT_P.n811 0.482824
R18453 VOUT_P.n867 VOUT_P.n866 0.482824
R18454 VOUT_P.n1755 VOUT_P.n1754 0.482824
R18455 VOUT_P.n1795 VOUT_P.n1794 0.482824
R18456 VOUT_P.n1858 VOUT_P.n1857 0.482824
R18457 VOUT_P.n774 VOUT_P.n773 0.453986
R18458 VOUT_P.n1773 VOUT_P.n1772 0.453986
R18459 VOUT_P.n1025 VOUT_P.n1024 0.4505
R18460 VOUT_P.n1017 VOUT_P.n1016 0.4505
R18461 VOUT_P.n1071 VOUT_P.n1070 0.4505
R18462 VOUT_P.n1021 VOUT_P.n1020 0.4505
R18463 VOUT_P.n1899 VOUT_P.n1898 0.447157
R18464 VOUT_P.n885 VOUT_P.n884 0.446728
R18465 VOUT_P.n738 VOUT_P.n737 0.441627
R18466 VOUT_P.n1737 VOUT_P.n1736 0.441627
R18467 VOUT_P.n830 VOUT_P.n829 0.440993
R18468 VOUT_P.n1813 VOUT_P.n1812 0.440993
R18469 VOUT_P.n849 VOUT_P.n848 0.427683
R18470 VOUT_P.n1817 VOUT_P.n1816 0.427683
R18471 VOUT_P.n734 VOUT_P.n733 0.427049
R18472 VOUT_P.n1727 VOUT_P.n1726 0.427049
R18473 VOUT_P.n794 VOUT_P.n793 0.41469
R18474 VOUT_P.n1777 VOUT_P.n1776 0.41469
R18475 VOUT_P.n258 VOUT_P.n257 0.395359
R18476 VOUT_P.n725 VOUT_P.n724 0.389021
R18477 VOUT_P.n747 VOUT_P.n746 0.389021
R18478 VOUT_P.n765 VOUT_P.n764 0.389021
R18479 VOUT_P.n803 VOUT_P.n802 0.389021
R18480 VOUT_P.n821 VOUT_P.n820 0.389021
R18481 VOUT_P.n858 VOUT_P.n857 0.389021
R18482 VOUT_P.n876 VOUT_P.n875 0.389021
R18483 VOUT_P.n1718 VOUT_P.n1717 0.389021
R18484 VOUT_P.n1746 VOUT_P.n1745 0.389021
R18485 VOUT_P.n1764 VOUT_P.n1763 0.389021
R18486 VOUT_P.n1786 VOUT_P.n1785 0.389021
R18487 VOUT_P.n1804 VOUT_P.n1803 0.389021
R18488 VOUT_P.n1838 VOUT_P.n1837 0.389021
R18489 VOUT_P.n1879 VOUT_P.n1878 0.389021
R18490 VOUT_P.n129 VOUT_P.n87 0.356063
R18491 VOUT_P.n1924 VOUT_P.n1923 0.356063
R18492 VOUT_P.n1906 VOUT_P.n1905 0.356063
R18493 VOUT_P.n956 VOUT_P.n955 0.336464
R18494 VOUT_P.n993 VOUT_P.n992 0.336464
R18495 VOUT_P.n559 VOUT_P.n558 0.336464
R18496 VOUT_P.n842 VOUT_P.n841 0.2705
R18497 VOUT_P.n899 VOUT_P.n898 0.2705
R18498 VOUT_P.n788 VOUT_P.n787 0.2705
R18499 VOUT_P.n120 VOUT_P.n119 0.231204
R18500 VOUT_P.n1914 VOUT_P.n1910 0.231204
R18501 VOUT_P.n930 VOUT_P.n927 0.191654
R18502 VOUT_P.n945 VOUT_P.n942 0.191654
R18503 VOUT_P.n550 VOUT_P.n549 0.191654
R18504 VOUT_P.n1042 VOUT_P.n1041 0.187374
R18505 VOUT_P.n1946 VOUT_P.n1945 0.186204
R18506 VOUT_P.n1561 VOUT_P.n1560 0.186204
R18507 VOUT_P.n1537 VOUT_P.n1536 0.186204
R18508 VOUT_P.n95 VOUT_P.n94 0.186204
R18509 VOUT_P.n110 VOUT_P.n109 0.186204
R18510 VOUT_P.n556 VOUT_P.n555 0.186204
R18511 VOUT_P.n1005 VOUT_P.n1004 0.186204
R18512 VOUT_P.n980 VOUT_P.n979 0.186204
R18513 VOUT_P.n967 VOUT_P.n966 0.186204
R18514 VOUT_P.n720 VOUT_P.n719 0.186204
R18515 VOUT_P.n729 VOUT_P.n728 0.186204
R18516 VOUT_P.n742 VOUT_P.n741 0.186204
R18517 VOUT_P.n751 VOUT_P.n750 0.186204
R18518 VOUT_P.n760 VOUT_P.n759 0.186204
R18519 VOUT_P.n769 VOUT_P.n768 0.186204
R18520 VOUT_P.n798 VOUT_P.n797 0.186204
R18521 VOUT_P.n807 VOUT_P.n806 0.186204
R18522 VOUT_P.n816 VOUT_P.n815 0.186204
R18523 VOUT_P.n825 VOUT_P.n824 0.186204
R18524 VOUT_P.n853 VOUT_P.n852 0.186204
R18525 VOUT_P.n862 VOUT_P.n861 0.186204
R18526 VOUT_P.n871 VOUT_P.n870 0.186204
R18527 VOUT_P.n880 VOUT_P.n879 0.186204
R18528 VOUT_P.n213 VOUT_P.n212 0.186204
R18529 VOUT_P.n224 VOUT_P.n223 0.186204
R18530 VOUT_P.n235 VOUT_P.n234 0.186204
R18531 VOUT_P.n272 VOUT_P.n271 0.186204
R18532 VOUT_P.n283 VOUT_P.n282 0.186204
R18533 VOUT_P.n294 VOUT_P.n293 0.186204
R18534 VOUT_P.n316 VOUT_P.n315 0.186204
R18535 VOUT_P.n327 VOUT_P.n326 0.186204
R18536 VOUT_P.n338 VOUT_P.n337 0.186204
R18537 VOUT_P.n369 VOUT_P.n368 0.186204
R18538 VOUT_P.n380 VOUT_P.n379 0.186204
R18539 VOUT_P.n391 VOUT_P.n390 0.186204
R18540 VOUT_P.n413 VOUT_P.n412 0.186204
R18541 VOUT_P.n424 VOUT_P.n423 0.186204
R18542 VOUT_P.n435 VOUT_P.n434 0.186204
R18543 VOUT_P.n461 VOUT_P.n460 0.186204
R18544 VOUT_P.n472 VOUT_P.n471 0.186204
R18545 VOUT_P.n483 VOUT_P.n482 0.186204
R18546 VOUT_P.n505 VOUT_P.n504 0.186204
R18547 VOUT_P.n516 VOUT_P.n515 0.186204
R18548 VOUT_P.n527 VOUT_P.n526 0.186204
R18549 VOUT_P.n182 VOUT_P.n181 0.186204
R18550 VOUT_P.n171 VOUT_P.n170 0.186204
R18551 VOUT_P.n152 VOUT_P.n151 0.186204
R18552 VOUT_P.n141 VOUT_P.n140 0.186204
R18553 VOUT_P.n26 VOUT_P.n25 0.186204
R18554 VOUT_P.n15 VOUT_P.n14 0.186204
R18555 VOUT_P.n56 VOUT_P.n55 0.186204
R18556 VOUT_P.n81 VOUT_P.n80 0.186204
R18557 VOUT_P.n1597 VOUT_P.n1596 0.186204
R18558 VOUT_P.n1593 VOUT_P.n1592 0.186204
R18559 VOUT_P.n1584 VOUT_P.n1583 0.186204
R18560 VOUT_P.n1579 VOUT_P.n1578 0.186204
R18561 VOUT_P.n1510 VOUT_P.n1509 0.186204
R18562 VOUT_P.n1506 VOUT_P.n1505 0.186204
R18563 VOUT_P.n1714 VOUT_P.n1713 0.186204
R18564 VOUT_P.n1723 VOUT_P.n1722 0.186204
R18565 VOUT_P.n1742 VOUT_P.n1741 0.186204
R18566 VOUT_P.n1751 VOUT_P.n1750 0.186204
R18567 VOUT_P.n1760 VOUT_P.n1759 0.186204
R18568 VOUT_P.n1769 VOUT_P.n1768 0.186204
R18569 VOUT_P.n1782 VOUT_P.n1781 0.186204
R18570 VOUT_P.n1791 VOUT_P.n1790 0.186204
R18571 VOUT_P.n1800 VOUT_P.n1799 0.186204
R18572 VOUT_P.n1809 VOUT_P.n1808 0.186204
R18573 VOUT_P.n1827 VOUT_P.n1826 0.186204
R18574 VOUT_P.n1849 VOUT_P.n1848 0.186204
R18575 VOUT_P.n1868 VOUT_P.n1867 0.186204
R18576 VOUT_P.n1890 VOUT_P.n1889 0.186204
R18577 VOUT_P.n1306 VOUT_P.n1305 0.186204
R18578 VOUT_P.n1310 VOUT_P.n1309 0.186204
R18579 VOUT_P.n1315 VOUT_P.n1314 0.186204
R18580 VOUT_P.n1333 VOUT_P.n1332 0.186204
R18581 VOUT_P.n1337 VOUT_P.n1336 0.186204
R18582 VOUT_P.n1342 VOUT_P.n1341 0.186204
R18583 VOUT_P.n1351 VOUT_P.n1350 0.186204
R18584 VOUT_P.n1355 VOUT_P.n1354 0.186204
R18585 VOUT_P.n1360 VOUT_P.n1359 0.186204
R18586 VOUT_P.n1374 VOUT_P.n1373 0.186204
R18587 VOUT_P.n1378 VOUT_P.n1377 0.186204
R18588 VOUT_P.n1383 VOUT_P.n1382 0.186204
R18589 VOUT_P.n1392 VOUT_P.n1391 0.186204
R18590 VOUT_P.n1396 VOUT_P.n1395 0.186204
R18591 VOUT_P.n1401 VOUT_P.n1400 0.186204
R18592 VOUT_P.n1415 VOUT_P.n1414 0.186204
R18593 VOUT_P.n1419 VOUT_P.n1418 0.186204
R18594 VOUT_P.n1424 VOUT_P.n1423 0.186204
R18595 VOUT_P.n1433 VOUT_P.n1432 0.186204
R18596 VOUT_P.n1437 VOUT_P.n1436 0.186204
R18597 VOUT_P.n1442 VOUT_P.n1441 0.186204
R18598 VOUT_P.n1126 VOUT_P.n1125 0.186204
R18599 VOUT_P.n1072 VOUT_P.n1071 0.180553
R18600 VOUT_P.n1065 VOUT_P.n1040 0.180553
R18601 VOUT_P.n1096 VOUT_P.n1028 0.180553
R18602 VOUT_P.n837 VOUT_P.n836 0.145641
R18603 VOUT_P.n894 VOUT_P.n893 0.145641
R18604 VOUT_P.n783 VOUT_P.n782 0.145641
R18605 VOUT_P.n961 VOUT_P.n960 0.109963
R18606 VOUT_P.n927 VOUT_P.n926 0.106363
R18607 VOUT_P.n942 VOUT_P.n941 0.106363
R18608 VOUT_P.n551 VOUT_P.n550 0.106363
R18609 VOUT_P.n125 VOUT_P.n124 0.106345
R18610 VOUT_P.n1568 VOUT_P.n1567 0.106345
R18611 VOUT_P.n1919 VOUT_P.n1918 0.106345
R18612 VOUT_P.n1454 VOUT_P.n1453 0.106345
R18613 VOUT_P.n1451 VOUT_P.n1450 0.101908
R18614 VOUT_P.n1935 VOUT_P.n1930 0.0992756
R18615 VOUT_P.n1895 VOUT_P.n1892 0.0992756
R18616 VOUT_P.n1886 VOUT_P.n1881 0.0992756
R18617 VOUT_P.n1875 VOUT_P.n1870 0.0992756
R18618 VOUT_P.n1864 VOUT_P.n1860 0.0992756
R18619 VOUT_P.n1854 VOUT_P.n1851 0.0992756
R18620 VOUT_P.n1845 VOUT_P.n1840 0.0992756
R18621 VOUT_P.n1834 VOUT_P.n1829 0.0992756
R18622 VOUT_P.n1823 VOUT_P.n1819 0.0992756
R18623 VOUT_P.n220 VOUT_P.n215 0.0992756
R18624 VOUT_P.n231 VOUT_P.n226 0.0992756
R18625 VOUT_P.n242 VOUT_P.n237 0.0992756
R18626 VOUT_P.n268 VOUT_P.n263 0.0992756
R18627 VOUT_P.n279 VOUT_P.n274 0.0992756
R18628 VOUT_P.n290 VOUT_P.n285 0.0992756
R18629 VOUT_P.n301 VOUT_P.n296 0.0992756
R18630 VOUT_P.n312 VOUT_P.n307 0.0992756
R18631 VOUT_P.n323 VOUT_P.n318 0.0992756
R18632 VOUT_P.n334 VOUT_P.n329 0.0992756
R18633 VOUT_P.n345 VOUT_P.n340 0.0992756
R18634 VOUT_P.n365 VOUT_P.n360 0.0992756
R18635 VOUT_P.n376 VOUT_P.n371 0.0992756
R18636 VOUT_P.n387 VOUT_P.n382 0.0992756
R18637 VOUT_P.n398 VOUT_P.n393 0.0992756
R18638 VOUT_P.n409 VOUT_P.n404 0.0992756
R18639 VOUT_P.n420 VOUT_P.n415 0.0992756
R18640 VOUT_P.n431 VOUT_P.n426 0.0992756
R18641 VOUT_P.n442 VOUT_P.n437 0.0992756
R18642 VOUT_P.n457 VOUT_P.n452 0.0992756
R18643 VOUT_P.n468 VOUT_P.n463 0.0992756
R18644 VOUT_P.n479 VOUT_P.n474 0.0992756
R18645 VOUT_P.n490 VOUT_P.n485 0.0992756
R18646 VOUT_P.n501 VOUT_P.n496 0.0992756
R18647 VOUT_P.n512 VOUT_P.n507 0.0992756
R18648 VOUT_P.n523 VOUT_P.n518 0.0992756
R18649 VOUT_P.n534 VOUT_P.n529 0.0992756
R18650 VOUT_P.n565 VOUT_P.n560 0.0992756
R18651 VOUT_P.n1903 VOUT_P.n1902 0.0982485
R18652 VOUT_P.n905 VOUT_P.n904 0.0978197
R18653 VOUT_P.n542 VOUT_P.n541 0.0973992
R18654 VOUT_P.n1093 VOUT_P.n1092 0.0890366
R18655 VOUT_P.n1062 VOUT_P.n1061 0.0890366
R18656 VOUT_P.n1502 VOUT_P.n1501 0.0832399
R18657 VOUT_P.n106 VOUT_P.n105 0.0832399
R18658 VOUT_P.n552 VOUT_P.n546 0.0832399
R18659 VOUT_P.n76 VOUT_P.n72 0.0832399
R18660 VOUT_P.n209 VOUT_P.n208 0.0831446
R18661 VOUT_P.n11 VOUT_P.n10 0.0826464
R18662 VOUT_P.n22 VOUT_P.n21 0.0826464
R18663 VOUT_P.n32 VOUT_P.n31 0.0826464
R18664 VOUT_P.n137 VOUT_P.n136 0.0826464
R18665 VOUT_P.n148 VOUT_P.n147 0.0826464
R18666 VOUT_P.n158 VOUT_P.n157 0.0826464
R18667 VOUT_P.n167 VOUT_P.n166 0.0826464
R18668 VOUT_P.n178 VOUT_P.n177 0.0826464
R18669 VOUT_P.n188 VOUT_P.n187 0.0826464
R18670 VOUT_P.n103 VOUT_P.n101 0.0824117
R18671 VOUT_P.n913 VOUT_P.n909 0.0824117
R18672 VOUT_P.n1301 VOUT_P.n1296 0.0823987
R18673 VOUT_P.n1289 VOUT_P.n1284 0.0823987
R18674 VOUT_P.n1115 VOUT_P.n1110 0.0823987
R18675 VOUT_P.n1709 VOUT_P.n1705 0.0823987
R18676 VOUT_P.n1698 VOUT_P.n1693 0.0823987
R18677 VOUT_P.n1688 VOUT_P.n1684 0.0823987
R18678 VOUT_P.n1677 VOUT_P.n1672 0.0823987
R18679 VOUT_P.n1667 VOUT_P.n1663 0.0823987
R18680 VOUT_P.n1656 VOUT_P.n1651 0.0823987
R18681 VOUT_P.n1646 VOUT_P.n1642 0.0823987
R18682 VOUT_P.n1635 VOUT_P.n1630 0.0823987
R18683 VOUT_P.n1625 VOUT_P.n1621 0.0823987
R18684 VOUT_P.n1614 VOUT_P.n1609 0.0823987
R18685 VOUT_P.n1462 VOUT_P.n1458 0.0823987
R18686 VOUT_P.n1472 VOUT_P.n1469 0.0823987
R18687 VOUT_P.n1483 VOUT_P.n1478 0.0823987
R18688 VOUT_P.n1492 VOUT_P.n1488 0.0823987
R18689 VOUT_P.n1556 VOUT_P.n1551 0.0823987
R18690 VOUT_P.n1526 VOUT_P.n1521 0.0823987
R18691 VOUT_P.n711 VOUT_P.n706 0.0823987
R18692 VOUT_P.n699 VOUT_P.n696 0.0823987
R18693 VOUT_P.n690 VOUT_P.n685 0.0823987
R18694 VOUT_P.n678 VOUT_P.n675 0.0823987
R18695 VOUT_P.n669 VOUT_P.n664 0.0823987
R18696 VOUT_P.n657 VOUT_P.n654 0.0823987
R18697 VOUT_P.n648 VOUT_P.n643 0.0823987
R18698 VOUT_P.n636 VOUT_P.n633 0.0823987
R18699 VOUT_P.n627 VOUT_P.n622 0.0823987
R18700 VOUT_P.n615 VOUT_P.n612 0.0823987
R18701 VOUT_P.n606 VOUT_P.n601 0.0823987
R18702 VOUT_P.n594 VOUT_P.n591 0.0823987
R18703 VOUT_P.n585 VOUT_P.n580 0.0823987
R18704 VOUT_P.n573 VOUT_P.n570 0.0823987
R18705 VOUT_P.n991 VOUT_P.n990 0.0823987
R18706 VOUT_P.n934 VOUT_P.n925 0.0823987
R18707 VOUT_P.n949 VOUT_P.n940 0.0823987
R18708 VOUT_P.n921 VOUT_P.n917 0.0823987
R18709 VOUT_P.n46 VOUT_P.n41 0.0823987
R18710 VOUT_P.n1277 VOUT_P.n1272 0.0823987
R18711 VOUT_P.n1265 VOUT_P.n1260 0.0823987
R18712 VOUT_P.n1253 VOUT_P.n1248 0.0823987
R18713 VOUT_P.n1241 VOUT_P.n1236 0.0823987
R18714 VOUT_P.n1229 VOUT_P.n1224 0.0823987
R18715 VOUT_P.n1217 VOUT_P.n1212 0.0823987
R18716 VOUT_P.n1205 VOUT_P.n1200 0.0823987
R18717 VOUT_P.n1193 VOUT_P.n1188 0.0823987
R18718 VOUT_P.n1181 VOUT_P.n1176 0.0823987
R18719 VOUT_P.n1169 VOUT_P.n1164 0.0823987
R18720 VOUT_P.n1157 VOUT_P.n1152 0.0823987
R18721 VOUT_P.n1145 VOUT_P.n1140 0.0823987
R18722 VOUT_P.n955 VOUT_P.n954 0.0748144
R18723 VOUT_P.n992 VOUT_P.n989 0.0748144
R18724 VOUT_P.n1550 VOUT_P.n1545 0.0712285
R18725 VOUT_P.n1532 VOUT_P.n1527 0.0712285
R18726 VOUT_P.n90 VOUT_P.n88 0.0712285
R18727 VOUT_P.n579 VOUT_P.n574 0.0712285
R18728 VOUT_P.n590 VOUT_P.n586 0.0712285
R18729 VOUT_P.n600 VOUT_P.n595 0.0712285
R18730 VOUT_P.n611 VOUT_P.n607 0.0712285
R18731 VOUT_P.n621 VOUT_P.n616 0.0712285
R18732 VOUT_P.n632 VOUT_P.n628 0.0712285
R18733 VOUT_P.n642 VOUT_P.n637 0.0712285
R18734 VOUT_P.n653 VOUT_P.n649 0.0712285
R18735 VOUT_P.n663 VOUT_P.n658 0.0712285
R18736 VOUT_P.n674 VOUT_P.n670 0.0712285
R18737 VOUT_P.n684 VOUT_P.n679 0.0712285
R18738 VOUT_P.n695 VOUT_P.n691 0.0712285
R18739 VOUT_P.n705 VOUT_P.n700 0.0712285
R18740 VOUT_P.n716 VOUT_P.n712 0.0712285
R18741 VOUT_P.n70 VOUT_P.n65 0.0712285
R18742 VOUT_P.n52 VOUT_P.n47 0.0712285
R18743 VOUT_P.n1487 VOUT_P.n1484 0.0712285
R18744 VOUT_P.n1498 VOUT_P.n1493 0.0712285
R18745 VOUT_P.n1477 VOUT_P.n1473 0.0712285
R18746 VOUT_P.n1468 VOUT_P.n1463 0.0712285
R18747 VOUT_P.n1608 VOUT_P.n1605 0.0712285
R18748 VOUT_P.n1620 VOUT_P.n1615 0.0712285
R18749 VOUT_P.n1629 VOUT_P.n1626 0.0712285
R18750 VOUT_P.n1641 VOUT_P.n1636 0.0712285
R18751 VOUT_P.n1650 VOUT_P.n1647 0.0712285
R18752 VOUT_P.n1662 VOUT_P.n1657 0.0712285
R18753 VOUT_P.n1671 VOUT_P.n1668 0.0712285
R18754 VOUT_P.n1683 VOUT_P.n1678 0.0712285
R18755 VOUT_P.n1692 VOUT_P.n1689 0.0712285
R18756 VOUT_P.n1704 VOUT_P.n1699 0.0712285
R18757 VOUT_P.n1139 VOUT_P.n1134 0.0712285
R18758 VOUT_P.n1151 VOUT_P.n1146 0.0712285
R18759 VOUT_P.n1163 VOUT_P.n1158 0.0712285
R18760 VOUT_P.n1175 VOUT_P.n1170 0.0712285
R18761 VOUT_P.n1187 VOUT_P.n1182 0.0712285
R18762 VOUT_P.n1199 VOUT_P.n1194 0.0712285
R18763 VOUT_P.n1211 VOUT_P.n1206 0.0712285
R18764 VOUT_P.n1223 VOUT_P.n1218 0.0712285
R18765 VOUT_P.n1235 VOUT_P.n1230 0.0712285
R18766 VOUT_P.n1247 VOUT_P.n1242 0.0712285
R18767 VOUT_P.n1259 VOUT_P.n1254 0.0712285
R18768 VOUT_P.n1271 VOUT_P.n1266 0.0712285
R18769 VOUT_P.n1283 VOUT_P.n1278 0.0712285
R18770 VOUT_P.n1121 VOUT_P.n1116 0.0712285
R18771 VOUT_P.n1295 VOUT_P.n1290 0.0712285
R18772 VOUT_P.n997 VOUT_P.n996 0.0709833
R18773 VOUT_P VOUT_P.n1989 0.0664984
R18774 VOUT_P.n1941 VOUT_P.n1940 0.0623855
R18775 VOUT_P.n1940 VOUT_P.n1939 0.0623855
R18776 VOUT_P.n962 VOUT_P.n951 0.0623855
R18777 VOUT_P.n951 VOUT_P.n950 0.0623855
R18778 VOUT_P.n997 VOUT_P.n985 0.0536862
R18779 VOUT_P.n1532 VOUT_P.n1531 0.0534597
R18780 VOUT_P.n1550 VOUT_P.n1549 0.0534597
R18781 VOUT_P.n90 VOUT_P.n89 0.0534597
R18782 VOUT_P.n716 VOUT_P.n715 0.0534597
R18783 VOUT_P.n705 VOUT_P.n704 0.0534597
R18784 VOUT_P.n695 VOUT_P.n694 0.0534597
R18785 VOUT_P.n684 VOUT_P.n683 0.0534597
R18786 VOUT_P.n674 VOUT_P.n673 0.0534597
R18787 VOUT_P.n663 VOUT_P.n662 0.0534597
R18788 VOUT_P.n653 VOUT_P.n652 0.0534597
R18789 VOUT_P.n642 VOUT_P.n641 0.0534597
R18790 VOUT_P.n632 VOUT_P.n631 0.0534597
R18791 VOUT_P.n621 VOUT_P.n620 0.0534597
R18792 VOUT_P.n611 VOUT_P.n610 0.0534597
R18793 VOUT_P.n600 VOUT_P.n599 0.0534597
R18794 VOUT_P.n590 VOUT_P.n589 0.0534597
R18795 VOUT_P.n579 VOUT_P.n578 0.0534597
R18796 VOUT_P.n52 VOUT_P.n51 0.0534597
R18797 VOUT_P.n70 VOUT_P.n69 0.0534597
R18798 VOUT_P.n1498 VOUT_P.n1497 0.0534597
R18799 VOUT_P.n1468 VOUT_P.n1467 0.0534597
R18800 VOUT_P.n1477 VOUT_P.n1476 0.0534597
R18801 VOUT_P.n1487 VOUT_P.n1486 0.0534597
R18802 VOUT_P.n1704 VOUT_P.n1703 0.0534597
R18803 VOUT_P.n1692 VOUT_P.n1691 0.0534597
R18804 VOUT_P.n1683 VOUT_P.n1682 0.0534597
R18805 VOUT_P.n1671 VOUT_P.n1670 0.0534597
R18806 VOUT_P.n1662 VOUT_P.n1661 0.0534597
R18807 VOUT_P.n1650 VOUT_P.n1649 0.0534597
R18808 VOUT_P.n1641 VOUT_P.n1640 0.0534597
R18809 VOUT_P.n1629 VOUT_P.n1628 0.0534597
R18810 VOUT_P.n1620 VOUT_P.n1619 0.0534597
R18811 VOUT_P.n1608 VOUT_P.n1607 0.0534597
R18812 VOUT_P.n1121 VOUT_P.n1120 0.0534597
R18813 VOUT_P.n1295 VOUT_P.n1294 0.0534597
R18814 VOUT_P.n1283 VOUT_P.n1282 0.0534597
R18815 VOUT_P.n1271 VOUT_P.n1270 0.0534597
R18816 VOUT_P.n1259 VOUT_P.n1258 0.0534597
R18817 VOUT_P.n1247 VOUT_P.n1246 0.0534597
R18818 VOUT_P.n1235 VOUT_P.n1234 0.0534597
R18819 VOUT_P.n1223 VOUT_P.n1222 0.0534597
R18820 VOUT_P.n1211 VOUT_P.n1210 0.0534597
R18821 VOUT_P.n1199 VOUT_P.n1198 0.0534597
R18822 VOUT_P.n1187 VOUT_P.n1186 0.0534597
R18823 VOUT_P.n1175 VOUT_P.n1174 0.0534597
R18824 VOUT_P.n1163 VOUT_P.n1162 0.0534597
R18825 VOUT_P.n1151 VOUT_P.n1150 0.0534597
R18826 VOUT_P.n1139 VOUT_P.n1138 0.0534597
R18827 VOUT_P.n11 VOUT_P.n9 0.0423164
R18828 VOUT_P.n22 VOUT_P.n20 0.0423164
R18829 VOUT_P.n32 VOUT_P.n30 0.0423164
R18830 VOUT_P.n137 VOUT_P.n135 0.0423164
R18831 VOUT_P.n148 VOUT_P.n146 0.0423164
R18832 VOUT_P.n158 VOUT_P.n156 0.0423164
R18833 VOUT_P.n167 VOUT_P.n165 0.0423164
R18834 VOUT_P.n178 VOUT_P.n176 0.0423164
R18835 VOUT_P.n188 VOUT_P.n186 0.0423164
R18836 VOUT_P.n208 VOUT_P.n207 0.0420655
R18837 VOUT_P.n1501 VOUT_P.n1500 0.0419676
R18838 VOUT_P.n105 VOUT_P.n104 0.0419676
R18839 VOUT_P.n546 VOUT_P.n545 0.0419676
R18840 VOUT_P.n72 VOUT_P.n71 0.0419676
R18841 VOUT_P.n1526 VOUT_P.n1525 0.0415773
R18842 VOUT_P.n1556 VOUT_P.n1555 0.0415773
R18843 VOUT_P.n949 VOUT_P.n948 0.0415773
R18844 VOUT_P.n934 VOUT_P.n933 0.0415773
R18845 VOUT_P.n921 VOUT_P.n920 0.0415773
R18846 VOUT_P.n573 VOUT_P.n572 0.0415773
R18847 VOUT_P.n585 VOUT_P.n584 0.0415773
R18848 VOUT_P.n594 VOUT_P.n593 0.0415773
R18849 VOUT_P.n606 VOUT_P.n605 0.0415773
R18850 VOUT_P.n615 VOUT_P.n614 0.0415773
R18851 VOUT_P.n627 VOUT_P.n626 0.0415773
R18852 VOUT_P.n636 VOUT_P.n635 0.0415773
R18853 VOUT_P.n648 VOUT_P.n647 0.0415773
R18854 VOUT_P.n657 VOUT_P.n656 0.0415773
R18855 VOUT_P.n669 VOUT_P.n668 0.0415773
R18856 VOUT_P.n678 VOUT_P.n677 0.0415773
R18857 VOUT_P.n690 VOUT_P.n689 0.0415773
R18858 VOUT_P.n699 VOUT_P.n698 0.0415773
R18859 VOUT_P.n711 VOUT_P.n710 0.0415773
R18860 VOUT_P.n46 VOUT_P.n45 0.0415773
R18861 VOUT_P.n1492 VOUT_P.n1491 0.0415773
R18862 VOUT_P.n1483 VOUT_P.n1482 0.0415773
R18863 VOUT_P.n1472 VOUT_P.n1471 0.0415773
R18864 VOUT_P.n1462 VOUT_P.n1461 0.0415773
R18865 VOUT_P.n1614 VOUT_P.n1613 0.0415773
R18866 VOUT_P.n1625 VOUT_P.n1624 0.0415773
R18867 VOUT_P.n1635 VOUT_P.n1634 0.0415773
R18868 VOUT_P.n1646 VOUT_P.n1645 0.0415773
R18869 VOUT_P.n1656 VOUT_P.n1655 0.0415773
R18870 VOUT_P.n1667 VOUT_P.n1666 0.0415773
R18871 VOUT_P.n1677 VOUT_P.n1676 0.0415773
R18872 VOUT_P.n1688 VOUT_P.n1687 0.0415773
R18873 VOUT_P.n1698 VOUT_P.n1697 0.0415773
R18874 VOUT_P.n1709 VOUT_P.n1708 0.0415773
R18875 VOUT_P.n1145 VOUT_P.n1144 0.0415773
R18876 VOUT_P.n1157 VOUT_P.n1156 0.0415773
R18877 VOUT_P.n1169 VOUT_P.n1168 0.0415773
R18878 VOUT_P.n1181 VOUT_P.n1180 0.0415773
R18879 VOUT_P.n1193 VOUT_P.n1192 0.0415773
R18880 VOUT_P.n1205 VOUT_P.n1204 0.0415773
R18881 VOUT_P.n1217 VOUT_P.n1216 0.0415773
R18882 VOUT_P.n1229 VOUT_P.n1228 0.0415773
R18883 VOUT_P.n1241 VOUT_P.n1240 0.0415773
R18884 VOUT_P.n1253 VOUT_P.n1252 0.0415773
R18885 VOUT_P.n1265 VOUT_P.n1264 0.0415773
R18886 VOUT_P.n1277 VOUT_P.n1276 0.0415773
R18887 VOUT_P.n1115 VOUT_P.n1114 0.0415773
R18888 VOUT_P.n1289 VOUT_P.n1288 0.0415773
R18889 VOUT_P.n1301 VOUT_P.n1300 0.0415773
R18890 VOUT_P.n103 VOUT_P.n102 0.0415636
R18891 VOUT_P.n913 VOUT_P.n912 0.0415636
R18892 VOUT_P.n116 VOUT_P.n115 0.0334577
R18893 VOUT_P.n1012 VOUT_P.n905 0.0334577
R18894 VOUT_P.n974 VOUT_P.n973 0.0334577
R18895 VOUT_P.n973 VOUT_P.n972 0.0334577
R18896 VOUT_P.n737 VOUT_P.n736 0.0334577
R18897 VOUT_P.n844 VOUT_P.n830 0.0334577
R18898 VOUT_P.n449 VOUT_P.n448 0.0334577
R18899 VOUT_P.n193 VOUT_P.n192 0.0334577
R18900 VOUT_P.n1776 VOUT_P.n1775 0.0334577
R18901 VOUT_P.n1816 VOUT_P.n1815 0.0334577
R18902 VOUT_P.n1092 VOUT_P.t225 0.0306947
R18903 VOUT_P.n1061 VOUT_P.t226 0.0285465
R18904 VOUT_P.n1935 VOUT_P.n1934 0.0254881
R18905 VOUT_P.n565 VOUT_P.n564 0.0254881
R18906 VOUT_P.n534 VOUT_P.n533 0.0254881
R18907 VOUT_P.n523 VOUT_P.n522 0.0254881
R18908 VOUT_P.n512 VOUT_P.n511 0.0254881
R18909 VOUT_P.n501 VOUT_P.n500 0.0254881
R18910 VOUT_P.n490 VOUT_P.n489 0.0254881
R18911 VOUT_P.n479 VOUT_P.n478 0.0254881
R18912 VOUT_P.n468 VOUT_P.n467 0.0254881
R18913 VOUT_P.n457 VOUT_P.n456 0.0254881
R18914 VOUT_P.n442 VOUT_P.n441 0.0254881
R18915 VOUT_P.n431 VOUT_P.n430 0.0254881
R18916 VOUT_P.n420 VOUT_P.n419 0.0254881
R18917 VOUT_P.n409 VOUT_P.n408 0.0254881
R18918 VOUT_P.n398 VOUT_P.n397 0.0254881
R18919 VOUT_P.n387 VOUT_P.n386 0.0254881
R18920 VOUT_P.n376 VOUT_P.n375 0.0254881
R18921 VOUT_P.n365 VOUT_P.n364 0.0254881
R18922 VOUT_P.n345 VOUT_P.n344 0.0254881
R18923 VOUT_P.n334 VOUT_P.n333 0.0254881
R18924 VOUT_P.n323 VOUT_P.n322 0.0254881
R18925 VOUT_P.n312 VOUT_P.n311 0.0254881
R18926 VOUT_P.n301 VOUT_P.n300 0.0254881
R18927 VOUT_P.n290 VOUT_P.n289 0.0254881
R18928 VOUT_P.n279 VOUT_P.n278 0.0254881
R18929 VOUT_P.n268 VOUT_P.n267 0.0254881
R18930 VOUT_P.n242 VOUT_P.n241 0.0254881
R18931 VOUT_P.n231 VOUT_P.n230 0.0254881
R18932 VOUT_P.n220 VOUT_P.n219 0.0254881
R18933 VOUT_P.n1823 VOUT_P.n1822 0.0254881
R18934 VOUT_P.n1834 VOUT_P.n1833 0.0254881
R18935 VOUT_P.n1845 VOUT_P.n1844 0.0254881
R18936 VOUT_P.n1854 VOUT_P.n1853 0.0254881
R18937 VOUT_P.n1864 VOUT_P.n1863 0.0254881
R18938 VOUT_P.n1875 VOUT_P.n1874 0.0254881
R18939 VOUT_P.n1886 VOUT_P.n1885 0.0254881
R18940 VOUT_P.n1895 VOUT_P.n1894 0.0254881
R18941 VOUT_P.n789 VOUT_P.n788 0.0235313
R18942 VOUT_P.n351 VOUT_P.n350 0.0235313
R18943 VOUT_P.n126 VOUT_P.n125 0.0235313
R18944 VOUT_P.n249 VOUT_P.n248 0.0235313
R18945 VOUT_P.n1367 VOUT_P.n1366 0.0235313
R18946 VOUT_P.n1408 VOUT_P.n1407 0.0235313
R18947 VOUT_P.n1449 VOUT_P.n1448 0.0235313
R18948 VOUT_P.n1900 VOUT_P.n1899 0.0234412
R18949 VOUT_P.n901 VOUT_P.n900 0.0228651
R18950 VOUT_P.n777 VOUT_P.n776 0.0228651
R18951 VOUT_P.n448 VOUT_P.n447 0.0228651
R18952 VOUT_P.n353 VOUT_P.n352 0.0228651
R18953 VOUT_P.n201 VOUT_P.n199 0.0228651
R18954 VOUT_P.n196 VOUT_P.n194 0.0228651
R18955 VOUT_P.n38 VOUT_P.n37 0.0228651
R18956 VOUT_P.n118 VOUT_P.n117 0.0228651
R18957 VOUT_P.n1517 VOUT_P.n1516 0.0228651
R18958 VOUT_P.n1569 VOUT_P.n1568 0.0228651
R18959 VOUT_P.n838 VOUT_P.n837 0.0228651
R18960 VOUT_P.n1814 VOUT_P.n1813 0.0228651
R18961 VOUT_P.n1729 VOUT_P.n1728 0.0228651
R18962 VOUT_P.n736 VOUT_P.n735 0.0228651
R18963 VOUT_P.n251 VOUT_P.n250 0.0228651
R18964 VOUT_P.n255 VOUT_P.n254 0.0228651
R18965 VOUT_P.n1731 VOUT_P.n1730 0.0228651
R18966 VOUT_P.n779 VOUT_P.n778 0.0228651
R18967 VOUT_P.n833 VOUT_P.n832 0.0228651
R18968 VOUT_P.n890 VOUT_P.n889 0.0228651
R18969 VOUT_P.n1918 VOUT_P.n1917 0.0228651
R18970 VOUT_P.n1921 VOUT_P.n1920 0.0228651
R18971 VOUT_P.n543 VOUT_P.n193 0.0228651
R18972 VOUT_P.n1925 VOUT_P.n1924 0.0228651
R18973 VOUT_P.n1100 VOUT_P.n1099 0.0228651
R18974 VOUT_P.n1455 VOUT_P.n1454 0.0228651
R18975 VOUT_P.n541 VOUT_P.n540 0.0211167
R18976 VOUT_P.n1067 VOUT_P.n1066 0.0195244
R18977 VOUT_P.n1068 VOUT_P.n1067 0.0195244
R18978 VOUT_P.n1069 VOUT_P.n1068 0.0195244
R18979 VOUT_P.n903 VOUT_P.n899 0.0179841
R18980 VOUT_P.n843 VOUT_P.n831 0.0179841
R18981 VOUT_P.n847 VOUT_P.n844 0.0179841
R18982 VOUT_P.n775 VOUT_P.n774 0.0179841
R18983 VOUT_P.n124 VOUT_P.n123 0.0179841
R18984 VOUT_P.n122 VOUT_P.n121 0.0179841
R18985 VOUT_P.n100 VOUT_P.n99 0.0179841
R18986 VOUT_P.n1542 VOUT_P.n1520 0.0179841
R18987 VOUT_P.n1519 VOUT_P.n1518 0.0179841
R18988 VOUT_P.n1572 VOUT_P.n1571 0.0179841
R18989 VOUT_P.n896 VOUT_P.n895 0.0179841
R18990 VOUT_P.n898 VOUT_P.n897 0.0179841
R18991 VOUT_P.n787 VOUT_P.n786 0.0179841
R18992 VOUT_P.n785 VOUT_P.n784 0.0179841
R18993 VOUT_P.n841 VOUT_P.n840 0.0179841
R18994 VOUT_P.n1774 VOUT_P.n1773 0.0179841
R18995 VOUT_P.n259 VOUT_P.n252 0.0179841
R18996 VOUT_P.n1323 VOUT_P.n1322 0.0179841
R18997 VOUT_P.n892 VOUT_P.n891 0.0179841
R18998 VOUT_P.n835 VOUT_P.n834 0.0179841
R18999 VOUT_P.n782 VOUT_P.n781 0.0179841
R19000 VOUT_P.n1320 VOUT_P.n1319 0.0179841
R19001 VOUT_P.n1326 VOUT_P.n1325 0.0179841
R19002 VOUT_P.n1131 VOUT_P.n1109 0.0179841
R19003 VOUT_P.n1908 VOUT_P.n1907 0.0179841
R19004 VOUT_P.n1910 VOUT_P.n1909 0.0179841
R19005 VOUT_P.n1916 VOUT_P.n1915 0.0179841
R19006 VOUT_P.n1012 VOUT_P.n1011 0.0179841
R19007 VOUT_P.n1952 VOUT_P.n1929 0.0179841
R19008 VOUT_P.n1603 VOUT_P.n1456 0.0179841
R19009 VOUT_P.n1108 VOUT_P.n1107 0.0179841
R19010 VOUT_P.n1098 VOUT_P.n1013 0.0179841
R19011 VOUT_P.n843 VOUT_P.n842 0.0177304
R19012 VOUT_P.n903 VOUT_P.n902 0.0177304
R19013 VOUT_P.n846 VOUT_P.n845 0.0177304
R19014 VOUT_P.n848 VOUT_P.n847 0.0177304
R19015 VOUT_P.n781 VOUT_P.n780 0.0177304
R19016 VOUT_P.n776 VOUT_P.n775 0.0177304
R19017 VOUT_P.n355 VOUT_P.n354 0.0177304
R19018 VOUT_P.n64 VOUT_P.n63 0.0177304
R19019 VOUT_P.n116 VOUT_P.n100 0.0177304
R19020 VOUT_P.n123 VOUT_P.n122 0.0177304
R19021 VOUT_P.n121 VOUT_P.n120 0.0177304
R19022 VOUT_P.n40 VOUT_P.n39 0.0177304
R19023 VOUT_P.n1571 VOUT_P.n1570 0.0177304
R19024 VOUT_P.n897 VOUT_P.n896 0.0177304
R19025 VOUT_P.n895 VOUT_P.n894 0.0177304
R19026 VOUT_P.n1775 VOUT_P.n1774 0.0177304
R19027 VOUT_P.n840 VOUT_P.n839 0.0177304
R19028 VOUT_P.n786 VOUT_P.n785 0.0177304
R19029 VOUT_P.n784 VOUT_P.n783 0.0177304
R19030 VOUT_P.n259 VOUT_P.n258 0.0177304
R19031 VOUT_P.n893 VOUT_P.n892 0.0177304
R19032 VOUT_P.n836 VOUT_P.n835 0.0177304
R19033 VOUT_P.n1321 VOUT_P.n1320 0.0177304
R19034 VOUT_P.n1011 VOUT_P.n1010 0.0177304
R19035 VOUT_P.n1915 VOUT_P.n1914 0.0177304
R19036 VOUT_P.n1909 VOUT_P.n1908 0.0177304
R19037 VOUT_P.n1907 VOUT_P.n1906 0.0177304
R19038 VOUT_P.n1952 VOUT_P.n1951 0.0177304
R19039 VOUT_P.n1905 VOUT_P.n1603 0.0177304
R19040 VOUT_P.n1107 VOUT_P.n1106 0.0177304
R19041 VOUT_P.n1098 VOUT_P.n1097 0.0177304
R19042 VOUT_P.n203 VOUT_P.n202 0.0174187
R19043 VOUT_P.n198 VOUT_P.n197 0.0174187
R19044 VOUT_P.n256 VOUT_P.n255 0.0174187
R19045 VOUT_P.n257 VOUT_P.n256 0.0174187
R19046 VOUT_P.n1922 VOUT_P.n1921 0.0174187
R19047 VOUT_P.n1923 VOUT_P.n1922 0.0174187
R19048 VOUT_P.n1566 VOUT_P.n1544 0.0173591
R19049 VOUT_P.n1913 VOUT_P.n1911 0.0173591
R19050 VOUT_P.n792 VOUT_P.n790 0.0173591
R19051 VOUT_P.n792 VOUT_P.n791 0.0173591
R19052 VOUT_P.n248 VOUT_P.n247 0.0173591
R19053 VOUT_P.n357 VOUT_P.n356 0.0173591
R19054 VOUT_P.n356 VOUT_P.n351 0.0173591
R19055 VOUT_P.n130 VOUT_P.n38 0.0173591
R19056 VOUT_P.n86 VOUT_P.n64 0.0173591
R19057 VOUT_P.n62 VOUT_P.n40 0.0173591
R19058 VOUT_P.n128 VOUT_P.n127 0.0173591
R19059 VOUT_P.n1543 VOUT_P.n1519 0.0173591
R19060 VOUT_P.n86 VOUT_P.n85 0.0173591
R19061 VOUT_P.n129 VOUT_P.n128 0.0173591
R19062 VOUT_P.n131 VOUT_P.n130 0.0173591
R19063 VOUT_P.n1567 VOUT_P.n1543 0.0173591
R19064 VOUT_P.n1566 VOUT_P.n1565 0.0173591
R19065 VOUT_P.n87 VOUT_P.n62 0.0173591
R19066 VOUT_P.n1904 VOUT_P.n1604 0.0173591
R19067 VOUT_P.n1574 VOUT_P.n1573 0.0173591
R19068 VOUT_P.n1573 VOUT_P.n1517 0.0173591
R19069 VOUT_P.n1735 VOUT_P.n1729 0.0173591
R19070 VOUT_P.n1734 VOUT_P.n1733 0.0173591
R19071 VOUT_P.n1733 VOUT_P.n1732 0.0173591
R19072 VOUT_P.n1736 VOUT_P.n1735 0.0173591
R19073 VOUT_P.n247 VOUT_P.n246 0.0173591
R19074 VOUT_P.n1327 VOUT_P.n1324 0.0173591
R19075 VOUT_P.n1366 VOUT_P.n1365 0.0173591
R19076 VOUT_P.n1407 VOUT_P.n1406 0.0173591
R19077 VOUT_P.n1448 VOUT_P.n1447 0.0173591
R19078 VOUT_P.n1452 VOUT_P.n1133 0.0173591
R19079 VOUT_P.n1324 VOUT_P.n1321 0.0173591
R19080 VOUT_P.n1447 VOUT_P.n1446 0.0173591
R19081 VOUT_P.n1406 VOUT_P.n1405 0.0173591
R19082 VOUT_P.n1365 VOUT_P.n1364 0.0173591
R19083 VOUT_P.n1953 VOUT_P.n1928 0.0173591
R19084 VOUT_P.n1132 VOUT_P.n1108 0.0173591
R19085 VOUT_P.n1104 VOUT_P.n1101 0.0173591
R19086 VOUT_P.n1453 VOUT_P.n1132 0.0173591
R19087 VOUT_P.n1913 VOUT_P.n1912 0.0173591
R19088 VOUT_P.n1928 VOUT_P.n1926 0.0173591
R19089 VOUT_P.n1904 VOUT_P.n1903 0.0173591
R19090 VOUT_P.n1452 VOUT_P.n1451 0.0173591
R19091 VOUT_P.n1105 VOUT_P.n1104 0.0173591
R19092 VOUT_P.n1967 VOUT_P.n1966 0.0171202
R19093 VOUT_P.n961 VOUT_P.n957 0.0167343
R19094 VOUT_P.n932 VOUT_P.n931 0.0167343
R19095 VOUT_P.n947 VOUT_P.n946 0.0167343
R19096 VOUT_P.n995 VOUT_P.n994 0.0167343
R19097 VOUT_P.n919 VOUT_P.n918 0.0167343
R19098 VOUT_P.n911 VOUT_P.n910 0.0167343
R19099 VOUT_P.n888 VOUT_P.n887 0.0161314
R19100 VOUT_P.n540 VOUT_P.n539 0.0147026
R19101 VOUT_P.n1085 VOUT_P.n1084 0.0136473
R19102 VOUT_P.n1084 VOUT_P.n1083 0.0136473
R19103 VOUT_P.n1986 VOUT_P.n1985 0.0131984
R19104 VOUT_P.n1985 VOUT_P.n1963 0.0131984
R19105 VOUT_P.n1901 VOUT_P.n1900 0.0130374
R19106 VOUT_P.n1959 VOUT_P.n1958 0.012898
R19107 VOUT_P.n1960 VOUT_P.n1959 0.012898
R19108 VOUT_P.n1902 VOUT_P.n1901 0.0127848
R19109 VOUT_P.n790 VOUT_P.n789 0.0122638
R19110 VOUT_P.n350 VOUT_P.n349 0.0122638
R19111 VOUT_P.n127 VOUT_P.n126 0.0122638
R19112 VOUT_P.n260 VOUT_P.n249 0.0122638
R19113 VOUT_P.n1368 VOUT_P.n1367 0.0122638
R19114 VOUT_P.n1409 VOUT_P.n1408 0.0122638
R19115 VOUT_P.n1450 VOUT_P.n1449 0.0122638
R19116 VOUT_P.n569 VOUT_P.n544 0.0122638
R19117 VOUT_P.n1602 VOUT_P.n1457 0.0122638
R19118 VOUT_P.n1103 VOUT_P.n1102 0.0119325
R19119 VOUT_P.n201 VOUT_P.n200 0.0119325
R19120 VOUT_P.n839 VOUT_P.n838 0.0119325
R19121 VOUT_P.n834 VOUT_P.n833 0.0119325
R19122 VOUT_P.n196 VOUT_P.n195 0.0119325
R19123 VOUT_P.n902 VOUT_P.n901 0.0119325
R19124 VOUT_P.n891 VOUT_P.n890 0.0119325
R19125 VOUT_P.n735 VOUT_P.n734 0.0119325
R19126 VOUT_P.n793 VOUT_P.n777 0.0119325
R19127 VOUT_P.n354 VOUT_P.n353 0.0119325
R19128 VOUT_P.n780 VOUT_P.n779 0.0119325
R19129 VOUT_P.n447 VOUT_P.n446 0.0119325
R19130 VOUT_P.n543 VOUT_P.n542 0.0119325
R19131 VOUT_P.n37 VOUT_P.n36 0.0119325
R19132 VOUT_P.n119 VOUT_P.n118 0.0119325
R19133 VOUT_P.n936 VOUT_P.n935 0.0119325
R19134 VOUT_P.n1570 VOUT_P.n1569 0.0119325
R19135 VOUT_P.n1516 VOUT_P.n1515 0.0119325
R19136 VOUT_P.n1728 VOUT_P.n1727 0.0119325
R19137 VOUT_P.n1815 VOUT_P.n1814 0.0119325
R19138 VOUT_P.n252 VOUT_P.n251 0.0119325
R19139 VOUT_P.n254 VOUT_P.n253 0.0119325
R19140 VOUT_P.n1732 VOUT_P.n1731 0.0119325
R19141 VOUT_P.n1926 VOUT_P.n1925 0.0119325
R19142 VOUT_P.n1920 VOUT_P.n1919 0.0119325
R19143 VOUT_P.n1917 VOUT_P.n1916 0.0119325
R19144 VOUT_P.n1456 VOUT_P.n1455 0.0119325
R19145 VOUT_P.n1101 VOUT_P.n1100 0.0119325
R19146 VOUT_P.n887 VOUT_P.n886 0.0118313
R19147 VOUT_P.n886 VOUT_P.n885 0.0118313
R19148 VOUT_P.n1059 VOUT_P.n1057 0.0110972
R19149 VOUT_P.n1063 VOUT_P.n1060 0.0110972
R19150 VOUT_P.n1094 VOUT_P.n1091 0.0110972
R19151 VOUT_P.n1063 VOUT_P.n1062 0.010845
R19152 VOUT_P.n1059 VOUT_P.n1058 0.010845
R19153 VOUT_P.n1053 VOUT_P.n1052 0.010845
R19154 VOUT_P.n1094 VOUT_P.n1093 0.010845
R19155 VOUT_P.n1087 VOUT_P.n1086 0.010845
R19156 VOUT_P.n1979 VOUT_P.n1978 0.0102276
R19157 VOUT_P.n1015 VOUT_P.n1014 0.00964634
R19158 VOUT_P.n1019 VOUT_P.n1018 0.00964634
R19159 VOUT_P.n1023 VOUT_P.n1022 0.00964634
R19160 VOUT_P.n1027 VOUT_P.n1026 0.00964634
R19161 VOUT_P.n1030 VOUT_P.n1029 0.00964634
R19162 VOUT_P.n1033 VOUT_P.n1032 0.00964634
R19163 VOUT_P.n1036 VOUT_P.n1035 0.00964634
R19164 VOUT_P.n1039 VOUT_P.n1038 0.00964634
R19165 VOUT_P.n1564 VOUT_P.n1563 0.00905634
R19166 VOUT_P.n1534 VOUT_P.n1533 0.00905634
R19167 VOUT_P.n98 VOUT_P.n97 0.00905634
R19168 VOUT_P.n109 VOUT_P.n108 0.00905634
R19169 VOUT_P.n555 VOUT_P.n554 0.00905634
R19170 VOUT_P.n999 VOUT_P.n998 0.00905634
R19171 VOUT_P.n719 VOUT_P.n718 0.00905634
R19172 VOUT_P.n728 VOUT_P.n727 0.00905634
R19173 VOUT_P.n741 VOUT_P.n740 0.00905634
R19174 VOUT_P.n750 VOUT_P.n749 0.00905634
R19175 VOUT_P.n759 VOUT_P.n758 0.00905634
R19176 VOUT_P.n768 VOUT_P.n767 0.00905634
R19177 VOUT_P.n797 VOUT_P.n796 0.00905634
R19178 VOUT_P.n806 VOUT_P.n805 0.00905634
R19179 VOUT_P.n815 VOUT_P.n814 0.00905634
R19180 VOUT_P.n824 VOUT_P.n823 0.00905634
R19181 VOUT_P.n852 VOUT_P.n851 0.00905634
R19182 VOUT_P.n861 VOUT_P.n860 0.00905634
R19183 VOUT_P.n870 VOUT_P.n869 0.00905634
R19184 VOUT_P.n879 VOUT_P.n878 0.00905634
R19185 VOUT_P.n212 VOUT_P.n211 0.00905634
R19186 VOUT_P.n14 VOUT_P.n13 0.00905634
R19187 VOUT_P.n55 VOUT_P.n54 0.00905634
R19188 VOUT_P.n82 VOUT_P.n81 0.00905634
R19189 VOUT_P.n1594 VOUT_P.n1593 0.00905634
R19190 VOUT_P.n1585 VOUT_P.n1584 0.00905634
R19191 VOUT_P.n1576 VOUT_P.n1575 0.00905634
R19192 VOUT_P.n1507 VOUT_P.n1506 0.00905634
R19193 VOUT_P.n1505 VOUT_P.n1504 0.00905634
R19194 VOUT_P.n1717 VOUT_P.n1716 0.00905634
R19195 VOUT_P.n1726 VOUT_P.n1725 0.00905634
R19196 VOUT_P.n1745 VOUT_P.n1744 0.00905634
R19197 VOUT_P.n1754 VOUT_P.n1753 0.00905634
R19198 VOUT_P.n1763 VOUT_P.n1762 0.00905634
R19199 VOUT_P.n1772 VOUT_P.n1771 0.00905634
R19200 VOUT_P.n1785 VOUT_P.n1784 0.00905634
R19201 VOUT_P.n1794 VOUT_P.n1793 0.00905634
R19202 VOUT_P.n1803 VOUT_P.n1802 0.00905634
R19203 VOUT_P.n1812 VOUT_P.n1811 0.00905634
R19204 VOUT_P.n1309 VOUT_P.n1308 0.00905634
R19205 VOUT_P.n1318 VOUT_P.n1317 0.00905634
R19206 VOUT_P.n1336 VOUT_P.n1335 0.00905634
R19207 VOUT_P.n1345 VOUT_P.n1344 0.00905634
R19208 VOUT_P.n1354 VOUT_P.n1353 0.00905634
R19209 VOUT_P.n1363 VOUT_P.n1362 0.00905634
R19210 VOUT_P.n1377 VOUT_P.n1376 0.00905634
R19211 VOUT_P.n1386 VOUT_P.n1385 0.00905634
R19212 VOUT_P.n1395 VOUT_P.n1394 0.00905634
R19213 VOUT_P.n1404 VOUT_P.n1403 0.00905634
R19214 VOUT_P.n1418 VOUT_P.n1417 0.00905634
R19215 VOUT_P.n1427 VOUT_P.n1426 0.00905634
R19216 VOUT_P.n1436 VOUT_P.n1435 0.00905634
R19217 VOUT_P.n1445 VOUT_P.n1444 0.00905634
R19218 VOUT_P.n1123 VOUT_P.n1122 0.00905634
R19219 VOUT_P.n7 VOUT_P.n0 0.00865331
R19220 VOUT_P.n904 VOUT_P.n888 0.00856444
R19221 VOUT_P.n1961 VOUT_P.n1960 0.00805034
R19222 VOUT_P.n1044 VOUT_P.n1043 0.008
R19223 VOUT_P.n1047 VOUT_P.n1046 0.008
R19224 VOUT_P.n1050 VOUT_P.n1049 0.008
R19225 VOUT_P.n1056 VOUT_P.n1055 0.008
R19226 VOUT_P.n1075 VOUT_P.n1074 0.008
R19227 VOUT_P.n1078 VOUT_P.n1077 0.008
R19228 VOUT_P.n1081 VOUT_P.n1080 0.008
R19229 VOUT_P.n1090 VOUT_P.n1089 0.008
R19230 VOUT_P.n1973 VOUT_P.n1972 0.00794621
R19231 VOUT_P.n539 VOUT_P.n538 0.00785132
R19232 VOUT_P.n1945 VOUT_P.n1944 0.00735609
R19233 VOUT_P.n1950 VOUT_P.n1949 0.00735609
R19234 VOUT_P.n568 VOUT_P.n567 0.00735609
R19235 VOUT_P.n966 VOUT_P.n965 0.00735609
R19236 VOUT_P.n528 VOUT_P.n527 0.00735609
R19237 VOUT_P.n517 VOUT_P.n516 0.00735609
R19238 VOUT_P.n506 VOUT_P.n505 0.00735609
R19239 VOUT_P.n495 VOUT_P.n494 0.00735609
R19240 VOUT_P.n484 VOUT_P.n483 0.00735609
R19241 VOUT_P.n473 VOUT_P.n472 0.00735609
R19242 VOUT_P.n462 VOUT_P.n461 0.00735609
R19243 VOUT_P.n451 VOUT_P.n450 0.00735609
R19244 VOUT_P.n436 VOUT_P.n435 0.00735609
R19245 VOUT_P.n425 VOUT_P.n424 0.00735609
R19246 VOUT_P.n414 VOUT_P.n413 0.00735609
R19247 VOUT_P.n403 VOUT_P.n402 0.00735609
R19248 VOUT_P.n392 VOUT_P.n391 0.00735609
R19249 VOUT_P.n381 VOUT_P.n380 0.00735609
R19250 VOUT_P.n370 VOUT_P.n369 0.00735609
R19251 VOUT_P.n359 VOUT_P.n358 0.00735609
R19252 VOUT_P.n339 VOUT_P.n338 0.00735609
R19253 VOUT_P.n328 VOUT_P.n327 0.00735609
R19254 VOUT_P.n317 VOUT_P.n316 0.00735609
R19255 VOUT_P.n306 VOUT_P.n305 0.00735609
R19256 VOUT_P.n295 VOUT_P.n294 0.00735609
R19257 VOUT_P.n284 VOUT_P.n283 0.00735609
R19258 VOUT_P.n273 VOUT_P.n272 0.00735609
R19259 VOUT_P.n262 VOUT_P.n261 0.00735609
R19260 VOUT_P.n236 VOUT_P.n235 0.00735609
R19261 VOUT_P.n225 VOUT_P.n224 0.00735609
R19262 VOUT_P.n214 VOUT_P.n213 0.00735609
R19263 VOUT_P.n1818 VOUT_P.n1817 0.00735609
R19264 VOUT_P.n1828 VOUT_P.n1827 0.00735609
R19265 VOUT_P.n1839 VOUT_P.n1838 0.00735609
R19266 VOUT_P.n1850 VOUT_P.n1849 0.00735609
R19267 VOUT_P.n1859 VOUT_P.n1858 0.00735609
R19268 VOUT_P.n1869 VOUT_P.n1868 0.00735609
R19269 VOUT_P.n1880 VOUT_P.n1879 0.00735609
R19270 VOUT_P.n1891 VOUT_P.n1890 0.00735609
R19271 VOUT_P.n1086 VOUT_P.n1085 0.00732364
R19272 VOUT_P.n1083 VOUT_P.n1082 0.00732364
R19273 VOUT_P.n1017 VOUT_P.n1015 0.00543902
R19274 VOUT_P.n1018 VOUT_P.n1017 0.00543902
R19275 VOUT_P.n1021 VOUT_P.n1019 0.00543902
R19276 VOUT_P.n1022 VOUT_P.n1021 0.00543902
R19277 VOUT_P.n1025 VOUT_P.n1023 0.00543902
R19278 VOUT_P.n1026 VOUT_P.n1025 0.00543902
R19279 VOUT_P.n1028 VOUT_P.n1027 0.00543902
R19280 VOUT_P.n1031 VOUT_P.n1030 0.00543902
R19281 VOUT_P.n1032 VOUT_P.n1031 0.00543902
R19282 VOUT_P.n1034 VOUT_P.n1033 0.00543902
R19283 VOUT_P.n1035 VOUT_P.n1034 0.00543902
R19284 VOUT_P.n1037 VOUT_P.n1036 0.00543902
R19285 VOUT_P.n1038 VOUT_P.n1037 0.00543902
R19286 VOUT_P.n1040 VOUT_P.n1039 0.00543902
R19287 VOUT_P.n1304 VOUT_P.n1303 0.00528925
R19288 VOUT_P.n1308 VOUT_P.n1307 0.00528925
R19289 VOUT_P.n1313 VOUT_P.n1312 0.00528925
R19290 VOUT_P.n1124 VOUT_P.n1123 0.00528925
R19291 VOUT_P.n1128 VOUT_P.n1127 0.00528925
R19292 VOUT_P.n1712 VOUT_P.n1711 0.00528925
R19293 VOUT_P.n1716 VOUT_P.n1715 0.00528925
R19294 VOUT_P.n1721 VOUT_P.n1720 0.00528925
R19295 VOUT_P.n1725 VOUT_P.n1724 0.00528925
R19296 VOUT_P.n1740 VOUT_P.n1739 0.00528925
R19297 VOUT_P.n1744 VOUT_P.n1743 0.00528925
R19298 VOUT_P.n1749 VOUT_P.n1748 0.00528925
R19299 VOUT_P.n1753 VOUT_P.n1752 0.00528925
R19300 VOUT_P.n1758 VOUT_P.n1757 0.00528925
R19301 VOUT_P.n1762 VOUT_P.n1761 0.00528925
R19302 VOUT_P.n1767 VOUT_P.n1766 0.00528925
R19303 VOUT_P.n1771 VOUT_P.n1770 0.00528925
R19304 VOUT_P.n1780 VOUT_P.n1779 0.00528925
R19305 VOUT_P.n1784 VOUT_P.n1783 0.00528925
R19306 VOUT_P.n1789 VOUT_P.n1788 0.00528925
R19307 VOUT_P.n1793 VOUT_P.n1792 0.00528925
R19308 VOUT_P.n1798 VOUT_P.n1797 0.00528925
R19309 VOUT_P.n1802 VOUT_P.n1801 0.00528925
R19310 VOUT_P.n1807 VOUT_P.n1806 0.00528925
R19311 VOUT_P.n1811 VOUT_P.n1810 0.00528925
R19312 VOUT_P.n1599 VOUT_P.n1598 0.00528925
R19313 VOUT_P.n1595 VOUT_P.n1594 0.00528925
R19314 VOUT_P.n1590 VOUT_P.n1589 0.00528925
R19315 VOUT_P.n1586 VOUT_P.n1585 0.00528925
R19316 VOUT_P.n1581 VOUT_P.n1580 0.00528925
R19317 VOUT_P.n1508 VOUT_P.n1507 0.00528925
R19318 VOUT_P.n1512 VOUT_P.n1511 0.00528925
R19319 VOUT_P.n1577 VOUT_P.n1576 0.00528925
R19320 VOUT_P.n1559 VOUT_P.n1558 0.00528925
R19321 VOUT_P.n1535 VOUT_P.n1534 0.00528925
R19322 VOUT_P.n1539 VOUT_P.n1538 0.00528925
R19323 VOUT_P.n1563 VOUT_P.n1562 0.00528925
R19324 VOUT_P.n718 VOUT_P.n717 0.00528925
R19325 VOUT_P.n723 VOUT_P.n722 0.00528925
R19326 VOUT_P.n727 VOUT_P.n726 0.00528925
R19327 VOUT_P.n732 VOUT_P.n731 0.00528925
R19328 VOUT_P.n740 VOUT_P.n739 0.00528925
R19329 VOUT_P.n745 VOUT_P.n744 0.00528925
R19330 VOUT_P.n749 VOUT_P.n748 0.00528925
R19331 VOUT_P.n754 VOUT_P.n753 0.00528925
R19332 VOUT_P.n758 VOUT_P.n757 0.00528925
R19333 VOUT_P.n763 VOUT_P.n762 0.00528925
R19334 VOUT_P.n767 VOUT_P.n766 0.00528925
R19335 VOUT_P.n772 VOUT_P.n771 0.00528925
R19336 VOUT_P.n796 VOUT_P.n795 0.00528925
R19337 VOUT_P.n801 VOUT_P.n800 0.00528925
R19338 VOUT_P.n805 VOUT_P.n804 0.00528925
R19339 VOUT_P.n810 VOUT_P.n809 0.00528925
R19340 VOUT_P.n814 VOUT_P.n813 0.00528925
R19341 VOUT_P.n819 VOUT_P.n818 0.00528925
R19342 VOUT_P.n823 VOUT_P.n822 0.00528925
R19343 VOUT_P.n828 VOUT_P.n827 0.00528925
R19344 VOUT_P.n851 VOUT_P.n850 0.00528925
R19345 VOUT_P.n856 VOUT_P.n855 0.00528925
R19346 VOUT_P.n860 VOUT_P.n859 0.00528925
R19347 VOUT_P.n865 VOUT_P.n864 0.00528925
R19348 VOUT_P.n869 VOUT_P.n868 0.00528925
R19349 VOUT_P.n874 VOUT_P.n873 0.00528925
R19350 VOUT_P.n878 VOUT_P.n877 0.00528925
R19351 VOUT_P.n883 VOUT_P.n882 0.00528925
R19352 VOUT_P.n93 VOUT_P.n92 0.00528925
R19353 VOUT_P.n978 VOUT_P.n977 0.00528925
R19354 VOUT_P.n97 VOUT_P.n96 0.00528925
R19355 VOUT_P.n970 VOUT_P.n969 0.00528925
R19356 VOUT_P.n113 VOUT_P.n112 0.00528925
R19357 VOUT_P.n1003 VOUT_P.n1002 0.00528925
R19358 VOUT_P.n1008 VOUT_P.n1007 0.00528925
R19359 VOUT_P.n54 VOUT_P.n53 0.00528925
R19360 VOUT_P.n59 VOUT_P.n58 0.00528925
R19361 VOUT_P.n83 VOUT_P.n82 0.00528925
R19362 VOUT_P.n79 VOUT_P.n78 0.00528925
R19363 VOUT_P.n1317 VOUT_P.n1316 0.00528925
R19364 VOUT_P.n1331 VOUT_P.n1330 0.00528925
R19365 VOUT_P.n1335 VOUT_P.n1334 0.00528925
R19366 VOUT_P.n1340 VOUT_P.n1339 0.00528925
R19367 VOUT_P.n1344 VOUT_P.n1343 0.00528925
R19368 VOUT_P.n1349 VOUT_P.n1348 0.00528925
R19369 VOUT_P.n1353 VOUT_P.n1352 0.00528925
R19370 VOUT_P.n1358 VOUT_P.n1357 0.00528925
R19371 VOUT_P.n1362 VOUT_P.n1361 0.00528925
R19372 VOUT_P.n1372 VOUT_P.n1371 0.00528925
R19373 VOUT_P.n1376 VOUT_P.n1375 0.00528925
R19374 VOUT_P.n1381 VOUT_P.n1380 0.00528925
R19375 VOUT_P.n1385 VOUT_P.n1384 0.00528925
R19376 VOUT_P.n1390 VOUT_P.n1389 0.00528925
R19377 VOUT_P.n1394 VOUT_P.n1393 0.00528925
R19378 VOUT_P.n1399 VOUT_P.n1398 0.00528925
R19379 VOUT_P.n1403 VOUT_P.n1402 0.00528925
R19380 VOUT_P.n1413 VOUT_P.n1412 0.00528925
R19381 VOUT_P.n1417 VOUT_P.n1416 0.00528925
R19382 VOUT_P.n1422 VOUT_P.n1421 0.00528925
R19383 VOUT_P.n1426 VOUT_P.n1425 0.00528925
R19384 VOUT_P.n1431 VOUT_P.n1430 0.00528925
R19385 VOUT_P.n1435 VOUT_P.n1434 0.00528925
R19386 VOUT_P.n1440 VOUT_P.n1439 0.00528925
R19387 VOUT_P.n1444 VOUT_P.n1443 0.00528925
R19388 VOUT_P.n1947 VOUT_P.n1946 0.00527411
R19389 VOUT_P.n1948 VOUT_P.n1947 0.00527411
R19390 VOUT_P.n1541 VOUT_P.n1540 0.00527411
R19391 VOUT_P.n1540 VOUT_P.n1539 0.00527411
R19392 VOUT_P.n1558 VOUT_P.n1557 0.00527411
R19393 VOUT_P.n111 VOUT_P.n110 0.00527411
R19394 VOUT_P.n92 VOUT_P.n91 0.00527411
R19395 VOUT_P.n112 VOUT_P.n111 0.00527411
R19396 VOUT_P.n557 VOUT_P.n556 0.00527411
R19397 VOUT_P.n566 VOUT_P.n557 0.00527411
R19398 VOUT_P.n1006 VOUT_P.n1005 0.00527411
R19399 VOUT_P.n1001 VOUT_P.n1000 0.00527411
R19400 VOUT_P.n981 VOUT_P.n980 0.00527411
R19401 VOUT_P.n976 VOUT_P.n975 0.00527411
R19402 VOUT_P.n968 VOUT_P.n967 0.00527411
R19403 VOUT_P.n1002 VOUT_P.n1001 0.00527411
R19404 VOUT_P.n977 VOUT_P.n976 0.00527411
R19405 VOUT_P.n969 VOUT_P.n968 0.00527411
R19406 VOUT_P.n998 VOUT_P.n981 0.00527411
R19407 VOUT_P.n1007 VOUT_P.n1006 0.00527411
R19408 VOUT_P.n721 VOUT_P.n720 0.00527411
R19409 VOUT_P.n730 VOUT_P.n729 0.00527411
R19410 VOUT_P.n743 VOUT_P.n742 0.00527411
R19411 VOUT_P.n752 VOUT_P.n751 0.00527411
R19412 VOUT_P.n761 VOUT_P.n760 0.00527411
R19413 VOUT_P.n770 VOUT_P.n769 0.00527411
R19414 VOUT_P.n799 VOUT_P.n798 0.00527411
R19415 VOUT_P.n808 VOUT_P.n807 0.00527411
R19416 VOUT_P.n817 VOUT_P.n816 0.00527411
R19417 VOUT_P.n826 VOUT_P.n825 0.00527411
R19418 VOUT_P.n854 VOUT_P.n853 0.00527411
R19419 VOUT_P.n863 VOUT_P.n862 0.00527411
R19420 VOUT_P.n872 VOUT_P.n871 0.00527411
R19421 VOUT_P.n881 VOUT_P.n880 0.00527411
R19422 VOUT_P.n882 VOUT_P.n881 0.00527411
R19423 VOUT_P.n873 VOUT_P.n872 0.00527411
R19424 VOUT_P.n864 VOUT_P.n863 0.00527411
R19425 VOUT_P.n855 VOUT_P.n854 0.00527411
R19426 VOUT_P.n827 VOUT_P.n826 0.00527411
R19427 VOUT_P.n818 VOUT_P.n817 0.00527411
R19428 VOUT_P.n809 VOUT_P.n808 0.00527411
R19429 VOUT_P.n800 VOUT_P.n799 0.00527411
R19430 VOUT_P.n771 VOUT_P.n770 0.00527411
R19431 VOUT_P.n762 VOUT_P.n761 0.00527411
R19432 VOUT_P.n753 VOUT_P.n752 0.00527411
R19433 VOUT_P.n744 VOUT_P.n743 0.00527411
R19434 VOUT_P.n731 VOUT_P.n730 0.00527411
R19435 VOUT_P.n722 VOUT_P.n721 0.00527411
R19436 VOUT_P.n223 VOUT_P.n222 0.00527411
R19437 VOUT_P.n234 VOUT_P.n233 0.00527411
R19438 VOUT_P.n245 VOUT_P.n244 0.00527411
R19439 VOUT_P.n271 VOUT_P.n270 0.00527411
R19440 VOUT_P.n282 VOUT_P.n281 0.00527411
R19441 VOUT_P.n293 VOUT_P.n292 0.00527411
R19442 VOUT_P.n304 VOUT_P.n303 0.00527411
R19443 VOUT_P.n315 VOUT_P.n314 0.00527411
R19444 VOUT_P.n326 VOUT_P.n325 0.00527411
R19445 VOUT_P.n337 VOUT_P.n336 0.00527411
R19446 VOUT_P.n348 VOUT_P.n347 0.00527411
R19447 VOUT_P.n368 VOUT_P.n367 0.00527411
R19448 VOUT_P.n379 VOUT_P.n378 0.00527411
R19449 VOUT_P.n390 VOUT_P.n389 0.00527411
R19450 VOUT_P.n401 VOUT_P.n400 0.00527411
R19451 VOUT_P.n412 VOUT_P.n411 0.00527411
R19452 VOUT_P.n423 VOUT_P.n422 0.00527411
R19453 VOUT_P.n434 VOUT_P.n433 0.00527411
R19454 VOUT_P.n445 VOUT_P.n444 0.00527411
R19455 VOUT_P.n460 VOUT_P.n459 0.00527411
R19456 VOUT_P.n471 VOUT_P.n470 0.00527411
R19457 VOUT_P.n482 VOUT_P.n481 0.00527411
R19458 VOUT_P.n493 VOUT_P.n492 0.00527411
R19459 VOUT_P.n504 VOUT_P.n503 0.00527411
R19460 VOUT_P.n515 VOUT_P.n514 0.00527411
R19461 VOUT_P.n526 VOUT_P.n525 0.00527411
R19462 VOUT_P.n537 VOUT_P.n536 0.00527411
R19463 VOUT_P.n536 VOUT_P.n535 0.00527411
R19464 VOUT_P.n525 VOUT_P.n524 0.00527411
R19465 VOUT_P.n514 VOUT_P.n513 0.00527411
R19466 VOUT_P.n503 VOUT_P.n502 0.00527411
R19467 VOUT_P.n492 VOUT_P.n491 0.00527411
R19468 VOUT_P.n481 VOUT_P.n480 0.00527411
R19469 VOUT_P.n470 VOUT_P.n469 0.00527411
R19470 VOUT_P.n459 VOUT_P.n458 0.00527411
R19471 VOUT_P.n444 VOUT_P.n443 0.00527411
R19472 VOUT_P.n433 VOUT_P.n432 0.00527411
R19473 VOUT_P.n422 VOUT_P.n421 0.00527411
R19474 VOUT_P.n411 VOUT_P.n410 0.00527411
R19475 VOUT_P.n400 VOUT_P.n399 0.00527411
R19476 VOUT_P.n389 VOUT_P.n388 0.00527411
R19477 VOUT_P.n378 VOUT_P.n377 0.00527411
R19478 VOUT_P.n367 VOUT_P.n366 0.00527411
R19479 VOUT_P.n347 VOUT_P.n346 0.00527411
R19480 VOUT_P.n336 VOUT_P.n335 0.00527411
R19481 VOUT_P.n325 VOUT_P.n324 0.00527411
R19482 VOUT_P.n314 VOUT_P.n313 0.00527411
R19483 VOUT_P.n303 VOUT_P.n302 0.00527411
R19484 VOUT_P.n292 VOUT_P.n291 0.00527411
R19485 VOUT_P.n281 VOUT_P.n280 0.00527411
R19486 VOUT_P.n270 VOUT_P.n269 0.00527411
R19487 VOUT_P.n244 VOUT_P.n243 0.00527411
R19488 VOUT_P.n233 VOUT_P.n232 0.00527411
R19489 VOUT_P.n222 VOUT_P.n221 0.00527411
R19490 VOUT_P.n190 VOUT_P.n189 0.00527411
R19491 VOUT_P.n183 VOUT_P.n182 0.00527411
R19492 VOUT_P.n180 VOUT_P.n179 0.00527411
R19493 VOUT_P.n172 VOUT_P.n171 0.00527411
R19494 VOUT_P.n169 VOUT_P.n168 0.00527411
R19495 VOUT_P.n163 VOUT_P.n162 0.00527411
R19496 VOUT_P.n160 VOUT_P.n159 0.00527411
R19497 VOUT_P.n153 VOUT_P.n152 0.00527411
R19498 VOUT_P.n150 VOUT_P.n149 0.00527411
R19499 VOUT_P.n142 VOUT_P.n141 0.00527411
R19500 VOUT_P.n139 VOUT_P.n138 0.00527411
R19501 VOUT_P.n133 VOUT_P.n132 0.00527411
R19502 VOUT_P.n34 VOUT_P.n33 0.00527411
R19503 VOUT_P.n27 VOUT_P.n26 0.00527411
R19504 VOUT_P.n24 VOUT_P.n23 0.00527411
R19505 VOUT_P.n16 VOUT_P.n15 0.00527411
R19506 VOUT_P.n25 VOUT_P.n24 0.00527411
R19507 VOUT_P.n23 VOUT_P.n16 0.00527411
R19508 VOUT_P.n35 VOUT_P.n34 0.00527411
R19509 VOUT_P.n33 VOUT_P.n27 0.00527411
R19510 VOUT_P.n140 VOUT_P.n139 0.00527411
R19511 VOUT_P.n138 VOUT_P.n133 0.00527411
R19512 VOUT_P.n151 VOUT_P.n150 0.00527411
R19513 VOUT_P.n149 VOUT_P.n142 0.00527411
R19514 VOUT_P.n161 VOUT_P.n160 0.00527411
R19515 VOUT_P.n159 VOUT_P.n153 0.00527411
R19516 VOUT_P.n170 VOUT_P.n169 0.00527411
R19517 VOUT_P.n168 VOUT_P.n163 0.00527411
R19518 VOUT_P.n181 VOUT_P.n180 0.00527411
R19519 VOUT_P.n179 VOUT_P.n172 0.00527411
R19520 VOUT_P.n191 VOUT_P.n190 0.00527411
R19521 VOUT_P.n189 VOUT_P.n183 0.00527411
R19522 VOUT_P.n57 VOUT_P.n56 0.00527411
R19523 VOUT_P.n58 VOUT_P.n57 0.00527411
R19524 VOUT_P.n1601 VOUT_P.n1600 0.00527411
R19525 VOUT_P.n1592 VOUT_P.n1591 0.00527411
R19526 VOUT_P.n1583 VOUT_P.n1582 0.00527411
R19527 VOUT_P.n1514 VOUT_P.n1513 0.00527411
R19528 VOUT_P.n1513 VOUT_P.n1512 0.00527411
R19529 VOUT_P.n1582 VOUT_P.n1581 0.00527411
R19530 VOUT_P.n1591 VOUT_P.n1590 0.00527411
R19531 VOUT_P.n1600 VOUT_P.n1599 0.00527411
R19532 VOUT_P.n1719 VOUT_P.n1718 0.00527411
R19533 VOUT_P.n1738 VOUT_P.n1737 0.00527411
R19534 VOUT_P.n1747 VOUT_P.n1746 0.00527411
R19535 VOUT_P.n1756 VOUT_P.n1755 0.00527411
R19536 VOUT_P.n1765 VOUT_P.n1764 0.00527411
R19537 VOUT_P.n1778 VOUT_P.n1777 0.00527411
R19538 VOUT_P.n1787 VOUT_P.n1786 0.00527411
R19539 VOUT_P.n1796 VOUT_P.n1795 0.00527411
R19540 VOUT_P.n1805 VOUT_P.n1804 0.00527411
R19541 VOUT_P.n1826 VOUT_P.n1825 0.00527411
R19542 VOUT_P.n1837 VOUT_P.n1836 0.00527411
R19543 VOUT_P.n1848 VOUT_P.n1847 0.00527411
R19544 VOUT_P.n1857 VOUT_P.n1856 0.00527411
R19545 VOUT_P.n1867 VOUT_P.n1866 0.00527411
R19546 VOUT_P.n1878 VOUT_P.n1877 0.00527411
R19547 VOUT_P.n1889 VOUT_P.n1888 0.00527411
R19548 VOUT_P.n1898 VOUT_P.n1897 0.00527411
R19549 VOUT_P.n1825 VOUT_P.n1824 0.00527411
R19550 VOUT_P.n1836 VOUT_P.n1835 0.00527411
R19551 VOUT_P.n1847 VOUT_P.n1846 0.00527411
R19552 VOUT_P.n1856 VOUT_P.n1855 0.00527411
R19553 VOUT_P.n1866 VOUT_P.n1865 0.00527411
R19554 VOUT_P.n1877 VOUT_P.n1876 0.00527411
R19555 VOUT_P.n1888 VOUT_P.n1887 0.00527411
R19556 VOUT_P.n1897 VOUT_P.n1896 0.00527411
R19557 VOUT_P.n1806 VOUT_P.n1805 0.00527411
R19558 VOUT_P.n1797 VOUT_P.n1796 0.00527411
R19559 VOUT_P.n1788 VOUT_P.n1787 0.00527411
R19560 VOUT_P.n1779 VOUT_P.n1778 0.00527411
R19561 VOUT_P.n1766 VOUT_P.n1765 0.00527411
R19562 VOUT_P.n1757 VOUT_P.n1756 0.00527411
R19563 VOUT_P.n1748 VOUT_P.n1747 0.00527411
R19564 VOUT_P.n1739 VOUT_P.n1738 0.00527411
R19565 VOUT_P.n1720 VOUT_P.n1719 0.00527411
R19566 VOUT_P.n1711 VOUT_P.n1710 0.00527411
R19567 VOUT_P.n1311 VOUT_P.n1310 0.00527411
R19568 VOUT_P.n1329 VOUT_P.n1328 0.00527411
R19569 VOUT_P.n1338 VOUT_P.n1337 0.00527411
R19570 VOUT_P.n1347 VOUT_P.n1346 0.00527411
R19571 VOUT_P.n1356 VOUT_P.n1355 0.00527411
R19572 VOUT_P.n1370 VOUT_P.n1369 0.00527411
R19573 VOUT_P.n1379 VOUT_P.n1378 0.00527411
R19574 VOUT_P.n1388 VOUT_P.n1387 0.00527411
R19575 VOUT_P.n1397 VOUT_P.n1396 0.00527411
R19576 VOUT_P.n1411 VOUT_P.n1410 0.00527411
R19577 VOUT_P.n1420 VOUT_P.n1419 0.00527411
R19578 VOUT_P.n1429 VOUT_P.n1428 0.00527411
R19579 VOUT_P.n1438 VOUT_P.n1437 0.00527411
R19580 VOUT_P.n1130 VOUT_P.n1129 0.00527411
R19581 VOUT_P.n1439 VOUT_P.n1438 0.00527411
R19582 VOUT_P.n1430 VOUT_P.n1429 0.00527411
R19583 VOUT_P.n1421 VOUT_P.n1420 0.00527411
R19584 VOUT_P.n1412 VOUT_P.n1411 0.00527411
R19585 VOUT_P.n1398 VOUT_P.n1397 0.00527411
R19586 VOUT_P.n1389 VOUT_P.n1388 0.00527411
R19587 VOUT_P.n1380 VOUT_P.n1379 0.00527411
R19588 VOUT_P.n1371 VOUT_P.n1370 0.00527411
R19589 VOUT_P.n1357 VOUT_P.n1356 0.00527411
R19590 VOUT_P.n1348 VOUT_P.n1347 0.00527411
R19591 VOUT_P.n1339 VOUT_P.n1338 0.00527411
R19592 VOUT_P.n1330 VOUT_P.n1329 0.00527411
R19593 VOUT_P.n1129 VOUT_P.n1128 0.00527411
R19594 VOUT_P.n1312 VOUT_P.n1311 0.00527411
R19595 VOUT_P.n1303 VOUT_P.n1302 0.00527411
R19596 VOUT_P.n1560 VOUT_P.n1559 0.00525899
R19597 VOUT_P.n1562 VOUT_P.n1561 0.00525899
R19598 VOUT_P.n1538 VOUT_P.n1537 0.00525899
R19599 VOUT_P.n1536 VOUT_P.n1535 0.00525899
R19600 VOUT_P.n94 VOUT_P.n93 0.00525899
R19601 VOUT_P.n96 VOUT_P.n95 0.00525899
R19602 VOUT_P.n114 VOUT_P.n113 0.00525899
R19603 VOUT_P.n1004 VOUT_P.n1003 0.00525899
R19604 VOUT_P.n979 VOUT_P.n978 0.00525899
R19605 VOUT_P.n971 VOUT_P.n970 0.00525899
R19606 VOUT_P.n1009 VOUT_P.n1008 0.00525899
R19607 VOUT_P.n724 VOUT_P.n723 0.00525899
R19608 VOUT_P.n726 VOUT_P.n725 0.00525899
R19609 VOUT_P.n733 VOUT_P.n732 0.00525899
R19610 VOUT_P.n739 VOUT_P.n738 0.00525899
R19611 VOUT_P.n746 VOUT_P.n745 0.00525899
R19612 VOUT_P.n748 VOUT_P.n747 0.00525899
R19613 VOUT_P.n755 VOUT_P.n754 0.00525899
R19614 VOUT_P.n757 VOUT_P.n756 0.00525899
R19615 VOUT_P.n764 VOUT_P.n763 0.00525899
R19616 VOUT_P.n766 VOUT_P.n765 0.00525899
R19617 VOUT_P.n773 VOUT_P.n772 0.00525899
R19618 VOUT_P.n795 VOUT_P.n794 0.00525899
R19619 VOUT_P.n802 VOUT_P.n801 0.00525899
R19620 VOUT_P.n804 VOUT_P.n803 0.00525899
R19621 VOUT_P.n811 VOUT_P.n810 0.00525899
R19622 VOUT_P.n813 VOUT_P.n812 0.00525899
R19623 VOUT_P.n820 VOUT_P.n819 0.00525899
R19624 VOUT_P.n822 VOUT_P.n821 0.00525899
R19625 VOUT_P.n829 VOUT_P.n828 0.00525899
R19626 VOUT_P.n850 VOUT_P.n849 0.00525899
R19627 VOUT_P.n857 VOUT_P.n856 0.00525899
R19628 VOUT_P.n859 VOUT_P.n858 0.00525899
R19629 VOUT_P.n866 VOUT_P.n865 0.00525899
R19630 VOUT_P.n868 VOUT_P.n867 0.00525899
R19631 VOUT_P.n875 VOUT_P.n874 0.00525899
R19632 VOUT_P.n877 VOUT_P.n876 0.00525899
R19633 VOUT_P.n884 VOUT_P.n883 0.00525899
R19634 VOUT_P.n60 VOUT_P.n59 0.00525899
R19635 VOUT_P.n84 VOUT_P.n83 0.00525899
R19636 VOUT_P.n80 VOUT_P.n79 0.00525899
R19637 VOUT_P.n1598 VOUT_P.n1597 0.00525899
R19638 VOUT_P.n1596 VOUT_P.n1595 0.00525899
R19639 VOUT_P.n1589 VOUT_P.n1588 0.00525899
R19640 VOUT_P.n1587 VOUT_P.n1586 0.00525899
R19641 VOUT_P.n1580 VOUT_P.n1579 0.00525899
R19642 VOUT_P.n1578 VOUT_P.n1577 0.00525899
R19643 VOUT_P.n1511 VOUT_P.n1510 0.00525899
R19644 VOUT_P.n1509 VOUT_P.n1508 0.00525899
R19645 VOUT_P.n1713 VOUT_P.n1712 0.00525899
R19646 VOUT_P.n1715 VOUT_P.n1714 0.00525899
R19647 VOUT_P.n1722 VOUT_P.n1721 0.00525899
R19648 VOUT_P.n1724 VOUT_P.n1723 0.00525899
R19649 VOUT_P.n1741 VOUT_P.n1740 0.00525899
R19650 VOUT_P.n1743 VOUT_P.n1742 0.00525899
R19651 VOUT_P.n1750 VOUT_P.n1749 0.00525899
R19652 VOUT_P.n1752 VOUT_P.n1751 0.00525899
R19653 VOUT_P.n1759 VOUT_P.n1758 0.00525899
R19654 VOUT_P.n1761 VOUT_P.n1760 0.00525899
R19655 VOUT_P.n1768 VOUT_P.n1767 0.00525899
R19656 VOUT_P.n1770 VOUT_P.n1769 0.00525899
R19657 VOUT_P.n1781 VOUT_P.n1780 0.00525899
R19658 VOUT_P.n1783 VOUT_P.n1782 0.00525899
R19659 VOUT_P.n1790 VOUT_P.n1789 0.00525899
R19660 VOUT_P.n1792 VOUT_P.n1791 0.00525899
R19661 VOUT_P.n1799 VOUT_P.n1798 0.00525899
R19662 VOUT_P.n1801 VOUT_P.n1800 0.00525899
R19663 VOUT_P.n1808 VOUT_P.n1807 0.00525899
R19664 VOUT_P.n1810 VOUT_P.n1809 0.00525899
R19665 VOUT_P.n1305 VOUT_P.n1304 0.00525899
R19666 VOUT_P.n1307 VOUT_P.n1306 0.00525899
R19667 VOUT_P.n1314 VOUT_P.n1313 0.00525899
R19668 VOUT_P.n1316 VOUT_P.n1315 0.00525899
R19669 VOUT_P.n1332 VOUT_P.n1331 0.00525899
R19670 VOUT_P.n1334 VOUT_P.n1333 0.00525899
R19671 VOUT_P.n1341 VOUT_P.n1340 0.00525899
R19672 VOUT_P.n1343 VOUT_P.n1342 0.00525899
R19673 VOUT_P.n1350 VOUT_P.n1349 0.00525899
R19674 VOUT_P.n1352 VOUT_P.n1351 0.00525899
R19675 VOUT_P.n1359 VOUT_P.n1358 0.00525899
R19676 VOUT_P.n1361 VOUT_P.n1360 0.00525899
R19677 VOUT_P.n1373 VOUT_P.n1372 0.00525899
R19678 VOUT_P.n1375 VOUT_P.n1374 0.00525899
R19679 VOUT_P.n1382 VOUT_P.n1381 0.00525899
R19680 VOUT_P.n1384 VOUT_P.n1383 0.00525899
R19681 VOUT_P.n1391 VOUT_P.n1390 0.00525899
R19682 VOUT_P.n1393 VOUT_P.n1392 0.00525899
R19683 VOUT_P.n1400 VOUT_P.n1399 0.00525899
R19684 VOUT_P.n1402 VOUT_P.n1401 0.00525899
R19685 VOUT_P.n1414 VOUT_P.n1413 0.00525899
R19686 VOUT_P.n1416 VOUT_P.n1415 0.00525899
R19687 VOUT_P.n1423 VOUT_P.n1422 0.00525899
R19688 VOUT_P.n1425 VOUT_P.n1424 0.00525899
R19689 VOUT_P.n1432 VOUT_P.n1431 0.00525899
R19690 VOUT_P.n1434 VOUT_P.n1433 0.00525899
R19691 VOUT_P.n1441 VOUT_P.n1440 0.00525899
R19692 VOUT_P.n1443 VOUT_P.n1442 0.00525899
R19693 VOUT_P.n1127 VOUT_P.n1126 0.00525899
R19694 VOUT_P.n1125 VOUT_P.n1124 0.00525899
R19695 VOUT_P.n5 VOUT_P.n4 0.00522947
R19696 VOUT_P.n6 VOUT_P.n5 0.00522947
R19697 VOUT_P.n1977 VOUT_P.n1976 0.00507926
R19698 VOUT_P.n3 VOUT_P.n1 0.00490313
R19699 VOUT_P.n1968 VOUT_P.n1967 0.00475992
R19700 VOUT_P.n1969 VOUT_P.n1968 0.00475992
R19701 VOUT_P.n1982 VOUT_P.n1981 0.00460338
R19702 VOUT_P.n1981 VOUT_P.n1980 0.00460338
R19703 VOUT_P.n1043 VOUT_P.n1042 0.00455
R19704 VOUT_P.n1045 VOUT_P.n1044 0.00455
R19705 VOUT_P.n1046 VOUT_P.n1045 0.00455
R19706 VOUT_P.n1048 VOUT_P.n1047 0.00455
R19707 VOUT_P.n1049 VOUT_P.n1048 0.00455
R19708 VOUT_P.n1054 VOUT_P.n1050 0.00455
R19709 VOUT_P.n1055 VOUT_P.n1054 0.00455
R19710 VOUT_P.n1064 VOUT_P.n1056 0.00455
R19711 VOUT_P.n1074 VOUT_P.n1073 0.00455
R19712 VOUT_P.n1076 VOUT_P.n1075 0.00455
R19713 VOUT_P.n1077 VOUT_P.n1076 0.00455
R19714 VOUT_P.n1079 VOUT_P.n1078 0.00455
R19715 VOUT_P.n1080 VOUT_P.n1079 0.00455
R19716 VOUT_P.n1088 VOUT_P.n1081 0.00455
R19717 VOUT_P.n1089 VOUT_P.n1088 0.00455
R19718 VOUT_P.n1095 VOUT_P.n1090 0.00455
R19719 VOUT_P.n1971 VOUT_P.n1970 0.00437476
R19720 VOUT_P.n1987 VOUT_P.n1986 0.0043197
R19721 VOUT_P.n1988 VOUT_P.n1987 0.0043197
R19722 VOUT_P.n1955 VOUT_P.n1954 0.00429028
R19723 VOUT_P.n1956 VOUT_P.n1955 0.00429028
R19724 VOUT_P.n1949 VOUT_P.n1948 0.00418876
R19725 VOUT_P.n1944 VOUT_P.n1943 0.00418876
R19726 VOUT_P.n567 VOUT_P.n566 0.00418876
R19727 VOUT_P.n965 VOUT_P.n964 0.00418876
R19728 VOUT_P.n221 VOUT_P.n214 0.00418876
R19729 VOUT_P.n232 VOUT_P.n225 0.00418876
R19730 VOUT_P.n243 VOUT_P.n236 0.00418876
R19731 VOUT_P.n269 VOUT_P.n262 0.00418876
R19732 VOUT_P.n280 VOUT_P.n273 0.00418876
R19733 VOUT_P.n291 VOUT_P.n284 0.00418876
R19734 VOUT_P.n302 VOUT_P.n295 0.00418876
R19735 VOUT_P.n313 VOUT_P.n306 0.00418876
R19736 VOUT_P.n324 VOUT_P.n317 0.00418876
R19737 VOUT_P.n335 VOUT_P.n328 0.00418876
R19738 VOUT_P.n346 VOUT_P.n339 0.00418876
R19739 VOUT_P.n366 VOUT_P.n359 0.00418876
R19740 VOUT_P.n377 VOUT_P.n370 0.00418876
R19741 VOUT_P.n388 VOUT_P.n381 0.00418876
R19742 VOUT_P.n399 VOUT_P.n392 0.00418876
R19743 VOUT_P.n410 VOUT_P.n403 0.00418876
R19744 VOUT_P.n421 VOUT_P.n414 0.00418876
R19745 VOUT_P.n432 VOUT_P.n425 0.00418876
R19746 VOUT_P.n443 VOUT_P.n436 0.00418876
R19747 VOUT_P.n458 VOUT_P.n451 0.00418876
R19748 VOUT_P.n469 VOUT_P.n462 0.00418876
R19749 VOUT_P.n480 VOUT_P.n473 0.00418876
R19750 VOUT_P.n491 VOUT_P.n484 0.00418876
R19751 VOUT_P.n502 VOUT_P.n495 0.00418876
R19752 VOUT_P.n513 VOUT_P.n506 0.00418876
R19753 VOUT_P.n524 VOUT_P.n517 0.00418876
R19754 VOUT_P.n535 VOUT_P.n528 0.00418876
R19755 VOUT_P.n1824 VOUT_P.n1818 0.00418876
R19756 VOUT_P.n1835 VOUT_P.n1828 0.00418876
R19757 VOUT_P.n1846 VOUT_P.n1839 0.00418876
R19758 VOUT_P.n1855 VOUT_P.n1850 0.00418876
R19759 VOUT_P.n1865 VOUT_P.n1859 0.00418876
R19760 VOUT_P.n1876 VOUT_P.n1869 0.00418876
R19761 VOUT_P.n1887 VOUT_P.n1880 0.00418876
R19762 VOUT_P.n1896 VOUT_P.n1891 0.00418876
R19763 VOUT_P.n13 VOUT_P.n12 0.00418126
R19764 VOUT_P.n1965 VOUT_P.n1964 0.00413371
R19765 VOUT_P.n1966 VOUT_P.n1965 0.00413371
R19766 VOUT_P.n78 VOUT_P.n77 0.00281899
R19767 VOUT_P.n1957 VOUT_P.n1956 0.00269512
R19768 VOUT_P.n1943 VOUT_P.n1942 0.00219433
R19769 VOUT_P.n964 VOUT_P.n963 0.00219433
R19770 VOUT_P.n108 VOUT_P.n107 0.00192237
R19771 VOUT_P.n554 VOUT_P.n553 0.00192237
R19772 VOUT_P.n1504 VOUT_P.n1503 0.00192237
R19773 VOUT_P.n211 VOUT_P.n210 0.00192078
R19774 VOUT_P.n1065 VOUT_P.n1064 0.00180358
R19775 VOUT_P.n1096 VOUT_P.n1095 0.00180358
R19776 VOUT_P.n1073 VOUT_P.n1072 0.00180358
R19777 VOUT_P.n1984 VOUT_P.n1969 0.00175436
R19778 VOUT_P.n1989 VOUT_P.n1988 0.00170805
R19779 VOUT_P.n1972 VOUT_P.n1971 0.00155675
R19780 VOUT_P.n1983 VOUT_P.n1982 0.00147033
R19781 VOUT_P.n1984 VOUT_P.n1983 0.00147033
R19782 VOUT_P.n1962 VOUT_P.n1961 0.001151
R19783 VOUT_P.n1963 VOUT_P.n1962 0.001151
R19784 VOUT_P.n3 VOUT_P.n2 0.00102838
R19785 VOUT_P.n1978 VOUT_P.n1977 0.00085225
R19786 VOUT_P.n7 VOUT_P.n6 0.000813589
R19787 Folded_Diff_Op_Amp_Layout_0.VOUT.n0 Folded_Diff_Op_Amp_Layout_0.VOUT.t1 3.46869
R19788 Folded_Diff_Op_Amp_Layout_0.VOUT.n0 Folded_Diff_Op_Amp_Layout_0.VOUT.t0 7.1411
R19789 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.VOUT.n0 9.35924
R19790 Folded_Diff_Op_Amp_Layout_0.VOUT.n3 Folded_Diff_Op_Amp_Layout_0.VOUT.n7 0.00773989
R19791 Folded_Diff_Op_Amp_Layout_0.VOUT.n1 Folded_Diff_Op_Amp_Layout_0.VOUT.n2 1.126
R19792 Folded_Diff_Op_Amp_Layout_0.VOUT.n8 Folded_Diff_Op_Amp_Layout_0.VOUT.n4 0.00582347
R19793 Folded_Diff_Op_Amp_Layout_0.VOUT.n1 Folded_Diff_Op_Amp_Layout_0.VOUT.n16 1.12675
R19794 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.VOUT.n1 0.111701
R19795 Folded_Diff_Op_Amp_Layout_0.VOUT.n8 Folded_Diff_Op_Amp_Layout_0.VOUT.n13 0.0236139
R19796 Folded_Diff_Op_Amp_Layout_0.VOUT.n16 Folded_Diff_Op_Amp_Layout_0.VOUT.n14 1.49801
R19797 Folded_Diff_Op_Amp_Layout_0.VOUT.n2 Folded_Diff_Op_Amp_Layout_0.VOUT.n8 1.49812
R19798 Folded_Diff_Op_Amp_Layout_0.VOUT.n3 Folded_Diff_Op_Amp_Layout_0.VOUT.n9 0.00773989
R19799 Folded_Diff_Op_Amp_Layout_0.VOUT.n15 Folded_Diff_Op_Amp_Layout_0.VOUT.n3 1.49801
R19800 Folded_Diff_Op_Amp_Layout_0.VOUT.n9 Folded_Diff_Op_Amp_Layout_0.VOUT.n10 0.00773989
R19801 Folded_Diff_Op_Amp_Layout_0.VOUT.n10 Folded_Diff_Op_Amp_Layout_0.VOUT.n44 5.09856
R19802 Folded_Diff_Op_Amp_Layout_0.VOUT.n42 Folded_Diff_Op_Amp_Layout_0.VOUT.n36 4.31354
R19803 Folded_Diff_Op_Amp_Layout_0.VOUT.n44 Folded_Diff_Op_Amp_Layout_0.VOUT.n42 0.626587
R19804 Folded_Diff_Op_Amp_Layout_0.VOUT.n44 Folded_Diff_Op_Amp_Layout_0.VOUT.t21 36.7201
R19805 Folded_Diff_Op_Amp_Layout_0.VOUT.n42 Folded_Diff_Op_Amp_Layout_0.VOUT.n43 14.2987
R19806 Folded_Diff_Op_Amp_Layout_0.VOUT.n43 Folded_Diff_Op_Amp_Layout_0.VOUT.t10 38.3255
R19807 Folded_Diff_Op_Amp_Layout_0.VOUT.n43 Folded_Diff_Op_Amp_Layout_0.VOUT.t8 17.4684
R19808 Folded_Diff_Op_Amp_Layout_0.VOUT.n41 Folded_Diff_Op_Amp_Layout_0.VOUT.n40 20.8576
R19809 Folded_Diff_Op_Amp_Layout_0.VOUT.n36 Folded_Diff_Op_Amp_Layout_0.VOUT.n41 19.8148
R19810 Folded_Diff_Op_Amp_Layout_0.VOUT.n41 Folded_Diff_Op_Amp_Layout_0.VOUT.t3 30.113
R19811 Folded_Diff_Op_Amp_Layout_0.VOUT.n40 Folded_Diff_Op_Amp_Layout_0.VOUT.t9 30.113
R19812 Folded_Diff_Op_Amp_Layout_0.VOUT.n40 Folded_Diff_Op_Amp_Layout_0.VOUT.n37 19.8148
R19813 Folded_Diff_Op_Amp_Layout_0.VOUT.n38 Folded_Diff_Op_Amp_Layout_0.VOUT.t18 37.0332
R19814 Folded_Diff_Op_Amp_Layout_0.VOUT.n37 Folded_Diff_Op_Amp_Layout_0.VOUT.n38 4.62659
R19815 Folded_Diff_Op_Amp_Layout_0.VOUT.n38 Folded_Diff_Op_Amp_Layout_0.VOUT.n39 14.2987
R19816 Folded_Diff_Op_Amp_Layout_0.VOUT.n39 Folded_Diff_Op_Amp_Layout_0.VOUT.t7 38.3255
R19817 Folded_Diff_Op_Amp_Layout_0.VOUT.n39 Folded_Diff_Op_Amp_Layout_0.VOUT.t29 17.4684
R19818 Folded_Diff_Op_Amp_Layout_0.VOUT.n37 Folded_Diff_Op_Amp_Layout_0.VOUT.t12 29.0701
R19819 Folded_Diff_Op_Amp_Layout_0.VOUT.n36 Folded_Diff_Op_Amp_Layout_0.VOUT.t23 29.0701
R19820 Folded_Diff_Op_Amp_Layout_0.VOUT.n2 Folded_Diff_Op_Amp_Layout_0.VOUT.n5 0.014
R19821 Folded_Diff_Op_Amp_Layout_0.VOUT.n2 Folded_Diff_Op_Amp_Layout_0.VOUT.n6 0.014
R19822 Folded_Diff_Op_Amp_Layout_0.VOUT.n6 Folded_Diff_Op_Amp_Layout_0.VOUT.n11 0.0134654
R19823 Folded_Diff_Op_Amp_Layout_0.VOUT.n16 Folded_Diff_Op_Amp_Layout_0.VOUT.n12 0.014
R19824 Folded_Diff_Op_Amp_Layout_0.VOUT.n16 Folded_Diff_Op_Amp_Layout_0.VOUT.n15 0.00549102
R19825 Folded_Diff_Op_Amp_Layout_0.VOUT.n17 Folded_Diff_Op_Amp_Layout_0.VOUT.n27 4.77125
R19826 Folded_Diff_Op_Amp_Layout_0.VOUT.n17 Folded_Diff_Op_Amp_Layout_0.VOUT.n18 4.17447
R19827 Folded_Diff_Op_Amp_Layout_0.VOUT.n5 Folded_Diff_Op_Amp_Layout_0.VOUT.n17 0.546814
R19828 Folded_Diff_Op_Amp_Layout_0.VOUT.n28 Folded_Diff_Op_Amp_Layout_0.VOUT.n30 4.31354
R19829 Folded_Diff_Op_Amp_Layout_0.VOUT.n27 Folded_Diff_Op_Amp_Layout_0.VOUT.n28 0.623815
R19830 Folded_Diff_Op_Amp_Layout_0.VOUT.n30 Folded_Diff_Op_Amp_Layout_0.VOUT.t28 34.9362
R19831 Folded_Diff_Op_Amp_Layout_0.VOUT.n30 Folded_Diff_Op_Amp_Layout_0.VOUT.n35 13.9445
R19832 Folded_Diff_Op_Amp_Layout_0.VOUT.n35 Folded_Diff_Op_Amp_Layout_0.VOUT.t6 36.2398
R19833 Folded_Diff_Op_Amp_Layout_0.VOUT.n35 Folded_Diff_Op_Amp_Layout_0.VOUT.n34 14.8868
R19834 Folded_Diff_Op_Amp_Layout_0.VOUT.n34 Folded_Diff_Op_Amp_Layout_0.VOUT.t16 36.2398
R19835 Folded_Diff_Op_Amp_Layout_0.VOUT.n34 Folded_Diff_Op_Amp_Layout_0.VOUT.n31 13.9445
R19836 Folded_Diff_Op_Amp_Layout_0.VOUT.n31 Folded_Diff_Op_Amp_Layout_0.VOUT.t17 34.9362
R19837 Folded_Diff_Op_Amp_Layout_0.VOUT.n32 Folded_Diff_Op_Amp_Layout_0.VOUT.t25 39.2493
R19838 Folded_Diff_Op_Amp_Layout_0.VOUT.n31 Folded_Diff_Op_Amp_Layout_0.VOUT.n32 4.62659
R19839 Folded_Diff_Op_Amp_Layout_0.VOUT.n32 Folded_Diff_Op_Amp_Layout_0.VOUT.n33 13.9076
R19840 Folded_Diff_Op_Amp_Layout_0.VOUT.n33 Folded_Diff_Op_Amp_Layout_0.VOUT.t20 36.5005
R19841 Folded_Diff_Op_Amp_Layout_0.VOUT.n33 Folded_Diff_Op_Amp_Layout_0.VOUT.t13 15.6434
R19842 Folded_Diff_Op_Amp_Layout_0.VOUT.n28 Folded_Diff_Op_Amp_Layout_0.VOUT.n29 13.9076
R19843 Folded_Diff_Op_Amp_Layout_0.VOUT.n29 Folded_Diff_Op_Amp_Layout_0.VOUT.t26 36.5005
R19844 Folded_Diff_Op_Amp_Layout_0.VOUT.n29 Folded_Diff_Op_Amp_Layout_0.VOUT.t24 15.6434
R19845 Folded_Diff_Op_Amp_Layout_0.VOUT.n27 Folded_Diff_Op_Amp_Layout_0.VOUT.t27 38.6755
R19846 Folded_Diff_Op_Amp_Layout_0.VOUT.n18 Folded_Diff_Op_Amp_Layout_0.VOUT.t14 37.8216
R19847 Folded_Diff_Op_Amp_Layout_0.VOUT.n18 Folded_Diff_Op_Amp_Layout_0.VOUT.n19 0.592658
R19848 Folded_Diff_Op_Amp_Layout_0.VOUT.n19 Folded_Diff_Op_Amp_Layout_0.VOUT.n21 4.31354
R19849 Folded_Diff_Op_Amp_Layout_0.VOUT.n21 Folded_Diff_Op_Amp_Layout_0.VOUT.t15 34.9362
R19850 Folded_Diff_Op_Amp_Layout_0.VOUT.n21 Folded_Diff_Op_Amp_Layout_0.VOUT.n26 13.9445
R19851 Folded_Diff_Op_Amp_Layout_0.VOUT.n26 Folded_Diff_Op_Amp_Layout_0.VOUT.t22 36.2398
R19852 Folded_Diff_Op_Amp_Layout_0.VOUT.n26 Folded_Diff_Op_Amp_Layout_0.VOUT.n25 14.8868
R19853 Folded_Diff_Op_Amp_Layout_0.VOUT.n25 Folded_Diff_Op_Amp_Layout_0.VOUT.t31 36.2398
R19854 Folded_Diff_Op_Amp_Layout_0.VOUT.n25 Folded_Diff_Op_Amp_Layout_0.VOUT.n22 13.9445
R19855 Folded_Diff_Op_Amp_Layout_0.VOUT.n22 Folded_Diff_Op_Amp_Layout_0.VOUT.t4 34.9362
R19856 Folded_Diff_Op_Amp_Layout_0.VOUT.n23 Folded_Diff_Op_Amp_Layout_0.VOUT.t11 39.2493
R19857 Folded_Diff_Op_Amp_Layout_0.VOUT.n22 Folded_Diff_Op_Amp_Layout_0.VOUT.n23 4.62659
R19858 Folded_Diff_Op_Amp_Layout_0.VOUT.n23 Folded_Diff_Op_Amp_Layout_0.VOUT.n24 13.9076
R19859 Folded_Diff_Op_Amp_Layout_0.VOUT.n24 Folded_Diff_Op_Amp_Layout_0.VOUT.t30 36.5005
R19860 Folded_Diff_Op_Amp_Layout_0.VOUT.n24 Folded_Diff_Op_Amp_Layout_0.VOUT.t19 15.6434
R19861 Folded_Diff_Op_Amp_Layout_0.VOUT.n19 Folded_Diff_Op_Amp_Layout_0.VOUT.n20 13.9076
R19862 Folded_Diff_Op_Amp_Layout_0.VOUT.n20 Folded_Diff_Op_Amp_Layout_0.VOUT.t5 36.5005
R19863 Folded_Diff_Op_Amp_Layout_0.VOUT.n20 Folded_Diff_Op_Amp_Layout_0.VOUT.t2 15.6434
R19864 Folded_Diff_Op_Amp_Layout_0.VCD.n184 Folded_Diff_Op_Amp_Layout_0.VCD.n183 4.27746
R19865 Folded_Diff_Op_Amp_Layout_0.VCD.n184 Folded_Diff_Op_Amp_Layout_0.VCD.n181 3.43224
R19866 Folded_Diff_Op_Amp_Layout_0.VCD.n186 Folded_Diff_Op_Amp_Layout_0.VCD.n185 2.39976
R19867 Folded_Diff_Op_Amp_Layout_0.VCD.n13 Folded_Diff_Op_Amp_Layout_0.VCD.n10 2.24691
R19868 Folded_Diff_Op_Amp_Layout_0.VCD.n22 Folded_Diff_Op_Amp_Layout_0.VCD.n19 2.24691
R19869 Folded_Diff_Op_Amp_Layout_0.VCD.n37 Folded_Diff_Op_Amp_Layout_0.VCD.n34 2.24691
R19870 Folded_Diff_Op_Amp_Layout_0.VCD.n46 Folded_Diff_Op_Amp_Layout_0.VCD.n43 2.24691
R19871 Folded_Diff_Op_Amp_Layout_0.VCD.n174 Folded_Diff_Op_Amp_Layout_0.VCD.n171 2.24691
R19872 Folded_Diff_Op_Amp_Layout_0.VCD.n103 Folded_Diff_Op_Amp_Layout_0.VCD.n102 2.15529
R19873 Folded_Diff_Op_Amp_Layout_0.VCD.n66 Folded_Diff_Op_Amp_Layout_0.VCD.t30 1.6385
R19874 Folded_Diff_Op_Amp_Layout_0.VCD.n66 Folded_Diff_Op_Amp_Layout_0.VCD.n65 1.6385
R19875 Folded_Diff_Op_Amp_Layout_0.VCD.n56 Folded_Diff_Op_Amp_Layout_0.VCD.t50 1.6385
R19876 Folded_Diff_Op_Amp_Layout_0.VCD.n56 Folded_Diff_Op_Amp_Layout_0.VCD.n55 1.6385
R19877 Folded_Diff_Op_Amp_Layout_0.VCD.n118 Folded_Diff_Op_Amp_Layout_0.VCD.t40 1.6385
R19878 Folded_Diff_Op_Amp_Layout_0.VCD.n118 Folded_Diff_Op_Amp_Layout_0.VCD.n117 1.6385
R19879 Folded_Diff_Op_Amp_Layout_0.VCD.n83 Folded_Diff_Op_Amp_Layout_0.VCD.t9 1.6385
R19880 Folded_Diff_Op_Amp_Layout_0.VCD.n83 Folded_Diff_Op_Amp_Layout_0.VCD.n82 1.6385
R19881 Folded_Diff_Op_Amp_Layout_0.VCD.n106 Folded_Diff_Op_Amp_Layout_0.VCD.t4 1.6385
R19882 Folded_Diff_Op_Amp_Layout_0.VCD.n106 Folded_Diff_Op_Amp_Layout_0.VCD.n105 1.6385
R19883 Folded_Diff_Op_Amp_Layout_0.VCD.n102 Folded_Diff_Op_Amp_Layout_0.VCD.t35 1.6385
R19884 Folded_Diff_Op_Amp_Layout_0.VCD.n102 Folded_Diff_Op_Amp_Layout_0.VCD.n101 1.6385
R19885 Folded_Diff_Op_Amp_Layout_0.VCD.n95 Folded_Diff_Op_Amp_Layout_0.VCD.t42 1.6385
R19886 Folded_Diff_Op_Amp_Layout_0.VCD.n95 Folded_Diff_Op_Amp_Layout_0.VCD.n94 1.6385
R19887 Folded_Diff_Op_Amp_Layout_0.VCD.n87 Folded_Diff_Op_Amp_Layout_0.VCD.t13 1.6385
R19888 Folded_Diff_Op_Amp_Layout_0.VCD.n87 Folded_Diff_Op_Amp_Layout_0.VCD.n86 1.6385
R19889 Folded_Diff_Op_Amp_Layout_0.VCD.n161 Folded_Diff_Op_Amp_Layout_0.VCD.t5 1.6385
R19890 Folded_Diff_Op_Amp_Layout_0.VCD.n161 Folded_Diff_Op_Amp_Layout_0.VCD.n160 1.6385
R19891 Folded_Diff_Op_Amp_Layout_0.VCD.n155 Folded_Diff_Op_Amp_Layout_0.VCD.t49 1.6385
R19892 Folded_Diff_Op_Amp_Layout_0.VCD.n155 Folded_Diff_Op_Amp_Layout_0.VCD.n154 1.6385
R19893 Folded_Diff_Op_Amp_Layout_0.VCD.n141 Folded_Diff_Op_Amp_Layout_0.VCD.t10 1.6385
R19894 Folded_Diff_Op_Amp_Layout_0.VCD.n141 Folded_Diff_Op_Amp_Layout_0.VCD.n140 1.6385
R19895 Folded_Diff_Op_Amp_Layout_0.VCD.n133 Folded_Diff_Op_Amp_Layout_0.VCD.t37 1.6385
R19896 Folded_Diff_Op_Amp_Layout_0.VCD.n133 Folded_Diff_Op_Amp_Layout_0.VCD.n132 1.6385
R19897 Folded_Diff_Op_Amp_Layout_0.VCD.n125 Folded_Diff_Op_Amp_Layout_0.VCD.t61 1.6385
R19898 Folded_Diff_Op_Amp_Layout_0.VCD.n125 Folded_Diff_Op_Amp_Layout_0.VCD.n124 1.6385
R19899 Folded_Diff_Op_Amp_Layout_0.VCD.n150 Folded_Diff_Op_Amp_Layout_0.VCD.t0 1.6385
R19900 Folded_Diff_Op_Amp_Layout_0.VCD.n150 Folded_Diff_Op_Amp_Layout_0.VCD.n149 1.6385
R19901 Folded_Diff_Op_Amp_Layout_0.VCD.n167 Folded_Diff_Op_Amp_Layout_0.VCD.t31 1.6385
R19902 Folded_Diff_Op_Amp_Layout_0.VCD.n167 Folded_Diff_Op_Amp_Layout_0.VCD.n166 1.6385
R19903 Folded_Diff_Op_Amp_Layout_0.VCD.n7 Folded_Diff_Op_Amp_Layout_0.VCD.t7 1.6385
R19904 Folded_Diff_Op_Amp_Layout_0.VCD.n7 Folded_Diff_Op_Amp_Layout_0.VCD.n6 1.6385
R19905 Folded_Diff_Op_Amp_Layout_0.VCD.n12 Folded_Diff_Op_Amp_Layout_0.VCD.t55 1.6385
R19906 Folded_Diff_Op_Amp_Layout_0.VCD.n12 Folded_Diff_Op_Amp_Layout_0.VCD.n11 1.6385
R19907 Folded_Diff_Op_Amp_Layout_0.VCD.n10 Folded_Diff_Op_Amp_Layout_0.VCD.t1 1.6385
R19908 Folded_Diff_Op_Amp_Layout_0.VCD.n10 Folded_Diff_Op_Amp_Layout_0.VCD.n9 1.6385
R19909 Folded_Diff_Op_Amp_Layout_0.VCD.n26 Folded_Diff_Op_Amp_Layout_0.VCD.t52 1.6385
R19910 Folded_Diff_Op_Amp_Layout_0.VCD.n26 Folded_Diff_Op_Amp_Layout_0.VCD.n25 1.6385
R19911 Folded_Diff_Op_Amp_Layout_0.VCD.n21 Folded_Diff_Op_Amp_Layout_0.VCD.t2 1.6385
R19912 Folded_Diff_Op_Amp_Layout_0.VCD.n21 Folded_Diff_Op_Amp_Layout_0.VCD.n20 1.6385
R19913 Folded_Diff_Op_Amp_Layout_0.VCD.n19 Folded_Diff_Op_Amp_Layout_0.VCD.t58 1.6385
R19914 Folded_Diff_Op_Amp_Layout_0.VCD.n19 Folded_Diff_Op_Amp_Layout_0.VCD.n18 1.6385
R19915 Folded_Diff_Op_Amp_Layout_0.VCD.n31 Folded_Diff_Op_Amp_Layout_0.VCD.t3 1.6385
R19916 Folded_Diff_Op_Amp_Layout_0.VCD.n31 Folded_Diff_Op_Amp_Layout_0.VCD.n30 1.6385
R19917 Folded_Diff_Op_Amp_Layout_0.VCD.n36 Folded_Diff_Op_Amp_Layout_0.VCD.t33 1.6385
R19918 Folded_Diff_Op_Amp_Layout_0.VCD.n36 Folded_Diff_Op_Amp_Layout_0.VCD.n35 1.6385
R19919 Folded_Diff_Op_Amp_Layout_0.VCD.n34 Folded_Diff_Op_Amp_Layout_0.VCD.t11 1.6385
R19920 Folded_Diff_Op_Amp_Layout_0.VCD.n34 Folded_Diff_Op_Amp_Layout_0.VCD.n33 1.6385
R19921 Folded_Diff_Op_Amp_Layout_0.VCD.n50 Folded_Diff_Op_Amp_Layout_0.VCD.t12 1.6385
R19922 Folded_Diff_Op_Amp_Layout_0.VCD.n50 Folded_Diff_Op_Amp_Layout_0.VCD.n49 1.6385
R19923 Folded_Diff_Op_Amp_Layout_0.VCD.n45 Folded_Diff_Op_Amp_Layout_0.VCD.t53 1.6385
R19924 Folded_Diff_Op_Amp_Layout_0.VCD.n45 Folded_Diff_Op_Amp_Layout_0.VCD.n44 1.6385
R19925 Folded_Diff_Op_Amp_Layout_0.VCD.n43 Folded_Diff_Op_Amp_Layout_0.VCD.t6 1.6385
R19926 Folded_Diff_Op_Amp_Layout_0.VCD.n43 Folded_Diff_Op_Amp_Layout_0.VCD.n42 1.6385
R19927 Folded_Diff_Op_Amp_Layout_0.VCD.n179 Folded_Diff_Op_Amp_Layout_0.VCD.t63 1.6385
R19928 Folded_Diff_Op_Amp_Layout_0.VCD.n179 Folded_Diff_Op_Amp_Layout_0.VCD.n178 1.6385
R19929 Folded_Diff_Op_Amp_Layout_0.VCD.n181 Folded_Diff_Op_Amp_Layout_0.VCD.t45 1.6385
R19930 Folded_Diff_Op_Amp_Layout_0.VCD.n181 Folded_Diff_Op_Amp_Layout_0.VCD.n180 1.6385
R19931 Folded_Diff_Op_Amp_Layout_0.VCD.n183 Folded_Diff_Op_Amp_Layout_0.VCD.t46 1.6385
R19932 Folded_Diff_Op_Amp_Layout_0.VCD.n183 Folded_Diff_Op_Amp_Layout_0.VCD.n182 1.6385
R19933 Folded_Diff_Op_Amp_Layout_0.VCD.n173 Folded_Diff_Op_Amp_Layout_0.VCD.t8 1.6385
R19934 Folded_Diff_Op_Amp_Layout_0.VCD.n173 Folded_Diff_Op_Amp_Layout_0.VCD.n172 1.6385
R19935 Folded_Diff_Op_Amp_Layout_0.VCD.n171 Folded_Diff_Op_Amp_Layout_0.VCD.t36 1.6385
R19936 Folded_Diff_Op_Amp_Layout_0.VCD.n171 Folded_Diff_Op_Amp_Layout_0.VCD.n170 1.6385
R19937 Folded_Diff_Op_Amp_Layout_0.VCD.n73 Folded_Diff_Op_Amp_Layout_0.VCD.t14 1.6385
R19938 Folded_Diff_Op_Amp_Layout_0.VCD.n73 Folded_Diff_Op_Amp_Layout_0.VCD.n72 1.6385
R19939 Folded_Diff_Op_Amp_Layout_0.VCD.n113 Folded_Diff_Op_Amp_Layout_0.VCD.n112 1.49763
R19940 Folded_Diff_Op_Amp_Layout_0.VCD.n13 Folded_Diff_Op_Amp_Layout_0.VCD.n12 1.46669
R19941 Folded_Diff_Op_Amp_Layout_0.VCD.n22 Folded_Diff_Op_Amp_Layout_0.VCD.n21 1.46669
R19942 Folded_Diff_Op_Amp_Layout_0.VCD.n37 Folded_Diff_Op_Amp_Layout_0.VCD.n36 1.46669
R19943 Folded_Diff_Op_Amp_Layout_0.VCD.n46 Folded_Diff_Op_Amp_Layout_0.VCD.n45 1.46669
R19944 Folded_Diff_Op_Amp_Layout_0.VCD.n174 Folded_Diff_Op_Amp_Layout_0.VCD.n173 1.46669
R19945 Folded_Diff_Op_Amp_Layout_0.VCD.n156 Folded_Diff_Op_Amp_Layout_0.VCD.n155 1.46648
R19946 Folded_Diff_Op_Amp_Layout_0.VCD.n4 Folded_Diff_Op_Amp_Layout_0.VCD.n17 1.2862
R19947 Folded_Diff_Op_Amp_Layout_0.VCD.n75 Folded_Diff_Op_Amp_Layout_0.VCD.n74 1.18907
R19948 Folded_Diff_Op_Amp_Layout_0.VCD.n163 Folded_Diff_Op_Amp_Layout_0.VCD.n162 1.18861
R19949 Folded_Diff_Op_Amp_Layout_0.VCD.n113 Folded_Diff_Op_Amp_Layout_0.VCD.n84 1.1885
R19950 Folded_Diff_Op_Amp_Layout_0.VCD.n152 Folded_Diff_Op_Amp_Layout_0.VCD.n151 1.1885
R19951 Folded_Diff_Op_Amp_Layout_0.VCD.n120 Folded_Diff_Op_Amp_Layout_0.VCD.n119 1.18813
R19952 Folded_Diff_Op_Amp_Layout_0.VCD.n108 Folded_Diff_Op_Amp_Layout_0.VCD.n107 1.18813
R19953 Folded_Diff_Op_Amp_Layout_0.VCD.n89 Folded_Diff_Op_Amp_Layout_0.VCD.n88 1.18813
R19954 Folded_Diff_Op_Amp_Layout_0.VCD.n143 Folded_Diff_Op_Amp_Layout_0.VCD.n142 1.18813
R19955 Folded_Diff_Op_Amp_Layout_0.VCD.n127 Folded_Diff_Op_Amp_Layout_0.VCD.n126 1.18813
R19956 Folded_Diff_Op_Amp_Layout_0.VCD.n68 Folded_Diff_Op_Amp_Layout_0.VCD.n67 1.18665
R19957 Folded_Diff_Op_Amp_Layout_0.VCD.n58 Folded_Diff_Op_Amp_Layout_0.VCD.n57 1.18665
R19958 Folded_Diff_Op_Amp_Layout_0.VCD.n97 Folded_Diff_Op_Amp_Layout_0.VCD.n96 1.18665
R19959 Folded_Diff_Op_Amp_Layout_0.VCD.n135 Folded_Diff_Op_Amp_Layout_0.VCD.n134 1.18665
R19960 Folded_Diff_Op_Amp_Layout_0.VCD.n169 Folded_Diff_Op_Amp_Layout_0.VCD.n168 1.18665
R19961 Folded_Diff_Op_Amp_Layout_0.VCD.n17 Folded_Diff_Op_Amp_Layout_0.VCD.n8 1.18665
R19962 Folded_Diff_Op_Amp_Layout_0.VCD.n41 Folded_Diff_Op_Amp_Layout_0.VCD.n32 1.18665
R19963 Folded_Diff_Op_Amp_Layout_0.VCD.n28 Folded_Diff_Op_Amp_Layout_0.VCD.n27 1.18614
R19964 Folded_Diff_Op_Amp_Layout_0.VCD.n52 Folded_Diff_Op_Amp_Layout_0.VCD.n51 1.18614
R19965 Folded_Diff_Op_Amp_Layout_0.VCD.n1 Folded_Diff_Op_Amp_Layout_0.VCD.n41 1.12572
R19966 Folded_Diff_Op_Amp_Layout_0.VCD.n0 Folded_Diff_Op_Amp_Layout_0.VCD.n177 1.10736
R19967 Folded_Diff_Op_Amp_Layout_0.VCD.n148 Folded_Diff_Op_Amp_Layout_0.VCD.n130 1.06662
R19968 Folded_Diff_Op_Amp_Layout_0.VCD.n185 Folded_Diff_Op_Amp_Layout_0.VCD.n184 1.02906
R19969 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VCD.n186 1.01399
R19970 Folded_Diff_Op_Amp_Layout_0.VCD.n185 Folded_Diff_Op_Amp_Layout_0.VCD.n179 0.927451
R19971 Folded_Diff_Op_Amp_Layout_0.VCD.n67 Folded_Diff_Op_Amp_Layout_0.VCD.n66 0.901687
R19972 Folded_Diff_Op_Amp_Layout_0.VCD.n57 Folded_Diff_Op_Amp_Layout_0.VCD.n56 0.901687
R19973 Folded_Diff_Op_Amp_Layout_0.VCD.n96 Folded_Diff_Op_Amp_Layout_0.VCD.n95 0.901687
R19974 Folded_Diff_Op_Amp_Layout_0.VCD.n162 Folded_Diff_Op_Amp_Layout_0.VCD.n161 0.901687
R19975 Folded_Diff_Op_Amp_Layout_0.VCD.n134 Folded_Diff_Op_Amp_Layout_0.VCD.n133 0.901687
R19976 Folded_Diff_Op_Amp_Layout_0.VCD.n168 Folded_Diff_Op_Amp_Layout_0.VCD.n167 0.901687
R19977 Folded_Diff_Op_Amp_Layout_0.VCD.n8 Folded_Diff_Op_Amp_Layout_0.VCD.n7 0.901687
R19978 Folded_Diff_Op_Amp_Layout_0.VCD.n32 Folded_Diff_Op_Amp_Layout_0.VCD.n31 0.901687
R19979 Folded_Diff_Op_Amp_Layout_0.VCD.n84 Folded_Diff_Op_Amp_Layout_0.VCD.n83 0.90147
R19980 Folded_Diff_Op_Amp_Layout_0.VCD.n151 Folded_Diff_Op_Amp_Layout_0.VCD.n150 0.90147
R19981 Folded_Diff_Op_Amp_Layout_0.VCD.n119 Folded_Diff_Op_Amp_Layout_0.VCD.n118 0.90147
R19982 Folded_Diff_Op_Amp_Layout_0.VCD.n107 Folded_Diff_Op_Amp_Layout_0.VCD.n106 0.90147
R19983 Folded_Diff_Op_Amp_Layout_0.VCD.n88 Folded_Diff_Op_Amp_Layout_0.VCD.n87 0.90147
R19984 Folded_Diff_Op_Amp_Layout_0.VCD.n142 Folded_Diff_Op_Amp_Layout_0.VCD.n141 0.90147
R19985 Folded_Diff_Op_Amp_Layout_0.VCD.n126 Folded_Diff_Op_Amp_Layout_0.VCD.n125 0.90147
R19986 Folded_Diff_Op_Amp_Layout_0.VCD.n27 Folded_Diff_Op_Amp_Layout_0.VCD.n26 0.90147
R19987 Folded_Diff_Op_Amp_Layout_0.VCD.n51 Folded_Diff_Op_Amp_Layout_0.VCD.n50 0.90147
R19988 Folded_Diff_Op_Amp_Layout_0.VCD.n74 Folded_Diff_Op_Amp_Layout_0.VCD.n73 0.901426
R19989 Folded_Diff_Op_Amp_Layout_0.VCD.n70 Folded_Diff_Op_Amp_Layout_0.VCD.n69 0.743266
R19990 Folded_Diff_Op_Amp_Layout_0.VCD.n100 Folded_Diff_Op_Amp_Layout_0.VCD.n98 0.727104
R19991 Folded_Diff_Op_Amp_Layout_0.VCD.n138 Folded_Diff_Op_Amp_Layout_0.VCD.n136 0.727104
R19992 Folded_Diff_Op_Amp_Layout_0.VCD.n61 Folded_Diff_Op_Amp_Layout_0.VCD.n59 0.727104
R19993 Folded_Diff_Op_Amp_Layout_0.VCD.n3 Folded_Diff_Op_Amp_Layout_0.VCD.n53 0.722779
R19994 Folded_Diff_Op_Amp_Layout_0.VCD.n5 Folded_Diff_Op_Amp_Layout_0.VCD.n29 0.722779
R19995 Folded_Diff_Op_Amp_Layout_0.VCD.n157 Folded_Diff_Op_Amp_Layout_0.VCD.n156 0.70619
R19996 Folded_Diff_Op_Amp_Layout_0.VCD.n14 Folded_Diff_Op_Amp_Layout_0.VCD.n13 0.693301
R19997 Folded_Diff_Op_Amp_Layout_0.VCD.n38 Folded_Diff_Op_Amp_Layout_0.VCD.n37 0.693301
R19998 Folded_Diff_Op_Amp_Layout_0.VCD.n156 Folded_Diff_Op_Amp_Layout_0.VCD.n153 0.689663
R19999 Folded_Diff_Op_Amp_Layout_0.VCD.n23 Folded_Diff_Op_Amp_Layout_0.VCD.n22 0.676871
R20000 Folded_Diff_Op_Amp_Layout_0.VCD.n47 Folded_Diff_Op_Amp_Layout_0.VCD.n46 0.676871
R20001 Folded_Diff_Op_Amp_Layout_0.VCD.n175 Folded_Diff_Op_Amp_Layout_0.VCD.n174 0.676871
R20002 Folded_Diff_Op_Amp_Layout_0.VCD.n110 Folded_Diff_Op_Amp_Layout_0.VCD.n109 0.631966
R20003 Folded_Diff_Op_Amp_Layout_0.VCD.n145 Folded_Diff_Op_Amp_Layout_0.VCD.n144 0.631966
R20004 Folded_Diff_Op_Amp_Layout_0.VCD.n63 Folded_Diff_Op_Amp_Layout_0.VCD.n76 0.616779
R20005 Folded_Diff_Op_Amp_Layout_0.VCD.n92 Folded_Diff_Op_Amp_Layout_0.VCD.n90 0.616779
R20006 Folded_Diff_Op_Amp_Layout_0.VCD.n122 Folded_Diff_Op_Amp_Layout_0.VCD.n121 0.616779
R20007 Folded_Diff_Op_Amp_Layout_0.VCD.n130 Folded_Diff_Op_Amp_Layout_0.VCD.n128 0.616779
R20008 Folded_Diff_Op_Amp_Layout_0.VCD.n115 Folded_Diff_Op_Amp_Layout_0.VCD.n114 0.598695
R20009 Folded_Diff_Op_Amp_Layout_0.VCD.n165 Folded_Diff_Op_Amp_Layout_0.VCD.n164 0.598695
R20010 Folded_Diff_Op_Amp_Layout_0.VCD.n186 Folded_Diff_Op_Amp_Layout_0.VCD.n0 0.499954
R20011 Folded_Diff_Op_Amp_Layout_0.VCD.n0 Folded_Diff_Op_Amp_Layout_0.VCD.n3 0.195441
R20012 Folded_Diff_Op_Amp_Layout_0.VCD.n112 Folded_Diff_Op_Amp_Layout_0.VCD.n92 0.187017
R20013 Folded_Diff_Op_Amp_Layout_0.VCD.n1 Folded_Diff_Op_Amp_Layout_0.VCD.n5 0.183654
R20014 Folded_Diff_Op_Amp_Layout_0.VCD.n2 Folded_Diff_Op_Amp_Layout_0.VCD.n1 0.160979
R20015 Folded_Diff_Op_Amp_Layout_0.VCD.n99 Folded_Diff_Op_Amp_Layout_0.VCD.n110 0.150125
R20016 Folded_Diff_Op_Amp_Layout_0.VCD.n91 Folded_Diff_Op_Amp_Layout_0.VCD.n111 0.150125
R20017 Folded_Diff_Op_Amp_Layout_0.VCD.n137 Folded_Diff_Op_Amp_Layout_0.VCD.n145 0.150125
R20018 Folded_Diff_Op_Amp_Layout_0.VCD.n129 Folded_Diff_Op_Amp_Layout_0.VCD.n146 0.150125
R20019 Folded_Diff_Op_Amp_Layout_0.VCD.n62 Folded_Diff_Op_Amp_Layout_0.VCD.n70 0.150125
R20020 Folded_Diff_Op_Amp_Layout_0.VCD.n60 Folded_Diff_Op_Amp_Layout_0.VCD.n77 0.150125
R20021 Folded_Diff_Op_Amp_Layout_0.VCD.n79 Folded_Diff_Op_Amp_Layout_0.VCD.n78 0.150125
R20022 Folded_Diff_Op_Amp_Layout_0.VCD.n152 Folded_Diff_Op_Amp_Layout_0.VCD.n148 0.0995747
R20023 Folded_Diff_Op_Amp_Layout_0.VCD.n177 Folded_Diff_Op_Amp_Layout_0.VCD.n176 0.0929251
R20024 Folded_Diff_Op_Amp_Layout_0.VCD.n17 Folded_Diff_Op_Amp_Layout_0.VCD.n16 0.0832399
R20025 Folded_Diff_Op_Amp_Layout_0.VCD.n41 Folded_Diff_Op_Amp_Layout_0.VCD.n40 0.0832399
R20026 Folded_Diff_Op_Amp_Layout_0.VCD.n113 Folded_Diff_Op_Amp_Layout_0.VCD.n81 0.0831446
R20027 Folded_Diff_Op_Amp_Layout_0.VCD.n69 Folded_Diff_Op_Amp_Layout_0.VCD.n64 0.0823987
R20028 Folded_Diff_Op_Amp_Layout_0.VCD.n59 Folded_Diff_Op_Amp_Layout_0.VCD.n54 0.0823987
R20029 Folded_Diff_Op_Amp_Layout_0.VCD.n98 Folded_Diff_Op_Amp_Layout_0.VCD.n93 0.0823987
R20030 Folded_Diff_Op_Amp_Layout_0.VCD.n136 Folded_Diff_Op_Amp_Layout_0.VCD.n131 0.0823987
R20031 Folded_Diff_Op_Amp_Layout_0.VCD.n159 Folded_Diff_Op_Amp_Layout_0.VCD.n158 0.0754039
R20032 Folded_Diff_Op_Amp_Layout_0.VCD.n90 Folded_Diff_Op_Amp_Layout_0.VCD.n85 0.0712285
R20033 Folded_Diff_Op_Amp_Layout_0.VCD.n109 Folded_Diff_Op_Amp_Layout_0.VCD.n104 0.0712285
R20034 Folded_Diff_Op_Amp_Layout_0.VCD.n128 Folded_Diff_Op_Amp_Layout_0.VCD.n123 0.0712285
R20035 Folded_Diff_Op_Amp_Layout_0.VCD.n144 Folded_Diff_Op_Amp_Layout_0.VCD.n139 0.0712285
R20036 Folded_Diff_Op_Amp_Layout_0.VCD.n121 Folded_Diff_Op_Amp_Layout_0.VCD.n116 0.0712285
R20037 Folded_Diff_Op_Amp_Layout_0.VCD.n76 Folded_Diff_Op_Amp_Layout_0.VCD.n71 0.0712285
R20038 Folded_Diff_Op_Amp_Layout_0.VCD.n53 Folded_Diff_Op_Amp_Layout_0.VCD.n52 0.0623678
R20039 Folded_Diff_Op_Amp_Layout_0.VCD.n29 Folded_Diff_Op_Amp_Layout_0.VCD.n28 0.0623678
R20040 Folded_Diff_Op_Amp_Layout_0.VCD.n29 Folded_Diff_Op_Amp_Layout_0.VCD.n24 0.0620327
R20041 Folded_Diff_Op_Amp_Layout_0.VCD.n53 Folded_Diff_Op_Amp_Layout_0.VCD.n48 0.0620327
R20042 Folded_Diff_Op_Amp_Layout_0.VCD.n109 Folded_Diff_Op_Amp_Layout_0.VCD.n108 0.0534597
R20043 Folded_Diff_Op_Amp_Layout_0.VCD.n90 Folded_Diff_Op_Amp_Layout_0.VCD.n89 0.0534597
R20044 Folded_Diff_Op_Amp_Layout_0.VCD.n144 Folded_Diff_Op_Amp_Layout_0.VCD.n143 0.0534597
R20045 Folded_Diff_Op_Amp_Layout_0.VCD.n128 Folded_Diff_Op_Amp_Layout_0.VCD.n127 0.0534597
R20046 Folded_Diff_Op_Amp_Layout_0.VCD.n121 Folded_Diff_Op_Amp_Layout_0.VCD.n120 0.0534597
R20047 Folded_Diff_Op_Amp_Layout_0.VCD.n76 Folded_Diff_Op_Amp_Layout_0.VCD.n75 0.0534597
R20048 Folded_Diff_Op_Amp_Layout_0.VCD.n163 Folded_Diff_Op_Amp_Layout_0.VCD.n159 0.0500104
R20049 Folded_Diff_Op_Amp_Layout_0.VCD.n81 Folded_Diff_Op_Amp_Layout_0.VCD.n80 0.0420655
R20050 Folded_Diff_Op_Amp_Layout_0.VCD.n16 Folded_Diff_Op_Amp_Layout_0.VCD.n15 0.0419676
R20051 Folded_Diff_Op_Amp_Layout_0.VCD.n40 Folded_Diff_Op_Amp_Layout_0.VCD.n39 0.0419676
R20052 Folded_Diff_Op_Amp_Layout_0.VCD.n98 Folded_Diff_Op_Amp_Layout_0.VCD.n97 0.0415773
R20053 Folded_Diff_Op_Amp_Layout_0.VCD.n136 Folded_Diff_Op_Amp_Layout_0.VCD.n135 0.0415773
R20054 Folded_Diff_Op_Amp_Layout_0.VCD.n59 Folded_Diff_Op_Amp_Layout_0.VCD.n58 0.0415773
R20055 Folded_Diff_Op_Amp_Layout_0.VCD.n69 Folded_Diff_Op_Amp_Layout_0.VCD.n68 0.0415773
R20056 Folded_Diff_Op_Amp_Layout_0.VCD.n104 Folded_Diff_Op_Amp_Layout_0.VCD.n103 0.0324737
R20057 Folded_Diff_Op_Amp_Layout_0.VCD.n114 Folded_Diff_Op_Amp_Layout_0.VCD.n113 0.0324737
R20058 Folded_Diff_Op_Amp_Layout_0.VCD.n116 Folded_Diff_Op_Amp_Layout_0.VCD.n115 0.0324737
R20059 Folded_Diff_Op_Amp_Layout_0.VCD.n153 Folded_Diff_Op_Amp_Layout_0.VCD.n152 0.0324737
R20060 Folded_Diff_Op_Amp_Layout_0.VCD.n24 Folded_Diff_Op_Amp_Layout_0.VCD.n23 0.0324737
R20061 Folded_Diff_Op_Amp_Layout_0.VCD.n48 Folded_Diff_Op_Amp_Layout_0.VCD.n47 0.0324737
R20062 Folded_Diff_Op_Amp_Layout_0.VCD.n169 Folded_Diff_Op_Amp_Layout_0.VCD.n165 0.0324737
R20063 Folded_Diff_Op_Amp_Layout_0.VCD.n176 Folded_Diff_Op_Amp_Layout_0.VCD.n175 0.0324737
R20064 Folded_Diff_Op_Amp_Layout_0.VCD.n164 Folded_Diff_Op_Amp_Layout_0.VCD.n163 0.0324737
R20065 Folded_Diff_Op_Amp_Layout_0.VCD.n177 Folded_Diff_Op_Amp_Layout_0.VCD.n169 0.0320039
R20066 Folded_Diff_Op_Amp_Layout_0.VCD.n148 Folded_Diff_Op_Amp_Layout_0.VCD.n147 0.0261793
R20067 Folded_Diff_Op_Amp_Layout_0.VCD.n39 Folded_Diff_Op_Amp_Layout_0.VCD.n38 0.0169302
R20068 Folded_Diff_Op_Amp_Layout_0.VCD.n15 Folded_Diff_Op_Amp_Layout_0.VCD.n14 0.0169302
R20069 Folded_Diff_Op_Amp_Layout_0.VCD.n158 Folded_Diff_Op_Amp_Layout_0.VCD.n157 0.0169302
R20070 Folded_Diff_Op_Amp_Layout_0.VCD.n63 Folded_Diff_Op_Amp_Layout_0.VCD.n62 0.016662
R20071 Folded_Diff_Op_Amp_Layout_0.VCD.n78 Folded_Diff_Op_Amp_Layout_0.VCD.n61 0.016662
R20072 Folded_Diff_Op_Amp_Layout_0.VCD.n111 Folded_Diff_Op_Amp_Layout_0.VCD.n100 0.016662
R20073 Folded_Diff_Op_Amp_Layout_0.VCD.n92 Folded_Diff_Op_Amp_Layout_0.VCD.n91 0.016662
R20074 Folded_Diff_Op_Amp_Layout_0.VCD.n146 Folded_Diff_Op_Amp_Layout_0.VCD.n138 0.016662
R20075 Folded_Diff_Op_Amp_Layout_0.VCD.n130 Folded_Diff_Op_Amp_Layout_0.VCD.n129 0.016662
R20076 Folded_Diff_Op_Amp_Layout_0.VCD.n61 Folded_Diff_Op_Amp_Layout_0.VCD.n60 0.0166619
R20077 Folded_Diff_Op_Amp_Layout_0.VCD.n100 Folded_Diff_Op_Amp_Layout_0.VCD.n99 0.0166619
R20078 Folded_Diff_Op_Amp_Layout_0.VCD.n138 Folded_Diff_Op_Amp_Layout_0.VCD.n137 0.0166619
R20079 Folded_Diff_Op_Amp_Layout_0.VCD.n5 Folded_Diff_Op_Amp_Layout_0.VCD.n4 0.016568
R20080 Folded_Diff_Op_Amp_Layout_0.VCD.n3 Folded_Diff_Op_Amp_Layout_0.VCD.n2 0.016568
R20081 Folded_Diff_Op_Amp_Layout_0.VCD.n77 Folded_Diff_Op_Amp_Layout_0.VCD.n63 0.0156875
R20082 Folded_Diff_Op_Amp_Layout_0.VCD.n122 Folded_Diff_Op_Amp_Layout_0.VCD.n79 0.0156875
R20083 Folded_Diff_Op_Amp_Layout_0.VCD.n159 Folded_Diff_Op_Amp_Layout_0.VCD.n122 1.05492
R20084 Folded_Diff_Op_Amp_Layout_0.VB1.n55 Folded_Diff_Op_Amp_Layout_0.VB1.t30 63.68
R20085 Folded_Diff_Op_Amp_Layout_0.VB1.n55 Folded_Diff_Op_Amp_Layout_0.VB1.t32 63.68
R20086 Folded_Diff_Op_Amp_Layout_0.VB1.n7 Folded_Diff_Op_Amp_Layout_0.VB1.t43 61.7898
R20087 Folded_Diff_Op_Amp_Layout_0.VB1.n10 Folded_Diff_Op_Amp_Layout_0.VB1.t42 61.7898
R20088 Folded_Diff_Op_Amp_Layout_0.VB1.n11 Folded_Diff_Op_Amp_Layout_0.VB1.t48 61.7898
R20089 Folded_Diff_Op_Amp_Layout_0.VB1.n12 Folded_Diff_Op_Amp_Layout_0.VB1.t35 61.7898
R20090 Folded_Diff_Op_Amp_Layout_0.VB1.n9 Folded_Diff_Op_Amp_Layout_0.VB1.t45 61.7898
R20091 Folded_Diff_Op_Amp_Layout_0.VB1.n5 Folded_Diff_Op_Amp_Layout_0.VB1.t63 61.7898
R20092 Folded_Diff_Op_Amp_Layout_0.VB1.n6 Folded_Diff_Op_Amp_Layout_0.VB1.t39 61.7898
R20093 Folded_Diff_Op_Amp_Layout_0.VB1.n8 Folded_Diff_Op_Amp_Layout_0.VB1.t60 61.7898
R20094 Folded_Diff_Op_Amp_Layout_0.VB1.n21 Folded_Diff_Op_Amp_Layout_0.VB1.t52 61.5291
R20095 Folded_Diff_Op_Amp_Layout_0.VB1.n22 Folded_Diff_Op_Amp_Layout_0.VB1.t62 61.5291
R20096 Folded_Diff_Op_Amp_Layout_0.VB1.n23 Folded_Diff_Op_Amp_Layout_0.VB1.t65 61.5291
R20097 Folded_Diff_Op_Amp_Layout_0.VB1.n24 Folded_Diff_Op_Amp_Layout_0.VB1.t61 61.5291
R20098 Folded_Diff_Op_Amp_Layout_0.VB1.n25 Folded_Diff_Op_Amp_Layout_0.VB1.t64 61.5291
R20099 Folded_Diff_Op_Amp_Layout_0.VB1.n26 Folded_Diff_Op_Amp_Layout_0.VB1.t41 61.5291
R20100 Folded_Diff_Op_Amp_Layout_0.VB1.n27 Folded_Diff_Op_Amp_Layout_0.VB1.t49 61.5291
R20101 Folded_Diff_Op_Amp_Layout_0.VB1.n13 Folded_Diff_Op_Amp_Layout_0.VB1.t55 60.6166
R20102 Folded_Diff_Op_Amp_Layout_0.VB1.n14 Folded_Diff_Op_Amp_Layout_0.VB1.t36 60.6166
R20103 Folded_Diff_Op_Amp_Layout_0.VB1.n15 Folded_Diff_Op_Amp_Layout_0.VB1.t38 60.6166
R20104 Folded_Diff_Op_Amp_Layout_0.VB1.n16 Folded_Diff_Op_Amp_Layout_0.VB1.t34 60.6166
R20105 Folded_Diff_Op_Amp_Layout_0.VB1.n17 Folded_Diff_Op_Amp_Layout_0.VB1.t37 60.6166
R20106 Folded_Diff_Op_Amp_Layout_0.VB1.n18 Folded_Diff_Op_Amp_Layout_0.VB1.t44 60.6166
R20107 Folded_Diff_Op_Amp_Layout_0.VB1.n20 Folded_Diff_Op_Amp_Layout_0.VB1.t54 60.6166
R20108 Folded_Diff_Op_Amp_Layout_0.VB1.n19 Folded_Diff_Op_Amp_Layout_0.VB1.t53 60.6166
R20109 Folded_Diff_Op_Amp_Layout_0.VB1.t51 Folded_Diff_Op_Amp_Layout_0.VB1.n20 58.7916
R20110 Folded_Diff_Op_Amp_Layout_0.VB1.n21 Folded_Diff_Op_Amp_Layout_0.VB1.t50 57.8791
R20111 Folded_Diff_Op_Amp_Layout_0.VB1.n22 Folded_Diff_Op_Amp_Layout_0.VB1.t57 57.8791
R20112 Folded_Diff_Op_Amp_Layout_0.VB1.n23 Folded_Diff_Op_Amp_Layout_0.VB1.t59 57.8791
R20113 Folded_Diff_Op_Amp_Layout_0.VB1.n24 Folded_Diff_Op_Amp_Layout_0.VB1.t56 57.8791
R20114 Folded_Diff_Op_Amp_Layout_0.VB1.n25 Folded_Diff_Op_Amp_Layout_0.VB1.t58 57.8791
R20115 Folded_Diff_Op_Amp_Layout_0.VB1.n26 Folded_Diff_Op_Amp_Layout_0.VB1.t40 57.8791
R20116 Folded_Diff_Op_Amp_Layout_0.VB1.n27 Folded_Diff_Op_Amp_Layout_0.VB1.t46 57.8791
R20117 Folded_Diff_Op_Amp_Layout_0.VB1.n28 Folded_Diff_Op_Amp_Layout_0.VB1.t47 57.8791
R20118 Folded_Diff_Op_Amp_Layout_0.VB1.t38 Folded_Diff_Op_Amp_Layout_0.VB1.n12 57.6184
R20119 Folded_Diff_Op_Amp_Layout_0.VB1.t34 Folded_Diff_Op_Amp_Layout_0.VB1.n9 57.6184
R20120 Folded_Diff_Op_Amp_Layout_0.VB1.t54 Folded_Diff_Op_Amp_Layout_0.VB1.n8 57.6184
R20121 Folded_Diff_Op_Amp_Layout_0.VB1.n30 Folded_Diff_Op_Amp_Layout_0.VB1.t51 56.0585
R20122 Folded_Diff_Op_Amp_Layout_0.VB1.n11 Folded_Diff_Op_Amp_Layout_0.VB1.n10 9.73383
R20123 Folded_Diff_Op_Amp_Layout_0.VB1.n12 Folded_Diff_Op_Amp_Layout_0.VB1.n11 9.73383
R20124 Folded_Diff_Op_Amp_Layout_0.VB1.n6 Folded_Diff_Op_Amp_Layout_0.VB1.n5 9.73383
R20125 Folded_Diff_Op_Amp_Layout_0.VB1.n7 Folded_Diff_Op_Amp_Layout_0.VB1.n6 9.73383
R20126 Folded_Diff_Op_Amp_Layout_0.VB1.n8 Folded_Diff_Op_Amp_Layout_0.VB1.n7 9.73383
R20127 Folded_Diff_Op_Amp_Layout_0.VB1.n14 Folded_Diff_Op_Amp_Layout_0.VB1.n13 9.73383
R20128 Folded_Diff_Op_Amp_Layout_0.VB1.n15 Folded_Diff_Op_Amp_Layout_0.VB1.n14 9.73383
R20129 Folded_Diff_Op_Amp_Layout_0.VB1.n16 Folded_Diff_Op_Amp_Layout_0.VB1.n15 9.73383
R20130 Folded_Diff_Op_Amp_Layout_0.VB1.n17 Folded_Diff_Op_Amp_Layout_0.VB1.n16 9.73383
R20131 Folded_Diff_Op_Amp_Layout_0.VB1.n18 Folded_Diff_Op_Amp_Layout_0.VB1.n17 9.73383
R20132 Folded_Diff_Op_Amp_Layout_0.VB1.n19 Folded_Diff_Op_Amp_Layout_0.VB1.n18 9.73383
R20133 Folded_Diff_Op_Amp_Layout_0.VB1.n20 Folded_Diff_Op_Amp_Layout_0.VB1.n19 9.73383
R20134 Folded_Diff_Op_Amp_Layout_0.VB1.n22 Folded_Diff_Op_Amp_Layout_0.VB1.n21 9.73383
R20135 Folded_Diff_Op_Amp_Layout_0.VB1.n23 Folded_Diff_Op_Amp_Layout_0.VB1.n22 9.73383
R20136 Folded_Diff_Op_Amp_Layout_0.VB1.n24 Folded_Diff_Op_Amp_Layout_0.VB1.n23 9.73383
R20137 Folded_Diff_Op_Amp_Layout_0.VB1.n25 Folded_Diff_Op_Amp_Layout_0.VB1.n24 9.73383
R20138 Folded_Diff_Op_Amp_Layout_0.VB1.n26 Folded_Diff_Op_Amp_Layout_0.VB1.n25 9.73383
R20139 Folded_Diff_Op_Amp_Layout_0.VB1.n27 Folded_Diff_Op_Amp_Layout_0.VB1.n26 9.73383
R20140 Folded_Diff_Op_Amp_Layout_0.VB1.n28 Folded_Diff_Op_Amp_Layout_0.VB1.n27 9.73383
R20141 Folded_Diff_Op_Amp_Layout_0.VB1.n43 Folded_Diff_Op_Amp_Layout_0.VB1.t13 6.32241
R20142 Folded_Diff_Op_Amp_Layout_0.VB1.n40 Folded_Diff_Op_Amp_Layout_0.VB1.n39 6.32241
R20143 Folded_Diff_Op_Amp_Layout_0.VB1.n63 Folded_Diff_Op_Amp_Layout_0.VB1.t6 6.32241
R20144 Folded_Diff_Op_Amp_Layout_0.VB1.n60 Folded_Diff_Op_Amp_Layout_0.VB1.n59 6.32241
R20145 Folded_Diff_Op_Amp_Layout_0.VB1.n80 Folded_Diff_Op_Amp_Layout_0.VB1.t20 6.32241
R20146 Folded_Diff_Op_Amp_Layout_0.VB1.n77 Folded_Diff_Op_Amp_Layout_0.VB1.n76 6.32241
R20147 Folded_Diff_Op_Amp_Layout_0.VB1.n71 Folded_Diff_Op_Amp_Layout_0.VB1.n56 5.64446
R20148 Folded_Diff_Op_Amp_Layout_0.VB1.n56 Folded_Diff_Op_Amp_Layout_0.VB1.n55 5.14084
R20149 Folded_Diff_Op_Amp_Layout_0.VB1.n47 Folded_Diff_Op_Amp_Layout_0.VB1.n46 4.39485
R20150 Folded_Diff_Op_Amp_Layout_0.VB1.n67 Folded_Diff_Op_Amp_Layout_0.VB1.n66 4.36159
R20151 Folded_Diff_Op_Amp_Layout_0.VB1.n84 Folded_Diff_Op_Amp_Layout_0.VB1.n83 4.36159
R20152 Folded_Diff_Op_Amp_Layout_0.VB1.n43 Folded_Diff_Op_Amp_Layout_0.VB1.n42 3.43224
R20153 Folded_Diff_Op_Amp_Layout_0.VB1.n40 Folded_Diff_Op_Amp_Layout_0.VB1.n38 3.43224
R20154 Folded_Diff_Op_Amp_Layout_0.VB1.n63 Folded_Diff_Op_Amp_Layout_0.VB1.n62 3.43224
R20155 Folded_Diff_Op_Amp_Layout_0.VB1.n60 Folded_Diff_Op_Amp_Layout_0.VB1.n58 3.43224
R20156 Folded_Diff_Op_Amp_Layout_0.VB1.n80 Folded_Diff_Op_Amp_Layout_0.VB1.n79 3.43224
R20157 Folded_Diff_Op_Amp_Layout_0.VB1.n77 Folded_Diff_Op_Amp_Layout_0.VB1.n75 3.43224
R20158 Folded_Diff_Op_Amp_Layout_0.VB1.n36 Folded_Diff_Op_Amp_Layout_0.VB1.n99 3.1965
R20159 Folded_Diff_Op_Amp_Layout_0.VB1.n34 Folded_Diff_Op_Amp_Layout_0.VB1.n30 2.8805
R20160 Folded_Diff_Op_Amp_Layout_0.VB1.n29 Folded_Diff_Op_Amp_Layout_0.VB1.n28 1.88633
R20161 Folded_Diff_Op_Amp_Layout_0.VB1.n95 Folded_Diff_Op_Amp_Layout_0.VB1.t21 1.6385
R20162 Folded_Diff_Op_Amp_Layout_0.VB1.n95 Folded_Diff_Op_Amp_Layout_0.VB1.n94 1.6385
R20163 Folded_Diff_Op_Amp_Layout_0.VB1.n46 Folded_Diff_Op_Amp_Layout_0.VB1.t24 1.6385
R20164 Folded_Diff_Op_Amp_Layout_0.VB1.n46 Folded_Diff_Op_Amp_Layout_0.VB1.n45 1.6385
R20165 Folded_Diff_Op_Amp_Layout_0.VB1.n42 Folded_Diff_Op_Amp_Layout_0.VB1.t22 1.6385
R20166 Folded_Diff_Op_Amp_Layout_0.VB1.n42 Folded_Diff_Op_Amp_Layout_0.VB1.n41 1.6385
R20167 Folded_Diff_Op_Amp_Layout_0.VB1.n38 Folded_Diff_Op_Amp_Layout_0.VB1.t8 1.6385
R20168 Folded_Diff_Op_Amp_Layout_0.VB1.n38 Folded_Diff_Op_Amp_Layout_0.VB1.n37 1.6385
R20169 Folded_Diff_Op_Amp_Layout_0.VB1.n51 Folded_Diff_Op_Amp_Layout_0.VB1.t5 1.6385
R20170 Folded_Diff_Op_Amp_Layout_0.VB1.n51 Folded_Diff_Op_Amp_Layout_0.VB1.n50 1.6385
R20171 Folded_Diff_Op_Amp_Layout_0.VB1.n66 Folded_Diff_Op_Amp_Layout_0.VB1.t11 1.6385
R20172 Folded_Diff_Op_Amp_Layout_0.VB1.n66 Folded_Diff_Op_Amp_Layout_0.VB1.n65 1.6385
R20173 Folded_Diff_Op_Amp_Layout_0.VB1.n62 Folded_Diff_Op_Amp_Layout_0.VB1.t15 1.6385
R20174 Folded_Diff_Op_Amp_Layout_0.VB1.n62 Folded_Diff_Op_Amp_Layout_0.VB1.n61 1.6385
R20175 Folded_Diff_Op_Amp_Layout_0.VB1.n58 Folded_Diff_Op_Amp_Layout_0.VB1.t3 1.6385
R20176 Folded_Diff_Op_Amp_Layout_0.VB1.n58 Folded_Diff_Op_Amp_Layout_0.VB1.n57 1.6385
R20177 Folded_Diff_Op_Amp_Layout_0.VB1.n83 Folded_Diff_Op_Amp_Layout_0.VB1.t1 1.6385
R20178 Folded_Diff_Op_Amp_Layout_0.VB1.n83 Folded_Diff_Op_Amp_Layout_0.VB1.n82 1.6385
R20179 Folded_Diff_Op_Amp_Layout_0.VB1.n79 Folded_Diff_Op_Amp_Layout_0.VB1.t0 1.6385
R20180 Folded_Diff_Op_Amp_Layout_0.VB1.n79 Folded_Diff_Op_Amp_Layout_0.VB1.n78 1.6385
R20181 Folded_Diff_Op_Amp_Layout_0.VB1.n75 Folded_Diff_Op_Amp_Layout_0.VB1.t16 1.6385
R20182 Folded_Diff_Op_Amp_Layout_0.VB1.n75 Folded_Diff_Op_Amp_Layout_0.VB1.n74 1.6385
R20183 Folded_Diff_Op_Amp_Layout_0.VB1.n89 Folded_Diff_Op_Amp_Layout_0.VB1.t26 1.6385
R20184 Folded_Diff_Op_Amp_Layout_0.VB1.n89 Folded_Diff_Op_Amp_Layout_0.VB1.n88 1.6385
R20185 Folded_Diff_Op_Amp_Layout_0.VB1.n3 Folded_Diff_Op_Amp_Layout_0.VB1.n93 1.50118
R20186 Folded_Diff_Op_Amp_Layout_0.VB1.n2 Folded_Diff_Op_Amp_Layout_0.VB1.n36 1.51249
R20187 Folded_Diff_Op_Amp_Layout_0.VB1.n92 Folded_Diff_Op_Amp_Layout_0.VB1.n91 1.49167
R20188 Folded_Diff_Op_Amp_Layout_0.VB1.n87 Folded_Diff_Op_Amp_Layout_0.VB1.n73 1.49167
R20189 Folded_Diff_Op_Amp_Layout_0.VB1.n3 Folded_Diff_Op_Amp_Layout_0.VB1.n98 1.48107
R20190 Folded_Diff_Op_Amp_Layout_0.VB1.n52 Folded_Diff_Op_Amp_Layout_0.VB1.n51 1.42054
R20191 Folded_Diff_Op_Amp_Layout_0.VB1.n96 Folded_Diff_Op_Amp_Layout_0.VB1.n95 1.42034
R20192 Folded_Diff_Op_Amp_Layout_0.VB1.n30 Folded_Diff_Op_Amp_Layout_0.VB1.n29 1.36152
R20193 Folded_Diff_Op_Amp_Layout_0.VB1.n91 Folded_Diff_Op_Amp_Layout_0.VB1.n90 1.17538
R20194 Folded_Diff_Op_Amp_Layout_0.VB1.n72 Folded_Diff_Op_Amp_Layout_0.VB1.n52 1.15277
R20195 Folded_Diff_Op_Amp_Layout_0.VB1.n97 Folded_Diff_Op_Amp_Layout_0.VB1.n96 1.15212
R20196 Folded_Diff_Op_Amp_Layout_0.VB1.n100 Folded_Diff_Op_Amp_Layout_0.VB1.n2 1.12725
R20197 Folded_Diff_Op_Amp_Layout_0.VB1.n100 Folded_Diff_Op_Amp_Layout_0.VB1.n0 1.12594
R20198 Folded_Diff_Op_Amp_Layout_0.VB1.n93 Folded_Diff_Op_Amp_Layout_0.VB1.n49 1.1255
R20199 Folded_Diff_Op_Amp_Layout_0.VB1.n70 Folded_Diff_Op_Amp_Layout_0.VB1.n69 1.1255
R20200 Folded_Diff_Op_Amp_Layout_0.VB1.n87 Folded_Diff_Op_Amp_Layout_0.VB1.n86 1.1255
R20201 Folded_Diff_Op_Amp_Layout_0.VB1.n68 Folded_Diff_Op_Amp_Layout_0.VB1.n67 1.07272
R20202 Folded_Diff_Op_Amp_Layout_0.VB1.n90 Folded_Diff_Op_Amp_Layout_0.VB1.n89 1.06259
R20203 Folded_Diff_Op_Amp_Layout_0.VB1.n85 Folded_Diff_Op_Amp_Layout_0.VB1.n84 1.05362
R20204 Folded_Diff_Op_Amp_Layout_0.VB1.n48 Folded_Diff_Op_Amp_Layout_0.VB1.n47 1.03946
R20205 Folded_Diff_Op_Amp_Layout_0.VB1.n4 Folded_Diff_Op_Amp_Layout_0.VB1.n34 4.74119
R20206 Folded_Diff_Op_Amp_Layout_0.VB1.n56 Folded_Diff_Op_Amp_Layout_0.VB1.n54 0.715901
R20207 Folded_Diff_Op_Amp_Layout_0.VB1.n54 Folded_Diff_Op_Amp_Layout_0.VB1.t33 0.4555
R20208 Folded_Diff_Op_Amp_Layout_0.VB1.n54 Folded_Diff_Op_Amp_Layout_0.VB1.n53 0.4555
R20209 Folded_Diff_Op_Amp_Layout_0.VB1.n44 Folded_Diff_Op_Amp_Layout_0.VB1.n43 0.337022
R20210 Folded_Diff_Op_Amp_Layout_0.VB1.n64 Folded_Diff_Op_Amp_Layout_0.VB1.n60 0.323326
R20211 Folded_Diff_Op_Amp_Layout_0.VB1.n81 Folded_Diff_Op_Amp_Layout_0.VB1.n77 0.323326
R20212 Folded_Diff_Op_Amp_Layout_0.VB1.n47 Folded_Diff_Op_Amp_Layout_0.VB1.n44 0.305717
R20213 Folded_Diff_Op_Amp_Layout_0.VB1.n67 Folded_Diff_Op_Amp_Layout_0.VB1.n64 0.305717
R20214 Folded_Diff_Op_Amp_Layout_0.VB1.n84 Folded_Diff_Op_Amp_Layout_0.VB1.n81 0.305717
R20215 Folded_Diff_Op_Amp_Layout_0.VB1.n64 Folded_Diff_Op_Amp_Layout_0.VB1.n63 0.303761
R20216 Folded_Diff_Op_Amp_Layout_0.VB1.n81 Folded_Diff_Op_Amp_Layout_0.VB1.n80 0.303761
R20217 Folded_Diff_Op_Amp_Layout_0.VB1.n44 Folded_Diff_Op_Amp_Layout_0.VB1.n40 0.290065
R20218 Folded_Diff_Op_Amp_Layout_0.VB1.n91 Folded_Diff_Op_Amp_Layout_0.VB1.n87 0.123658
R20219 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VB1.n100 0.110882
R20220 Folded_Diff_Op_Amp_Layout_0.VB1.n71 Folded_Diff_Op_Amp_Layout_0.VB1.n70 0.0929251
R20221 Folded_Diff_Op_Amp_Layout_0.VB1.n33 Folded_Diff_Op_Amp_Layout_0.VB1.n32 0.0656316
R20222 Folded_Diff_Op_Amp_Layout_0.VB1.n98 Folded_Diff_Op_Amp_Layout_0.VB1.n97 0.0423089
R20223 Folded_Diff_Op_Amp_Layout_0.VB1.n93 Folded_Diff_Op_Amp_Layout_0.VB1.n92 0.0324737
R20224 Folded_Diff_Op_Amp_Layout_0.VB1.n73 Folded_Diff_Op_Amp_Layout_0.VB1.n72 0.0324737
R20225 Folded_Diff_Op_Amp_Layout_0.VB1.n86 Folded_Diff_Op_Amp_Layout_0.VB1.n85 0.0324737
R20226 Folded_Diff_Op_Amp_Layout_0.VB1.n72 Folded_Diff_Op_Amp_Layout_0.VB1.n71 0.0320039
R20227 Folded_Diff_Op_Amp_Layout_0.VB1.n34 Folded_Diff_Op_Amp_Layout_0.VB1.n33 0.0301053
R20228 Folded_Diff_Op_Amp_Layout_0.VB1.n32 Folded_Diff_Op_Amp_Layout_0.VB1.n31 0.0289211
R20229 Folded_Diff_Op_Amp_Layout_0.VB1.n0 Folded_Diff_Op_Amp_Layout_0.VB1.n4 0.0222197
R20230 Folded_Diff_Op_Amp_Layout_0.VB1.n0 Folded_Diff_Op_Amp_Layout_0.VB1.n35 0.0207053
R20231 Folded_Diff_Op_Amp_Layout_0.VB1.n99 Folded_Diff_Op_Amp_Layout_0.VB1.n3 0.0201085
R20232 Folded_Diff_Op_Amp_Layout_0.VB1.n49 Folded_Diff_Op_Amp_Layout_0.VB1.n48 0.014283
R20233 Folded_Diff_Op_Amp_Layout_0.VB1.n69 Folded_Diff_Op_Amp_Layout_0.VB1.n68 0.014283
R20234 Folded_Diff_Op_Amp_Layout_0.VB1.n2 Folded_Diff_Op_Amp_Layout_0.VB1.n1 0.0127309
R20235 Folded_Diff_Op_Amp_Layout_0.VB2.n20 Folded_Diff_Op_Amp_Layout_0.VB2.t62 62.1809
R20236 Folded_Diff_Op_Amp_Layout_0.VB2.n21 Folded_Diff_Op_Amp_Layout_0.VB2.t38 62.1809
R20237 Folded_Diff_Op_Amp_Layout_0.VB2.n22 Folded_Diff_Op_Amp_Layout_0.VB2.t40 62.1809
R20238 Folded_Diff_Op_Amp_Layout_0.VB2.n23 Folded_Diff_Op_Amp_Layout_0.VB2.t34 62.1809
R20239 Folded_Diff_Op_Amp_Layout_0.VB2.n24 Folded_Diff_Op_Amp_Layout_0.VB2.t56 62.1809
R20240 Folded_Diff_Op_Amp_Layout_0.VB2.n25 Folded_Diff_Op_Amp_Layout_0.VB2.t45 62.1809
R20241 Folded_Diff_Op_Amp_Layout_0.VB2.n26 Folded_Diff_Op_Amp_Layout_0.VB2.t47 62.1809
R20242 Folded_Diff_Op_Amp_Layout_0.VB2.n11 Folded_Diff_Op_Amp_Layout_0.VB2.t64 61.6594
R20243 Folded_Diff_Op_Amp_Layout_0.VB2.n12 Folded_Diff_Op_Amp_Layout_0.VB2.t48 61.6594
R20244 Folded_Diff_Op_Amp_Layout_0.VB2.n13 Folded_Diff_Op_Amp_Layout_0.VB2.t50 61.6594
R20245 Folded_Diff_Op_Amp_Layout_0.VB2.n14 Folded_Diff_Op_Amp_Layout_0.VB2.t46 61.6594
R20246 Folded_Diff_Op_Amp_Layout_0.VB2.n15 Folded_Diff_Op_Amp_Layout_0.VB2.t61 61.6594
R20247 Folded_Diff_Op_Amp_Layout_0.VB2.n16 Folded_Diff_Op_Amp_Layout_0.VB2.t54 61.6594
R20248 Folded_Diff_Op_Amp_Layout_0.VB2.n18 Folded_Diff_Op_Amp_Layout_0.VB2.t52 61.6594
R20249 Folded_Diff_Op_Amp_Layout_0.VB2.n17 Folded_Diff_Op_Amp_Layout_0.VB2.t57 61.6594
R20250 Folded_Diff_Op_Amp_Layout_0.VB2.n4 Folded_Diff_Op_Amp_Layout_0.VB2.t58 59.8344
R20251 Folded_Diff_Op_Amp_Layout_0.VB2.n9 Folded_Diff_Op_Amp_Layout_0.VB2.t67 59.8344
R20252 Folded_Diff_Op_Amp_Layout_0.VB2.n10 Folded_Diff_Op_Amp_Layout_0.VB2.t55 59.8344
R20253 Folded_Diff_Op_Amp_Layout_0.VB2.n8 Folded_Diff_Op_Amp_Layout_0.VB2.t70 59.8344
R20254 Folded_Diff_Op_Amp_Layout_0.VB2.n5 Folded_Diff_Op_Amp_Layout_0.VB2.t53 59.8344
R20255 Folded_Diff_Op_Amp_Layout_0.VB2.n6 Folded_Diff_Op_Amp_Layout_0.VB2.t63 59.8344
R20256 Folded_Diff_Op_Amp_Layout_0.VB2.n7 Folded_Diff_Op_Amp_Layout_0.VB2.t69 59.8344
R20257 Folded_Diff_Op_Amp_Layout_0.VB2.n3 Folded_Diff_Op_Amp_Layout_0.VB2.t68 59.8344
R20258 Folded_Diff_Op_Amp_Layout_0.VB2.t48 Folded_Diff_Op_Amp_Layout_0.VB2.n10 59.5737
R20259 Folded_Diff_Op_Amp_Layout_0.VB2.t50 Folded_Diff_Op_Amp_Layout_0.VB2.n8 59.5737
R20260 Folded_Diff_Op_Amp_Layout_0.VB2.t54 Folded_Diff_Op_Amp_Layout_0.VB2.n7 59.5737
R20261 Folded_Diff_Op_Amp_Layout_0.VB2.t52 Folded_Diff_Op_Amp_Layout_0.VB2.n3 59.5737
R20262 Folded_Diff_Op_Amp_Layout_0.VB2.t57 Folded_Diff_Op_Amp_Layout_0.VB2.n4 59.5737
R20263 Folded_Diff_Op_Amp_Layout_0.VB2.t41 Folded_Diff_Op_Amp_Layout_0.VB2.n18 57.7487
R20264 Folded_Diff_Op_Amp_Layout_0.VB2.n20 Folded_Diff_Op_Amp_Layout_0.VB2.t60 57.2273
R20265 Folded_Diff_Op_Amp_Layout_0.VB2.n21 Folded_Diff_Op_Amp_Layout_0.VB2.t73 57.2273
R20266 Folded_Diff_Op_Amp_Layout_0.VB2.n22 Folded_Diff_Op_Amp_Layout_0.VB2.t35 57.2273
R20267 Folded_Diff_Op_Amp_Layout_0.VB2.n23 Folded_Diff_Op_Amp_Layout_0.VB2.t72 57.2273
R20268 Folded_Diff_Op_Amp_Layout_0.VB2.n24 Folded_Diff_Op_Amp_Layout_0.VB2.t49 57.2273
R20269 Folded_Diff_Op_Amp_Layout_0.VB2.n25 Folded_Diff_Op_Amp_Layout_0.VB2.t39 57.2273
R20270 Folded_Diff_Op_Amp_Layout_0.VB2.n26 Folded_Diff_Op_Amp_Layout_0.VB2.t42 57.2273
R20271 Folded_Diff_Op_Amp_Layout_0.VB2.n27 Folded_Diff_Op_Amp_Layout_0.VB2.t36 57.2273
R20272 Folded_Diff_Op_Amp_Layout_0.VB2.n19 Folded_Diff_Op_Amp_Layout_0.VB2.t41 56.8812
R20273 Folded_Diff_Op_Amp_Layout_0.VB2.n51 Folded_Diff_Op_Amp_Layout_0.VB2.t26 31.4166
R20274 Folded_Diff_Op_Amp_Layout_0.VB2.n63 Folded_Diff_Op_Amp_Layout_0.VB2.t44 26.7169
R20275 Folded_Diff_Op_Amp_Layout_0.VB2.n64 Folded_Diff_Op_Amp_Layout_0.VB2.n63 20.8576
R20276 Folded_Diff_Op_Amp_Layout_0.VB2.n65 Folded_Diff_Op_Amp_Layout_0.VB2.n64 20.8576
R20277 Folded_Diff_Op_Amp_Layout_0.VB2.n66 Folded_Diff_Op_Amp_Layout_0.VB2.n65 20.8576
R20278 Folded_Diff_Op_Amp_Layout_0.VB2.n67 Folded_Diff_Op_Amp_Layout_0.VB2.n66 20.8576
R20279 Folded_Diff_Op_Amp_Layout_0.VB2.n68 Folded_Diff_Op_Amp_Layout_0.VB2.n67 20.8576
R20280 Folded_Diff_Op_Amp_Layout_0.VB2.n70 Folded_Diff_Op_Amp_Layout_0.VB2.n69 20.8576
R20281 Folded_Diff_Op_Amp_Layout_0.VB2.n54 Folded_Diff_Op_Amp_Layout_0.VB2.n53 19.8148
R20282 Folded_Diff_Op_Amp_Layout_0.VB2.n44 Folded_Diff_Op_Amp_Layout_0.VB2.n43 19.8148
R20283 Folded_Diff_Op_Amp_Layout_0.VB2.n71 Folded_Diff_Op_Amp_Layout_0.VB2.n68 19.8148
R20284 Folded_Diff_Op_Amp_Layout_0.VB2.n71 Folded_Diff_Op_Amp_Layout_0.VB2.n70 19.8148
R20285 Folded_Diff_Op_Amp_Layout_0.VB2.n44 Folded_Diff_Op_Amp_Layout_0.VB2.n42 19.8148
R20286 Folded_Diff_Op_Amp_Layout_0.VB2.n10 Folded_Diff_Op_Amp_Layout_0.VB2.n9 17.5205
R20287 Folded_Diff_Op_Amp_Layout_0.VB2.n7 Folded_Diff_Op_Amp_Layout_0.VB2.n6 17.5205
R20288 Folded_Diff_Op_Amp_Layout_0.VB2.n12 Folded_Diff_Op_Amp_Layout_0.VB2.n11 17.5205
R20289 Folded_Diff_Op_Amp_Layout_0.VB2.n14 Folded_Diff_Op_Amp_Layout_0.VB2.n13 17.5205
R20290 Folded_Diff_Op_Amp_Layout_0.VB2.n16 Folded_Diff_Op_Amp_Layout_0.VB2.n15 17.5205
R20291 Folded_Diff_Op_Amp_Layout_0.VB2.n18 Folded_Diff_Op_Amp_Layout_0.VB2.n17 17.5205
R20292 Folded_Diff_Op_Amp_Layout_0.VB2.n21 Folded_Diff_Op_Amp_Layout_0.VB2.n20 17.5205
R20293 Folded_Diff_Op_Amp_Layout_0.VB2.n23 Folded_Diff_Op_Amp_Layout_0.VB2.n22 17.5205
R20294 Folded_Diff_Op_Amp_Layout_0.VB2.n25 Folded_Diff_Op_Amp_Layout_0.VB2.n24 17.5205
R20295 Folded_Diff_Op_Amp_Layout_0.VB2.n27 Folded_Diff_Op_Amp_Layout_0.VB2.n26 17.5205
R20296 Folded_Diff_Op_Amp_Layout_0.VB2.n43 Folded_Diff_Op_Amp_Layout_0.VB2.t24 11.6023
R20297 Folded_Diff_Op_Amp_Layout_0.VB2.n53 Folded_Diff_Op_Amp_Layout_0.VB2.t8 11.6023
R20298 Folded_Diff_Op_Amp_Layout_0.VB2.n63 Folded_Diff_Op_Amp_Layout_0.VB2.t16 11.6023
R20299 Folded_Diff_Op_Amp_Layout_0.VB2.n64 Folded_Diff_Op_Amp_Layout_0.VB2.t2 11.6023
R20300 Folded_Diff_Op_Amp_Layout_0.VB2.n65 Folded_Diff_Op_Amp_Layout_0.VB2.t18 11.6023
R20301 Folded_Diff_Op_Amp_Layout_0.VB2.n66 Folded_Diff_Op_Amp_Layout_0.VB2.t6 11.6023
R20302 Folded_Diff_Op_Amp_Layout_0.VB2.n67 Folded_Diff_Op_Amp_Layout_0.VB2.t12 11.6023
R20303 Folded_Diff_Op_Amp_Layout_0.VB2.n68 Folded_Diff_Op_Amp_Layout_0.VB2.t4 11.6023
R20304 Folded_Diff_Op_Amp_Layout_0.VB2.n70 Folded_Diff_Op_Amp_Layout_0.VB2.t28 11.6023
R20305 Folded_Diff_Op_Amp_Layout_0.VB2.n69 Folded_Diff_Op_Amp_Layout_0.VB2.t20 11.6023
R20306 Folded_Diff_Op_Amp_Layout_0.VB2.n42 Folded_Diff_Op_Amp_Layout_0.VB2.t30 11.6023
R20307 Folded_Diff_Op_Amp_Layout_0.VB2.n71 Folded_Diff_Op_Amp_Layout_0.VB2.t22 10.5594
R20308 Folded_Diff_Op_Amp_Layout_0.VB2.n51 Folded_Diff_Op_Amp_Layout_0.VB2.t10 10.5594
R20309 Folded_Diff_Op_Amp_Layout_0.VB2.n54 Folded_Diff_Op_Amp_Layout_0.VB2.t0 10.5594
R20310 Folded_Diff_Op_Amp_Layout_0.VB2.n44 Folded_Diff_Op_Amp_Layout_0.VB2.t14 10.5594
R20311 Folded_Diff_Op_Amp_Layout_0.VB2.n6 Folded_Diff_Op_Amp_Layout_0.VB2.n5 9.73383
R20312 Folded_Diff_Op_Amp_Layout_0.VB2.n13 Folded_Diff_Op_Amp_Layout_0.VB2.n12 9.73383
R20313 Folded_Diff_Op_Amp_Layout_0.VB2.n15 Folded_Diff_Op_Amp_Layout_0.VB2.n14 9.73383
R20314 Folded_Diff_Op_Amp_Layout_0.VB2.n17 Folded_Diff_Op_Amp_Layout_0.VB2.n16 9.73383
R20315 Folded_Diff_Op_Amp_Layout_0.VB2.n22 Folded_Diff_Op_Amp_Layout_0.VB2.n21 9.73383
R20316 Folded_Diff_Op_Amp_Layout_0.VB2.n24 Folded_Diff_Op_Amp_Layout_0.VB2.n23 9.73383
R20317 Folded_Diff_Op_Amp_Layout_0.VB2.n26 Folded_Diff_Op_Amp_Layout_0.VB2.n25 9.73383
R20318 Folded_Diff_Op_Amp_Layout_0.VB2.n77 Folded_Diff_Op_Amp_Layout_0.VB2.n75 5.92029
R20319 Folded_Diff_Op_Amp_Layout_0.VB2.n0 Folded_Diff_Op_Amp_Layout_0.VB2.n80 4.48545
R20320 Folded_Diff_Op_Amp_Layout_0.VB2.n58 Folded_Diff_Op_Amp_Layout_0.VB2.n44 4.0005
R20321 Folded_Diff_Op_Amp_Layout_0.VB2.n55 Folded_Diff_Op_Amp_Layout_0.VB2.n54 4.0005
R20322 Folded_Diff_Op_Amp_Layout_0.VB2.n52 Folded_Diff_Op_Amp_Layout_0.VB2.n51 4.0005
R20323 Folded_Diff_Op_Amp_Layout_0.VB2.n72 Folded_Diff_Op_Amp_Layout_0.VB2.n71 4.0005
R20324 Folded_Diff_Op_Amp_Layout_0.VB2.n29 Folded_Diff_Op_Amp_Layout_0.VB2.n28 3.91467
R20325 Folded_Diff_Op_Amp_Layout_0.VB2.n35 Folded_Diff_Op_Amp_Layout_0.VB2.t17 3.6405
R20326 Folded_Diff_Op_Amp_Layout_0.VB2.n35 Folded_Diff_Op_Amp_Layout_0.VB2.n34 3.6405
R20327 Folded_Diff_Op_Amp_Layout_0.VB2.n37 Folded_Diff_Op_Amp_Layout_0.VB2.t19 3.6405
R20328 Folded_Diff_Op_Amp_Layout_0.VB2.n37 Folded_Diff_Op_Amp_Layout_0.VB2.n36 3.6405
R20329 Folded_Diff_Op_Amp_Layout_0.VB2.n39 Folded_Diff_Op_Amp_Layout_0.VB2.t13 3.6405
R20330 Folded_Diff_Op_Amp_Layout_0.VB2.n39 Folded_Diff_Op_Amp_Layout_0.VB2.n38 3.6405
R20331 Folded_Diff_Op_Amp_Layout_0.VB2.n41 Folded_Diff_Op_Amp_Layout_0.VB2.t21 3.6405
R20332 Folded_Diff_Op_Amp_Layout_0.VB2.n41 Folded_Diff_Op_Amp_Layout_0.VB2.n40 3.6405
R20333 Folded_Diff_Op_Amp_Layout_0.VB2.n46 Folded_Diff_Op_Amp_Layout_0.VB2.t15 3.6405
R20334 Folded_Diff_Op_Amp_Layout_0.VB2.n46 Folded_Diff_Op_Amp_Layout_0.VB2.n45 3.6405
R20335 Folded_Diff_Op_Amp_Layout_0.VB2.n48 Folded_Diff_Op_Amp_Layout_0.VB2.t9 3.6405
R20336 Folded_Diff_Op_Amp_Layout_0.VB2.n48 Folded_Diff_Op_Amp_Layout_0.VB2.n47 3.6405
R20337 Folded_Diff_Op_Amp_Layout_0.VB2.n50 Folded_Diff_Op_Amp_Layout_0.VB2.t11 3.6405
R20338 Folded_Diff_Op_Amp_Layout_0.VB2.n50 Folded_Diff_Op_Amp_Layout_0.VB2.n49 3.6405
R20339 Folded_Diff_Op_Amp_Layout_0.VB2.n61 Folded_Diff_Op_Amp_Layout_0.VB2.t23 3.6405
R20340 Folded_Diff_Op_Amp_Layout_0.VB2.n61 Folded_Diff_Op_Amp_Layout_0.VB2.n60 3.6405
R20341 Folded_Diff_Op_Amp_Layout_0.VB2.n52 Folded_Diff_Op_Amp_Layout_0.VB2.n50 2.94093
R20342 Folded_Diff_Op_Amp_Layout_0.VB2.n32 Folded_Diff_Op_Amp_Layout_0.VB2.n19 2.8805
R20343 Folded_Diff_Op_Amp_Layout_0.VB2.n75 Folded_Diff_Op_Amp_Layout_0.VB2.n35 2.80007
R20344 Folded_Diff_Op_Amp_Layout_0.VB2.n74 Folded_Diff_Op_Amp_Layout_0.VB2.n37 2.78441
R20345 Folded_Diff_Op_Amp_Layout_0.VB2.n73 Folded_Diff_Op_Amp_Layout_0.VB2.n39 2.78441
R20346 Folded_Diff_Op_Amp_Layout_0.VB2.n59 Folded_Diff_Op_Amp_Layout_0.VB2.n41 2.78441
R20347 Folded_Diff_Op_Amp_Layout_0.VB2.n57 Folded_Diff_Op_Amp_Layout_0.VB2.n46 2.78441
R20348 Folded_Diff_Op_Amp_Layout_0.VB2.n56 Folded_Diff_Op_Amp_Layout_0.VB2.n48 2.78441
R20349 Folded_Diff_Op_Amp_Layout_0.VB2.n62 Folded_Diff_Op_Amp_Layout_0.VB2.n61 2.78441
R20350 Folded_Diff_Op_Amp_Layout_0.VB2.n78 Folded_Diff_Op_Amp_Layout_0.VB2.t32 2.53976
R20351 Folded_Diff_Op_Amp_Layout_0.VB2.n28 Folded_Diff_Op_Amp_Layout_0.VB2.n27 1.643
R20352 Folded_Diff_Op_Amp_Layout_0.VB2.n81 Folded_Diff_Op_Amp_Layout_0.VB2.n0 2.62476
R20353 Folded_Diff_Op_Amp_Layout_0.VB2.n79 Folded_Diff_Op_Amp_Layout_0.VB2.n78 1.18731
R20354 Folded_Diff_Op_Amp_Layout_0.VB2.n81 Folded_Diff_Op_Amp_Layout_0.VB2.n2 1.12594
R20355 Folded_Diff_Op_Amp_Layout_0.VB2.n74 Folded_Diff_Op_Amp_Layout_0.VB2.n73 0.626587
R20356 Folded_Diff_Op_Amp_Layout_0.VB2.n62 Folded_Diff_Op_Amp_Layout_0.VB2.n59 0.626587
R20357 Folded_Diff_Op_Amp_Layout_0.VB2.n57 Folded_Diff_Op_Amp_Layout_0.VB2.n56 0.626587
R20358 Folded_Diff_Op_Amp_Layout_0.VB2.n75 Folded_Diff_Op_Amp_Layout_0.VB2.n74 0.552239
R20359 Folded_Diff_Op_Amp_Layout_0.VB2.n73 Folded_Diff_Op_Amp_Layout_0.VB2.n72 0.470065
R20360 Folded_Diff_Op_Amp_Layout_0.VB2.n59 Folded_Diff_Op_Amp_Layout_0.VB2.n58 0.470065
R20361 Folded_Diff_Op_Amp_Layout_0.VB2.n55 Folded_Diff_Op_Amp_Layout_0.VB2.n52 0.313543
R20362 Folded_Diff_Op_Amp_Layout_0.VB2.n72 Folded_Diff_Op_Amp_Layout_0.VB2.n62 0.157022
R20363 Folded_Diff_Op_Amp_Layout_0.VB2.n58 Folded_Diff_Op_Amp_Layout_0.VB2.n57 0.157022
R20364 Folded_Diff_Op_Amp_Layout_0.VB2.n56 Folded_Diff_Op_Amp_Layout_0.VB2.n55 0.157022
R20365 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB2.n81 0.110882
R20366 Folded_Diff_Op_Amp_Layout_0.VB2.n77 Folded_Diff_Op_Amp_Layout_0.VB2.n76 0.0832399
R20367 Folded_Diff_Op_Amp_Layout_0.VB2.n31 Folded_Diff_Op_Amp_Layout_0.VB2.n30 0.0656316
R20368 Folded_Diff_Op_Amp_Layout_0.VB2.n79 Folded_Diff_Op_Amp_Layout_0.VB2.n77 0.0419676
R20369 Folded_Diff_Op_Amp_Layout_0.VB2.n32 Folded_Diff_Op_Amp_Layout_0.VB2.n31 0.0301053
R20370 Folded_Diff_Op_Amp_Layout_0.VB2.n30 Folded_Diff_Op_Amp_Layout_0.VB2.n29 0.0289211
R20371 Folded_Diff_Op_Amp_Layout_0.VB2.n2 Folded_Diff_Op_Amp_Layout_0.VB2.n1 0.0279452
R20372 Folded_Diff_Op_Amp_Layout_0.VB2.n80 Folded_Diff_Op_Amp_Layout_0.VB2.n79 0.0169282
R20373 Folded_Diff_Op_Amp_Layout_0.VB2.n2 Folded_Diff_Op_Amp_Layout_0.VB2.n32 7.26386
R20374 Folded_Diff_Op_Amp_Layout_0.VB2.n0 Folded_Diff_Op_Amp_Layout_0.VB2.n33 0.0761302
R20375 Folded_Diff_Op_Amp_Layout_0.IB2.n16 Folded_Diff_Op_Amp_Layout_0.IB2.t12 7.0505
R20376 Folded_Diff_Op_Amp_Layout_0.IB2.n15 Folded_Diff_Op_Amp_Layout_0.IB2.t3 3.6405
R20377 Folded_Diff_Op_Amp_Layout_0.IB2.n15 Folded_Diff_Op_Amp_Layout_0.IB2.n14 3.6405
R20378 Folded_Diff_Op_Amp_Layout_0.IB2.n13 Folded_Diff_Op_Amp_Layout_0.IB2.t6 3.6405
R20379 Folded_Diff_Op_Amp_Layout_0.IB2.n13 Folded_Diff_Op_Amp_Layout_0.IB2.n12 3.6405
R20380 Folded_Diff_Op_Amp_Layout_0.IB2.n11 Folded_Diff_Op_Amp_Layout_0.IB2.t10 3.6405
R20381 Folded_Diff_Op_Amp_Layout_0.IB2.n11 Folded_Diff_Op_Amp_Layout_0.IB2.n10 3.6405
R20382 Folded_Diff_Op_Amp_Layout_0.IB2.n9 Folded_Diff_Op_Amp_Layout_0.IB2.t16 3.6405
R20383 Folded_Diff_Op_Amp_Layout_0.IB2.n9 Folded_Diff_Op_Amp_Layout_0.IB2.n8 3.6405
R20384 Folded_Diff_Op_Amp_Layout_0.IB2.n1 Folded_Diff_Op_Amp_Layout_0.IB2.t5 3.6405
R20385 Folded_Diff_Op_Amp_Layout_0.IB2.n1 Folded_Diff_Op_Amp_Layout_0.IB2.n0 3.6405
R20386 Folded_Diff_Op_Amp_Layout_0.IB2.n3 Folded_Diff_Op_Amp_Layout_0.IB2.t13 3.6405
R20387 Folded_Diff_Op_Amp_Layout_0.IB2.n3 Folded_Diff_Op_Amp_Layout_0.IB2.n2 3.6405
R20388 Folded_Diff_Op_Amp_Layout_0.IB2.n5 Folded_Diff_Op_Amp_Layout_0.IB2.t0 3.6405
R20389 Folded_Diff_Op_Amp_Layout_0.IB2.n5 Folded_Diff_Op_Amp_Layout_0.IB2.n4 3.6405
R20390 Folded_Diff_Op_Amp_Layout_0.IB2.n21 Folded_Diff_Op_Amp_Layout_0.IB2.t15 3.6405
R20391 Folded_Diff_Op_Amp_Layout_0.IB2.n21 Folded_Diff_Op_Amp_Layout_0.IB2.n20 3.6405
R20392 Folded_Diff_Op_Amp_Layout_0.IB2.n6 Folded_Diff_Op_Amp_Layout_0.IB2.n5 3.4105
R20393 Folded_Diff_Op_Amp_Layout_0.IB2.n16 Folded_Diff_Op_Amp_Layout_0.IB2.n15 2.78441
R20394 Folded_Diff_Op_Amp_Layout_0.IB2.n17 Folded_Diff_Op_Amp_Layout_0.IB2.n13 2.78441
R20395 Folded_Diff_Op_Amp_Layout_0.IB2.n18 Folded_Diff_Op_Amp_Layout_0.IB2.n11 2.78441
R20396 Folded_Diff_Op_Amp_Layout_0.IB2.n19 Folded_Diff_Op_Amp_Layout_0.IB2.n9 2.78441
R20397 Folded_Diff_Op_Amp_Layout_0.IB2.n7 Folded_Diff_Op_Amp_Layout_0.IB2.n1 2.78441
R20398 Folded_Diff_Op_Amp_Layout_0.IB2.n6 Folded_Diff_Op_Amp_Layout_0.IB2.n3 2.78441
R20399 Folded_Diff_Op_Amp_Layout_0.IB2.n22 Folded_Diff_Op_Amp_Layout_0.IB2.n21 2.78441
R20400 Folded_Diff_Op_Amp_Layout_0.IB2.n7 Folded_Diff_Op_Amp_Layout_0.IB2.n6 0.626587
R20401 Folded_Diff_Op_Amp_Layout_0.IB2.n22 Folded_Diff_Op_Amp_Layout_0.IB2.n19 0.626587
R20402 Folded_Diff_Op_Amp_Layout_0.IB2.n19 Folded_Diff_Op_Amp_Layout_0.IB2.n18 0.626587
R20403 Folded_Diff_Op_Amp_Layout_0.IB2.n18 Folded_Diff_Op_Amp_Layout_0.IB2.n17 0.626587
R20404 Folded_Diff_Op_Amp_Layout_0.IB2.n17 Folded_Diff_Op_Amp_Layout_0.IB2.n16 0.626587
R20405 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.IB2.n7 0.503326
R20406 Folded_Diff_Op_Amp_Layout_0.IB2 Folded_Diff_Op_Amp_Layout_0.IB2.n22 0.123761
R20407 Folded_Diff_Op_Amp_Layout_0.IBIAS.t19 Folded_Diff_Op_Amp_Layout_0.IBIAS.t35 49.6666
R20408 Folded_Diff_Op_Amp_Layout_0.IBIAS.t18 Folded_Diff_Op_Amp_Layout_0.IBIAS.t19 49.6666
R20409 Folded_Diff_Op_Amp_Layout_0.IBIAS.t36 Folded_Diff_Op_Amp_Layout_0.IBIAS.t18 49.6666
R20410 Folded_Diff_Op_Amp_Layout_0.IBIAS.t33 Folded_Diff_Op_Amp_Layout_0.IBIAS.t14 49.6666
R20411 Folded_Diff_Op_Amp_Layout_0.IBIAS.t32 Folded_Diff_Op_Amp_Layout_0.IBIAS.t33 49.6666
R20412 Folded_Diff_Op_Amp_Layout_0.IBIAS.t17 Folded_Diff_Op_Amp_Layout_0.IBIAS.t32 49.6666
R20413 Folded_Diff_Op_Amp_Layout_0.IBIAS.t40 Folded_Diff_Op_Amp_Layout_0.IBIAS.t20 49.6666
R20414 Folded_Diff_Op_Amp_Layout_0.IBIAS.t39 Folded_Diff_Op_Amp_Layout_0.IBIAS.t40 49.6666
R20415 Folded_Diff_Op_Amp_Layout_0.IBIAS.t24 Folded_Diff_Op_Amp_Layout_0.IBIAS.t39 49.6666
R20416 Folded_Diff_Op_Amp_Layout_0.IBIAS.t44 Folded_Diff_Op_Amp_Layout_0.IBIAS.t25 49.6666
R20417 Folded_Diff_Op_Amp_Layout_0.IBIAS.t42 Folded_Diff_Op_Amp_Layout_0.IBIAS.t44 49.6666
R20418 Folded_Diff_Op_Amp_Layout_0.IBIAS.t28 Folded_Diff_Op_Amp_Layout_0.IBIAS.t42 49.6666
R20419 Folded_Diff_Op_Amp_Layout_0.IBIAS.t43 Folded_Diff_Op_Amp_Layout_0.IBIAS.t22 49.6666
R20420 Folded_Diff_Op_Amp_Layout_0.IBIAS.t41 Folded_Diff_Op_Amp_Layout_0.IBIAS.t43 49.6666
R20421 Folded_Diff_Op_Amp_Layout_0.IBIAS.t26 Folded_Diff_Op_Amp_Layout_0.IBIAS.t41 49.6666
R20422 Folded_Diff_Op_Amp_Layout_0.IBIAS.t13 Folded_Diff_Op_Amp_Layout_0.IBIAS.t27 49.6666
R20423 Folded_Diff_Op_Amp_Layout_0.IBIAS.t12 Folded_Diff_Op_Amp_Layout_0.IBIAS.t13 49.6666
R20424 Folded_Diff_Op_Amp_Layout_0.IBIAS.t29 Folded_Diff_Op_Amp_Layout_0.IBIAS.t12 49.6666
R20425 Folded_Diff_Op_Amp_Layout_0.IBIAS.t16 Folded_Diff_Op_Amp_Layout_0.IBIAS.t30 49.6666
R20426 Folded_Diff_Op_Amp_Layout_0.IBIAS.t15 Folded_Diff_Op_Amp_Layout_0.IBIAS.t16 49.6666
R20427 Folded_Diff_Op_Amp_Layout_0.IBIAS.t31 Folded_Diff_Op_Amp_Layout_0.IBIAS.t15 49.6666
R20428 Folded_Diff_Op_Amp_Layout_0.IBIAS.t23 Folded_Diff_Op_Amp_Layout_0.IBIAS.t37 49.6666
R20429 Folded_Diff_Op_Amp_Layout_0.IBIAS.t21 Folded_Diff_Op_Amp_Layout_0.IBIAS.t23 49.6666
R20430 Folded_Diff_Op_Amp_Layout_0.IBIAS.t38 Folded_Diff_Op_Amp_Layout_0.IBIAS.t21 49.6666
R20431 Folded_Diff_Op_Amp_Layout_0.IBIAS.n31 Folded_Diff_Op_Amp_Layout_0.IBIAS.t8 45.8862
R20432 Folded_Diff_Op_Amp_Layout_0.IBIAS.n22 Folded_Diff_Op_Amp_Layout_0.IBIAS.t4 39.6291
R20433 Folded_Diff_Op_Amp_Layout_0.IBIAS.n7 Folded_Diff_Op_Amp_Layout_0.IBIAS.t36 35.7835
R20434 Folded_Diff_Op_Amp_Layout_0.IBIAS.n28 Folded_Diff_Op_Amp_Layout_0.IBIAS.t2 31.8076
R20435 Folded_Diff_Op_Amp_Layout_0.IBIAS.n24 Folded_Diff_Op_Amp_Layout_0.IBIAS.t0 31.8076
R20436 Folded_Diff_Op_Amp_Layout_0.IBIAS.n31 Folded_Diff_Op_Amp_Layout_0.IBIAS.t6 31.8076
R20437 Folded_Diff_Op_Amp_Layout_0.IBIAS.n5 Folded_Diff_Op_Amp_Layout_0.IBIAS.t38 22.1612
R20438 Folded_Diff_Op_Amp_Layout_0.IBIAS.n7 Folded_Diff_Op_Amp_Layout_0.IBIAS.t17 21.705
R20439 Folded_Diff_Op_Amp_Layout_0.IBIAS.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS.t24 21.705
R20440 Folded_Diff_Op_Amp_Layout_0.IBIAS.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS.t28 21.705
R20441 Folded_Diff_Op_Amp_Layout_0.IBIAS.n10 Folded_Diff_Op_Amp_Layout_0.IBIAS.t26 21.705
R20442 Folded_Diff_Op_Amp_Layout_0.IBIAS.n11 Folded_Diff_Op_Amp_Layout_0.IBIAS.t29 21.705
R20443 Folded_Diff_Op_Amp_Layout_0.IBIAS.n12 Folded_Diff_Op_Amp_Layout_0.IBIAS.t31 21.705
R20444 Folded_Diff_Op_Amp_Layout_0.IBIAS.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS.n7 14.0791
R20445 Folded_Diff_Op_Amp_Layout_0.IBIAS.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS.n8 14.0791
R20446 Folded_Diff_Op_Amp_Layout_0.IBIAS.n10 Folded_Diff_Op_Amp_Layout_0.IBIAS.n9 14.0791
R20447 Folded_Diff_Op_Amp_Layout_0.IBIAS.n11 Folded_Diff_Op_Amp_Layout_0.IBIAS.n10 14.0791
R20448 Folded_Diff_Op_Amp_Layout_0.IBIAS.n12 Folded_Diff_Op_Amp_Layout_0.IBIAS.n11 14.0791
R20449 Folded_Diff_Op_Amp_Layout_0.IBIAS.n13 Folded_Diff_Op_Amp_Layout_0.IBIAS.n12 6.84425
R20450 Folded_Diff_Op_Amp_Layout_0.IBIAS.n16 Folded_Diff_Op_Amp_Layout_0.IBIAS.n18 6.27404
R20451 Folded_Diff_Op_Amp_Layout_0.IBIAS.n23 Folded_Diff_Op_Amp_Layout_0.IBIAS.t5 4.52093
R20452 Folded_Diff_Op_Amp_Layout_0.IBIAS.n30 Folded_Diff_Op_Amp_Layout_0.IBIAS.n19 4.0005
R20453 Folded_Diff_Op_Amp_Layout_0.IBIAS.n29 Folded_Diff_Op_Amp_Layout_0.IBIAS.n28 4.0005
R20454 Folded_Diff_Op_Amp_Layout_0.IBIAS.n2 Folded_Diff_Op_Amp_Layout_0.IBIAS.n27 4.0005
R20455 Folded_Diff_Op_Amp_Layout_0.IBIAS.n26 Folded_Diff_Op_Amp_Layout_0.IBIAS.n25 4.0005
R20456 Folded_Diff_Op_Amp_Layout_0.IBIAS.n23 Folded_Diff_Op_Amp_Layout_0.IBIAS.n22 4.0005
R20457 Folded_Diff_Op_Amp_Layout_0.IBIAS.n33 Folded_Diff_Op_Amp_Layout_0.IBIAS.n32 4.0005
R20458 Folded_Diff_Op_Amp_Layout_0.IBIAS.n2 Folded_Diff_Op_Amp_Layout_0.IBIAS.n21 3.61985
R20459 Folded_Diff_Op_Amp_Layout_0.IBIAS.n14 Folded_Diff_Op_Amp_Layout_0.IBIAS.n13 2.8805
R20460 Folded_Diff_Op_Amp_Layout_0.IBIAS.n6 Folded_Diff_Op_Amp_Layout_0.IBIAS.n5 2.8805
R20461 Folded_Diff_Op_Amp_Layout_0.IBIAS.n18 Folded_Diff_Op_Amp_Layout_0.IBIAS.t10 1.6385
R20462 Folded_Diff_Op_Amp_Layout_0.IBIAS.n18 Folded_Diff_Op_Amp_Layout_0.IBIAS.n17 1.6385
R20463 Folded_Diff_Op_Amp_Layout_0.IBIAS.n39 Folded_Diff_Op_Amp_Layout_0.IBIAS.n38 1.34737
R20464 Folded_Diff_Op_Amp_Layout_0.IBIAS.n40 Folded_Diff_Op_Amp_Layout_0.IBIAS.n39 1.14222
R20465 Folded_Diff_Op_Amp_Layout_0.IBIAS.n45 Folded_Diff_Op_Amp_Layout_0.IBIAS.n44 1.1403
R20466 Folded_Diff_Op_Amp_Layout_0.IBIAS.n36 Folded_Diff_Op_Amp_Layout_0.IBIAS.n35 1.1255
R20467 Folded_Diff_Op_Amp_Layout_0.IBIAS.n44 Folded_Diff_Op_Amp_Layout_0.IBIAS.n43 0.718974
R20468 Folded_Diff_Op_Amp_Layout_0.IBIAS.n43 Folded_Diff_Op_Amp_Layout_0.IBIAS.n1 0.631893
R20469 Folded_Diff_Op_Amp_Layout_0.IBIAS.n0 Folded_Diff_Op_Amp_Layout_0.IBIAS.n41 0.616779
R20470 Folded_Diff_Op_Amp_Layout_0.IBIAS.n32 Folded_Diff_Op_Amp_Layout_0.IBIAS.n31 0.521929
R20471 Folded_Diff_Op_Amp_Layout_0.IBIAS.n25 Folded_Diff_Op_Amp_Layout_0.IBIAS.n24 0.521929
R20472 Folded_Diff_Op_Amp_Layout_0.IBIAS.n34 Folded_Diff_Op_Amp_Layout_0.IBIAS.n33 0.500676
R20473 Folded_Diff_Op_Amp_Layout_0.IBIAS.n21 Folded_Diff_Op_Amp_Layout_0.IBIAS.t3 0.4555
R20474 Folded_Diff_Op_Amp_Layout_0.IBIAS.n21 Folded_Diff_Op_Amp_Layout_0.IBIAS.n20 0.4555
R20475 Folded_Diff_Op_Amp_Layout_0.IBIAS.n38 Folded_Diff_Op_Amp_Layout_0.IBIAS.t9 0.4555
R20476 Folded_Diff_Op_Amp_Layout_0.IBIAS.n38 Folded_Diff_Op_Amp_Layout_0.IBIAS.n37 0.4555
R20477 Folded_Diff_Op_Amp_Layout_0.IBIAS.n33 Folded_Diff_Op_Amp_Layout_0.IBIAS.n30 0.203978
R20478 Folded_Diff_Op_Amp_Layout_0.IBIAS.n30 Folded_Diff_Op_Amp_Layout_0.IBIAS.n29 0.203978
R20479 Folded_Diff_Op_Amp_Layout_0.IBIAS.n29 Folded_Diff_Op_Amp_Layout_0.IBIAS.n2 0.203978
R20480 Folded_Diff_Op_Amp_Layout_0.IBIAS.n26 Folded_Diff_Op_Amp_Layout_0.IBIAS.n23 0.203978
R20481 Folded_Diff_Op_Amp_Layout_0.IBIAS.n2 Folded_Diff_Op_Amp_Layout_0.IBIAS.n26 0.203978
R20482 Folded_Diff_Op_Amp_Layout_0.IBIAS.n45 Folded_Diff_Op_Amp_Layout_0.IBIAS.n3 0.0887019
R20483 Folded_Diff_Op_Amp_Layout_0.IBIAS.n41 Folded_Diff_Op_Amp_Layout_0.IBIAS.n36 0.0712285
R20484 Folded_Diff_Op_Amp_Layout_0.IBIAS.n15 Folded_Diff_Op_Amp_Layout_0.IBIAS.n14 0.062564
R20485 Folded_Diff_Op_Amp_Layout_0.IBIAS.n15 Folded_Diff_Op_Amp_Layout_0.IBIAS.n6 0.0620381
R20486 Folded_Diff_Op_Amp_Layout_0.IBIAS.n41 Folded_Diff_Op_Amp_Layout_0.IBIAS.n40 0.0534597
R20487 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.IBIAS.n45 0.0311329
R20488 Folded_Diff_Op_Amp_Layout_0.IBIAS.n44 Folded_Diff_Op_Amp_Layout_0.IBIAS.n4 0.0286073
R20489 Folded_Diff_Op_Amp_Layout_0.IBIAS.n43 Folded_Diff_Op_Amp_Layout_0.IBIAS.n42 0.0250648
R20490 Folded_Diff_Op_Amp_Layout_0.IBIAS.n0 Folded_Diff_Op_Amp_Layout_0.IBIAS.n16 0.016662
R20491 Folded_Diff_Op_Amp_Layout_0.IBIAS.n35 Folded_Diff_Op_Amp_Layout_0.IBIAS.n34 0.0157844
R20492 Folded_Diff_Op_Amp_Layout_0.IBIAS.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS.n0 3.83721
R20493 Folded_Diff_Op_Amp_Layout_0.IBIAS.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS.n15 0.549
R20494 Folded_Diff_Op_Amp_Layout_0.BD.n8 Folded_Diff_Op_Amp_Layout_0.BD.n7 4.81137
R20495 Folded_Diff_Op_Amp_Layout_0.BD.n13 Folded_Diff_Op_Amp_Layout_0.BD.n12 4.81137
R20496 Folded_Diff_Op_Amp_Layout_0.BD.n18 Folded_Diff_Op_Amp_Layout_0.BD.n17 4.81137
R20497 Folded_Diff_Op_Amp_Layout_0.BD.n136 Folded_Diff_Op_Amp_Layout_0.BD.n135 4.09137
R20498 Folded_Diff_Op_Amp_Layout_0.BD.n125 Folded_Diff_Op_Amp_Layout_0.BD.n124 4.09137
R20499 Folded_Diff_Op_Amp_Layout_0.BD.n147 Folded_Diff_Op_Amp_Layout_0.BD.n144 4.09137
R20500 Folded_Diff_Op_Amp_Layout_0.BD.n166 Folded_Diff_Op_Amp_Layout_0.BD.n165 4.04637
R20501 Folded_Diff_Op_Amp_Layout_0.BD.n198 Folded_Diff_Op_Amp_Layout_0.BD.n197 4.04637
R20502 Folded_Diff_Op_Amp_Layout_0.BD.n86 Folded_Diff_Op_Amp_Layout_0.BD.n85 4.04637
R20503 Folded_Diff_Op_Amp_Layout_0.BD.n50 Folded_Diff_Op_Amp_Layout_0.BD.n49 4.04637
R20504 Folded_Diff_Op_Amp_Layout_0.BD.n167 Folded_Diff_Op_Amp_Layout_0.BD.n161 3.42028
R20505 Folded_Diff_Op_Amp_Layout_0.BD.n166 Folded_Diff_Op_Amp_Layout_0.BD.n163 3.42028
R20506 Folded_Diff_Op_Amp_Layout_0.BD.n199 Folded_Diff_Op_Amp_Layout_0.BD.n193 3.42028
R20507 Folded_Diff_Op_Amp_Layout_0.BD.n198 Folded_Diff_Op_Amp_Layout_0.BD.n195 3.42028
R20508 Folded_Diff_Op_Amp_Layout_0.BD.n87 Folded_Diff_Op_Amp_Layout_0.BD.n81 3.42028
R20509 Folded_Diff_Op_Amp_Layout_0.BD.n86 Folded_Diff_Op_Amp_Layout_0.BD.n83 3.42028
R20510 Folded_Diff_Op_Amp_Layout_0.BD.n51 Folded_Diff_Op_Amp_Layout_0.BD.n45 3.42028
R20511 Folded_Diff_Op_Amp_Layout_0.BD.n50 Folded_Diff_Op_Amp_Layout_0.BD.n47 3.42028
R20512 Folded_Diff_Op_Amp_Layout_0.BD.n136 Folded_Diff_Op_Amp_Layout_0.BD.n133 2.6005
R20513 Folded_Diff_Op_Amp_Layout_0.BD.n137 Folded_Diff_Op_Amp_Layout_0.BD.n131 2.6005
R20514 Folded_Diff_Op_Amp_Layout_0.BD.n138 Folded_Diff_Op_Amp_Layout_0.BD.n129 2.6005
R20515 Folded_Diff_Op_Amp_Layout_0.BD.n125 Folded_Diff_Op_Amp_Layout_0.BD.n122 2.6005
R20516 Folded_Diff_Op_Amp_Layout_0.BD.n126 Folded_Diff_Op_Amp_Layout_0.BD.n120 2.6005
R20517 Folded_Diff_Op_Amp_Layout_0.BD.n127 Folded_Diff_Op_Amp_Layout_0.BD.n118 2.6005
R20518 Folded_Diff_Op_Amp_Layout_0.BD.n8 Folded_Diff_Op_Amp_Layout_0.BD.n5 2.6005
R20519 Folded_Diff_Op_Amp_Layout_0.BD.n13 Folded_Diff_Op_Amp_Layout_0.BD.n10 2.6005
R20520 Folded_Diff_Op_Amp_Layout_0.BD.n18 Folded_Diff_Op_Amp_Layout_0.BD.n15 2.6005
R20521 Folded_Diff_Op_Amp_Layout_0.BD.n23 Folded_Diff_Op_Amp_Layout_0.BD.n22 2.6005
R20522 Folded_Diff_Op_Amp_Layout_0.BD.n75 Folded_Diff_Op_Amp_Layout_0.BD.n43 2.6005
R20523 Folded_Diff_Op_Amp_Layout_0.BD.n148 Folded_Diff_Op_Amp_Layout_0.BD.n142 2.6005
R20524 Folded_Diff_Op_Amp_Layout_0.BD.n149 Folded_Diff_Op_Amp_Layout_0.BD.n140 2.6005
R20525 Folded_Diff_Op_Amp_Layout_0.BD.n147 Folded_Diff_Op_Amp_Layout_0.BD.n146 2.6005
R20526 Folded_Diff_Op_Amp_Layout_0.BD.n24 Folded_Diff_Op_Amp_Layout_0.BD.n23 1.79659
R20527 Folded_Diff_Op_Amp_Layout_0.BD.n155 Folded_Diff_Op_Amp_Layout_0.BD.n154 1.64287
R20528 Folded_Diff_Op_Amp_Layout_0.BD.n150 Folded_Diff_Op_Amp_Layout_0.BD.n138 1.5442
R20529 Folded_Diff_Op_Amp_Layout_0.BD.n79 Folded_Diff_Op_Amp_Layout_0.BD.n41 1.54399
R20530 Folded_Diff_Op_Amp_Layout_0.BD.n0 Folded_Diff_Op_Amp_Layout_0.BD.n191 1.50472
R20531 Folded_Diff_Op_Amp_Layout_0.BD.n203 Folded_Diff_Op_Amp_Layout_0.BD.n202 1.50128
R20532 Folded_Diff_Op_Amp_Layout_0.BD.n210 Folded_Diff_Op_Amp_Layout_0.BD.n209 1.49812
R20533 Folded_Diff_Op_Amp_Layout_0.BD.n3 Folded_Diff_Op_Amp_Layout_0.BD.n2 1.49812
R20534 Folded_Diff_Op_Amp_Layout_0.BD.n109 Folded_Diff_Op_Amp_Layout_0.BD.n38 1.49812
R20535 Folded_Diff_Op_Amp_Layout_0.BD.n210 Folded_Diff_Op_Amp_Layout_0.BD.n206 1.49801
R20536 Folded_Diff_Op_Amp_Layout_0.BD.n184 Folded_Diff_Op_Amp_Layout_0.BD.n183 1.49801
R20537 Folded_Diff_Op_Amp_Layout_0.BD.n116 Folded_Diff_Op_Amp_Layout_0.BD.n115 1.49801
R20538 Folded_Diff_Op_Amp_Layout_0.BD.n138 Folded_Diff_Op_Amp_Layout_0.BD.n137 1.49137
R20539 Folded_Diff_Op_Amp_Layout_0.BD.n137 Folded_Diff_Op_Amp_Layout_0.BD.n136 1.49137
R20540 Folded_Diff_Op_Amp_Layout_0.BD.n127 Folded_Diff_Op_Amp_Layout_0.BD.n126 1.49137
R20541 Folded_Diff_Op_Amp_Layout_0.BD.n126 Folded_Diff_Op_Amp_Layout_0.BD.n125 1.49137
R20542 Folded_Diff_Op_Amp_Layout_0.BD.n149 Folded_Diff_Op_Amp_Layout_0.BD.n148 1.49137
R20543 Folded_Diff_Op_Amp_Layout_0.BD.n148 Folded_Diff_Op_Amp_Layout_0.BD.n147 1.49137
R20544 Folded_Diff_Op_Amp_Layout_0.BD.n0 Folded_Diff_Op_Amp_Layout_0.BD.n187 1.48107
R20545 Folded_Diff_Op_Amp_Layout_0.BD.n19 Folded_Diff_Op_Amp_Layout_0.BD.n18 1.44637
R20546 Folded_Diff_Op_Amp_Layout_0.BD.n23 Folded_Diff_Op_Amp_Layout_0.BD.n20 1.44637
R20547 Folded_Diff_Op_Amp_Layout_0.BD.n179 Folded_Diff_Op_Amp_Layout_0.BD.n159 1.36943
R20548 Folded_Diff_Op_Amp_Layout_0.BD.n179 Folded_Diff_Op_Amp_Layout_0.BD.n178 1.33886
R20549 Folded_Diff_Op_Amp_Layout_0.BD.n152 Folded_Diff_Op_Amp_Layout_0.BD.n151 1.28649
R20550 Folded_Diff_Op_Amp_Layout_0.BD.n72 Folded_Diff_Op_Amp_Layout_0.BD.n71 1.26677
R20551 Folded_Diff_Op_Amp_Layout_0.BD.n30 Folded_Diff_Op_Amp_Layout_0.BD.n29 1.17988
R20552 Folded_Diff_Op_Amp_Layout_0.BD.n58 Folded_Diff_Op_Amp_Layout_0.BD.n57 1.16583
R20553 Folded_Diff_Op_Amp_Layout_0.BD.n174 Folded_Diff_Op_Amp_Layout_0.BD.n173 1.1658
R20554 Folded_Diff_Op_Amp_Layout_0.BD.n191 Folded_Diff_Op_Amp_Layout_0.BD.n190 1.1658
R20555 Folded_Diff_Op_Amp_Layout_0.BD.n94 Folded_Diff_Op_Amp_Layout_0.BD.n93 1.1658
R20556 Folded_Diff_Op_Amp_Layout_0.BD.n72 Folded_Diff_Op_Amp_Layout_0.BD.n69 1.14125
R20557 Folded_Diff_Op_Amp_Layout_0.BD.n211 Folded_Diff_Op_Amp_Layout_0.BD.n210 1.12725
R20558 Folded_Diff_Op_Amp_Layout_0.BD.n211 Folded_Diff_Op_Amp_Layout_0.BD.n185 1.12594
R20559 Folded_Diff_Op_Amp_Layout_0.BD.n26 Folded_Diff_Op_Amp_Layout_0.BD.n25 1.1255
R20560 Folded_Diff_Op_Amp_Layout_0.BD.n170 Folded_Diff_Op_Amp_Layout_0.BD.n169 1.1255
R20561 Folded_Diff_Op_Amp_Layout_0.BD.n202 Folded_Diff_Op_Amp_Layout_0.BD.n201 1.1255
R20562 Folded_Diff_Op_Amp_Layout_0.BD.n90 Folded_Diff_Op_Amp_Layout_0.BD.n89 1.1255
R20563 Folded_Diff_Op_Amp_Layout_0.BD.n54 Folded_Diff_Op_Amp_Layout_0.BD.n53 1.1255
R20564 Folded_Diff_Op_Amp_Layout_0.BD.n73 Folded_Diff_Op_Amp_Layout_0.BD.n68 1.1255
R20565 Folded_Diff_Op_Amp_Layout_0.BD.n105 Folded_Diff_Op_Amp_Layout_0.BD.n104 1.1255
R20566 Folded_Diff_Op_Amp_Layout_0.BD.n78 Folded_Diff_Op_Amp_Layout_0.BD.n77 1.1255
R20567 Folded_Diff_Op_Amp_Layout_0.BD.n75 Folded_Diff_Op_Amp_Layout_0.BD.n74 1.11357
R20568 Folded_Diff_Op_Amp_Layout_0.BD.n103 Folded_Diff_Op_Amp_Layout_0.BD.n102 1.10736
R20569 Folded_Diff_Op_Amp_Layout_0.BD.n67 Folded_Diff_Op_Amp_Layout_0.BD.n66 1.10736
R20570 Folded_Diff_Op_Amp_Layout_0.BD.n76 Folded_Diff_Op_Amp_Layout_0.BD.n75 1.01985
R20571 Folded_Diff_Op_Amp_Layout_0.BD.n173 Folded_Diff_Op_Amp_Layout_0.BD.n172 1.00677
R20572 Folded_Diff_Op_Amp_Layout_0.BD.n190 Folded_Diff_Op_Amp_Layout_0.BD.n189 1.00677
R20573 Folded_Diff_Op_Amp_Layout_0.BD.n93 Folded_Diff_Op_Amp_Layout_0.BD.n92 1.00677
R20574 Folded_Diff_Op_Amp_Layout_0.BD.n107 Folded_Diff_Op_Amp_Layout_0.BD.n106 0.984698
R20575 Folded_Diff_Op_Amp_Layout_0.BD.n52 Folded_Diff_Op_Amp_Layout_0.BD.n51 0.968978
R20576 Folded_Diff_Op_Amp_Layout_0.BD.n57 Folded_Diff_Op_Amp_Layout_0.BD.n56 0.966825
R20577 Folded_Diff_Op_Amp_Layout_0.BD.n29 Folded_Diff_Op_Amp_Layout_0.BD.n28 0.963628
R20578 Folded_Diff_Op_Amp_Layout_0.BD.n151 Folded_Diff_Op_Amp_Layout_0.BD.n150 0.845717
R20579 Folded_Diff_Op_Amp_Layout_0.BD.n20 Folded_Diff_Op_Amp_Layout_0.BD.n8 0.820283
R20580 Folded_Diff_Op_Amp_Layout_0.BD.n19 Folded_Diff_Op_Amp_Layout_0.BD.n13 0.820283
R20581 Folded_Diff_Op_Amp_Layout_0.BD.n168 Folded_Diff_Op_Amp_Layout_0.BD.n167 0.773326
R20582 Folded_Diff_Op_Amp_Layout_0.BD.n200 Folded_Diff_Op_Amp_Layout_0.BD.n199 0.773326
R20583 Folded_Diff_Op_Amp_Layout_0.BD.n88 Folded_Diff_Op_Amp_Layout_0.BD.n87 0.773326
R20584 Folded_Diff_Op_Amp_Layout_0.BD.n99 Folded_Diff_Op_Amp_Layout_0.BD.n98 0.761
R20585 Folded_Diff_Op_Amp_Layout_0.BD.n63 Folded_Diff_Op_Amp_Layout_0.BD.n62 0.761
R20586 Folded_Diff_Op_Amp_Layout_0.BD.n35 Folded_Diff_Op_Amp_Layout_0.BD.n34 0.760312
R20587 Folded_Diff_Op_Amp_Layout_0.BD.n205 Folded_Diff_Op_Amp_Layout_0.BD.n204 0.760312
R20588 Folded_Diff_Op_Amp_Layout_0.BD.n157 Folded_Diff_Op_Amp_Layout_0.BD.n156 0.7505
R20589 Folded_Diff_Op_Amp_Layout_0.BD.n109 Folded_Diff_Op_Amp_Layout_0.BD.n108 0.7505
R20590 Folded_Diff_Op_Amp_Layout_0.BD.n151 Folded_Diff_Op_Amp_Layout_0.BD.n127 0.698978
R20591 Folded_Diff_Op_Amp_Layout_0.BD.n150 Folded_Diff_Op_Amp_Layout_0.BD.n149 0.698978
R20592 Folded_Diff_Op_Amp_Layout_0.BD.n20 Folded_Diff_Op_Amp_Layout_0.BD.n19 0.626587
R20593 Folded_Diff_Op_Amp_Layout_0.BD.n167 Folded_Diff_Op_Amp_Layout_0.BD.n166 0.626587
R20594 Folded_Diff_Op_Amp_Layout_0.BD.n199 Folded_Diff_Op_Amp_Layout_0.BD.n198 0.626587
R20595 Folded_Diff_Op_Amp_Layout_0.BD.n87 Folded_Diff_Op_Amp_Layout_0.BD.n86 0.626587
R20596 Folded_Diff_Op_Amp_Layout_0.BD.n51 Folded_Diff_Op_Amp_Layout_0.BD.n50 0.626587
R20597 Folded_Diff_Op_Amp_Layout_0.BD.n33 Folded_Diff_Op_Amp_Layout_0.BD.n31 0.616779
R20598 Folded_Diff_Op_Amp_Layout_0.BD.n177 Folded_Diff_Op_Amp_Layout_0.BD.n175 0.616779
R20599 Folded_Diff_Op_Amp_Layout_0.BD.n97 Folded_Diff_Op_Amp_Layout_0.BD.n95 0.616779
R20600 Folded_Diff_Op_Amp_Layout_0.BD.n61 Folded_Diff_Op_Amp_Layout_0.BD.n59 0.616779
R20601 Folded_Diff_Op_Amp_Layout_0.BD.n180 Folded_Diff_Op_Amp_Layout_0.BD.n179 0.585272
R20602 Folded_Diff_Op_Amp_Layout_0.BD.n140 Folded_Diff_Op_Amp_Layout_0.BD.t21 0.58197
R20603 Folded_Diff_Op_Amp_Layout_0.BD.n140 Folded_Diff_Op_Amp_Layout_0.BD.n139 0.58197
R20604 Folded_Diff_Op_Amp_Layout_0.BD.n142 Folded_Diff_Op_Amp_Layout_0.BD.t1 0.58197
R20605 Folded_Diff_Op_Amp_Layout_0.BD.n142 Folded_Diff_Op_Amp_Layout_0.BD.n141 0.58197
R20606 Folded_Diff_Op_Amp_Layout_0.BD.n144 Folded_Diff_Op_Amp_Layout_0.BD.t17 0.58197
R20607 Folded_Diff_Op_Amp_Layout_0.BD.n144 Folded_Diff_Op_Amp_Layout_0.BD.n143 0.58197
R20608 Folded_Diff_Op_Amp_Layout_0.BD.n129 Folded_Diff_Op_Amp_Layout_0.BD.t13 0.58197
R20609 Folded_Diff_Op_Amp_Layout_0.BD.n129 Folded_Diff_Op_Amp_Layout_0.BD.n128 0.58197
R20610 Folded_Diff_Op_Amp_Layout_0.BD.n131 Folded_Diff_Op_Amp_Layout_0.BD.t27 0.58197
R20611 Folded_Diff_Op_Amp_Layout_0.BD.n131 Folded_Diff_Op_Amp_Layout_0.BD.n130 0.58197
R20612 Folded_Diff_Op_Amp_Layout_0.BD.n133 Folded_Diff_Op_Amp_Layout_0.BD.t28 0.58197
R20613 Folded_Diff_Op_Amp_Layout_0.BD.n133 Folded_Diff_Op_Amp_Layout_0.BD.n132 0.58197
R20614 Folded_Diff_Op_Amp_Layout_0.BD.n135 Folded_Diff_Op_Amp_Layout_0.BD.t12 0.58197
R20615 Folded_Diff_Op_Amp_Layout_0.BD.n135 Folded_Diff_Op_Amp_Layout_0.BD.n134 0.58197
R20616 Folded_Diff_Op_Amp_Layout_0.BD.n118 Folded_Diff_Op_Amp_Layout_0.BD.t23 0.58197
R20617 Folded_Diff_Op_Amp_Layout_0.BD.n118 Folded_Diff_Op_Amp_Layout_0.BD.n117 0.58197
R20618 Folded_Diff_Op_Amp_Layout_0.BD.n120 Folded_Diff_Op_Amp_Layout_0.BD.t4 0.58197
R20619 Folded_Diff_Op_Amp_Layout_0.BD.n120 Folded_Diff_Op_Amp_Layout_0.BD.n119 0.58197
R20620 Folded_Diff_Op_Amp_Layout_0.BD.n122 Folded_Diff_Op_Amp_Layout_0.BD.t5 0.58197
R20621 Folded_Diff_Op_Amp_Layout_0.BD.n122 Folded_Diff_Op_Amp_Layout_0.BD.n121 0.58197
R20622 Folded_Diff_Op_Amp_Layout_0.BD.n124 Folded_Diff_Op_Amp_Layout_0.BD.t19 0.58197
R20623 Folded_Diff_Op_Amp_Layout_0.BD.n124 Folded_Diff_Op_Amp_Layout_0.BD.n123 0.58197
R20624 Folded_Diff_Op_Amp_Layout_0.BD.n154 Folded_Diff_Op_Amp_Layout_0.BD.t9 0.58197
R20625 Folded_Diff_Op_Amp_Layout_0.BD.n154 Folded_Diff_Op_Amp_Layout_0.BD.n153 0.58197
R20626 Folded_Diff_Op_Amp_Layout_0.BD.n41 Folded_Diff_Op_Amp_Layout_0.BD.t24 0.58197
R20627 Folded_Diff_Op_Amp_Layout_0.BD.n41 Folded_Diff_Op_Amp_Layout_0.BD.n40 0.58197
R20628 Folded_Diff_Op_Amp_Layout_0.BD.n43 Folded_Diff_Op_Amp_Layout_0.BD.t25 0.58197
R20629 Folded_Diff_Op_Amp_Layout_0.BD.n43 Folded_Diff_Op_Amp_Layout_0.BD.n42 0.58197
R20630 Folded_Diff_Op_Amp_Layout_0.BD.n71 Folded_Diff_Op_Amp_Layout_0.BD.t8 0.58197
R20631 Folded_Diff_Op_Amp_Layout_0.BD.n71 Folded_Diff_Op_Amp_Layout_0.BD.n70 0.58197
R20632 Folded_Diff_Op_Amp_Layout_0.BD.n146 Folded_Diff_Op_Amp_Layout_0.BD.t3 0.58197
R20633 Folded_Diff_Op_Amp_Layout_0.BD.n146 Folded_Diff_Op_Amp_Layout_0.BD.n145 0.58197
R20634 Folded_Diff_Op_Amp_Layout_0.BD.n22 Folded_Diff_Op_Amp_Layout_0.BD.t42 0.485833
R20635 Folded_Diff_Op_Amp_Layout_0.BD.n22 Folded_Diff_Op_Amp_Layout_0.BD.n21 0.485833
R20636 Folded_Diff_Op_Amp_Layout_0.BD.n5 Folded_Diff_Op_Amp_Layout_0.BD.t56 0.485833
R20637 Folded_Diff_Op_Amp_Layout_0.BD.n5 Folded_Diff_Op_Amp_Layout_0.BD.n4 0.485833
R20638 Folded_Diff_Op_Amp_Layout_0.BD.n7 Folded_Diff_Op_Amp_Layout_0.BD.t59 0.485833
R20639 Folded_Diff_Op_Amp_Layout_0.BD.n7 Folded_Diff_Op_Amp_Layout_0.BD.n6 0.485833
R20640 Folded_Diff_Op_Amp_Layout_0.BD.n10 Folded_Diff_Op_Amp_Layout_0.BD.t70 0.485833
R20641 Folded_Diff_Op_Amp_Layout_0.BD.n10 Folded_Diff_Op_Amp_Layout_0.BD.n9 0.485833
R20642 Folded_Diff_Op_Amp_Layout_0.BD.n12 Folded_Diff_Op_Amp_Layout_0.BD.t36 0.485833
R20643 Folded_Diff_Op_Amp_Layout_0.BD.n12 Folded_Diff_Op_Amp_Layout_0.BD.n11 0.485833
R20644 Folded_Diff_Op_Amp_Layout_0.BD.n15 Folded_Diff_Op_Amp_Layout_0.BD.t61 0.485833
R20645 Folded_Diff_Op_Amp_Layout_0.BD.n15 Folded_Diff_Op_Amp_Layout_0.BD.n14 0.485833
R20646 Folded_Diff_Op_Amp_Layout_0.BD.n17 Folded_Diff_Op_Amp_Layout_0.BD.t51 0.485833
R20647 Folded_Diff_Op_Amp_Layout_0.BD.n17 Folded_Diff_Op_Amp_Layout_0.BD.n16 0.485833
R20648 Folded_Diff_Op_Amp_Layout_0.BD.n28 Folded_Diff_Op_Amp_Layout_0.BD.t74 0.485833
R20649 Folded_Diff_Op_Amp_Layout_0.BD.n28 Folded_Diff_Op_Amp_Layout_0.BD.n27 0.485833
R20650 Folded_Diff_Op_Amp_Layout_0.BD.n161 Folded_Diff_Op_Amp_Layout_0.BD.t41 0.485833
R20651 Folded_Diff_Op_Amp_Layout_0.BD.n161 Folded_Diff_Op_Amp_Layout_0.BD.n160 0.485833
R20652 Folded_Diff_Op_Amp_Layout_0.BD.n163 Folded_Diff_Op_Amp_Layout_0.BD.t55 0.485833
R20653 Folded_Diff_Op_Amp_Layout_0.BD.n163 Folded_Diff_Op_Amp_Layout_0.BD.n162 0.485833
R20654 Folded_Diff_Op_Amp_Layout_0.BD.n165 Folded_Diff_Op_Amp_Layout_0.BD.t34 0.485833
R20655 Folded_Diff_Op_Amp_Layout_0.BD.n165 Folded_Diff_Op_Amp_Layout_0.BD.n164 0.485833
R20656 Folded_Diff_Op_Amp_Layout_0.BD.n172 Folded_Diff_Op_Amp_Layout_0.BD.t66 0.485833
R20657 Folded_Diff_Op_Amp_Layout_0.BD.n172 Folded_Diff_Op_Amp_Layout_0.BD.n171 0.485833
R20658 Folded_Diff_Op_Amp_Layout_0.BD.n193 Folded_Diff_Op_Amp_Layout_0.BD.t65 0.485833
R20659 Folded_Diff_Op_Amp_Layout_0.BD.n193 Folded_Diff_Op_Amp_Layout_0.BD.n192 0.485833
R20660 Folded_Diff_Op_Amp_Layout_0.BD.n195 Folded_Diff_Op_Amp_Layout_0.BD.t40 0.485833
R20661 Folded_Diff_Op_Amp_Layout_0.BD.n195 Folded_Diff_Op_Amp_Layout_0.BD.n194 0.485833
R20662 Folded_Diff_Op_Amp_Layout_0.BD.n197 Folded_Diff_Op_Amp_Layout_0.BD.t50 0.485833
R20663 Folded_Diff_Op_Amp_Layout_0.BD.n197 Folded_Diff_Op_Amp_Layout_0.BD.n196 0.485833
R20664 Folded_Diff_Op_Amp_Layout_0.BD.n189 Folded_Diff_Op_Amp_Layout_0.BD.t69 0.485833
R20665 Folded_Diff_Op_Amp_Layout_0.BD.n189 Folded_Diff_Op_Amp_Layout_0.BD.n188 0.485833
R20666 Folded_Diff_Op_Amp_Layout_0.BD.n81 Folded_Diff_Op_Amp_Layout_0.BD.t72 0.485833
R20667 Folded_Diff_Op_Amp_Layout_0.BD.n81 Folded_Diff_Op_Amp_Layout_0.BD.n80 0.485833
R20668 Folded_Diff_Op_Amp_Layout_0.BD.n83 Folded_Diff_Op_Amp_Layout_0.BD.t58 0.485833
R20669 Folded_Diff_Op_Amp_Layout_0.BD.n83 Folded_Diff_Op_Amp_Layout_0.BD.n82 0.485833
R20670 Folded_Diff_Op_Amp_Layout_0.BD.n85 Folded_Diff_Op_Amp_Layout_0.BD.t33 0.485833
R20671 Folded_Diff_Op_Amp_Layout_0.BD.n85 Folded_Diff_Op_Amp_Layout_0.BD.n84 0.485833
R20672 Folded_Diff_Op_Amp_Layout_0.BD.n92 Folded_Diff_Op_Amp_Layout_0.BD.t46 0.485833
R20673 Folded_Diff_Op_Amp_Layout_0.BD.n92 Folded_Diff_Op_Amp_Layout_0.BD.n91 0.485833
R20674 Folded_Diff_Op_Amp_Layout_0.BD.n45 Folded_Diff_Op_Amp_Layout_0.BD.t44 0.485833
R20675 Folded_Diff_Op_Amp_Layout_0.BD.n45 Folded_Diff_Op_Amp_Layout_0.BD.n44 0.485833
R20676 Folded_Diff_Op_Amp_Layout_0.BD.n47 Folded_Diff_Op_Amp_Layout_0.BD.t71 0.485833
R20677 Folded_Diff_Op_Amp_Layout_0.BD.n47 Folded_Diff_Op_Amp_Layout_0.BD.n46 0.485833
R20678 Folded_Diff_Op_Amp_Layout_0.BD.n49 Folded_Diff_Op_Amp_Layout_0.BD.t62 0.485833
R20679 Folded_Diff_Op_Amp_Layout_0.BD.n49 Folded_Diff_Op_Amp_Layout_0.BD.n48 0.485833
R20680 Folded_Diff_Op_Amp_Layout_0.BD.n56 Folded_Diff_Op_Amp_Layout_0.BD.t38 0.485833
R20681 Folded_Diff_Op_Amp_Layout_0.BD.n56 Folded_Diff_Op_Amp_Layout_0.BD.n55 0.485833
R20682 Folded_Diff_Op_Amp_Layout_0.BD.n25 Folded_Diff_Op_Amp_Layout_0.BD.n24 0.3155
R20683 Folded_Diff_Op_Amp_Layout_0.BD.n53 Folded_Diff_Op_Amp_Layout_0.BD.n52 0.252891
R20684 Folded_Diff_Op_Amp_Layout_0.BD.n108 Folded_Diff_Op_Amp_Layout_0.BD.n107 0.213196
R20685 Folded_Diff_Op_Amp_Layout_0.BD.n106 Folded_Diff_Op_Amp_Layout_0.BD.n105 0.204046
R20686 Folded_Diff_Op_Amp_Layout_0.BD.n78 Folded_Diff_Op_Amp_Layout_0.BD.n76 0.137457
R20687 Folded_Diff_Op_Amp_Layout_0.BD.n73 Folded_Diff_Op_Amp_Layout_0.BD.n72 0.109357
R20688 Folded_Diff_Op_Amp_Layout_0.BD.n156 Folded_Diff_Op_Amp_Layout_0.BD.n152 0.097556
R20689 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.BD.n211 0.0906317
R20690 Folded_Diff_Op_Amp_Layout_0.BD.n31 Folded_Diff_Op_Amp_Layout_0.BD.n26 0.0712285
R20691 Folded_Diff_Op_Amp_Layout_0.BD.n175 Folded_Diff_Op_Amp_Layout_0.BD.n170 0.0712285
R20692 Folded_Diff_Op_Amp_Layout_0.BD.n95 Folded_Diff_Op_Amp_Layout_0.BD.n90 0.0712285
R20693 Folded_Diff_Op_Amp_Layout_0.BD.n59 Folded_Diff_Op_Amp_Layout_0.BD.n54 0.0712285
R20694 Folded_Diff_Op_Amp_Layout_0.BD.n74 Folded_Diff_Op_Amp_Layout_0.BD.n73 0.0698213
R20695 Folded_Diff_Op_Amp_Layout_0.BD.n79 Folded_Diff_Op_Amp_Layout_0.BD.n78 0.0624212
R20696 Folded_Diff_Op_Amp_Layout_0.BD.n105 Folded_Diff_Op_Amp_Layout_0.BD.n79 0.0620608
R20697 Folded_Diff_Op_Amp_Layout_0.BD.n169 Folded_Diff_Op_Amp_Layout_0.BD.n168 0.0572391
R20698 Folded_Diff_Op_Amp_Layout_0.BD.n201 Folded_Diff_Op_Amp_Layout_0.BD.n200 0.0572391
R20699 Folded_Diff_Op_Amp_Layout_0.BD.n89 Folded_Diff_Op_Amp_Layout_0.BD.n88 0.0572391
R20700 Folded_Diff_Op_Amp_Layout_0.BD.n31 Folded_Diff_Op_Amp_Layout_0.BD.n30 0.0534597
R20701 Folded_Diff_Op_Amp_Layout_0.BD.n175 Folded_Diff_Op_Amp_Layout_0.BD.n174 0.0534597
R20702 Folded_Diff_Op_Amp_Layout_0.BD.n95 Folded_Diff_Op_Amp_Layout_0.BD.n94 0.0534597
R20703 Folded_Diff_Op_Amp_Layout_0.BD.n59 Folded_Diff_Op_Amp_Layout_0.BD.n58 0.0534597
R20704 Folded_Diff_Op_Amp_Layout_0.BD.n156 Folded_Diff_Op_Amp_Layout_0.BD.n155 0.0364864
R20705 Folded_Diff_Op_Amp_Layout_0.BD.n104 Folded_Diff_Op_Amp_Layout_0.BD.n103 0.0320039
R20706 Folded_Diff_Op_Amp_Layout_0.BD.n68 Folded_Diff_Op_Amp_Layout_0.BD.n67 0.0320039
R20707 Folded_Diff_Op_Amp_Layout_0.BD.n113 Folded_Diff_Op_Amp_Layout_0.BD.n112 0.0229474
R20708 Folded_Diff_Op_Amp_Layout_0.BD.n116 Folded_Diff_Op_Amp_Layout_0.BD.n111 0.0229474
R20709 Folded_Diff_Op_Amp_Layout_0.BD.n34 Folded_Diff_Op_Amp_Layout_0.BD.n33 0.0156875
R20710 Folded_Diff_Op_Amp_Layout_0.BD.n178 Folded_Diff_Op_Amp_Layout_0.BD.n177 0.0156875
R20711 Folded_Diff_Op_Amp_Layout_0.BD.n98 Folded_Diff_Op_Amp_Layout_0.BD.n97 0.0156875
R20712 Folded_Diff_Op_Amp_Layout_0.BD.n62 Folded_Diff_Op_Amp_Layout_0.BD.n61 0.0156875
R20713 Folded_Diff_Op_Amp_Layout_0.BD.n115 Folded_Diff_Op_Amp_Layout_0.BD.n114 0.014
R20714 Folded_Diff_Op_Amp_Layout_0.BD.n183 Folded_Diff_Op_Amp_Layout_0.BD.n182 0.014
R20715 Folded_Diff_Op_Amp_Layout_0.BD.n2 Folded_Diff_Op_Amp_Layout_0.BD.n1 0.014
R20716 Folded_Diff_Op_Amp_Layout_0.BD.n210 Folded_Diff_Op_Amp_Layout_0.BD.n186 0.014
R20717 Folded_Diff_Op_Amp_Layout_0.BD.n210 Folded_Diff_Op_Amp_Layout_0.BD.n208 0.014
R20718 Folded_Diff_Op_Amp_Layout_0.BD.n110 Folded_Diff_Op_Amp_Layout_0.BD.n109 0.014
R20719 Folded_Diff_Op_Amp_Layout_0.BD.n109 Folded_Diff_Op_Amp_Layout_0.BD.n39 0.014
R20720 Folded_Diff_Op_Amp_Layout_0.BD.n208 Folded_Diff_Op_Amp_Layout_0.BD.n207 0.0134654
R20721 Folded_Diff_Op_Amp_Layout_0.BD.n182 Folded_Diff_Op_Amp_Layout_0.BD.n181 0.0134654
R20722 Folded_Diff_Op_Amp_Layout_0.BD.n111 Folded_Diff_Op_Amp_Layout_0.BD.n110 0.0134654
R20723 Folded_Diff_Op_Amp_Layout_0.BD.n204 Folded_Diff_Op_Amp_Layout_0.BD.n203 0.0117561
R20724 Folded_Diff_Op_Amp_Layout_0.BD.n100 Folded_Diff_Op_Amp_Layout_0.BD.n99 0.0111023
R20725 Folded_Diff_Op_Amp_Layout_0.BD.n64 Folded_Diff_Op_Amp_Layout_0.BD.n63 0.0111023
R20726 Folded_Diff_Op_Amp_Layout_0.BD.n184 Folded_Diff_Op_Amp_Layout_0.BD.n180 0.00998204
R20727 Folded_Diff_Op_Amp_Layout_0.BD.n206 Folded_Diff_Op_Amp_Layout_0.BD.n205 0.00998204
R20728 Folded_Diff_Op_Amp_Layout_0.BD.n203 Folded_Diff_Op_Amp_Layout_0.BD.n0 0.00983809
R20729 Folded_Diff_Op_Amp_Layout_0.BD.n33 Folded_Diff_Op_Amp_Layout_0.BD.n32 0.00860784
R20730 Folded_Diff_Op_Amp_Layout_0.BD.n177 Folded_Diff_Op_Amp_Layout_0.BD.n176 0.00860784
R20731 Folded_Diff_Op_Amp_Layout_0.BD.n97 Folded_Diff_Op_Amp_Layout_0.BD.n96 0.00860784
R20732 Folded_Diff_Op_Amp_Layout_0.BD.n61 Folded_Diff_Op_Amp_Layout_0.BD.n60 0.00860784
R20733 Folded_Diff_Op_Amp_Layout_0.BD.n37 Folded_Diff_Op_Amp_Layout_0.BD.n36 0.00773989
R20734 Folded_Diff_Op_Amp_Layout_0.BD.n159 Folded_Diff_Op_Amp_Layout_0.BD.n158 0.00773989
R20735 Folded_Diff_Op_Amp_Layout_0.BD.n36 Folded_Diff_Op_Amp_Layout_0.BD.n35 0.00773989
R20736 Folded_Diff_Op_Amp_Layout_0.BD.n158 Folded_Diff_Op_Amp_Layout_0.BD.n157 0.00773989
R20737 Folded_Diff_Op_Amp_Layout_0.BD.n102 Folded_Diff_Op_Amp_Layout_0.BD.n100 0.00605114
R20738 Folded_Diff_Op_Amp_Layout_0.BD.n66 Folded_Diff_Op_Amp_Layout_0.BD.n64 0.00605114
R20739 Folded_Diff_Op_Amp_Layout_0.BD.n185 Folded_Diff_Op_Amp_Layout_0.BD.n3 0.00582347
R20740 Folded_Diff_Op_Amp_Layout_0.BD.n38 Folded_Diff_Op_Amp_Layout_0.BD.n37 0.00582347
R20741 Folded_Diff_Op_Amp_Layout_0.BD.n115 Folded_Diff_Op_Amp_Layout_0.BD.n113 0.00549102
R20742 Folded_Diff_Op_Amp_Layout_0.BD.n185 Folded_Diff_Op_Amp_Layout_0.BD.n184 0.00549102
R20743 Folded_Diff_Op_Amp_Layout_0.BD.n157 Folded_Diff_Op_Amp_Layout_0.BD.n116 0.00549102
R20744 Folded_Diff_Op_Amp_Layout_0.BD.n102 Folded_Diff_Op_Amp_Layout_0.BD.n101 0.005061
R20745 Folded_Diff_Op_Amp_Layout_0.BD.n66 Folded_Diff_Op_Amp_Layout_0.BD.n65 0.005061
R20746 Folded_Diff_Op_Amp_Layout_0.OUT2.t44 Folded_Diff_Op_Amp_Layout_0.OUT2.t88 122.014
R20747 Folded_Diff_Op_Amp_Layout_0.OUT2.t90 Folded_Diff_Op_Amp_Layout_0.OUT2.t70 122.014
R20748 Folded_Diff_Op_Amp_Layout_0.OUT2.t61 Folded_Diff_Op_Amp_Layout_0.OUT2.t50 122.014
R20749 Folded_Diff_Op_Amp_Layout_0.OUT2.t66 Folded_Diff_Op_Amp_Layout_0.OUT2.t97 122.014
R20750 Folded_Diff_Op_Amp_Layout_0.OUT2.t81 Folded_Diff_Op_Amp_Layout_0.OUT2.t101 122.014
R20751 Folded_Diff_Op_Amp_Layout_0.OUT2.t86 Folded_Diff_Op_Amp_Layout_0.OUT2.t68 122.014
R20752 Folded_Diff_Op_Amp_Layout_0.OUT2.t105 Folded_Diff_Op_Amp_Layout_0.OUT2.t72 122.014
R20753 Folded_Diff_Op_Amp_Layout_0.OUT2.t52 Folded_Diff_Op_Amp_Layout_0.OUT2.t92 122.014
R20754 Folded_Diff_Op_Amp_Layout_0.OUT2.t47 Folded_Diff_Op_Amp_Layout_0.OUT2.t59 122.014
R20755 Folded_Diff_Op_Amp_Layout_0.OUT2.t41 Folded_Diff_Op_Amp_Layout_0.OUT2.t94 122.014
R20756 Folded_Diff_Op_Amp_Layout_0.OUT2.t63 Folded_Diff_Op_Amp_Layout_0.OUT2.t95 122.014
R20757 Folded_Diff_Op_Amp_Layout_0.OUT2.t58 Folded_Diff_Op_Amp_Layout_0.OUT2.t102 122.014
R20758 Folded_Diff_Op_Amp_Layout_0.OUT2.n57 Folded_Diff_Op_Amp_Layout_0.OUT2.t67 63.548
R20759 Folded_Diff_Op_Amp_Layout_0.OUT2.n77 Folded_Diff_Op_Amp_Layout_0.OUT2.t75 63.548
R20760 Folded_Diff_Op_Amp_Layout_0.OUT2.n49 Folded_Diff_Op_Amp_Layout_0.OUT2.t57 63.548
R20761 Folded_Diff_Op_Amp_Layout_0.OUT2.n69 Folded_Diff_Op_Amp_Layout_0.OUT2.t37 63.548
R20762 Folded_Diff_Op_Amp_Layout_0.OUT2.n35 Folded_Diff_Op_Amp_Layout_0.OUT2.t77 63.548
R20763 Folded_Diff_Op_Amp_Layout_0.OUT2.n28 Folded_Diff_Op_Amp_Layout_0.OUT2.t49 63.548
R20764 Folded_Diff_Op_Amp_Layout_0.OUT2.n41 Folded_Diff_Op_Amp_Layout_0.OUT2.t82 62.5719
R20765 Folded_Diff_Op_Amp_Layout_0.OUT2.n42 Folded_Diff_Op_Amp_Layout_0.OUT2.t106 62.5719
R20766 Folded_Diff_Op_Amp_Layout_0.OUT2.n43 Folded_Diff_Op_Amp_Layout_0.OUT2.t98 62.5719
R20767 Folded_Diff_Op_Amp_Layout_0.OUT2.n44 Folded_Diff_Op_Amp_Layout_0.OUT2.t56 62.5719
R20768 Folded_Diff_Op_Amp_Layout_0.OUT2.n60 Folded_Diff_Op_Amp_Layout_0.OUT2.t90 62.5719
R20769 Folded_Diff_Op_Amp_Layout_0.OUT2.n58 Folded_Diff_Op_Amp_Layout_0.OUT2.t89 62.5719
R20770 Folded_Diff_Op_Amp_Layout_0.OUT2.n56 Folded_Diff_Op_Amp_Layout_0.OUT2.t66 62.5719
R20771 Folded_Diff_Op_Amp_Layout_0.OUT2.n74 Folded_Diff_Op_Amp_Layout_0.OUT2.t86 62.5719
R20772 Folded_Diff_Op_Amp_Layout_0.OUT2.n75 Folded_Diff_Op_Amp_Layout_0.OUT2.t107 62.5719
R20773 Folded_Diff_Op_Amp_Layout_0.OUT2.n76 Folded_Diff_Op_Amp_Layout_0.OUT2.t52 62.5719
R20774 Folded_Diff_Op_Amp_Layout_0.OUT2.n52 Folded_Diff_Op_Amp_Layout_0.OUT2.t73 62.5719
R20775 Folded_Diff_Op_Amp_Layout_0.OUT2.n50 Folded_Diff_Op_Amp_Layout_0.OUT2.t64 62.5719
R20776 Folded_Diff_Op_Amp_Layout_0.OUT2.n48 Folded_Diff_Op_Amp_Layout_0.OUT2.t103 62.5719
R20777 Folded_Diff_Op_Amp_Layout_0.OUT2.n66 Folded_Diff_Op_Amp_Layout_0.OUT2.t71 62.5719
R20778 Folded_Diff_Op_Amp_Layout_0.OUT2.n67 Folded_Diff_Op_Amp_Layout_0.OUT2.t42 62.5719
R20779 Folded_Diff_Op_Amp_Layout_0.OUT2.n68 Folded_Diff_Op_Amp_Layout_0.OUT2.t96 62.5719
R20780 Folded_Diff_Op_Amp_Layout_0.OUT2.n45 Folded_Diff_Op_Amp_Layout_0.OUT2.t60 62.5719
R20781 Folded_Diff_Op_Amp_Layout_0.OUT2.n46 Folded_Diff_Op_Amp_Layout_0.OUT2.t46 62.5719
R20782 Folded_Diff_Op_Amp_Layout_0.OUT2.n38 Folded_Diff_Op_Amp_Layout_0.OUT2.t41 62.5719
R20783 Folded_Diff_Op_Amp_Layout_0.OUT2.n36 Folded_Diff_Op_Amp_Layout_0.OUT2.t91 62.5719
R20784 Folded_Diff_Op_Amp_Layout_0.OUT2.n34 Folded_Diff_Op_Amp_Layout_0.OUT2.t58 62.5719
R20785 Folded_Diff_Op_Amp_Layout_0.OUT2.n31 Folded_Diff_Op_Amp_Layout_0.OUT2.t99 62.5719
R20786 Folded_Diff_Op_Amp_Layout_0.OUT2.n29 Folded_Diff_Op_Amp_Layout_0.OUT2.t48 62.5719
R20787 Folded_Diff_Op_Amp_Layout_0.OUT2.n27 Folded_Diff_Op_Amp_Layout_0.OUT2.t39 62.5719
R20788 Folded_Diff_Op_Amp_Layout_0.OUT2.n80 Folded_Diff_Op_Amp_Layout_0.OUT2.t84 61.8074
R20789 Folded_Diff_Op_Amp_Layout_0.OUT2.n72 Folded_Diff_Op_Amp_Layout_0.OUT2.t62 61.8074
R20790 Folded_Diff_Op_Amp_Layout_0.OUT2.n62 Folded_Diff_Op_Amp_Layout_0.OUT2.t80 61.8072
R20791 Folded_Diff_Op_Amp_Layout_0.OUT2.n54 Folded_Diff_Op_Amp_Layout_0.OUT2.t76 61.8072
R20792 Folded_Diff_Op_Amp_Layout_0.OUT2.n40 Folded_Diff_Op_Amp_Layout_0.OUT2.t85 61.8072
R20793 Folded_Diff_Op_Amp_Layout_0.OUT2.n33 Folded_Diff_Op_Amp_Layout_0.OUT2.t51 61.8072
R20794 Folded_Diff_Op_Amp_Layout_0.OUT2.n41 Folded_Diff_Op_Amp_Layout_0.OUT2.t87 41.7148
R20795 Folded_Diff_Op_Amp_Layout_0.OUT2.n42 Folded_Diff_Op_Amp_Layout_0.OUT2.t43 41.7148
R20796 Folded_Diff_Op_Amp_Layout_0.OUT2.n43 Folded_Diff_Op_Amp_Layout_0.OUT2.t74 41.7148
R20797 Folded_Diff_Op_Amp_Layout_0.OUT2.n44 Folded_Diff_Op_Amp_Layout_0.OUT2.t54 41.7148
R20798 Folded_Diff_Op_Amp_Layout_0.OUT2.n60 Folded_Diff_Op_Amp_Layout_0.OUT2.t44 41.7148
R20799 Folded_Diff_Op_Amp_Layout_0.OUT2.n58 Folded_Diff_Op_Amp_Layout_0.OUT2.t40 41.7148
R20800 Folded_Diff_Op_Amp_Layout_0.OUT2.n56 Folded_Diff_Op_Amp_Layout_0.OUT2.t61 41.7148
R20801 Folded_Diff_Op_Amp_Layout_0.OUT2.n74 Folded_Diff_Op_Amp_Layout_0.OUT2.t81 41.7148
R20802 Folded_Diff_Op_Amp_Layout_0.OUT2.n75 Folded_Diff_Op_Amp_Layout_0.OUT2.t104 41.7148
R20803 Folded_Diff_Op_Amp_Layout_0.OUT2.n76 Folded_Diff_Op_Amp_Layout_0.OUT2.t105 41.7148
R20804 Folded_Diff_Op_Amp_Layout_0.OUT2.n52 Folded_Diff_Op_Amp_Layout_0.OUT2.t93 41.7148
R20805 Folded_Diff_Op_Amp_Layout_0.OUT2.n50 Folded_Diff_Op_Amp_Layout_0.OUT2.t79 41.7148
R20806 Folded_Diff_Op_Amp_Layout_0.OUT2.n48 Folded_Diff_Op_Amp_Layout_0.OUT2.t53 41.7148
R20807 Folded_Diff_Op_Amp_Layout_0.OUT2.n66 Folded_Diff_Op_Amp_Layout_0.OUT2.t36 41.7148
R20808 Folded_Diff_Op_Amp_Layout_0.OUT2.n67 Folded_Diff_Op_Amp_Layout_0.OUT2.t69 41.7148
R20809 Folded_Diff_Op_Amp_Layout_0.OUT2.n68 Folded_Diff_Op_Amp_Layout_0.OUT2.t78 41.7148
R20810 Folded_Diff_Op_Amp_Layout_0.OUT2.n45 Folded_Diff_Op_Amp_Layout_0.OUT2.t83 41.7148
R20811 Folded_Diff_Op_Amp_Layout_0.OUT2.n46 Folded_Diff_Op_Amp_Layout_0.OUT2.t38 41.7148
R20812 Folded_Diff_Op_Amp_Layout_0.OUT2.n38 Folded_Diff_Op_Amp_Layout_0.OUT2.t47 41.7148
R20813 Folded_Diff_Op_Amp_Layout_0.OUT2.n36 Folded_Diff_Op_Amp_Layout_0.OUT2.t45 41.7148
R20814 Folded_Diff_Op_Amp_Layout_0.OUT2.n34 Folded_Diff_Op_Amp_Layout_0.OUT2.t63 41.7148
R20815 Folded_Diff_Op_Amp_Layout_0.OUT2.n31 Folded_Diff_Op_Amp_Layout_0.OUT2.t65 41.7148
R20816 Folded_Diff_Op_Amp_Layout_0.OUT2.n29 Folded_Diff_Op_Amp_Layout_0.OUT2.t55 41.7148
R20817 Folded_Diff_Op_Amp_Layout_0.OUT2.n27 Folded_Diff_Op_Amp_Layout_0.OUT2.t100 41.7148
R20818 Folded_Diff_Op_Amp_Layout_0.OUT2.n47 Folded_Diff_Op_Amp_Layout_0.OUT2.n46 17.2118
R20819 Folded_Diff_Op_Amp_Layout_0.OUT2.n61 Folded_Diff_Op_Amp_Layout_0.OUT2.n60 15.9934
R20820 Folded_Diff_Op_Amp_Layout_0.OUT2.n57 Folded_Diff_Op_Amp_Layout_0.OUT2.n56 15.9934
R20821 Folded_Diff_Op_Amp_Layout_0.OUT2.n79 Folded_Diff_Op_Amp_Layout_0.OUT2.n74 15.9934
R20822 Folded_Diff_Op_Amp_Layout_0.OUT2.n77 Folded_Diff_Op_Amp_Layout_0.OUT2.n76 15.9934
R20823 Folded_Diff_Op_Amp_Layout_0.OUT2.n53 Folded_Diff_Op_Amp_Layout_0.OUT2.n52 15.9934
R20824 Folded_Diff_Op_Amp_Layout_0.OUT2.n49 Folded_Diff_Op_Amp_Layout_0.OUT2.n48 15.9934
R20825 Folded_Diff_Op_Amp_Layout_0.OUT2.n71 Folded_Diff_Op_Amp_Layout_0.OUT2.n66 15.9934
R20826 Folded_Diff_Op_Amp_Layout_0.OUT2.n69 Folded_Diff_Op_Amp_Layout_0.OUT2.n68 15.9934
R20827 Folded_Diff_Op_Amp_Layout_0.OUT2.n39 Folded_Diff_Op_Amp_Layout_0.OUT2.n38 15.9934
R20828 Folded_Diff_Op_Amp_Layout_0.OUT2.n35 Folded_Diff_Op_Amp_Layout_0.OUT2.n34 15.9934
R20829 Folded_Diff_Op_Amp_Layout_0.OUT2.n32 Folded_Diff_Op_Amp_Layout_0.OUT2.n31 15.9934
R20830 Folded_Diff_Op_Amp_Layout_0.OUT2.n28 Folded_Diff_Op_Amp_Layout_0.OUT2.n27 15.9934
R20831 Folded_Diff_Op_Amp_Layout_0.OUT2.n84 Folded_Diff_Op_Amp_Layout_0.OUT2.n44 14.8788
R20832 Folded_Diff_Op_Amp_Layout_0.OUT2.n86 Folded_Diff_Op_Amp_Layout_0.OUT2.n42 14.8788
R20833 Folded_Diff_Op_Amp_Layout_0.OUT2.n47 Folded_Diff_Op_Amp_Layout_0.OUT2.n45 14.8786
R20834 Folded_Diff_Op_Amp_Layout_0.OUT2.n85 Folded_Diff_Op_Amp_Layout_0.OUT2.n43 14.8786
R20835 Folded_Diff_Op_Amp_Layout_0.OUT2.n87 Folded_Diff_Op_Amp_Layout_0.OUT2.n41 14.8786
R20836 Folded_Diff_Op_Amp_Layout_0.OUT2.n59 Folded_Diff_Op_Amp_Layout_0.OUT2.n58 13.9076
R20837 Folded_Diff_Op_Amp_Layout_0.OUT2.n78 Folded_Diff_Op_Amp_Layout_0.OUT2.n75 13.9076
R20838 Folded_Diff_Op_Amp_Layout_0.OUT2.n51 Folded_Diff_Op_Amp_Layout_0.OUT2.n50 13.9076
R20839 Folded_Diff_Op_Amp_Layout_0.OUT2.n70 Folded_Diff_Op_Amp_Layout_0.OUT2.n67 13.9076
R20840 Folded_Diff_Op_Amp_Layout_0.OUT2.n37 Folded_Diff_Op_Amp_Layout_0.OUT2.n36 13.9076
R20841 Folded_Diff_Op_Amp_Layout_0.OUT2.n30 Folded_Diff_Op_Amp_Layout_0.OUT2.n29 13.9076
R20842 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.OUT2.n89 8.55615
R20843 Folded_Diff_Op_Amp_Layout_0.OUT2.n86 Folded_Diff_Op_Amp_Layout_0.OUT2.n85 8.51465
R20844 Folded_Diff_Op_Amp_Layout_0.OUT2.n88 Folded_Diff_Op_Amp_Layout_0.OUT2.n87 7.59746
R20845 Folded_Diff_Op_Amp_Layout_0.OUT2.n23 Folded_Diff_Op_Amp_Layout_0.OUT2.t19 6.49823
R20846 Folded_Diff_Op_Amp_Layout_0.OUT2.n23 Folded_Diff_Op_Amp_Layout_0.OUT2.t14 6.4095
R20847 Folded_Diff_Op_Amp_Layout_0.OUT2.n82 Folded_Diff_Op_Amp_Layout_0.OUT2.n73 5.57576
R20848 Folded_Diff_Op_Amp_Layout_0.OUT2.n64 Folded_Diff_Op_Amp_Layout_0.OUT2.n55 5.57576
R20849 Folded_Diff_Op_Amp_Layout_0.OUT2.n89 Folded_Diff_Op_Amp_Layout_0.OUT2.n88 5.57576
R20850 Folded_Diff_Op_Amp_Layout_0.OUT2.n102 Folded_Diff_Op_Amp_Layout_0.OUT2.n101 5.40577
R20851 Folded_Diff_Op_Amp_Layout_0.OUT2.n99 Folded_Diff_Op_Amp_Layout_0.OUT2.t16 5.40577
R20852 Folded_Diff_Op_Amp_Layout_0.OUT2.n98 Folded_Diff_Op_Amp_Layout_0.OUT2.n97 5.40577
R20853 Folded_Diff_Op_Amp_Layout_0.OUT2.n88 Folded_Diff_Op_Amp_Layout_0.OUT2.n40 5.19114
R20854 Folded_Diff_Op_Amp_Layout_0.OUT2.n111 Folded_Diff_Op_Amp_Layout_0.OUT2.t6 5.08295
R20855 Folded_Diff_Op_Amp_Layout_0.OUT2.n93 Folded_Diff_Op_Amp_Layout_0.OUT2.t7 4.9949
R20856 Folded_Diff_Op_Amp_Layout_0.OUT2.n208 Folded_Diff_Op_Amp_Layout_0.OUT2.t3 4.9949
R20857 Folded_Diff_Op_Amp_Layout_0.OUT2.n140 Folded_Diff_Op_Amp_Layout_0.OUT2.n139 4.66184
R20858 Folded_Diff_Op_Amp_Layout_0.OUT2.n118 Folded_Diff_Op_Amp_Layout_0.OUT2.t28 4.66184
R20859 Folded_Diff_Op_Amp_Layout_0.OUT2.n83 Folded_Diff_Op_Amp_Layout_0.OUT2.n82 4.46734
R20860 Folded_Diff_Op_Amp_Layout_0.OUT2.n65 Folded_Diff_Op_Amp_Layout_0.OUT2.n64 4.46734
R20861 Folded_Diff_Op_Amp_Layout_0.OUT2.n95 Folded_Diff_Op_Amp_Layout_0.OUT2.n91 4.36882
R20862 Folded_Diff_Op_Amp_Layout_0.OUT2.n94 Folded_Diff_Op_Amp_Layout_0.OUT2.t9 4.36882
R20863 Folded_Diff_Op_Amp_Layout_0.OUT2.n93 Folded_Diff_Op_Amp_Layout_0.OUT2.n92 4.36882
R20864 Folded_Diff_Op_Amp_Layout_0.OUT2.n206 Folded_Diff_Op_Amp_Layout_0.OUT2.t2 4.36882
R20865 Folded_Diff_Op_Amp_Layout_0.OUT2.n208 Folded_Diff_Op_Amp_Layout_0.OUT2.n207 4.36882
R20866 Folded_Diff_Op_Amp_Layout_0.OUT2.n168 Folded_Diff_Op_Amp_Layout_0.OUT2.n167 4.10662
R20867 Folded_Diff_Op_Amp_Layout_0.OUT2.n133 Folded_Diff_Op_Amp_Layout_0.OUT2.n132 4.05775
R20868 Folded_Diff_Op_Amp_Layout_0.OUT2.n102 Folded_Diff_Op_Amp_Layout_0.OUT2.n100 3.71925
R20869 Folded_Diff_Op_Amp_Layout_0.OUT2.n99 Folded_Diff_Op_Amp_Layout_0.OUT2.t1 3.71925
R20870 Folded_Diff_Op_Amp_Layout_0.OUT2.n98 Folded_Diff_Op_Amp_Layout_0.OUT2.n96 3.71925
R20871 Folded_Diff_Op_Amp_Layout_0.OUT2.n65 Folded_Diff_Op_Amp_Layout_0.OUT2.n47 3.13062
R20872 Folded_Diff_Op_Amp_Layout_0.OUT2.n84 Folded_Diff_Op_Amp_Layout_0.OUT2.n83 3.12979
R20873 Folded_Diff_Op_Amp_Layout_0.OUT2.n55 Folded_Diff_Op_Amp_Layout_0.OUT2.n54 2.94114
R20874 Folded_Diff_Op_Amp_Layout_0.OUT2.n63 Folded_Diff_Op_Amp_Layout_0.OUT2.n62 2.94114
R20875 Folded_Diff_Op_Amp_Layout_0.OUT2.n73 Folded_Diff_Op_Amp_Layout_0.OUT2.n72 2.94095
R20876 Folded_Diff_Op_Amp_Layout_0.OUT2.n81 Folded_Diff_Op_Amp_Layout_0.OUT2.n80 2.94095
R20877 Folded_Diff_Op_Amp_Layout_0.OUT2.n89 Folded_Diff_Op_Amp_Layout_0.OUT2.n33 2.94051
R20878 Folded_Diff_Op_Amp_Layout_0.OUT2.n154 Folded_Diff_Op_Amp_Layout_0.OUT2.n200 2.63228
R20879 Folded_Diff_Op_Amp_Layout_0.OUT2.n22 Folded_Diff_Op_Amp_Layout_0.OUT2.t15 2.4095
R20880 Folded_Diff_Op_Amp_Layout_0.OUT2.n82 Folded_Diff_Op_Amp_Layout_0.OUT2.n81 2.2505
R20881 Folded_Diff_Op_Amp_Layout_0.OUT2.n64 Folded_Diff_Op_Amp_Layout_0.OUT2.n63 2.2505
R20882 Folded_Diff_Op_Amp_Layout_0.OUT2.n6 Folded_Diff_Op_Amp_Layout_0.OUT2.n5 2.24736
R20883 Folded_Diff_Op_Amp_Layout_0.OUT2.n25 Folded_Diff_Op_Amp_Layout_0.OUT2.n22 2.11382
R20884 Folded_Diff_Op_Amp_Layout_0.OUT2.n103 Folded_Diff_Op_Amp_Layout_0.OUT2.n102 1.77702
R20885 Folded_Diff_Op_Amp_Layout_0.OUT2.n202 Folded_Diff_Op_Amp_Layout_0.OUT2.n204 1.76122
R20886 Folded_Diff_Op_Amp_Layout_0.OUT2.n18 Folded_Diff_Op_Amp_Layout_0.OUT2.n198 1.52544
R20887 Folded_Diff_Op_Amp_Layout_0.OUT2.n171 Folded_Diff_Op_Amp_Layout_0.OUT2.n157 1.48953
R20888 Folded_Diff_Op_Amp_Layout_0.OUT2.n189 Folded_Diff_Op_Amp_Layout_0.OUT2.n188 1.48953
R20889 Folded_Diff_Op_Amp_Layout_0.OUT2.n191 Folded_Diff_Op_Amp_Layout_0.OUT2.n152 1.48953
R20890 Folded_Diff_Op_Amp_Layout_0.OUT2.n192 Folded_Diff_Op_Amp_Layout_0.OUT2.n151 1.48953
R20891 Folded_Diff_Op_Amp_Layout_0.OUT2.n154 Folded_Diff_Op_Amp_Layout_0.OUT2.n153 1.48107
R20892 Folded_Diff_Op_Amp_Layout_0.OUT2.n202 Folded_Diff_Op_Amp_Layout_0.OUT2.n206 1.34243
R20893 Folded_Diff_Op_Amp_Layout_0.OUT2.n165 Folded_Diff_Op_Amp_Layout_0.OUT2.n21 1.35922
R20894 Folded_Diff_Op_Amp_Layout_0.OUT2.n145 Folded_Diff_Op_Amp_Layout_0.OUT2.n144 1.30811
R20895 Folded_Diff_Op_Amp_Layout_0.OUT2.n122 Folded_Diff_Op_Amp_Layout_0.OUT2.n121 1.30811
R20896 Folded_Diff_Op_Amp_Layout_0.OUT2.n110 Folded_Diff_Op_Amp_Layout_0.OUT2.n109 1.28725
R20897 Folded_Diff_Op_Amp_Layout_0.OUT2.n184 Folded_Diff_Op_Amp_Layout_0.OUT2.n183 1.19489
R20898 Folded_Diff_Op_Amp_Layout_0.OUT2.n85 Folded_Diff_Op_Amp_Layout_0.OUT2.n84 1.18503
R20899 Folded_Diff_Op_Amp_Layout_0.OUT2.n87 Folded_Diff_Op_Amp_Layout_0.OUT2.n86 1.18503
R20900 Folded_Diff_Op_Amp_Layout_0.OUT2.n176 Folded_Diff_Op_Amp_Layout_0.OUT2.n175 1.17841
R20901 Folded_Diff_Op_Amp_Layout_0.OUT2.n130 Folded_Diff_Op_Amp_Layout_0.OUT2.n129 1.16567
R20902 Folded_Diff_Op_Amp_Layout_0.OUT2.n15 Folded_Diff_Op_Amp_Layout_0.OUT2.n14 1.16484
R20903 Folded_Diff_Op_Amp_Layout_0.OUT2.n4 Folded_Diff_Op_Amp_Layout_0.OUT2.n3 1.1643
R20904 Folded_Diff_Op_Amp_Layout_0.OUT2.n146 Folded_Diff_Op_Amp_Layout_0.OUT2.n145 1.14175
R20905 Folded_Diff_Op_Amp_Layout_0.OUT2.n123 Folded_Diff_Op_Amp_Layout_0.OUT2.n122 1.14175
R20906 Folded_Diff_Op_Amp_Layout_0.OUT2.n94 Folded_Diff_Op_Amp_Layout_0.OUT2.n93 1.12746
R20907 Folded_Diff_Op_Amp_Layout_0.OUT2.n206 Folded_Diff_Op_Amp_Layout_0.OUT2.n208 1.12746
R20908 Folded_Diff_Op_Amp_Layout_0.OUT2.n142 Folded_Diff_Op_Amp_Layout_0.OUT2.n141 1.1255
R20909 Folded_Diff_Op_Amp_Layout_0.OUT2.n120 Folded_Diff_Op_Amp_Layout_0.OUT2.n119 1.1255
R20910 Folded_Diff_Op_Amp_Layout_0.OUT2.n108 Folded_Diff_Op_Amp_Layout_0.OUT2.n107 1.1255
R20911 Folded_Diff_Op_Amp_Layout_0.OUT2.n113 Folded_Diff_Op_Amp_Layout_0.OUT2.n112 1.1255
R20912 Folded_Diff_Op_Amp_Layout_0.OUT2.n135 Folded_Diff_Op_Amp_Layout_0.OUT2.n134 1.1255
R20913 Folded_Diff_Op_Amp_Layout_0.OUT2.n26 Folded_Diff_Op_Amp_Layout_0.OUT2.n21 1.12145
R20914 Folded_Diff_Op_Amp_Layout_0.OUT2.n167 Folded_Diff_Op_Amp_Layout_0.OUT2.n166 1.1318
R20915 Folded_Diff_Op_Amp_Layout_0.OUT2.n17 Folded_Diff_Op_Amp_Layout_0.OUT2.n16 1.10737
R20916 Folded_Diff_Op_Amp_Layout_0.OUT2.n3 Folded_Diff_Op_Amp_Layout_0.OUT2.n2 1.00262
R20917 Folded_Diff_Op_Amp_Layout_0.OUT2.n14 Folded_Diff_Op_Amp_Layout_0.OUT2.n13 1.00232
R20918 Folded_Diff_Op_Amp_Layout_0.OUT2.n129 Folded_Diff_Op_Amp_Layout_0.OUT2.n128 0.995607
R20919 Folded_Diff_Op_Amp_Layout_0.OUT2.n194 Folded_Diff_Op_Amp_Layout_0.OUT2.n117 0.978961
R20920 Folded_Diff_Op_Amp_Layout_0.OUT2.n18 Folded_Diff_Op_Amp_Layout_0.OUT2.n90 0.917563
R20921 Folded_Diff_Op_Amp_Layout_0.OUT2.n6 Folded_Diff_Op_Amp_Layout_0.OUT2.n4 0.911329
R20922 Folded_Diff_Op_Amp_Layout_0.OUT2.n105 Folded_Diff_Op_Amp_Layout_0.OUT2.n104 0.877022
R20923 Folded_Diff_Op_Amp_Layout_0.OUT2.n195 Folded_Diff_Op_Amp_Layout_0.OUT2.n194 0.857314
R20924 Folded_Diff_Op_Amp_Layout_0.OUT2.n183 Folded_Diff_Op_Amp_Layout_0.OUT2.n182 0.824494
R20925 Folded_Diff_Op_Amp_Layout_0.OUT2.n175 Folded_Diff_Op_Amp_Layout_0.OUT2.n174 0.824494
R20926 Folded_Diff_Op_Amp_Layout_0.OUT2.n171 Folded_Diff_Op_Amp_Layout_0.OUT2.n170 4.05954
R20927 Folded_Diff_Op_Amp_Layout_0.OUT2.n186 Folded_Diff_Op_Amp_Layout_0.OUT2.n185 0.743266
R20928 Folded_Diff_Op_Amp_Layout_0.OUT2.n188 Folded_Diff_Op_Amp_Layout_0.OUT2.n187 0.72825
R20929 Folded_Diff_Op_Amp_Layout_0.OUT2.n138 Folded_Diff_Op_Amp_Layout_0.OUT2.n136 0.727104
R20930 Folded_Diff_Op_Amp_Layout_0.OUT2.n103 Folded_Diff_Op_Amp_Layout_0.OUT2.n99 0.650065
R20931 Folded_Diff_Op_Amp_Layout_0.OUT2.n104 Folded_Diff_Op_Amp_Layout_0.OUT2.n98 0.650065
R20932 Folded_Diff_Op_Amp_Layout_0.OUT2.n148 Folded_Diff_Op_Amp_Layout_0.OUT2.n147 0.631966
R20933 Folded_Diff_Op_Amp_Layout_0.OUT2.n95 Folded_Diff_Op_Amp_Layout_0.OUT2.n94 0.626587
R20934 Folded_Diff_Op_Amp_Layout_0.OUT2.n104 Folded_Diff_Op_Amp_Layout_0.OUT2.n103 0.626587
R20935 Folded_Diff_Op_Amp_Layout_0.OUT2.n59 Folded_Diff_Op_Amp_Layout_0.OUT2.n57 0.626587
R20936 Folded_Diff_Op_Amp_Layout_0.OUT2.n61 Folded_Diff_Op_Amp_Layout_0.OUT2.n59 0.626587
R20937 Folded_Diff_Op_Amp_Layout_0.OUT2.n79 Folded_Diff_Op_Amp_Layout_0.OUT2.n78 0.626587
R20938 Folded_Diff_Op_Amp_Layout_0.OUT2.n78 Folded_Diff_Op_Amp_Layout_0.OUT2.n77 0.626587
R20939 Folded_Diff_Op_Amp_Layout_0.OUT2.n51 Folded_Diff_Op_Amp_Layout_0.OUT2.n49 0.626587
R20940 Folded_Diff_Op_Amp_Layout_0.OUT2.n53 Folded_Diff_Op_Amp_Layout_0.OUT2.n51 0.626587
R20941 Folded_Diff_Op_Amp_Layout_0.OUT2.n71 Folded_Diff_Op_Amp_Layout_0.OUT2.n70 0.626587
R20942 Folded_Diff_Op_Amp_Layout_0.OUT2.n70 Folded_Diff_Op_Amp_Layout_0.OUT2.n69 0.626587
R20943 Folded_Diff_Op_Amp_Layout_0.OUT2.n37 Folded_Diff_Op_Amp_Layout_0.OUT2.n35 0.626587
R20944 Folded_Diff_Op_Amp_Layout_0.OUT2.n39 Folded_Diff_Op_Amp_Layout_0.OUT2.n37 0.626587
R20945 Folded_Diff_Op_Amp_Layout_0.OUT2.n30 Folded_Diff_Op_Amp_Layout_0.OUT2.n28 0.626587
R20946 Folded_Diff_Op_Amp_Layout_0.OUT2.n32 Folded_Diff_Op_Amp_Layout_0.OUT2.n30 0.626587
R20947 Folded_Diff_Op_Amp_Layout_0.OUT2.n126 Folded_Diff_Op_Amp_Layout_0.OUT2.n124 0.616779
R20948 Folded_Diff_Op_Amp_Layout_0.OUT2.n116 Folded_Diff_Op_Amp_Layout_0.OUT2.n114 0.616779
R20949 Folded_Diff_Op_Amp_Layout_0.OUT2.n179 Folded_Diff_Op_Amp_Layout_0.OUT2.n177 0.616779
R20950 Folded_Diff_Op_Amp_Layout_0.OUT2.n144 Folded_Diff_Op_Amp_Layout_0.OUT2.n143 0.58197
R20951 Folded_Diff_Op_Amp_Layout_0.OUT2.n121 Folded_Diff_Op_Amp_Layout_0.OUT2.t30 0.58197
R20952 Folded_Diff_Op_Amp_Layout_0.OUT2.n13 Folded_Diff_Op_Amp_Layout_0.OUT2.t27 0.58197
R20953 Folded_Diff_Op_Amp_Layout_0.OUT2.n13 Folded_Diff_Op_Amp_Layout_0.OUT2.n12 0.58197
R20954 Folded_Diff_Op_Amp_Layout_0.OUT2.n2 Folded_Diff_Op_Amp_Layout_0.OUT2.t26 0.58197
R20955 Folded_Diff_Op_Amp_Layout_0.OUT2.n2 Folded_Diff_Op_Amp_Layout_0.OUT2.n1 0.58197
R20956 Folded_Diff_Op_Amp_Layout_0.OUT2.n182 Folded_Diff_Op_Amp_Layout_0.OUT2.t25 0.58197
R20957 Folded_Diff_Op_Amp_Layout_0.OUT2.n182 Folded_Diff_Op_Amp_Layout_0.OUT2.n181 0.58197
R20958 Folded_Diff_Op_Amp_Layout_0.OUT2.n174 Folded_Diff_Op_Amp_Layout_0.OUT2.t31 0.58197
R20959 Folded_Diff_Op_Amp_Layout_0.OUT2.n174 Folded_Diff_Op_Amp_Layout_0.OUT2.n173 0.58197
R20960 Folded_Diff_Op_Amp_Layout_0.OUT2.n132 Folded_Diff_Op_Amp_Layout_0.OUT2.t29 0.58197
R20961 Folded_Diff_Op_Amp_Layout_0.OUT2.n132 Folded_Diff_Op_Amp_Layout_0.OUT2.n131 0.58197
R20962 Folded_Diff_Op_Amp_Layout_0.OUT2.n128 Folded_Diff_Op_Amp_Layout_0.OUT2.t32 0.58197
R20963 Folded_Diff_Op_Amp_Layout_0.OUT2.n128 Folded_Diff_Op_Amp_Layout_0.OUT2.n127 0.58197
R20964 Folded_Diff_Op_Amp_Layout_0.OUT2.n109 Folded_Diff_Op_Amp_Layout_0.OUT2.t12 0.56925
R20965 Folded_Diff_Op_Amp_Layout_0.OUT2.n204 Folded_Diff_Op_Amp_Layout_0.OUT2.n205 0.56925
R20966 Folded_Diff_Op_Amp_Layout_0.OUT2.n106 Folded_Diff_Op_Amp_Layout_0.OUT2.n105 0.532674
R20967 Folded_Diff_Op_Amp_Layout_0.OUT2.n191 Folded_Diff_Op_Amp_Layout_0.OUT2.n190 0.527875
R20968 Folded_Diff_Op_Amp_Layout_0.OUT2.n156 Folded_Diff_Op_Amp_Layout_0.OUT2.n155 0.4875
R20969 Folded_Diff_Op_Amp_Layout_0.OUT2.n151 Folded_Diff_Op_Amp_Layout_0.OUT2.n150 0.47625
R20970 Folded_Diff_Op_Amp_Layout_0.OUT2.n83 Folded_Diff_Op_Amp_Layout_0.OUT2.n65 0.475368
R20971 Folded_Diff_Op_Amp_Layout_0.OUT2.n8 Folded_Diff_Op_Amp_Layout_0.OUT2.n7 0.474125
R20972 Folded_Diff_Op_Amp_Layout_0.OUT2.n178 Folded_Diff_Op_Amp_Layout_0.OUT2.n186 0.474125
R20973 Folded_Diff_Op_Amp_Layout_0.OUT2.n137 Folded_Diff_Op_Amp_Layout_0.OUT2.n148 0.474125
R20974 Folded_Diff_Op_Amp_Layout_0.OUT2.n125 Folded_Diff_Op_Amp_Layout_0.OUT2.n149 0.474125
R20975 Folded_Diff_Op_Amp_Layout_0.OUT2.n33 Folded_Diff_Op_Amp_Layout_0.OUT2.n32 0.279824
R20976 Folded_Diff_Op_Amp_Layout_0.OUT2.n62 Folded_Diff_Op_Amp_Layout_0.OUT2.n61 0.279823
R20977 Folded_Diff_Op_Amp_Layout_0.OUT2.n54 Folded_Diff_Op_Amp_Layout_0.OUT2.n53 0.279823
R20978 Folded_Diff_Op_Amp_Layout_0.OUT2.n40 Folded_Diff_Op_Amp_Layout_0.OUT2.n39 0.279823
R20979 Folded_Diff_Op_Amp_Layout_0.OUT2.n80 Folded_Diff_Op_Amp_Layout_0.OUT2.n79 0.279615
R20980 Folded_Diff_Op_Amp_Layout_0.OUT2.n72 Folded_Diff_Op_Amp_Layout_0.OUT2.n71 0.279615
R20981 Folded_Diff_Op_Amp_Layout_0.OUT2.n112 Folded_Diff_Op_Amp_Layout_0.OUT2.n111 0.239196
R20982 Folded_Diff_Op_Amp_Layout_0.OUT2.n194 Folded_Diff_Op_Amp_Layout_0.OUT2.n193 0.238721
R20983 Folded_Diff_Op_Amp_Layout_0.OUT2.n105 Folded_Diff_Op_Amp_Layout_0.OUT2.n95 0.207891
R20984 Folded_Diff_Op_Amp_Layout_0.OUT2.n200 Folded_Diff_Op_Amp_Layout_0.OUT2.n202 0.19908
R20985 Folded_Diff_Op_Amp_Layout_0.OUT2.n107 Folded_Diff_Op_Amp_Layout_0.OUT2.n106 0.190283
R20986 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.OUT2.n199 0.0999375
R20987 Folded_Diff_Op_Amp_Layout_0.OUT2.n200 Folded_Diff_Op_Amp_Layout_0.OUT2.n203 0.0935118
R20988 Folded_Diff_Op_Amp_Layout_0.OUT2.n16 Folded_Diff_Op_Amp_Layout_0.OUT2.n10 0.106801
R20989 Folded_Diff_Op_Amp_Layout_0.OUT2.n136 Folded_Diff_Op_Amp_Layout_0.OUT2.n130 0.0823987
R20990 Folded_Diff_Op_Amp_Layout_0.OUT2.n185 Folded_Diff_Op_Amp_Layout_0.OUT2.n180 0.0823987
R20991 Folded_Diff_Op_Amp_Layout_0.OUT2.n14 Folded_Diff_Op_Amp_Layout_0.OUT2.n11 0.0790912
R20992 Folded_Diff_Op_Amp_Layout_0.OUT2.n3 Folded_Diff_Op_Amp_Layout_0.OUT2.n0 0.0786471
R20993 Folded_Diff_Op_Amp_Layout_0.OUT2.n114 Folded_Diff_Op_Amp_Layout_0.OUT2.n108 0.0712285
R20994 Folded_Diff_Op_Amp_Layout_0.OUT2.n177 Folded_Diff_Op_Amp_Layout_0.OUT2.n172 0.0712285
R20995 Folded_Diff_Op_Amp_Layout_0.OUT2.n124 Folded_Diff_Op_Amp_Layout_0.OUT2.n120 0.0712285
R20996 Folded_Diff_Op_Amp_Layout_0.OUT2.n147 Folded_Diff_Op_Amp_Layout_0.OUT2.n142 0.0712285
R20997 Folded_Diff_Op_Amp_Layout_0.OUT2.n24 Folded_Diff_Op_Amp_Layout_0.OUT2.n23 0.0603944
R20998 Folded_Diff_Op_Amp_Layout_0.OUT2.n112 Folded_Diff_Op_Amp_Layout_0.OUT2.n110 0.0568678
R20999 Folded_Diff_Op_Amp_Layout_0.OUT2.n114 Folded_Diff_Op_Amp_Layout_0.OUT2.n113 0.0534597
R21000 Folded_Diff_Op_Amp_Layout_0.OUT2.n177 Folded_Diff_Op_Amp_Layout_0.OUT2.n176 0.0534597
R21001 Folded_Diff_Op_Amp_Layout_0.OUT2.n147 Folded_Diff_Op_Amp_Layout_0.OUT2.n146 0.0534597
R21002 Folded_Diff_Op_Amp_Layout_0.OUT2.n124 Folded_Diff_Op_Amp_Layout_0.OUT2.n123 0.0534597
R21003 Folded_Diff_Op_Amp_Layout_0.OUT2.n134 Folded_Diff_Op_Amp_Layout_0.OUT2.n133 0.0419474
R21004 Folded_Diff_Op_Amp_Layout_0.OUT2.n185 Folded_Diff_Op_Amp_Layout_0.OUT2.n184 0.0415773
R21005 Folded_Diff_Op_Amp_Layout_0.OUT2.n136 Folded_Diff_Op_Amp_Layout_0.OUT2.n135 0.0415773
R21006 Folded_Diff_Op_Amp_Layout_0.OUT2.n189 Folded_Diff_Op_Amp_Layout_0.OUT2.n171 0.0354016
R21007 Folded_Diff_Op_Amp_Layout_0.OUT2.n192 Folded_Diff_Op_Amp_Layout_0.OUT2.n191 0.0354016
R21008 Folded_Diff_Op_Amp_Layout_0.OUT2.n16 Folded_Diff_Op_Amp_Layout_0.OUT2.n15 0.0319869
R21009 Folded_Diff_Op_Amp_Layout_0.OUT2.n26 Folded_Diff_Op_Amp_Layout_0.OUT2.n19 0.0296151
R21010 Folded_Diff_Op_Amp_Layout_0.OUT2.n203 Folded_Diff_Op_Amp_Layout_0.OUT2.n201 0.0230949
R21011 Folded_Diff_Op_Amp_Layout_0.OUT2.n18 Folded_Diff_Op_Amp_Layout_0.OUT2.n197 0.0229474
R21012 Folded_Diff_Op_Amp_Layout_0.OUT2.n160 Folded_Diff_Op_Amp_Layout_0.OUT2.n159 0.0228651
R21013 Folded_Diff_Op_Amp_Layout_0.OUT2.n141 Folded_Diff_Op_Amp_Layout_0.OUT2.n140 0.0201463
R21014 Folded_Diff_Op_Amp_Layout_0.OUT2.n119 Folded_Diff_Op_Amp_Layout_0.OUT2.n118 0.0201463
R21015 Folded_Diff_Op_Amp_Layout_0.OUT2.n157 Folded_Diff_Op_Amp_Layout_0.OUT2.n156 0.0182008
R21016 Folded_Diff_Op_Amp_Layout_0.OUT2.n190 Folded_Diff_Op_Amp_Layout_0.OUT2.n189 0.0182008
R21017 Folded_Diff_Op_Amp_Layout_0.OUT2.n193 Folded_Diff_Op_Amp_Layout_0.OUT2.n192 0.0182008
R21018 Folded_Diff_Op_Amp_Layout_0.OUT2.n165 Folded_Diff_Op_Amp_Layout_0.OUT2.n164 0.0179841
R21019 Folded_Diff_Op_Amp_Layout_0.OUT2.n167 Folded_Diff_Op_Amp_Layout_0.OUT2.n165 0.0177304
R21020 Folded_Diff_Op_Amp_Layout_0.OUT2.n162 Folded_Diff_Op_Amp_Layout_0.OUT2.n161 0.0173591
R21021 Folded_Diff_Op_Amp_Layout_0.OUT2.n164 Folded_Diff_Op_Amp_Layout_0.OUT2.n163 0.0173591
R21022 Folded_Diff_Op_Amp_Layout_0.OUT2.n163 Folded_Diff_Op_Amp_Layout_0.OUT2.n162 0.0173591
R21023 Folded_Diff_Op_Amp_Layout_0.OUT2.n161 Folded_Diff_Op_Amp_Layout_0.OUT2.n160 0.0173591
R21024 Folded_Diff_Op_Amp_Layout_0.OUT2.n19 Folded_Diff_Op_Amp_Layout_0.OUT2.t0 3.89253
R21025 Folded_Diff_Op_Amp_Layout_0.OUT2.n26 Folded_Diff_Op_Amp_Layout_0.OUT2.n25 0.0289893
R21026 Folded_Diff_Op_Amp_Layout_0.OUT2.n117 Folded_Diff_Op_Amp_Layout_0.OUT2.n116 0.016662
R21027 Folded_Diff_Op_Amp_Layout_0.OUT2.n149 Folded_Diff_Op_Amp_Layout_0.OUT2.n138 0.016662
R21028 Folded_Diff_Op_Amp_Layout_0.OUT2.n126 Folded_Diff_Op_Amp_Layout_0.OUT2.n125 0.016662
R21029 Folded_Diff_Op_Amp_Layout_0.OUT2.n179 Folded_Diff_Op_Amp_Layout_0.OUT2.n178 0.016662
R21030 Folded_Diff_Op_Amp_Layout_0.OUT2.n138 Folded_Diff_Op_Amp_Layout_0.OUT2.n137 0.0166619
R21031 Folded_Diff_Op_Amp_Layout_0.OUT2.n170 Folded_Diff_Op_Amp_Layout_0.OUT2.n169 0.0163451
R21032 Folded_Diff_Op_Amp_Layout_0.OUT2.n116 Folded_Diff_Op_Amp_Layout_0.OUT2.n115 0.0156875
R21033 Folded_Diff_Op_Amp_Layout_0.OUT2.n7 Folded_Diff_Op_Amp_Layout_0.OUT2.n6 0.0156875
R21034 Folded_Diff_Op_Amp_Layout_0.OUT2.n155 Folded_Diff_Op_Amp_Layout_0.OUT2.n154 0.0156875
R21035 Folded_Diff_Op_Amp_Layout_0.OUT2.n187 Folded_Diff_Op_Amp_Layout_0.OUT2.n179 0.0156875
R21036 Folded_Diff_Op_Amp_Layout_0.OUT2.n150 Folded_Diff_Op_Amp_Layout_0.OUT2.n126 0.0156875
R21037 Folded_Diff_Op_Amp_Layout_0.OUT2.n196 Folded_Diff_Op_Amp_Layout_0.OUT2.n5 0.014
R21038 Folded_Diff_Op_Amp_Layout_0.OUT2.n5 Folded_Diff_Op_Amp_Layout_0.OUT2.n195 0.014
R21039 Folded_Diff_Op_Amp_Layout_0.OUT2.n197 Folded_Diff_Op_Amp_Layout_0.OUT2.n196 0.0134654
R21040 Folded_Diff_Op_Amp_Layout_0.OUT2.n159 Folded_Diff_Op_Amp_Layout_0.OUT2.n158 0.0119325
R21041 Folded_Diff_Op_Amp_Layout_0.OUT2.n25 Folded_Diff_Op_Amp_Layout_0.OUT2.n24 0.0200461
R21042 Folded_Diff_Op_Amp_Layout_0.OUT2.n199 Folded_Diff_Op_Amp_Layout_0.OUT2.n18 0.0199708
R21043 Folded_Diff_Op_Amp_Layout_0.OUT2.n17 Folded_Diff_Op_Amp_Layout_0.OUT2.n9 0.014159
R21044 Folded_Diff_Op_Amp_Layout_0.OUT2.n169 Folded_Diff_Op_Amp_Layout_0.OUT2.n168 0.0112521
R21045 Folded_Diff_Op_Amp_Layout_0.OUT2.n17 Folded_Diff_Op_Amp_Layout_0.OUT2.n8 0.0111023
R21046 Folded_Diff_Op_Amp_Layout_0.OUT2.n21 Folded_Diff_Op_Amp_Layout_0.OUT2.n20 0.010845
R21047 Folded_Diff_Op_Amp_Layout_0.VPD.n70 Folded_Diff_Op_Amp_Layout_0.VPD.t20 5.22731
R21048 Folded_Diff_Op_Amp_Layout_0.VPD.n64 Folded_Diff_Op_Amp_Layout_0.VPD.n63 5.20893
R21049 Folded_Diff_Op_Amp_Layout_0.VPD.n61 Folded_Diff_Op_Amp_Layout_0.VPD.t23 5.20893
R21050 Folded_Diff_Op_Amp_Layout_0.VPD.n60 Folded_Diff_Op_Amp_Layout_0.VPD.n59 5.20893
R21051 Folded_Diff_Op_Amp_Layout_0.VPD.n30 Folded_Diff_Op_Amp_Layout_0.VPD.n29 5.11385
R21052 Folded_Diff_Op_Amp_Layout_0.VPD.n47 Folded_Diff_Op_Amp_Layout_0.VPD.t7 5.11385
R21053 Folded_Diff_Op_Amp_Layout_0.VPD.n55 Folded_Diff_Op_Amp_Layout_0.VPD.t22 4.55153
R21054 Folded_Diff_Op_Amp_Layout_0.VPD.n95 Folded_Diff_Op_Amp_Layout_0.VPD.t27 4.55153
R21055 Folded_Diff_Op_Amp_Layout_0.VPD.n36 Folded_Diff_Op_Amp_Layout_0.VPD.n35 4.53238
R21056 Folded_Diff_Op_Amp_Layout_0.VPD.n57 Folded_Diff_Op_Amp_Layout_0.VPD.n53 3.92545
R21057 Folded_Diff_Op_Amp_Layout_0.VPD.n56 Folded_Diff_Op_Amp_Layout_0.VPD.t17 3.92545
R21058 Folded_Diff_Op_Amp_Layout_0.VPD.n55 Folded_Diff_Op_Amp_Layout_0.VPD.n54 3.92545
R21059 Folded_Diff_Op_Amp_Layout_0.VPD.n96 Folded_Diff_Op_Amp_Layout_0.VPD.t30 3.92545
R21060 Folded_Diff_Op_Amp_Layout_0.VPD.n95 Folded_Diff_Op_Amp_Layout_0.VPD.n94 3.92545
R21061 Folded_Diff_Op_Amp_Layout_0.VPD.n64 Folded_Diff_Op_Amp_Layout_0.VPD.n62 3.18197
R21062 Folded_Diff_Op_Amp_Layout_0.VPD.n61 Folded_Diff_Op_Amp_Layout_0.VPD.t21 3.18197
R21063 Folded_Diff_Op_Amp_Layout_0.VPD.n60 Folded_Diff_Op_Amp_Layout_0.VPD.n58 3.18197
R21064 Folded_Diff_Op_Amp_Layout_0.VPD.n127 Folded_Diff_Op_Amp_Layout_0.VPD.n126 2.26288
R21065 Folded_Diff_Op_Amp_Layout_0.VPD.n65 Folded_Diff_Op_Amp_Layout_0.VPD.n64 1.87093
R21066 Folded_Diff_Op_Amp_Layout_0.VPD.n70 Folded_Diff_Op_Amp_Layout_0.VPD.n69 1.55818
R21067 Folded_Diff_Op_Amp_Layout_0.VPD.n24 Folded_Diff_Op_Amp_Layout_0.VPD.n23 1.49812
R21068 Folded_Diff_Op_Amp_Layout_0.VPD.n138 Folded_Diff_Op_Amp_Layout_0.VPD.n137 1.49801
R21069 Folded_Diff_Op_Amp_Layout_0.VPD.n97 Folded_Diff_Op_Amp_Layout_0.VPD.n96 1.276
R21070 Folded_Diff_Op_Amp_Layout_0.VPD.n5 Folded_Diff_Op_Amp_Layout_0.VPD.n4 1.19453
R21071 Folded_Diff_Op_Amp_Layout_0.VPD.n16 Folded_Diff_Op_Amp_Layout_0.VPD.n15 1.19453
R21072 Folded_Diff_Op_Amp_Layout_0.VPD.n27 Folded_Diff_Op_Amp_Layout_0.VPD.n26 1.18339
R21073 Folded_Diff_Op_Amp_Layout_0.VPD.n45 Folded_Diff_Op_Amp_Layout_0.VPD.n44 1.18339
R21074 Folded_Diff_Op_Amp_Layout_0.VPD.n41 Folded_Diff_Op_Amp_Layout_0.VPD.n40 1.18329
R21075 Folded_Diff_Op_Amp_Layout_0.VPD.n92 Folded_Diff_Op_Amp_Layout_0.VPD.n91 1.18328
R21076 Folded_Diff_Op_Amp_Layout_0.VPD.n110 Folded_Diff_Op_Amp_Layout_0.VPD.n109 1.17867
R21077 Folded_Diff_Op_Amp_Layout_0.VPD.n121 Folded_Diff_Op_Amp_Layout_0.VPD.n120 1.17867
R21078 Folded_Diff_Op_Amp_Layout_0.VPD.n42 Folded_Diff_Op_Amp_Layout_0.VPD.n41 1.17343
R21079 Folded_Diff_Op_Amp_Layout_0.VPD.n28 Folded_Diff_Op_Amp_Layout_0.VPD.n27 1.17279
R21080 Folded_Diff_Op_Amp_Layout_0.VPD.n46 Folded_Diff_Op_Amp_Layout_0.VPD.n45 1.17279
R21081 Folded_Diff_Op_Amp_Layout_0.VPD.n93 Folded_Diff_Op_Amp_Layout_0.VPD.n92 1.17279
R21082 Folded_Diff_Op_Amp_Layout_0.VPD.n56 Folded_Diff_Op_Amp_Layout_0.VPD.n55 1.12746
R21083 Folded_Diff_Op_Amp_Layout_0.VPD.n96 Folded_Diff_Op_Amp_Layout_0.VPD.n95 1.12746
R21084 Folded_Diff_Op_Amp_Layout_0.VPD.n75 Folded_Diff_Op_Amp_Layout_0.VPD.n74 1.13842
R21085 Folded_Diff_Op_Amp_Layout_0.VPD.n32 Folded_Diff_Op_Amp_Layout_0.VPD.n31 1.1255
R21086 Folded_Diff_Op_Amp_Layout_0.VPD.n49 Folded_Diff_Op_Amp_Layout_0.VPD.n48 1.1255
R21087 Folded_Diff_Op_Amp_Layout_0.VPD.n74 Folded_Diff_Op_Amp_Layout_0.VPD.n73 1.1255
R21088 Folded_Diff_Op_Amp_Layout_0.VPD.n139 Folded_Diff_Op_Amp_Layout_0.VPD.n138 1.1255
R21089 Folded_Diff_Op_Amp_Layout_0.VPD.n99 Folded_Diff_Op_Amp_Layout_0.VPD.n98 1.1255
R21090 Folded_Diff_Op_Amp_Layout_0.VPD.n38 Folded_Diff_Op_Amp_Layout_0.VPD.n37 1.1255
R21091 Folded_Diff_Op_Amp_Layout_0.VPD.n127 Folded_Diff_Op_Amp_Layout_0.VPD.n89 0.926774
R21092 Folded_Diff_Op_Amp_Layout_0.VPD.n67 Folded_Diff_Op_Amp_Layout_0.VPD.n66 0.877022
R21093 Folded_Diff_Op_Amp_Layout_0.VPD.n105 Folded_Diff_Op_Amp_Layout_0.VPD.n104 0.87575
R21094 Folded_Diff_Op_Amp_Layout_0.VPD.n109 Folded_Diff_Op_Amp_Layout_0.VPD.n108 0.824494
R21095 Folded_Diff_Op_Amp_Layout_0.VPD.n120 Folded_Diff_Op_Amp_Layout_0.VPD.n119 0.824494
R21096 Folded_Diff_Op_Amp_Layout_0.VPD.n4 Folded_Diff_Op_Amp_Layout_0.VPD.n3 0.824332
R21097 Folded_Diff_Op_Amp_Layout_0.VPD.n15 Folded_Diff_Op_Amp_Layout_0.VPD.n14 0.824332
R21098 Folded_Diff_Op_Amp_Layout_0.VPD.n65 Folded_Diff_Op_Amp_Layout_0.VPD.n61 0.743978
R21099 Folded_Diff_Op_Amp_Layout_0.VPD.n66 Folded_Diff_Op_Amp_Layout_0.VPD.n60 0.743978
R21100 Folded_Diff_Op_Amp_Layout_0.VPD.n19 Folded_Diff_Op_Amp_Layout_0.VPD.n18 0.727916
R21101 Folded_Diff_Op_Amp_Layout_0.VPD.n113 Folded_Diff_Op_Amp_Layout_0.VPD.n112 0.727916
R21102 Folded_Diff_Op_Amp_Layout_0.VPD.n124 Folded_Diff_Op_Amp_Layout_0.VPD.n123 0.727916
R21103 Folded_Diff_Op_Amp_Layout_0.VPD.n83 Folded_Diff_Op_Amp_Layout_0.VPD.n43 0.727104
R21104 Folded_Diff_Op_Amp_Layout_0.VPD.n57 Folded_Diff_Op_Amp_Layout_0.VPD.n56 0.626587
R21105 Folded_Diff_Op_Amp_Layout_0.VPD.n66 Folded_Diff_Op_Amp_Layout_0.VPD.n65 0.626587
R21106 Folded_Diff_Op_Amp_Layout_0.VPD.n77 Folded_Diff_Op_Amp_Layout_0.VPD.n76 0.62375
R21107 Folded_Diff_Op_Amp_Layout_0.VPD.n87 Folded_Diff_Op_Amp_Layout_0.VPD.n33 0.616779
R21108 Folded_Diff_Op_Amp_Layout_0.VPD.n78 Folded_Diff_Op_Amp_Layout_0.VPD.n50 0.616779
R21109 Folded_Diff_Op_Amp_Layout_0.VPD.n8 Folded_Diff_Op_Amp_Layout_0.VPD.n6 0.616779
R21110 Folded_Diff_Op_Amp_Layout_0.VPD.n102 Folded_Diff_Op_Amp_Layout_0.VPD.n100 0.616779
R21111 Folded_Diff_Op_Amp_Layout_0.VPD.n26 Folded_Diff_Op_Amp_Layout_0.VPD.n25 0.58197
R21112 Folded_Diff_Op_Amp_Layout_0.VPD.n44 Folded_Diff_Op_Amp_Layout_0.VPD.t5 0.58197
R21113 Folded_Diff_Op_Amp_Layout_0.VPD.n69 Folded_Diff_Op_Amp_Layout_0.VPD.t19 0.58197
R21114 Folded_Diff_Op_Amp_Layout_0.VPD.n3 Folded_Diff_Op_Amp_Layout_0.VPD.t12 0.58197
R21115 Folded_Diff_Op_Amp_Layout_0.VPD.n3 Folded_Diff_Op_Amp_Layout_0.VPD.n2 0.58197
R21116 Folded_Diff_Op_Amp_Layout_0.VPD.n14 Folded_Diff_Op_Amp_Layout_0.VPD.t8 0.58197
R21117 Folded_Diff_Op_Amp_Layout_0.VPD.n14 Folded_Diff_Op_Amp_Layout_0.VPD.n13 0.58197
R21118 Folded_Diff_Op_Amp_Layout_0.VPD.n91 Folded_Diff_Op_Amp_Layout_0.VPD.n90 0.58197
R21119 Folded_Diff_Op_Amp_Layout_0.VPD.n108 Folded_Diff_Op_Amp_Layout_0.VPD.t11 0.58197
R21120 Folded_Diff_Op_Amp_Layout_0.VPD.n108 Folded_Diff_Op_Amp_Layout_0.VPD.n107 0.58197
R21121 Folded_Diff_Op_Amp_Layout_0.VPD.n119 Folded_Diff_Op_Amp_Layout_0.VPD.t3 0.58197
R21122 Folded_Diff_Op_Amp_Layout_0.VPD.n119 Folded_Diff_Op_Amp_Layout_0.VPD.n118 0.58197
R21123 Folded_Diff_Op_Amp_Layout_0.VPD.n35 Folded_Diff_Op_Amp_Layout_0.VPD.t1 0.58197
R21124 Folded_Diff_Op_Amp_Layout_0.VPD.n35 Folded_Diff_Op_Amp_Layout_0.VPD.n34 0.58197
R21125 Folded_Diff_Op_Amp_Layout_0.VPD.n40 Folded_Diff_Op_Amp_Layout_0.VPD.t15 0.58197
R21126 Folded_Diff_Op_Amp_Layout_0.VPD.n40 Folded_Diff_Op_Amp_Layout_0.VPD.n39 0.58197
R21127 Folded_Diff_Op_Amp_Layout_0.VPD.n22 Folded_Diff_Op_Amp_Layout_0.VPD.n21 0.53025
R21128 Folded_Diff_Op_Amp_Layout_0.VPD.n68 Folded_Diff_Op_Amp_Layout_0.VPD.n67 0.442674
R21129 Folded_Diff_Op_Amp_Layout_0.VPD.n67 Folded_Diff_Op_Amp_Layout_0.VPD.n57 0.3605
R21130 Folded_Diff_Op_Amp_Layout_0.VPD.n98 Folded_Diff_Op_Amp_Layout_0.VPD.n97 0.330999
R21131 Folded_Diff_Op_Amp_Layout_0.VPD.n11 Folded_Diff_Op_Amp_Layout_0.VPD.n10 0.330125
R21132 Folded_Diff_Op_Amp_Layout_0.VPD.n116 Folded_Diff_Op_Amp_Layout_0.VPD.n115 0.330125
R21133 Folded_Diff_Op_Amp_Layout_0.VPD.n86 Folded_Diff_Op_Amp_Layout_0.VPD.n85 0.330125
R21134 Folded_Diff_Op_Amp_Layout_0.VPD.n81 Folded_Diff_Op_Amp_Layout_0.VPD.n80 0.330125
R21135 Folded_Diff_Op_Amp_Layout_0.VPD.n31 Folded_Diff_Op_Amp_Layout_0.VPD.n30 0.32803
R21136 Folded_Diff_Op_Amp_Layout_0.VPD.n48 Folded_Diff_Op_Amp_Layout_0.VPD.n47 0.32803
R21137 Folded_Diff_Op_Amp_Layout_0.VPD.n37 Folded_Diff_Op_Amp_Layout_0.VPD.n36 0.32803
R21138 Folded_Diff_Op_Amp_Layout_0.VPD.n128 Folded_Diff_Op_Amp_Layout_0.VPD.n127 0.323011
R21139 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VPD.n139 0.29625
R21140 Folded_Diff_Op_Amp_Layout_0.VPD.n71 Folded_Diff_Op_Amp_Layout_0.VPD.n70 0.201042
R21141 Folded_Diff_Op_Amp_Layout_0.VPD.n72 Folded_Diff_Op_Amp_Layout_0.VPD.n71 0.0953821
R21142 Folded_Diff_Op_Amp_Layout_0.VPD.n74 Folded_Diff_Op_Amp_Layout_0.VPD.n52 0.0832399
R21143 Folded_Diff_Op_Amp_Layout_0.VPD.n18 Folded_Diff_Op_Amp_Layout_0.VPD.n17 0.0826464
R21144 Folded_Diff_Op_Amp_Layout_0.VPD.n112 Folded_Diff_Op_Amp_Layout_0.VPD.n111 0.0826464
R21145 Folded_Diff_Op_Amp_Layout_0.VPD.n123 Folded_Diff_Op_Amp_Layout_0.VPD.n122 0.0826464
R21146 Folded_Diff_Op_Amp_Layout_0.VPD.n43 Folded_Diff_Op_Amp_Layout_0.VPD.n38 0.0823987
R21147 Folded_Diff_Op_Amp_Layout_0.VPD.n6 Folded_Diff_Op_Amp_Layout_0.VPD.n1 0.0712285
R21148 Folded_Diff_Op_Amp_Layout_0.VPD.n100 Folded_Diff_Op_Amp_Layout_0.VPD.n93 0.0712285
R21149 Folded_Diff_Op_Amp_Layout_0.VPD.n50 Folded_Diff_Op_Amp_Layout_0.VPD.n46 0.0712285
R21150 Folded_Diff_Op_Amp_Layout_0.VPD.n33 Folded_Diff_Op_Amp_Layout_0.VPD.n28 0.0712285
R21151 Folded_Diff_Op_Amp_Layout_0.VPD.n73 Folded_Diff_Op_Amp_Layout_0.VPD.n68 0.0552826
R21152 Folded_Diff_Op_Amp_Layout_0.VPD.n6 Folded_Diff_Op_Amp_Layout_0.VPD.n5 0.0534597
R21153 Folded_Diff_Op_Amp_Layout_0.VPD.n100 Folded_Diff_Op_Amp_Layout_0.VPD.n99 0.0534597
R21154 Folded_Diff_Op_Amp_Layout_0.VPD.n33 Folded_Diff_Op_Amp_Layout_0.VPD.n32 0.0534597
R21155 Folded_Diff_Op_Amp_Layout_0.VPD.n50 Folded_Diff_Op_Amp_Layout_0.VPD.n49 0.0534597
R21156 Folded_Diff_Op_Amp_Layout_0.VPD.n18 Folded_Diff_Op_Amp_Layout_0.VPD.n16 0.0423164
R21157 Folded_Diff_Op_Amp_Layout_0.VPD.n112 Folded_Diff_Op_Amp_Layout_0.VPD.n110 0.0423164
R21158 Folded_Diff_Op_Amp_Layout_0.VPD.n123 Folded_Diff_Op_Amp_Layout_0.VPD.n121 0.0423164
R21159 Folded_Diff_Op_Amp_Layout_0.VPD.n52 Folded_Diff_Op_Amp_Layout_0.VPD.n51 0.0419676
R21160 Folded_Diff_Op_Amp_Layout_0.VPD.n43 Folded_Diff_Op_Amp_Layout_0.VPD.n42 0.0415773
R21161 Folded_Diff_Op_Amp_Layout_0.VPD.n73 Folded_Diff_Op_Amp_Layout_0.VPD.n72 0.0293873
R21162 Folded_Diff_Op_Amp_Layout_0.VPD.n135 Folded_Diff_Op_Amp_Layout_0.VPD.n134 0.0229474
R21163 Folded_Diff_Op_Amp_Layout_0.VPD.n8 Folded_Diff_Op_Amp_Layout_0.VPD.n7 0.0156875
R21164 Folded_Diff_Op_Amp_Layout_0.VPD.n102 Folded_Diff_Op_Amp_Layout_0.VPD.n101 0.0156875
R21165 Folded_Diff_Op_Amp_Layout_0.VPD.n87 Folded_Diff_Op_Amp_Layout_0.VPD.n86 0.0156875
R21166 Folded_Diff_Op_Amp_Layout_0.VPD.n78 Folded_Diff_Op_Amp_Layout_0.VPD.n77 0.0156875
R21167 Folded_Diff_Op_Amp_Layout_0.VPD.n23 Folded_Diff_Op_Amp_Layout_0.VPD.n22 0.014
R21168 Folded_Diff_Op_Amp_Layout_0.VPD.n138 Folded_Diff_Op_Amp_Layout_0.VPD.n133 0.014
R21169 Folded_Diff_Op_Amp_Layout_0.VPD.n131 Folded_Diff_Op_Amp_Layout_0.VPD.n130 0.014
R21170 Folded_Diff_Op_Amp_Layout_0.VPD.n133 Folded_Diff_Op_Amp_Layout_0.VPD.n132 0.0134654
R21171 Folded_Diff_Op_Amp_Layout_0.VPD.n132 Folded_Diff_Op_Amp_Layout_0.VPD.n131 0.0134654
R21172 Folded_Diff_Op_Amp_Layout_0.VPD.n88 Folded_Diff_Op_Amp_Layout_0.VPD.n87 0.00860784
R21173 Folded_Diff_Op_Amp_Layout_0.VPD.n83 Folded_Diff_Op_Amp_Layout_0.VPD.n82 0.00860784
R21174 Folded_Diff_Op_Amp_Layout_0.VPD.n79 Folded_Diff_Op_Amp_Layout_0.VPD.n78 0.00860784
R21175 Folded_Diff_Op_Amp_Layout_0.VPD.n9 Folded_Diff_Op_Amp_Layout_0.VPD.n8 0.00860784
R21176 Folded_Diff_Op_Amp_Layout_0.VPD.n103 Folded_Diff_Op_Amp_Layout_0.VPD.n102 0.00860784
R21177 Folded_Diff_Op_Amp_Layout_0.VPD.n20 Folded_Diff_Op_Amp_Layout_0.VPD.n19 0.00858096
R21178 Folded_Diff_Op_Amp_Layout_0.VPD.n12 Folded_Diff_Op_Amp_Layout_0.VPD.n11 0.00858096
R21179 Folded_Diff_Op_Amp_Layout_0.VPD.n21 Folded_Diff_Op_Amp_Layout_0.VPD.n20 0.00858096
R21180 Folded_Diff_Op_Amp_Layout_0.VPD.n19 Folded_Diff_Op_Amp_Layout_0.VPD.n12 0.00858096
R21181 Folded_Diff_Op_Amp_Layout_0.VPD.n125 Folded_Diff_Op_Amp_Layout_0.VPD.n124 0.00858096
R21182 Folded_Diff_Op_Amp_Layout_0.VPD.n117 Folded_Diff_Op_Amp_Layout_0.VPD.n116 0.00858096
R21183 Folded_Diff_Op_Amp_Layout_0.VPD.n114 Folded_Diff_Op_Amp_Layout_0.VPD.n113 0.00858096
R21184 Folded_Diff_Op_Amp_Layout_0.VPD.n106 Folded_Diff_Op_Amp_Layout_0.VPD.n105 0.00858096
R21185 Folded_Diff_Op_Amp_Layout_0.VPD.n126 Folded_Diff_Op_Amp_Layout_0.VPD.n125 0.00858096
R21186 Folded_Diff_Op_Amp_Layout_0.VPD.n124 Folded_Diff_Op_Amp_Layout_0.VPD.n117 0.00858096
R21187 Folded_Diff_Op_Amp_Layout_0.VPD.n115 Folded_Diff_Op_Amp_Layout_0.VPD.n114 0.00858096
R21188 Folded_Diff_Op_Amp_Layout_0.VPD.n113 Folded_Diff_Op_Amp_Layout_0.VPD.n106 0.00858096
R21189 Folded_Diff_Op_Amp_Layout_0.VPD.n85 Folded_Diff_Op_Amp_Layout_0.VPD.n84 0.00858096
R21190 Folded_Diff_Op_Amp_Layout_0.VPD.n84 Folded_Diff_Op_Amp_Layout_0.VPD.n83 0.00858096
R21191 Folded_Diff_Op_Amp_Layout_0.VPD.n10 Folded_Diff_Op_Amp_Layout_0.VPD.n9 0.00855417
R21192 Folded_Diff_Op_Amp_Layout_0.VPD.n104 Folded_Diff_Op_Amp_Layout_0.VPD.n103 0.00855417
R21193 Folded_Diff_Op_Amp_Layout_0.VPD.n89 Folded_Diff_Op_Amp_Layout_0.VPD.n88 0.00855417
R21194 Folded_Diff_Op_Amp_Layout_0.VPD.n82 Folded_Diff_Op_Amp_Layout_0.VPD.n81 0.00855417
R21195 Folded_Diff_Op_Amp_Layout_0.VPD.n80 Folded_Diff_Op_Amp_Layout_0.VPD.n79 0.00855417
R21196 Folded_Diff_Op_Amp_Layout_0.VPD.n76 Folded_Diff_Op_Amp_Layout_0.VPD.n75 0.00855417
R21197 Folded_Diff_Op_Amp_Layout_0.VPD.n23 Folded_Diff_Op_Amp_Layout_0.VPD.n0 0.00773989
R21198 Folded_Diff_Op_Amp_Layout_0.VPD.n129 Folded_Diff_Op_Amp_Layout_0.VPD.n128 0.00773989
R21199 Folded_Diff_Op_Amp_Layout_0.VPD.n130 Folded_Diff_Op_Amp_Layout_0.VPD.n129 0.00773989
R21200 Folded_Diff_Op_Amp_Layout_0.VPD.n138 Folded_Diff_Op_Amp_Layout_0.VPD.n24 0.00582347
R21201 Folded_Diff_Op_Amp_Layout_0.VPD.n137 Folded_Diff_Op_Amp_Layout_0.VPD.n136 0.00549102
R21202 Folded_Diff_Op_Amp_Layout_0.VPD.n136 Folded_Diff_Op_Amp_Layout_0.VPD.n135 0.00549102
R21203 Folded_Diff_Op_Amp_Layout_0.VND.n11 Folded_Diff_Op_Amp_Layout_0.VND.t24 5.20893
R21204 Folded_Diff_Op_Amp_Layout_0.VND.n14 Folded_Diff_Op_Amp_Layout_0.VND.n12 5.20893
R21205 Folded_Diff_Op_Amp_Layout_0.VND.n15 Folded_Diff_Op_Amp_Layout_0.VND.t21 5.20893
R21206 Folded_Diff_Op_Amp_Layout_0.VND.n2 Folded_Diff_Op_Amp_Layout_0.VND.n1 5.11992
R21207 Folded_Diff_Op_Amp_Layout_0.VND.n8 Folded_Diff_Op_Amp_Layout_0.VND.n7 5.0524
R21208 Folded_Diff_Op_Amp_Layout_0.VND.n102 Folded_Diff_Op_Amp_Layout_0.VND.n101 5.0524
R21209 Folded_Diff_Op_Amp_Layout_0.VND.n37 Folded_Diff_Op_Amp_Layout_0.VND.n36 4.53845
R21210 Folded_Diff_Op_Amp_Layout_0.VND.n52 Folded_Diff_Op_Amp_Layout_0.VND.n51 4.53845
R21211 Folded_Diff_Op_Amp_Layout_0.VND.n10 Folded_Diff_Op_Amp_Layout_0.VND.t20 4.17588
R21212 Folded_Diff_Op_Amp_Layout_0.VND.n8 Folded_Diff_Op_Amp_Layout_0.VND.t25 3.92545
R21213 Folded_Diff_Op_Amp_Layout_0.VND.n9 Folded_Diff_Op_Amp_Layout_0.VND.n6 3.92545
R21214 Folded_Diff_Op_Amp_Layout_0.VND.n102 Folded_Diff_Op_Amp_Layout_0.VND.t19 3.92545
R21215 Folded_Diff_Op_Amp_Layout_0.VND.n103 Folded_Diff_Op_Amp_Layout_0.VND.n100 3.92545
R21216 Folded_Diff_Op_Amp_Layout_0.VND.n11 Folded_Diff_Op_Amp_Layout_0.VND.t29 3.18197
R21217 Folded_Diff_Op_Amp_Layout_0.VND.n14 Folded_Diff_Op_Amp_Layout_0.VND.n13 3.18197
R21218 Folded_Diff_Op_Amp_Layout_0.VND.n15 Folded_Diff_Op_Amp_Layout_0.VND.t27 3.18197
R21219 Folded_Diff_Op_Amp_Layout_0.VND.n21 Folded_Diff_Op_Amp_Layout_0.VND.n20 2.40175
R21220 Folded_Diff_Op_Amp_Layout_0.VND.n88 Folded_Diff_Op_Amp_Layout_0.VND.n87 1.65012
R21221 Folded_Diff_Op_Amp_Layout_0.VND.n139 Folded_Diff_Op_Amp_Layout_0.VND.n138 1.58409
R21222 Folded_Diff_Op_Amp_Layout_0.VND.n123 Folded_Diff_Op_Amp_Layout_0.VND.t3 1.58409
R21223 Folded_Diff_Op_Amp_Layout_0.VND.n107 Folded_Diff_Op_Amp_Layout_0.VND.t18 1.58402
R21224 Folded_Diff_Op_Amp_Layout_0.VND.n0 Folded_Diff_Op_Amp_Layout_0.VND.n146 1.50852
R21225 Folded_Diff_Op_Amp_Layout_0.VND.n114 Folded_Diff_Op_Amp_Layout_0.VND.n113 1.4964
R21226 Folded_Diff_Op_Amp_Layout_0.VND.n114 Folded_Diff_Op_Amp_Layout_0.VND.n109 1.48461
R21227 Folded_Diff_Op_Amp_Layout_0.VND.n60 Folded_Diff_Op_Amp_Layout_0.VND.t9 1.40773
R21228 Folded_Diff_Op_Amp_Layout_0.VND.n81 Folded_Diff_Op_Amp_Layout_0.VND.n80 1.40773
R21229 Folded_Diff_Op_Amp_Layout_0.VND.n16 Folded_Diff_Op_Amp_Layout_0.VND.n15 1.37007
R21230 Folded_Diff_Op_Amp_Layout_0.VND.n89 Folded_Diff_Op_Amp_Layout_0.VND.n88 1.35681
R21231 Folded_Diff_Op_Amp_Layout_0.VND.n104 Folded_Diff_Op_Amp_Layout_0.VND.n103 1.26302
R21232 Folded_Diff_Op_Amp_Layout_0.VND.n88 Folded_Diff_Op_Amp_Layout_0.VND.n58 1.25459
R21233 Folded_Diff_Op_Amp_Layout_0.VND.n61 Folded_Diff_Op_Amp_Layout_0.VND.n60 1.19469
R21234 Folded_Diff_Op_Amp_Layout_0.VND.n82 Folded_Diff_Op_Amp_Layout_0.VND.n81 1.19469
R21235 Folded_Diff_Op_Amp_Layout_0.VND.n72 Folded_Diff_Op_Amp_Layout_0.VND.n71 1.19441
R21236 Folded_Diff_Op_Amp_Layout_0.VND.n33 Folded_Diff_Op_Amp_Layout_0.VND.n32 1.18273
R21237 Folded_Diff_Op_Amp_Layout_0.VND.n48 Folded_Diff_Op_Amp_Layout_0.VND.n47 1.18273
R21238 Folded_Diff_Op_Amp_Layout_0.VND.n150 Folded_Diff_Op_Amp_Layout_0.VND.n90 1.1775
R21239 Folded_Diff_Op_Amp_Layout_0.VND.n34 Folded_Diff_Op_Amp_Layout_0.VND.n33 1.17276
R21240 Folded_Diff_Op_Amp_Layout_0.VND.n49 Folded_Diff_Op_Amp_Layout_0.VND.n48 1.17276
R21241 Folded_Diff_Op_Amp_Layout_0.VND.n140 Folded_Diff_Op_Amp_Layout_0.VND.n139 1.1643
R21242 Folded_Diff_Op_Amp_Layout_0.VND.n98 Folded_Diff_Op_Amp_Layout_0.VND.n97 1.1643
R21243 Folded_Diff_Op_Amp_Layout_0.VND.n124 Folded_Diff_Op_Amp_Layout_0.VND.n123 1.1643
R21244 Folded_Diff_Op_Amp_Layout_0.VND.n108 Folded_Diff_Op_Amp_Layout_0.VND.n107 1.1643
R21245 Folded_Diff_Op_Amp_Layout_0.VND.n17 Folded_Diff_Op_Amp_Layout_0.VND.n16 1.12746
R21246 Folded_Diff_Op_Amp_Layout_0.VND.n5 Folded_Diff_Op_Amp_Layout_0.VND.n4 1.1255
R21247 Folded_Diff_Op_Amp_Layout_0.VND.n23 Folded_Diff_Op_Amp_Layout_0.VND.n22 1.1255
R21248 Folded_Diff_Op_Amp_Layout_0.VND.n39 Folded_Diff_Op_Amp_Layout_0.VND.n38 1.1255
R21249 Folded_Diff_Op_Amp_Layout_0.VND.n150 Folded_Diff_Op_Amp_Layout_0.VND.n0 1.1255
R21250 Folded_Diff_Op_Amp_Layout_0.VND.n54 Folded_Diff_Op_Amp_Layout_0.VND.n53 1.1255
R21251 Folded_Diff_Op_Amp_Layout_0.VND.n126 Folded_Diff_Op_Amp_Layout_0.VND.n125 1.10737
R21252 Folded_Diff_Op_Amp_Layout_0.VND.n142 Folded_Diff_Op_Amp_Layout_0.VND.n141 1.10737
R21253 Folded_Diff_Op_Amp_Layout_0.VND.n97 Folded_Diff_Op_Amp_Layout_0.VND.n96 1.00262
R21254 Folded_Diff_Op_Amp_Layout_0.VND.n130 Folded_Diff_Op_Amp_Layout_0.VND.n99 0.88565
R21255 Folded_Diff_Op_Amp_Layout_0.VND.n10 Folded_Diff_Op_Amp_Layout_0.VND.n9 0.877022
R21256 Folded_Diff_Op_Amp_Layout_0.VND.n29 Folded_Diff_Op_Amp_Layout_0.VND.n28 0.87575
R21257 Folded_Diff_Op_Amp_Layout_0.VND.n71 Folded_Diff_Op_Amp_Layout_0.VND.n70 0.825944
R21258 Folded_Diff_Op_Amp_Layout_0.VND.n17 Folded_Diff_Op_Amp_Layout_0.VND.n11 0.743978
R21259 Folded_Diff_Op_Amp_Layout_0.VND.n16 Folded_Diff_Op_Amp_Layout_0.VND.n14 0.743978
R21260 Folded_Diff_Op_Amp_Layout_0.VND.n41 Folded_Diff_Op_Amp_Layout_0.VND.n40 0.727916
R21261 Folded_Diff_Op_Amp_Layout_0.VND.n56 Folded_Diff_Op_Amp_Layout_0.VND.n55 0.727916
R21262 Folded_Diff_Op_Amp_Layout_0.VND.n75 Folded_Diff_Op_Amp_Layout_0.VND.n74 0.727916
R21263 Folded_Diff_Op_Amp_Layout_0.VND.n85 Folded_Diff_Op_Amp_Layout_0.VND.n84 0.727916
R21264 Folded_Diff_Op_Amp_Layout_0.VND.n9 Folded_Diff_Op_Amp_Layout_0.VND.n8 0.626587
R21265 Folded_Diff_Op_Amp_Layout_0.VND.n18 Folded_Diff_Op_Amp_Layout_0.VND.n17 0.626587
R21266 Folded_Diff_Op_Amp_Layout_0.VND.n103 Folded_Diff_Op_Amp_Layout_0.VND.n102 0.626587
R21267 Folded_Diff_Op_Amp_Layout_0.VND.n117 Folded_Diff_Op_Amp_Layout_0.VND.n116 0.62375
R21268 Folded_Diff_Op_Amp_Layout_0.VND.n26 Folded_Diff_Op_Amp_Layout_0.VND.n24 0.616779
R21269 Folded_Diff_Op_Amp_Layout_0.VND.n64 Folded_Diff_Op_Amp_Layout_0.VND.n62 0.616779
R21270 Folded_Diff_Op_Amp_Layout_0.VND.n20 Folded_Diff_Op_Amp_Layout_0.VND.n19 0.58197
R21271 Folded_Diff_Op_Amp_Layout_0.VND.n36 Folded_Diff_Op_Amp_Layout_0.VND.t11 0.58197
R21272 Folded_Diff_Op_Amp_Layout_0.VND.n36 Folded_Diff_Op_Amp_Layout_0.VND.n35 0.58197
R21273 Folded_Diff_Op_Amp_Layout_0.VND.n32 Folded_Diff_Op_Amp_Layout_0.VND.t13 0.58197
R21274 Folded_Diff_Op_Amp_Layout_0.VND.n32 Folded_Diff_Op_Amp_Layout_0.VND.n31 0.58197
R21275 Folded_Diff_Op_Amp_Layout_0.VND.n96 Folded_Diff_Op_Amp_Layout_0.VND.t10 0.58197
R21276 Folded_Diff_Op_Amp_Layout_0.VND.n96 Folded_Diff_Op_Amp_Layout_0.VND.n95 0.58197
R21277 Folded_Diff_Op_Amp_Layout_0.VND.n70 Folded_Diff_Op_Amp_Layout_0.VND.t5 0.58197
R21278 Folded_Diff_Op_Amp_Layout_0.VND.n70 Folded_Diff_Op_Amp_Layout_0.VND.n69 0.58197
R21279 Folded_Diff_Op_Amp_Layout_0.VND.n47 Folded_Diff_Op_Amp_Layout_0.VND.t2 0.58197
R21280 Folded_Diff_Op_Amp_Layout_0.VND.n47 Folded_Diff_Op_Amp_Layout_0.VND.n46 0.58197
R21281 Folded_Diff_Op_Amp_Layout_0.VND.n51 Folded_Diff_Op_Amp_Layout_0.VND.t15 0.58197
R21282 Folded_Diff_Op_Amp_Layout_0.VND.n51 Folded_Diff_Op_Amp_Layout_0.VND.n50 0.58197
R21283 Folded_Diff_Op_Amp_Layout_0.VND.n145 Folded_Diff_Op_Amp_Layout_0.VND.n144 0.497625
R21284 Folded_Diff_Op_Amp_Layout_0.VND.n18 Folded_Diff_Op_Amp_Layout_0.VND.n10 0.3605
R21285 Folded_Diff_Op_Amp_Layout_0.VND.n4 Folded_Diff_Op_Amp_Layout_0.VND.n2 0.341925
R21286 Folded_Diff_Op_Amp_Layout_0.VND.n38 Folded_Diff_Op_Amp_Layout_0.VND.n37 0.341925
R21287 Folded_Diff_Op_Amp_Layout_0.VND.n53 Folded_Diff_Op_Amp_Layout_0.VND.n52 0.341925
R21288 Folded_Diff_Op_Amp_Layout_0.VND.n132 Folded_Diff_Op_Amp_Layout_0.VND.n131 0.330125
R21289 Folded_Diff_Op_Amp_Layout_0.VND.n129 Folded_Diff_Op_Amp_Layout_0.VND.n128 0.330125
R21290 Folded_Diff_Op_Amp_Layout_0.VND.n78 Folded_Diff_Op_Amp_Layout_0.VND.n77 0.330125
R21291 Folded_Diff_Op_Amp_Layout_0.VND.n67 Folded_Diff_Op_Amp_Layout_0.VND.n66 0.330125
R21292 Folded_Diff_Op_Amp_Layout_0.VND.n44 Folded_Diff_Op_Amp_Layout_0.VND.n43 0.330125
R21293 Folded_Diff_Op_Amp_Layout_0.VND.n21 Folded_Diff_Op_Amp_Layout_0.VND.n18 0.206051
R21294 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VND.n150 0.09825
R21295 Folded_Diff_Op_Amp_Layout_0.VND.n99 Folded_Diff_Op_Amp_Layout_0.VND.n93 0.0936537
R21296 Folded_Diff_Op_Amp_Layout_0.VND.n141 Folded_Diff_Op_Amp_Layout_0.VND.n136 0.0880141
R21297 Folded_Diff_Op_Amp_Layout_0.VND.n125 Folded_Diff_Op_Amp_Layout_0.VND.n121 0.0880141
R21298 Folded_Diff_Op_Amp_Layout_0.VND.n40 Folded_Diff_Op_Amp_Layout_0.VND.n39 0.0826464
R21299 Folded_Diff_Op_Amp_Layout_0.VND.n55 Folded_Diff_Op_Amp_Layout_0.VND.n54 0.0826464
R21300 Folded_Diff_Op_Amp_Layout_0.VND.n74 Folded_Diff_Op_Amp_Layout_0.VND.n73 0.0826464
R21301 Folded_Diff_Op_Amp_Layout_0.VND.n84 Folded_Diff_Op_Amp_Layout_0.VND.n83 0.0826464
R21302 Folded_Diff_Op_Amp_Layout_0.VND.n107 Folded_Diff_Op_Amp_Layout_0.VND.n106 0.0786497
R21303 Folded_Diff_Op_Amp_Layout_0.VND.n139 Folded_Diff_Op_Amp_Layout_0.VND.n137 0.0786471
R21304 Folded_Diff_Op_Amp_Layout_0.VND.n97 Folded_Diff_Op_Amp_Layout_0.VND.n94 0.0786471
R21305 Folded_Diff_Op_Amp_Layout_0.VND.n123 Folded_Diff_Op_Amp_Layout_0.VND.n122 0.0786471
R21306 Folded_Diff_Op_Amp_Layout_0.VND.n62 Folded_Diff_Op_Amp_Layout_0.VND.n59 0.0712285
R21307 Folded_Diff_Op_Amp_Layout_0.VND.n24 Folded_Diff_Op_Amp_Layout_0.VND.n5 0.0712285
R21308 Folded_Diff_Op_Amp_Layout_0.VND.n62 Folded_Diff_Op_Amp_Layout_0.VND.n61 0.0534597
R21309 Folded_Diff_Op_Amp_Layout_0.VND.n24 Folded_Diff_Op_Amp_Layout_0.VND.n23 0.0534597
R21310 Folded_Diff_Op_Amp_Layout_0.VND.n40 Folded_Diff_Op_Amp_Layout_0.VND.n34 0.0423164
R21311 Folded_Diff_Op_Amp_Layout_0.VND.n55 Folded_Diff_Op_Amp_Layout_0.VND.n49 0.0423164
R21312 Folded_Diff_Op_Amp_Layout_0.VND.n74 Folded_Diff_Op_Amp_Layout_0.VND.n72 0.0423164
R21313 Folded_Diff_Op_Amp_Layout_0.VND.n84 Folded_Diff_Op_Amp_Layout_0.VND.n82 0.0423164
R21314 Folded_Diff_Op_Amp_Layout_0.VND.n109 Folded_Diff_Op_Amp_Layout_0.VND.n108 0.0420655
R21315 Folded_Diff_Op_Amp_Layout_0.VND.n141 Folded_Diff_Op_Amp_Layout_0.VND.n140 0.0319869
R21316 Folded_Diff_Op_Amp_Layout_0.VND.n125 Folded_Diff_Op_Amp_Layout_0.VND.n124 0.0319869
R21317 Folded_Diff_Op_Amp_Layout_0.VND.n4 Folded_Diff_Op_Amp_Layout_0.VND.n3 0.0293873
R21318 Folded_Diff_Op_Amp_Layout_0.VND.n99 Folded_Diff_Op_Amp_Layout_0.VND.n98 0.0261793
R21319 Folded_Diff_Op_Amp_Layout_0.VND.n105 Folded_Diff_Op_Amp_Layout_0.VND.n104 0.0253684
R21320 Folded_Diff_Op_Amp_Layout_0.VND.n22 Folded_Diff_Op_Amp_Layout_0.VND.n21 0.022679
R21321 Folded_Diff_Op_Amp_Layout_0.VND.n148 Folded_Diff_Op_Amp_Layout_0.VND.n147 0.0207053
R21322 Folded_Diff_Op_Amp_Layout_0.VND.n0 Folded_Diff_Op_Amp_Layout_0.VND.n149 0.0171572
R21323 Folded_Diff_Op_Amp_Layout_0.VND.n131 Folded_Diff_Op_Amp_Layout_0.VND.n130 0.0156875
R21324 Folded_Diff_Op_Amp_Layout_0.VND.n130 Folded_Diff_Op_Amp_Layout_0.VND.n129 0.0156875
R21325 Folded_Diff_Op_Amp_Layout_0.VND.n64 Folded_Diff_Op_Amp_Layout_0.VND.n63 0.0156875
R21326 Folded_Diff_Op_Amp_Layout_0.VND.n26 Folded_Diff_Op_Amp_Layout_0.VND.n25 0.0156875
R21327 Folded_Diff_Op_Amp_Layout_0.VND.n90 Folded_Diff_Op_Amp_Layout_0.VND.n89 0.014
R21328 Folded_Diff_Op_Amp_Layout_0.VND.n149 Folded_Diff_Op_Amp_Layout_0.VND.n148 0.0134654
R21329 Folded_Diff_Op_Amp_Layout_0.VND.n135 Folded_Diff_Op_Amp_Layout_0.VND.n134 0.0133659
R21330 Folded_Diff_Op_Amp_Layout_0.VND.n120 Folded_Diff_Op_Amp_Layout_0.VND.n119 0.0133659
R21331 Folded_Diff_Op_Amp_Layout_0.VND.n133 Folded_Diff_Op_Amp_Layout_0.VND.n132 0.0111023
R21332 Folded_Diff_Op_Amp_Layout_0.VND.n118 Folded_Diff_Op_Amp_Layout_0.VND.n117 0.0111023
R21333 Folded_Diff_Op_Amp_Layout_0.VND.n113 Folded_Diff_Op_Amp_Layout_0.VND.n112 0.00958206
R21334 Folded_Diff_Op_Amp_Layout_0.VND.n27 Folded_Diff_Op_Amp_Layout_0.VND.n26 0.00860784
R21335 Folded_Diff_Op_Amp_Layout_0.VND.n143 Folded_Diff_Op_Amp_Layout_0.VND.n142 0.00860784
R21336 Folded_Diff_Op_Amp_Layout_0.VND.n127 Folded_Diff_Op_Amp_Layout_0.VND.n126 0.00860784
R21337 Folded_Diff_Op_Amp_Layout_0.VND.n65 Folded_Diff_Op_Amp_Layout_0.VND.n64 0.00860784
R21338 Folded_Diff_Op_Amp_Layout_0.VND.n116 Folded_Diff_Op_Amp_Layout_0.VND.n115 0.00858096
R21339 Folded_Diff_Op_Amp_Layout_0.VND.n115 Folded_Diff_Op_Amp_Layout_0.VND.n114 0.00858096
R21340 Folded_Diff_Op_Amp_Layout_0.VND.n114 Folded_Diff_Op_Amp_Layout_0.VND.n110 0.00858096
R21341 Folded_Diff_Op_Amp_Layout_0.VND.n86 Folded_Diff_Op_Amp_Layout_0.VND.n85 0.00858096
R21342 Folded_Diff_Op_Amp_Layout_0.VND.n79 Folded_Diff_Op_Amp_Layout_0.VND.n78 0.00858096
R21343 Folded_Diff_Op_Amp_Layout_0.VND.n76 Folded_Diff_Op_Amp_Layout_0.VND.n75 0.00858096
R21344 Folded_Diff_Op_Amp_Layout_0.VND.n68 Folded_Diff_Op_Amp_Layout_0.VND.n67 0.00858096
R21345 Folded_Diff_Op_Amp_Layout_0.VND.n87 Folded_Diff_Op_Amp_Layout_0.VND.n86 0.00858096
R21346 Folded_Diff_Op_Amp_Layout_0.VND.n85 Folded_Diff_Op_Amp_Layout_0.VND.n79 0.00858096
R21347 Folded_Diff_Op_Amp_Layout_0.VND.n77 Folded_Diff_Op_Amp_Layout_0.VND.n76 0.00858096
R21348 Folded_Diff_Op_Amp_Layout_0.VND.n75 Folded_Diff_Op_Amp_Layout_0.VND.n68 0.00858096
R21349 Folded_Diff_Op_Amp_Layout_0.VND.n57 Folded_Diff_Op_Amp_Layout_0.VND.n56 0.00858096
R21350 Folded_Diff_Op_Amp_Layout_0.VND.n45 Folded_Diff_Op_Amp_Layout_0.VND.n44 0.00858096
R21351 Folded_Diff_Op_Amp_Layout_0.VND.n42 Folded_Diff_Op_Amp_Layout_0.VND.n41 0.00858096
R21352 Folded_Diff_Op_Amp_Layout_0.VND.n30 Folded_Diff_Op_Amp_Layout_0.VND.n29 0.00858096
R21353 Folded_Diff_Op_Amp_Layout_0.VND.n58 Folded_Diff_Op_Amp_Layout_0.VND.n57 0.00858096
R21354 Folded_Diff_Op_Amp_Layout_0.VND.n56 Folded_Diff_Op_Amp_Layout_0.VND.n45 0.00858096
R21355 Folded_Diff_Op_Amp_Layout_0.VND.n43 Folded_Diff_Op_Amp_Layout_0.VND.n42 0.00858096
R21356 Folded_Diff_Op_Amp_Layout_0.VND.n41 Folded_Diff_Op_Amp_Layout_0.VND.n30 0.00858096
R21357 Folded_Diff_Op_Amp_Layout_0.VND.n144 Folded_Diff_Op_Amp_Layout_0.VND.n143 0.00855417
R21358 Folded_Diff_Op_Amp_Layout_0.VND.n128 Folded_Diff_Op_Amp_Layout_0.VND.n127 0.00855417
R21359 Folded_Diff_Op_Amp_Layout_0.VND.n66 Folded_Diff_Op_Amp_Layout_0.VND.n65 0.00855417
R21360 Folded_Diff_Op_Amp_Layout_0.VND.n28 Folded_Diff_Op_Amp_Layout_0.VND.n27 0.00855417
R21361 Folded_Diff_Op_Amp_Layout_0.VND.n146 Folded_Diff_Op_Amp_Layout_0.VND.n145 0.00773989
R21362 Folded_Diff_Op_Amp_Layout_0.VND.n136 Folded_Diff_Op_Amp_Layout_0.VND.n135 0.00642105
R21363 Folded_Diff_Op_Amp_Layout_0.VND.n93 Folded_Diff_Op_Amp_Layout_0.VND.n92 0.00642105
R21364 Folded_Diff_Op_Amp_Layout_0.VND.n121 Folded_Diff_Op_Amp_Layout_0.VND.n120 0.00642105
R21365 Folded_Diff_Op_Amp_Layout_0.VND.n106 Folded_Diff_Op_Amp_Layout_0.VND.n105 0.00642105
R21366 Folded_Diff_Op_Amp_Layout_0.VND.n112 Folded_Diff_Op_Amp_Layout_0.VND.n111 0.00642105
R21367 Folded_Diff_Op_Amp_Layout_0.VND.n126 Folded_Diff_Op_Amp_Layout_0.VND.n118 0.00605114
R21368 Folded_Diff_Op_Amp_Layout_0.VND.n142 Folded_Diff_Op_Amp_Layout_0.VND.n133 0.00605114
R21369 Folded_Diff_Op_Amp_Layout_0.VND.n92 Folded_Diff_Op_Amp_Layout_0.VND.n91 0.00551512
R21370 VCM1.n12 VCM1.t4 43.4933
R21371 VCM1.n46 VCM1.t19 39.2493
R21372 VCM1.n27 VCM1.t29 38.9885
R21373 VCM1.n33 VCM1.t0 38.877
R21374 VCM1.n52 VCM1.t22 38.6755
R21375 VCM1.n11 VCM1.t5 37.5555
R21376 VCM1.n25 VCM1.t21 36.7612
R21377 VCM1.n26 VCM1.t17 36.7612
R21378 VCM1.n38 VCM1.t26 36.5005
R21379 VCM1.n36 VCM1.t23 36.5005
R21380 VCM1.n44 VCM1.t13 36.5005
R21381 VCM1.n45 VCM1.t7 36.5005
R21382 VCM1.n48 VCM1.t10 36.2398
R21383 VCM1.n49 VCM1.t3 36.2398
R21384 VCM1.n30 VCM1.t9 35.9791
R21385 VCM1.n47 VCM1.t12 34.9362
R21386 VCM1.n50 VCM1.t24 34.9362
R21387 VCM1.n31 VCM1.t2 34.6755
R21388 VCM1.n29 VCM1.t16 32.0684
R21389 VCM1.n13 VCM1.t27 31.938
R21390 VCM1.n14 VCM1.t15 31.938
R21391 VCM1.n15 VCM1.t6 31.0255
R21392 VCM1.n12 VCM1.t28 31.0255
R21393 VCM1.n28 VCM1.t18 31.0255
R21394 VCM1.n14 VCM1.n13 20.8576
R21395 VCM1.n13 VCM1.n12 19.8148
R21396 VCM1.n15 VCM1.n14 19.8148
R21397 VCM1.n29 VCM1.n28 19.8148
R21398 VCM1.n30 VCM1.n29 18.5368
R21399 VCM1.n25 VCM1.t20 15.9041
R21400 VCM1.n26 VCM1.t8 15.9041
R21401 VCM1.n37 VCM1.n36 15.7269
R21402 VCM1.n38 VCM1.t25 15.6434
R21403 VCM1.n36 VCM1.t14 15.6434
R21404 VCM1.n44 VCM1.t11 15.6434
R21405 VCM1.n45 VCM1.t1 15.6434
R21406 VCM1.n49 VCM1.n48 14.8868
R21407 VCM1.n18 VCM1 14.8432
R21408 VCM1.n31 VCM1.n30 13.9445
R21409 VCM1.n48 VCM1.n47 13.9445
R21410 VCM1.n50 VCM1.n49 13.9445
R21411 VCM1.n32 VCM1.n25 13.9076
R21412 VCM1.n27 VCM1.n26 13.9076
R21413 VCM1.n51 VCM1.n44 13.9076
R21414 VCM1.n46 VCM1.n45 13.9076
R21415 VCM1.n39 VCM1.n38 11.2018
R21416 VCM1.n54 VCM1.n33 5.43841
R21417 VCM1.n16 VCM1.n15 4.8863
R21418 VCM1.n28 VCM1.n27 4.62659
R21419 VCM1.n47 VCM1.n46 4.62659
R21420 VCM1.n32 VCM1.n31 4.31354
R21421 VCM1.n51 VCM1.n50 4.31354
R21422 VCM1.n53 VCM1.n52 3.38239
R21423 VCM1.n53 VCM1.n43 2.39553
R21424 VCM1.n41 VCM1.n39 1.50178
R21425 VCM1.n56 VCM1.n24 1.49801
R21426 VCM1.n8 VCM1.n7 1.49801
R21427 VCM1.n18 VCM1.n17 1.49774
R21428 VCM1.n17 VCM1.n16 1.49456
R21429 VCM1.n54 VCM1.n53 1.24481
R21430 VCM1.n57 VCM1.n56 1.12725
R21431 VCM1.n57 VCM1.n3 1.12594
R21432 VCM1.n43 VCM1.n42 1.12411
R21433 VCM1.n52 VCM1.n51 0.623652
R21434 VCM1.n55 VCM1.n54 0.582814
R21435 VCM1.n21 VCM1.n20 0.582
R21436 VCM1.n33 VCM1.n32 0.36637
R21437 VCM1 VCM1.n57 0.100194
R21438 VCM1.n17 VCM1.n10 0.0301053
R21439 VCM1.n39 VCM1.n37 0.0301053
R21440 VCM1.n6 VCM1.n5 0.0207053
R21441 VCM1.n42 VCM1.n35 0.0206316
R21442 VCM1.n20 VCM1.n19 0.0156875
R21443 VCM1.n17 VCM1.n9 0.0152105
R21444 VCM1.n3 VCM1.n2 0.014
R21445 VCM1.n56 VCM1.n55 0.014
R21446 VCM1.n2 VCM1.n1 0.0134654
R21447 VCM1.n16 VCM1.n11 0.0111568
R21448 VCM1.n24 VCM1.n21 0.00998204
R21449 VCM1.n42 VCM1.n41 0.00808664
R21450 VCM1.n3 VCM1.n0 0.00773989
R21451 VCM1.n7 VCM1.n6 0.00773989
R21452 VCM1.n7 VCM1.n4 0.00773989
R21453 VCM1.n23 VCM1.n22 0.00773989
R21454 VCM1.n19 VCM1.n18 0.00638348
R21455 VCM1.n56 VCM1.n8 0.00549102
R21456 VCM1.n24 VCM1.n23 0.00549102
R21457 VCM1.n43 VCM1.n34 0.00503958
R21458 VCM1.n41 VCM1.n40 0.00455447
R21459 Folded_Diff_Op_Amp_Layout_0.VBM.n58 Folded_Diff_Op_Amp_Layout_0.VBM.t30 63.68
R21460 Folded_Diff_Op_Amp_Layout_0.VBM.n58 Folded_Diff_Op_Amp_Layout_0.VBM.t32 63.68
R21461 Folded_Diff_Op_Amp_Layout_0.VBM.n19 Folded_Diff_Op_Amp_Layout_0.VBM.t10 6.32241
R21462 Folded_Diff_Op_Amp_Layout_0.VBM.n16 Folded_Diff_Op_Amp_Layout_0.VBM.n15 6.32241
R21463 Folded_Diff_Op_Amp_Layout_0.VBM.n42 Folded_Diff_Op_Amp_Layout_0.VBM.n41 6.32241
R21464 Folded_Diff_Op_Amp_Layout_0.VBM.n34 Folded_Diff_Op_Amp_Layout_0.VBM.n33 6.32241
R21465 Folded_Diff_Op_Amp_Layout_0.VBM.n12 Folded_Diff_Op_Amp_Layout_0.VBM.n11 5.47432
R21466 Folded_Diff_Op_Amp_Layout_0.VBM.n59 Folded_Diff_Op_Amp_Layout_0.VBM.n58 5.14084
R21467 Folded_Diff_Op_Amp_Layout_0.VBM.n48 Folded_Diff_Op_Amp_Layout_0.VBM.n30 4.38115
R21468 Folded_Diff_Op_Amp_Layout_0.VBM.n23 Folded_Diff_Op_Amp_Layout_0.VBM.n22 4.38115
R21469 Folded_Diff_Op_Amp_Layout_0.VBM.n53 Folded_Diff_Op_Amp_Layout_0.VBM.n52 3.83266
R21470 Folded_Diff_Op_Amp_Layout_0.VBM.n60 Folded_Diff_Op_Amp_Layout_0.VBM.n59 3.74876
R21471 Folded_Diff_Op_Amp_Layout_0.VBM.n19 Folded_Diff_Op_Amp_Layout_0.VBM.n18 3.43224
R21472 Folded_Diff_Op_Amp_Layout_0.VBM.n16 Folded_Diff_Op_Amp_Layout_0.VBM.n14 3.43224
R21473 Folded_Diff_Op_Amp_Layout_0.VBM.n43 Folded_Diff_Op_Amp_Layout_0.VBM.n38 3.43224
R21474 Folded_Diff_Op_Amp_Layout_0.VBM.n42 Folded_Diff_Op_Amp_Layout_0.VBM.n40 3.43224
R21475 Folded_Diff_Op_Amp_Layout_0.VBM.n46 Folded_Diff_Op_Amp_Layout_0.VBM.n36 3.43224
R21476 Folded_Diff_Op_Amp_Layout_0.VBM.n34 Folded_Diff_Op_Amp_Layout_0.VBM.n32 3.43224
R21477 Folded_Diff_Op_Amp_Layout_0.VBM.n45 Folded_Diff_Op_Amp_Layout_0.VBM.n44 2.72313
R21478 Folded_Diff_Op_Amp_Layout_0.VBM.n45 Folded_Diff_Op_Amp_Layout_0.VBM.t0 2.56499
R21479 Folded_Diff_Op_Amp_Layout_0.VBM.n44 Folded_Diff_Op_Amp_Layout_0.VBM.t25 2.56298
R21480 Folded_Diff_Op_Amp_Layout_0.VBM.n26 Folded_Diff_Op_Amp_Layout_0.VBM.n12 2.12306
R21481 Folded_Diff_Op_Amp_Layout_0.VBM.n30 Folded_Diff_Op_Amp_Layout_0.VBM.t8 1.6385
R21482 Folded_Diff_Op_Amp_Layout_0.VBM.n30 Folded_Diff_Op_Amp_Layout_0.VBM.n29 1.6385
R21483 Folded_Diff_Op_Amp_Layout_0.VBM.n6 Folded_Diff_Op_Amp_Layout_0.VBM.t22 1.6385
R21484 Folded_Diff_Op_Amp_Layout_0.VBM.n6 Folded_Diff_Op_Amp_Layout_0.VBM.n5 1.6385
R21485 Folded_Diff_Op_Amp_Layout_0.VBM.n22 Folded_Diff_Op_Amp_Layout_0.VBM.t16 1.6385
R21486 Folded_Diff_Op_Amp_Layout_0.VBM.n22 Folded_Diff_Op_Amp_Layout_0.VBM.n21 1.6385
R21487 Folded_Diff_Op_Amp_Layout_0.VBM.n18 Folded_Diff_Op_Amp_Layout_0.VBM.t19 1.6385
R21488 Folded_Diff_Op_Amp_Layout_0.VBM.n18 Folded_Diff_Op_Amp_Layout_0.VBM.n17 1.6385
R21489 Folded_Diff_Op_Amp_Layout_0.VBM.n14 Folded_Diff_Op_Amp_Layout_0.VBM.t5 1.6385
R21490 Folded_Diff_Op_Amp_Layout_0.VBM.n14 Folded_Diff_Op_Amp_Layout_0.VBM.n13 1.6385
R21491 Folded_Diff_Op_Amp_Layout_0.VBM.n9 Folded_Diff_Op_Amp_Layout_0.VBM.t6 1.6385
R21492 Folded_Diff_Op_Amp_Layout_0.VBM.n9 Folded_Diff_Op_Amp_Layout_0.VBM.n8 1.6385
R21493 Folded_Diff_Op_Amp_Layout_0.VBM.n11 Folded_Diff_Op_Amp_Layout_0.VBM.t3 1.6385
R21494 Folded_Diff_Op_Amp_Layout_0.VBM.n11 Folded_Diff_Op_Amp_Layout_0.VBM.n10 1.6385
R21495 Folded_Diff_Op_Amp_Layout_0.VBM.n2 Folded_Diff_Op_Amp_Layout_0.VBM.t12 1.6385
R21496 Folded_Diff_Op_Amp_Layout_0.VBM.n2 Folded_Diff_Op_Amp_Layout_0.VBM.n1 1.6385
R21497 Folded_Diff_Op_Amp_Layout_0.VBM.n38 Folded_Diff_Op_Amp_Layout_0.VBM.t2 1.6385
R21498 Folded_Diff_Op_Amp_Layout_0.VBM.n38 Folded_Diff_Op_Amp_Layout_0.VBM.n37 1.6385
R21499 Folded_Diff_Op_Amp_Layout_0.VBM.n40 Folded_Diff_Op_Amp_Layout_0.VBM.t23 1.6385
R21500 Folded_Diff_Op_Amp_Layout_0.VBM.n40 Folded_Diff_Op_Amp_Layout_0.VBM.n39 1.6385
R21501 Folded_Diff_Op_Amp_Layout_0.VBM.n36 Folded_Diff_Op_Amp_Layout_0.VBM.t13 1.6385
R21502 Folded_Diff_Op_Amp_Layout_0.VBM.n36 Folded_Diff_Op_Amp_Layout_0.VBM.n35 1.6385
R21503 Folded_Diff_Op_Amp_Layout_0.VBM.n32 Folded_Diff_Op_Amp_Layout_0.VBM.t27 1.6385
R21504 Folded_Diff_Op_Amp_Layout_0.VBM.n32 Folded_Diff_Op_Amp_Layout_0.VBM.n31 1.6385
R21505 Folded_Diff_Op_Amp_Layout_0.VBM.n61 Folded_Diff_Op_Amp_Layout_0.VBM.n55 1.51694
R21506 Folded_Diff_Op_Amp_Layout_0.VBM.n61 Folded_Diff_Op_Amp_Layout_0.VBM.n53 1.49812
R21507 Folded_Diff_Op_Amp_Layout_0.VBM.n28 Folded_Diff_Op_Amp_Layout_0.VBM.n27 1.4921
R21508 Folded_Diff_Op_Amp_Layout_0.VBM.n44 Folded_Diff_Op_Amp_Layout_0.VBM.n43 1.44185
R21509 Folded_Diff_Op_Amp_Layout_0.VBM.n46 Folded_Diff_Op_Amp_Layout_0.VBM.n45 1.43911
R21510 Folded_Diff_Op_Amp_Layout_0.VBM.n3 Folded_Diff_Op_Amp_Layout_0.VBM.n2 1.42063
R21511 Folded_Diff_Op_Amp_Layout_0.VBM.n7 Folded_Diff_Op_Amp_Layout_0.VBM.n6 1.42054
R21512 Folded_Diff_Op_Amp_Layout_0.VBM.n27 Folded_Diff_Op_Amp_Layout_0.VBM.n7 1.15277
R21513 Folded_Diff_Op_Amp_Layout_0.VBM.n4 Folded_Diff_Op_Amp_Layout_0.VBM.n3 1.15212
R21514 Folded_Diff_Op_Amp_Layout_0.VBM.n62 Folded_Diff_Op_Amp_Layout_0.VBM.n61 1.1255
R21515 Folded_Diff_Op_Amp_Layout_0.VBM.n26 Folded_Diff_Op_Amp_Layout_0.VBM.n25 1.1255
R21516 Folded_Diff_Op_Amp_Layout_0.VBM.n51 Folded_Diff_Op_Amp_Layout_0.VBM.n50 1.1255
R21517 Folded_Diff_Op_Amp_Layout_0.VBM.n24 Folded_Diff_Op_Amp_Layout_0.VBM.n23 1.05315
R21518 Folded_Diff_Op_Amp_Layout_0.VBM.n49 Folded_Diff_Op_Amp_Layout_0.VBM.n48 1.05315
R21519 Folded_Diff_Op_Amp_Layout_0.VBM.n12 Folded_Diff_Op_Amp_Layout_0.VBM.n9 0.926316
R21520 Folded_Diff_Op_Amp_Layout_0.VBM.n59 Folded_Diff_Op_Amp_Layout_0.VBM.n57 0.715901
R21521 Folded_Diff_Op_Amp_Layout_0.VBM.n43 Folded_Diff_Op_Amp_Layout_0.VBM.n42 0.626587
R21522 Folded_Diff_Op_Amp_Layout_0.VBM.n57 Folded_Diff_Op_Amp_Layout_0.VBM.t33 0.4555
R21523 Folded_Diff_Op_Amp_Layout_0.VBM.n57 Folded_Diff_Op_Amp_Layout_0.VBM.n56 0.4555
R21524 Folded_Diff_Op_Amp_Layout_0.VBM.n20 Folded_Diff_Op_Amp_Layout_0.VBM.n16 0.323326
R21525 Folded_Diff_Op_Amp_Layout_0.VBM.n47 Folded_Diff_Op_Amp_Layout_0.VBM.n34 0.323326
R21526 Folded_Diff_Op_Amp_Layout_0.VBM.n23 Folded_Diff_Op_Amp_Layout_0.VBM.n20 0.305717
R21527 Folded_Diff_Op_Amp_Layout_0.VBM.n48 Folded_Diff_Op_Amp_Layout_0.VBM.n47 0.305717
R21528 Folded_Diff_Op_Amp_Layout_0.VBM.n20 Folded_Diff_Op_Amp_Layout_0.VBM.n19 0.303761
R21529 Folded_Diff_Op_Amp_Layout_0.VBM.n47 Folded_Diff_Op_Amp_Layout_0.VBM.n46 0.303761
R21530 Folded_Diff_Op_Amp_Layout_0.VBM.n27 Folded_Diff_Op_Amp_Layout_0.VBM.n26 0.123658
R21531 Folded_Diff_Op_Amp_Layout_0.VBM Folded_Diff_Op_Amp_Layout_0.VBM.n62 0.09825
R21532 Folded_Diff_Op_Amp_Layout_0.VBM.n52 Folded_Diff_Op_Amp_Layout_0.VBM.n51 0.0929251
R21533 Folded_Diff_Op_Amp_Layout_0.VBM.n51 Folded_Diff_Op_Amp_Layout_0.VBM.n28 0.0324737
R21534 Folded_Diff_Op_Amp_Layout_0.VBM.n52 Folded_Diff_Op_Amp_Layout_0.VBM.n4 0.0320039
R21535 Folded_Diff_Op_Amp_Layout_0.VBM.n53 Folded_Diff_Op_Amp_Layout_0.VBM.n54 0.0236139
R21536 Folded_Diff_Op_Amp_Layout_0.VBM.n25 Folded_Diff_Op_Amp_Layout_0.VBM.n24 0.014283
R21537 Folded_Diff_Op_Amp_Layout_0.VBM.n50 Folded_Diff_Op_Amp_Layout_0.VBM.n49 0.014283
R21538 Folded_Diff_Op_Amp_Layout_0.VBM.n61 Folded_Diff_Op_Amp_Layout_0.VBM.n0 0.014
R21539 Folded_Diff_Op_Amp_Layout_0.VBM.n61 Folded_Diff_Op_Amp_Layout_0.VBM.n60 0.0679038
R21540 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t0 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t2 95.9434
R21541 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t8 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t9 95.9434
R21542 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t5 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t8 95.9434
R21543 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t6 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t5 95.9434
R21544 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t11 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t12 95.9434
R21545 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t7 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t11 95.9434
R21546 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t10 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t7 95.9434
R21547 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n14 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t10 51.7088
R21548 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t0 48.1313
R21549 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n12 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t6 46.538
R21550 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n10 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n9 11.0519
R21551 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t3 4.7685
R21552 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n8 4.67159
R21553 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t1 3.3285
R21554 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n0 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n13 2.8805
R21555 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n14 2.8805
R21556 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n11 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n10 2.8805
R21557 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n16 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n4 6.88768
R21558 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n3 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n15 1.5039
R21559 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n2 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n7 1.14437
R21560 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n6 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n5 1.1255
R21561 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n3 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n16 1.11782
R21562 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n4 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n2 0.894961
R21563 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n15 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n1 0.893721
R21564 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n4 Folded_Diff_Op_Amp_Layout_0.IBIAS4.t4 3.97269
R21565 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n13 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n12 0.507444
R21566 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n0 0.128441
R21567 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n0 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n11 0.127911
R21568 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n2 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n6 0.125253
R21569 Folded_Diff_Op_Amp_Layout_0.IBIAS4 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n3 0.118134
R21570 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n16 Folded_Diff_Op_Amp_Layout_0.IBIAS4.n17 0.0459619
R21571 Folded_Diff_Op_Amp_Layout_0.IB4.n36 Folded_Diff_Op_Amp_Layout_0.IB4.t21 22.0465
R21572 Folded_Diff_Op_Amp_Layout_0.IB4.n29 Folded_Diff_Op_Amp_Layout_0.IB4.t6 14.9532
R21573 Folded_Diff_Op_Amp_Layout_0.IB4.n37 Folded_Diff_Op_Amp_Layout_0.IB4.n36 11.0965
R21574 Folded_Diff_Op_Amp_Layout_0.IB4.n38 Folded_Diff_Op_Amp_Layout_0.IB4.n37 11.0965
R21575 Folded_Diff_Op_Amp_Layout_0.IB4.n39 Folded_Diff_Op_Amp_Layout_0.IB4.n38 11.0965
R21576 Folded_Diff_Op_Amp_Layout_0.IB4.n43 Folded_Diff_Op_Amp_Layout_0.IB4.n42 11.0965
R21577 Folded_Diff_Op_Amp_Layout_0.IB4.n31 Folded_Diff_Op_Amp_Layout_0.IB4.n30 11.0965
R21578 Folded_Diff_Op_Amp_Layout_0.IB4.n36 Folded_Diff_Op_Amp_Layout_0.IB4.t19 10.9505
R21579 Folded_Diff_Op_Amp_Layout_0.IB4.n37 Folded_Diff_Op_Amp_Layout_0.IB4.t22 10.9505
R21580 Folded_Diff_Op_Amp_Layout_0.IB4.n38 Folded_Diff_Op_Amp_Layout_0.IB4.t25 10.9505
R21581 Folded_Diff_Op_Amp_Layout_0.IB4.n39 Folded_Diff_Op_Amp_Layout_0.IB4.t23 10.9505
R21582 Folded_Diff_Op_Amp_Layout_0.IB4.n42 Folded_Diff_Op_Amp_Layout_0.IB4.t0 10.9505
R21583 Folded_Diff_Op_Amp_Layout_0.IB4.n43 Folded_Diff_Op_Amp_Layout_0.IB4.t4 10.9505
R21584 Folded_Diff_Op_Amp_Layout_0.IB4.n31 Folded_Diff_Op_Amp_Layout_0.IB4.t8 10.9505
R21585 Folded_Diff_Op_Amp_Layout_0.IB4.n30 Folded_Diff_Op_Amp_Layout_0.IB4.t2 10.9505
R21586 Folded_Diff_Op_Amp_Layout_0.IB4.n41 Folded_Diff_Op_Amp_Layout_0.IB4.n39 8.67659
R21587 Folded_Diff_Op_Amp_Layout_0.IB4.n41 Folded_Diff_Op_Amp_Layout_0.IB4.n40 5.29669
R21588 Folded_Diff_Op_Amp_Layout_0.IB4.n29 Folded_Diff_Op_Amp_Layout_0.IB4.n28 4.47769
R21589 Folded_Diff_Op_Amp_Layout_0.IB4.n12 Folded_Diff_Op_Amp_Layout_0.IB4.n9 4.0405
R21590 Folded_Diff_Op_Amp_Layout_0.IB4.n30 Folded_Diff_Op_Amp_Layout_0.IB4.n29 4.00459
R21591 Folded_Diff_Op_Amp_Layout_0.IB4.n42 Folded_Diff_Op_Amp_Layout_0.IB4.n41 4.00315
R21592 Folded_Diff_Op_Amp_Layout_0.IB4.n48 Folded_Diff_Op_Amp_Layout_0.IB4.n35 3.85876
R21593 Folded_Diff_Op_Amp_Layout_0.IB4.n33 Folded_Diff_Op_Amp_Layout_0.IB4.n32 2.8805
R21594 Folded_Diff_Op_Amp_Layout_0.IB4.n45 Folded_Diff_Op_Amp_Layout_0.IB4.n44 2.8805
R21595 Folded_Diff_Op_Amp_Layout_0.IB4.n48 Folded_Diff_Op_Amp_Layout_0.IB4.n47 2.8805
R21596 Folded_Diff_Op_Amp_Layout_0.IB4.n13 Folded_Diff_Op_Amp_Layout_0.IB4.n7 2.6005
R21597 Folded_Diff_Op_Amp_Layout_0.IB4.n12 Folded_Diff_Op_Amp_Layout_0.IB4.n11 2.6005
R21598 Folded_Diff_Op_Amp_Layout_0.IB4.n44 Folded_Diff_Op_Amp_Layout_0.IB4.n43 1.7525
R21599 Folded_Diff_Op_Amp_Layout_0.IB4.n32 Folded_Diff_Op_Amp_Layout_0.IB4.n31 1.7525
R21600 Folded_Diff_Op_Amp_Layout_0.IB4.n13 Folded_Diff_Op_Amp_Layout_0.IB4.n12 1.4405
R21601 Folded_Diff_Op_Amp_Layout_0.IB4.n50 Folded_Diff_Op_Amp_Layout_0.IB4.n49 1.38361
R21602 Folded_Diff_Op_Amp_Layout_0.IB4.n3 Folded_Diff_Op_Amp_Layout_0.IB4.n2 1.26725
R21603 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IB4.n0 1.20885
R21604 Folded_Diff_Op_Amp_Layout_0.IB4.n4 Folded_Diff_Op_Amp_Layout_0.IB4.n3 1.14126
R21605 Folded_Diff_Op_Amp_Layout_0.IB4.n16 Folded_Diff_Op_Amp_Layout_0.IB4.n15 1.1255
R21606 Folded_Diff_Op_Amp_Layout_0.IB4.n19 Folded_Diff_Op_Amp_Layout_0.IB4.n18 1.1255
R21607 Folded_Diff_Op_Amp_Layout_0.IB4.n25 Folded_Diff_Op_Amp_Layout_0.IB4.n23 1.11801
R21608 Folded_Diff_Op_Amp_Layout_0.IB4.n51 Folded_Diff_Op_Amp_Layout_0.IB4.n50 1.11782
R21609 Folded_Diff_Op_Amp_Layout_0.IB4 Folded_Diff_Op_Amp_Layout_0.IB4.n52 1.07796
R21610 Folded_Diff_Op_Amp_Layout_0.IB4.n14 Folded_Diff_Op_Amp_Layout_0.IB4.n13 0.906819
R21611 Folded_Diff_Op_Amp_Layout_0.IB4.n0 Folded_Diff_Op_Amp_Layout_0.IB4.n5 0.88565
R21612 Folded_Diff_Op_Amp_Layout_0.IB4.n0 Folded_Diff_Op_Amp_Layout_0.IB4.n20 0.884803
R21613 Folded_Diff_Op_Amp_Layout_0.IB4.n35 Folded_Diff_Op_Amp_Layout_0.IB4.t5 0.8195
R21614 Folded_Diff_Op_Amp_Layout_0.IB4.n35 Folded_Diff_Op_Amp_Layout_0.IB4.n34 0.8195
R21615 Folded_Diff_Op_Amp_Layout_0.IB4.n28 Folded_Diff_Op_Amp_Layout_0.IB4.t3 0.8195
R21616 Folded_Diff_Op_Amp_Layout_0.IB4.n28 Folded_Diff_Op_Amp_Layout_0.IB4.n27 0.8195
R21617 Folded_Diff_Op_Amp_Layout_0.IB4.n7 Folded_Diff_Op_Amp_Layout_0.IB4.t14 0.607167
R21618 Folded_Diff_Op_Amp_Layout_0.IB4.n7 Folded_Diff_Op_Amp_Layout_0.IB4.n6 0.607167
R21619 Folded_Diff_Op_Amp_Layout_0.IB4.n9 Folded_Diff_Op_Amp_Layout_0.IB4.t16 0.607167
R21620 Folded_Diff_Op_Amp_Layout_0.IB4.n9 Folded_Diff_Op_Amp_Layout_0.IB4.n8 0.607167
R21621 Folded_Diff_Op_Amp_Layout_0.IB4.n2 Folded_Diff_Op_Amp_Layout_0.IB4.t13 0.607167
R21622 Folded_Diff_Op_Amp_Layout_0.IB4.n2 Folded_Diff_Op_Amp_Layout_0.IB4.n1 0.607167
R21623 Folded_Diff_Op_Amp_Layout_0.IB4.n11 Folded_Diff_Op_Amp_Layout_0.IB4.t17 0.607167
R21624 Folded_Diff_Op_Amp_Layout_0.IB4.n11 Folded_Diff_Op_Amp_Layout_0.IB4.n10 0.607167
R21625 Folded_Diff_Op_Amp_Layout_0.IB4.n48 Folded_Diff_Op_Amp_Layout_0.IB4.n46 0.0996189
R21626 Folded_Diff_Op_Amp_Layout_0.IB4.n20 Folded_Diff_Op_Amp_Layout_0.IB4.n16 0.0740848
R21627 Folded_Diff_Op_Amp_Layout_0.IB4.n49 Folded_Diff_Op_Amp_Layout_0.IB4.n48 0.0710322
R21628 Folded_Diff_Op_Amp_Layout_0.IB4.n49 Folded_Diff_Op_Amp_Layout_0.IB4.n33 0.0535557
R21629 Folded_Diff_Op_Amp_Layout_0.IB4.n20 Folded_Diff_Op_Amp_Layout_0.IB4.n19 0.0503537
R21630 Folded_Diff_Op_Amp_Layout_0.IB4.n25 Folded_Diff_Op_Amp_Layout_0.IB4.n24 0.0334577
R21631 Folded_Diff_Op_Amp_Layout_0.IB4.n18 Folded_Diff_Op_Amp_Layout_0.IB4.n17 0.0293873
R21632 Folded_Diff_Op_Amp_Layout_0.IB4.n46 Folded_Diff_Op_Amp_Layout_0.IB4.n45 0.0269989
R21633 Folded_Diff_Op_Amp_Layout_0.IB4.n5 Folded_Diff_Op_Amp_Layout_0.IB4.n4 0.0261793
R21634 Folded_Diff_Op_Amp_Layout_0.IB4.n15 Folded_Diff_Op_Amp_Layout_0.IB4.n14 0.0185116
R21635 Folded_Diff_Op_Amp_Layout_0.IB4.n23 Folded_Diff_Op_Amp_Layout_0.IB4.n21 0.0179841
R21636 Folded_Diff_Op_Amp_Layout_0.IB4.n50 Folded_Diff_Op_Amp_Layout_0.IB4.n26 0.0179841
R21637 Folded_Diff_Op_Amp_Layout_0.IB4.n23 Folded_Diff_Op_Amp_Layout_0.IB4.n22 0.0177304
R21638 Folded_Diff_Op_Amp_Layout_0.IB4.n51 Folded_Diff_Op_Amp_Layout_0.IB4.n25 0.0173591
R21639 Folded_Diff_Op_Amp_Layout_0.IB4.n52 Folded_Diff_Op_Amp_Layout_0.IB4.n51 0.0173591
R21640 a_25284_4817.t0 a_25284_4817.t1 13.3663
R21641 a_24108_3715.t0 a_24108_3715.t1 13.4632
R21642 Folded_Diff_Op_Amp_Layout_0.IVS.t80 Folded_Diff_Op_Amp_Layout_0.IVS.t79 19.5645
R21643 Folded_Diff_Op_Amp_Layout_0.IVS.t76 Folded_Diff_Op_Amp_Layout_0.IVS.t90 19.5645
R21644 Folded_Diff_Op_Amp_Layout_0.IVS.t82 Folded_Diff_Op_Amp_Layout_0.IVS.t81 19.5645
R21645 Folded_Diff_Op_Amp_Layout_0.IVS.t89 Folded_Diff_Op_Amp_Layout_0.IVS.t87 19.5645
R21646 Folded_Diff_Op_Amp_Layout_0.IVS.t85 Folded_Diff_Op_Amp_Layout_0.IVS.t83 19.5645
R21647 Folded_Diff_Op_Amp_Layout_0.IVS.t42 Folded_Diff_Op_Amp_Layout_0.IVS.t44 19.5645
R21648 Folded_Diff_Op_Amp_Layout_0.IVS.t50 Folded_Diff_Op_Amp_Layout_0.IVS.t52 19.5645
R21649 Folded_Diff_Op_Amp_Layout_0.IVS.t38 Folded_Diff_Op_Amp_Layout_0.IVS.t40 19.5645
R21650 Folded_Diff_Op_Amp_Layout_0.IVS.t46 Folded_Diff_Op_Amp_Layout_0.IVS.t48 19.5645
R21651 Folded_Diff_Op_Amp_Layout_0.IVS.t54 Folded_Diff_Op_Amp_Layout_0.IVS.t56 19.5645
R21652 Folded_Diff_Op_Amp_Layout_0.IVS.n28 Folded_Diff_Op_Amp_Layout_0.IVS.t54 13.4939
R21653 Folded_Diff_Op_Amp_Layout_0.IVS.n46 Folded_Diff_Op_Amp_Layout_0.IVS.n45 11.0965
R21654 Folded_Diff_Op_Amp_Layout_0.IVS.n45 Folded_Diff_Op_Amp_Layout_0.IVS.n44 11.0965
R21655 Folded_Diff_Op_Amp_Layout_0.IVS.n44 Folded_Diff_Op_Amp_Layout_0.IVS.n43 11.0965
R21656 Folded_Diff_Op_Amp_Layout_0.IVS.n38 Folded_Diff_Op_Amp_Layout_0.IVS.n37 11.0965
R21657 Folded_Diff_Op_Amp_Layout_0.IVS.n30 Folded_Diff_Op_Amp_Layout_0.IVS.n29 11.0965
R21658 Folded_Diff_Op_Amp_Layout_0.IVS.n18 Folded_Diff_Op_Amp_Layout_0.IVS.t80 10.987
R21659 Folded_Diff_Op_Amp_Layout_0.IVS.n46 Folded_Diff_Op_Amp_Layout_0.IVS.t76 9.4905
R21660 Folded_Diff_Op_Amp_Layout_0.IVS.n45 Folded_Diff_Op_Amp_Layout_0.IVS.t82 9.4905
R21661 Folded_Diff_Op_Amp_Layout_0.IVS.n44 Folded_Diff_Op_Amp_Layout_0.IVS.t89 9.4905
R21662 Folded_Diff_Op_Amp_Layout_0.IVS.n43 Folded_Diff_Op_Amp_Layout_0.IVS.t85 9.4905
R21663 Folded_Diff_Op_Amp_Layout_0.IVS.n38 Folded_Diff_Op_Amp_Layout_0.IVS.t42 9.4905
R21664 Folded_Diff_Op_Amp_Layout_0.IVS.n37 Folded_Diff_Op_Amp_Layout_0.IVS.t50 9.4905
R21665 Folded_Diff_Op_Amp_Layout_0.IVS.n30 Folded_Diff_Op_Amp_Layout_0.IVS.t38 9.4905
R21666 Folded_Diff_Op_Amp_Layout_0.IVS.n29 Folded_Diff_Op_Amp_Layout_0.IVS.t46 9.4905
R21667 Folded_Diff_Op_Amp_Layout_0.IVS.n43 Folded_Diff_Op_Amp_Layout_0.IVS.n42 8.67515
R21668 Folded_Diff_Op_Amp_Layout_0.IVS.n41 Folded_Diff_Op_Amp_Layout_0.IVS.n39 5.0182
R21669 Folded_Diff_Op_Amp_Layout_0.IVS.n35 Folded_Diff_Op_Amp_Layout_0.IVS.n32 4.1992
R21670 Folded_Diff_Op_Amp_Layout_0.IVS.n27 Folded_Diff_Op_Amp_Layout_0.IVS.n24 4.1992
R21671 Folded_Diff_Op_Amp_Layout_0.IVS.n92 Folded_Diff_Op_Amp_Layout_0.IVS.n89 4.0405
R21672 Folded_Diff_Op_Amp_Layout_0.IVS.n108 Folded_Diff_Op_Amp_Layout_0.IVS.n111 4.0405
R21673 Folded_Diff_Op_Amp_Layout_0.IVS.n75 Folded_Diff_Op_Amp_Layout_0.IVS.n72 4.0405
R21674 Folded_Diff_Op_Amp_Layout_0.IVS.n117 Folded_Diff_Op_Amp_Layout_0.IVS.n120 4.0405
R21675 Folded_Diff_Op_Amp_Layout_0.IVS.n126 Folded_Diff_Op_Amp_Layout_0.IVS.n129 4.0405
R21676 Folded_Diff_Op_Amp_Layout_0.IVS.n134 Folded_Diff_Op_Amp_Layout_0.IVS.n137 4.0405
R21677 Folded_Diff_Op_Amp_Layout_0.IVS.n143 Folded_Diff_Op_Amp_Layout_0.IVS.n146 4.0405
R21678 Folded_Diff_Op_Amp_Layout_0.IVS.n42 Folded_Diff_Op_Amp_Layout_0.IVS.n38 4.00459
R21679 Folded_Diff_Op_Amp_Layout_0.IVS.n36 Folded_Diff_Op_Amp_Layout_0.IVS.n30 4.00459
R21680 Folded_Diff_Op_Amp_Layout_0.IVS.n37 Folded_Diff_Op_Amp_Layout_0.IVS.n36 4.00315
R21681 Folded_Diff_Op_Amp_Layout_0.IVS.n29 Folded_Diff_Op_Amp_Layout_0.IVS.n28 4.00314
R21682 Folded_Diff_Op_Amp_Layout_0.IVS.n41 Folded_Diff_Op_Amp_Layout_0.IVS.n40 3.9695
R21683 Folded_Diff_Op_Amp_Layout_0.IVS.n35 Folded_Diff_Op_Amp_Layout_0.IVS.n34 3.1505
R21684 Folded_Diff_Op_Amp_Layout_0.IVS.n27 Folded_Diff_Op_Amp_Layout_0.IVS.n26 3.1505
R21685 Folded_Diff_Op_Amp_Layout_0.IVS.n95 Folded_Diff_Op_Amp_Layout_0.IVS.n94 2.6005
R21686 Folded_Diff_Op_Amp_Layout_0.IVS.n92 Folded_Diff_Op_Amp_Layout_0.IVS.n91 2.6005
R21687 Folded_Diff_Op_Amp_Layout_0.IVS.n108 Folded_Diff_Op_Amp_Layout_0.IVS.n109 2.6005
R21688 Folded_Diff_Op_Amp_Layout_0.IVS.n105 Folded_Diff_Op_Amp_Layout_0.IVS.n106 2.6005
R21689 Folded_Diff_Op_Amp_Layout_0.IVS.n75 Folded_Diff_Op_Amp_Layout_0.IVS.n74 2.6005
R21690 Folded_Diff_Op_Amp_Layout_0.IVS.n78 Folded_Diff_Op_Amp_Layout_0.IVS.n77 2.6005
R21691 Folded_Diff_Op_Amp_Layout_0.IVS.n117 Folded_Diff_Op_Amp_Layout_0.IVS.n118 2.6005
R21692 Folded_Diff_Op_Amp_Layout_0.IVS.n114 Folded_Diff_Op_Amp_Layout_0.IVS.n115 2.6005
R21693 Folded_Diff_Op_Amp_Layout_0.IVS.n126 Folded_Diff_Op_Amp_Layout_0.IVS.n127 2.6005
R21694 Folded_Diff_Op_Amp_Layout_0.IVS.n123 Folded_Diff_Op_Amp_Layout_0.IVS.n124 2.6005
R21695 Folded_Diff_Op_Amp_Layout_0.IVS.n134 Folded_Diff_Op_Amp_Layout_0.IVS.n135 2.6005
R21696 Folded_Diff_Op_Amp_Layout_0.IVS.n131 Folded_Diff_Op_Amp_Layout_0.IVS.n132 2.6005
R21697 Folded_Diff_Op_Amp_Layout_0.IVS.n143 Folded_Diff_Op_Amp_Layout_0.IVS.n144 2.6005
R21698 Folded_Diff_Op_Amp_Layout_0.IVS.n140 Folded_Diff_Op_Amp_Layout_0.IVS.n141 2.6005
R21699 Folded_Diff_Op_Amp_Layout_0.IVS.n0 Folded_Diff_Op_Amp_Layout_0.IVS.n67 3.547
R21700 Folded_Diff_Op_Amp_Layout_0.IVS.n10 Folded_Diff_Op_Amp_Layout_0.IVS.n60 2.40398
R21701 Folded_Diff_Op_Amp_Layout_0.IVS.n11 Folded_Diff_Op_Amp_Layout_0.IVS.n57 2.40398
R21702 Folded_Diff_Op_Amp_Layout_0.IVS.n12 Folded_Diff_Op_Amp_Layout_0.IVS.n86 2.40398
R21703 Folded_Diff_Op_Amp_Layout_0.IVS.n13 Folded_Diff_Op_Amp_Layout_0.IVS.n49 2.40398
R21704 Folded_Diff_Op_Amp_Layout_0.IVS.n14 Folded_Diff_Op_Amp_Layout_0.IVS.n99 2.40398
R21705 Folded_Diff_Op_Amp_Layout_0.IVS.n22 Folded_Diff_Op_Amp_Layout_0.IVS.n46 4.95069
R21706 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IVS.n22 1.71232
R21707 Folded_Diff_Op_Amp_Layout_0.IVS.n79 Folded_Diff_Op_Amp_Layout_0.IVS.n70 1.58214
R21708 Folded_Diff_Op_Amp_Layout_0.IVS.n22 Folded_Diff_Op_Amp_Layout_0.IVS.n17 1.49924
R21709 Folded_Diff_Op_Amp_Layout_0.IVS.n95 Folded_Diff_Op_Amp_Layout_0.IVS.n92 1.4405
R21710 Folded_Diff_Op_Amp_Layout_0.IVS.n105 Folded_Diff_Op_Amp_Layout_0.IVS.n108 1.4405
R21711 Folded_Diff_Op_Amp_Layout_0.IVS.n78 Folded_Diff_Op_Amp_Layout_0.IVS.n75 1.4405
R21712 Folded_Diff_Op_Amp_Layout_0.IVS.n114 Folded_Diff_Op_Amp_Layout_0.IVS.n117 1.4405
R21713 Folded_Diff_Op_Amp_Layout_0.IVS.n123 Folded_Diff_Op_Amp_Layout_0.IVS.n126 1.4405
R21714 Folded_Diff_Op_Amp_Layout_0.IVS.n131 Folded_Diff_Op_Amp_Layout_0.IVS.n134 1.4405
R21715 Folded_Diff_Op_Amp_Layout_0.IVS.n140 Folded_Diff_Op_Amp_Layout_0.IVS.n143 1.4405
R21716 Folded_Diff_Op_Amp_Layout_0.IVS.n19 Folded_Diff_Op_Amp_Layout_0.IVS.n20 1.4405
R21717 Folded_Diff_Op_Amp_Layout_0.IVS.n17 Folded_Diff_Op_Amp_Layout_0.IVS.n18 1.4405
R21718 Folded_Diff_Op_Amp_Layout_0.IVS.n79 Folded_Diff_Op_Amp_Layout_0.IVS.n78 1.36839
R21719 Folded_Diff_Op_Amp_Layout_0.IVS.n62 Folded_Diff_Op_Amp_Layout_0.IVS.n101 1.32
R21720 Folded_Diff_Op_Amp_Layout_0.IVS.n51 Folded_Diff_Op_Amp_Layout_0.IVS.n100 1.32
R21721 Folded_Diff_Op_Amp_Layout_0.IVS.n96 Folded_Diff_Op_Amp_Layout_0.IVS.n95 1.6095
R21722 Folded_Diff_Op_Amp_Layout_0.IVS.n104 Folded_Diff_Op_Amp_Layout_0.IVS.n105 1.30464
R21723 Folded_Diff_Op_Amp_Layout_0.IVS.n113 Folded_Diff_Op_Amp_Layout_0.IVS.n114 1.30464
R21724 Folded_Diff_Op_Amp_Layout_0.IVS.n122 Folded_Diff_Op_Amp_Layout_0.IVS.n123 1.30464
R21725 Folded_Diff_Op_Amp_Layout_0.IVS.n139 Folded_Diff_Op_Amp_Layout_0.IVS.n140 1.30464
R21726 Folded_Diff_Op_Amp_Layout_0.IVS.n42 Folded_Diff_Op_Amp_Layout_0.IVS.n41 1.24943
R21727 Folded_Diff_Op_Amp_Layout_0.IVS.n36 Folded_Diff_Op_Amp_Layout_0.IVS.n35 1.24943
R21728 Folded_Diff_Op_Amp_Layout_0.IVS.n28 Folded_Diff_Op_Amp_Layout_0.IVS.n27 1.24937
R21729 Folded_Diff_Op_Amp_Layout_0.IVS.n65 Folded_Diff_Op_Amp_Layout_0.IVS.n102 1.24927
R21730 Folded_Diff_Op_Amp_Layout_0.IVS.n54 Folded_Diff_Op_Amp_Layout_0.IVS.n103 1.24927
R21731 Folded_Diff_Op_Amp_Layout_0.IVS.n81 Folded_Diff_Op_Amp_Layout_0.IVS.n80 1.1255
R21732 Folded_Diff_Op_Amp_Layout_0.IVS.n61 Folded_Diff_Op_Amp_Layout_0.IVS.n10 1.1255
R21733 Folded_Diff_Op_Amp_Layout_0.IVS.n1 Folded_Diff_Op_Amp_Layout_0.IVS.n11 1.1255
R21734 Folded_Diff_Op_Amp_Layout_0.IVS.n6 Folded_Diff_Op_Amp_Layout_0.IVS.n12 2.03653
R21735 Folded_Diff_Op_Amp_Layout_0.IVS.n50 Folded_Diff_Op_Amp_Layout_0.IVS.n13 1.1255
R21736 Folded_Diff_Op_Amp_Layout_0.IVS.n2 Folded_Diff_Op_Amp_Layout_0.IVS.n96 1.1255
R21737 Folded_Diff_Op_Amp_Layout_0.IVS.n4 Folded_Diff_Op_Amp_Layout_0.IVS.n9 1.1255
R21738 Folded_Diff_Op_Amp_Layout_0.IVS.n3 Folded_Diff_Op_Amp_Layout_0.IVS.n14 1.1255
R21739 Folded_Diff_Op_Amp_Layout_0.IVS.n5 Folded_Diff_Op_Amp_Layout_0.IVS.n3 0.885413
R21740 Folded_Diff_Op_Amp_Layout_0.IVS.n15 Folded_Diff_Op_Amp_Layout_0.IVS.n4 0.885412
R21741 Folded_Diff_Op_Amp_Layout_0.IVS.n6 Folded_Diff_Op_Amp_Layout_0.IVS.n131 3.53561
R21742 Folded_Diff_Op_Amp_Layout_0.IVS.n26 Folded_Diff_Op_Amp_Layout_0.IVS.t47 0.8195
R21743 Folded_Diff_Op_Amp_Layout_0.IVS.n26 Folded_Diff_Op_Amp_Layout_0.IVS.n25 0.8195
R21744 Folded_Diff_Op_Amp_Layout_0.IVS.n34 Folded_Diff_Op_Amp_Layout_0.IVS.t51 0.8195
R21745 Folded_Diff_Op_Amp_Layout_0.IVS.n34 Folded_Diff_Op_Amp_Layout_0.IVS.n33 0.8195
R21746 Folded_Diff_Op_Amp_Layout_0.IVS.n32 Folded_Diff_Op_Amp_Layout_0.IVS.t53 0.8195
R21747 Folded_Diff_Op_Amp_Layout_0.IVS.n32 Folded_Diff_Op_Amp_Layout_0.IVS.n31 0.8195
R21748 Folded_Diff_Op_Amp_Layout_0.IVS.n24 Folded_Diff_Op_Amp_Layout_0.IVS.t49 0.8195
R21749 Folded_Diff_Op_Amp_Layout_0.IVS.n24 Folded_Diff_Op_Amp_Layout_0.IVS.n23 0.8195
R21750 Folded_Diff_Op_Amp_Layout_0.IVS.n68 Folded_Diff_Op_Amp_Layout_0.IVS.n0 0.736713
R21751 Folded_Diff_Op_Amp_Layout_0.IVS.n8 Folded_Diff_Op_Amp_Layout_0.IVS.n1 0.727165
R21752 Folded_Diff_Op_Amp_Layout_0.IVS.n7 Folded_Diff_Op_Amp_Layout_0.IVS.n62 0.616779
R21753 Folded_Diff_Op_Amp_Layout_0.IVS.n16 Folded_Diff_Op_Amp_Layout_0.IVS.n51 0.616779
R21754 Folded_Diff_Op_Amp_Layout_0.IVS.n89 Folded_Diff_Op_Amp_Layout_0.IVS.t24 0.607167
R21755 Folded_Diff_Op_Amp_Layout_0.IVS.n89 Folded_Diff_Op_Amp_Layout_0.IVS.n88 0.607167
R21756 Folded_Diff_Op_Amp_Layout_0.IVS.n91 Folded_Diff_Op_Amp_Layout_0.IVS.t23 0.607167
R21757 Folded_Diff_Op_Amp_Layout_0.IVS.n91 Folded_Diff_Op_Amp_Layout_0.IVS.n90 0.607167
R21758 Folded_Diff_Op_Amp_Layout_0.IVS.n94 Folded_Diff_Op_Amp_Layout_0.IVS.t3 0.607167
R21759 Folded_Diff_Op_Amp_Layout_0.IVS.n94 Folded_Diff_Op_Amp_Layout_0.IVS.n93 0.607167
R21760 Folded_Diff_Op_Amp_Layout_0.IVS.n99 Folded_Diff_Op_Amp_Layout_0.IVS.t63 0.607167
R21761 Folded_Diff_Op_Amp_Layout_0.IVS.n99 Folded_Diff_Op_Amp_Layout_0.IVS.n98 0.607167
R21762 Folded_Diff_Op_Amp_Layout_0.IVS.n67 Folded_Diff_Op_Amp_Layout_0.IVS.t26 0.607167
R21763 Folded_Diff_Op_Amp_Layout_0.IVS.n67 Folded_Diff_Op_Amp_Layout_0.IVS.n66 0.607167
R21764 Folded_Diff_Op_Amp_Layout_0.IVS.n106 Folded_Diff_Op_Amp_Layout_0.IVS.t61 0.607167
R21765 Folded_Diff_Op_Amp_Layout_0.IVS.n106 Folded_Diff_Op_Amp_Layout_0.IVS.n107 0.607167
R21766 Folded_Diff_Op_Amp_Layout_0.IVS.n109 Folded_Diff_Op_Amp_Layout_0.IVS.t37 0.607167
R21767 Folded_Diff_Op_Amp_Layout_0.IVS.n109 Folded_Diff_Op_Amp_Layout_0.IVS.n110 0.607167
R21768 Folded_Diff_Op_Amp_Layout_0.IVS.n111 Folded_Diff_Op_Amp_Layout_0.IVS.t18 0.607167
R21769 Folded_Diff_Op_Amp_Layout_0.IVS.n111 Folded_Diff_Op_Amp_Layout_0.IVS.n112 0.607167
R21770 Folded_Diff_Op_Amp_Layout_0.IVS.n70 Folded_Diff_Op_Amp_Layout_0.IVS.t66 0.607167
R21771 Folded_Diff_Op_Amp_Layout_0.IVS.n70 Folded_Diff_Op_Amp_Layout_0.IVS.n69 0.607167
R21772 Folded_Diff_Op_Amp_Layout_0.IVS.n77 Folded_Diff_Op_Amp_Layout_0.IVS.t27 0.607167
R21773 Folded_Diff_Op_Amp_Layout_0.IVS.n77 Folded_Diff_Op_Amp_Layout_0.IVS.n76 0.607167
R21774 Folded_Diff_Op_Amp_Layout_0.IVS.n74 Folded_Diff_Op_Amp_Layout_0.IVS.t69 0.607167
R21775 Folded_Diff_Op_Amp_Layout_0.IVS.n74 Folded_Diff_Op_Amp_Layout_0.IVS.n73 0.607167
R21776 Folded_Diff_Op_Amp_Layout_0.IVS.n72 Folded_Diff_Op_Amp_Layout_0.IVS.t70 0.607167
R21777 Folded_Diff_Op_Amp_Layout_0.IVS.n72 Folded_Diff_Op_Amp_Layout_0.IVS.n71 0.607167
R21778 Folded_Diff_Op_Amp_Layout_0.IVS.n60 Folded_Diff_Op_Amp_Layout_0.IVS.t14 0.607167
R21779 Folded_Diff_Op_Amp_Layout_0.IVS.n60 Folded_Diff_Op_Amp_Layout_0.IVS.n59 0.607167
R21780 Folded_Diff_Op_Amp_Layout_0.IVS.n115 Folded_Diff_Op_Amp_Layout_0.IVS.t72 0.607167
R21781 Folded_Diff_Op_Amp_Layout_0.IVS.n115 Folded_Diff_Op_Amp_Layout_0.IVS.n116 0.607167
R21782 Folded_Diff_Op_Amp_Layout_0.IVS.n118 Folded_Diff_Op_Amp_Layout_0.IVS.t0 0.607167
R21783 Folded_Diff_Op_Amp_Layout_0.IVS.n118 Folded_Diff_Op_Amp_Layout_0.IVS.n119 0.607167
R21784 Folded_Diff_Op_Amp_Layout_0.IVS.n120 Folded_Diff_Op_Amp_Layout_0.IVS.t1 0.607167
R21785 Folded_Diff_Op_Amp_Layout_0.IVS.n120 Folded_Diff_Op_Amp_Layout_0.IVS.n121 0.607167
R21786 Folded_Diff_Op_Amp_Layout_0.IVS.n57 Folded_Diff_Op_Amp_Layout_0.IVS.t62 0.607167
R21787 Folded_Diff_Op_Amp_Layout_0.IVS.n57 Folded_Diff_Op_Amp_Layout_0.IVS.n56 0.607167
R21788 Folded_Diff_Op_Amp_Layout_0.IVS.n124 Folded_Diff_Op_Amp_Layout_0.IVS.t2 0.607167
R21789 Folded_Diff_Op_Amp_Layout_0.IVS.n124 Folded_Diff_Op_Amp_Layout_0.IVS.n125 0.607167
R21790 Folded_Diff_Op_Amp_Layout_0.IVS.n127 Folded_Diff_Op_Amp_Layout_0.IVS.t21 0.607167
R21791 Folded_Diff_Op_Amp_Layout_0.IVS.n127 Folded_Diff_Op_Amp_Layout_0.IVS.n128 0.607167
R21792 Folded_Diff_Op_Amp_Layout_0.IVS.n129 Folded_Diff_Op_Amp_Layout_0.IVS.t22 0.607167
R21793 Folded_Diff_Op_Amp_Layout_0.IVS.n129 Folded_Diff_Op_Amp_Layout_0.IVS.n130 0.607167
R21794 Folded_Diff_Op_Amp_Layout_0.IVS.n86 Folded_Diff_Op_Amp_Layout_0.IVS.t25 0.607167
R21795 Folded_Diff_Op_Amp_Layout_0.IVS.n86 Folded_Diff_Op_Amp_Layout_0.IVS.n85 0.607167
R21796 Folded_Diff_Op_Amp_Layout_0.IVS.n132 Folded_Diff_Op_Amp_Layout_0.IVS.t60 0.607167
R21797 Folded_Diff_Op_Amp_Layout_0.IVS.n132 Folded_Diff_Op_Amp_Layout_0.IVS.n133 0.607167
R21798 Folded_Diff_Op_Amp_Layout_0.IVS.n135 Folded_Diff_Op_Amp_Layout_0.IVS.t36 0.607167
R21799 Folded_Diff_Op_Amp_Layout_0.IVS.n135 Folded_Diff_Op_Amp_Layout_0.IVS.n136 0.607167
R21800 Folded_Diff_Op_Amp_Layout_0.IVS.n137 Folded_Diff_Op_Amp_Layout_0.IVS.t17 0.607167
R21801 Folded_Diff_Op_Amp_Layout_0.IVS.n137 Folded_Diff_Op_Amp_Layout_0.IVS.n138 0.607167
R21802 Folded_Diff_Op_Amp_Layout_0.IVS.n49 Folded_Diff_Op_Amp_Layout_0.IVS.t71 0.607167
R21803 Folded_Diff_Op_Amp_Layout_0.IVS.n49 Folded_Diff_Op_Amp_Layout_0.IVS.n48 0.607167
R21804 Folded_Diff_Op_Amp_Layout_0.IVS.n141 Folded_Diff_Op_Amp_Layout_0.IVS.t19 0.607167
R21805 Folded_Diff_Op_Amp_Layout_0.IVS.n141 Folded_Diff_Op_Amp_Layout_0.IVS.n142 0.607167
R21806 Folded_Diff_Op_Amp_Layout_0.IVS.n144 Folded_Diff_Op_Amp_Layout_0.IVS.t12 0.607167
R21807 Folded_Diff_Op_Amp_Layout_0.IVS.n144 Folded_Diff_Op_Amp_Layout_0.IVS.n145 0.607167
R21808 Folded_Diff_Op_Amp_Layout_0.IVS.n146 Folded_Diff_Op_Amp_Layout_0.IVS.t13 0.607167
R21809 Folded_Diff_Op_Amp_Layout_0.IVS.n146 Folded_Diff_Op_Amp_Layout_0.IVS.n147 0.607167
R21810 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IVS.n5 0.402965
R21811 Folded_Diff_Op_Amp_Layout_0.IVS.n13 Folded_Diff_Op_Amp_Layout_0.IVS.n47 0.21657
R21812 Folded_Diff_Op_Amp_Layout_0.IVS.n12 Folded_Diff_Op_Amp_Layout_0.IVS.n84 0.21657
R21813 Folded_Diff_Op_Amp_Layout_0.IVS.n11 Folded_Diff_Op_Amp_Layout_0.IVS.n55 0.21657
R21814 Folded_Diff_Op_Amp_Layout_0.IVS.n10 Folded_Diff_Op_Amp_Layout_0.IVS.n58 0.21657
R21815 Folded_Diff_Op_Amp_Layout_0.IVS.n9 Folded_Diff_Op_Amp_Layout_0.IVS.n83 0.198558
R21816 Folded_Diff_Op_Amp_Layout_0.IVS.n102 Folded_Diff_Op_Amp_Layout_0.IVS.n104 0.181594
R21817 Folded_Diff_Op_Amp_Layout_0.IVS.n101 Folded_Diff_Op_Amp_Layout_0.IVS.n113 0.181594
R21818 Folded_Diff_Op_Amp_Layout_0.IVS.n103 Folded_Diff_Op_Amp_Layout_0.IVS.n122 0.181594
R21819 Folded_Diff_Op_Amp_Layout_0.IVS.n100 Folded_Diff_Op_Amp_Layout_0.IVS.n139 0.181594
R21820 Folded_Diff_Op_Amp_Layout_0.IVS.n3 Folded_Diff_Op_Amp_Layout_0.IVS.n2 0.125253
R21821 Folded_Diff_Op_Amp_Layout_0.IVS.n5 Folded_Diff_Op_Amp_Layout_0.IVS.n16 0.114434
R21822 Folded_Diff_Op_Amp_Layout_0.IVS.n80 Folded_Diff_Op_Amp_Layout_0.IVS.n79 0.114284
R21823 Folded_Diff_Op_Amp_Layout_0.IVS.n16 Folded_Diff_Op_Amp_Layout_0.IVS.n6 0.11344
R21824 Folded_Diff_Op_Amp_Layout_0.IVS.n14 Folded_Diff_Op_Amp_Layout_0.IVS.n97 0.113394
R21825 Folded_Diff_Op_Amp_Layout_0.IVS.n6 Folded_Diff_Op_Amp_Layout_0.IVS.n8 0.103892
R21826 Folded_Diff_Op_Amp_Layout_0.IVS.n8 Folded_Diff_Op_Amp_Layout_0.IVS.n7 0.10389
R21827 Folded_Diff_Op_Amp_Layout_0.IVS.n7 Folded_Diff_Op_Amp_Layout_0.IVS.n15 0.0953406
R21828 Folded_Diff_Op_Amp_Layout_0.IVS.n15 Folded_Diff_Op_Amp_Layout_0.IVS.n68 0.0943399
R21829 Folded_Diff_Op_Amp_Layout_0.IVS.n9 Folded_Diff_Op_Amp_Layout_0.IVS.n82 0.0800906
R21830 Folded_Diff_Op_Amp_Layout_0.IVS.n65 Folded_Diff_Op_Amp_Layout_0.IVS.n64 0.0625655
R21831 Folded_Diff_Op_Amp_Layout_0.IVS.n54 Folded_Diff_Op_Amp_Layout_0.IVS.n53 0.0625655
R21832 Folded_Diff_Op_Amp_Layout_0.IVS.n64 Folded_Diff_Op_Amp_Layout_0.IVS.n63 0.0625188
R21833 Folded_Diff_Op_Amp_Layout_0.IVS.n53 Folded_Diff_Op_Amp_Layout_0.IVS.n52 0.0625188
R21834 Folded_Diff_Op_Amp_Layout_0.IVS.n4 Folded_Diff_Op_Amp_Layout_0.IVS.n81 0.249023
R21835 Folded_Diff_Op_Amp_Layout_0.IVS.n2 Folded_Diff_Op_Amp_Layout_0.IVS.n87 0.125422
R21836 Folded_Diff_Op_Amp_Layout_0.IVS.n1 Folded_Diff_Op_Amp_Layout_0.IVS.n54 0.124472
R21837 Folded_Diff_Op_Amp_Layout_0.IVS.n0 Folded_Diff_Op_Amp_Layout_0.IVS.n65 0.124472
R21838 Folded_Diff_Op_Amp_Layout_0.IVS.n62 Folded_Diff_Op_Amp_Layout_0.IVS.n61 0.0534597
R21839 Folded_Diff_Op_Amp_Layout_0.IVS.n51 Folded_Diff_Op_Amp_Layout_0.IVS.n50 0.0534597
R21840 Folded_Diff_Op_Amp_Layout_0.IVS.n17 Folded_Diff_Op_Amp_Layout_0.IVS.n19 0.0492192
R21841 Folded_Diff_Op_Amp_Layout_0.IVS.n22 Folded_Diff_Op_Amp_Layout_0.IVS.n21 0.0471546
R21842 Folded_Diff_Op_Amp_Layout_0.IBS.n4 Folded_Diff_Op_Amp_Layout_0.IBS.t10 15.4765
R21843 Folded_Diff_Op_Amp_Layout_0.IBS.n5 Folded_Diff_Op_Amp_Layout_0.IBS.n4 11.0965
R21844 Folded_Diff_Op_Amp_Layout_0.IBS Folded_Diff_Op_Amp_Layout_0.IBS.n1 8.10022
R21845 Folded_Diff_Op_Amp_Layout_0.IBS.n3 Folded_Diff_Op_Amp_Layout_0.IBS.t3 7.191
R21846 Folded_Diff_Op_Amp_Layout_0.IBS.n16 Folded_Diff_Op_Amp_Layout_0.IBS.t8 4.76941
R21847 Folded_Diff_Op_Amp_Layout_0.IBS.n6 Folded_Diff_Op_Amp_Layout_0.IBS.n5 4.49
R21848 Folded_Diff_Op_Amp_Layout_0.IBS.n4 Folded_Diff_Op_Amp_Layout_0.IBS.t11 4.3805
R21849 Folded_Diff_Op_Amp_Layout_0.IBS.n5 Folded_Diff_Op_Amp_Layout_0.IBS.t5 4.3805
R21850 Folded_Diff_Op_Amp_Layout_0.IBS.n16 Folded_Diff_Op_Amp_Layout_0.IBS.n15 3.4692
R21851 Folded_Diff_Op_Amp_Layout_0.IBS.n2 Folded_Diff_Op_Amp_Layout_0.IBS.n9 3.42896
R21852 Folded_Diff_Op_Amp_Layout_0.IBS.n9 Folded_Diff_Op_Amp_Layout_0.IBS.t4 1.6385
R21853 Folded_Diff_Op_Amp_Layout_0.IBS.n9 Folded_Diff_Op_Amp_Layout_0.IBS.n8 1.6385
R21854 Folded_Diff_Op_Amp_Layout_0.IBS.n17 Folded_Diff_Op_Amp_Layout_0.IBS.n16 1.6365
R21855 Folded_Diff_Op_Amp_Layout_0.IBS Folded_Diff_Op_Amp_Layout_0.IBS.n10 1.61193
R21856 Folded_Diff_Op_Amp_Layout_0.IBS.n13 Folded_Diff_Op_Amp_Layout_0.IBS.n12 1.18193
R21857 Folded_Diff_Op_Amp_Layout_0.IBS.n1 Folded_Diff_Op_Amp_Layout_0.IBS.n13 1.17273
R21858 Folded_Diff_Op_Amp_Layout_0.IBS.n7 Folded_Diff_Op_Amp_Layout_0.IBS.n6 1.14565
R21859 Folded_Diff_Op_Amp_Layout_0.IBS.n7 Folded_Diff_Op_Amp_Layout_0.IBS.n3 1.14531
R21860 Folded_Diff_Op_Amp_Layout_0.IBS.n0 Folded_Diff_Op_Amp_Layout_0.IBS.n18 1.1255
R21861 Folded_Diff_Op_Amp_Layout_0.IBS.n2 Folded_Diff_Op_Amp_Layout_0.IBS.n7 0.869271
R21862 Folded_Diff_Op_Amp_Layout_0.IBS.n18 Folded_Diff_Op_Amp_Layout_0.IBS.n17 0.546716
R21863 Folded_Diff_Op_Amp_Layout_0.IBS.n15 Folded_Diff_Op_Amp_Layout_0.IBS.t1 0.4555
R21864 Folded_Diff_Op_Amp_Layout_0.IBS.n15 Folded_Diff_Op_Amp_Layout_0.IBS.n14 0.4555
R21865 Folded_Diff_Op_Amp_Layout_0.IBS.n12 Folded_Diff_Op_Amp_Layout_0.IBS.t0 0.4555
R21866 Folded_Diff_Op_Amp_Layout_0.IBS.n12 Folded_Diff_Op_Amp_Layout_0.IBS.n11 0.4555
R21867 Folded_Diff_Op_Amp_Layout_0.IBS.n1 Folded_Diff_Op_Amp_Layout_0.IBS.n0 0.125254
R21868 Folded_Diff_Op_Amp_Layout_0.IBS.n10 Folded_Diff_Op_Amp_Layout_0.IBS.n2 0.259993
R21869 a_24836_4817.t0 a_24836_4817.t1 13.4632
R21870 a_26012_3715.t0 a_26012_3715.t1 13.3663
R21871 Folded_Diff_Op_Amp_Layout_0.VBIASN.n16 Folded_Diff_Op_Amp_Layout_0.VBIASN.t12 25.1953
R21872 Folded_Diff_Op_Amp_Layout_0.VBIASN.n9 Folded_Diff_Op_Amp_Layout_0.VBIASN.n8 14.0791
R21873 Folded_Diff_Op_Amp_Layout_0.VBIASN.n10 Folded_Diff_Op_Amp_Layout_0.VBIASN.n9 14.0791
R21874 Folded_Diff_Op_Amp_Layout_0.VBIASN.n11 Folded_Diff_Op_Amp_Layout_0.VBIASN.n10 14.0791
R21875 Folded_Diff_Op_Amp_Layout_0.VBIASN.n12 Folded_Diff_Op_Amp_Layout_0.VBIASN.n11 14.0791
R21876 Folded_Diff_Op_Amp_Layout_0.VBIASN.n13 Folded_Diff_Op_Amp_Layout_0.VBIASN.n12 14.0791
R21877 Folded_Diff_Op_Amp_Layout_0.VBIASN.n14 Folded_Diff_Op_Amp_Layout_0.VBIASN.n13 14.0791
R21878 Folded_Diff_Op_Amp_Layout_0.VBIASN.n3 Folded_Diff_Op_Amp_Layout_0.VBIASN.t5 13.5278
R21879 Folded_Diff_Op_Amp_Layout_0.VBIASN.n7 Folded_Diff_Op_Amp_Layout_0.VBIASN.t3 11.2226
R21880 Folded_Diff_Op_Amp_Layout_0.VBIASN.n15 Folded_Diff_Op_Amp_Layout_0.VBIASN.n14 8.47371
R21881 Folded_Diff_Op_Amp_Layout_0.VBIASN.n14 Folded_Diff_Op_Amp_Layout_0.VBIASN.t10 7.82193
R21882 Folded_Diff_Op_Amp_Layout_0.VBIASN.n13 Folded_Diff_Op_Amp_Layout_0.VBIASN.t9 7.82193
R21883 Folded_Diff_Op_Amp_Layout_0.VBIASN.n12 Folded_Diff_Op_Amp_Layout_0.VBIASN.t11 7.82193
R21884 Folded_Diff_Op_Amp_Layout_0.VBIASN.n11 Folded_Diff_Op_Amp_Layout_0.VBIASN.t8 7.82193
R21885 Folded_Diff_Op_Amp_Layout_0.VBIASN.n10 Folded_Diff_Op_Amp_Layout_0.VBIASN.t7 7.82193
R21886 Folded_Diff_Op_Amp_Layout_0.VBIASN.n9 Folded_Diff_Op_Amp_Layout_0.VBIASN.t13 7.82193
R21887 Folded_Diff_Op_Amp_Layout_0.VBIASN.n8 Folded_Diff_Op_Amp_Layout_0.VBIASN.t1 7.82193
R21888 Folded_Diff_Op_Amp_Layout_0.VBIASN.n3 Folded_Diff_Op_Amp_Layout_0.VBIASN.n15 4.48087
R21889 Folded_Diff_Op_Amp_Layout_0.VBIASN.n7 Folded_Diff_Op_Amp_Layout_0.VBIASN.n6 3.82142
R21890 Folded_Diff_Op_Amp_Layout_0.VBIASN.n8 Folded_Diff_Op_Amp_Layout_0.VBIASN.n7 3.3996
R21891 Folded_Diff_Op_Amp_Layout_0.VBIASN.n0 Folded_Diff_Op_Amp_Layout_0.VBIASN.n2 3.2818
R21892 Folded_Diff_Op_Amp_Layout_0.VBIASN Folded_Diff_Op_Amp_Layout_0.VBIASN.n0 2.27678
R21893 Folded_Diff_Op_Amp_Layout_0.VBIASN.n6 Folded_Diff_Op_Amp_Layout_0.VBIASN.t4 1.6385
R21894 Folded_Diff_Op_Amp_Layout_0.VBIASN.n6 Folded_Diff_Op_Amp_Layout_0.VBIASN.n5 1.6385
R21895 Folded_Diff_Op_Amp_Layout_0.VBIASN.n0 Folded_Diff_Op_Amp_Layout_0.VBIASN.n17 1.48953
R21896 Folded_Diff_Op_Amp_Layout_0.VBIASN.n4 Folded_Diff_Op_Amp_Layout_0.VBIASN.t0 1.47411
R21897 Folded_Diff_Op_Amp_Layout_0.VBIASN.n16 Folded_Diff_Op_Amp_Layout_0.VBIASN.n3 1.27179
R21898 Folded_Diff_Op_Amp_Layout_0.VBIASN.n2 Folded_Diff_Op_Amp_Layout_0.VBIASN.n4 1.16684
R21899 Folded_Diff_Op_Amp_Layout_0.VBIASN.n0 Folded_Diff_Op_Amp_Layout_0.VBIASN.n16 0.313311
R21900 Folded_Diff_Op_Amp_Layout_0.VBIASN.n2 Folded_Diff_Op_Amp_Layout_0.VBIASN.n1 0.124429
R21901 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t13 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t0 82.1255
R21902 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n3 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t4 49.4342
R21903 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n13 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t2 42.7576
R21904 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t12 42.7576
R21905 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t0 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n3 29.7219
R21906 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n13 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t3 28.6791
R21907 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n10 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t14 28.6791
R21908 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t10 28.6791
R21909 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t7 28.6791
R21910 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n7 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t8 28.6791
R21911 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n6 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t6 28.6791
R21912 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n5 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t5 28.6791
R21913 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t11 28.6791
R21914 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n4 Folded_Diff_Op_Amp_Layout_0.IBIAS1.t13 28.6791
R21915 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n4 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n1 14.0791
R21916 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n5 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n4 14.0791
R21917 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n6 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n5 14.0791
R21918 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n7 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n6 14.0791
R21919 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n7 14.0791
R21920 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n8 14.0791
R21921 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n10 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n9 14.0791
R21922 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n3 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n2 8.09246
R21923 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n11 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n10 7.3005
R21924 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n12 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n11 2.8805
R21925 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n14 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n13 2.8805
R21926 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n0 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n12 1.50421
R21927 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n0 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n14 1.50283
R21928 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n0 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n15 1.48384
R21929 Folded_Diff_Op_Amp_Layout_0.IBIAS1 Folded_Diff_Op_Amp_Layout_0.IBIAS1.n0 1.05318
R21930 VIN_N1 VIN_N1.t0 5.04285
R21931 a_n5986_5540.t0 a_n5986_5540.t1 14.4367
R21932 a_29734_1647.t0 a_29734_1647.t1 9.25328
R21933 a_n5706_9350.t0 a_n5706_9350.t1 13.5425
R21934 a_n6266_8788.t0 a_n6266_8788.t1 13.5425
R21935 filter_res_magic_0.R7_R8_R10_C filter_res_magic_0.R7_R8_R10_C.t0 4.51219
R21936 a_n6826_5540.t0 a_n6826_5540.t1 13.5425
R21937 Folded_Diff_Op_Amp_Layout_0.VB4.n58 Folded_Diff_Op_Amp_Layout_0.VB4.t67 52.1434
R21938 Folded_Diff_Op_Amp_Layout_0.VB4.n57 Folded_Diff_Op_Amp_Layout_0.VB4.t68 52.1434
R21939 Folded_Diff_Op_Amp_Layout_0.VB4.n56 Folded_Diff_Op_Amp_Layout_0.VB4.t84 52.1434
R21940 Folded_Diff_Op_Amp_Layout_0.VB4.n55 Folded_Diff_Op_Amp_Layout_0.VB4.t89 52.1434
R21941 Folded_Diff_Op_Amp_Layout_0.VB4.n54 Folded_Diff_Op_Amp_Layout_0.VB4.t41 52.1434
R21942 Folded_Diff_Op_Amp_Layout_0.VB4.n53 Folded_Diff_Op_Amp_Layout_0.VB4.t37 52.1434
R21943 Folded_Diff_Op_Amp_Layout_0.VB4.n52 Folded_Diff_Op_Amp_Layout_0.VB4.t40 52.1434
R21944 Folded_Diff_Op_Amp_Layout_0.VB4.t79 Folded_Diff_Op_Amp_Layout_0.VB4.n12 51.2309
R21945 Folded_Diff_Op_Amp_Layout_0.VB4.t94 Folded_Diff_Op_Amp_Layout_0.VB4.n16 51.2309
R21946 Folded_Diff_Op_Amp_Layout_0.VB4.t48 Folded_Diff_Op_Amp_Layout_0.VB4.n17 51.2309
R21947 Folded_Diff_Op_Amp_Layout_0.VB4.t63 Folded_Diff_Op_Amp_Layout_0.VB4.n31 51.2309
R21948 Folded_Diff_Op_Amp_Layout_0.VB4.t56 Folded_Diff_Op_Amp_Layout_0.VB4.n13 50.188
R21949 Folded_Diff_Op_Amp_Layout_0.VB4.t69 Folded_Diff_Op_Amp_Layout_0.VB4.n21 50.188
R21950 Folded_Diff_Op_Amp_Layout_0.VB4.t33 Folded_Diff_Op_Amp_Layout_0.VB4.n32 50.188
R21951 Folded_Diff_Op_Amp_Layout_0.VB4.t60 Folded_Diff_Op_Amp_Layout_0.VB4.n36 50.188
R21952 Folded_Diff_Op_Amp_Layout_0.VB4.t46 Folded_Diff_Op_Amp_Layout_0.VB4.n51 49.6666
R21953 Folded_Diff_Op_Amp_Layout_0.VB4.t97 Folded_Diff_Op_Amp_Layout_0.VB4.n28 48.8844
R21954 Folded_Diff_Op_Amp_Layout_0.VB4.t70 Folded_Diff_Op_Amp_Layout_0.VB4.n42 48.8844
R21955 Folded_Diff_Op_Amp_Layout_0.VB4.t88 Folded_Diff_Op_Amp_Layout_0.VB4.n43 48.8844
R21956 Folded_Diff_Op_Amp_Layout_0.VB4.t42 Folded_Diff_Op_Amp_Layout_0.VB4.n23 48.6237
R21957 Folded_Diff_Op_Amp_Layout_0.VB4.t95 Folded_Diff_Op_Amp_Layout_0.VB4.n25 48.6237
R21958 Folded_Diff_Op_Amp_Layout_0.VB4.t77 Folded_Diff_Op_Amp_Layout_0.VB4.n34 48.6237
R21959 Folded_Diff_Op_Amp_Layout_0.VB4.t45 Folded_Diff_Op_Amp_Layout_0.VB4.n38 48.6237
R21960 Folded_Diff_Op_Amp_Layout_0.VB4.n23 Folded_Diff_Op_Amp_Layout_0.VB4.t56 48.1023
R21961 Folded_Diff_Op_Amp_Layout_0.VB4.n22 Folded_Diff_Op_Amp_Layout_0.VB4.t69 48.1023
R21962 Folded_Diff_Op_Amp_Layout_0.VB4.n25 Folded_Diff_Op_Amp_Layout_0.VB4.t36 48.1023
R21963 Folded_Diff_Op_Amp_Layout_0.VB4.n24 Folded_Diff_Op_Amp_Layout_0.VB4.t53 48.1023
R21964 Folded_Diff_Op_Amp_Layout_0.VB4.n34 Folded_Diff_Op_Amp_Layout_0.VB4.t87 48.1023
R21965 Folded_Diff_Op_Amp_Layout_0.VB4.n33 Folded_Diff_Op_Amp_Layout_0.VB4.t33 48.1023
R21966 Folded_Diff_Op_Amp_Layout_0.VB4.n37 Folded_Diff_Op_Amp_Layout_0.VB4.t99 48.1023
R21967 Folded_Diff_Op_Amp_Layout_0.VB4.n38 Folded_Diff_Op_Amp_Layout_0.VB4.t60 48.1023
R21968 Folded_Diff_Op_Amp_Layout_0.VB4.n28 Folded_Diff_Op_Amp_Layout_0.VB4.t42 47.8416
R21969 Folded_Diff_Op_Amp_Layout_0.VB4.n27 Folded_Diff_Op_Amp_Layout_0.VB4.t59 47.8416
R21970 Folded_Diff_Op_Amp_Layout_0.VB4.n26 Folded_Diff_Op_Amp_Layout_0.VB4.t95 47.8416
R21971 Folded_Diff_Op_Amp_Layout_0.VB4.n42 Folded_Diff_Op_Amp_Layout_0.VB4.t39 47.8416
R21972 Folded_Diff_Op_Amp_Layout_0.VB4.n41 Folded_Diff_Op_Amp_Layout_0.VB4.t77 47.8416
R21973 Folded_Diff_Op_Amp_Layout_0.VB4.n40 Folded_Diff_Op_Amp_Layout_0.VB4.t93 47.8416
R21974 Folded_Diff_Op_Amp_Layout_0.VB4.n39 Folded_Diff_Op_Amp_Layout_0.VB4.t45 47.8416
R21975 Folded_Diff_Op_Amp_Layout_0.VB4.n43 Folded_Diff_Op_Amp_Layout_0.VB4.t81 47.8416
R21976 Folded_Diff_Op_Amp_Layout_0.VB4.n61 Folded_Diff_Op_Amp_Layout_0.VB4.t46 47.3393
R21977 Folded_Diff_Op_Amp_Layout_0.VB4.n51 Folded_Diff_Op_Amp_Layout_0.VB4.t97 47.0594
R21978 Folded_Diff_Op_Amp_Layout_0.VB4.n50 Folded_Diff_Op_Amp_Layout_0.VB4.t47 47.0594
R21979 Folded_Diff_Op_Amp_Layout_0.VB4.n49 Folded_Diff_Op_Amp_Layout_0.VB4.t49 47.0594
R21980 Folded_Diff_Op_Amp_Layout_0.VB4.n48 Folded_Diff_Op_Amp_Layout_0.VB4.t70 47.0594
R21981 Folded_Diff_Op_Amp_Layout_0.VB4.n47 Folded_Diff_Op_Amp_Layout_0.VB4.t72 47.0594
R21982 Folded_Diff_Op_Amp_Layout_0.VB4.n46 Folded_Diff_Op_Amp_Layout_0.VB4.t90 47.0594
R21983 Folded_Diff_Op_Amp_Layout_0.VB4.n44 Folded_Diff_Op_Amp_Layout_0.VB4.t88 47.0594
R21984 Folded_Diff_Op_Amp_Layout_0.VB4.n45 Folded_Diff_Op_Amp_Layout_0.VB4.t83 47.0594
R21985 Folded_Diff_Op_Amp_Layout_0.VB4.n13 Folded_Diff_Op_Amp_Layout_0.VB4.t79 46.538
R21986 Folded_Diff_Op_Amp_Layout_0.VB4.n21 Folded_Diff_Op_Amp_Layout_0.VB4.t94 46.538
R21987 Folded_Diff_Op_Amp_Layout_0.VB4.n20 Folded_Diff_Op_Amp_Layout_0.VB4.t64 46.538
R21988 Folded_Diff_Op_Amp_Layout_0.VB4.n19 Folded_Diff_Op_Amp_Layout_0.VB4.t76 46.538
R21989 Folded_Diff_Op_Amp_Layout_0.VB4.n18 Folded_Diff_Op_Amp_Layout_0.VB4.t48 46.538
R21990 Folded_Diff_Op_Amp_Layout_0.VB4.n32 Folded_Diff_Op_Amp_Layout_0.VB4.t63 46.538
R21991 Folded_Diff_Op_Amp_Layout_0.VB4.n36 Folded_Diff_Op_Amp_Layout_0.VB4.t80 46.538
R21992 Folded_Diff_Op_Amp_Layout_0.VB4.n35 Folded_Diff_Op_Amp_Layout_0.VB4.t52 46.538
R21993 Folded_Diff_Op_Amp_Layout_0.VB4.t92 Folded_Diff_Op_Amp_Layout_0.VB4.n11 45.8862
R21994 Folded_Diff_Op_Amp_Layout_0.VB4.n12 Folded_Diff_Op_Amp_Layout_0.VB4.t92 45.4951
R21995 Folded_Diff_Op_Amp_Layout_0.VB4.n16 Folded_Diff_Op_Amp_Layout_0.VB4.t35 45.4951
R21996 Folded_Diff_Op_Amp_Layout_0.VB4.n15 Folded_Diff_Op_Amp_Layout_0.VB4.t74 45.4951
R21997 Folded_Diff_Op_Amp_Layout_0.VB4.n14 Folded_Diff_Op_Amp_Layout_0.VB4.t86 45.4951
R21998 Folded_Diff_Op_Amp_Layout_0.VB4.n17 Folded_Diff_Op_Amp_Layout_0.VB4.t61 45.4951
R21999 Folded_Diff_Op_Amp_Layout_0.VB4.n31 Folded_Diff_Op_Amp_Layout_0.VB4.t73 45.4951
R22000 Folded_Diff_Op_Amp_Layout_0.VB4.n29 Folded_Diff_Op_Amp_Layout_0.VB4.t65 45.4951
R22001 Folded_Diff_Op_Amp_Layout_0.VB4.n30 Folded_Diff_Op_Amp_Layout_0.VB4.t98 45.4951
R22002 Folded_Diff_Op_Amp_Layout_0.VB4.n5 Folded_Diff_Op_Amp_Layout_0.VB4.t62 45.2344
R22003 Folded_Diff_Op_Amp_Layout_0.VB4.n11 Folded_Diff_Op_Amp_Layout_0.VB4.t58 45.2344
R22004 Folded_Diff_Op_Amp_Layout_0.VB4.n10 Folded_Diff_Op_Amp_Layout_0.VB4.t71 45.2344
R22005 Folded_Diff_Op_Amp_Layout_0.VB4.n9 Folded_Diff_Op_Amp_Layout_0.VB4.t38 45.2344
R22006 Folded_Diff_Op_Amp_Layout_0.VB4.n8 Folded_Diff_Op_Amp_Layout_0.VB4.t55 45.2344
R22007 Folded_Diff_Op_Amp_Layout_0.VB4.n7 Folded_Diff_Op_Amp_Layout_0.VB4.t91 45.2344
R22008 Folded_Diff_Op_Amp_Layout_0.VB4.n6 Folded_Diff_Op_Amp_Layout_0.VB4.t34 45.2344
R22009 Folded_Diff_Op_Amp_Layout_0.VB4.n4 Folded_Diff_Op_Amp_Layout_0.VB4.t100 45.2344
R22010 Folded_Diff_Op_Amp_Layout_0.VB4.n58 Folded_Diff_Op_Amp_Layout_0.VB4.t54 44.5826
R22011 Folded_Diff_Op_Amp_Layout_0.VB4.n57 Folded_Diff_Op_Amp_Layout_0.VB4.t57 44.5826
R22012 Folded_Diff_Op_Amp_Layout_0.VB4.n56 Folded_Diff_Op_Amp_Layout_0.VB4.t75 44.5826
R22013 Folded_Diff_Op_Amp_Layout_0.VB4.n55 Folded_Diff_Op_Amp_Layout_0.VB4.t78 44.5826
R22014 Folded_Diff_Op_Amp_Layout_0.VB4.n54 Folded_Diff_Op_Amp_Layout_0.VB4.t102 44.5826
R22015 Folded_Diff_Op_Amp_Layout_0.VB4.n53 Folded_Diff_Op_Amp_Layout_0.VB4.t96 44.5826
R22016 Folded_Diff_Op_Amp_Layout_0.VB4.n52 Folded_Diff_Op_Amp_Layout_0.VB4.t101 44.5826
R22017 Folded_Diff_Op_Amp_Layout_0.VB4.n59 Folded_Diff_Op_Amp_Layout_0.VB4.t32 44.5826
R22018 Folded_Diff_Op_Amp_Layout_0.VB4.n117 Folded_Diff_Op_Amp_Layout_0.VB4.t8 17.0773
R22019 Folded_Diff_Op_Amp_Layout_0.VB4.n115 Folded_Diff_Op_Amp_Layout_0.VB4.t30 17.0773
R22020 Folded_Diff_Op_Amp_Layout_0.VB4.n121 Folded_Diff_Op_Amp_Layout_0.VB4.t10 17.0773
R22021 Folded_Diff_Op_Amp_Layout_0.VB4.n105 Folded_Diff_Op_Amp_Layout_0.VB4.t16 17.0773
R22022 Folded_Diff_Op_Amp_Layout_0.VB4.n102 Folded_Diff_Op_Amp_Layout_0.VB4.t18 17.0773
R22023 Folded_Diff_Op_Amp_Layout_0.VB4.n100 Folded_Diff_Op_Amp_Layout_0.VB4.t28 17.0773
R22024 Folded_Diff_Op_Amp_Layout_0.VB4.n97 Folded_Diff_Op_Amp_Layout_0.VB4.t24 17.0773
R22025 Folded_Diff_Op_Amp_Layout_0.VB4.n95 Folded_Diff_Op_Amp_Layout_0.VB4.t26 17.0773
R22026 Folded_Diff_Op_Amp_Layout_0.VB4.n92 Folded_Diff_Op_Amp_Layout_0.VB4.t4 17.0773
R22027 Folded_Diff_Op_Amp_Layout_0.VB4.n90 Folded_Diff_Op_Amp_Layout_0.VB4.t6 17.0773
R22028 Folded_Diff_Op_Amp_Layout_0.VB4.n87 Folded_Diff_Op_Amp_Layout_0.VB4.t14 17.0773
R22029 Folded_Diff_Op_Amp_Layout_0.VB4.n85 Folded_Diff_Op_Amp_Layout_0.VB4.t22 17.0773
R22030 Folded_Diff_Op_Amp_Layout_0.VB4.n82 Folded_Diff_Op_Amp_Layout_0.VB4.t12 17.0773
R22031 Folded_Diff_Op_Amp_Layout_0.VB4.n80 Folded_Diff_Op_Amp_Layout_0.VB4.t20 17.0773
R22032 Folded_Diff_Op_Amp_Layout_0.VB4.n6 Folded_Diff_Op_Amp_Layout_0.VB4.n5 9.73383
R22033 Folded_Diff_Op_Amp_Layout_0.VB4.n5 Folded_Diff_Op_Amp_Layout_0.VB4.n4 9.73383
R22034 Folded_Diff_Op_Amp_Layout_0.VB4.n16 Folded_Diff_Op_Amp_Layout_0.VB4.n15 9.73383
R22035 Folded_Diff_Op_Amp_Layout_0.VB4.n15 Folded_Diff_Op_Amp_Layout_0.VB4.n14 9.73383
R22036 Folded_Diff_Op_Amp_Layout_0.VB4.n31 Folded_Diff_Op_Amp_Layout_0.VB4.n30 9.73383
R22037 Folded_Diff_Op_Amp_Layout_0.VB4.n30 Folded_Diff_Op_Amp_Layout_0.VB4.n29 9.73383
R22038 Folded_Diff_Op_Amp_Layout_0.VB4.n21 Folded_Diff_Op_Amp_Layout_0.VB4.n20 9.73383
R22039 Folded_Diff_Op_Amp_Layout_0.VB4.n20 Folded_Diff_Op_Amp_Layout_0.VB4.n19 9.73383
R22040 Folded_Diff_Op_Amp_Layout_0.VB4.n19 Folded_Diff_Op_Amp_Layout_0.VB4.n18 9.73383
R22041 Folded_Diff_Op_Amp_Layout_0.VB4.n36 Folded_Diff_Op_Amp_Layout_0.VB4.n35 9.73383
R22042 Folded_Diff_Op_Amp_Layout_0.VB4.n23 Folded_Diff_Op_Amp_Layout_0.VB4.n22 9.73383
R22043 Folded_Diff_Op_Amp_Layout_0.VB4.n25 Folded_Diff_Op_Amp_Layout_0.VB4.n24 9.73383
R22044 Folded_Diff_Op_Amp_Layout_0.VB4.n34 Folded_Diff_Op_Amp_Layout_0.VB4.n33 9.73383
R22045 Folded_Diff_Op_Amp_Layout_0.VB4.n38 Folded_Diff_Op_Amp_Layout_0.VB4.n37 9.73383
R22046 Folded_Diff_Op_Amp_Layout_0.VB4.n28 Folded_Diff_Op_Amp_Layout_0.VB4.n27 9.73383
R22047 Folded_Diff_Op_Amp_Layout_0.VB4.n27 Folded_Diff_Op_Amp_Layout_0.VB4.n26 9.73383
R22048 Folded_Diff_Op_Amp_Layout_0.VB4.n42 Folded_Diff_Op_Amp_Layout_0.VB4.n41 9.73383
R22049 Folded_Diff_Op_Amp_Layout_0.VB4.n41 Folded_Diff_Op_Amp_Layout_0.VB4.n40 9.73383
R22050 Folded_Diff_Op_Amp_Layout_0.VB4.n40 Folded_Diff_Op_Amp_Layout_0.VB4.n39 9.73383
R22051 Folded_Diff_Op_Amp_Layout_0.VB4.n51 Folded_Diff_Op_Amp_Layout_0.VB4.n50 9.73383
R22052 Folded_Diff_Op_Amp_Layout_0.VB4.n50 Folded_Diff_Op_Amp_Layout_0.VB4.n49 9.73383
R22053 Folded_Diff_Op_Amp_Layout_0.VB4.n49 Folded_Diff_Op_Amp_Layout_0.VB4.n48 9.73383
R22054 Folded_Diff_Op_Amp_Layout_0.VB4.n48 Folded_Diff_Op_Amp_Layout_0.VB4.n47 9.73383
R22055 Folded_Diff_Op_Amp_Layout_0.VB4.n47 Folded_Diff_Op_Amp_Layout_0.VB4.n46 9.73383
R22056 Folded_Diff_Op_Amp_Layout_0.VB4.n46 Folded_Diff_Op_Amp_Layout_0.VB4.n45 9.73383
R22057 Folded_Diff_Op_Amp_Layout_0.VB4.n45 Folded_Diff_Op_Amp_Layout_0.VB4.n44 9.73383
R22058 Folded_Diff_Op_Amp_Layout_0.VB4.n59 Folded_Diff_Op_Amp_Layout_0.VB4.n58 9.73383
R22059 Folded_Diff_Op_Amp_Layout_0.VB4.n58 Folded_Diff_Op_Amp_Layout_0.VB4.n57 9.73383
R22060 Folded_Diff_Op_Amp_Layout_0.VB4.n57 Folded_Diff_Op_Amp_Layout_0.VB4.n56 9.73383
R22061 Folded_Diff_Op_Amp_Layout_0.VB4.n56 Folded_Diff_Op_Amp_Layout_0.VB4.n55 9.73383
R22062 Folded_Diff_Op_Amp_Layout_0.VB4.n55 Folded_Diff_Op_Amp_Layout_0.VB4.n54 9.73383
R22063 Folded_Diff_Op_Amp_Layout_0.VB4.n54 Folded_Diff_Op_Amp_Layout_0.VB4.n53 9.73383
R22064 Folded_Diff_Op_Amp_Layout_0.VB4.n53 Folded_Diff_Op_Amp_Layout_0.VB4.n52 9.73383
R22065 Folded_Diff_Op_Amp_Layout_0.VB4.n7 Folded_Diff_Op_Amp_Layout_0.VB4.n6 9.28449
R22066 Folded_Diff_Op_Amp_Layout_0.VB4.n11 Folded_Diff_Op_Amp_Layout_0.VB4.n10 7.16614
R22067 Folded_Diff_Op_Amp_Layout_0.VB4.n10 Folded_Diff_Op_Amp_Layout_0.VB4.n9 7.16614
R22068 Folded_Diff_Op_Amp_Layout_0.VB4.n9 Folded_Diff_Op_Amp_Layout_0.VB4.n8 7.16614
R22069 Folded_Diff_Op_Amp_Layout_0.VB4.n8 Folded_Diff_Op_Amp_Layout_0.VB4.n7 7.16614
R22070 Folded_Diff_Op_Amp_Layout_0.VB4.n64 Folded_Diff_Op_Amp_Layout_0.VB4.n63 6.78515
R22071 Folded_Diff_Op_Amp_Layout_0.VB4.n111 Folded_Diff_Op_Amp_Layout_0.VB4.t3 5.69633
R22072 Folded_Diff_Op_Amp_Layout_0.VB4.n81 Folded_Diff_Op_Amp_Layout_0.VB4.n79 5.22676
R22073 Folded_Diff_Op_Amp_Layout_0.VB4.n0 Folded_Diff_Op_Amp_Layout_0.VB4.n122 4.5005
R22074 Folded_Diff_Op_Amp_Layout_0.VB4.n81 Folded_Diff_Op_Amp_Layout_0.VB4.n80 4.0005
R22075 Folded_Diff_Op_Amp_Layout_0.VB4.n83 Folded_Diff_Op_Amp_Layout_0.VB4.n82 4.0005
R22076 Folded_Diff_Op_Amp_Layout_0.VB4.n86 Folded_Diff_Op_Amp_Layout_0.VB4.n85 4.0005
R22077 Folded_Diff_Op_Amp_Layout_0.VB4.n88 Folded_Diff_Op_Amp_Layout_0.VB4.n87 4.0005
R22078 Folded_Diff_Op_Amp_Layout_0.VB4.n91 Folded_Diff_Op_Amp_Layout_0.VB4.n90 4.0005
R22079 Folded_Diff_Op_Amp_Layout_0.VB4.n93 Folded_Diff_Op_Amp_Layout_0.VB4.n92 4.0005
R22080 Folded_Diff_Op_Amp_Layout_0.VB4.n96 Folded_Diff_Op_Amp_Layout_0.VB4.n95 4.0005
R22081 Folded_Diff_Op_Amp_Layout_0.VB4.n98 Folded_Diff_Op_Amp_Layout_0.VB4.n97 4.0005
R22082 Folded_Diff_Op_Amp_Layout_0.VB4.n101 Folded_Diff_Op_Amp_Layout_0.VB4.n100 4.0005
R22083 Folded_Diff_Op_Amp_Layout_0.VB4.n103 Folded_Diff_Op_Amp_Layout_0.VB4.n102 4.0005
R22084 Folded_Diff_Op_Amp_Layout_0.VB4.n106 Folded_Diff_Op_Amp_Layout_0.VB4.n105 4.0005
R22085 Folded_Diff_Op_Amp_Layout_0.VB4.n0 Folded_Diff_Op_Amp_Layout_0.VB4.n121 4.0005
R22086 Folded_Diff_Op_Amp_Layout_0.VB4.n116 Folded_Diff_Op_Amp_Layout_0.VB4.n115 4.0005
R22087 Folded_Diff_Op_Amp_Layout_0.VB4.n118 Folded_Diff_Op_Amp_Layout_0.VB4.n117 4.0005
R22088 Folded_Diff_Op_Amp_Layout_0.VB4.n119 Folded_Diff_Op_Amp_Layout_0.VB4.n108 3.43224
R22089 Folded_Diff_Op_Amp_Layout_0.VB4.n104 Folded_Diff_Op_Amp_Layout_0.VB4.n70 3.43224
R22090 Folded_Diff_Op_Amp_Layout_0.VB4.n99 Folded_Diff_Op_Amp_Layout_0.VB4.n72 3.43224
R22091 Folded_Diff_Op_Amp_Layout_0.VB4.n94 Folded_Diff_Op_Amp_Layout_0.VB4.n74 3.43224
R22092 Folded_Diff_Op_Amp_Layout_0.VB4.n89 Folded_Diff_Op_Amp_Layout_0.VB4.n76 3.43224
R22093 Folded_Diff_Op_Amp_Layout_0.VB4.n84 Folded_Diff_Op_Amp_Layout_0.VB4.n78 3.43224
R22094 Folded_Diff_Op_Amp_Layout_0.VB4.n111 Folded_Diff_Op_Amp_Layout_0.VB4.n110 3.43224
R22095 Folded_Diff_Op_Amp_Layout_0.VB4.n114 Folded_Diff_Op_Amp_Layout_0.VB4.n113 3.1505
R22096 Folded_Diff_Op_Amp_Layout_0.VB4.n67 Folded_Diff_Op_Amp_Layout_0.VB4.n62 2.8805
R22097 Folded_Diff_Op_Amp_Layout_0.VB4.n61 Folded_Diff_Op_Amp_Layout_0.VB4.n60 2.82317
R22098 Folded_Diff_Op_Amp_Layout_0.VB4.n108 Folded_Diff_Op_Amp_Layout_0.VB4.t11 1.6385
R22099 Folded_Diff_Op_Amp_Layout_0.VB4.n108 Folded_Diff_Op_Amp_Layout_0.VB4.n107 1.6385
R22100 Folded_Diff_Op_Amp_Layout_0.VB4.n70 Folded_Diff_Op_Amp_Layout_0.VB4.t19 1.6385
R22101 Folded_Diff_Op_Amp_Layout_0.VB4.n70 Folded_Diff_Op_Amp_Layout_0.VB4.n69 1.6385
R22102 Folded_Diff_Op_Amp_Layout_0.VB4.n72 Folded_Diff_Op_Amp_Layout_0.VB4.t25 1.6385
R22103 Folded_Diff_Op_Amp_Layout_0.VB4.n72 Folded_Diff_Op_Amp_Layout_0.VB4.n71 1.6385
R22104 Folded_Diff_Op_Amp_Layout_0.VB4.n74 Folded_Diff_Op_Amp_Layout_0.VB4.t5 1.6385
R22105 Folded_Diff_Op_Amp_Layout_0.VB4.n74 Folded_Diff_Op_Amp_Layout_0.VB4.n73 1.6385
R22106 Folded_Diff_Op_Amp_Layout_0.VB4.n76 Folded_Diff_Op_Amp_Layout_0.VB4.t15 1.6385
R22107 Folded_Diff_Op_Amp_Layout_0.VB4.n76 Folded_Diff_Op_Amp_Layout_0.VB4.n75 1.6385
R22108 Folded_Diff_Op_Amp_Layout_0.VB4.n78 Folded_Diff_Op_Amp_Layout_0.VB4.t13 1.6385
R22109 Folded_Diff_Op_Amp_Layout_0.VB4.n78 Folded_Diff_Op_Amp_Layout_0.VB4.n77 1.6385
R22110 Folded_Diff_Op_Amp_Layout_0.VB4.n110 Folded_Diff_Op_Amp_Layout_0.VB4.t1 1.6385
R22111 Folded_Diff_Op_Amp_Layout_0.VB4.n110 Folded_Diff_Op_Amp_Layout_0.VB4.n109 1.6385
R22112 Folded_Diff_Op_Amp_Layout_0.VB4.n113 Folded_Diff_Op_Amp_Layout_0.VB4.t31 1.6385
R22113 Folded_Diff_Op_Amp_Layout_0.VB4.n113 Folded_Diff_Op_Amp_Layout_0.VB4.n112 1.6385
R22114 Folded_Diff_Op_Amp_Layout_0.VB4.n121 Folded_Diff_Op_Amp_Layout_0.VB4.n120 1.31856
R22115 Folded_Diff_Op_Amp_Layout_0.VB4.n62 Folded_Diff_Op_Amp_Layout_0.VB4.n61 1.18887
R22116 Folded_Diff_Op_Amp_Layout_0.VB4.n123 Folded_Diff_Op_Amp_Layout_0.VB4.n2 1.12594
R22117 Folded_Diff_Op_Amp_Layout_0.VB4.n123 Folded_Diff_Op_Amp_Layout_0.VB4.n3 6.85581
R22118 Folded_Diff_Op_Amp_Layout_0.VB4.n114 Folded_Diff_Op_Amp_Layout_0.VB4.n111 0.908326
R22119 Folded_Diff_Op_Amp_Layout_0.VB4.n1 Folded_Diff_Op_Amp_Layout_0.VB4.n67 4.23366
R22120 Folded_Diff_Op_Amp_Layout_0.VB4.n60 Folded_Diff_Op_Amp_Layout_0.VB4.n59 0.548
R22121 Folded_Diff_Op_Amp_Layout_0.VB4.n116 Folded_Diff_Op_Amp_Layout_0.VB4.n114 0.438761
R22122 Folded_Diff_Op_Amp_Layout_0.VB4.n83 Folded_Diff_Op_Amp_Layout_0.VB4.n81 0.313543
R22123 Folded_Diff_Op_Amp_Layout_0.VB4.n88 Folded_Diff_Op_Amp_Layout_0.VB4.n86 0.313543
R22124 Folded_Diff_Op_Amp_Layout_0.VB4.n93 Folded_Diff_Op_Amp_Layout_0.VB4.n91 0.313543
R22125 Folded_Diff_Op_Amp_Layout_0.VB4.n98 Folded_Diff_Op_Amp_Layout_0.VB4.n96 0.313543
R22126 Folded_Diff_Op_Amp_Layout_0.VB4.n103 Folded_Diff_Op_Amp_Layout_0.VB4.n101 0.313543
R22127 Folded_Diff_Op_Amp_Layout_0.VB4.n118 Folded_Diff_Op_Amp_Layout_0.VB4.n116 0.313543
R22128 Folded_Diff_Op_Amp_Layout_0.VB4.n3 Folded_Diff_Op_Amp_Layout_0.VB4.n106 0.202326
R22129 Folded_Diff_Op_Amp_Layout_0.VB4.n84 Folded_Diff_Op_Amp_Layout_0.VB4.n83 0.157022
R22130 Folded_Diff_Op_Amp_Layout_0.VB4.n86 Folded_Diff_Op_Amp_Layout_0.VB4.n84 0.157022
R22131 Folded_Diff_Op_Amp_Layout_0.VB4.n89 Folded_Diff_Op_Amp_Layout_0.VB4.n88 0.157022
R22132 Folded_Diff_Op_Amp_Layout_0.VB4.n91 Folded_Diff_Op_Amp_Layout_0.VB4.n89 0.157022
R22133 Folded_Diff_Op_Amp_Layout_0.VB4.n94 Folded_Diff_Op_Amp_Layout_0.VB4.n93 0.157022
R22134 Folded_Diff_Op_Amp_Layout_0.VB4.n96 Folded_Diff_Op_Amp_Layout_0.VB4.n94 0.157022
R22135 Folded_Diff_Op_Amp_Layout_0.VB4.n99 Folded_Diff_Op_Amp_Layout_0.VB4.n98 0.157022
R22136 Folded_Diff_Op_Amp_Layout_0.VB4.n101 Folded_Diff_Op_Amp_Layout_0.VB4.n99 0.157022
R22137 Folded_Diff_Op_Amp_Layout_0.VB4.n104 Folded_Diff_Op_Amp_Layout_0.VB4.n103 0.157022
R22138 Folded_Diff_Op_Amp_Layout_0.VB4.n106 Folded_Diff_Op_Amp_Layout_0.VB4.n104 0.157022
R22139 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB4.n123 0.112007
R22140 Folded_Diff_Op_Amp_Layout_0.VB4.n119 Folded_Diff_Op_Amp_Layout_0.VB4.n118 0.104587
R22141 Folded_Diff_Op_Amp_Layout_0.VB4.n66 Folded_Diff_Op_Amp_Layout_0.VB4.n65 0.0656316
R22142 Folded_Diff_Op_Amp_Layout_0.VB4.n0 Folded_Diff_Op_Amp_Layout_0.VB4.n119 0.034
R22143 Folded_Diff_Op_Amp_Layout_0.VB4.n67 Folded_Diff_Op_Amp_Layout_0.VB4.n66 0.0301053
R22144 Folded_Diff_Op_Amp_Layout_0.VB4.n65 Folded_Diff_Op_Amp_Layout_0.VB4.n64 0.0289211
R22145 Folded_Diff_Op_Amp_Layout_0.VB4.n3 Folded_Diff_Op_Amp_Layout_0.VB4.n0 0.025
R22146 Folded_Diff_Op_Amp_Layout_0.VB4.n2 Folded_Diff_Op_Amp_Layout_0.VB4.n1 0.0222197
R22147 Folded_Diff_Op_Amp_Layout_0.VB4.n2 Folded_Diff_Op_Amp_Layout_0.VB4.n68 0.0207053
R22148 Folded_Diff_Op_Amp_Layout_0.IND.n311 Folded_Diff_Op_Amp_Layout_0.IND.t68 4.62366
R22149 Folded_Diff_Op_Amp_Layout_0.IND.n337 Folded_Diff_Op_Amp_Layout_0.IND.n336 4.62366
R22150 Folded_Diff_Op_Amp_Layout_0.IND.n56 Folded_Diff_Op_Amp_Layout_0.IND.n55 4.37688
R22151 Folded_Diff_Op_Amp_Layout_0.IND.n110 Folded_Diff_Op_Amp_Layout_0.IND.n109 4.34373
R22152 Folded_Diff_Op_Amp_Layout_0.IND.n96 Folded_Diff_Op_Amp_Layout_0.IND.n95 4.34373
R22153 Folded_Diff_Op_Amp_Layout_0.IND.n62 Folded_Diff_Op_Amp_Layout_0.IND.n61 4.34007
R22154 Folded_Diff_Op_Amp_Layout_0.IND.n323 Folded_Diff_Op_Amp_Layout_0.IND.n322 4.13833
R22155 Folded_Diff_Op_Amp_Layout_0.IND.n306 Folded_Diff_Op_Amp_Layout_0.IND.n305 2.31142
R22156 Folded_Diff_Op_Amp_Layout_0.IND.n431 Folded_Diff_Op_Amp_Layout_0.IND.n430 1.66567
R22157 Folded_Diff_Op_Amp_Layout_0.IND.n455 Folded_Diff_Op_Amp_Layout_0.IND.t3 1.66567
R22158 Folded_Diff_Op_Amp_Layout_0.IND.n358 Folded_Diff_Op_Amp_Layout_0.IND.n356 1.6654
R22159 Folded_Diff_Op_Amp_Layout_0.IND.n383 Folded_Diff_Op_Amp_Layout_0.IND.t25 1.6654
R22160 Folded_Diff_Op_Amp_Layout_0.IND.n218 Folded_Diff_Op_Amp_Layout_0.IND.t2 1.66411
R22161 Folded_Diff_Op_Amp_Layout_0.IND.n168 Folded_Diff_Op_Amp_Layout_0.IND.n166 1.66411
R22162 Folded_Diff_Op_Amp_Layout_0.IND.n424 Folded_Diff_Op_Amp_Layout_0.IND.n421 1.49812
R22163 Folded_Diff_Op_Amp_Layout_0.IND.n465 Folded_Diff_Op_Amp_Layout_0.IND.n464 1.49801
R22164 Folded_Diff_Op_Amp_Layout_0.IND.n91 Folded_Diff_Op_Amp_Layout_0.IND.n90 1.49201
R22165 Folded_Diff_Op_Amp_Layout_0.IND.n80 Folded_Diff_Op_Amp_Layout_0.IND.t9 1.49201
R22166 Folded_Diff_Op_Amp_Layout_0.IND.n291 Folded_Diff_Op_Amp_Layout_0.IND.n290 1.49175
R22167 Folded_Diff_Op_Amp_Layout_0.IND.n280 Folded_Diff_Op_Amp_Layout_0.IND.t62 1.49175
R22168 Folded_Diff_Op_Amp_Layout_0.IND.n183 Folded_Diff_Op_Amp_Layout_0.IND.n182 1.49048
R22169 Folded_Diff_Op_Amp_Layout_0.IND.n172 Folded_Diff_Op_Amp_Layout_0.IND.t38 1.49048
R22170 Folded_Diff_Op_Amp_Layout_0.IND.n106 Folded_Diff_Op_Amp_Layout_0.IND.n105 1.47245
R22171 Folded_Diff_Op_Amp_Layout_0.IND.n101 Folded_Diff_Op_Amp_Layout_0.IND.n100 1.47245
R22172 Folded_Diff_Op_Amp_Layout_0.IND.n52 Folded_Diff_Op_Amp_Layout_0.IND.n51 1.46565
R22173 Folded_Diff_Op_Amp_Layout_0.IND.n2 Folded_Diff_Op_Amp_Layout_0.IND.n1 1.31982
R22174 Folded_Diff_Op_Amp_Layout_0.IND.n13 Folded_Diff_Op_Amp_Layout_0.IND.t71 1.31982
R22175 Folded_Diff_Op_Amp_Layout_0.IND.n142 Folded_Diff_Op_Amp_Layout_0.IND.t56 1.31982
R22176 Folded_Diff_Op_Amp_Layout_0.IND.n138 Folded_Diff_Op_Amp_Layout_0.IND.n137 1.31982
R22177 Folded_Diff_Op_Amp_Layout_0.IND.n252 Folded_Diff_Op_Amp_Layout_0.IND.n251 1.23423
R22178 Folded_Diff_Op_Amp_Layout_0.IND.n396 Folded_Diff_Op_Amp_Layout_0.IND.n395 1.19479
R22179 Folded_Diff_Op_Amp_Layout_0.IND.n287 Folded_Diff_Op_Amp_Layout_0.IND.n286 1.19462
R22180 Folded_Diff_Op_Amp_Layout_0.IND.n92 Folded_Diff_Op_Amp_Layout_0.IND.n91 1.19459
R22181 Folded_Diff_Op_Amp_Layout_0.IND.n81 Folded_Diff_Op_Amp_Layout_0.IND.n80 1.19459
R22182 Folded_Diff_Op_Amp_Layout_0.IND.n179 Folded_Diff_Op_Amp_Layout_0.IND.n178 1.19439
R22183 Folded_Diff_Op_Amp_Layout_0.IND.n9 Folded_Diff_Op_Amp_Layout_0.IND.n8 1.19395
R22184 Folded_Diff_Op_Amp_Layout_0.IND.n154 Folded_Diff_Op_Amp_Layout_0.IND.n153 1.19395
R22185 Folded_Diff_Op_Amp_Layout_0.IND.n143 Folded_Diff_Op_Amp_Layout_0.IND.n142 1.19393
R22186 Folded_Diff_Op_Amp_Layout_0.IND.n87 Folded_Diff_Op_Amp_Layout_0.IND.n86 1.17958
R22187 Folded_Diff_Op_Amp_Layout_0.IND.n269 Folded_Diff_Op_Amp_Layout_0.IND.n268 1.17929
R22188 Folded_Diff_Op_Amp_Layout_0.IND.n44 Folded_Diff_Op_Amp_Layout_0.IND.n43 1.17929
R22189 Folded_Diff_Op_Amp_Layout_0.IND.n292 Folded_Diff_Op_Amp_Layout_0.IND.n291 1.17924
R22190 Folded_Diff_Op_Amp_Layout_0.IND.n281 Folded_Diff_Op_Amp_Layout_0.IND.n280 1.17924
R22191 Folded_Diff_Op_Amp_Layout_0.IND.n184 Folded_Diff_Op_Amp_Layout_0.IND.n183 1.17917
R22192 Folded_Diff_Op_Amp_Layout_0.IND.n173 Folded_Diff_Op_Amp_Layout_0.IND.n172 1.17917
R22193 Folded_Diff_Op_Amp_Layout_0.IND.n402 Folded_Diff_Op_Amp_Layout_0.IND.n401 1.17907
R22194 Folded_Diff_Op_Amp_Layout_0.IND.n258 Folded_Diff_Op_Amp_Layout_0.IND.n257 1.17902
R22195 Folded_Diff_Op_Amp_Layout_0.IND.n33 Folded_Diff_Op_Amp_Layout_0.IND.n32 1.17902
R22196 Folded_Diff_Op_Amp_Layout_0.IND.n3 Folded_Diff_Op_Amp_Layout_0.IND.n2 1.1787
R22197 Folded_Diff_Op_Amp_Layout_0.IND.n14 Folded_Diff_Op_Amp_Layout_0.IND.n13 1.1787
R22198 Folded_Diff_Op_Amp_Layout_0.IND.n139 Folded_Diff_Op_Amp_Layout_0.IND.n138 1.1787
R22199 Folded_Diff_Op_Amp_Layout_0.IND.n467 Folded_Diff_Op_Amp_Layout_0.IND.n418 1.1775
R22200 Folded_Diff_Op_Amp_Layout_0.IND.n211 Folded_Diff_Op_Amp_Layout_0.IND.n210 1.16728
R22201 Folded_Diff_Op_Amp_Layout_0.IND.n235 Folded_Diff_Op_Amp_Layout_0.IND.n234 1.16675
R22202 Folded_Diff_Op_Amp_Layout_0.IND.n247 Folded_Diff_Op_Amp_Layout_0.IND.n246 1.16675
R22203 Folded_Diff_Op_Amp_Layout_0.IND.n374 Folded_Diff_Op_Amp_Layout_0.IND.n373 1.16675
R22204 Folded_Diff_Op_Amp_Layout_0.IND.n68 Folded_Diff_Op_Amp_Layout_0.IND.n67 1.16667
R22205 Folded_Diff_Op_Amp_Layout_0.IND.n219 Folded_Diff_Op_Amp_Layout_0.IND.n218 1.16641
R22206 Folded_Diff_Op_Amp_Layout_0.IND.n169 Folded_Diff_Op_Amp_Layout_0.IND.n168 1.16641
R22207 Folded_Diff_Op_Amp_Layout_0.IND.n445 Folded_Diff_Op_Amp_Layout_0.IND.n444 1.16617
R22208 Folded_Diff_Op_Amp_Layout_0.IND.n359 Folded_Diff_Op_Amp_Layout_0.IND.n358 1.16588
R22209 Folded_Diff_Op_Amp_Layout_0.IND.n384 Folded_Diff_Op_Amp_Layout_0.IND.n383 1.16588
R22210 Folded_Diff_Op_Amp_Layout_0.IND.n310 Folded_Diff_Op_Amp_Layout_0.IND.n309 1.1658
R22211 Folded_Diff_Op_Amp_Layout_0.IND.n329 Folded_Diff_Op_Amp_Layout_0.IND.n328 1.1658
R22212 Folded_Diff_Op_Amp_Layout_0.IND.n343 Folded_Diff_Op_Amp_Layout_0.IND.n342 1.1658
R22213 Folded_Diff_Op_Amp_Layout_0.IND.n432 Folded_Diff_Op_Amp_Layout_0.IND.n431 1.1656
R22214 Folded_Diff_Op_Amp_Layout_0.IND.n456 Folded_Diff_Op_Amp_Layout_0.IND.n455 1.1656
R22215 Folded_Diff_Op_Amp_Layout_0.IND.n278 Folded_Diff_Op_Amp_Layout_0.IND.n135 1.1515
R22216 Folded_Diff_Op_Amp_Layout_0.IND.n351 Folded_Diff_Op_Amp_Layout_0.IND.n78 1.1515
R22217 Folded_Diff_Op_Amp_Layout_0.IND.n415 Folded_Diff_Op_Amp_Layout_0.IND.n28 1.1515
R22218 Folded_Diff_Op_Amp_Layout_0.IND.n107 Folded_Diff_Op_Amp_Layout_0.IND.n106 1.14066
R22219 Folded_Diff_Op_Amp_Layout_0.IND.n102 Folded_Diff_Op_Amp_Layout_0.IND.n101 1.14066
R22220 Folded_Diff_Op_Amp_Layout_0.IND.n53 Folded_Diff_Op_Amp_Layout_0.IND.n52 1.14059
R22221 Folded_Diff_Op_Amp_Layout_0.IND.n15 Folded_Diff_Op_Amp_Layout_0.IND.n14 1.12717
R22222 Folded_Diff_Op_Amp_Layout_0.IND.n236 Folded_Diff_Op_Amp_Layout_0.IND.n235 1.1257
R22223 Folded_Diff_Op_Amp_Layout_0.IND.n375 Folded_Diff_Op_Amp_Layout_0.IND.n374 1.1257
R22224 Folded_Diff_Op_Amp_Layout_0.IND.n212 Folded_Diff_Op_Amp_Layout_0.IND.n211 1.1257
R22225 Folded_Diff_Op_Amp_Layout_0.IND.n112 Folded_Diff_Op_Amp_Layout_0.IND.n111 1.1255
R22226 Folded_Diff_Op_Amp_Layout_0.IND.n98 Folded_Diff_Op_Amp_Layout_0.IND.n97 1.1255
R22227 Folded_Diff_Op_Amp_Layout_0.IND.n313 Folded_Diff_Op_Amp_Layout_0.IND.n312 1.1255
R22228 Folded_Diff_Op_Amp_Layout_0.IND.n325 Folded_Diff_Op_Amp_Layout_0.IND.n324 1.1255
R22229 Folded_Diff_Op_Amp_Layout_0.IND.n339 Folded_Diff_Op_Amp_Layout_0.IND.n338 1.1255
R22230 Folded_Diff_Op_Amp_Layout_0.IND.n58 Folded_Diff_Op_Amp_Layout_0.IND.n57 1.1255
R22231 Folded_Diff_Op_Amp_Layout_0.IND.n64 Folded_Diff_Op_Amp_Layout_0.IND.n63 1.1255
R22232 Folded_Diff_Op_Amp_Layout_0.IND.n467 Folded_Diff_Op_Amp_Layout_0.IND.n466 1.1255
R22233 Folded_Diff_Op_Amp_Layout_0.IND.n414 Folded_Diff_Op_Amp_Layout_0.IND.n413 1.1255
R22234 Folded_Diff_Op_Amp_Layout_0.IND.n350 Folded_Diff_Op_Amp_Layout_0.IND.n349 1.1255
R22235 Folded_Diff_Op_Amp_Layout_0.IND.n277 Folded_Diff_Op_Amp_Layout_0.IND.n276 1.1255
R22236 Folded_Diff_Op_Amp_Layout_0.IND.n447 Folded_Diff_Op_Amp_Layout_0.IND.n446 1.10737
R22237 Folded_Diff_Op_Amp_Layout_0.IND.n249 Folded_Diff_Op_Amp_Layout_0.IND.n248 1.1073
R22238 Folded_Diff_Op_Amp_Layout_0.IND.n361 Folded_Diff_Op_Amp_Layout_0.IND.n360 1.1073
R22239 Folded_Diff_Op_Amp_Layout_0.IND.n386 Folded_Diff_Op_Amp_Layout_0.IND.n385 1.1073
R22240 Folded_Diff_Op_Amp_Layout_0.IND.n201 Folded_Diff_Op_Amp_Layout_0.IND.n170 1.1073
R22241 Folded_Diff_Op_Amp_Layout_0.IND.n221 Folded_Diff_Op_Amp_Layout_0.IND.n220 1.1073
R22242 Folded_Diff_Op_Amp_Layout_0.IND.n444 Folded_Diff_Op_Amp_Layout_0.IND.n443 1.09663
R22243 Folded_Diff_Op_Amp_Layout_0.IND.n234 Folded_Diff_Op_Amp_Layout_0.IND.n232 1.09644
R22244 Folded_Diff_Op_Amp_Layout_0.IND.n246 Folded_Diff_Op_Amp_Layout_0.IND.n245 1.09644
R22245 Folded_Diff_Op_Amp_Layout_0.IND.n373 Folded_Diff_Op_Amp_Layout_0.IND.n371 1.09644
R22246 Folded_Diff_Op_Amp_Layout_0.IND.n210 Folded_Diff_Op_Amp_Layout_0.IND.n208 1.09514
R22247 Folded_Diff_Op_Amp_Layout_0.IND.n67 Folded_Diff_Op_Amp_Layout_0.IND.n66 1.08656
R22248 Folded_Diff_Op_Amp_Layout_0.IND.n389 Folded_Diff_Op_Amp_Layout_0.IND.n388 1.05423
R22249 Folded_Diff_Op_Amp_Layout_0.IND.n390 Folded_Diff_Op_Amp_Layout_0.IND.n49 1.05265
R22250 Folded_Diff_Op_Amp_Layout_0.IND.n252 Folded_Diff_Op_Amp_Layout_0.IND.n224 1.0087
R22251 Folded_Diff_Op_Amp_Layout_0.IND.n309 Folded_Diff_Op_Amp_Layout_0.IND.n308 1.00677
R22252 Folded_Diff_Op_Amp_Layout_0.IND.n328 Folded_Diff_Op_Amp_Layout_0.IND.n327 1.00677
R22253 Folded_Diff_Op_Amp_Layout_0.IND.n342 Folded_Diff_Op_Amp_Layout_0.IND.n341 1.00677
R22254 Folded_Diff_Op_Amp_Layout_0.IND.n286 Folded_Diff_Op_Amp_Layout_0.IND.n285 0.922998
R22255 Folded_Diff_Op_Amp_Layout_0.IND.n86 Folded_Diff_Op_Amp_Layout_0.IND.n85 0.922926
R22256 Folded_Diff_Op_Amp_Layout_0.IND.n178 Folded_Diff_Op_Amp_Layout_0.IND.n177 0.92139
R22257 Folded_Diff_Op_Amp_Layout_0.IND.n401 Folded_Diff_Op_Amp_Layout_0.IND.n400 0.920264
R22258 Folded_Diff_Op_Amp_Layout_0.IND.n395 Folded_Diff_Op_Amp_Layout_0.IND.n394 0.920264
R22259 Folded_Diff_Op_Amp_Layout_0.IND.n434 Folded_Diff_Op_Amp_Layout_0.IND.n433 0.88565
R22260 Folded_Diff_Op_Amp_Layout_0.IND.n458 Folded_Diff_Op_Amp_Layout_0.IND.n457 0.88565
R22261 Folded_Diff_Op_Amp_Layout_0.IND.n268 Folded_Diff_Op_Amp_Layout_0.IND.n267 0.834379
R22262 Folded_Diff_Op_Amp_Layout_0.IND.n43 Folded_Diff_Op_Amp_Layout_0.IND.n42 0.834379
R22263 Folded_Diff_Op_Amp_Layout_0.IND.n257 Folded_Diff_Op_Amp_Layout_0.IND.n256 0.834365
R22264 Folded_Diff_Op_Amp_Layout_0.IND.n32 Folded_Diff_Op_Amp_Layout_0.IND.n31 0.834365
R22265 Folded_Diff_Op_Amp_Layout_0.IND.n8 Folded_Diff_Op_Amp_Layout_0.IND.n7 0.834193
R22266 Folded_Diff_Op_Amp_Layout_0.IND.n153 Folded_Diff_Op_Amp_Layout_0.IND.n152 0.834193
R22267 Folded_Diff_Op_Amp_Layout_0.IND.n122 Folded_Diff_Op_Amp_Layout_0.IND.n121 0.759312
R22268 Folded_Diff_Op_Amp_Layout_0.IND.n272 Folded_Diff_Op_Amp_Layout_0.IND.n271 0.727916
R22269 Folded_Diff_Op_Amp_Layout_0.IND.n331 Folded_Diff_Op_Amp_Layout_0.IND.n330 0.727916
R22270 Folded_Diff_Op_Amp_Layout_0.IND.n345 Folded_Diff_Op_Amp_Layout_0.IND.n344 0.727916
R22271 Folded_Diff_Op_Amp_Layout_0.IND.n47 Folded_Diff_Op_Amp_Layout_0.IND.n46 0.727916
R22272 Folded_Diff_Op_Amp_Layout_0.IND.n157 Folded_Diff_Op_Amp_Layout_0.IND.n156 0.727916
R22273 Folded_Diff_Op_Amp_Layout_0.IND.n119 Folded_Diff_Op_Amp_Layout_0.IND.n103 0.727104
R22274 Folded_Diff_Op_Amp_Layout_0.IND.n128 Folded_Diff_Op_Amp_Layout_0.IND.n88 0.727104
R22275 Folded_Diff_Op_Amp_Layout_0.IND.n299 Folded_Diff_Op_Amp_Layout_0.IND.n288 0.727104
R22276 Folded_Diff_Op_Amp_Layout_0.IND.n71 Folded_Diff_Op_Amp_Layout_0.IND.n69 0.727104
R22277 Folded_Diff_Op_Amp_Layout_0.IND.n25 Folded_Diff_Op_Amp_Layout_0.IND.n4 0.727104
R22278 Folded_Diff_Op_Amp_Layout_0.IND.n409 Folded_Diff_Op_Amp_Layout_0.IND.n397 0.727104
R22279 Folded_Diff_Op_Amp_Layout_0.IND.n162 Folded_Diff_Op_Amp_Layout_0.IND.n140 0.727104
R22280 Folded_Diff_Op_Amp_Layout_0.IND.n187 Folded_Diff_Op_Amp_Layout_0.IND.n185 0.727104
R22281 Folded_Diff_Op_Amp_Layout_0.IND.n196 Folded_Diff_Op_Amp_Layout_0.IND.n174 0.727104
R22282 Folded_Diff_Op_Amp_Layout_0.IND.n306 Folded_Diff_Op_Amp_Layout_0.IND.n278 0.656743
R22283 Folded_Diff_Op_Amp_Layout_0.IND.n78 Folded_Diff_Op_Amp_Layout_0.IND.n77 0.650188
R22284 Folded_Diff_Op_Amp_Layout_0.IND.n412 Folded_Diff_Op_Amp_Layout_0.IND.n411 0.650188
R22285 Folded_Diff_Op_Amp_Layout_0.IND.n192 Folded_Diff_Op_Amp_Layout_0.IND.n180 0.616779
R22286 Folded_Diff_Op_Amp_Layout_0.IND.n261 Folded_Diff_Op_Amp_Layout_0.IND.n259 0.616779
R22287 Folded_Diff_Op_Amp_Layout_0.IND.n115 Folded_Diff_Op_Amp_Layout_0.IND.n113 0.616779
R22288 Folded_Diff_Op_Amp_Layout_0.IND.n124 Folded_Diff_Op_Amp_Layout_0.IND.n93 0.616779
R22289 Folded_Diff_Op_Amp_Layout_0.IND.n133 Folded_Diff_Op_Amp_Layout_0.IND.n82 0.616779
R22290 Folded_Diff_Op_Amp_Layout_0.IND.n295 Folded_Diff_Op_Amp_Layout_0.IND.n293 0.616779
R22291 Folded_Diff_Op_Amp_Layout_0.IND.n304 Folded_Diff_Op_Amp_Layout_0.IND.n282 0.616779
R22292 Folded_Diff_Op_Amp_Layout_0.IND.n316 Folded_Diff_Op_Amp_Layout_0.IND.n314 0.616779
R22293 Folded_Diff_Op_Amp_Layout_0.IND.n76 Folded_Diff_Op_Amp_Layout_0.IND.n59 0.616779
R22294 Folded_Diff_Op_Amp_Layout_0.IND.n36 Folded_Diff_Op_Amp_Layout_0.IND.n34 0.616779
R22295 Folded_Diff_Op_Amp_Layout_0.IND.n20 Folded_Diff_Op_Amp_Layout_0.IND.n10 0.616779
R22296 Folded_Diff_Op_Amp_Layout_0.IND.n405 Folded_Diff_Op_Amp_Layout_0.IND.n403 0.616779
R22297 Folded_Diff_Op_Amp_Layout_0.IND.n146 Folded_Diff_Op_Amp_Layout_0.IND.n144 0.616779
R22298 Folded_Diff_Op_Amp_Layout_0.IND.n177 Folded_Diff_Op_Amp_Layout_0.IND.t41 0.56925
R22299 Folded_Diff_Op_Amp_Layout_0.IND.n177 Folded_Diff_Op_Amp_Layout_0.IND.n176 0.56925
R22300 Folded_Diff_Op_Amp_Layout_0.IND.n208 Folded_Diff_Op_Amp_Layout_0.IND.t13 0.56925
R22301 Folded_Diff_Op_Amp_Layout_0.IND.n208 Folded_Diff_Op_Amp_Layout_0.IND.n207 0.56925
R22302 Folded_Diff_Op_Amp_Layout_0.IND.n232 Folded_Diff_Op_Amp_Layout_0.IND.t20 0.56925
R22303 Folded_Diff_Op_Amp_Layout_0.IND.n232 Folded_Diff_Op_Amp_Layout_0.IND.n231 0.56925
R22304 Folded_Diff_Op_Amp_Layout_0.IND.n245 Folded_Diff_Op_Amp_Layout_0.IND.t28 0.56925
R22305 Folded_Diff_Op_Amp_Layout_0.IND.n245 Folded_Diff_Op_Amp_Layout_0.IND.n244 0.56925
R22306 Folded_Diff_Op_Amp_Layout_0.IND.n105 Folded_Diff_Op_Amp_Layout_0.IND.t0 0.56925
R22307 Folded_Diff_Op_Amp_Layout_0.IND.n105 Folded_Diff_Op_Amp_Layout_0.IND.n104 0.56925
R22308 Folded_Diff_Op_Amp_Layout_0.IND.n109 Folded_Diff_Op_Amp_Layout_0.IND.t42 0.56925
R22309 Folded_Diff_Op_Amp_Layout_0.IND.n109 Folded_Diff_Op_Amp_Layout_0.IND.n108 0.56925
R22310 Folded_Diff_Op_Amp_Layout_0.IND.n100 Folded_Diff_Op_Amp_Layout_0.IND.t1 0.56925
R22311 Folded_Diff_Op_Amp_Layout_0.IND.n100 Folded_Diff_Op_Amp_Layout_0.IND.n99 0.56925
R22312 Folded_Diff_Op_Amp_Layout_0.IND.n95 Folded_Diff_Op_Amp_Layout_0.IND.t44 0.56925
R22313 Folded_Diff_Op_Amp_Layout_0.IND.n95 Folded_Diff_Op_Amp_Layout_0.IND.n94 0.56925
R22314 Folded_Diff_Op_Amp_Layout_0.IND.n85 Folded_Diff_Op_Amp_Layout_0.IND.t17 0.56925
R22315 Folded_Diff_Op_Amp_Layout_0.IND.n85 Folded_Diff_Op_Amp_Layout_0.IND.n84 0.56925
R22316 Folded_Diff_Op_Amp_Layout_0.IND.n285 Folded_Diff_Op_Amp_Layout_0.IND.t34 0.56925
R22317 Folded_Diff_Op_Amp_Layout_0.IND.n285 Folded_Diff_Op_Amp_Layout_0.IND.n284 0.56925
R22318 Folded_Diff_Op_Amp_Layout_0.IND.n66 Folded_Diff_Op_Amp_Layout_0.IND.t18 0.56925
R22319 Folded_Diff_Op_Amp_Layout_0.IND.n66 Folded_Diff_Op_Amp_Layout_0.IND.n65 0.56925
R22320 Folded_Diff_Op_Amp_Layout_0.IND.n61 Folded_Diff_Op_Amp_Layout_0.IND.t22 0.56925
R22321 Folded_Diff_Op_Amp_Layout_0.IND.n61 Folded_Diff_Op_Amp_Layout_0.IND.n60 0.56925
R22322 Folded_Diff_Op_Amp_Layout_0.IND.n51 Folded_Diff_Op_Amp_Layout_0.IND.t32 0.56925
R22323 Folded_Diff_Op_Amp_Layout_0.IND.n51 Folded_Diff_Op_Amp_Layout_0.IND.n50 0.56925
R22324 Folded_Diff_Op_Amp_Layout_0.IND.n55 Folded_Diff_Op_Amp_Layout_0.IND.t7 0.56925
R22325 Folded_Diff_Op_Amp_Layout_0.IND.n55 Folded_Diff_Op_Amp_Layout_0.IND.n54 0.56925
R22326 Folded_Diff_Op_Amp_Layout_0.IND.n371 Folded_Diff_Op_Amp_Layout_0.IND.t12 0.56925
R22327 Folded_Diff_Op_Amp_Layout_0.IND.n371 Folded_Diff_Op_Amp_Layout_0.IND.n370 0.56925
R22328 Folded_Diff_Op_Amp_Layout_0.IND.n400 Folded_Diff_Op_Amp_Layout_0.IND.t31 0.56925
R22329 Folded_Diff_Op_Amp_Layout_0.IND.n400 Folded_Diff_Op_Amp_Layout_0.IND.n399 0.56925
R22330 Folded_Diff_Op_Amp_Layout_0.IND.n394 Folded_Diff_Op_Amp_Layout_0.IND.t15 0.56925
R22331 Folded_Diff_Op_Amp_Layout_0.IND.n394 Folded_Diff_Op_Amp_Layout_0.IND.n393 0.56925
R22332 Folded_Diff_Op_Amp_Layout_0.IND.n443 Folded_Diff_Op_Amp_Layout_0.IND.t24 0.56925
R22333 Folded_Diff_Op_Amp_Layout_0.IND.n443 Folded_Diff_Op_Amp_Layout_0.IND.n442 0.56925
R22334 Folded_Diff_Op_Amp_Layout_0.IND.n224 Folded_Diff_Op_Amp_Layout_0.IND.n223 0.516159
R22335 Folded_Diff_Op_Amp_Layout_0.IND.n199 Folded_Diff_Op_Amp_Layout_0.IND.n198 0.507313
R22336 Folded_Diff_Op_Amp_Layout_0.IND.n256 Folded_Diff_Op_Amp_Layout_0.IND.t47 0.485833
R22337 Folded_Diff_Op_Amp_Layout_0.IND.n256 Folded_Diff_Op_Amp_Layout_0.IND.n255 0.485833
R22338 Folded_Diff_Op_Amp_Layout_0.IND.n267 Folded_Diff_Op_Amp_Layout_0.IND.t51 0.485833
R22339 Folded_Diff_Op_Amp_Layout_0.IND.n267 Folded_Diff_Op_Amp_Layout_0.IND.n266 0.485833
R22340 Folded_Diff_Op_Amp_Layout_0.IND.n308 Folded_Diff_Op_Amp_Layout_0.IND.t59 0.485833
R22341 Folded_Diff_Op_Amp_Layout_0.IND.n327 Folded_Diff_Op_Amp_Layout_0.IND.t50 0.485833
R22342 Folded_Diff_Op_Amp_Layout_0.IND.n327 Folded_Diff_Op_Amp_Layout_0.IND.n326 0.485833
R22343 Folded_Diff_Op_Amp_Layout_0.IND.n322 Folded_Diff_Op_Amp_Layout_0.IND.t54 0.485833
R22344 Folded_Diff_Op_Amp_Layout_0.IND.n322 Folded_Diff_Op_Amp_Layout_0.IND.n321 0.485833
R22345 Folded_Diff_Op_Amp_Layout_0.IND.n341 Folded_Diff_Op_Amp_Layout_0.IND.n340 0.485833
R22346 Folded_Diff_Op_Amp_Layout_0.IND.n31 Folded_Diff_Op_Amp_Layout_0.IND.t55 0.485833
R22347 Folded_Diff_Op_Amp_Layout_0.IND.n31 Folded_Diff_Op_Amp_Layout_0.IND.n30 0.485833
R22348 Folded_Diff_Op_Amp_Layout_0.IND.n42 Folded_Diff_Op_Amp_Layout_0.IND.t49 0.485833
R22349 Folded_Diff_Op_Amp_Layout_0.IND.n42 Folded_Diff_Op_Amp_Layout_0.IND.n41 0.485833
R22350 Folded_Diff_Op_Amp_Layout_0.IND.n7 Folded_Diff_Op_Amp_Layout_0.IND.t64 0.485833
R22351 Folded_Diff_Op_Amp_Layout_0.IND.n7 Folded_Diff_Op_Amp_Layout_0.IND.n6 0.485833
R22352 Folded_Diff_Op_Amp_Layout_0.IND.n152 Folded_Diff_Op_Amp_Layout_0.IND.t67 0.485833
R22353 Folded_Diff_Op_Amp_Layout_0.IND.n152 Folded_Diff_Op_Amp_Layout_0.IND.n151 0.485833
R22354 Folded_Diff_Op_Amp_Layout_0.IND.n460 Folded_Diff_Op_Amp_Layout_0.IND.n459 0.475688
R22355 Folded_Diff_Op_Amp_Layout_0.IND.n117 Folded_Diff_Op_Amp_Layout_0.IND.n116 0.474125
R22356 Folded_Diff_Op_Amp_Layout_0.IND.n297 Folded_Diff_Op_Amp_Layout_0.IND.n296 0.474125
R22357 Folded_Diff_Op_Amp_Layout_0.IND.n302 Folded_Diff_Op_Amp_Layout_0.IND.n301 0.474125
R22358 Folded_Diff_Op_Amp_Layout_0.IND.n190 Folded_Diff_Op_Amp_Layout_0.IND.n189 0.474125
R22359 Folded_Diff_Op_Amp_Layout_0.IND.n194 Folded_Diff_Op_Amp_Layout_0.IND.n193 0.474125
R22360 Folded_Diff_Op_Amp_Layout_0.IND.n275 Folded_Diff_Op_Amp_Layout_0.IND.n274 0.470187
R22361 Folded_Diff_Op_Amp_Layout_0.IND.n135 Folded_Diff_Op_Amp_Layout_0.IND.n134 0.470187
R22362 Folded_Diff_Op_Amp_Layout_0.IND.n389 Folded_Diff_Op_Amp_Layout_0.IND.n351 0.419368
R22363 Folded_Diff_Op_Amp_Layout_0.IND.n253 Folded_Diff_Op_Amp_Layout_0.IND.n252 0.395709
R22364 Folded_Diff_Op_Amp_Layout_0.IND.n390 Folded_Diff_Op_Amp_Layout_0.IND.n389 0.390055
R22365 Folded_Diff_Op_Amp_Layout_0.IND.n416 Folded_Diff_Op_Amp_Layout_0.IND.n415 0.368687
R22366 Folded_Diff_Op_Amp_Layout_0.IND.n224 Folded_Diff_Op_Amp_Layout_0.IND.n164 0.336564
R22367 Folded_Diff_Op_Amp_Layout_0.IND.n264 Folded_Diff_Op_Amp_Layout_0.IND.n263 0.330687
R22368 Folded_Diff_Op_Amp_Layout_0.IND.n39 Folded_Diff_Op_Amp_Layout_0.IND.n38 0.330687
R22369 Folded_Diff_Op_Amp_Layout_0.IND.n238 Folded_Diff_Op_Amp_Layout_0.IND.n237 0.330125
R22370 Folded_Diff_Op_Amp_Layout_0.IND.n126 Folded_Diff_Op_Amp_Layout_0.IND.n125 0.330125
R22371 Folded_Diff_Op_Amp_Layout_0.IND.n131 Folded_Diff_Op_Amp_Layout_0.IND.n130 0.330125
R22372 Folded_Diff_Op_Amp_Layout_0.IND.n334 Folded_Diff_Op_Amp_Layout_0.IND.n333 0.330125
R22373 Folded_Diff_Op_Amp_Layout_0.IND.n319 Folded_Diff_Op_Amp_Layout_0.IND.n318 0.330125
R22374 Folded_Diff_Op_Amp_Layout_0.IND.n74 Folded_Diff_Op_Amp_Layout_0.IND.n73 0.330125
R22375 Folded_Diff_Op_Amp_Layout_0.IND.n364 Folded_Diff_Op_Amp_Layout_0.IND.n363 0.330125
R22376 Folded_Diff_Op_Amp_Layout_0.IND.n377 Folded_Diff_Op_Amp_Layout_0.IND.n376 0.330125
R22377 Folded_Diff_Op_Amp_Layout_0.IND.n23 Folded_Diff_Op_Amp_Layout_0.IND.n22 0.330125
R22378 Folded_Diff_Op_Amp_Layout_0.IND.n19 Folded_Diff_Op_Amp_Layout_0.IND.n18 0.330125
R22379 Folded_Diff_Op_Amp_Layout_0.IND.n407 Folded_Diff_Op_Amp_Layout_0.IND.n406 0.330125
R22380 Folded_Diff_Op_Amp_Layout_0.IND.n436 Folded_Diff_Op_Amp_Layout_0.IND.n435 0.330125
R22381 Folded_Diff_Op_Amp_Layout_0.IND.n450 Folded_Diff_Op_Amp_Layout_0.IND.n449 0.330125
R22382 Folded_Diff_Op_Amp_Layout_0.IND.n160 Folded_Diff_Op_Amp_Layout_0.IND.n159 0.330125
R22383 Folded_Diff_Op_Amp_Layout_0.IND.n149 Folded_Diff_Op_Amp_Layout_0.IND.n148 0.330125
R22384 Folded_Diff_Op_Amp_Layout_0.IND.n204 Folded_Diff_Op_Amp_Layout_0.IND.n203 0.330125
R22385 Folded_Diff_Op_Amp_Layout_0.IND.n214 Folded_Diff_Op_Amp_Layout_0.IND.n213 0.330125
R22386 Folded_Diff_Op_Amp_Layout_0.IND.n348 Folded_Diff_Op_Amp_Layout_0.IND.n347 0.29075
R22387 Folded_Diff_Op_Amp_Layout_0.IND.n28 Folded_Diff_Op_Amp_Layout_0.IND.n27 0.29075
R22388 Folded_Diff_Op_Amp_Layout_0.IND.n391 Folded_Diff_Op_Amp_Layout_0.IND.n390 0.262189
R22389 Folded_Diff_Op_Amp_Layout_0.IND.n307 Folded_Diff_Op_Amp_Layout_0.IND.n306 0.203334
R22390 Folded_Diff_Op_Amp_Layout_0.IND.n457 Folded_Diff_Op_Amp_Layout_0.IND.n453 0.0936537
R22391 Folded_Diff_Op_Amp_Layout_0.IND.n433 Folded_Diff_Op_Amp_Layout_0.IND.n428 0.0936537
R22392 Folded_Diff_Op_Amp_Layout_0.IND.n220 Folded_Diff_Op_Amp_Layout_0.IND.n216 0.108032
R22393 Folded_Diff_Op_Amp_Layout_0.IND.n170 Folded_Diff_Op_Amp_Layout_0.IND.n165 0.108032
R22394 Folded_Diff_Op_Amp_Layout_0.IND.n248 Folded_Diff_Op_Amp_Layout_0.IND.n242 0.0886741
R22395 Folded_Diff_Op_Amp_Layout_0.IND.n360 Folded_Diff_Op_Amp_Layout_0.IND.n355 0.0886741
R22396 Folded_Diff_Op_Amp_Layout_0.IND.n385 Folded_Diff_Op_Amp_Layout_0.IND.n381 0.0886741
R22397 Folded_Diff_Op_Amp_Layout_0.IND.n446 Folded_Diff_Op_Amp_Layout_0.IND.n440 0.0880141
R22398 Folded_Diff_Op_Amp_Layout_0.IND.n14 Folded_Diff_Op_Amp_Layout_0.IND.n12 0.0832399
R22399 Folded_Diff_Op_Amp_Layout_0.IND.n271 Folded_Diff_Op_Amp_Layout_0.IND.n270 0.0826464
R22400 Folded_Diff_Op_Amp_Layout_0.IND.n330 Folded_Diff_Op_Amp_Layout_0.IND.n329 0.0826464
R22401 Folded_Diff_Op_Amp_Layout_0.IND.n344 Folded_Diff_Op_Amp_Layout_0.IND.n343 0.0826464
R22402 Folded_Diff_Op_Amp_Layout_0.IND.n46 Folded_Diff_Op_Amp_Layout_0.IND.n45 0.0826464
R22403 Folded_Diff_Op_Amp_Layout_0.IND.n156 Folded_Diff_Op_Amp_Layout_0.IND.n155 0.0826464
R22404 Folded_Diff_Op_Amp_Layout_0.IND.n185 Folded_Diff_Op_Amp_Layout_0.IND.n181 0.0823987
R22405 Folded_Diff_Op_Amp_Layout_0.IND.n174 Folded_Diff_Op_Amp_Layout_0.IND.n171 0.0823987
R22406 Folded_Diff_Op_Amp_Layout_0.IND.n103 Folded_Diff_Op_Amp_Layout_0.IND.n98 0.0823987
R22407 Folded_Diff_Op_Amp_Layout_0.IND.n88 Folded_Diff_Op_Amp_Layout_0.IND.n83 0.0823987
R22408 Folded_Diff_Op_Amp_Layout_0.IND.n288 Folded_Diff_Op_Amp_Layout_0.IND.n283 0.0823987
R22409 Folded_Diff_Op_Amp_Layout_0.IND.n69 Folded_Diff_Op_Amp_Layout_0.IND.n64 0.0823987
R22410 Folded_Diff_Op_Amp_Layout_0.IND.n4 Folded_Diff_Op_Amp_Layout_0.IND.n0 0.0823987
R22411 Folded_Diff_Op_Amp_Layout_0.IND.n397 Folded_Diff_Op_Amp_Layout_0.IND.n392 0.0823987
R22412 Folded_Diff_Op_Amp_Layout_0.IND.n140 Folded_Diff_Op_Amp_Layout_0.IND.n136 0.0823987
R22413 Folded_Diff_Op_Amp_Layout_0.IND.n210 Folded_Diff_Op_Amp_Layout_0.IND.n209 0.0801656
R22414 Folded_Diff_Op_Amp_Layout_0.IND.n218 Folded_Diff_Op_Amp_Layout_0.IND.n217 0.0800575
R22415 Folded_Diff_Op_Amp_Layout_0.IND.n168 Folded_Diff_Op_Amp_Layout_0.IND.n167 0.0800575
R22416 Folded_Diff_Op_Amp_Layout_0.IND.n234 Folded_Diff_Op_Amp_Layout_0.IND.n233 0.0784141
R22417 Folded_Diff_Op_Amp_Layout_0.IND.n246 Folded_Diff_Op_Amp_Layout_0.IND.n243 0.0784141
R22418 Folded_Diff_Op_Amp_Layout_0.IND.n373 Folded_Diff_Op_Amp_Layout_0.IND.n372 0.0784141
R22419 Folded_Diff_Op_Amp_Layout_0.IND.n358 Folded_Diff_Op_Amp_Layout_0.IND.n357 0.0783056
R22420 Folded_Diff_Op_Amp_Layout_0.IND.n383 Folded_Diff_Op_Amp_Layout_0.IND.n382 0.0783056
R22421 Folded_Diff_Op_Amp_Layout_0.IND.n444 Folded_Diff_Op_Amp_Layout_0.IND.n441 0.0778549
R22422 Folded_Diff_Op_Amp_Layout_0.IND.n431 Folded_Diff_Op_Amp_Layout_0.IND.n429 0.0774429
R22423 Folded_Diff_Op_Amp_Layout_0.IND.n455 Folded_Diff_Op_Amp_Layout_0.IND.n454 0.0774429
R22424 Folded_Diff_Op_Amp_Layout_0.IND.n259 Folded_Diff_Op_Amp_Layout_0.IND.n254 0.0712285
R22425 Folded_Diff_Op_Amp_Layout_0.IND.n82 Folded_Diff_Op_Amp_Layout_0.IND.n79 0.0712285
R22426 Folded_Diff_Op_Amp_Layout_0.IND.n93 Folded_Diff_Op_Amp_Layout_0.IND.n89 0.0712285
R22427 Folded_Diff_Op_Amp_Layout_0.IND.n113 Folded_Diff_Op_Amp_Layout_0.IND.n107 0.0712285
R22428 Folded_Diff_Op_Amp_Layout_0.IND.n282 Folded_Diff_Op_Amp_Layout_0.IND.n279 0.0712285
R22429 Folded_Diff_Op_Amp_Layout_0.IND.n293 Folded_Diff_Op_Amp_Layout_0.IND.n289 0.0712285
R22430 Folded_Diff_Op_Amp_Layout_0.IND.n314 Folded_Diff_Op_Amp_Layout_0.IND.n310 0.0712285
R22431 Folded_Diff_Op_Amp_Layout_0.IND.n59 Folded_Diff_Op_Amp_Layout_0.IND.n53 0.0712285
R22432 Folded_Diff_Op_Amp_Layout_0.IND.n34 Folded_Diff_Op_Amp_Layout_0.IND.n29 0.0712285
R22433 Folded_Diff_Op_Amp_Layout_0.IND.n10 Folded_Diff_Op_Amp_Layout_0.IND.n5 0.0712285
R22434 Folded_Diff_Op_Amp_Layout_0.IND.n403 Folded_Diff_Op_Amp_Layout_0.IND.n398 0.0712285
R22435 Folded_Diff_Op_Amp_Layout_0.IND.n144 Folded_Diff_Op_Amp_Layout_0.IND.n141 0.0712285
R22436 Folded_Diff_Op_Amp_Layout_0.IND.n180 Folded_Diff_Op_Amp_Layout_0.IND.n175 0.0712285
R22437 Folded_Diff_Op_Amp_Layout_0.IND.n63 Folded_Diff_Op_Amp_Layout_0.IND.n62 0.0631087
R22438 Folded_Diff_Op_Amp_Layout_0.IND.n211 Folded_Diff_Op_Amp_Layout_0.IND.n206 0.129868
R22439 Folded_Diff_Op_Amp_Layout_0.IND.n235 Folded_Diff_Op_Amp_Layout_0.IND.n230 0.0623855
R22440 Folded_Diff_Op_Amp_Layout_0.IND.n374 Folded_Diff_Op_Amp_Layout_0.IND.n369 0.0623855
R22441 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.IND.n467 0.058875
R22442 Folded_Diff_Op_Amp_Layout_0.IND.n230 Folded_Diff_Op_Amp_Layout_0.IND.n229 0.0576486
R22443 Folded_Diff_Op_Amp_Layout_0.IND.n369 Folded_Diff_Op_Amp_Layout_0.IND.n368 0.0576486
R22444 Folded_Diff_Op_Amp_Layout_0.IND.n312 Folded_Diff_Op_Amp_Layout_0.IND.n311 0.0572391
R22445 Folded_Diff_Op_Amp_Layout_0.IND.n324 Folded_Diff_Op_Amp_Layout_0.IND.n323 0.0572391
R22446 Folded_Diff_Op_Amp_Layout_0.IND.n338 Folded_Diff_Op_Amp_Layout_0.IND.n337 0.0572391
R22447 Folded_Diff_Op_Amp_Layout_0.IND.n259 Folded_Diff_Op_Amp_Layout_0.IND.n258 0.0534597
R22448 Folded_Diff_Op_Amp_Layout_0.IND.n113 Folded_Diff_Op_Amp_Layout_0.IND.n112 0.0534597
R22449 Folded_Diff_Op_Amp_Layout_0.IND.n93 Folded_Diff_Op_Amp_Layout_0.IND.n92 0.0534597
R22450 Folded_Diff_Op_Amp_Layout_0.IND.n82 Folded_Diff_Op_Amp_Layout_0.IND.n81 0.0534597
R22451 Folded_Diff_Op_Amp_Layout_0.IND.n293 Folded_Diff_Op_Amp_Layout_0.IND.n292 0.0534597
R22452 Folded_Diff_Op_Amp_Layout_0.IND.n282 Folded_Diff_Op_Amp_Layout_0.IND.n281 0.0534597
R22453 Folded_Diff_Op_Amp_Layout_0.IND.n314 Folded_Diff_Op_Amp_Layout_0.IND.n313 0.0534597
R22454 Folded_Diff_Op_Amp_Layout_0.IND.n59 Folded_Diff_Op_Amp_Layout_0.IND.n58 0.0534597
R22455 Folded_Diff_Op_Amp_Layout_0.IND.n34 Folded_Diff_Op_Amp_Layout_0.IND.n33 0.0534597
R22456 Folded_Diff_Op_Amp_Layout_0.IND.n10 Folded_Diff_Op_Amp_Layout_0.IND.n9 0.0534597
R22457 Folded_Diff_Op_Amp_Layout_0.IND.n403 Folded_Diff_Op_Amp_Layout_0.IND.n402 0.0534597
R22458 Folded_Diff_Op_Amp_Layout_0.IND.n144 Folded_Diff_Op_Amp_Layout_0.IND.n143 0.0534597
R22459 Folded_Diff_Op_Amp_Layout_0.IND.n180 Folded_Diff_Op_Amp_Layout_0.IND.n179 0.0534597
R22460 Folded_Diff_Op_Amp_Layout_0.IND.n415 Folded_Diff_Op_Amp_Layout_0.IND.n414 0.0525
R22461 Folded_Diff_Op_Amp_Layout_0.IND.n414 Folded_Diff_Op_Amp_Layout_0.IND.n391 0.0525
R22462 Folded_Diff_Op_Amp_Layout_0.IND.n351 Folded_Diff_Op_Amp_Layout_0.IND.n350 0.0525
R22463 Folded_Diff_Op_Amp_Layout_0.IND.n350 Folded_Diff_Op_Amp_Layout_0.IND.n307 0.0525
R22464 Folded_Diff_Op_Amp_Layout_0.IND.n278 Folded_Diff_Op_Amp_Layout_0.IND.n277 0.0525
R22465 Folded_Diff_Op_Amp_Layout_0.IND.n277 Folded_Diff_Op_Amp_Layout_0.IND.n253 0.0525
R22466 Folded_Diff_Op_Amp_Layout_0.IND.n271 Folded_Diff_Op_Amp_Layout_0.IND.n269 0.0423164
R22467 Folded_Diff_Op_Amp_Layout_0.IND.n330 Folded_Diff_Op_Amp_Layout_0.IND.n325 0.0423164
R22468 Folded_Diff_Op_Amp_Layout_0.IND.n344 Folded_Diff_Op_Amp_Layout_0.IND.n339 0.0423164
R22469 Folded_Diff_Op_Amp_Layout_0.IND.n46 Folded_Diff_Op_Amp_Layout_0.IND.n44 0.0423164
R22470 Folded_Diff_Op_Amp_Layout_0.IND.n156 Folded_Diff_Op_Amp_Layout_0.IND.n154 0.0423164
R22471 Folded_Diff_Op_Amp_Layout_0.IND.n12 Folded_Diff_Op_Amp_Layout_0.IND.n11 0.0419676
R22472 Folded_Diff_Op_Amp_Layout_0.IND.n88 Folded_Diff_Op_Amp_Layout_0.IND.n87 0.0415773
R22473 Folded_Diff_Op_Amp_Layout_0.IND.n103 Folded_Diff_Op_Amp_Layout_0.IND.n102 0.0415773
R22474 Folded_Diff_Op_Amp_Layout_0.IND.n288 Folded_Diff_Op_Amp_Layout_0.IND.n287 0.0415773
R22475 Folded_Diff_Op_Amp_Layout_0.IND.n69 Folded_Diff_Op_Amp_Layout_0.IND.n68 0.0415773
R22476 Folded_Diff_Op_Amp_Layout_0.IND.n4 Folded_Diff_Op_Amp_Layout_0.IND.n3 0.0415773
R22477 Folded_Diff_Op_Amp_Layout_0.IND.n397 Folded_Diff_Op_Amp_Layout_0.IND.n396 0.0415773
R22478 Folded_Diff_Op_Amp_Layout_0.IND.n140 Folded_Diff_Op_Amp_Layout_0.IND.n139 0.0415773
R22479 Folded_Diff_Op_Amp_Layout_0.IND.n174 Folded_Diff_Op_Amp_Layout_0.IND.n173 0.0415773
R22480 Folded_Diff_Op_Amp_Layout_0.IND.n185 Folded_Diff_Op_Amp_Layout_0.IND.n184 0.0415773
R22481 Folded_Diff_Op_Amp_Layout_0.IND.n248 Folded_Diff_Op_Amp_Layout_0.IND.n247 0.032498
R22482 Folded_Diff_Op_Amp_Layout_0.IND.n385 Folded_Diff_Op_Amp_Layout_0.IND.n384 0.032498
R22483 Folded_Diff_Op_Amp_Layout_0.IND.n360 Folded_Diff_Op_Amp_Layout_0.IND.n359 0.032498
R22484 Folded_Diff_Op_Amp_Layout_0.IND.n220 Folded_Diff_Op_Amp_Layout_0.IND.n219 0.032498
R22485 Folded_Diff_Op_Amp_Layout_0.IND.n170 Folded_Diff_Op_Amp_Layout_0.IND.n169 0.032498
R22486 Folded_Diff_Op_Amp_Layout_0.IND.n446 Folded_Diff_Op_Amp_Layout_0.IND.n445 0.0319869
R22487 Folded_Diff_Op_Amp_Layout_0.IND.n57 Folded_Diff_Op_Amp_Layout_0.IND.n56 0.0269366
R22488 Folded_Diff_Op_Amp_Layout_0.IND.n276 Folded_Diff_Op_Amp_Layout_0.IND.n275 0.0265
R22489 Folded_Diff_Op_Amp_Layout_0.IND.n349 Folded_Diff_Op_Amp_Layout_0.IND.n348 0.0265
R22490 Folded_Diff_Op_Amp_Layout_0.IND.n413 Folded_Diff_Op_Amp_Layout_0.IND.n412 0.0265
R22491 Folded_Diff_Op_Amp_Layout_0.IND.n457 Folded_Diff_Op_Amp_Layout_0.IND.n456 0.0261793
R22492 Folded_Diff_Op_Amp_Layout_0.IND.n433 Folded_Diff_Op_Amp_Layout_0.IND.n432 0.0261793
R22493 Folded_Diff_Op_Amp_Layout_0.IND.n424 Folded_Diff_Op_Amp_Layout_0.IND.n423 0.0236139
R22494 Folded_Diff_Op_Amp_Layout_0.IND.n423 Folded_Diff_Op_Amp_Layout_0.IND.n422 0.0207053
R22495 Folded_Diff_Op_Amp_Layout_0.IND.n111 Folded_Diff_Op_Amp_Layout_0.IND.n110 0.0191828
R22496 Folded_Diff_Op_Amp_Layout_0.IND.n97 Folded_Diff_Op_Amp_Layout_0.IND.n96 0.0191828
R22497 Folded_Diff_Op_Amp_Layout_0.IND.n226 Folded_Diff_Op_Amp_Layout_0.IND.n225 0.0156875
R22498 Folded_Diff_Op_Amp_Layout_0.IND.n261 Folded_Diff_Op_Amp_Layout_0.IND.n260 0.0156875
R22499 Folded_Diff_Op_Amp_Layout_0.IND.n116 Folded_Diff_Op_Amp_Layout_0.IND.n115 0.0156875
R22500 Folded_Diff_Op_Amp_Layout_0.IND.n125 Folded_Diff_Op_Amp_Layout_0.IND.n124 0.0156875
R22501 Folded_Diff_Op_Amp_Layout_0.IND.n134 Folded_Diff_Op_Amp_Layout_0.IND.n133 0.0156875
R22502 Folded_Diff_Op_Amp_Layout_0.IND.n296 Folded_Diff_Op_Amp_Layout_0.IND.n295 0.0156875
R22503 Folded_Diff_Op_Amp_Layout_0.IND.n305 Folded_Diff_Op_Amp_Layout_0.IND.n304 0.0156875
R22504 Folded_Diff_Op_Amp_Layout_0.IND.n316 Folded_Diff_Op_Amp_Layout_0.IND.n315 0.0156875
R22505 Folded_Diff_Op_Amp_Layout_0.IND.n77 Folded_Diff_Op_Amp_Layout_0.IND.n76 0.0156875
R22506 Folded_Diff_Op_Amp_Layout_0.IND.n365 Folded_Diff_Op_Amp_Layout_0.IND.n364 0.0156875
R22507 Folded_Diff_Op_Amp_Layout_0.IND.n36 Folded_Diff_Op_Amp_Layout_0.IND.n35 0.0156875
R22508 Folded_Diff_Op_Amp_Layout_0.IND.n20 Folded_Diff_Op_Amp_Layout_0.IND.n19 0.0156875
R22509 Folded_Diff_Op_Amp_Layout_0.IND.n406 Folded_Diff_Op_Amp_Layout_0.IND.n405 0.0156875
R22510 Folded_Diff_Op_Amp_Layout_0.IND.n434 Folded_Diff_Op_Amp_Layout_0.IND.n425 0.0156875
R22511 Folded_Diff_Op_Amp_Layout_0.IND.n435 Folded_Diff_Op_Amp_Layout_0.IND.n434 0.0156875
R22512 Folded_Diff_Op_Amp_Layout_0.IND.n458 Folded_Diff_Op_Amp_Layout_0.IND.n450 0.0156875
R22513 Folded_Diff_Op_Amp_Layout_0.IND.n459 Folded_Diff_Op_Amp_Layout_0.IND.n458 0.0156875
R22514 Folded_Diff_Op_Amp_Layout_0.IND.n146 Folded_Diff_Op_Amp_Layout_0.IND.n145 0.0156875
R22515 Folded_Diff_Op_Amp_Layout_0.IND.n193 Folded_Diff_Op_Amp_Layout_0.IND.n192 0.0156875
R22516 Folded_Diff_Op_Amp_Layout_0.IND.n205 Folded_Diff_Op_Amp_Layout_0.IND.n204 0.0156875
R22517 Folded_Diff_Op_Amp_Layout_0.IND.n464 Folded_Diff_Op_Amp_Layout_0.IND.n463 0.014
R22518 Folded_Diff_Op_Amp_Layout_0.IND.n421 Folded_Diff_Op_Amp_Layout_0.IND.n419 0.014
R22519 Folded_Diff_Op_Amp_Layout_0.IND.n421 Folded_Diff_Op_Amp_Layout_0.IND.n420 0.014
R22520 Folded_Diff_Op_Amp_Layout_0.IND.n241 Folded_Diff_Op_Amp_Layout_0.IND.n240 0.0139513
R22521 Folded_Diff_Op_Amp_Layout_0.IND.n380 Folded_Diff_Op_Amp_Layout_0.IND.n379 0.0139513
R22522 Folded_Diff_Op_Amp_Layout_0.IND.n354 Folded_Diff_Op_Amp_Layout_0.IND.n353 0.0139513
R22523 Folded_Diff_Op_Amp_Layout_0.IND.n463 Folded_Diff_Op_Amp_Layout_0.IND.n462 0.0134654
R22524 Folded_Diff_Op_Amp_Layout_0.IND.n439 Folded_Diff_Op_Amp_Layout_0.IND.n438 0.0133659
R22525 Folded_Diff_Op_Amp_Layout_0.IND.n237 Folded_Diff_Op_Amp_Layout_0.IND.n236 0.0123533
R22526 Folded_Diff_Op_Amp_Layout_0.IND.n376 Folded_Diff_Op_Amp_Layout_0.IND.n375 0.0123533
R22527 Folded_Diff_Op_Amp_Layout_0.IND.n213 Folded_Diff_Op_Amp_Layout_0.IND.n212 0.0123533
R22528 Folded_Diff_Op_Amp_Layout_0.IND.n251 Folded_Diff_Op_Amp_Layout_0.IND.n250 0.0111023
R22529 Folded_Diff_Op_Amp_Layout_0.IND.n363 Folded_Diff_Op_Amp_Layout_0.IND.n362 0.0111023
R22530 Folded_Diff_Op_Amp_Layout_0.IND.n388 Folded_Diff_Op_Amp_Layout_0.IND.n387 0.0111023
R22531 Folded_Diff_Op_Amp_Layout_0.IND.n449 Folded_Diff_Op_Amp_Layout_0.IND.n448 0.0111023
R22532 Folded_Diff_Op_Amp_Layout_0.IND.n223 Folded_Diff_Op_Amp_Layout_0.IND.n222 0.0111023
R22533 Folded_Diff_Op_Amp_Layout_0.IND.n203 Folded_Diff_Op_Amp_Layout_0.IND.n202 0.0111023
R22534 Folded_Diff_Op_Amp_Layout_0.IND.n461 Folded_Diff_Op_Amp_Layout_0.IND.n460 0.00998204
R22535 Folded_Diff_Op_Amp_Layout_0.IND.n188 Folded_Diff_Op_Amp_Layout_0.IND.n187 0.00860784
R22536 Folded_Diff_Op_Amp_Layout_0.IND.n192 Folded_Diff_Op_Amp_Layout_0.IND.n191 0.00860784
R22537 Folded_Diff_Op_Amp_Layout_0.IND.n197 Folded_Diff_Op_Amp_Layout_0.IND.n196 0.00860784
R22538 Folded_Diff_Op_Amp_Layout_0.IND.n201 Folded_Diff_Op_Amp_Layout_0.IND.n200 0.00860784
R22539 Folded_Diff_Op_Amp_Layout_0.IND.n221 Folded_Diff_Op_Amp_Layout_0.IND.n215 0.00860784
R22540 Folded_Diff_Op_Amp_Layout_0.IND.n249 Folded_Diff_Op_Amp_Layout_0.IND.n239 0.00860784
R22541 Folded_Diff_Op_Amp_Layout_0.IND.n262 Folded_Diff_Op_Amp_Layout_0.IND.n261 0.00860784
R22542 Folded_Diff_Op_Amp_Layout_0.IND.n115 Folded_Diff_Op_Amp_Layout_0.IND.n114 0.00860784
R22543 Folded_Diff_Op_Amp_Layout_0.IND.n120 Folded_Diff_Op_Amp_Layout_0.IND.n119 0.00860784
R22544 Folded_Diff_Op_Amp_Layout_0.IND.n124 Folded_Diff_Op_Amp_Layout_0.IND.n123 0.00860784
R22545 Folded_Diff_Op_Amp_Layout_0.IND.n129 Folded_Diff_Op_Amp_Layout_0.IND.n128 0.00860784
R22546 Folded_Diff_Op_Amp_Layout_0.IND.n133 Folded_Diff_Op_Amp_Layout_0.IND.n132 0.00860784
R22547 Folded_Diff_Op_Amp_Layout_0.IND.n295 Folded_Diff_Op_Amp_Layout_0.IND.n294 0.00860784
R22548 Folded_Diff_Op_Amp_Layout_0.IND.n300 Folded_Diff_Op_Amp_Layout_0.IND.n299 0.00860784
R22549 Folded_Diff_Op_Amp_Layout_0.IND.n304 Folded_Diff_Op_Amp_Layout_0.IND.n303 0.00860784
R22550 Folded_Diff_Op_Amp_Layout_0.IND.n317 Folded_Diff_Op_Amp_Layout_0.IND.n316 0.00860784
R22551 Folded_Diff_Op_Amp_Layout_0.IND.n72 Folded_Diff_Op_Amp_Layout_0.IND.n71 0.00860784
R22552 Folded_Diff_Op_Amp_Layout_0.IND.n76 Folded_Diff_Op_Amp_Layout_0.IND.n75 0.00860784
R22553 Folded_Diff_Op_Amp_Layout_0.IND.n361 Folded_Diff_Op_Amp_Layout_0.IND.n352 0.00860784
R22554 Folded_Diff_Op_Amp_Layout_0.IND.n386 Folded_Diff_Op_Amp_Layout_0.IND.n378 0.00860784
R22555 Folded_Diff_Op_Amp_Layout_0.IND.n37 Folded_Diff_Op_Amp_Layout_0.IND.n36 0.00860784
R22556 Folded_Diff_Op_Amp_Layout_0.IND.n25 Folded_Diff_Op_Amp_Layout_0.IND.n24 0.00860784
R22557 Folded_Diff_Op_Amp_Layout_0.IND.n21 Folded_Diff_Op_Amp_Layout_0.IND.n20 0.00860784
R22558 Folded_Diff_Op_Amp_Layout_0.IND.n17 Folded_Diff_Op_Amp_Layout_0.IND.n16 0.00860784
R22559 Folded_Diff_Op_Amp_Layout_0.IND.n405 Folded_Diff_Op_Amp_Layout_0.IND.n404 0.00860784
R22560 Folded_Diff_Op_Amp_Layout_0.IND.n410 Folded_Diff_Op_Amp_Layout_0.IND.n409 0.00860784
R22561 Folded_Diff_Op_Amp_Layout_0.IND.n447 Folded_Diff_Op_Amp_Layout_0.IND.n437 0.00860784
R22562 Folded_Diff_Op_Amp_Layout_0.IND.n147 Folded_Diff_Op_Amp_Layout_0.IND.n146 0.00860784
R22563 Folded_Diff_Op_Amp_Layout_0.IND.n162 Folded_Diff_Op_Amp_Layout_0.IND.n161 0.00860784
R22564 Folded_Diff_Op_Amp_Layout_0.IND.n273 Folded_Diff_Op_Amp_Layout_0.IND.n272 0.00858096
R22565 Folded_Diff_Op_Amp_Layout_0.IND.n265 Folded_Diff_Op_Amp_Layout_0.IND.n264 0.00858096
R22566 Folded_Diff_Op_Amp_Layout_0.IND.n274 Folded_Diff_Op_Amp_Layout_0.IND.n273 0.00858096
R22567 Folded_Diff_Op_Amp_Layout_0.IND.n272 Folded_Diff_Op_Amp_Layout_0.IND.n265 0.00858096
R22568 Folded_Diff_Op_Amp_Layout_0.IND.n118 Folded_Diff_Op_Amp_Layout_0.IND.n117 0.00858096
R22569 Folded_Diff_Op_Amp_Layout_0.IND.n127 Folded_Diff_Op_Amp_Layout_0.IND.n126 0.00858096
R22570 Folded_Diff_Op_Amp_Layout_0.IND.n128 Folded_Diff_Op_Amp_Layout_0.IND.n127 0.00858096
R22571 Folded_Diff_Op_Amp_Layout_0.IND.n119 Folded_Diff_Op_Amp_Layout_0.IND.n118 0.00858096
R22572 Folded_Diff_Op_Amp_Layout_0.IND.n298 Folded_Diff_Op_Amp_Layout_0.IND.n297 0.00858096
R22573 Folded_Diff_Op_Amp_Layout_0.IND.n299 Folded_Diff_Op_Amp_Layout_0.IND.n298 0.00858096
R22574 Folded_Diff_Op_Amp_Layout_0.IND.n346 Folded_Diff_Op_Amp_Layout_0.IND.n345 0.00858096
R22575 Folded_Diff_Op_Amp_Layout_0.IND.n335 Folded_Diff_Op_Amp_Layout_0.IND.n334 0.00858096
R22576 Folded_Diff_Op_Amp_Layout_0.IND.n332 Folded_Diff_Op_Amp_Layout_0.IND.n331 0.00858096
R22577 Folded_Diff_Op_Amp_Layout_0.IND.n320 Folded_Diff_Op_Amp_Layout_0.IND.n319 0.00858096
R22578 Folded_Diff_Op_Amp_Layout_0.IND.n347 Folded_Diff_Op_Amp_Layout_0.IND.n346 0.00858096
R22579 Folded_Diff_Op_Amp_Layout_0.IND.n345 Folded_Diff_Op_Amp_Layout_0.IND.n335 0.00858096
R22580 Folded_Diff_Op_Amp_Layout_0.IND.n333 Folded_Diff_Op_Amp_Layout_0.IND.n332 0.00858096
R22581 Folded_Diff_Op_Amp_Layout_0.IND.n331 Folded_Diff_Op_Amp_Layout_0.IND.n320 0.00858096
R22582 Folded_Diff_Op_Amp_Layout_0.IND.n71 Folded_Diff_Op_Amp_Layout_0.IND.n70 0.00858096
R22583 Folded_Diff_Op_Amp_Layout_0.IND.n48 Folded_Diff_Op_Amp_Layout_0.IND.n47 0.00858096
R22584 Folded_Diff_Op_Amp_Layout_0.IND.n40 Folded_Diff_Op_Amp_Layout_0.IND.n39 0.00858096
R22585 Folded_Diff_Op_Amp_Layout_0.IND.n49 Folded_Diff_Op_Amp_Layout_0.IND.n48 0.00858096
R22586 Folded_Diff_Op_Amp_Layout_0.IND.n47 Folded_Diff_Op_Amp_Layout_0.IND.n40 0.00858096
R22587 Folded_Diff_Op_Amp_Layout_0.IND.n27 Folded_Diff_Op_Amp_Layout_0.IND.n26 0.00858096
R22588 Folded_Diff_Op_Amp_Layout_0.IND.n26 Folded_Diff_Op_Amp_Layout_0.IND.n25 0.00858096
R22589 Folded_Diff_Op_Amp_Layout_0.IND.n408 Folded_Diff_Op_Amp_Layout_0.IND.n407 0.00858096
R22590 Folded_Diff_Op_Amp_Layout_0.IND.n409 Folded_Diff_Op_Amp_Layout_0.IND.n408 0.00858096
R22591 Folded_Diff_Op_Amp_Layout_0.IND.n164 Folded_Diff_Op_Amp_Layout_0.IND.n163 0.00858096
R22592 Folded_Diff_Op_Amp_Layout_0.IND.n158 Folded_Diff_Op_Amp_Layout_0.IND.n157 0.00858096
R22593 Folded_Diff_Op_Amp_Layout_0.IND.n150 Folded_Diff_Op_Amp_Layout_0.IND.n149 0.00858096
R22594 Folded_Diff_Op_Amp_Layout_0.IND.n163 Folded_Diff_Op_Amp_Layout_0.IND.n162 0.00858096
R22595 Folded_Diff_Op_Amp_Layout_0.IND.n159 Folded_Diff_Op_Amp_Layout_0.IND.n158 0.00858096
R22596 Folded_Diff_Op_Amp_Layout_0.IND.n157 Folded_Diff_Op_Amp_Layout_0.IND.n150 0.00858096
R22597 Folded_Diff_Op_Amp_Layout_0.IND.n195 Folded_Diff_Op_Amp_Layout_0.IND.n194 0.00858096
R22598 Folded_Diff_Op_Amp_Layout_0.IND.n196 Folded_Diff_Op_Amp_Layout_0.IND.n195 0.00858096
R22599 Folded_Diff_Op_Amp_Layout_0.IND.n187 Folded_Diff_Op_Amp_Layout_0.IND.n186 0.00858096
R22600 Folded_Diff_Op_Amp_Layout_0.IND.n239 Folded_Diff_Op_Amp_Layout_0.IND.n238 0.00855417
R22601 Folded_Diff_Op_Amp_Layout_0.IND.n263 Folded_Diff_Op_Amp_Layout_0.IND.n262 0.00855417
R22602 Folded_Diff_Op_Amp_Layout_0.IND.n121 Folded_Diff_Op_Amp_Layout_0.IND.n120 0.00855417
R22603 Folded_Diff_Op_Amp_Layout_0.IND.n123 Folded_Diff_Op_Amp_Layout_0.IND.n122 0.00855417
R22604 Folded_Diff_Op_Amp_Layout_0.IND.n130 Folded_Diff_Op_Amp_Layout_0.IND.n129 0.00855417
R22605 Folded_Diff_Op_Amp_Layout_0.IND.n132 Folded_Diff_Op_Amp_Layout_0.IND.n131 0.00855417
R22606 Folded_Diff_Op_Amp_Layout_0.IND.n301 Folded_Diff_Op_Amp_Layout_0.IND.n300 0.00855417
R22607 Folded_Diff_Op_Amp_Layout_0.IND.n303 Folded_Diff_Op_Amp_Layout_0.IND.n302 0.00855417
R22608 Folded_Diff_Op_Amp_Layout_0.IND.n318 Folded_Diff_Op_Amp_Layout_0.IND.n317 0.00855417
R22609 Folded_Diff_Op_Amp_Layout_0.IND.n73 Folded_Diff_Op_Amp_Layout_0.IND.n72 0.00855417
R22610 Folded_Diff_Op_Amp_Layout_0.IND.n75 Folded_Diff_Op_Amp_Layout_0.IND.n74 0.00855417
R22611 Folded_Diff_Op_Amp_Layout_0.IND.n378 Folded_Diff_Op_Amp_Layout_0.IND.n377 0.00855417
R22612 Folded_Diff_Op_Amp_Layout_0.IND.n38 Folded_Diff_Op_Amp_Layout_0.IND.n37 0.00855417
R22613 Folded_Diff_Op_Amp_Layout_0.IND.n24 Folded_Diff_Op_Amp_Layout_0.IND.n23 0.00855417
R22614 Folded_Diff_Op_Amp_Layout_0.IND.n22 Folded_Diff_Op_Amp_Layout_0.IND.n21 0.00855417
R22615 Folded_Diff_Op_Amp_Layout_0.IND.n18 Folded_Diff_Op_Amp_Layout_0.IND.n17 0.00855417
R22616 Folded_Diff_Op_Amp_Layout_0.IND.n411 Folded_Diff_Op_Amp_Layout_0.IND.n410 0.00855417
R22617 Folded_Diff_Op_Amp_Layout_0.IND.n437 Folded_Diff_Op_Amp_Layout_0.IND.n436 0.00855417
R22618 Folded_Diff_Op_Amp_Layout_0.IND.n161 Folded_Diff_Op_Amp_Layout_0.IND.n160 0.00855417
R22619 Folded_Diff_Op_Amp_Layout_0.IND.n148 Folded_Diff_Op_Amp_Layout_0.IND.n147 0.00855417
R22620 Folded_Diff_Op_Amp_Layout_0.IND.n189 Folded_Diff_Op_Amp_Layout_0.IND.n188 0.00855417
R22621 Folded_Diff_Op_Amp_Layout_0.IND.n191 Folded_Diff_Op_Amp_Layout_0.IND.n190 0.00855417
R22622 Folded_Diff_Op_Amp_Layout_0.IND.n198 Folded_Diff_Op_Amp_Layout_0.IND.n197 0.00855417
R22623 Folded_Diff_Op_Amp_Layout_0.IND.n200 Folded_Diff_Op_Amp_Layout_0.IND.n199 0.00855417
R22624 Folded_Diff_Op_Amp_Layout_0.IND.n215 Folded_Diff_Op_Amp_Layout_0.IND.n214 0.00855417
R22625 Folded_Diff_Op_Amp_Layout_0.IND.n417 Folded_Diff_Op_Amp_Layout_0.IND.n416 0.00773989
R22626 Folded_Diff_Op_Amp_Layout_0.IND.n418 Folded_Diff_Op_Amp_Layout_0.IND.n417 0.00773989
R22627 Folded_Diff_Op_Amp_Layout_0.IND.n428 Folded_Diff_Op_Amp_Layout_0.IND.n427 0.00642105
R22628 Folded_Diff_Op_Amp_Layout_0.IND.n440 Folded_Diff_Op_Amp_Layout_0.IND.n439 0.00642105
R22629 Folded_Diff_Op_Amp_Layout_0.IND.n453 Folded_Diff_Op_Amp_Layout_0.IND.n452 0.00642105
R22630 Folded_Diff_Op_Amp_Layout_0.IND.n250 Folded_Diff_Op_Amp_Layout_0.IND.n249 0.00605114
R22631 Folded_Diff_Op_Amp_Layout_0.IND.n387 Folded_Diff_Op_Amp_Layout_0.IND.n386 0.00605114
R22632 Folded_Diff_Op_Amp_Layout_0.IND.n362 Folded_Diff_Op_Amp_Layout_0.IND.n361 0.00605114
R22633 Folded_Diff_Op_Amp_Layout_0.IND.n448 Folded_Diff_Op_Amp_Layout_0.IND.n447 0.00605114
R22634 Folded_Diff_Op_Amp_Layout_0.IND.n202 Folded_Diff_Op_Amp_Layout_0.IND.n201 0.00605114
R22635 Folded_Diff_Op_Amp_Layout_0.IND.n222 Folded_Diff_Op_Amp_Layout_0.IND.n221 0.00605114
R22636 Folded_Diff_Op_Amp_Layout_0.IND.n466 Folded_Diff_Op_Amp_Layout_0.IND.n424 0.00582347
R22637 Folded_Diff_Op_Amp_Layout_0.IND.n228 Folded_Diff_Op_Amp_Layout_0.IND.n227 0.00570918
R22638 Folded_Diff_Op_Amp_Layout_0.IND.n367 Folded_Diff_Op_Amp_Layout_0.IND.n366 0.00570918
R22639 Folded_Diff_Op_Amp_Layout_0.IND.n452 Folded_Diff_Op_Amp_Layout_0.IND.n451 0.00551512
R22640 Folded_Diff_Op_Amp_Layout_0.IND.n427 Folded_Diff_Op_Amp_Layout_0.IND.n426 0.00551512
R22641 Folded_Diff_Op_Amp_Layout_0.IND.n464 Folded_Diff_Op_Amp_Layout_0.IND.n461 0.00549102
R22642 Folded_Diff_Op_Amp_Layout_0.IND.n466 Folded_Diff_Op_Amp_Layout_0.IND.n465 0.00549102
R22643 Folded_Diff_Op_Amp_Layout_0.IND.n229 Folded_Diff_Op_Amp_Layout_0.IND.n228 0.00523684
R22644 Folded_Diff_Op_Amp_Layout_0.IND.n242 Folded_Diff_Op_Amp_Layout_0.IND.n241 0.00523684
R22645 Folded_Diff_Op_Amp_Layout_0.IND.n355 Folded_Diff_Op_Amp_Layout_0.IND.n354 0.00523684
R22646 Folded_Diff_Op_Amp_Layout_0.IND.n368 Folded_Diff_Op_Amp_Layout_0.IND.n367 0.00523684
R22647 Folded_Diff_Op_Amp_Layout_0.IND.n381 Folded_Diff_Op_Amp_Layout_0.IND.n380 0.00523684
R22648 Folded_Diff_Op_Amp_Layout_0.IND.n236 Folded_Diff_Op_Amp_Layout_0.IND.n226 0.00479588
R22649 Folded_Diff_Op_Amp_Layout_0.IND.n375 Folded_Diff_Op_Amp_Layout_0.IND.n365 0.00479588
R22650 Folded_Diff_Op_Amp_Layout_0.IND.n212 Folded_Diff_Op_Amp_Layout_0.IND.n205 0.00479588
R22651 Folded_Diff_Op_Amp_Layout_0.IND.n16 Folded_Diff_Op_Amp_Layout_0.IND.n15 0.00364318
R22652 VOUT_OPAMP_P.t27 VOUT_OPAMP_P.t11 147.304
R22653 VOUT_OPAMP_P.t26 VOUT_OPAMP_P.t21 147.304
R22654 VOUT_OPAMP_P.t13 VOUT_OPAMP_P.t23 147.304
R22655 VOUT_OPAMP_P.t30 VOUT_OPAMP_P.t16 147.304
R22656 VOUT_OPAMP_P.n49 VOUT_OPAMP_P.t18 75.0919
R22657 VOUT_OPAMP_P.n17 VOUT_OPAMP_P.t19 74.8891
R22658 VOUT_OPAMP_P.n54 VOUT_OPAMP_P.t8 73.3458
R22659 VOUT_OPAMP_P.n22 VOUT_OPAMP_P.t12 73.143
R22660 VOUT_OPAMP_P.n52 VOUT_OPAMP_P.t26 72.3487
R22661 VOUT_OPAMP_P.n50 VOUT_OPAMP_P.t20 72.3487
R22662 VOUT_OPAMP_P.n48 VOUT_OPAMP_P.t30 72.3487
R22663 VOUT_OPAMP_P.n40 VOUT_OPAMP_P.t14 72.3487
R22664 VOUT_OPAMP_P.n37 VOUT_OPAMP_P.t17 72.3487
R22665 VOUT_OPAMP_P.n20 VOUT_OPAMP_P.t7 72.3487
R22666 VOUT_OPAMP_P.n18 VOUT_OPAMP_P.t29 72.3487
R22667 VOUT_OPAMP_P.n16 VOUT_OPAMP_P.t28 72.3487
R22668 VOUT_OPAMP_P.n52 VOUT_OPAMP_P.t27 51.4916
R22669 VOUT_OPAMP_P.n50 VOUT_OPAMP_P.t25 51.4916
R22670 VOUT_OPAMP_P.n48 VOUT_OPAMP_P.t13 51.4916
R22671 VOUT_OPAMP_P.n40 VOUT_OPAMP_P.t15 51.4916
R22672 VOUT_OPAMP_P.n37 VOUT_OPAMP_P.t24 51.4916
R22673 VOUT_OPAMP_P.n20 VOUT_OPAMP_P.t22 51.4916
R22674 VOUT_OPAMP_P.n18 VOUT_OPAMP_P.t10 51.4916
R22675 VOUT_OPAMP_P.n16 VOUT_OPAMP_P.t9 51.4916
R22676 VOUT_OPAMP_P.n21 VOUT_OPAMP_P.n20 20.1648
R22677 VOUT_OPAMP_P.n17 VOUT_OPAMP_P.n16 20.1648
R22678 VOUT_OPAMP_P.n53 VOUT_OPAMP_P.n52 19.9041
R22679 VOUT_OPAMP_P.n49 VOUT_OPAMP_P.n48 19.9041
R22680 VOUT_OPAMP_P.n51 VOUT_OPAMP_P.n50 15.6747
R22681 VOUT_OPAMP_P.n19 VOUT_OPAMP_P.n18 15.4719
R22682 VOUT_OPAMP_P.n38 VOUT_OPAMP_P.n37 15.1167
R22683 VOUT_OPAMP_P.n41 VOUT_OPAMP_P.n40 12.7876
R22684 VOUT_OPAMP_P.n86 VOUT_OPAMP_P.t4 6.55774
R22685 VOUT_OPAMP_P.n88 VOUT_OPAMP_P.t6 6.43045
R22686 VOUT_OPAMP_P.n87 VOUT_OPAMP_P.t3 6.42009
R22687 VOUT_OPAMP_P.n86 VOUT_OPAMP_P.t2 6.4095
R22688 VOUT_OPAMP_P.n56 VOUT_OPAMP_P.n55 4.52696
R22689 VOUT_OPAMP_P.n31 VOUT_OPAMP_P.n11 4.51065
R22690 VOUT_OPAMP_P.n28 VOUT_OPAMP_P.n15 4.50858
R22691 VOUT_OPAMP_P.n57 VOUT_OPAMP_P.n46 4.50855
R22692 VOUT_OPAMP_P.n59 VOUT_OPAMP_P.n58 4.5005
R22693 VOUT_OPAMP_P.n61 VOUT_OPAMP_P.n60 4.5005
R22694 VOUT_OPAMP_P.n23 VOUT_OPAMP_P.n14 4.5005
R22695 VOUT_OPAMP_P.n29 VOUT_OPAMP_P.n28 4.5005
R22696 VOUT_OPAMP_P.n64 VOUT_OPAMP_P.n12 4.5005
R22697 VOUT_OPAMP_P.n64 VOUT_OPAMP_P.n32 4.5005
R22698 VOUT_OPAMP_P.n69 VOUT_OPAMP_P.n33 4.5005
R22699 VOUT_OPAMP_P.n69 VOUT_OPAMP_P.n30 4.5005
R22700 VOUT_OPAMP_P.n66 VOUT_OPAMP_P.n12 4.5005
R22701 VOUT_OPAMP_P.n66 VOUT_OPAMP_P.n65 4.5005
R22702 VOUT_OPAMP_P.n65 VOUT_OPAMP_P.n64 4.5005
R22703 VOUT_OPAMP_P.n81 VOUT_OPAMP_P.n80 2.82778
R22704 VOUT_OPAMP_P.n2 VOUT_OPAMP_P.t1 2.73276
R22705 VOUT_OPAMP_P.n62 VOUT_OPAMP_P.n44 2.48131
R22706 VOUT_OPAMP_P.n2 VOUT_OPAMP_P.t0 2.40975
R22707 VOUT_OPAMP_P.n60 VOUT_OPAMP_P.n59 2.34524
R22708 VOUT_OPAMP_P.n24 VOUT_OPAMP_P.n23 2.34524
R22709 VOUT_OPAMP_P.n41 VOUT_OPAMP_P.n39 2.26226
R22710 VOUT_OPAMP_P.n60 VOUT_OPAMP_P.n46 2.25517
R22711 VOUT_OPAMP_P.n44 VOUT_OPAMP_P.n43 2.251
R22712 VOUT_OPAMP_P.n90 VOUT_OPAMP_P.n89 2.2505
R22713 VOUT_OPAMP_P.n24 VOUT_OPAMP_P.n15 2.24721
R22714 VOUT_OPAMP_P.n66 VOUT_OPAMP_P.n35 2.24477
R22715 VOUT_OPAMP_P.n67 VOUT_OPAMP_P.n11 2.24477
R22716 VOUT_OPAMP_P.n43 VOUT_OPAMP_P.n38 2.24392
R22717 VOUT_OPAMP_P.n42 VOUT_OPAMP_P.n41 2.24362
R22718 VOUT_OPAMP_P.n26 VOUT_OPAMP_P.n25 2.23629
R22719 VOUT_OPAMP_P.n80 VOUT_OPAMP_P.t5 2.1905
R22720 VOUT_OPAMP_P.n65 VOUT_OPAMP_P.n62 1.8554
R22721 VOUT_OPAMP_P.n42 VOUT_OPAMP_P.n36 1.55989
R22722 VOUT_OPAMP_P.n27 VOUT_OPAMP_P.n26 1.50595
R22723 VOUT_OPAMP_P.n24 VOUT_OPAMP_P.n13 1.50128
R22724 VOUT_OPAMP_P.n39 VOUT_OPAMP_P.n36 1.49987
R22725 VOUT_OPAMP_P.n69 VOUT_OPAMP_P.n31 1.49812
R22726 VOUT_OPAMP_P.n69 VOUT_OPAMP_P.n68 1.49812
R22727 VOUT_OPAMP_P.n34 VOUT_OPAMP_P.n11 1.49801
R22728 VOUT_OPAMP_P.n64 VOUT_OPAMP_P.n63 1.49801
R22729 VOUT_OPAMP_P.n57 VOUT_OPAMP_P.n45 1.49763
R22730 VOUT_OPAMP_P.n1 VOUT_OPAMP_P.n0 1.4964
R22731 VOUT_OPAMP_P.n4 VOUT_OPAMP_P.n3 1.49069
R22732 VOUT_OPAMP_P.n70 VOUT_OPAMP_P.n11 1.15313
R22733 VOUT_OPAMP_P.n70 VOUT_OPAMP_P.n69 1.15091
R22734 VOUT_OPAMP_P.n6 VOUT_OPAMP_P.n5 1.14993
R22735 VOUT_OPAMP_P.n6 VOUT_OPAMP_P.n1 1.14978
R22736 VOUT_OPAMP_P.n74 VOUT_OPAMP_P.n73 1.11304
R22737 VOUT_OPAMP_P.n55 VOUT_OPAMP_P.n47 1.1073
R22738 VOUT_OPAMP_P.n62 VOUT_OPAMP_P.n61 1.09079
R22739 VOUT_OPAMP_P.n27 VOUT_OPAMP_P.n22 0.901569
R22740 VOUT_OPAMP_P.n56 VOUT_OPAMP_P.n54 0.897484
R22741 VOUT_OPAMP_P VOUT_OPAMP_P.n90 0.878717
R22742 VOUT_OPAMP_P VOUT_OPAMP_P.n75 0.728695
R22743 VOUT_OPAMP_P.n7 VOUT_OPAMP_P.n6 0.691886
R22744 VOUT_OPAMP_P.n51 VOUT_OPAMP_P.n49 0.626587
R22745 VOUT_OPAMP_P.n53 VOUT_OPAMP_P.n51 0.626587
R22746 VOUT_OPAMP_P.n19 VOUT_OPAMP_P.n17 0.626587
R22747 VOUT_OPAMP_P.n21 VOUT_OPAMP_P.n19 0.626587
R22748 VOUT_OPAMP_P.n30 VOUT_OPAMP_P.n29 0.51225
R22749 VOUT_OPAMP_P.n71 VOUT_OPAMP_P 0.488719
R22750 VOUT_OPAMP_P.n89 VOUT_OPAMP_P.n88 0.245262
R22751 VOUT_OPAMP_P.n54 VOUT_OPAMP_P.n53 0.239196
R22752 VOUT_OPAMP_P.n22 VOUT_OPAMP_P.n21 0.239196
R22753 VOUT_OPAMP_P.n87 VOUT_OPAMP_P.n86 0.212047
R22754 VOUT_OPAMP_P.n81 VOUT_OPAMP_P.n79 0.141929
R22755 VOUT_OPAMP_P.n83 VOUT_OPAMP_P.n82 0.121357
R22756 VOUT_OPAMP_P.n88 VOUT_OPAMP_P.n87 0.0830882
R22757 VOUT_OPAMP_P.n58 VOUT_OPAMP_P.n47 0.0649899
R22758 VOUT_OPAMP_P.n25 VOUT_OPAMP_P.n24 0.0623855
R22759 VOUT_OPAMP_P.n3 VOUT_OPAMP_P.n2 0.0608233
R22760 VOUT_OPAMP_P.n74 VOUT_OPAMP_P.n10 0.0553537
R22761 VOUT_OPAMP_P.n10 VOUT_OPAMP_P.n9 0.0550978
R22762 VOUT_OPAMP_P.n8 VOUT_OPAMP_P.n7 0.0537258
R22763 VOUT_OPAMP_P.n79 VOUT_OPAMP_P.n78 0.051948
R22764 VOUT_OPAMP_P VOUT_OPAMP_P.n70 0.0432915
R22765 VOUT_OPAMP_P.n25 VOUT_OPAMP_P.n14 0.0339644
R22766 VOUT_OPAMP_P.n60 VOUT_OPAMP_P.n47 0.032498
R22767 VOUT_OPAMP_P.n59 VOUT_OPAMP_P.n54 0.0289211
R22768 VOUT_OPAMP_P.n58 VOUT_OPAMP_P.n57 0.0289211
R22769 VOUT_OPAMP_P.n23 VOUT_OPAMP_P.n22 0.0289211
R22770 VOUT_OPAMP_P.n28 VOUT_OPAMP_P.n14 0.0289211
R22771 VOUT_OPAMP_P.n9 VOUT_OPAMP_P.n8 0.0276709
R22772 VOUT_OPAMP_P.n75 VOUT_OPAMP_P.n74 0.0276709
R22773 VOUT_OPAMP_P.n68 VOUT_OPAMP_P.n67 0.0236139
R22774 VOUT_OPAMP_P.n63 VOUT_OPAMP_P.n35 0.0229474
R22775 VOUT_OPAMP_P.n83 VOUT_OPAMP_P.n81 0.0210714
R22776 VOUT_OPAMP_P.n5 VOUT_OPAMP_P.n4 0.0164591
R22777 VOUT_OPAMP_P.n43 VOUT_OPAMP_P.n42 0.0157541
R22778 VOUT_OPAMP_P.n41 VOUT_OPAMP_P.n38 0.0151658
R22779 VOUT_OPAMP_P.n69 VOUT_OPAMP_P.n12 0.014
R22780 VOUT_OPAMP_P.n69 VOUT_OPAMP_P.n32 0.014
R22781 VOUT_OPAMP_P.n65 VOUT_OPAMP_P.n11 0.014
R22782 VOUT_OPAMP_P.n64 VOUT_OPAMP_P.n33 0.014
R22783 VOUT_OPAMP_P.n67 VOUT_OPAMP_P.n33 0.0134654
R22784 VOUT_OPAMP_P.n35 VOUT_OPAMP_P.n32 0.0134654
R22785 VOUT_OPAMP_P.n73 VOUT_OPAMP_P.n72 0.0122123
R22786 VOUT_OPAMP_P.n29 VOUT_OPAMP_P.n13 0.0117561
R22787 VOUT_OPAMP_P.n72 VOUT_OPAMP_P.n71 0.0113904
R22788 VOUT_OPAMP_P.n61 VOUT_OPAMP_P.n45 0.0111023
R22789 VOUT_OPAMP_P.n90 VOUT_OPAMP_P.n77 0.0108185
R22790 VOUT_OPAMP_P.n34 VOUT_OPAMP_P.n30 0.00998204
R22791 VOUT_OPAMP_P.n55 VOUT_OPAMP_P.n46 0.00860784
R22792 VOUT_OPAMP_P.n44 VOUT_OPAMP_P.n36 0.00859375
R22793 VOUT_OPAMP_P.n26 VOUT_OPAMP_P.n15 0.00858096
R22794 VOUT_OPAMP_P.n85 VOUT_OPAMP_P.n84 0.00764286
R22795 VOUT_OPAMP_P.n57 VOUT_OPAMP_P.n56 0.00685938
R22796 VOUT_OPAMP_P.n26 VOUT_OPAMP_P.n13 0.00639619
R22797 VOUT_OPAMP_P.n77 VOUT_OPAMP_P.n76 0.00623248
R22798 VOUT_OPAMP_P.n43 VOUT_OPAMP_P.n39 0.00621251
R22799 VOUT_OPAMP_P.n55 VOUT_OPAMP_P.n45 0.00605114
R22800 VOUT_OPAMP_P.n68 VOUT_OPAMP_P.n66 0.00582347
R22801 VOUT_OPAMP_P.n64 VOUT_OPAMP_P.n31 0.00582347
R22802 VOUT_OPAMP_P.n63 VOUT_OPAMP_P.n11 0.00549102
R22803 VOUT_OPAMP_P.n66 VOUT_OPAMP_P.n34 0.00549102
R22804 VOUT_OPAMP_P.n28 VOUT_OPAMP_P.n27 0.00400424
R22805 VOUT_OPAMP_P.n84 VOUT_OPAMP_P.n83 0.00240476
R22806 VOUT_OPAMP_P.n89 VOUT_OPAMP_P.n85 0.00192857
R22807 Folded_Diff_Op_Amp_Layout_0.IPD.n301 Folded_Diff_Op_Amp_Layout_0.IPD.n300 5.29686
R22808 Folded_Diff_Op_Amp_Layout_0.IPD.n282 Folded_Diff_Op_Amp_Layout_0.IPD.t35 5.29686
R22809 Folded_Diff_Op_Amp_Layout_0.IPD.n167 Folded_Diff_Op_Amp_Layout_0.IPD.n166 4.97729
R22810 Folded_Diff_Op_Amp_Layout_0.IPD.n148 Folded_Diff_Op_Amp_Layout_0.IPD.t60 4.97729
R22811 Folded_Diff_Op_Amp_Layout_0.IPD.n37 Folded_Diff_Op_Amp_Layout_0.IPD.n36 4.86858
R22812 Folded_Diff_Op_Amp_Layout_0.IPD.n288 Folded_Diff_Op_Amp_Layout_0.IPD.n287 4.72811
R22813 Folded_Diff_Op_Amp_Layout_0.IPD.n52 Folded_Diff_Op_Amp_Layout_0.IPD.n51 4.71629
R22814 Folded_Diff_Op_Amp_Layout_0.IPD.n154 Folded_Diff_Op_Amp_Layout_0.IPD.n153 4.40854
R22815 Folded_Diff_Op_Amp_Layout_0.IPD.n277 Folded_Diff_Op_Amp_Layout_0.IPD.n276 2.41042
R22816 Folded_Diff_Op_Amp_Layout_0.IPD.n351 Folded_Diff_Op_Amp_Layout_0.IPD.n349 1.6654
R22817 Folded_Diff_Op_Amp_Layout_0.IPD.n376 Folded_Diff_Op_Amp_Layout_0.IPD.t39 1.6654
R22818 Folded_Diff_Op_Amp_Layout_0.IPD.n33 Folded_Diff_Op_Amp_Layout_0.IPD.n32 1.64142
R22819 Folded_Diff_Op_Amp_Layout_0.IPD.n438 Folded_Diff_Op_Amp_Layout_0.IPD.n434 1.49801
R22820 Folded_Diff_Op_Amp_Layout_0.IPD.n410 Folded_Diff_Op_Amp_Layout_0.IPD.n409 1.49801
R22821 Folded_Diff_Op_Amp_Layout_0.IPD.n229 Folded_Diff_Op_Amp_Layout_0.IPD.n228 1.48953
R22822 Folded_Diff_Op_Amp_Layout_0.IPD.n321 Folded_Diff_Op_Amp_Layout_0.IPD.n30 1.48953
R22823 Folded_Diff_Op_Amp_Layout_0.IPD.n343 Folded_Diff_Op_Amp_Layout_0.IPD.n342 1.48953
R22824 Folded_Diff_Op_Amp_Layout_0.IPD.n142 Folded_Diff_Op_Amp_Layout_0.IPD.n141 1.47785
R22825 Folded_Diff_Op_Amp_Layout_0.IPD.n131 Folded_Diff_Op_Amp_Layout_0.IPD.t52 1.47785
R22826 Folded_Diff_Op_Amp_Layout_0.IPD.n203 Folded_Diff_Op_Amp_Layout_0.IPD.t22 1.31982
R22827 Folded_Diff_Op_Amp_Layout_0.IPD.n199 Folded_Diff_Op_Amp_Layout_0.IPD.n198 1.31982
R22828 Folded_Diff_Op_Amp_Layout_0.IPD.n6 Folded_Diff_Op_Amp_Layout_0.IPD.t18 1.30711
R22829 Folded_Diff_Op_Amp_Layout_0.IPD.n2 Folded_Diff_Op_Amp_Layout_0.IPD.n1 1.30711
R22830 Folded_Diff_Op_Amp_Layout_0.IPD.n298 Folded_Diff_Op_Amp_Layout_0.IPD.n297 1.28973
R22831 Folded_Diff_Op_Amp_Layout_0.IPD.n293 Folded_Diff_Op_Amp_Layout_0.IPD.n292 1.28973
R22832 Folded_Diff_Op_Amp_Layout_0.IPD.n280 Folded_Diff_Op_Amp_Layout_0.IPD.n279 1.28973
R22833 Folded_Diff_Op_Amp_Layout_0.IPD.n138 Folded_Diff_Op_Amp_Layout_0.IPD.n137 1.19571
R22834 Folded_Diff_Op_Amp_Layout_0.IPD.n332 Folded_Diff_Op_Amp_Layout_0.IPD.n331 1.19534
R22835 Folded_Diff_Op_Amp_Layout_0.IPD.n396 Folded_Diff_Op_Amp_Layout_0.IPD.n395 1.19519
R22836 Folded_Diff_Op_Amp_Layout_0.IPD.n18 Folded_Diff_Op_Amp_Layout_0.IPD.n17 1.19509
R22837 Folded_Diff_Op_Amp_Layout_0.IPD.n7 Folded_Diff_Op_Amp_Layout_0.IPD.n6 1.19506
R22838 Folded_Diff_Op_Amp_Layout_0.IPD.n71 Folded_Diff_Op_Amp_Layout_0.IPD.n70 1.19466
R22839 Folded_Diff_Op_Amp_Layout_0.IPD.n261 Folded_Diff_Op_Amp_Layout_0.IPD.n260 1.19444
R22840 Folded_Diff_Op_Amp_Layout_0.IPD.n420 Folded_Diff_Op_Amp_Layout_0.IPD.n419 1.1943
R22841 Folded_Diff_Op_Amp_Layout_0.IPD.n215 Folded_Diff_Op_Amp_Layout_0.IPD.n214 1.19395
R22842 Folded_Diff_Op_Amp_Layout_0.IPD.n204 Folded_Diff_Op_Amp_Layout_0.IPD.n203 1.19393
R22843 Folded_Diff_Op_Amp_Layout_0.IPD.n49 Folded_Diff_Op_Amp_Layout_0.IPD.n48 1.18349
R22844 Folded_Diff_Op_Amp_Layout_0.IPD.n267 Folded_Diff_Op_Amp_Layout_0.IPD.n266 1.17941
R22845 Folded_Diff_Op_Amp_Layout_0.IPD.n122 Folded_Diff_Op_Amp_Layout_0.IPD.n121 1.17929
R22846 Folded_Diff_Op_Amp_Layout_0.IPD.n415 Folded_Diff_Op_Amp_Layout_0.IPD.n414 1.17902
R22847 Folded_Diff_Op_Amp_Layout_0.IPD.n111 Folded_Diff_Op_Amp_Layout_0.IPD.n110 1.17902
R22848 Folded_Diff_Op_Amp_Layout_0.IPD.n65 Folded_Diff_Op_Amp_Layout_0.IPD.n64 1.17891
R22849 Folded_Diff_Op_Amp_Layout_0.IPD.n200 Folded_Diff_Op_Amp_Layout_0.IPD.n199 1.1787
R22850 Folded_Diff_Op_Amp_Layout_0.IPD.n326 Folded_Diff_Op_Amp_Layout_0.IPD.n325 1.1782
R22851 Folded_Diff_Op_Amp_Layout_0.IPD.n143 Folded_Diff_Op_Amp_Layout_0.IPD.n142 1.17812
R22852 Folded_Diff_Op_Amp_Layout_0.IPD.n132 Folded_Diff_Op_Amp_Layout_0.IPD.n131 1.17812
R22853 Folded_Diff_Op_Amp_Layout_0.IPD.n390 Folded_Diff_Op_Amp_Layout_0.IPD.n389 1.17768
R22854 Folded_Diff_Op_Amp_Layout_0.IPD.n3 Folded_Diff_Op_Amp_Layout_0.IPD.n2 1.17753
R22855 Folded_Diff_Op_Amp_Layout_0.IPD.n439 Folded_Diff_Op_Amp_Layout_0.IPD.n385 1.1775
R22856 Folded_Diff_Op_Amp_Layout_0.IPD.n299 Folded_Diff_Op_Amp_Layout_0.IPD.n298 1.17428
R22857 Folded_Diff_Op_Amp_Layout_0.IPD.n294 Folded_Diff_Op_Amp_Layout_0.IPD.n293 1.17428
R22858 Folded_Diff_Op_Amp_Layout_0.IPD.n281 Folded_Diff_Op_Amp_Layout_0.IPD.n280 1.17428
R22859 Folded_Diff_Op_Amp_Layout_0.IPD.n367 Folded_Diff_Op_Amp_Layout_0.IPD.n366 1.16675
R22860 Folded_Diff_Op_Amp_Layout_0.IPD.n165 Folded_Diff_Op_Amp_Layout_0.IPD.n164 1.16619
R22861 Folded_Diff_Op_Amp_Layout_0.IPD.n160 Folded_Diff_Op_Amp_Layout_0.IPD.n159 1.16619
R22862 Folded_Diff_Op_Amp_Layout_0.IPD.n147 Folded_Diff_Op_Amp_Layout_0.IPD.n146 1.16619
R22863 Folded_Diff_Op_Amp_Layout_0.IPD.n239 Folded_Diff_Op_Amp_Layout_0.IPD.n238 1.16617
R22864 Folded_Diff_Op_Amp_Layout_0.IPD.n352 Folded_Diff_Op_Amp_Layout_0.IPD.n351 1.16588
R22865 Folded_Diff_Op_Amp_Layout_0.IPD.n377 Folded_Diff_Op_Amp_Layout_0.IPD.n376 1.16588
R22866 Folded_Diff_Op_Amp_Layout_0.IPD.n81 Folded_Diff_Op_Amp_Layout_0.IPD.n80 1.16562
R22867 Folded_Diff_Op_Amp_Layout_0.IPD.n252 Folded_Diff_Op_Amp_Layout_0.IPD.n251 1.1656
R22868 Folded_Diff_Op_Amp_Layout_0.IPD.n94 Folded_Diff_Op_Amp_Layout_0.IPD.n93 1.16506
R22869 Folded_Diff_Op_Amp_Layout_0.IPD.n320 Folded_Diff_Op_Amp_Layout_0.IPD.n60 1.1515
R22870 Folded_Diff_Op_Amp_Layout_0.IPD.n34 Folded_Diff_Op_Amp_Layout_0.IPD.n33 1.14576
R22871 Folded_Diff_Op_Amp_Layout_0.IPD.n368 Folded_Diff_Op_Amp_Layout_0.IPD.n367 1.1257
R22872 Folded_Diff_Op_Amp_Layout_0.IPD.n39 Folded_Diff_Op_Amp_Layout_0.IPD.n38 1.1255
R22873 Folded_Diff_Op_Amp_Layout_0.IPD.n54 Folded_Diff_Op_Amp_Layout_0.IPD.n53 1.1255
R22874 Folded_Diff_Op_Amp_Layout_0.IPD.n303 Folded_Diff_Op_Amp_Layout_0.IPD.n302 1.1255
R22875 Folded_Diff_Op_Amp_Layout_0.IPD.n284 Folded_Diff_Op_Amp_Layout_0.IPD.n283 1.1255
R22876 Folded_Diff_Op_Amp_Layout_0.IPD.n290 Folded_Diff_Op_Amp_Layout_0.IPD.n289 1.1255
R22877 Folded_Diff_Op_Amp_Layout_0.IPD.n169 Folded_Diff_Op_Amp_Layout_0.IPD.n168 1.1255
R22878 Folded_Diff_Op_Amp_Layout_0.IPD.n156 Folded_Diff_Op_Amp_Layout_0.IPD.n155 1.1255
R22879 Folded_Diff_Op_Amp_Layout_0.IPD.n150 Folded_Diff_Op_Amp_Layout_0.IPD.n149 1.1255
R22880 Folded_Diff_Op_Amp_Layout_0.IPD.n319 Folded_Diff_Op_Amp_Layout_0.IPD.n318 1.1255
R22881 Folded_Diff_Op_Amp_Layout_0.IPD.n439 Folded_Diff_Op_Amp_Layout_0.IPD.n438 1.1255
R22882 Folded_Diff_Op_Amp_Layout_0.IPD.n241 Folded_Diff_Op_Amp_Layout_0.IPD.n240 1.10737
R22883 Folded_Diff_Op_Amp_Layout_0.IPD.n83 Folded_Diff_Op_Amp_Layout_0.IPD.n82 1.10737
R22884 Folded_Diff_Op_Amp_Layout_0.IPD.n354 Folded_Diff_Op_Amp_Layout_0.IPD.n353 1.1073
R22885 Folded_Diff_Op_Amp_Layout_0.IPD.n379 Folded_Diff_Op_Amp_Layout_0.IPD.n378 1.1073
R22886 Folded_Diff_Op_Amp_Layout_0.IPD.n93 Folded_Diff_Op_Amp_Layout_0.IPD.n92 1.09806
R22887 Folded_Diff_Op_Amp_Layout_0.IPD.n80 Folded_Diff_Op_Amp_Layout_0.IPD.n79 1.09777
R22888 Folded_Diff_Op_Amp_Layout_0.IPD.n251 Folded_Diff_Op_Amp_Layout_0.IPD.n250 1.09692
R22889 Folded_Diff_Op_Amp_Layout_0.IPD.n238 Folded_Diff_Op_Amp_Layout_0.IPD.n237 1.09663
R22890 Folded_Diff_Op_Amp_Layout_0.IPD.n366 Folded_Diff_Op_Amp_Layout_0.IPD.n364 1.09644
R22891 Folded_Diff_Op_Amp_Layout_0.IPD.n256 Folded_Diff_Op_Amp_Layout_0.IPD.n255 1.08123
R22892 Folded_Diff_Op_Amp_Layout_0.IPD.n164 Folded_Diff_Op_Amp_Layout_0.IPD.n163 1.07378
R22893 Folded_Diff_Op_Amp_Layout_0.IPD.n159 Folded_Diff_Op_Amp_Layout_0.IPD.n158 1.07378
R22894 Folded_Diff_Op_Amp_Layout_0.IPD.n146 Folded_Diff_Op_Amp_Layout_0.IPD.n145 1.07378
R22895 Folded_Diff_Op_Amp_Layout_0.IPD.n98 Folded_Diff_Op_Amp_Layout_0.IPD.n97 0.939312
R22896 Folded_Diff_Op_Amp_Layout_0.IPD.n70 Folded_Diff_Op_Amp_Layout_0.IPD.n69 0.922529
R22897 Folded_Diff_Op_Amp_Layout_0.IPD.n64 Folded_Diff_Op_Amp_Layout_0.IPD.n63 0.922508
R22898 Folded_Diff_Op_Amp_Layout_0.IPD.n266 Folded_Diff_Op_Amp_Layout_0.IPD.n265 0.920678
R22899 Folded_Diff_Op_Amp_Layout_0.IPD.n260 Folded_Diff_Op_Amp_Layout_0.IPD.n259 0.920678
R22900 Folded_Diff_Op_Amp_Layout_0.IPD.n331 Folded_Diff_Op_Amp_Layout_0.IPD.n330 0.913532
R22901 Folded_Diff_Op_Amp_Layout_0.IPD.n325 Folded_Diff_Op_Amp_Layout_0.IPD.n324 0.913527
R22902 Folded_Diff_Op_Amp_Layout_0.IPD.n395 Folded_Diff_Op_Amp_Layout_0.IPD.n394 0.911021
R22903 Folded_Diff_Op_Amp_Layout_0.IPD.n389 Folded_Diff_Op_Amp_Layout_0.IPD.n388 0.911021
R22904 Folded_Diff_Op_Amp_Layout_0.IPD.n137 Folded_Diff_Op_Amp_Layout_0.IPD.n136 0.909101
R22905 Folded_Diff_Op_Amp_Layout_0.IPD.n382 Folded_Diff_Op_Amp_Layout_0.IPD.n381 0.901232
R22906 Folded_Diff_Op_Amp_Layout_0.IPD.n254 Folded_Diff_Op_Amp_Layout_0.IPD.n253 0.88565
R22907 Folded_Diff_Op_Amp_Layout_0.IPD.n96 Folded_Diff_Op_Amp_Layout_0.IPD.n95 0.88565
R22908 Folded_Diff_Op_Amp_Layout_0.IPD.n424 Folded_Diff_Op_Amp_Layout_0.IPD.n422 0.88565
R22909 Folded_Diff_Op_Amp_Layout_0.IPD.n121 Folded_Diff_Op_Amp_Layout_0.IPD.n120 0.834379
R22910 Folded_Diff_Op_Amp_Layout_0.IPD.n414 Folded_Diff_Op_Amp_Layout_0.IPD.n413 0.834365
R22911 Folded_Diff_Op_Amp_Layout_0.IPD.n110 Folded_Diff_Op_Amp_Layout_0.IPD.n109 0.834365
R22912 Folded_Diff_Op_Amp_Layout_0.IPD.n419 Folded_Diff_Op_Amp_Layout_0.IPD.n418 0.834251
R22913 Folded_Diff_Op_Amp_Layout_0.IPD.n214 Folded_Diff_Op_Amp_Layout_0.IPD.n213 0.834193
R22914 Folded_Diff_Op_Amp_Layout_0.IPD.n17 Folded_Diff_Op_Amp_Layout_0.IPD.n16 0.821487
R22915 Folded_Diff_Op_Amp_Layout_0.IPD.n21 Folded_Diff_Op_Amp_Layout_0.IPD.n20 0.727916
R22916 Folded_Diff_Op_Amp_Layout_0.IPD.n57 Folded_Diff_Op_Amp_Layout_0.IPD.n56 0.727916
R22917 Folded_Diff_Op_Amp_Layout_0.IPD.n218 Folded_Diff_Op_Amp_Layout_0.IPD.n217 0.727916
R22918 Folded_Diff_Op_Amp_Layout_0.IPD.n125 Folded_Diff_Op_Amp_Layout_0.IPD.n124 0.727916
R22919 Folded_Diff_Op_Amp_Layout_0.IPD.n26 Folded_Diff_Op_Amp_Layout_0.IPD.n4 0.727104
R22920 Folded_Diff_Op_Amp_Layout_0.IPD.n335 Folded_Diff_Op_Amp_Layout_0.IPD.n333 0.727104
R22921 Folded_Diff_Op_Amp_Layout_0.IPD.n310 Folded_Diff_Op_Amp_Layout_0.IPD.n295 0.727104
R22922 Folded_Diff_Op_Amp_Layout_0.IPD.n270 Folded_Diff_Op_Amp_Layout_0.IPD.n268 0.727104
R22923 Folded_Diff_Op_Amp_Layout_0.IPD.n223 Folded_Diff_Op_Amp_Layout_0.IPD.n201 0.727104
R22924 Folded_Diff_Op_Amp_Layout_0.IPD.n172 Folded_Diff_Op_Amp_Layout_0.IPD.n170 0.727104
R22925 Folded_Diff_Op_Amp_Layout_0.IPD.n181 Folded_Diff_Op_Amp_Layout_0.IPD.n151 0.727104
R22926 Folded_Diff_Op_Amp_Layout_0.IPD.n190 Folded_Diff_Op_Amp_Layout_0.IPD.n139 0.727104
R22927 Folded_Diff_Op_Amp_Layout_0.IPD.n100 Folded_Diff_Op_Amp_Layout_0.IPD.n72 0.727104
R22928 Folded_Diff_Op_Amp_Layout_0.IPD.n403 Folded_Diff_Op_Amp_Layout_0.IPD.n391 0.727104
R22929 Folded_Diff_Op_Amp_Layout_0.IPD.n129 Folded_Diff_Op_Amp_Layout_0.IPD.n128 0.691748
R22930 Folded_Diff_Op_Amp_Layout_0.IPD.n128 Folded_Diff_Op_Amp_Layout_0.IPD.n127 0.648341
R22931 Folded_Diff_Op_Amp_Layout_0.IPD.n278 Folded_Diff_Op_Amp_Layout_0.IPD.n277 0.632522
R22932 Folded_Diff_Op_Amp_Layout_0.IPD.n431 Folded_Diff_Op_Amp_Layout_0.IPD.n430 0.628687
R22933 Folded_Diff_Op_Amp_Layout_0.IPD.n60 Folded_Diff_Op_Amp_Layout_0.IPD.n59 0.623188
R22934 Folded_Diff_Op_Amp_Layout_0.IPD.n428 Folded_Diff_Op_Amp_Layout_0.IPD.n416 0.616779
R22935 Folded_Diff_Op_Amp_Layout_0.IPD.n10 Folded_Diff_Op_Amp_Layout_0.IPD.n8 0.616779
R22936 Folded_Diff_Op_Amp_Layout_0.IPD.n340 Folded_Diff_Op_Amp_Layout_0.IPD.n327 0.616779
R22937 Folded_Diff_Op_Amp_Layout_0.IPD.n42 Folded_Diff_Op_Amp_Layout_0.IPD.n40 0.616779
R22938 Folded_Diff_Op_Amp_Layout_0.IPD.n306 Folded_Diff_Op_Amp_Layout_0.IPD.n304 0.616779
R22939 Folded_Diff_Op_Amp_Layout_0.IPD.n315 Folded_Diff_Op_Amp_Layout_0.IPD.n285 0.616779
R22940 Folded_Diff_Op_Amp_Layout_0.IPD.n275 Folded_Diff_Op_Amp_Layout_0.IPD.n262 0.616779
R22941 Folded_Diff_Op_Amp_Layout_0.IPD.n207 Folded_Diff_Op_Amp_Layout_0.IPD.n205 0.616779
R22942 Folded_Diff_Op_Amp_Layout_0.IPD.n177 Folded_Diff_Op_Amp_Layout_0.IPD.n161 0.616779
R22943 Folded_Diff_Op_Amp_Layout_0.IPD.n186 Folded_Diff_Op_Amp_Layout_0.IPD.n144 0.616779
R22944 Folded_Diff_Op_Amp_Layout_0.IPD.n195 Folded_Diff_Op_Amp_Layout_0.IPD.n133 0.616779
R22945 Folded_Diff_Op_Amp_Layout_0.IPD.n114 Folded_Diff_Op_Amp_Layout_0.IPD.n112 0.616779
R22946 Folded_Diff_Op_Amp_Layout_0.IPD.n105 Folded_Diff_Op_Amp_Layout_0.IPD.n66 0.616779
R22947 Folded_Diff_Op_Amp_Layout_0.IPD.n399 Folded_Diff_Op_Amp_Layout_0.IPD.n397 0.616779
R22948 Folded_Diff_Op_Amp_Layout_0.IPD.n364 Folded_Diff_Op_Amp_Layout_0.IPD.t32 0.56925
R22949 Folded_Diff_Op_Amp_Layout_0.IPD.n364 Folded_Diff_Op_Amp_Layout_0.IPD.n363 0.56925
R22950 Folded_Diff_Op_Amp_Layout_0.IPD.n330 Folded_Diff_Op_Amp_Layout_0.IPD.t27 0.56925
R22951 Folded_Diff_Op_Amp_Layout_0.IPD.n330 Folded_Diff_Op_Amp_Layout_0.IPD.n329 0.56925
R22952 Folded_Diff_Op_Amp_Layout_0.IPD.n324 Folded_Diff_Op_Amp_Layout_0.IPD.t41 0.56925
R22953 Folded_Diff_Op_Amp_Layout_0.IPD.n324 Folded_Diff_Op_Amp_Layout_0.IPD.n323 0.56925
R22954 Folded_Diff_Op_Amp_Layout_0.IPD.n297 Folded_Diff_Op_Amp_Layout_0.IPD.n296 0.56925
R22955 Folded_Diff_Op_Amp_Layout_0.IPD.n292 Folded_Diff_Op_Amp_Layout_0.IPD.t47 0.56925
R22956 Folded_Diff_Op_Amp_Layout_0.IPD.n292 Folded_Diff_Op_Amp_Layout_0.IPD.n291 0.56925
R22957 Folded_Diff_Op_Amp_Layout_0.IPD.n287 Folded_Diff_Op_Amp_Layout_0.IPD.t53 0.56925
R22958 Folded_Diff_Op_Amp_Layout_0.IPD.n287 Folded_Diff_Op_Amp_Layout_0.IPD.n286 0.56925
R22959 Folded_Diff_Op_Amp_Layout_0.IPD.n279 Folded_Diff_Op_Amp_Layout_0.IPD.t25 0.56925
R22960 Folded_Diff_Op_Amp_Layout_0.IPD.n265 Folded_Diff_Op_Amp_Layout_0.IPD.t71 0.56925
R22961 Folded_Diff_Op_Amp_Layout_0.IPD.n265 Folded_Diff_Op_Amp_Layout_0.IPD.n264 0.56925
R22962 Folded_Diff_Op_Amp_Layout_0.IPD.n259 Folded_Diff_Op_Amp_Layout_0.IPD.t59 0.56925
R22963 Folded_Diff_Op_Amp_Layout_0.IPD.n259 Folded_Diff_Op_Amp_Layout_0.IPD.n258 0.56925
R22964 Folded_Diff_Op_Amp_Layout_0.IPD.n237 Folded_Diff_Op_Amp_Layout_0.IPD.t49 0.56925
R22965 Folded_Diff_Op_Amp_Layout_0.IPD.n237 Folded_Diff_Op_Amp_Layout_0.IPD.n236 0.56925
R22966 Folded_Diff_Op_Amp_Layout_0.IPD.n250 Folded_Diff_Op_Amp_Layout_0.IPD.t29 0.56925
R22967 Folded_Diff_Op_Amp_Layout_0.IPD.n250 Folded_Diff_Op_Amp_Layout_0.IPD.n249 0.56925
R22968 Folded_Diff_Op_Amp_Layout_0.IPD.n163 Folded_Diff_Op_Amp_Layout_0.IPD.n162 0.56925
R22969 Folded_Diff_Op_Amp_Layout_0.IPD.n153 Folded_Diff_Op_Amp_Layout_0.IPD.t63 0.56925
R22970 Folded_Diff_Op_Amp_Layout_0.IPD.n153 Folded_Diff_Op_Amp_Layout_0.IPD.n152 0.56925
R22971 Folded_Diff_Op_Amp_Layout_0.IPD.n158 Folded_Diff_Op_Amp_Layout_0.IPD.t68 0.56925
R22972 Folded_Diff_Op_Amp_Layout_0.IPD.n158 Folded_Diff_Op_Amp_Layout_0.IPD.n157 0.56925
R22973 Folded_Diff_Op_Amp_Layout_0.IPD.n145 Folded_Diff_Op_Amp_Layout_0.IPD.t70 0.56925
R22974 Folded_Diff_Op_Amp_Layout_0.IPD.n136 Folded_Diff_Op_Amp_Layout_0.IPD.t33 0.56925
R22975 Folded_Diff_Op_Amp_Layout_0.IPD.n136 Folded_Diff_Op_Amp_Layout_0.IPD.n135 0.56925
R22976 Folded_Diff_Op_Amp_Layout_0.IPD.n79 Folded_Diff_Op_Amp_Layout_0.IPD.t65 0.56925
R22977 Folded_Diff_Op_Amp_Layout_0.IPD.n79 Folded_Diff_Op_Amp_Layout_0.IPD.n78 0.56925
R22978 Folded_Diff_Op_Amp_Layout_0.IPD.n92 Folded_Diff_Op_Amp_Layout_0.IPD.t66 0.56925
R22979 Folded_Diff_Op_Amp_Layout_0.IPD.n92 Folded_Diff_Op_Amp_Layout_0.IPD.n91 0.56925
R22980 Folded_Diff_Op_Amp_Layout_0.IPD.n69 Folded_Diff_Op_Amp_Layout_0.IPD.t46 0.56925
R22981 Folded_Diff_Op_Amp_Layout_0.IPD.n69 Folded_Diff_Op_Amp_Layout_0.IPD.n68 0.56925
R22982 Folded_Diff_Op_Amp_Layout_0.IPD.n63 Folded_Diff_Op_Amp_Layout_0.IPD.t24 0.56925
R22983 Folded_Diff_Op_Amp_Layout_0.IPD.n63 Folded_Diff_Op_Amp_Layout_0.IPD.n62 0.56925
R22984 Folded_Diff_Op_Amp_Layout_0.IPD.n394 Folded_Diff_Op_Amp_Layout_0.IPD.t38 0.56925
R22985 Folded_Diff_Op_Amp_Layout_0.IPD.n394 Folded_Diff_Op_Amp_Layout_0.IPD.n393 0.56925
R22986 Folded_Diff_Op_Amp_Layout_0.IPD.n388 Folded_Diff_Op_Amp_Layout_0.IPD.t55 0.56925
R22987 Folded_Diff_Op_Amp_Layout_0.IPD.n388 Folded_Diff_Op_Amp_Layout_0.IPD.n387 0.56925
R22988 Folded_Diff_Op_Amp_Layout_0.IPD.n256 Folded_Diff_Op_Amp_Layout_0.IPD.n230 0.526243
R22989 Folded_Diff_Op_Amp_Layout_0.IPD.n128 Folded_Diff_Op_Amp_Layout_0.IPD.n106 0.524913
R22990 Folded_Diff_Op_Amp_Layout_0.IPD.n342 Folded_Diff_Op_Amp_Layout_0.IPD.n341 0.516188
R22991 Folded_Diff_Op_Amp_Layout_0.IPD.n184 Folded_Diff_Op_Amp_Layout_0.IPD.n183 0.507313
R22992 Folded_Diff_Op_Amp_Layout_0.IPD.n406 Folded_Diff_Op_Amp_Layout_0.IPD.n405 0.502687
R22993 Folded_Diff_Op_Amp_Layout_0.IPD.n383 Folded_Diff_Op_Amp_Layout_0.IPD.n382 0.500334
R22994 Folded_Diff_Op_Amp_Layout_0.IPD.n413 Folded_Diff_Op_Amp_Layout_0.IPD.t2 0.485833
R22995 Folded_Diff_Op_Amp_Layout_0.IPD.n413 Folded_Diff_Op_Amp_Layout_0.IPD.n412 0.485833
R22996 Folded_Diff_Op_Amp_Layout_0.IPD.n16 Folded_Diff_Op_Amp_Layout_0.IPD.t1 0.485833
R22997 Folded_Diff_Op_Amp_Layout_0.IPD.n16 Folded_Diff_Op_Amp_Layout_0.IPD.n15 0.485833
R22998 Folded_Diff_Op_Amp_Layout_0.IPD.n32 Folded_Diff_Op_Amp_Layout_0.IPD.t9 0.485833
R22999 Folded_Diff_Op_Amp_Layout_0.IPD.n32 Folded_Diff_Op_Amp_Layout_0.IPD.n31 0.485833
R23000 Folded_Diff_Op_Amp_Layout_0.IPD.n36 Folded_Diff_Op_Amp_Layout_0.IPD.t4 0.485833
R23001 Folded_Diff_Op_Amp_Layout_0.IPD.n36 Folded_Diff_Op_Amp_Layout_0.IPD.n35 0.485833
R23002 Folded_Diff_Op_Amp_Layout_0.IPD.n48 Folded_Diff_Op_Amp_Layout_0.IPD.t14 0.485833
R23003 Folded_Diff_Op_Amp_Layout_0.IPD.n48 Folded_Diff_Op_Amp_Layout_0.IPD.n47 0.485833
R23004 Folded_Diff_Op_Amp_Layout_0.IPD.n51 Folded_Diff_Op_Amp_Layout_0.IPD.t0 0.485833
R23005 Folded_Diff_Op_Amp_Layout_0.IPD.n51 Folded_Diff_Op_Amp_Layout_0.IPD.n50 0.485833
R23006 Folded_Diff_Op_Amp_Layout_0.IPD.n213 Folded_Diff_Op_Amp_Layout_0.IPD.t10 0.485833
R23007 Folded_Diff_Op_Amp_Layout_0.IPD.n213 Folded_Diff_Op_Amp_Layout_0.IPD.n212 0.485833
R23008 Folded_Diff_Op_Amp_Layout_0.IPD.n109 Folded_Diff_Op_Amp_Layout_0.IPD.t16 0.485833
R23009 Folded_Diff_Op_Amp_Layout_0.IPD.n109 Folded_Diff_Op_Amp_Layout_0.IPD.n108 0.485833
R23010 Folded_Diff_Op_Amp_Layout_0.IPD.n120 Folded_Diff_Op_Amp_Layout_0.IPD.t13 0.485833
R23011 Folded_Diff_Op_Amp_Layout_0.IPD.n120 Folded_Diff_Op_Amp_Layout_0.IPD.n119 0.485833
R23012 Folded_Diff_Op_Amp_Layout_0.IPD.n418 Folded_Diff_Op_Amp_Layout_0.IPD.t23 0.485833
R23013 Folded_Diff_Op_Amp_Layout_0.IPD.n418 Folded_Diff_Op_Amp_Layout_0.IPD.n417 0.485833
R23014 Folded_Diff_Op_Amp_Layout_0.IPD.n273 Folded_Diff_Op_Amp_Layout_0.IPD.n272 0.474125
R23015 Folded_Diff_Op_Amp_Layout_0.IPD.n175 Folded_Diff_Op_Amp_Layout_0.IPD.n174 0.474125
R23016 Folded_Diff_Op_Amp_Layout_0.IPD.n179 Folded_Diff_Op_Amp_Layout_0.IPD.n178 0.474125
R23017 Folded_Diff_Op_Amp_Layout_0.IPD.n86 Folded_Diff_Op_Amp_Layout_0.IPD.n85 0.474125
R23018 Folded_Diff_Op_Amp_Layout_0.IPD.n29 Folded_Diff_Op_Amp_Layout_0.IPD.n28 0.46275
R23019 Folded_Diff_Op_Amp_Layout_0.IPD.n226 Folded_Diff_Op_Amp_Layout_0.IPD.n225 0.46275
R23020 Folded_Diff_Op_Amp_Layout_0.IPD.n53 Folded_Diff_Op_Amp_Layout_0.IPD.n52 0.447377
R23021 Folded_Diff_Op_Amp_Layout_0.IPD.n321 Folded_Diff_Op_Amp_Layout_0.IPD.n320 0.352375
R23022 Folded_Diff_Op_Amp_Layout_0.IPD.n228 Folded_Diff_Op_Amp_Layout_0.IPD.n196 0.336187
R23023 Folded_Diff_Op_Amp_Layout_0.IPD.n45 Folded_Diff_Op_Amp_Layout_0.IPD.n44 0.330687
R23024 Folded_Diff_Op_Amp_Layout_0.IPD.n117 Folded_Diff_Op_Amp_Layout_0.IPD.n116 0.330687
R23025 Folded_Diff_Op_Amp_Layout_0.IPD.n427 Folded_Diff_Op_Amp_Layout_0.IPD.n426 0.330687
R23026 Folded_Diff_Op_Amp_Layout_0.IPD.n357 Folded_Diff_Op_Amp_Layout_0.IPD.n356 0.330125
R23027 Folded_Diff_Op_Amp_Layout_0.IPD.n370 Folded_Diff_Op_Amp_Layout_0.IPD.n369 0.330125
R23028 Folded_Diff_Op_Amp_Layout_0.IPD.n24 Folded_Diff_Op_Amp_Layout_0.IPD.n23 0.330125
R23029 Folded_Diff_Op_Amp_Layout_0.IPD.n13 Folded_Diff_Op_Amp_Layout_0.IPD.n12 0.330125
R23030 Folded_Diff_Op_Amp_Layout_0.IPD.n338 Folded_Diff_Op_Amp_Layout_0.IPD.n337 0.330125
R23031 Folded_Diff_Op_Amp_Layout_0.IPD.n308 Folded_Diff_Op_Amp_Layout_0.IPD.n307 0.330125
R23032 Folded_Diff_Op_Amp_Layout_0.IPD.n313 Folded_Diff_Op_Amp_Layout_0.IPD.n312 0.330125
R23033 Folded_Diff_Op_Amp_Layout_0.IPD.n244 Folded_Diff_Op_Amp_Layout_0.IPD.n243 0.330125
R23034 Folded_Diff_Op_Amp_Layout_0.IPD.n221 Folded_Diff_Op_Amp_Layout_0.IPD.n220 0.330125
R23035 Folded_Diff_Op_Amp_Layout_0.IPD.n210 Folded_Diff_Op_Amp_Layout_0.IPD.n209 0.330125
R23036 Folded_Diff_Op_Amp_Layout_0.IPD.n188 Folded_Diff_Op_Amp_Layout_0.IPD.n187 0.330125
R23037 Folded_Diff_Op_Amp_Layout_0.IPD.n193 Folded_Diff_Op_Amp_Layout_0.IPD.n192 0.330125
R23038 Folded_Diff_Op_Amp_Layout_0.IPD.n103 Folded_Diff_Op_Amp_Layout_0.IPD.n102 0.330125
R23039 Folded_Diff_Op_Amp_Layout_0.IPD.n401 Folded_Diff_Op_Amp_Layout_0.IPD.n400 0.330125
R23040 Folded_Diff_Op_Amp_Layout_0.IPD.n317 Folded_Diff_Op_Amp_Layout_0.IPD.n316 0.317187
R23041 Folded_Diff_Op_Amp_Layout_0.IPD.n38 Folded_Diff_Op_Amp_Layout_0.IPD.n37 0.269474
R23042 Folded_Diff_Op_Amp_Layout_0.IPD.n382 Folded_Diff_Op_Amp_Layout_0.IPD.n344 0.268618
R23043 Folded_Diff_Op_Amp_Layout_0.IPD.n277 Folded_Diff_Op_Amp_Layout_0.IPD.n256 0.248389
R23044 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.IPD.n439 0.241687
R23045 Folded_Diff_Op_Amp_Layout_0.IPD.n302 Folded_Diff_Op_Amp_Layout_0.IPD.n301 0.235932
R23046 Folded_Diff_Op_Amp_Layout_0.IPD.n289 Folded_Diff_Op_Amp_Layout_0.IPD.n288 0.235932
R23047 Folded_Diff_Op_Amp_Layout_0.IPD.n283 Folded_Diff_Op_Amp_Layout_0.IPD.n282 0.235932
R23048 Folded_Diff_Op_Amp_Layout_0.IPD.n168 Folded_Diff_Op_Amp_Layout_0.IPD.n167 0.12963
R23049 Folded_Diff_Op_Amp_Layout_0.IPD.n155 Folded_Diff_Op_Amp_Layout_0.IPD.n154 0.12963
R23050 Folded_Diff_Op_Amp_Layout_0.IPD.n149 Folded_Diff_Op_Amp_Layout_0.IPD.n148 0.12963
R23051 Folded_Diff_Op_Amp_Layout_0.IPD.n422 Folded_Diff_Op_Amp_Layout_0.IPD.n421 0.0995747
R23052 Folded_Diff_Op_Amp_Layout_0.IPD.n253 Folded_Diff_Op_Amp_Layout_0.IPD.n247 0.0936537
R23053 Folded_Diff_Op_Amp_Layout_0.IPD.n95 Folded_Diff_Op_Amp_Layout_0.IPD.n89 0.0912853
R23054 Folded_Diff_Op_Amp_Layout_0.IPD.n353 Folded_Diff_Op_Amp_Layout_0.IPD.n348 0.0886741
R23055 Folded_Diff_Op_Amp_Layout_0.IPD.n378 Folded_Diff_Op_Amp_Layout_0.IPD.n374 0.0886741
R23056 Folded_Diff_Op_Amp_Layout_0.IPD.n240 Folded_Diff_Op_Amp_Layout_0.IPD.n234 0.0880141
R23057 Folded_Diff_Op_Amp_Layout_0.IPD.n82 Folded_Diff_Op_Amp_Layout_0.IPD.n76 0.0856456
R23058 Folded_Diff_Op_Amp_Layout_0.IPD.n20 Folded_Diff_Op_Amp_Layout_0.IPD.n19 0.0826464
R23059 Folded_Diff_Op_Amp_Layout_0.IPD.n56 Folded_Diff_Op_Amp_Layout_0.IPD.n55 0.0826464
R23060 Folded_Diff_Op_Amp_Layout_0.IPD.n217 Folded_Diff_Op_Amp_Layout_0.IPD.n216 0.0826464
R23061 Folded_Diff_Op_Amp_Layout_0.IPD.n124 Folded_Diff_Op_Amp_Layout_0.IPD.n123 0.0826464
R23062 Folded_Diff_Op_Amp_Layout_0.IPD.n4 Folded_Diff_Op_Amp_Layout_0.IPD.n0 0.0823987
R23063 Folded_Diff_Op_Amp_Layout_0.IPD.n333 Folded_Diff_Op_Amp_Layout_0.IPD.n328 0.0823987
R23064 Folded_Diff_Op_Amp_Layout_0.IPD.n295 Folded_Diff_Op_Amp_Layout_0.IPD.n290 0.0823987
R23065 Folded_Diff_Op_Amp_Layout_0.IPD.n268 Folded_Diff_Op_Amp_Layout_0.IPD.n263 0.0823987
R23066 Folded_Diff_Op_Amp_Layout_0.IPD.n201 Folded_Diff_Op_Amp_Layout_0.IPD.n197 0.0823987
R23067 Folded_Diff_Op_Amp_Layout_0.IPD.n170 Folded_Diff_Op_Amp_Layout_0.IPD.n165 0.0823987
R23068 Folded_Diff_Op_Amp_Layout_0.IPD.n151 Folded_Diff_Op_Amp_Layout_0.IPD.n147 0.0823987
R23069 Folded_Diff_Op_Amp_Layout_0.IPD.n139 Folded_Diff_Op_Amp_Layout_0.IPD.n134 0.0823987
R23070 Folded_Diff_Op_Amp_Layout_0.IPD.n72 Folded_Diff_Op_Amp_Layout_0.IPD.n67 0.0823987
R23071 Folded_Diff_Op_Amp_Layout_0.IPD.n391 Folded_Diff_Op_Amp_Layout_0.IPD.n386 0.0823987
R23072 Folded_Diff_Op_Amp_Layout_0.IPD.n366 Folded_Diff_Op_Amp_Layout_0.IPD.n365 0.0784141
R23073 Folded_Diff_Op_Amp_Layout_0.IPD.n351 Folded_Diff_Op_Amp_Layout_0.IPD.n350 0.0783056
R23074 Folded_Diff_Op_Amp_Layout_0.IPD.n376 Folded_Diff_Op_Amp_Layout_0.IPD.n375 0.0783056
R23075 Folded_Diff_Op_Amp_Layout_0.IPD.n238 Folded_Diff_Op_Amp_Layout_0.IPD.n235 0.0778549
R23076 Folded_Diff_Op_Amp_Layout_0.IPD.n251 Folded_Diff_Op_Amp_Layout_0.IPD.n248 0.0774429
R23077 Folded_Diff_Op_Amp_Layout_0.IPD.n53 Folded_Diff_Op_Amp_Layout_0.IPD.n49 0.0761444
R23078 Folded_Diff_Op_Amp_Layout_0.IPD.n80 Folded_Diff_Op_Amp_Layout_0.IPD.n77 0.0761073
R23079 Folded_Diff_Op_Amp_Layout_0.IPD.n93 Folded_Diff_Op_Amp_Layout_0.IPD.n90 0.0756955
R23080 Folded_Diff_Op_Amp_Layout_0.IPD.n8 Folded_Diff_Op_Amp_Layout_0.IPD.n5 0.0712285
R23081 Folded_Diff_Op_Amp_Layout_0.IPD.n327 Folded_Diff_Op_Amp_Layout_0.IPD.n322 0.0712285
R23082 Folded_Diff_Op_Amp_Layout_0.IPD.n40 Folded_Diff_Op_Amp_Layout_0.IPD.n34 0.0712285
R23083 Folded_Diff_Op_Amp_Layout_0.IPD.n285 Folded_Diff_Op_Amp_Layout_0.IPD.n281 0.0712285
R23084 Folded_Diff_Op_Amp_Layout_0.IPD.n304 Folded_Diff_Op_Amp_Layout_0.IPD.n299 0.0712285
R23085 Folded_Diff_Op_Amp_Layout_0.IPD.n262 Folded_Diff_Op_Amp_Layout_0.IPD.n257 0.0712285
R23086 Folded_Diff_Op_Amp_Layout_0.IPD.n205 Folded_Diff_Op_Amp_Layout_0.IPD.n202 0.0712285
R23087 Folded_Diff_Op_Amp_Layout_0.IPD.n133 Folded_Diff_Op_Amp_Layout_0.IPD.n130 0.0712285
R23088 Folded_Diff_Op_Amp_Layout_0.IPD.n144 Folded_Diff_Op_Amp_Layout_0.IPD.n140 0.0712285
R23089 Folded_Diff_Op_Amp_Layout_0.IPD.n161 Folded_Diff_Op_Amp_Layout_0.IPD.n156 0.0712285
R23090 Folded_Diff_Op_Amp_Layout_0.IPD.n112 Folded_Diff_Op_Amp_Layout_0.IPD.n107 0.0712285
R23091 Folded_Diff_Op_Amp_Layout_0.IPD.n66 Folded_Diff_Op_Amp_Layout_0.IPD.n61 0.0712285
R23092 Folded_Diff_Op_Amp_Layout_0.IPD.n397 Folded_Diff_Op_Amp_Layout_0.IPD.n392 0.0712285
R23093 Folded_Diff_Op_Amp_Layout_0.IPD.n416 Folded_Diff_Op_Amp_Layout_0.IPD.n411 0.0712285
R23094 Folded_Diff_Op_Amp_Layout_0.IPD.n367 Folded_Diff_Op_Amp_Layout_0.IPD.n362 0.0623855
R23095 Folded_Diff_Op_Amp_Layout_0.IPD.n362 Folded_Diff_Op_Amp_Layout_0.IPD.n361 0.0576486
R23096 Folded_Diff_Op_Amp_Layout_0.IPD.n8 Folded_Diff_Op_Amp_Layout_0.IPD.n7 0.0534597
R23097 Folded_Diff_Op_Amp_Layout_0.IPD.n327 Folded_Diff_Op_Amp_Layout_0.IPD.n326 0.0534597
R23098 Folded_Diff_Op_Amp_Layout_0.IPD.n40 Folded_Diff_Op_Amp_Layout_0.IPD.n39 0.0534597
R23099 Folded_Diff_Op_Amp_Layout_0.IPD.n304 Folded_Diff_Op_Amp_Layout_0.IPD.n303 0.0534597
R23100 Folded_Diff_Op_Amp_Layout_0.IPD.n285 Folded_Diff_Op_Amp_Layout_0.IPD.n284 0.0534597
R23101 Folded_Diff_Op_Amp_Layout_0.IPD.n262 Folded_Diff_Op_Amp_Layout_0.IPD.n261 0.0534597
R23102 Folded_Diff_Op_Amp_Layout_0.IPD.n205 Folded_Diff_Op_Amp_Layout_0.IPD.n204 0.0534597
R23103 Folded_Diff_Op_Amp_Layout_0.IPD.n161 Folded_Diff_Op_Amp_Layout_0.IPD.n160 0.0534597
R23104 Folded_Diff_Op_Amp_Layout_0.IPD.n144 Folded_Diff_Op_Amp_Layout_0.IPD.n143 0.0534597
R23105 Folded_Diff_Op_Amp_Layout_0.IPD.n133 Folded_Diff_Op_Amp_Layout_0.IPD.n132 0.0534597
R23106 Folded_Diff_Op_Amp_Layout_0.IPD.n112 Folded_Diff_Op_Amp_Layout_0.IPD.n111 0.0534597
R23107 Folded_Diff_Op_Amp_Layout_0.IPD.n66 Folded_Diff_Op_Amp_Layout_0.IPD.n65 0.0534597
R23108 Folded_Diff_Op_Amp_Layout_0.IPD.n397 Folded_Diff_Op_Amp_Layout_0.IPD.n396 0.0534597
R23109 Folded_Diff_Op_Amp_Layout_0.IPD.n416 Folded_Diff_Op_Amp_Layout_0.IPD.n415 0.0534597
R23110 Folded_Diff_Op_Amp_Layout_0.IPD.n320 Folded_Diff_Op_Amp_Layout_0.IPD.n319 0.0525
R23111 Folded_Diff_Op_Amp_Layout_0.IPD.n319 Folded_Diff_Op_Amp_Layout_0.IPD.n278 0.0525
R23112 Folded_Diff_Op_Amp_Layout_0.IPD.n20 Folded_Diff_Op_Amp_Layout_0.IPD.n18 0.0423164
R23113 Folded_Diff_Op_Amp_Layout_0.IPD.n56 Folded_Diff_Op_Amp_Layout_0.IPD.n54 0.0423164
R23114 Folded_Diff_Op_Amp_Layout_0.IPD.n217 Folded_Diff_Op_Amp_Layout_0.IPD.n215 0.0423164
R23115 Folded_Diff_Op_Amp_Layout_0.IPD.n124 Folded_Diff_Op_Amp_Layout_0.IPD.n122 0.0423164
R23116 Folded_Diff_Op_Amp_Layout_0.IPD.n4 Folded_Diff_Op_Amp_Layout_0.IPD.n3 0.0415773
R23117 Folded_Diff_Op_Amp_Layout_0.IPD.n333 Folded_Diff_Op_Amp_Layout_0.IPD.n332 0.0415773
R23118 Folded_Diff_Op_Amp_Layout_0.IPD.n295 Folded_Diff_Op_Amp_Layout_0.IPD.n294 0.0415773
R23119 Folded_Diff_Op_Amp_Layout_0.IPD.n268 Folded_Diff_Op_Amp_Layout_0.IPD.n267 0.0415773
R23120 Folded_Diff_Op_Amp_Layout_0.IPD.n201 Folded_Diff_Op_Amp_Layout_0.IPD.n200 0.0415773
R23121 Folded_Diff_Op_Amp_Layout_0.IPD.n139 Folded_Diff_Op_Amp_Layout_0.IPD.n138 0.0415773
R23122 Folded_Diff_Op_Amp_Layout_0.IPD.n151 Folded_Diff_Op_Amp_Layout_0.IPD.n150 0.0415773
R23123 Folded_Diff_Op_Amp_Layout_0.IPD.n170 Folded_Diff_Op_Amp_Layout_0.IPD.n169 0.0415773
R23124 Folded_Diff_Op_Amp_Layout_0.IPD.n72 Folded_Diff_Op_Amp_Layout_0.IPD.n71 0.0415773
R23125 Folded_Diff_Op_Amp_Layout_0.IPD.n391 Folded_Diff_Op_Amp_Layout_0.IPD.n390 0.0415773
R23126 Folded_Diff_Op_Amp_Layout_0.IPD.n228 Folded_Diff_Op_Amp_Layout_0.IPD.n227 0.0354016
R23127 Folded_Diff_Op_Amp_Layout_0.IPD.n229 Folded_Diff_Op_Amp_Layout_0.IPD.n129 0.0354016
R23128 Folded_Diff_Op_Amp_Layout_0.IPD.n343 Folded_Diff_Op_Amp_Layout_0.IPD.n321 0.0354016
R23129 Folded_Diff_Op_Amp_Layout_0.IPD.n378 Folded_Diff_Op_Amp_Layout_0.IPD.n377 0.032498
R23130 Folded_Diff_Op_Amp_Layout_0.IPD.n353 Folded_Diff_Op_Amp_Layout_0.IPD.n352 0.032498
R23131 Folded_Diff_Op_Amp_Layout_0.IPD.n240 Folded_Diff_Op_Amp_Layout_0.IPD.n239 0.0319869
R23132 Folded_Diff_Op_Amp_Layout_0.IPD.n82 Folded_Diff_Op_Amp_Layout_0.IPD.n81 0.0319869
R23133 Folded_Diff_Op_Amp_Layout_0.IPD.n318 Folded_Diff_Op_Amp_Layout_0.IPD.n317 0.0265
R23134 Folded_Diff_Op_Amp_Layout_0.IPD.n253 Folded_Diff_Op_Amp_Layout_0.IPD.n252 0.0261793
R23135 Folded_Diff_Op_Amp_Layout_0.IPD.n95 Folded_Diff_Op_Amp_Layout_0.IPD.n94 0.0261793
R23136 Folded_Diff_Op_Amp_Layout_0.IPD.n422 Folded_Diff_Op_Amp_Layout_0.IPD.n420 0.0261793
R23137 Folded_Diff_Op_Amp_Layout_0.IPD.n436 Folded_Diff_Op_Amp_Layout_0.IPD.n435 0.0207053
R23138 Folded_Diff_Op_Amp_Layout_0.IPD.n408 Folded_Diff_Op_Amp_Layout_0.IPD.n407 0.0207053
R23139 Folded_Diff_Op_Amp_Layout_0.IPD.n30 Folded_Diff_Op_Amp_Layout_0.IPD.n29 0.0182008
R23140 Folded_Diff_Op_Amp_Layout_0.IPD.n227 Folded_Diff_Op_Amp_Layout_0.IPD.n226 0.0182008
R23141 Folded_Diff_Op_Amp_Layout_0.IPD.n230 Folded_Diff_Op_Amp_Layout_0.IPD.n229 0.0182008
R23142 Folded_Diff_Op_Amp_Layout_0.IPD.n344 Folded_Diff_Op_Amp_Layout_0.IPD.n343 0.0182008
R23143 Folded_Diff_Op_Amp_Layout_0.IPD.n358 Folded_Diff_Op_Amp_Layout_0.IPD.n357 0.0156875
R23144 Folded_Diff_Op_Amp_Layout_0.IPD.n10 Folded_Diff_Op_Amp_Layout_0.IPD.n9 0.0156875
R23145 Folded_Diff_Op_Amp_Layout_0.IPD.n341 Folded_Diff_Op_Amp_Layout_0.IPD.n340 0.0156875
R23146 Folded_Diff_Op_Amp_Layout_0.IPD.n42 Folded_Diff_Op_Amp_Layout_0.IPD.n41 0.0156875
R23147 Folded_Diff_Op_Amp_Layout_0.IPD.n307 Folded_Diff_Op_Amp_Layout_0.IPD.n306 0.0156875
R23148 Folded_Diff_Op_Amp_Layout_0.IPD.n316 Folded_Diff_Op_Amp_Layout_0.IPD.n315 0.0156875
R23149 Folded_Diff_Op_Amp_Layout_0.IPD.n276 Folded_Diff_Op_Amp_Layout_0.IPD.n275 0.0156875
R23150 Folded_Diff_Op_Amp_Layout_0.IPD.n254 Folded_Diff_Op_Amp_Layout_0.IPD.n244 0.0156875
R23151 Folded_Diff_Op_Amp_Layout_0.IPD.n255 Folded_Diff_Op_Amp_Layout_0.IPD.n254 0.0156875
R23152 Folded_Diff_Op_Amp_Layout_0.IPD.n207 Folded_Diff_Op_Amp_Layout_0.IPD.n206 0.0156875
R23153 Folded_Diff_Op_Amp_Layout_0.IPD.n178 Folded_Diff_Op_Amp_Layout_0.IPD.n177 0.0156875
R23154 Folded_Diff_Op_Amp_Layout_0.IPD.n187 Folded_Diff_Op_Amp_Layout_0.IPD.n186 0.0156875
R23155 Folded_Diff_Op_Amp_Layout_0.IPD.n196 Folded_Diff_Op_Amp_Layout_0.IPD.n195 0.0156875
R23156 Folded_Diff_Op_Amp_Layout_0.IPD.n114 Folded_Diff_Op_Amp_Layout_0.IPD.n113 0.0156875
R23157 Folded_Diff_Op_Amp_Layout_0.IPD.n96 Folded_Diff_Op_Amp_Layout_0.IPD.n86 0.0156875
R23158 Folded_Diff_Op_Amp_Layout_0.IPD.n97 Folded_Diff_Op_Amp_Layout_0.IPD.n96 0.0156875
R23159 Folded_Diff_Op_Amp_Layout_0.IPD.n106 Folded_Diff_Op_Amp_Layout_0.IPD.n105 0.0156875
R23160 Folded_Diff_Op_Amp_Layout_0.IPD.n400 Folded_Diff_Op_Amp_Layout_0.IPD.n399 0.0156875
R23161 Folded_Diff_Op_Amp_Layout_0.IPD.n428 Folded_Diff_Op_Amp_Layout_0.IPD.n427 0.0156875
R23162 Folded_Diff_Op_Amp_Layout_0.IPD.n438 Folded_Diff_Op_Amp_Layout_0.IPD.n437 0.014
R23163 Folded_Diff_Op_Amp_Layout_0.IPD.n409 Folded_Diff_Op_Amp_Layout_0.IPD.n406 0.014
R23164 Folded_Diff_Op_Amp_Layout_0.IPD.n373 Folded_Diff_Op_Amp_Layout_0.IPD.n372 0.0139513
R23165 Folded_Diff_Op_Amp_Layout_0.IPD.n347 Folded_Diff_Op_Amp_Layout_0.IPD.n346 0.0139513
R23166 Folded_Diff_Op_Amp_Layout_0.IPD.n437 Folded_Diff_Op_Amp_Layout_0.IPD.n436 0.0134654
R23167 Folded_Diff_Op_Amp_Layout_0.IPD.n233 Folded_Diff_Op_Amp_Layout_0.IPD.n232 0.0133659
R23168 Folded_Diff_Op_Amp_Layout_0.IPD.n369 Folded_Diff_Op_Amp_Layout_0.IPD.n368 0.0123533
R23169 Folded_Diff_Op_Amp_Layout_0.IPD.n75 Folded_Diff_Op_Amp_Layout_0.IPD.n74 0.012194
R23170 Folded_Diff_Op_Amp_Layout_0.IPD.n356 Folded_Diff_Op_Amp_Layout_0.IPD.n355 0.0111023
R23171 Folded_Diff_Op_Amp_Layout_0.IPD.n381 Folded_Diff_Op_Amp_Layout_0.IPD.n380 0.0111023
R23172 Folded_Diff_Op_Amp_Layout_0.IPD.n243 Folded_Diff_Op_Amp_Layout_0.IPD.n242 0.0111023
R23173 Folded_Diff_Op_Amp_Layout_0.IPD.n85 Folded_Diff_Op_Amp_Layout_0.IPD.n84 0.0111023
R23174 Folded_Diff_Op_Amp_Layout_0.IPD.n426 Folded_Diff_Op_Amp_Layout_0.IPD.n425 0.0111023
R23175 Folded_Diff_Op_Amp_Layout_0.IPD.n434 Folded_Diff_Op_Amp_Layout_0.IPD.n431 0.00998204
R23176 Folded_Diff_Op_Amp_Layout_0.IPD.n76 Folded_Diff_Op_Amp_Layout_0.IPD.n75 0.00878947
R23177 Folded_Diff_Op_Amp_Layout_0.IPD.n89 Folded_Diff_Op_Amp_Layout_0.IPD.n88 0.00878947
R23178 Folded_Diff_Op_Amp_Layout_0.IPD.n429 Folded_Diff_Op_Amp_Layout_0.IPD.n428 0.00860784
R23179 Folded_Diff_Op_Amp_Layout_0.IPD.n354 Folded_Diff_Op_Amp_Layout_0.IPD.n345 0.00860784
R23180 Folded_Diff_Op_Amp_Layout_0.IPD.n379 Folded_Diff_Op_Amp_Layout_0.IPD.n371 0.00860784
R23181 Folded_Diff_Op_Amp_Layout_0.IPD.n11 Folded_Diff_Op_Amp_Layout_0.IPD.n10 0.00860784
R23182 Folded_Diff_Op_Amp_Layout_0.IPD.n26 Folded_Diff_Op_Amp_Layout_0.IPD.n25 0.00860784
R23183 Folded_Diff_Op_Amp_Layout_0.IPD.n336 Folded_Diff_Op_Amp_Layout_0.IPD.n335 0.00860784
R23184 Folded_Diff_Op_Amp_Layout_0.IPD.n340 Folded_Diff_Op_Amp_Layout_0.IPD.n339 0.00860784
R23185 Folded_Diff_Op_Amp_Layout_0.IPD.n43 Folded_Diff_Op_Amp_Layout_0.IPD.n42 0.00860784
R23186 Folded_Diff_Op_Amp_Layout_0.IPD.n306 Folded_Diff_Op_Amp_Layout_0.IPD.n305 0.00860784
R23187 Folded_Diff_Op_Amp_Layout_0.IPD.n311 Folded_Diff_Op_Amp_Layout_0.IPD.n310 0.00860784
R23188 Folded_Diff_Op_Amp_Layout_0.IPD.n315 Folded_Diff_Op_Amp_Layout_0.IPD.n314 0.00860784
R23189 Folded_Diff_Op_Amp_Layout_0.IPD.n271 Folded_Diff_Op_Amp_Layout_0.IPD.n270 0.00860784
R23190 Folded_Diff_Op_Amp_Layout_0.IPD.n275 Folded_Diff_Op_Amp_Layout_0.IPD.n274 0.00860784
R23191 Folded_Diff_Op_Amp_Layout_0.IPD.n241 Folded_Diff_Op_Amp_Layout_0.IPD.n231 0.00860784
R23192 Folded_Diff_Op_Amp_Layout_0.IPD.n208 Folded_Diff_Op_Amp_Layout_0.IPD.n207 0.00860784
R23193 Folded_Diff_Op_Amp_Layout_0.IPD.n223 Folded_Diff_Op_Amp_Layout_0.IPD.n222 0.00860784
R23194 Folded_Diff_Op_Amp_Layout_0.IPD.n173 Folded_Diff_Op_Amp_Layout_0.IPD.n172 0.00860784
R23195 Folded_Diff_Op_Amp_Layout_0.IPD.n177 Folded_Diff_Op_Amp_Layout_0.IPD.n176 0.00860784
R23196 Folded_Diff_Op_Amp_Layout_0.IPD.n182 Folded_Diff_Op_Amp_Layout_0.IPD.n181 0.00860784
R23197 Folded_Diff_Op_Amp_Layout_0.IPD.n186 Folded_Diff_Op_Amp_Layout_0.IPD.n185 0.00860784
R23198 Folded_Diff_Op_Amp_Layout_0.IPD.n191 Folded_Diff_Op_Amp_Layout_0.IPD.n190 0.00860784
R23199 Folded_Diff_Op_Amp_Layout_0.IPD.n195 Folded_Diff_Op_Amp_Layout_0.IPD.n194 0.00860784
R23200 Folded_Diff_Op_Amp_Layout_0.IPD.n115 Folded_Diff_Op_Amp_Layout_0.IPD.n114 0.00860784
R23201 Folded_Diff_Op_Amp_Layout_0.IPD.n83 Folded_Diff_Op_Amp_Layout_0.IPD.n73 0.00860784
R23202 Folded_Diff_Op_Amp_Layout_0.IPD.n101 Folded_Diff_Op_Amp_Layout_0.IPD.n100 0.00860784
R23203 Folded_Diff_Op_Amp_Layout_0.IPD.n105 Folded_Diff_Op_Amp_Layout_0.IPD.n104 0.00860784
R23204 Folded_Diff_Op_Amp_Layout_0.IPD.n399 Folded_Diff_Op_Amp_Layout_0.IPD.n398 0.00860784
R23205 Folded_Diff_Op_Amp_Layout_0.IPD.n404 Folded_Diff_Op_Amp_Layout_0.IPD.n403 0.00860784
R23206 Folded_Diff_Op_Amp_Layout_0.IPD.n424 Folded_Diff_Op_Amp_Layout_0.IPD.n423 0.00860784
R23207 Folded_Diff_Op_Amp_Layout_0.IPD.n28 Folded_Diff_Op_Amp_Layout_0.IPD.n27 0.00858096
R23208 Folded_Diff_Op_Amp_Layout_0.IPD.n22 Folded_Diff_Op_Amp_Layout_0.IPD.n21 0.00858096
R23209 Folded_Diff_Op_Amp_Layout_0.IPD.n14 Folded_Diff_Op_Amp_Layout_0.IPD.n13 0.00858096
R23210 Folded_Diff_Op_Amp_Layout_0.IPD.n27 Folded_Diff_Op_Amp_Layout_0.IPD.n26 0.00858096
R23211 Folded_Diff_Op_Amp_Layout_0.IPD.n23 Folded_Diff_Op_Amp_Layout_0.IPD.n22 0.00858096
R23212 Folded_Diff_Op_Amp_Layout_0.IPD.n21 Folded_Diff_Op_Amp_Layout_0.IPD.n14 0.00858096
R23213 Folded_Diff_Op_Amp_Layout_0.IPD.n335 Folded_Diff_Op_Amp_Layout_0.IPD.n334 0.00858096
R23214 Folded_Diff_Op_Amp_Layout_0.IPD.n58 Folded_Diff_Op_Amp_Layout_0.IPD.n57 0.00858096
R23215 Folded_Diff_Op_Amp_Layout_0.IPD.n46 Folded_Diff_Op_Amp_Layout_0.IPD.n45 0.00858096
R23216 Folded_Diff_Op_Amp_Layout_0.IPD.n59 Folded_Diff_Op_Amp_Layout_0.IPD.n58 0.00858096
R23217 Folded_Diff_Op_Amp_Layout_0.IPD.n57 Folded_Diff_Op_Amp_Layout_0.IPD.n46 0.00858096
R23218 Folded_Diff_Op_Amp_Layout_0.IPD.n309 Folded_Diff_Op_Amp_Layout_0.IPD.n308 0.00858096
R23219 Folded_Diff_Op_Amp_Layout_0.IPD.n310 Folded_Diff_Op_Amp_Layout_0.IPD.n309 0.00858096
R23220 Folded_Diff_Op_Amp_Layout_0.IPD.n270 Folded_Diff_Op_Amp_Layout_0.IPD.n269 0.00858096
R23221 Folded_Diff_Op_Amp_Layout_0.IPD.n225 Folded_Diff_Op_Amp_Layout_0.IPD.n224 0.00858096
R23222 Folded_Diff_Op_Amp_Layout_0.IPD.n219 Folded_Diff_Op_Amp_Layout_0.IPD.n218 0.00858096
R23223 Folded_Diff_Op_Amp_Layout_0.IPD.n211 Folded_Diff_Op_Amp_Layout_0.IPD.n210 0.00858096
R23224 Folded_Diff_Op_Amp_Layout_0.IPD.n224 Folded_Diff_Op_Amp_Layout_0.IPD.n223 0.00858096
R23225 Folded_Diff_Op_Amp_Layout_0.IPD.n220 Folded_Diff_Op_Amp_Layout_0.IPD.n219 0.00858096
R23226 Folded_Diff_Op_Amp_Layout_0.IPD.n218 Folded_Diff_Op_Amp_Layout_0.IPD.n211 0.00858096
R23227 Folded_Diff_Op_Amp_Layout_0.IPD.n180 Folded_Diff_Op_Amp_Layout_0.IPD.n179 0.00858096
R23228 Folded_Diff_Op_Amp_Layout_0.IPD.n189 Folded_Diff_Op_Amp_Layout_0.IPD.n188 0.00858096
R23229 Folded_Diff_Op_Amp_Layout_0.IPD.n190 Folded_Diff_Op_Amp_Layout_0.IPD.n189 0.00858096
R23230 Folded_Diff_Op_Amp_Layout_0.IPD.n181 Folded_Diff_Op_Amp_Layout_0.IPD.n180 0.00858096
R23231 Folded_Diff_Op_Amp_Layout_0.IPD.n172 Folded_Diff_Op_Amp_Layout_0.IPD.n171 0.00858096
R23232 Folded_Diff_Op_Amp_Layout_0.IPD.n126 Folded_Diff_Op_Amp_Layout_0.IPD.n125 0.00858096
R23233 Folded_Diff_Op_Amp_Layout_0.IPD.n118 Folded_Diff_Op_Amp_Layout_0.IPD.n117 0.00858096
R23234 Folded_Diff_Op_Amp_Layout_0.IPD.n127 Folded_Diff_Op_Amp_Layout_0.IPD.n126 0.00858096
R23235 Folded_Diff_Op_Amp_Layout_0.IPD.n125 Folded_Diff_Op_Amp_Layout_0.IPD.n118 0.00858096
R23236 Folded_Diff_Op_Amp_Layout_0.IPD.n99 Folded_Diff_Op_Amp_Layout_0.IPD.n98 0.00858096
R23237 Folded_Diff_Op_Amp_Layout_0.IPD.n100 Folded_Diff_Op_Amp_Layout_0.IPD.n99 0.00858096
R23238 Folded_Diff_Op_Amp_Layout_0.IPD.n402 Folded_Diff_Op_Amp_Layout_0.IPD.n401 0.00858096
R23239 Folded_Diff_Op_Amp_Layout_0.IPD.n403 Folded_Diff_Op_Amp_Layout_0.IPD.n402 0.00858096
R23240 Folded_Diff_Op_Amp_Layout_0.IPD.n371 Folded_Diff_Op_Amp_Layout_0.IPD.n370 0.00855417
R23241 Folded_Diff_Op_Amp_Layout_0.IPD.n25 Folded_Diff_Op_Amp_Layout_0.IPD.n24 0.00855417
R23242 Folded_Diff_Op_Amp_Layout_0.IPD.n12 Folded_Diff_Op_Amp_Layout_0.IPD.n11 0.00855417
R23243 Folded_Diff_Op_Amp_Layout_0.IPD.n337 Folded_Diff_Op_Amp_Layout_0.IPD.n336 0.00855417
R23244 Folded_Diff_Op_Amp_Layout_0.IPD.n339 Folded_Diff_Op_Amp_Layout_0.IPD.n338 0.00855417
R23245 Folded_Diff_Op_Amp_Layout_0.IPD.n44 Folded_Diff_Op_Amp_Layout_0.IPD.n43 0.00855417
R23246 Folded_Diff_Op_Amp_Layout_0.IPD.n312 Folded_Diff_Op_Amp_Layout_0.IPD.n311 0.00855417
R23247 Folded_Diff_Op_Amp_Layout_0.IPD.n314 Folded_Diff_Op_Amp_Layout_0.IPD.n313 0.00855417
R23248 Folded_Diff_Op_Amp_Layout_0.IPD.n272 Folded_Diff_Op_Amp_Layout_0.IPD.n271 0.00855417
R23249 Folded_Diff_Op_Amp_Layout_0.IPD.n274 Folded_Diff_Op_Amp_Layout_0.IPD.n273 0.00855417
R23250 Folded_Diff_Op_Amp_Layout_0.IPD.n222 Folded_Diff_Op_Amp_Layout_0.IPD.n221 0.00855417
R23251 Folded_Diff_Op_Amp_Layout_0.IPD.n209 Folded_Diff_Op_Amp_Layout_0.IPD.n208 0.00855417
R23252 Folded_Diff_Op_Amp_Layout_0.IPD.n174 Folded_Diff_Op_Amp_Layout_0.IPD.n173 0.00855417
R23253 Folded_Diff_Op_Amp_Layout_0.IPD.n176 Folded_Diff_Op_Amp_Layout_0.IPD.n175 0.00855417
R23254 Folded_Diff_Op_Amp_Layout_0.IPD.n183 Folded_Diff_Op_Amp_Layout_0.IPD.n182 0.00855417
R23255 Folded_Diff_Op_Amp_Layout_0.IPD.n185 Folded_Diff_Op_Amp_Layout_0.IPD.n184 0.00855417
R23256 Folded_Diff_Op_Amp_Layout_0.IPD.n192 Folded_Diff_Op_Amp_Layout_0.IPD.n191 0.00855417
R23257 Folded_Diff_Op_Amp_Layout_0.IPD.n194 Folded_Diff_Op_Amp_Layout_0.IPD.n193 0.00855417
R23258 Folded_Diff_Op_Amp_Layout_0.IPD.n116 Folded_Diff_Op_Amp_Layout_0.IPD.n115 0.00855417
R23259 Folded_Diff_Op_Amp_Layout_0.IPD.n102 Folded_Diff_Op_Amp_Layout_0.IPD.n101 0.00855417
R23260 Folded_Diff_Op_Amp_Layout_0.IPD.n104 Folded_Diff_Op_Amp_Layout_0.IPD.n103 0.00855417
R23261 Folded_Diff_Op_Amp_Layout_0.IPD.n405 Folded_Diff_Op_Amp_Layout_0.IPD.n404 0.00855417
R23262 Folded_Diff_Op_Amp_Layout_0.IPD.n430 Folded_Diff_Op_Amp_Layout_0.IPD.n429 0.00855417
R23263 Folded_Diff_Op_Amp_Layout_0.IPD.n384 Folded_Diff_Op_Amp_Layout_0.IPD.n383 0.00773989
R23264 Folded_Diff_Op_Amp_Layout_0.IPD.n409 Folded_Diff_Op_Amp_Layout_0.IPD.n408 0.00773989
R23265 Folded_Diff_Op_Amp_Layout_0.IPD.n433 Folded_Diff_Op_Amp_Layout_0.IPD.n432 0.00773989
R23266 Folded_Diff_Op_Amp_Layout_0.IPD.n385 Folded_Diff_Op_Amp_Layout_0.IPD.n384 0.00773989
R23267 Folded_Diff_Op_Amp_Layout_0.IPD.n234 Folded_Diff_Op_Amp_Layout_0.IPD.n233 0.00642105
R23268 Folded_Diff_Op_Amp_Layout_0.IPD.n247 Folded_Diff_Op_Amp_Layout_0.IPD.n246 0.00642105
R23269 Folded_Diff_Op_Amp_Layout_0.IPD.n380 Folded_Diff_Op_Amp_Layout_0.IPD.n379 0.00605114
R23270 Folded_Diff_Op_Amp_Layout_0.IPD.n355 Folded_Diff_Op_Amp_Layout_0.IPD.n354 0.00605114
R23271 Folded_Diff_Op_Amp_Layout_0.IPD.n242 Folded_Diff_Op_Amp_Layout_0.IPD.n241 0.00605114
R23272 Folded_Diff_Op_Amp_Layout_0.IPD.n84 Folded_Diff_Op_Amp_Layout_0.IPD.n83 0.00605114
R23273 Folded_Diff_Op_Amp_Layout_0.IPD.n425 Folded_Diff_Op_Amp_Layout_0.IPD.n424 0.00605114
R23274 Folded_Diff_Op_Amp_Layout_0.IPD.n360 Folded_Diff_Op_Amp_Layout_0.IPD.n359 0.00570918
R23275 Folded_Diff_Op_Amp_Layout_0.IPD.n246 Folded_Diff_Op_Amp_Layout_0.IPD.n245 0.00551512
R23276 Folded_Diff_Op_Amp_Layout_0.IPD.n438 Folded_Diff_Op_Amp_Layout_0.IPD.n410 0.00549102
R23277 Folded_Diff_Op_Amp_Layout_0.IPD.n434 Folded_Diff_Op_Amp_Layout_0.IPD.n433 0.00549102
R23278 Folded_Diff_Op_Amp_Layout_0.IPD.n348 Folded_Diff_Op_Amp_Layout_0.IPD.n347 0.00523684
R23279 Folded_Diff_Op_Amp_Layout_0.IPD.n361 Folded_Diff_Op_Amp_Layout_0.IPD.n360 0.00523684
R23280 Folded_Diff_Op_Amp_Layout_0.IPD.n374 Folded_Diff_Op_Amp_Layout_0.IPD.n373 0.00523684
R23281 Folded_Diff_Op_Amp_Layout_0.IPD.n88 Folded_Diff_Op_Amp_Layout_0.IPD.n87 0.0051267
R23282 Folded_Diff_Op_Amp_Layout_0.IPD.n368 Folded_Diff_Op_Amp_Layout_0.IPD.n358 0.00479588
R23283 VOUT_OPAMP_N.t19 VOUT_OPAMP_N.t22 147.304
R23284 VOUT_OPAMP_N.t11 VOUT_OPAMP_N.t15 147.304
R23285 VOUT_OPAMP_N.t24 VOUT_OPAMP_N.t14 147.304
R23286 VOUT_OPAMP_N.t20 VOUT_OPAMP_N.t27 147.304
R23287 VOUT_OPAMP_N.n13 VOUT_OPAMP_N.t13 75.2545
R23288 VOUT_OPAMP_N.n24 VOUT_OPAMP_N.t25 75.1498
R23289 VOUT_OPAMP_N.n43 VOUT_OPAMP_N.t24 75.0919
R23290 VOUT_OPAMP_N.n30 VOUT_OPAMP_N.t17 73.4037
R23291 VOUT_OPAMP_N.n49 VOUT_OPAMP_N.t20 73.3458
R23292 VOUT_OPAMP_N.n14 VOUT_OPAMP_N.t30 72.8823
R23293 VOUT_OPAMP_N.n46 VOUT_OPAMP_N.t16 72.3487
R23294 VOUT_OPAMP_N.n44 VOUT_OPAMP_N.t11 72.3487
R23295 VOUT_OPAMP_N.n42 VOUT_OPAMP_N.t10 72.3487
R23296 VOUT_OPAMP_N.n27 VOUT_OPAMP_N.t8 72.3487
R23297 VOUT_OPAMP_N.n25 VOUT_OPAMP_N.t26 72.3487
R23298 VOUT_OPAMP_N.n23 VOUT_OPAMP_N.t12 72.3487
R23299 VOUT_OPAMP_N.n12 VOUT_OPAMP_N.t23 72.3487
R23300 VOUT_OPAMP_N.n46 VOUT_OPAMP_N.t29 51.4916
R23301 VOUT_OPAMP_N.n44 VOUT_OPAMP_N.t19 51.4916
R23302 VOUT_OPAMP_N.n42 VOUT_OPAMP_N.t18 51.4916
R23303 VOUT_OPAMP_N.n27 VOUT_OPAMP_N.t9 51.4916
R23304 VOUT_OPAMP_N.n25 VOUT_OPAMP_N.t7 51.4916
R23305 VOUT_OPAMP_N.n23 VOUT_OPAMP_N.t21 51.4916
R23306 VOUT_OPAMP_N.n12 VOUT_OPAMP_N.t28 51.4916
R23307 VOUT_OPAMP_N.n47 VOUT_OPAMP_N.n46 19.9041
R23308 VOUT_OPAMP_N.n43 VOUT_OPAMP_N.n42 19.9041
R23309 VOUT_OPAMP_N.n28 VOUT_OPAMP_N.n27 19.9041
R23310 VOUT_OPAMP_N.n24 VOUT_OPAMP_N.n23 19.9041
R23311 VOUT_OPAMP_N.n45 VOUT_OPAMP_N.n44 15.6747
R23312 VOUT_OPAMP_N.n26 VOUT_OPAMP_N.n25 15.6747
R23313 VOUT_OPAMP_N.n13 VOUT_OPAMP_N.n12 15.2112
R23314 VOUT_OPAMP_N.n68 VOUT_OPAMP_N.t0 6.52638
R23315 VOUT_OPAMP_N.n70 VOUT_OPAMP_N.t1 6.43144
R23316 VOUT_OPAMP_N.n69 VOUT_OPAMP_N.t3 6.43144
R23317 VOUT_OPAMP_N.n68 VOUT_OPAMP_N.t4 6.43144
R23318 VOUT_OPAMP_N.n71 VOUT_OPAMP_N.t2 3.18927
R23319 VOUT_OPAMP_N.n57 VOUT_OPAMP_N.n38 2.82762
R23320 VOUT_OPAMP_N.n63 VOUT_OPAMP_N.t5 2.73371
R23321 VOUT_OPAMP_N.n63 VOUT_OPAMP_N.t6 2.4088
R23322 VOUT_OPAMP_N.n66 VOUT_OPAMP_N.n65 2.2579
R23323 VOUT_OPAMP_N VOUT_OPAMP_N.n67 1.65759
R23324 VOUT_OPAMP_N.n50 VOUT_OPAMP_N.n49 1.5005
R23325 VOUT_OPAMP_N.n9 VOUT_OPAMP_N.n3 1.49812
R23326 VOUT_OPAMP_N.n9 VOUT_OPAMP_N.n8 1.49812
R23327 VOUT_OPAMP_N.n59 VOUT_OPAMP_N.n21 1.49801
R23328 VOUT_OPAMP_N.n65 VOUT_OPAMP_N.n61 1.4964
R23329 VOUT_OPAMP_N.n64 VOUT_OPAMP_N.n62 1.49069
R23330 VOUT_OPAMP_N.n58 VOUT_OPAMP_N.n57 1.21977
R23331 VOUT_OPAMP_N.n72 VOUT_OPAMP_N.n71 1.19823
R23332 VOUT_OPAMP_N.n67 VOUT_OPAMP_N.n66 1.14993
R23333 VOUT_OPAMP_N.n67 VOUT_OPAMP_N.n61 1.14978
R23334 VOUT_OPAMP_N.n18 VOUT_OPAMP_N.n17 1.14692
R23335 VOUT_OPAMP_N.n60 VOUT_OPAMP_N.n59 1.12675
R23336 VOUT_OPAMP_N.n60 VOUT_OPAMP_N.n9 1.126
R23337 VOUT_OPAMP_N.n16 VOUT_OPAMP_N.n15 1.12272
R23338 VOUT_OPAMP_N.n54 VOUT_OPAMP_N.n53 1.1073
R23339 VOUT_OPAMP_N.n36 VOUT_OPAMP_N.n35 1.1073
R23340 VOUT_OPAMP_N.n57 VOUT_OPAMP_N.n56 0.933295
R23341 VOUT_OPAMP_N.n15 VOUT_OPAMP_N.n13 0.90419
R23342 VOUT_OPAMP_N.n31 VOUT_OPAMP_N.n30 0.897484
R23343 VOUT_OPAMP_N.n45 VOUT_OPAMP_N.n43 0.626587
R23344 VOUT_OPAMP_N.n47 VOUT_OPAMP_N.n45 0.626587
R23345 VOUT_OPAMP_N.n26 VOUT_OPAMP_N.n24 0.626587
R23346 VOUT_OPAMP_N.n28 VOUT_OPAMP_N.n26 0.626587
R23347 VOUT_OPAMP_N VOUT_OPAMP_N.n72 0.391851
R23348 VOUT_OPAMP_N.n20 VOUT_OPAMP_N.n19 0.366019
R23349 VOUT_OPAMP_N.n71 VOUT_OPAMP_N.n70 0.302215
R23350 VOUT_OPAMP_N.n69 VOUT_OPAMP_N.n68 0.289625
R23351 VOUT_OPAMP_N.n72 VOUT_OPAMP_N 0.24757
R23352 VOUT_OPAMP_N.n49 VOUT_OPAMP_N.n47 0.239196
R23353 VOUT_OPAMP_N.n30 VOUT_OPAMP_N.n28 0.239196
R23354 VOUT_OPAMP_N VOUT_OPAMP_N.n60 0.112826
R23355 VOUT_OPAMP_N.n70 VOUT_OPAMP_N.n69 0.069461
R23356 VOUT_OPAMP_N.n35 VOUT_OPAMP_N.n33 0.0649899
R23357 VOUT_OPAMP_N.n53 VOUT_OPAMP_N.n51 0.0638057
R23358 VOUT_OPAMP_N.n64 VOUT_OPAMP_N.n63 0.0608233
R23359 VOUT_OPAMP_N.n53 VOUT_OPAMP_N.n52 0.032498
R23360 VOUT_OPAMP_N.n35 VOUT_OPAMP_N.n34 0.032498
R23361 VOUT_OPAMP_N.n62 VOUT_OPAMP_N.n61 0.0319182
R23362 VOUT_OPAMP_N.n16 VOUT_OPAMP_N.n11 0.0301053
R23363 VOUT_OPAMP_N.n30 VOUT_OPAMP_N.n29 0.0289211
R23364 VOUT_OPAMP_N.n33 VOUT_OPAMP_N.n32 0.0289211
R23365 VOUT_OPAMP_N.n49 VOUT_OPAMP_N.n48 0.0277368
R23366 VOUT_OPAMP_N.n51 VOUT_OPAMP_N.n50 0.0277368
R23367 VOUT_OPAMP_N.n8 VOUT_OPAMP_N.n7 0.0236139
R23368 VOUT_OPAMP_N.n17 VOUT_OPAMP_N.n16 0.0220754
R23369 VOUT_OPAMP_N.n66 VOUT_OPAMP_N.n62 0.0164591
R23370 VOUT_OPAMP_N.n41 VOUT_OPAMP_N.n40 0.0151213
R23371 VOUT_OPAMP_N.n65 VOUT_OPAMP_N.n64 0.0147941
R23372 VOUT_OPAMP_N.n9 VOUT_OPAMP_N.n0 0.014
R23373 VOUT_OPAMP_N.n9 VOUT_OPAMP_N.n5 0.014
R23374 VOUT_OPAMP_N.n59 VOUT_OPAMP_N.n58 0.014
R23375 VOUT_OPAMP_N.n2 VOUT_OPAMP_N.n1 0.014
R23376 VOUT_OPAMP_N.n5 VOUT_OPAMP_N.n4 0.0134654
R23377 VOUT_OPAMP_N.n56 VOUT_OPAMP_N.n55 0.0111023
R23378 VOUT_OPAMP_N.n38 VOUT_OPAMP_N.n37 0.0111023
R23379 VOUT_OPAMP_N.n21 VOUT_OPAMP_N.n20 0.00998204
R23380 VOUT_OPAMP_N.n54 VOUT_OPAMP_N.n39 0.00860784
R23381 VOUT_OPAMP_N.n36 VOUT_OPAMP_N.n22 0.00860784
R23382 VOUT_OPAMP_N.n15 VOUT_OPAMP_N.n14 0.00845754
R23383 VOUT_OPAMP_N.n32 VOUT_OPAMP_N.n31 0.00685938
R23384 VOUT_OPAMP_N.n19 VOUT_OPAMP_N.n18 0.00638348
R23385 VOUT_OPAMP_N.n55 VOUT_OPAMP_N.n54 0.00605114
R23386 VOUT_OPAMP_N.n37 VOUT_OPAMP_N.n36 0.00605114
R23387 VOUT_OPAMP_N.n8 VOUT_OPAMP_N.n6 0.00582347
R23388 VOUT_OPAMP_N.n3 VOUT_OPAMP_N.n2 0.00582347
R23389 VOUT_OPAMP_N.n59 VOUT_OPAMP_N.n10 0.00549102
R23390 VOUT_OPAMP_N.n50 VOUT_OPAMP_N.n41 0.00286842
R23391 Folded_Diff_Op_Amp_Layout_0.IB5.n12 Folded_Diff_Op_Amp_Layout_0.IB5.t0 37.9344
R23392 Folded_Diff_Op_Amp_Layout_0.IB5.n10 Folded_Diff_Op_Amp_Layout_0.IB5.t6 37.9344
R23393 Folded_Diff_Op_Amp_Layout_0.IB5.n12 Folded_Diff_Op_Amp_Layout_0.IB5.t2 17.0773
R23394 Folded_Diff_Op_Amp_Layout_0.IB5.n10 Folded_Diff_Op_Amp_Layout_0.IB5.t4 17.0773
R23395 Folded_Diff_Op_Amp_Layout_0.IB5.n6 Folded_Diff_Op_Amp_Layout_0.IB5.n5 5.57726
R23396 Folded_Diff_Op_Amp_Layout_0.IB5.n11 Folded_Diff_Op_Amp_Layout_0.IB5.n10 4.0005
R23397 Folded_Diff_Op_Amp_Layout_0.IB5.n13 Folded_Diff_Op_Amp_Layout_0.IB5.n12 4.0005
R23398 Folded_Diff_Op_Amp_Layout_0.IB5.n11 Folded_Diff_Op_Amp_Layout_0.IB5.n9 3.58876
R23399 Folded_Diff_Op_Amp_Layout_0.IB5 Folded_Diff_Op_Amp_Layout_0.IB5.n7 2.80542
R23400 Folded_Diff_Op_Amp_Layout_0.IB5 Folded_Diff_Op_Amp_Layout_0.IB5.n22 1.8225
R23401 Folded_Diff_Op_Amp_Layout_0.IB5.n18 Folded_Diff_Op_Amp_Layout_0.IB5.t3 1.6385
R23402 Folded_Diff_Op_Amp_Layout_0.IB5.n18 Folded_Diff_Op_Amp_Layout_0.IB5.n17 1.6385
R23403 Folded_Diff_Op_Amp_Layout_0.IB5.n9 Folded_Diff_Op_Amp_Layout_0.IB5.t7 1.6385
R23404 Folded_Diff_Op_Amp_Layout_0.IB5.n9 Folded_Diff_Op_Amp_Layout_0.IB5.n8 1.6385
R23405 Folded_Diff_Op_Amp_Layout_0.IB5.n2 Folded_Diff_Op_Amp_Layout_0.IB5.n1 1.34776
R23406 Folded_Diff_Op_Amp_Layout_0.IB5.n20 Folded_Diff_Op_Amp_Layout_0.IB5.n19 1.17795
R23407 Folded_Diff_Op_Amp_Layout_0.IB5.n3 Folded_Diff_Op_Amp_Layout_0.IB5.n2 1.14195
R23408 Folded_Diff_Op_Amp_Layout_0.IB5.n16 Folded_Diff_Op_Amp_Layout_0.IB5.n15 1.1255
R23409 Folded_Diff_Op_Amp_Layout_0.IB5.n19 Folded_Diff_Op_Amp_Layout_0.IB5.n18 1.06216
R23410 Folded_Diff_Op_Amp_Layout_0.IB5.n22 Folded_Diff_Op_Amp_Layout_0.IB5.n21 0.631966
R23411 Folded_Diff_Op_Amp_Layout_0.IB5.n5 Folded_Diff_Op_Amp_Layout_0.IB5.t10 0.4555
R23412 Folded_Diff_Op_Amp_Layout_0.IB5.n5 Folded_Diff_Op_Amp_Layout_0.IB5.n4 0.4555
R23413 Folded_Diff_Op_Amp_Layout_0.IB5.n1 Folded_Diff_Op_Amp_Layout_0.IB5.t8 0.4555
R23414 Folded_Diff_Op_Amp_Layout_0.IB5.n1 Folded_Diff_Op_Amp_Layout_0.IB5.n0 0.4555
R23415 Folded_Diff_Op_Amp_Layout_0.IB5.n13 Folded_Diff_Op_Amp_Layout_0.IB5.n11 0.313543
R23416 Folded_Diff_Op_Amp_Layout_0.IB5.n14 Folded_Diff_Op_Amp_Layout_0.IB5.n13 0.281106
R23417 Folded_Diff_Op_Amp_Layout_0.IB5.n7 Folded_Diff_Op_Amp_Layout_0.IB5.n6 0.0929251
R23418 Folded_Diff_Op_Amp_Layout_0.IB5.n21 Folded_Diff_Op_Amp_Layout_0.IB5.n16 0.0712285
R23419 Folded_Diff_Op_Amp_Layout_0.IB5.n21 Folded_Diff_Op_Amp_Layout_0.IB5.n20 0.0534597
R23420 Folded_Diff_Op_Amp_Layout_0.IB5.n15 Folded_Diff_Op_Amp_Layout_0.IB5.n14 0.0407632
R23421 Folded_Diff_Op_Amp_Layout_0.IB5.n7 Folded_Diff_Op_Amp_Layout_0.IB5.n3 0.0320039
R23422 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t47 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t55 95.9434
R23423 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t66 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t47 95.9434
R23424 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t67 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t66 95.9434
R23425 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t42 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t54 95.9434
R23426 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t61 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t42 95.9434
R23427 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t62 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t61 95.9434
R23428 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t33 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t38 95.9434
R23429 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t44 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t33 95.9434
R23430 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t46 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t44 95.9434
R23431 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t80 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t26 95.9434
R23432 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t34 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t80 95.9434
R23433 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t35 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t34 95.9434
R23434 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t75 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t23 95.9434
R23435 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t29 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t75 95.9434
R23436 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t31 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t29 95.9434
R23437 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t51 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t63 95.9434
R23438 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t76 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t51 95.9434
R23439 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t78 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t76 95.9434
R23440 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t49 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t57 95.9434
R23441 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t69 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t49 95.9434
R23442 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t72 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t69 95.9434
R23443 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t41 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t53 95.9434
R23444 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t59 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t41 95.9434
R23445 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t60 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t59 95.9434
R23446 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t32 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t37 95.9434
R23447 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t43 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t32 95.9434
R23448 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t45 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t43 95.9434
R23449 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t27 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t36 95.9434
R23450 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t39 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t27 95.9434
R23451 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t40 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t39 95.9434
R23452 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t74 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t22 95.9434
R23453 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t28 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t74 95.9434
R23454 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t30 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t28 95.9434
R23455 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t65 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t21 95.9434
R23456 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t24 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t65 95.9434
R23457 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t25 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t24 95.9434
R23458 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t48 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t56 95.9434
R23459 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t68 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t48 95.9434
R23460 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t70 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t68 95.9434
R23461 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t52 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t64 95.9434
R23462 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t77 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t52 95.9434
R23463 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t79 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t77 95.9434
R23464 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t10 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t4 95.9434
R23465 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t2 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t10 95.9434
R23466 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t0 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t2 95.9434
R23467 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t14 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t12 95.9434
R23468 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t8 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t14 95.9434
R23469 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t6 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t8 95.9434
R23470 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n50 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t67 65.3674
R23471 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n44 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t6 57.2563
R23472 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n50 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t62 49.1451
R23473 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n51 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t46 49.1451
R23474 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n52 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t35 49.1451
R23475 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n53 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t31 49.1451
R23476 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n54 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t78 49.1451
R23477 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n55 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t72 49.1451
R23478 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n56 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t60 49.1451
R23479 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n57 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t45 49.1451
R23480 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n58 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t40 49.1451
R23481 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n59 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t30 49.1451
R23482 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n60 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t25 49.1451
R23483 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n61 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t70 49.1451
R23484 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n62 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t79 49.1451
R23485 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n63 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t0 49.1451
R23486 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n62 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n63 16.2227
R23487 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n61 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n62 16.2227
R23488 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n60 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n61 16.2227
R23489 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n59 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n58 16.2227
R23490 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n58 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n57 16.2227
R23491 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n57 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n56 16.2227
R23492 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n56 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n55 16.2227
R23493 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n55 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n54 16.2227
R23494 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n54 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n53 16.2227
R23495 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n53 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n52 16.2227
R23496 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n52 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n51 16.2227
R23497 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n51 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n50 16.2227
R23498 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n63 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n44 8.11161
R23499 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t17 5.63646
R23500 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n8 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n7 4.81746
R23501 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n44 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n64 4.80854
R23502 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n43 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n70 4.0405
R23503 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n47 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n60 2.94078
R23504 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n48 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n47 2.8805
R23505 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n46 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n45 2.8805
R23506 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n45 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n59 2.738
R23507 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n67 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n68 2.6005
R23508 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n64 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n65 2.6005
R23509 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n43 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n42 2.6005
R23510 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n24 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n48 1.68759
R23511 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n27 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n26 1.52353
R23512 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n64 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n67 1.4405
R23513 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n67 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n43 1.4405
R23514 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n33 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n32 1.28809
R23515 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n2 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n35 1.14402
R23516 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n34 1.1255
R23517 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n3 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n10 1.1255
R23518 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n41 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n40 1.11801
R23519 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n15 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n11 1.11801
R23520 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n38 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n37 1.11782
R23521 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n29 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n28 1.11782
R23522 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n26 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n25 1.11782
R23523 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n32 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t18 0.8195
R23524 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n32 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n31 0.8195
R23525 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n7 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t19 0.8195
R23526 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n7 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n6 0.8195
R23527 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n65 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t7 0.607167
R23528 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n65 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n66 0.607167
R23529 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n68 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t9 0.607167
R23530 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n68 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n69 0.607167
R23531 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n70 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t13 0.607167
R23532 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n70 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n71 0.607167
R23533 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n42 Folded_Diff_Op_Amp_Layout_0.IBIAS3.t15 0.607167
R23534 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n42 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n72 0.607167
R23535 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n37 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n2 0.576345
R23536 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n9 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n8 0.211804
R23537 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n3 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n29 0.209193
R23538 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n10 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n9 0.121804
R23539 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n41 0.0917676
R23540 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n48 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n49 0.0834892
R23541 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n34 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n33 0.061035
R23542 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n49 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n46 0.0416511
R23543 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n2 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n1 0.0249014
R23544 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n20 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n19 0.0228651
R23545 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n22 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n21 0.0228651
R23546 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n40 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n39 0.0179841
R23547 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n14 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n13 0.0179841
R23548 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n29 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n15 0.0179841
R23549 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n19 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n18 0.0179841
R23550 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n5 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n4 0.0177304
R23551 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n15 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n14 0.0177304
R23552 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n13 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n12 0.0177304
R23553 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n18 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n17 0.0177304
R23554 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n1 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n0 0.0176127
R23555 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n38 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n5 0.0173591
R23556 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n37 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n36 0.0173591
R23557 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n41 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n38 0.0173591
R23558 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n28 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n16 0.0173591
R23559 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n28 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n27 0.0173591
R23560 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n25 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n23 0.0173591
R23561 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n25 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n24 0.0173591
R23562 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n0 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n30 0.0163451
R23563 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n26 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n20 0.0119325
R23564 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n23 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n22 0.0119325
R23565 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n30 Folded_Diff_Op_Amp_Layout_0.IBIAS3.n3 0.0105038
R23566 a_29734_3659.n4 a_29734_3659.n0 2.11607
R23567 a_29734_3659.n1 a_29734_3659.n2 0.3755
R23568 a_29734_3659.n0 a_29734_3659.n5 0.00704942
R23569 a_29734_3659.t0 a_29734_3659.n4 2.4095
R23570 a_29734_3659.n11 a_29734_3659.n12 0.2255
R23571 a_29734_3659.n2 a_29734_3659.n13 0.2255
R23572 a_29734_3659.n14 a_29734_3659.n15 0.2255
R23573 a_29734_3659.n18 a_29734_3659.n14 0.00133482
R23574 a_29734_3659.n52 a_29734_3659.n53 1.4369
R23575 a_29734_3659.n8 a_29734_3659.n7 0.00183414
R23576 a_29734_3659.n52 a_29734_3659.n48 0.011643
R23577 a_29734_3659.n49 a_29734_3659.n8 0.00104878
R23578 a_29734_3659.n21 a_29734_3659.n49 0.00489024
R23579 a_29734_3659.n25 a_29734_3659.n21 0.00964634
R23580 a_29734_3659.n9 a_29734_3659.n25 0.00543902
R23581 a_29734_3659.n23 a_29734_3659.n9 0.00543902
R23582 a_29734_3659.n29 a_29734_3659.n23 0.00964634
R23583 a_29734_3659.n11 a_29734_3659.n29 0.00543902
R23584 a_29734_3659.n27 a_29734_3659.n11 0.00543902
R23585 a_29734_3659.n34 a_29734_3659.n27 0.00964634
R23586 a_29734_3659.n2 a_29734_3659.n34 0.00543902
R23587 a_29734_3659.n2 a_29734_3659.n16 0.00543902
R23588 a_29734_3659.n55 a_29734_3659.n32 0.00470732
R23589 a_29734_3659.n14 a_29734_3659.n55 0.00123171
R23590 a_29734_3659.n51 a_29734_3659.t3 6.46072
R23591 a_29734_3659.n6 a_29734_3659.n51 0.0350732
R23592 a_29734_3659.n50 a_29734_3659.n6 0.00470732
R23593 a_29734_3659.n48 a_29734_3659.n50 0.00104878
R23594 a_29734_3659.n19 a_29734_3659.n52 0.0107893
R23595 a_29734_3659.n54 a_29734_3659.n19 0.00745122
R23596 a_29734_3659.n20 a_29734_3659.n54 0.0125732
R23597 a_29734_3659.n3 a_29734_3659.n20 0.0174535
R23598 a_29734_3659.n1 a_29734_3659.n3 0.00356683
R23599 a_29734_3659.n0 a_29734_3659.n1 0.0142296
R23600 a_29734_3659.n5 a_29734_3659.n18 0.376453
R23601 a_29734_3659.n53 a_29734_3659.t2 2.4095
R23602 a_29734_3659.n51 a_29734_3659.t1 6.4095
R23603 a_29734_3659.n39 a_29734_3659.n37 0.0102304
R23604 a_29734_3659.n43 a_29734_3659.n45 0.0101264
R23605 a_29734_3659.n7 a_29734_3659.n22 0.185497
R23606 a_29734_3659.n22 a_29734_3659.n26 0.00964634
R23607 a_29734_3659.n26 a_29734_3659.n10 0.00543902
R23608 a_29734_3659.n10 a_29734_3659.n24 0.00543902
R23609 a_29734_3659.n12 a_29734_3659.n30 0.00543902
R23610 a_29734_3659.n35 a_29734_3659.n28 0.00964634
R23611 a_29734_3659.n13 a_29734_3659.n35 0.00543902
R23612 a_29734_3659.n13 a_29734_3659.n17 0.00543902
R23613 a_29734_3659.n15 a_29734_3659.n33 0.00543902
R23614 a_29734_3659.n15 a_29734_3659.n31 0.00543902
R23615 a_29734_3659.n31 a_29734_3659.n36 0.246171
R23616 a_29734_3659.n36 a_29734_3659.n38 0.0195244
R23617 a_29734_3659.n38 a_29734_3659.n40 0.0195244
R23618 a_29734_3659.n40 a_29734_3659.n43 0.245024
R23619 a_29734_3659.n41 a_29734_3659.n39 0.0195244
R23620 a_29734_3659.n45 a_29734_3659.n41 0.0195244
R23621 a_29734_3659.n37 a_29734_3659.n42 0.231891
R23622 a_29734_3659.n42 a_29734_3659.n44 0.00895528
R23623 a_29734_3659.n44 a_29734_3659.n46 0.00895528
R23624 a_29734_3659.n47 a_29734_3659.t4 2.2505
R23625 a_29734_3659.n46 a_29734_3659.n47 0.105743
R23626 a_29734_3659.n47 a_29734_3659.t5 2.38861
R23627 a_n5986_9350.t0 a_n5986_9350.t1 14.4367
R23628 VIN_P1 VIN_P1.t0 5.25526
R23629 a_n7106_6102.t0 a_n7106_6102.t1 14.32
R23630 Folded_Diff_Op_Amp_Layout_0.VB3.n61 Folded_Diff_Op_Amp_Layout_0.VB3.t43 51.5034
R23631 Folded_Diff_Op_Amp_Layout_0.VB3.n60 Folded_Diff_Op_Amp_Layout_0.VB3.t20 50.3184
R23632 Folded_Diff_Op_Amp_Layout_0.VB3.n59 Folded_Diff_Op_Amp_Layout_0.VB3.t33 50.3184
R23633 Folded_Diff_Op_Amp_Layout_0.VB3.n58 Folded_Diff_Op_Amp_Layout_0.VB3.t24 50.3184
R23634 Folded_Diff_Op_Amp_Layout_0.VB3.n57 Folded_Diff_Op_Amp_Layout_0.VB3.t38 50.3184
R23635 Folded_Diff_Op_Amp_Layout_0.VB3.n56 Folded_Diff_Op_Amp_Layout_0.VB3.t22 50.3184
R23636 Folded_Diff_Op_Amp_Layout_0.VB3.n55 Folded_Diff_Op_Amp_Layout_0.VB3.t34 50.3184
R23637 Folded_Diff_Op_Amp_Layout_0.VB3.n54 Folded_Diff_Op_Amp_Layout_0.VB3.t41 50.3184
R23638 Folded_Diff_Op_Amp_Layout_0.VB3.n47 Folded_Diff_Op_Amp_Layout_0.VB3.t44 50.3184
R23639 Folded_Diff_Op_Amp_Layout_0.VB3.n39 Folded_Diff_Op_Amp_Layout_0.VB3.t29 50.3184
R23640 Folded_Diff_Op_Amp_Layout_0.VB3.n38 Folded_Diff_Op_Amp_Layout_0.VB3.t21 50.3184
R23641 Folded_Diff_Op_Amp_Layout_0.VB3.n43 Folded_Diff_Op_Amp_Layout_0.VB3.t16 50.3184
R23642 Folded_Diff_Op_Amp_Layout_0.VB3.n42 Folded_Diff_Op_Amp_Layout_0.VB3.t52 50.3184
R23643 Folded_Diff_Op_Amp_Layout_0.VB3.n44 Folded_Diff_Op_Amp_Layout_0.VB3.t26 50.3184
R23644 Folded_Diff_Op_Amp_Layout_0.VB3.n41 Folded_Diff_Op_Amp_Layout_0.VB3.t19 50.3184
R23645 Folded_Diff_Op_Amp_Layout_0.VB3.n45 Folded_Diff_Op_Amp_Layout_0.VB3.t18 50.3184
R23646 Folded_Diff_Op_Amp_Layout_0.VB3.n40 Folded_Diff_Op_Amp_Layout_0.VB3.t36 50.3184
R23647 Folded_Diff_Op_Amp_Layout_0.VB3.n50 Folded_Diff_Op_Amp_Layout_0.VB3.t31 50.3184
R23648 Folded_Diff_Op_Amp_Layout_0.VB3.n49 Folded_Diff_Op_Amp_Layout_0.VB3.t46 50.3184
R23649 Folded_Diff_Op_Amp_Layout_0.VB3.n53 Folded_Diff_Op_Amp_Layout_0.VB3.t17 50.3184
R23650 Folded_Diff_Op_Amp_Layout_0.VB3.n48 Folded_Diff_Op_Amp_Layout_0.VB3.t35 50.3184
R23651 Folded_Diff_Op_Amp_Layout_0.VB3.n51 Folded_Diff_Op_Amp_Layout_0.VB3.t39 50.3184
R23652 Folded_Diff_Op_Amp_Layout_0.VB3.n46 Folded_Diff_Op_Amp_Layout_0.VB3.t51 50.3184
R23653 Folded_Diff_Op_Amp_Layout_0.VB3.n52 Folded_Diff_Op_Amp_Layout_0.VB3.t28 50.3184
R23654 Folded_Diff_Op_Amp_Layout_0.VB3.n61 Folded_Diff_Op_Amp_Layout_0.VB3.t37 48.2728
R23655 Folded_Diff_Op_Amp_Layout_0.VB3.t43 Folded_Diff_Op_Amp_Layout_0.VB3.n39 46.4076
R23656 Folded_Diff_Op_Amp_Layout_0.VB3.n60 Folded_Diff_Op_Amp_Layout_0.VB3.t25 46.4076
R23657 Folded_Diff_Op_Amp_Layout_0.VB3.t25 Folded_Diff_Op_Amp_Layout_0.VB3.n43 46.4076
R23658 Folded_Diff_Op_Amp_Layout_0.VB3.n59 Folded_Diff_Op_Amp_Layout_0.VB3.t40 46.4076
R23659 Folded_Diff_Op_Amp_Layout_0.VB3.t40 Folded_Diff_Op_Amp_Layout_0.VB3.n44 46.4076
R23660 Folded_Diff_Op_Amp_Layout_0.VB3.n58 Folded_Diff_Op_Amp_Layout_0.VB3.t30 46.4076
R23661 Folded_Diff_Op_Amp_Layout_0.VB3.t30 Folded_Diff_Op_Amp_Layout_0.VB3.n45 46.4076
R23662 Folded_Diff_Op_Amp_Layout_0.VB3.n57 Folded_Diff_Op_Amp_Layout_0.VB3.t45 46.4076
R23663 Folded_Diff_Op_Amp_Layout_0.VB3.t45 Folded_Diff_Op_Amp_Layout_0.VB3.n50 46.4076
R23664 Folded_Diff_Op_Amp_Layout_0.VB3.n56 Folded_Diff_Op_Amp_Layout_0.VB3.t27 46.4076
R23665 Folded_Diff_Op_Amp_Layout_0.VB3.t27 Folded_Diff_Op_Amp_Layout_0.VB3.n53 46.4076
R23666 Folded_Diff_Op_Amp_Layout_0.VB3.n55 Folded_Diff_Op_Amp_Layout_0.VB3.t42 46.4076
R23667 Folded_Diff_Op_Amp_Layout_0.VB3.t29 Folded_Diff_Op_Amp_Layout_0.VB3.n38 46.4076
R23668 Folded_Diff_Op_Amp_Layout_0.VB3.t16 Folded_Diff_Op_Amp_Layout_0.VB3.n42 46.4076
R23669 Folded_Diff_Op_Amp_Layout_0.VB3.t31 Folded_Diff_Op_Amp_Layout_0.VB3.n49 46.4076
R23670 Folded_Diff_Op_Amp_Layout_0.VB3.n54 Folded_Diff_Op_Amp_Layout_0.VB3.t49 46.4076
R23671 Folded_Diff_Op_Amp_Layout_0.VB3.n34 Folded_Diff_Op_Amp_Layout_0.VB3.t8 20.6621
R23672 Folded_Diff_Op_Amp_Layout_0.VB3.n17 Folded_Diff_Op_Amp_Layout_0.VB3.t48 20.0755
R23673 Folded_Diff_Op_Amp_Layout_0.VB3.n61 Folded_Diff_Op_Amp_Layout_0.VB3.n60 18.9805
R23674 Folded_Diff_Op_Amp_Layout_0.VB3.n41 Folded_Diff_Op_Amp_Layout_0.VB3.n40 17.5205
R23675 Folded_Diff_Op_Amp_Layout_0.VB3.n49 Folded_Diff_Op_Amp_Layout_0.VB3.n48 17.5205
R23676 Folded_Diff_Op_Amp_Layout_0.VB3.n47 Folded_Diff_Op_Amp_Layout_0.VB3.n46 17.5205
R23677 Folded_Diff_Op_Amp_Layout_0.VB3.n52 Folded_Diff_Op_Amp_Layout_0.VB3.n51 17.5205
R23678 Folded_Diff_Op_Amp_Layout_0.VB3.n59 Folded_Diff_Op_Amp_Layout_0.VB3.n58 17.5205
R23679 Folded_Diff_Op_Amp_Layout_0.VB3.n57 Folded_Diff_Op_Amp_Layout_0.VB3.n56 17.5205
R23680 Folded_Diff_Op_Amp_Layout_0.VB3.n55 Folded_Diff_Op_Amp_Layout_0.VB3.n54 17.5205
R23681 Folded_Diff_Op_Amp_Layout_0.VB3.n17 Folded_Diff_Op_Amp_Layout_0.VB3.t10 15.6434
R23682 Folded_Diff_Op_Amp_Layout_0.VB3.n20 Folded_Diff_Op_Amp_Layout_0.VB3.t4 15.6434
R23683 Folded_Diff_Op_Amp_Layout_0.VB3.n23 Folded_Diff_Op_Amp_Layout_0.VB3.t12 15.6434
R23684 Folded_Diff_Op_Amp_Layout_0.VB3.n26 Folded_Diff_Op_Amp_Layout_0.VB3.t2 15.6434
R23685 Folded_Diff_Op_Amp_Layout_0.VB3.n30 Folded_Diff_Op_Amp_Layout_0.VB3.t0 15.6434
R23686 Folded_Diff_Op_Amp_Layout_0.VB3.n36 Folded_Diff_Op_Amp_Layout_0.VB3.t6 15.6434
R23687 Folded_Diff_Op_Amp_Layout_0.VB3.n42 Folded_Diff_Op_Amp_Layout_0.VB3.n41 9.73383
R23688 Folded_Diff_Op_Amp_Layout_0.VB3.n48 Folded_Diff_Op_Amp_Layout_0.VB3.n47 9.73383
R23689 Folded_Diff_Op_Amp_Layout_0.VB3.n53 Folded_Diff_Op_Amp_Layout_0.VB3.n52 9.73383
R23690 Folded_Diff_Op_Amp_Layout_0.VB3.n60 Folded_Diff_Op_Amp_Layout_0.VB3.n59 9.73383
R23691 Folded_Diff_Op_Amp_Layout_0.VB3.n58 Folded_Diff_Op_Amp_Layout_0.VB3.n57 9.73383
R23692 Folded_Diff_Op_Amp_Layout_0.VB3.n56 Folded_Diff_Op_Amp_Layout_0.VB3.n55 9.73383
R23693 Folded_Diff_Op_Amp_Layout_0.VB3.n2 Folded_Diff_Op_Amp_Layout_0.VB3.n10 7.46311
R23694 Folded_Diff_Op_Amp_Layout_0.VB3.n1 Folded_Diff_Op_Amp_Layout_0.VB3.n33 5.31813
R23695 Folded_Diff_Op_Amp_Layout_0.VB3.n27 Folded_Diff_Op_Amp_Layout_0.VB3.n26 5.21479
R23696 Folded_Diff_Op_Amp_Layout_0.VB3.n24 Folded_Diff_Op_Amp_Layout_0.VB3.n23 5.21479
R23697 Folded_Diff_Op_Amp_Layout_0.VB3.n21 Folded_Diff_Op_Amp_Layout_0.VB3.n20 5.21479
R23698 Folded_Diff_Op_Amp_Layout_0.VB3.n18 Folded_Diff_Op_Amp_Layout_0.VB3.n17 5.21479
R23699 Folded_Diff_Op_Amp_Layout_0.VB3.n1 Folded_Diff_Op_Amp_Layout_0.VB3.n37 4.5005
R23700 Folded_Diff_Op_Amp_Layout_0.VB3.n31 Folded_Diff_Op_Amp_Layout_0.VB3.n30 4.04157
R23701 Folded_Diff_Op_Amp_Layout_0.VB3.n28 Folded_Diff_Op_Amp_Layout_0.VB3.n27 4.0005
R23702 Folded_Diff_Op_Amp_Layout_0.VB3.n25 Folded_Diff_Op_Amp_Layout_0.VB3.n24 4.0005
R23703 Folded_Diff_Op_Amp_Layout_0.VB3.n22 Folded_Diff_Op_Amp_Layout_0.VB3.n21 4.0005
R23704 Folded_Diff_Op_Amp_Layout_0.VB3.n19 Folded_Diff_Op_Amp_Layout_0.VB3.n18 4.0005
R23705 Folded_Diff_Op_Amp_Layout_0.VB3.n1 Folded_Diff_Op_Amp_Layout_0.VB3.n35 4.0005
R23706 Folded_Diff_Op_Amp_Layout_0.VB3.n4 Folded_Diff_Op_Amp_Layout_0.VB3.n32 4.0005
R23707 Folded_Diff_Op_Amp_Layout_0.VB3.n37 Folded_Diff_Op_Amp_Layout_0.VB3.n36 3.91121
R23708 Folded_Diff_Op_Amp_Layout_0.VB3.n4 Folded_Diff_Op_Amp_Layout_0.VB3.n12 3.43224
R23709 Folded_Diff_Op_Amp_Layout_0.VB3.n19 Folded_Diff_Op_Amp_Layout_0.VB3.n16 3.43224
R23710 Folded_Diff_Op_Amp_Layout_0.VB3.n25 Folded_Diff_Op_Amp_Layout_0.VB3.n14 3.43224
R23711 Folded_Diff_Op_Amp_Layout_0.VB3.n62 Folded_Diff_Op_Amp_Layout_0.VB3.n61 11.085
R23712 Folded_Diff_Op_Amp_Layout_0.VB3.n2 Folded_Diff_Op_Amp_Layout_0.VB3.n4 1.695
R23713 Folded_Diff_Op_Amp_Layout_0.VB3.n3 Folded_Diff_Op_Amp_Layout_0.VB3.n1 1.688
R23714 Folded_Diff_Op_Amp_Layout_0.VB3.n12 Folded_Diff_Op_Amp_Layout_0.VB3.t7 1.6385
R23715 Folded_Diff_Op_Amp_Layout_0.VB3.n12 Folded_Diff_Op_Amp_Layout_0.VB3.n11 1.6385
R23716 Folded_Diff_Op_Amp_Layout_0.VB3.n16 Folded_Diff_Op_Amp_Layout_0.VB3.t5 1.6385
R23717 Folded_Diff_Op_Amp_Layout_0.VB3.n16 Folded_Diff_Op_Amp_Layout_0.VB3.n15 1.6385
R23718 Folded_Diff_Op_Amp_Layout_0.VB3.n14 Folded_Diff_Op_Amp_Layout_0.VB3.t3 1.6385
R23719 Folded_Diff_Op_Amp_Layout_0.VB3.n14 Folded_Diff_Op_Amp_Layout_0.VB3.n13 1.6385
R23720 Folded_Diff_Op_Amp_Layout_0.VB3.n10 Folded_Diff_Op_Amp_Layout_0.VB3.n7 1.19119
R23721 Folded_Diff_Op_Amp_Layout_0.VB3.n32 Folded_Diff_Op_Amp_Layout_0.VB3.n31 1.17371
R23722 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VB3.n62 1.05764
R23723 Folded_Diff_Op_Amp_Layout_0.VB3.n7 Folded_Diff_Op_Amp_Layout_0.VB3.n6 0.813264
R23724 Folded_Diff_Op_Amp_Layout_0.VB3.n62 Folded_Diff_Op_Amp_Layout_0.VB3.n3 0.806689
R23725 Folded_Diff_Op_Amp_Layout_0.VB3.n6 Folded_Diff_Op_Amp_Layout_0.VB3.t14 0.4555
R23726 Folded_Diff_Op_Amp_Layout_0.VB3.n6 Folded_Diff_Op_Amp_Layout_0.VB3.n5 0.4555
R23727 Folded_Diff_Op_Amp_Layout_0.VB3.n32 Folded_Diff_Op_Amp_Layout_0.VB3.n29 0.326393
R23728 Folded_Diff_Op_Amp_Layout_0.VB3.n28 Folded_Diff_Op_Amp_Layout_0.VB3.n25 0.253132
R23729 Folded_Diff_Op_Amp_Layout_0.VB3.n25 Folded_Diff_Op_Amp_Layout_0.VB3.n22 0.253132
R23730 Folded_Diff_Op_Amp_Layout_0.VB3.n22 Folded_Diff_Op_Amp_Layout_0.VB3.n19 0.253132
R23731 Folded_Diff_Op_Amp_Layout_0.VB3.n4 Folded_Diff_Op_Amp_Layout_0.VB3.n28 0.227237
R23732 Folded_Diff_Op_Amp_Layout_0.VB3.n35 Folded_Diff_Op_Amp_Layout_0.VB3.n34 0.196036
R23733 Folded_Diff_Op_Amp_Layout_0.VB3.n1 Folded_Diff_Op_Amp_Layout_0.VB3.n0 0.0740526
R23734 Folded_Diff_Op_Amp_Layout_0.VB3.n3 Folded_Diff_Op_Amp_Layout_0.VB3.n2 0.066
R23735 Folded_Diff_Op_Amp_Layout_0.VB3.n10 Folded_Diff_Op_Amp_Layout_0.VB3.n9 0.0623855
R23736 Folded_Diff_Op_Amp_Layout_0.VB3.n9 Folded_Diff_Op_Amp_Layout_0.VB3.n8 0.0623855
R23737 a_24556_2845.t0 a_24556_2845.t1 13.3663
R23738 a_24836_1743.t0 a_24836_1743.t1 13.4632
R23739 a_n6826_9350.t0 a_n6826_9350.t1 13.5425
R23740 a_n7106_8433.n0 a_n7106_8433.t0 7.26507
R23741 a_n7106_8433.n4 a_n7106_8433.t1 3.89298
R23742 a_n7106_8433.t3 a_n7106_8433.n5 3.06722
R23743 a_n7106_8433.n4 a_n7106_8433.n0 2.47036
R23744 a_n7106_8433.n3 a_n7106_8433.t2 2.3
R23745 a_n7106_8433.t4 a_n7106_8433.n1 1.1255
R23746 a_n7106_8433.t4 a_n7106_8433.n2 1.1255
R23747 a_n7106_8433.t4 a_n7106_8433.n4 2.42357
R23748 a_n7106_8433.n0 a_n7106_8433.n3 1.75717
R23749 a_n7106_8433.n5 a_n7106_8433.t4 0.607547
R23750 a_n6546_6102.t0 a_n6546_6102.t1 14.6442
R23751 a_n5426_5540.t0 a_n5426_5540.t1 8.92051
R23752 a_26292_4817.t0 a_26292_4817.t1 13.4632
R23753 a_26740_4817.t0 a_26740_4817.t1 13.3663
R23754 a_27020_3715.t0 a_27020_3715.t1 11.9264
R23755 a_n6266_10267.t0 a_n6266_10267.t1 13.5444
R23756 a_n5706_9705.t0 a_n5706_9705.t1 13.5425
R23757 a_n7106_8788.t0 a_n7106_8788.t1 14.32
R23758 a_n5146_6102.t0 a_n5146_6102.t1 13.5425
R23759 a_n4866_5185.t0 a_n4866_5185.t1 10.1673
R23760 a_n5426_9350.t0 a_n5426_9350.t1 8.88572
R23761 a_n6546_8788.t0 a_n6546_8788.t1 14.6442
R23762 a_24108_2845.t0 a_24108_2845.t1 13.4632
R23763 Folded_Diff_Op_Amp_Layout_0.IB3.n9 Folded_Diff_Op_Amp_Layout_0.IB3.n8 4.05833
R23764 Folded_Diff_Op_Amp_Layout_0.IB3.n4 Folded_Diff_Op_Amp_Layout_0.IB3.n3 4.05833
R23765 Folded_Diff_Op_Amp_Layout_0.IB3.n4 Folded_Diff_Op_Amp_Layout_0.IB3.n1 3.43224
R23766 Folded_Diff_Op_Amp_Layout_0.IB3.n9 Folded_Diff_Op_Amp_Layout_0.IB3.n6 3.43224
R23767 Folded_Diff_Op_Amp_Layout_0.IB3.n1 Folded_Diff_Op_Amp_Layout_0.IB3.t5 1.6385
R23768 Folded_Diff_Op_Amp_Layout_0.IB3.n1 Folded_Diff_Op_Amp_Layout_0.IB3.n0 1.6385
R23769 Folded_Diff_Op_Amp_Layout_0.IB3.n6 Folded_Diff_Op_Amp_Layout_0.IB3.t4 1.6385
R23770 Folded_Diff_Op_Amp_Layout_0.IB3.n6 Folded_Diff_Op_Amp_Layout_0.IB3.n5 1.6385
R23771 Folded_Diff_Op_Amp_Layout_0.IB3.n8 Folded_Diff_Op_Amp_Layout_0.IB3.t1 1.6385
R23772 Folded_Diff_Op_Amp_Layout_0.IB3.n8 Folded_Diff_Op_Amp_Layout_0.IB3.n7 1.6385
R23773 Folded_Diff_Op_Amp_Layout_0.IB3.n3 Folded_Diff_Op_Amp_Layout_0.IB3.t0 1.6385
R23774 Folded_Diff_Op_Amp_Layout_0.IB3.n3 Folded_Diff_Op_Amp_Layout_0.IB3.n2 1.6385
R23775 Folded_Diff_Op_Amp_Layout_0.IB3 Folded_Diff_Op_Amp_Layout_0.IB3.n4 0.313543
R23776 Folded_Diff_Op_Amp_Layout_0.IB3 Folded_Diff_Op_Amp_Layout_0.IB3.n9 0.313543
R23777 a_n5426_10267.t0 a_n5426_10267.t1 13.5425
R23778 a_n4866_9705.t0 a_n4866_9705.t1 10.1324
R23779 a_n7106_9350.t2 a_n7106_9350.t3 5.9203
R23780 a_n7106_9350.t2 a_n7106_9350.t1 4.57473
R23781 a_n7106_9350.t0 a_n7106_9350.t2 3.89251
R23782 a_n6826_9705.t0 a_n6826_9705.t1 13.5425
R23783 a_n5146_8788.t0 a_n5146_8788.t1 13.5425
R23784 a_n5706_5540.t0 a_n5706_5540.t1 13.5425
R23785 filter_res_magic_0.R3_R7.t6 filter_res_magic_0.R3_R7.t7 5.14152
R23786 filter_res_magic_0.R3_R7.n2 filter_res_magic_0.R3_R7.t0 4.72867
R23787 filter_res_magic_0.R3_R7.n2 filter_res_magic_0.R3_R7.t1 3.99183
R23788 filter_res_magic_0.R3_R7.t3 filter_res_magic_0.R3_R7.n6 2.88446
R23789 filter_res_magic_0.R3_R7.n0 filter_res_magic_0.R3_R7.t5 2.27001
R23790 filter_res_magic_0.R3_R7.n6 filter_res_magic_0.R3_R7.t4 2.25756
R23791 filter_res_magic_0.R3_R7.n5 filter_res_magic_0.R3_R7.t2 2.25756
R23792 filter_res_magic_0.R3_R7.n4 filter_res_magic_0.R3_R7.n3 1.77718
R23793 filter_res_magic_0.R3_R7.n6 filter_res_magic_0.R3_R7.n5 1.44088
R23794 filter_res_magic_0.R3_R7.n4 filter_res_magic_0.R3_R7.n1 1.14805
R23795 filter_res_magic_0.R3_R7.n0 filter_res_magic_0.R3_R7.n4 0.6705
R23796 filter_res_magic_0.R3_R7.t6 filter_res_magic_0.R3_R7.t3 0.663092
R23797 filter_res_magic_0.R3_R7.n5 filter_res_magic_0.R3_R7.n0 0.582009
R23798 filter_res_magic_0.R3_R7 filter_res_magic_0.R3_R7.n2 0.299466
R23799 filter_res_magic_0.R3_R7.n3 filter_res_magic_0.R3_R7 0.152486
R23800 a_n6546_10267.t0 a_n6546_10267.t1 13.5425
R23801 a_n5986_9705.t0 a_n5986_9705.t1 13.5425
R23802 a_n6266_6102.t0 a_n6266_6102.t1 13.5425
R23803 a_n5986_7019.t0 a_n5986_7019.t1 12.9821
R23804 a_n5706_6457.t0 a_n5706_6457.t1 12.9821
R23805 a_n5146_10267.t0 a_n5146_10267.t1 13.5444
R23806 a_n5706_5185.t0 a_n5706_5185.t1 13.5425
R23807 a_n6266_4623.t0 a_n6266_4623.t1 13.5444
R23808 a_n7106_9705.t0 a_n7106_9705.t1 13.5444
R23809 a_25564_2845.t0 a_25564_2845.t1 13.4632
R23810 a_25284_1743.t0 a_25284_1743.t1 13.3663
R23811 a_n7106_7019.t0 a_n7106_7019.t1 12.9821
R23812 a_n6826_6457.t0 a_n6826_6457.t1 12.9821
R23813 a_n5426_4623.t0 a_n5426_4623.t1 13.5425
R23814 a_26292_1743.t0 a_26292_1743.t1 13.4632
R23815 a_n5706_8433.t0 a_n5706_8433.t1 12.9667
R23816 a_n5986_7871.t0 a_n5986_7871.t1 13.0109
R23817 a_26740_1743.t0 a_26740_1743.t1 13.3663
R23818 a_n6826_5185.t0 a_n6826_5185.t1 13.5425
R23819 a_n6266_6457.t0 a_n6266_6457.t1 12.9821
R23820 a_n5426_7019.t0 a_n5426_7019.t1 12.9821
R23821 a_n5986_5185.t0 a_n5986_5185.t1 13.5425
R23822 a_n6546_4623.t0 a_n6546_4623.t1 13.5425
R23823 a_n6826_8433.t0 a_n6826_8433.t1 12.9821
R23824 a_n7106_7871.t0 a_n7106_7871.t1 12.9821
R23825 a_26012_2845.t0 a_26012_2845.t1 13.3663
R23826 a_n6546_7019.t0 a_n6546_7019.t1 12.9821
R23827 a_n6266_8433.t0 a_n6266_8433.t1 12.98
R23828 a_n5146_4623.t0 a_n5146_4623.t1 13.5444
R23829 a_n5426_7871.t0 a_n5426_7871.t1 12.9667
R23830 a_n7106_5185.t0 a_n7106_5185.t1 13.5444
R23831 a_n6546_7871.t0 a_n6546_7871.t1 12.9821
R23832 a_27020_2845.t0 a_27020_2845.t1 13.3199
R23833 a_24556_3715.t0 a_24556_3715.t1 13.3663
R23834 a_25564_3715.t0 a_25564_3715.t1 13.4632
C0 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB4 1.68f
C1 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.OUT2 0.655f
C2 VOUT_OPAMP_N VOUT_OPAMP_P 3.52f
C3 VOUT_OPAMP_P VIN_P1 0.0407f
C4 Folded_Diff_Op_Amp_Layout_0.IND VOUT_P 0.00521f
C5 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.IB5 0.178f
C6 Folded_Diff_Op_Amp_Layout_0.OUT1 VCM1 0.00957f
C7 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IBIAS 0.95f
C8 Folded_Diff_Op_Amp_Layout_0.IBIAS3 VDD 9.66f
C9 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VND 0.998f
C10 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB1 0.656f
C11 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VPD 5.35f
C12 Folded_Diff_Op_Amp_Layout_0.IB3 VCM1 6.71e-19
C13 Folded_Diff_Op_Amp_Layout_0.IBIAS VCM1 0.935f
C14 VDD VIN_N1 0.667f
C15 Folded_Diff_Op_Amp_Layout_0.IBS Folded_Diff_Op_Amp_Layout_0.IB5 0.854f
C16 Folded_Diff_Op_Amp_Layout_0.IBIAS1 Folded_Diff_Op_Amp_Layout_0.VBIASN 0.559f
C17 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IVS 1.2f
C18 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.VB1 1.84f
C19 Folded_Diff_Op_Amp_Layout_0.VOUT VDD 2.29f
C20 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.BD 9.48f
C21 filter_res_magic_0.R7_R8_R10_C VDD 1.03f
C22 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.OUT1 0.00709f
C23 filter_res_magic_0.R7_R8_R10_C VOUT_N 0.00657f
C24 Folded_Diff_Op_Amp_Layout_0.IBS VCM1 0.124f
C25 Folded_Diff_Op_Amp_Layout_0.IND VCM1 8.4e-20
C26 filter_res_magic_0.R3_R7 VDD 0.931f
C27 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.VCD 0.929f
C28 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.IBIAS4 0.0154f
C29 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.IBS 0.292f
C30 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.VB4 0.185f
C31 Folded_Diff_Op_Amp_Layout_0.OUT2 VDD 12.2f
C32 Folded_Diff_Op_Amp_Layout_0.OUT2 VOUT_N 7.55f
C33 VOUT_OPAMP_N VIN_N1 0.0413f
C34 VDD VOUT_P 87.9f
C35 VOUT_N VOUT_P 0.112p
C36 Folded_Diff_Op_Amp_Layout_0.IB4 VDD 2.94f
C37 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VBM 0.00633f
C38 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VOUT 0.594f
C39 Folded_Diff_Op_Amp_Layout_0.VPD Folded_Diff_Op_Amp_Layout_0.VB1 0.946f
C40 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.IBS 0.029f
C41 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB4 1.39f
C42 filter_res_magic_0.R7_R8_R10_C VOUT_OPAMP_N 6.07e-19
C43 filter_res_magic_0.R7_R8_R10_C VIN_P1 0.992f
C44 filter_res_magic_0.R3_R7 VOUT_OPAMP_N 0.349f
C45 Folded_Diff_Op_Amp_Layout_0.IB5 Folded_Diff_Op_Amp_Layout_0.IB2 0.00262f
C46 Folded_Diff_Op_Amp_Layout_0.VBIASN Folded_Diff_Op_Amp_Layout_0.IBIAS4 0.155f
C47 VOUT_OPAMP_P VOUT_P 0.964f
C48 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.IBIAS1 0.196f
C49 filter_res_magic_0.R3_R7 VIN_P1 0.189f
C50 Folded_Diff_Op_Amp_Layout_0.IB5 VDD 1.28f
C51 Folded_Diff_Op_Amp_Layout_0.BD VDD 8.89f
C52 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VND 6.12f
C53 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB3 1.58f
C54 Folded_Diff_Op_Amp_Layout_0.BD VOUT_N 0.102f
C55 VOUT_OPAMP_N VOUT_P 5.46f
C56 VDD VCM1 1.08f
C57 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS4 0.0575f
C58 Folded_Diff_Op_Amp_Layout_0.IBIAS1 Folded_Diff_Op_Amp_Layout_0.IBS 0.361f
C59 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.IB2 0.0224f
C60 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.IBIAS3 0.063f
C61 Folded_Diff_Op_Amp_Layout_0.VBM Folded_Diff_Op_Amp_Layout_0.VBIASN 0.174f
C62 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.IB5 0.124f
C63 Folded_Diff_Op_Amp_Layout_0.VB1 VDD 9.95f
C64 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_P 4.97f
C65 Folded_Diff_Op_Amp_Layout_0.VB1 VOUT_N 4.8e-19
C66 Folded_Diff_Op_Amp_Layout_0.VCD VCM1 1.27f
C67 filter_res_magic_0.R7_R8_R10_C VIN_N1 0.504f
C68 VOUT_OPAMP_P VCM1 0.0688f
C69 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.IB5 0.562f
C70 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VBIASN 1.23f
C71 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.IBIAS3 0.00232f
C72 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VCD 7.56f
C73 filter_res_magic_0.R3_R7 VIN_N1 0.73f
C74 Folded_Diff_Op_Amp_Layout_0.BD VOUT_OPAMP_N 4.52f
C75 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB2 8.26e-20
C76 Folded_Diff_Op_Amp_Layout_0.VB4 VDD 0.72f
C77 Folded_Diff_Op_Amp_Layout_0.VB4 VOUT_N 0.0256f
C78 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IB4 1.33f
C79 VOUT_OPAMP_N VCM1 0.343f
C80 Folded_Diff_Op_Amp_Layout_0.VB3 VCM1 0.267f
C81 filter_res_magic_0.R7_R8_R10_C filter_res_magic_0.R3_R7 1.5f
C82 Folded_Diff_Op_Amp_Layout_0.IVS VDD 17.6f
C83 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VPD 10.7f
C84 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VOUT 0.0466f
C85 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VB1 0.553f
C86 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VCD 0.697f
C87 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.IB4 0.376f
C88 Folded_Diff_Op_Amp_Layout_0.IBIAS1 Folded_Diff_Op_Amp_Layout_0.IB2 0.0416f
C89 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.VBM 0.235f
C90 Folded_Diff_Op_Amp_Layout_0.IBIAS1 VDD 4.43f
C91 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB3 0.388f
C92 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB2 1.45f
C93 filter_res_magic_0.R3_R7 VOUT_P 0.562f
C94 Folded_Diff_Op_Amp_Layout_0.OUT2 VOUT_P 4.06f
C95 Folded_Diff_Op_Amp_Layout_0.VBM Folded_Diff_Op_Amp_Layout_0.IBS 0.409f
C96 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.IB3 0.0152f
C97 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.VB2 0.0347f
C98 VIN_N1 VCM1 0.27f
C99 Folded_Diff_Op_Amp_Layout_0.VND VDD 9.42f
C100 Folded_Diff_Op_Amp_Layout_0.VND VOUT_N 0.00416f
C101 Folded_Diff_Op_Amp_Layout_0.VOUT VCM1 2.45f
C102 filter_res_magic_0.R7_R8_R10_C VCM1 0.0163f
C103 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.IBS 1.95f
C104 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.IBIAS1 0.0776f
C105 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VOUT 6.79f
C106 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.OUT1 0.874f
C107 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB2 2.07e-20
C108 filter_res_magic_0.R3_R7 VCM1 1.25f
C109 Folded_Diff_Op_Amp_Layout_0.BD VOUT_P 0.0197f
C110 Folded_Diff_Op_Amp_Layout_0.VBIASN Folded_Diff_Op_Amp_Layout_0.IB3 3.45e-20
C111 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IVS 2.78f
C112 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.VBIASN 0.317f
C113 Folded_Diff_Op_Amp_Layout_0.OUT2 VCM1 0.00142f
C114 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.IBIAS 0.0029f
C115 Folded_Diff_Op_Amp_Layout_0.IBIAS4 VDD 3.94f
C116 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB1 0.3f
C117 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.IBIAS2 0.431f
C118 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VOUT 0.0396f
C119 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VPD 0.982f
C120 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VND 2.36e-19
C121 VOUT_P VCM1 0.282f
C122 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.IB4 0.0425f
C123 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.IVS 0.0183f
C124 Folded_Diff_Op_Amp_Layout_0.VBM Folded_Diff_Op_Amp_Layout_0.IB2 0.0221f
C125 Folded_Diff_Op_Amp_Layout_0.IBS Folded_Diff_Op_Amp_Layout_0.VBIASN 1.95f
C126 Folded_Diff_Op_Amp_Layout_0.VBM VDD 1.58f
C127 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.IPD 14.3f
C128 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.OUT2 0.00296f
C129 Folded_Diff_Op_Amp_Layout_0.BD VCM1 1.38e-19
C130 Folded_Diff_Op_Amp_Layout_0.VB4 VOUT_P 0.00195f
C131 Folded_Diff_Op_Amp_Layout_0.VBM Folded_Diff_Op_Amp_Layout_0.VCD 7.59f
C132 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.IB5 0.53f
C133 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.IB2 2.01f
C134 Folded_Diff_Op_Amp_Layout_0.VB2 VDD 12.7f
C135 Folded_Diff_Op_Amp_Layout_0.VB2 VOUT_N 4.8e-19
C136 Folded_Diff_Op_Amp_Layout_0.IVS Folded_Diff_Op_Amp_Layout_0.IB4 1.15f
C137 Folded_Diff_Op_Amp_Layout_0.VB1 VCM1 1.11f
C138 filter_res_magic_0.R7_R8_R10_C m3_n10442_12259# 0.0764f
C139 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.IB5 0.719f
C140 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VCD 0.0792f
C141 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VBM 0.0534f
C142 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.OUT1 4.85f
C143 Folded_Diff_Op_Amp_Layout_0.VBIASN Folded_Diff_Op_Amp_Layout_0.IB2 0.0176f
C144 Folded_Diff_Op_Amp_Layout_0.IBS Folded_Diff_Op_Amp_Layout_0.IB3 0.00347f
C145 Folded_Diff_Op_Amp_Layout_0.IBIAS3 Folded_Diff_Op_Amp_Layout_0.IBIAS4 0.739f
C146 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.IBS 0.597f
C147 Folded_Diff_Op_Amp_Layout_0.VB4 VCM1 0.814f
C148 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.IBIAS 0.00217f
C149 Folded_Diff_Op_Amp_Layout_0.VBIASN VDD 1.45f
C150 Folded_Diff_Op_Amp_Layout_0.IPD VDD 2.94f
C151 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB1 0.193f
C152 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VPD 0.748f
C153 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VND 1.17f
C154 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB3 0.619f
C155 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_N 0.239f
C156 Folded_Diff_Op_Amp_Layout_0.VND VOUT_P 0.00173f
C157 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.VBIASN 0.391f
C158 Folded_Diff_Op_Amp_Layout_0.IBIAS1 Folded_Diff_Op_Amp_Layout_0.IB5 0.186f
C159 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.IBIAS4 0.0051f
C160 Folded_Diff_Op_Amp_Layout_0.IBIAS2 VDD 0.142p
C161 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_P 0.59f
C162 Folded_Diff_Op_Amp_Layout_0.IBIAS2 VOUT_N 14.4f
C163 Folded_Diff_Op_Amp_Layout_0.IBIAS1 VCM1 0.0208f
C164 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VBIASN 0.285f
C165 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.VBM 0.542f
C166 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.IBIAS1 0.0893f
C167 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.VB3 0.53f
C168 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_OPAMP_N 0.486f
C169 Folded_Diff_Op_Amp_Layout_0.OUT1 VDD 8.72f
C170 Folded_Diff_Op_Amp_Layout_0.OUT1 VOUT_N 5.21f
C171 Folded_Diff_Op_Amp_Layout_0.IBIAS4 Folded_Diff_Op_Amp_Layout_0.IB4 0.949f
C172 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.IB2 0.0141f
C173 Folded_Diff_Op_Amp_Layout_0.IBIAS VDD 10.1f
C174 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VOUT 0.149f
C175 Folded_Diff_Op_Amp_Layout_0.VND Folded_Diff_Op_Amp_Layout_0.VB1 0.78f
C176 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.VCD 0.515f
C177 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.IB3 5.9e-19
C178 Folded_Diff_Op_Amp_Layout_0.IBIAS VOUT_OPAMP_P 0.216f
C179 Folded_Diff_Op_Amp_Layout_0.IBS VDD 2.11f
C180 Folded_Diff_Op_Amp_Layout_0.IND VDD 7.04f
C181 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.VB2 1.03f
C182 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VB3 1.2f
C183 Folded_Diff_Op_Amp_Layout_0.IND VOUT_N 0.613f
C184 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.IB4 0.00218f
C185 Folded_Diff_Op_Amp_Layout_0.VCD Folded_Diff_Op_Amp_Layout_0.IBS 0.0309f
C186 Folded_Diff_Op_Amp_Layout_0.IBIAS VOUT_OPAMP_N 0.281f
C187 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.IB3 1.09f
C188 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.VB3 0.656f
C189 Folded_Diff_Op_Amp_Layout_0.VBM Folded_Diff_Op_Amp_Layout_0.IB5 0.101f
C190 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IBIAS3 1.68f
C191 Folded_Diff_Op_Amp_Layout_0.VPD VDD 10.7f
C192 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_P 0.571f
C193 Folded_Diff_Op_Amp_Layout_0.VPD VOUT_N 5.25e-19
C194 Folded_Diff_Op_Amp_Layout_0.VBM VCM1 6.49f
C195 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.IBIAS3 0.00364f
C196 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.VOUT 0.00234f
C197 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.IB5 0.004f
C198 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.IBS 1.14f
C199 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VBM 2.6f
C200 Folded_Diff_Op_Amp_Layout_0.IPD Folded_Diff_Op_Amp_Layout_0.OUT2 5.04f
C201 Folded_Diff_Op_Amp_Layout_0.IND Folded_Diff_Op_Amp_Layout_0.VB3 0.576f
C202 Folded_Diff_Op_Amp_Layout_0.IND VOUT_OPAMP_N 0.716f
C203 Folded_Diff_Op_Amp_Layout_0.IPD VOUT_P 0.0039f
C204 Folded_Diff_Op_Amp_Layout_0.IBIAS4 Folded_Diff_Op_Amp_Layout_0.IVS 0.393f
C205 Folded_Diff_Op_Amp_Layout_0.VBIASN Folded_Diff_Op_Amp_Layout_0.IB4 0.0856f
C206 Folded_Diff_Op_Amp_Layout_0.VB2 VCM1 5.28e-19
C207 Folded_Diff_Op_Amp_Layout_0.IB2 VDD 0.845f
C208 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VBM 0.525f
C209 Folded_Diff_Op_Amp_Layout_0.OUT2 Folded_Diff_Op_Amp_Layout_0.IBIAS2 5.16e-19
C210 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.VOUT 1.63f
C211 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.VB1 0.191f
C212 VDD VOUT_N 91.5f
C213 Folded_Diff_Op_Amp_Layout_0.IBIAS2 VOUT_P 16.4f
C214 Folded_Diff_Op_Amp_Layout_0.IB5 Folded_Diff_Op_Amp_Layout_0.VBIASN 1.08f
C215 Folded_Diff_Op_Amp_Layout_0.IBIAS Folded_Diff_Op_Amp_Layout_0.VOUT 0.352f
C216 Folded_Diff_Op_Amp_Layout_0.IBIAS2 Folded_Diff_Op_Amp_Layout_0.IB4 0.725f
C217 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.IB3 1.55e-19
C218 Folded_Diff_Op_Amp_Layout_0.VCD VDD 0.0177f
C219 Folded_Diff_Op_Amp_Layout_0.BD Folded_Diff_Op_Amp_Layout_0.IPD 9.31f
C220 VDD VOUT_OPAMP_P 9.52f
C221 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.OUT2 30.1f
C222 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VB2 0.0126f
C223 VOUT_OPAMP_P VOUT_N 4.45f
C224 Folded_Diff_Op_Amp_Layout_0.IBIAS filter_res_magic_0.R3_R7 0.287f
C225 Folded_Diff_Op_Amp_Layout_0.VBIASN VCM1 0.0164f
C226 Folded_Diff_Op_Amp_Layout_0.IPD VCM1 1.19e-19
C227 Folded_Diff_Op_Amp_Layout_0.OUT1 VOUT_P 5.73f
C228 Folded_Diff_Op_Amp_Layout_0.OUT1 Folded_Diff_Op_Amp_Layout_0.IB4 0.0172f
C229 Folded_Diff_Op_Amp_Layout_0.VBM Folded_Diff_Op_Amp_Layout_0.IBIAS1 0.243f
C230 Folded_Diff_Op_Amp_Layout_0.VOUT Folded_Diff_Op_Amp_Layout_0.IBS 0.0174f
C231 Folded_Diff_Op_Amp_Layout_0.VB1 Folded_Diff_Op_Amp_Layout_0.VBIASN 0.128f
C232 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.IVS 0.0083f
C233 Folded_Diff_Op_Amp_Layout_0.VB3 VDD 0.946f
C234 VDD VOUT_OPAMP_N 10.1f
C235 VOUT_OPAMP_N VOUT_N 2.75f
C236 VDD VIN_P1 0.654f
C237 Folded_Diff_Op_Amp_Layout_0.IBIAS VOUT_P 0.163f
C238 Folded_Diff_Op_Amp_Layout_0.VB2 Folded_Diff_Op_Amp_Layout_0.IBIAS1 0.0175f
C239 Folded_Diff_Op_Amp_Layout_0.VB3 Folded_Diff_Op_Amp_Layout_0.VCD 0.713f
C240 Folded_Diff_Op_Amp_Layout_0.VB4 Folded_Diff_Op_Amp_Layout_0.VBIASN 0.108f
.ends

