magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -1991 -3127 4457 2666
<< nwell >>
rect 152 484 2433 666
rect 2152 -484 2433 484
<< psubdiff >>
rect 664 -1057 1679 -1042
rect 664 -1103 973 -1057
rect 1489 -1103 1679 -1057
rect 664 -1121 1679 -1103
<< nsubdiff >>
rect 192 603 2406 642
rect 192 557 938 603
rect 1548 557 2406 603
rect 192 524 2406 557
<< psubdiffcont >>
rect 973 -1103 1489 -1057
<< nsubdiffcont >>
rect 938 557 1548 603
<< polysilicon >>
rect 326 398 870 442
rect 974 398 1518 442
rect 94 -15 181 -10
rect 94 -29 251 -15
rect 94 -75 118 -29
rect 164 -46 251 -29
rect 164 -75 654 -46
rect 94 -86 654 -75
rect 758 -86 870 86
rect 974 40 1086 86
rect 974 -25 1174 40
rect 974 -71 1047 -25
rect 1093 -71 1174 -25
rect 1866 18 1978 86
rect 2106 18 2190 20
rect 1866 1 2190 18
rect 1866 -45 2122 1
rect 2168 -45 2190 1
rect 1866 -61 2190 -45
rect 974 -86 1174 -71
rect 94 -92 251 -86
rect 1086 -94 1174 -86
rect 1434 -99 1762 -63
rect 1866 -86 1978 -61
rect 2106 -63 2190 -61
rect 758 -447 870 -398
rect 1434 -410 1546 -334
rect 67 -469 870 -447
rect 67 -515 89 -469
rect 135 -484 870 -469
rect 1129 -463 1241 -446
rect 135 -515 377 -484
rect 67 -532 377 -515
rect 1129 -509 1162 -463
rect 1208 -509 1241 -463
rect 1129 -532 1241 -509
rect 1345 -470 1546 -410
rect 1861 -405 2321 -375
rect 1861 -451 1880 -405
rect 1926 -431 2321 -405
rect 1926 -451 1947 -431
rect 1861 -469 1947 -451
rect 1345 -516 1377 -470
rect 1423 -486 1546 -470
rect 1423 -516 1457 -486
rect 1345 -532 1457 -516
rect 2209 -532 2321 -431
rect 67 -535 265 -532
rect 481 -981 593 -841
rect 697 -848 809 -800
rect 913 -848 1025 -800
rect 697 -870 1025 -848
rect 697 -916 725 -870
rect 771 -885 1025 -870
rect 1129 -868 1241 -841
rect 771 -916 809 -885
rect 697 -933 809 -916
rect 1129 -914 1153 -868
rect 1199 -914 1241 -868
rect 1129 -981 1241 -914
rect 481 -1019 1241 -981
rect 1345 -981 1457 -841
rect 1561 -868 1889 -841
rect 1561 -914 1584 -868
rect 1630 -877 1889 -868
rect 1630 -914 1673 -877
rect 1561 -933 1673 -914
rect 1993 -981 2105 -841
rect 1345 -1019 2105 -981
<< polycontact >>
rect 118 -75 164 -29
rect 1047 -71 1093 -25
rect 2122 -45 2168 1
rect 89 -515 135 -469
rect 1162 -509 1208 -463
rect 1880 -451 1926 -405
rect 1377 -516 1423 -470
rect 725 -916 771 -870
rect 1153 -914 1199 -868
rect 1584 -914 1630 -868
<< metal1 >>
rect 192 603 2406 642
rect 192 557 938 603
rect 1548 557 2406 603
rect 192 524 2406 557
rect 251 444 297 524
rect 251 398 729 444
rect 251 341 297 398
rect 683 341 729 398
rect 1115 398 1593 444
rect 1115 341 1161 398
rect 1547 341 1593 398
rect 1791 341 1837 524
rect 94 -25 175 -10
rect 22 -26 175 -25
rect 22 -78 115 -26
rect 167 -78 175 -26
rect 94 -90 175 -78
rect 251 -40 297 143
rect 467 86 513 143
rect 899 86 945 143
rect 1331 86 1377 143
rect 467 40 1377 86
rect 251 -86 729 -40
rect 251 -143 297 -86
rect 683 -143 729 -86
rect 899 -143 945 40
rect 1023 -20 1123 -7
rect 1547 -19 1593 143
rect 1023 -72 1043 -20
rect 1095 -72 1123 -20
rect 1023 -83 1123 -72
rect 1230 -73 1593 -19
rect 1023 -94 1077 -83
rect 1230 -238 1284 -73
rect 1791 -143 1837 143
rect 2007 -143 2053 143
rect 2106 1 2285 18
rect 2106 -45 2122 1
rect 2168 -45 2285 1
rect 2106 -61 2285 -45
rect 442 -268 538 -264
rect 442 -320 464 -268
rect 516 -320 538 -268
rect 442 -332 538 -320
rect 1014 -322 1144 -276
rect 1161 -292 1284 -238
rect 1356 -286 1427 -271
rect 1014 -398 1060 -322
rect 1356 -338 1361 -286
rect 1413 -338 1427 -286
rect 1356 -354 1427 -338
rect 1767 -286 1837 -271
rect 1767 -338 1781 -286
rect 1833 -338 1837 -286
rect 190 -444 1060 -398
rect 1575 -401 1621 -341
rect 1767 -354 1837 -338
rect 2007 -353 2396 -307
rect 1866 -401 1943 -398
rect 1575 -405 1943 -401
rect 67 -463 142 -447
rect 9 -469 142 -463
rect 9 -515 89 -469
rect 135 -515 142 -469
rect 9 -521 142 -515
rect 67 -535 142 -521
rect 190 -586 236 -444
rect 1142 -460 1229 -447
rect 1575 -448 1880 -405
rect 1142 -512 1159 -460
rect 1211 -512 1229 -460
rect 1142 -525 1229 -512
rect 1361 -467 1440 -453
rect 1361 -519 1374 -467
rect 1426 -519 1440 -467
rect 1361 -533 1440 -519
rect 813 -576 910 -563
rect 813 -628 835 -576
rect 887 -628 910 -576
rect 1702 -586 1748 -448
rect 1861 -451 1880 -448
rect 1926 -451 1943 -405
rect 1861 -457 1943 -451
rect 2350 -442 2396 -353
rect 2350 -488 2457 -442
rect 2350 -586 2396 -488
rect 813 -641 910 -628
rect 622 -732 689 -716
rect 622 -784 623 -732
rect 675 -784 689 -732
rect 190 -869 236 -787
rect 180 -881 260 -869
rect 180 -933 194 -881
rect 246 -933 260 -881
rect 180 -948 260 -933
rect 406 -1037 452 -784
rect 622 -799 689 -784
rect 1031 -731 1107 -718
rect 1031 -783 1043 -731
rect 1095 -783 1107 -731
rect 1031 -796 1107 -783
rect 1476 -732 1555 -711
rect 1476 -784 1487 -732
rect 1539 -784 1555 -732
rect 703 -865 791 -851
rect 703 -917 721 -865
rect 773 -917 791 -865
rect 703 -932 791 -917
rect 1132 -865 1220 -851
rect 1132 -917 1150 -865
rect 1202 -917 1220 -865
rect 1132 -931 1220 -917
rect 1270 -1037 1316 -784
rect 1476 -799 1555 -784
rect 1889 -731 1987 -711
rect 1889 -783 1913 -731
rect 1965 -783 1987 -731
rect 1889 -797 1987 -783
rect 1563 -865 1651 -850
rect 1563 -917 1581 -865
rect 1633 -917 1651 -865
rect 1563 -930 1651 -917
rect 2134 -1037 2180 -784
rect 178 -1057 2456 -1037
rect 178 -1103 973 -1057
rect 1489 -1103 2456 -1057
rect 178 -1127 2456 -1103
<< via1 >>
rect 115 -29 167 -26
rect 115 -75 118 -29
rect 118 -75 164 -29
rect 164 -75 167 -29
rect 115 -78 167 -75
rect 1043 -25 1095 -20
rect 1043 -71 1047 -25
rect 1047 -71 1093 -25
rect 1093 -71 1095 -25
rect 1043 -72 1095 -71
rect 464 -320 516 -268
rect 1361 -338 1413 -286
rect 1781 -338 1833 -286
rect 1159 -463 1211 -460
rect 1159 -509 1162 -463
rect 1162 -509 1208 -463
rect 1208 -509 1211 -463
rect 1159 -512 1211 -509
rect 1374 -470 1426 -467
rect 1374 -516 1377 -470
rect 1377 -516 1423 -470
rect 1423 -516 1426 -470
rect 1374 -519 1426 -516
rect 835 -628 887 -576
rect 623 -784 675 -732
rect 194 -933 246 -881
rect 1043 -783 1095 -731
rect 1487 -784 1539 -732
rect 721 -870 773 -865
rect 721 -916 725 -870
rect 725 -916 771 -870
rect 771 -916 773 -870
rect 721 -917 773 -916
rect 1150 -868 1202 -865
rect 1150 -914 1153 -868
rect 1153 -914 1199 -868
rect 1199 -914 1202 -868
rect 1150 -917 1202 -914
rect 1913 -783 1965 -731
rect 1581 -868 1633 -865
rect 1581 -914 1584 -868
rect 1584 -914 1630 -868
rect 1630 -914 1633 -868
rect 1581 -917 1633 -914
<< metal2 >>
rect 175 -15 251 -10
rect 1023 -15 1123 3
rect 100 -20 1123 -15
rect 100 -26 1043 -20
rect 100 -78 115 -26
rect 167 -72 1043 -26
rect 1095 -72 1123 -20
rect 167 -78 1123 -72
rect 100 -86 251 -78
rect 175 -90 251 -86
rect 1023 -94 1123 -78
rect 442 -268 538 -264
rect 442 -320 464 -268
rect 516 -320 538 -268
rect 442 -332 538 -320
rect 454 -450 526 -332
rect 1037 -446 1095 -94
rect 1356 -286 1837 -271
rect 1356 -338 1361 -286
rect 1413 -338 1781 -286
rect 1833 -338 1837 -286
rect 1356 -354 1837 -338
rect 454 -506 898 -450
rect 825 -563 898 -506
rect 1037 -460 1241 -446
rect 1037 -512 1159 -460
rect 1211 -512 1241 -460
rect 1037 -528 1241 -512
rect 1361 -465 1440 -453
rect 1361 -521 1372 -465
rect 1428 -521 1440 -465
rect 1361 -533 1440 -521
rect 813 -576 910 -563
rect 813 -632 834 -576
rect 890 -632 910 -576
rect 813 -641 910 -632
rect 609 -728 689 -716
rect 1031 -728 1115 -718
rect 609 -731 1115 -728
rect 609 -732 1043 -731
rect 609 -784 623 -732
rect 675 -783 1043 -732
rect 1095 -783 1115 -731
rect 675 -784 1115 -783
rect 609 -786 1115 -784
rect 609 -799 689 -786
rect 1031 -796 1115 -786
rect 1473 -731 1987 -711
rect 1473 -732 1913 -731
rect 1473 -784 1487 -732
rect 1539 -783 1913 -732
rect 1965 -783 1987 -731
rect 1539 -784 1987 -783
rect 1473 -797 1987 -784
rect 1473 -799 1972 -797
rect 730 -859 791 -851
rect 712 -863 791 -859
rect 248 -865 791 -863
rect 248 -869 721 -865
rect 180 -881 721 -869
rect 180 -933 194 -881
rect 246 -917 721 -881
rect 773 -917 791 -865
rect 246 -932 791 -917
rect 1132 -863 1220 -851
rect 1563 -863 1651 -856
rect 1132 -865 1651 -863
rect 1132 -917 1150 -865
rect 1202 -917 1581 -865
rect 1633 -917 1651 -865
rect 1132 -919 1651 -917
rect 1132 -931 1220 -919
rect 1563 -930 1651 -919
rect 246 -933 779 -932
rect 180 -948 260 -933
<< via2 >>
rect 1372 -467 1428 -465
rect 1372 -519 1374 -467
rect 1374 -519 1426 -467
rect 1426 -519 1428 -467
rect 1372 -521 1428 -519
rect 834 -628 835 -576
rect 835 -628 887 -576
rect 887 -628 890 -576
rect 834 -632 890 -628
<< metal3 >>
rect 813 -465 1457 -453
rect 813 -521 1372 -465
rect 1428 -521 1457 -465
rect 813 -535 1457 -521
rect 813 -576 910 -535
rect 813 -632 834 -576
rect 890 -632 910 -576
rect 813 -641 910 -632
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_0
timestamp 1713185578
transform 1 0 321 0 1 -688
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_1
timestamp 1713185578
transform 1 0 537 0 1 -688
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_2
timestamp 1713185578
transform 1 0 1185 0 1 -688
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_3
timestamp 1713185578
transform 1 0 1401 0 1 -688
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_4
timestamp 1713185578
transform 1 0 2049 0 1 -688
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_5
timestamp 1713185578
transform 1 0 2265 0 1 -688
box -168 -180 168 180
use nmos_3p3_F2UGVV  nmos_3p3_F2UGVV_0
timestamp 1713185578
transform 1 0 861 0 1 -688
box -276 -180 276 180
use nmos_3p3_F2UGVV  nmos_3p3_F2UGVV_1
timestamp 1713185578
transform 1 0 1725 0 1 -688
box -276 -180 276 180
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_0
timestamp 1713185578
transform 1 0 814 0 1 242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_1
timestamp 1713185578
transform 1 0 382 0 1 242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_2
timestamp 1713185578
transform 1 0 382 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_3
timestamp 1713185578
transform 1 0 1030 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_4
timestamp 1713185578
transform 1 0 814 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_5
timestamp 1713185578
transform 1 0 598 0 1 242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_6
timestamp 1713185578
transform 1 0 1922 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_7
timestamp 1713185578
transform 1 0 1706 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_8
timestamp 1713185578
transform 1 0 598 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_9
timestamp 1713185578
transform 1 0 1490 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_10
timestamp 1713185578
transform 1 0 1030 0 1 242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_11
timestamp 1713185578
transform 1 0 1246 0 1 242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_12
timestamp 1713185578
transform 1 0 1462 0 1 242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_13
timestamp 1713185578
transform 1 0 1922 0 1 242
box -230 -242 230 242
<< labels >>
flabel nsubdiffcont 1245 581 1245 581 0 FreeSans 750 0 0 0 VDD
flabel psubdiffcont 1229 -1083 1229 -1083 0 FreeSans 750 0 0 0 VSS
flabel metal1 s 40 -49 40 -49 0 FreeSans 250 0 0 0 CLK
port 1 nsew
flabel metal1 s 22 -498 22 -498 0 FreeSans 250 0 0 0 D
port 2 nsew
flabel metal1 s 2428 -466 2428 -466 0 FreeSans 750 0 0 0 Q
port 3 nsew
flabel metal1 s 2250 -25 2250 -25 0 FreeSans 750 0 0 0 QB
port 4 nsew
<< end >>
