** sch_path: /home/shahid/GF180Projects/Top_test/top/xschem/VCO_TB.sch
**.subckt VCO_TB OUT OUTB
*.opin OUT
*.opin OUTB
VCNTL VCONT GND 1.075
.save i(vcntl)
V2 VDD GND PWL( 0 0 100n 0 100.001n 3.3)
.save i(v2)
VCNTL1 VSS GND 0
.save i(vcntl1)
V1 EN GND 3.3
.save i(v1)
x1 VDD EN OUT OUTB VCONT VSS VCO_PEX
**** begin user architecture code


.include VCO_PEX.spice
.control
set color0=white
set color1=black

save all
tran 10p 200n
plot v(OUT) v(OUTB)+4
write VCO_TB.raw
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
