magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1682 -1022 1022 1022
<< metal4 >>
rect -679 14 19 19
rect -679 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 19 14
rect -679 -19 19 -14
<< via4 >>
rect -674 -14 -646 14
rect -608 -14 -580 14
rect -542 -14 -514 14
rect -476 -14 -448 14
rect -410 -14 -382 14
rect -344 -14 -316 14
rect -278 -14 -250 14
rect -212 -14 -184 14
rect -146 -14 -118 14
rect -80 -14 -52 14
rect -14 -14 14 14
<< metal5 >>
rect -682 14 22 22
rect -682 -14 -674 14
rect -646 -14 -608 14
rect -580 -14 -542 14
rect -514 -14 -476 14
rect -448 -14 -410 14
rect -382 -14 -344 14
rect -316 -14 -278 14
rect -250 -14 -212 14
rect -184 -14 -146 14
rect -118 -14 -80 14
rect -52 -14 -14 14
rect 14 -14 22 14
rect -682 -22 22 -14
<< end >>
