magic
tech gf180mcuC
magscale 1 10
timestamp 1693223404
<< nwell >>
rect 11880 4374 11981 4464
rect 9432 3387 12398 3389
rect 3198 3117 6016 3315
rect 9432 3135 12407 3387
rect 5394 3028 6015 3117
rect 11641 3036 12407 3135
rect 5395 3026 5797 3028
rect 11643 3023 12407 3036
rect 217 2206 622 2377
rect 217 2090 2160 2206
rect 403 1995 2160 2090
rect 6247 2158 9356 2261
rect 6247 2097 9667 2158
rect 6247 1996 9356 2097
rect 9064 1995 9356 1996
rect 9064 1986 9288 1995
<< nsubdiff >>
rect 4380 3135 5428 3250
rect 655 2095 922 2177
rect 1225 2110 1561 2168
rect 6733 2068 9206 2213
rect 7749 2012 7832 2068
rect 8313 2037 8396 2068
<< metal1 >>
rect -258 5173 6745 5409
rect 8567 5253 12153 5432
rect -258 3104 -41 5173
rect 5822 4702 5917 4721
rect 5822 4612 5835 4702
rect 5901 4612 5917 4702
rect 5822 4590 5917 4612
rect 6472 4588 6745 5173
rect 8569 4588 8848 5253
rect 11869 4935 11969 4947
rect 11869 4880 11902 4935
rect 11958 4880 11969 4935
rect 11869 4868 11969 4880
rect 6098 4514 6231 4521
rect 6098 4421 6114 4514
rect 6212 4421 6231 4514
rect 6098 4410 6231 4421
rect 6472 4345 8848 4588
rect 9045 4532 9233 4588
rect 9045 4402 9084 4532
rect 9210 4402 9233 4532
rect 9045 4361 9233 4402
rect 9421 4455 11997 4493
rect 9421 4386 11890 4455
rect 11966 4386 11997 4455
rect 6375 4166 8978 4345
rect 9421 4338 11997 4386
rect 8739 4163 8848 4166
rect 11860 3845 11934 3853
rect 8682 3824 8759 3836
rect 8682 3762 8696 3824
rect 8748 3762 8759 3824
rect 11860 3793 11869 3845
rect 11926 3793 11934 3845
rect 12464 3803 12584 3804
rect 11860 3779 11934 3793
rect 8682 3750 8759 3762
rect 12288 3731 12584 3803
rect 9432 3387 12398 3389
rect 6246 3331 8822 3376
rect 6004 3323 8822 3331
rect 6004 3315 8681 3323
rect 3198 3254 8681 3315
rect 8757 3254 8822 3323
rect 3198 3221 8822 3254
rect 3198 3117 6277 3221
rect 9432 3135 12407 3387
rect -258 3085 2167 3104
rect -258 2975 -131 3085
rect -24 2975 2167 3085
rect 5394 3033 6277 3117
rect 11641 3036 12407 3135
rect 5394 3028 6015 3033
rect 5395 3026 5797 3028
rect 11643 3023 12407 3036
rect -258 2964 2167 2975
rect -171 2952 9 2964
rect -283 2658 302 2772
rect 8676 2739 8753 2748
rect 8676 2674 8688 2739
rect 8742 2674 8753 2739
rect 9523 2698 9635 2709
rect 9523 2689 9541 2698
rect 8676 2662 8753 2674
rect -283 1693 -177 2658
rect 9095 2621 9541 2689
rect 9617 2621 9635 2698
rect 12464 2634 12584 3731
rect 6031 2602 6138 2611
rect 6031 2586 6040 2602
rect 5740 2528 6040 2586
rect 6031 2521 6040 2528
rect 6130 2521 6138 2602
rect 9095 2604 9635 2621
rect 9095 2595 9634 2604
rect 11955 2576 12584 2634
rect 11987 2536 12584 2576
rect 6031 2504 6138 2521
rect 217 2206 622 2377
rect 217 2090 2160 2206
rect 403 1995 2160 2090
rect 6247 2158 9356 2261
rect 6247 2097 9667 2158
rect 6247 1996 9356 2097
rect 9140 1995 9356 1996
rect -283 1661 204 1693
rect -283 1587 206 1661
rect -155 1383 25 1408
rect -155 1273 -131 1383
rect -24 1382 25 1383
rect -24 1336 51 1382
rect -24 1285 56 1336
rect -24 1273 25 1285
rect -155 1256 25 1273
rect 12306 127 12448 2315
rect 6024 113 12448 127
rect 237 -108 12448 113
rect 237 -109 12407 -108
rect 237 -117 6680 -109
rect 237 -123 6130 -117
<< via1 >>
rect 5835 4612 5901 4702
rect 11902 4880 11958 4935
rect 10849 4785 10908 4837
rect 6114 4421 6212 4514
rect 9084 4402 9210 4532
rect 11890 4386 11966 4455
rect 8696 3762 8748 3824
rect 11869 3793 11926 3845
rect 7677 3668 7730 3720
rect 8681 3254 8757 3323
rect -131 2975 -24 3085
rect 8688 2674 8742 2739
rect 9541 2621 9617 2698
rect 6040 2521 6130 2602
rect -131 1273 -24 1383
<< metal2 >>
rect 11869 4935 11969 4947
rect 11869 4880 11902 4935
rect 11958 4880 11969 4935
rect 11869 4868 11969 4880
rect 10833 4846 10936 4851
rect 10833 4776 10844 4846
rect 10926 4776 10936 4846
rect 10833 4766 10936 4776
rect 5822 4702 5917 4721
rect 5822 4693 5835 4702
rect 5204 4637 5835 4693
rect 5204 4584 5260 4637
rect 5822 4612 5835 4637
rect 5901 4612 5917 4702
rect 5822 4590 5917 4612
rect 9045 4532 9233 4588
rect 6098 4514 6231 4521
rect 6098 4421 6114 4514
rect 6212 4421 6231 4514
rect 6098 4410 6231 4421
rect -171 3085 9 3104
rect -171 2975 -131 3085
rect -24 2975 9 3085
rect -171 2952 9 2975
rect 6108 2955 6208 4410
rect 9045 4402 9084 4532
rect 9210 4402 9233 4532
rect 11898 4464 11954 4868
rect 9045 4361 9233 4402
rect 11880 4455 11981 4464
rect 11880 4386 11890 4455
rect 11966 4386 11981 4455
rect 11880 4374 11981 4386
rect 9512 3896 9649 3952
rect 8682 3824 8759 3836
rect 8682 3762 8696 3824
rect 8748 3762 8759 3824
rect 8682 3750 8759 3762
rect 7660 3721 7762 3725
rect 7660 3645 7671 3721
rect 7740 3645 7762 3721
rect 7660 3639 7762 3645
rect 8689 3332 8752 3750
rect 8668 3323 8771 3332
rect 8668 3254 8681 3323
rect 8757 3254 8771 3323
rect 8668 3239 8771 3254
rect -121 1408 -35 2952
rect 6108 2871 6474 2955
rect 8689 2750 8752 3239
rect 8676 2739 8753 2750
rect 8676 2674 8688 2739
rect 8742 2674 8753 2739
rect 8676 2664 8753 2674
rect 9512 2709 9619 3896
rect 11898 3853 11954 4374
rect 11860 3845 11954 3853
rect 11860 3793 11869 3845
rect 11926 3793 11954 3845
rect 11860 3785 11954 3793
rect 11860 3782 11934 3785
rect 9512 2698 9635 2709
rect 9512 2621 9541 2698
rect 9617 2621 9635 2698
rect 6031 2602 6138 2611
rect 9512 2604 9635 2621
rect 9512 2603 9619 2604
rect 9535 2602 9617 2603
rect 6031 2586 6040 2602
rect 6015 2521 6040 2586
rect 6130 2521 6138 2602
rect 6015 2504 6138 2521
rect -155 1383 25 1408
rect -155 1273 -131 1383
rect -24 1273 25 1383
rect -155 1256 25 1273
rect 6015 1257 6120 2504
rect 6015 1142 7059 1257
rect 1475 632 1561 639
rect 1475 562 1481 632
rect 1550 562 1561 632
rect 1475 556 1561 562
rect 7705 633 7799 639
rect 7705 560 7716 633
rect 7792 585 7799 633
rect 7792 560 7803 585
rect 7705 556 7803 560
rect 7709 502 7803 556
<< via2 >>
rect 10844 4837 10926 4846
rect 10844 4785 10849 4837
rect 10849 4785 10908 4837
rect 10908 4785 10926 4837
rect 10844 4776 10926 4785
rect 9088 4410 9204 4515
rect 7671 3720 7740 3721
rect 7671 3668 7677 3720
rect 7677 3668 7730 3720
rect 7730 3668 7740 3720
rect 7671 3645 7740 3668
rect 1481 562 1550 632
rect 7716 560 7792 633
<< metal3 >>
rect 2805 672 2908 4862
rect 10833 4846 11004 4851
rect 10833 4776 10844 4846
rect 10926 4776 11004 4846
rect 10833 4766 11004 4776
rect 9045 4515 9233 4588
rect 9045 4410 9088 4515
rect 9204 4410 9233 4515
rect 9045 4361 9233 4410
rect 9089 3725 9191 4361
rect 10892 3725 11004 4766
rect 7660 3721 11004 3725
rect 7660 3645 7671 3721
rect 7740 3645 11004 3721
rect 7660 3639 11004 3645
rect 7684 3590 11004 3639
rect 7686 3535 11004 3590
rect 7686 672 7813 3535
rect 1475 633 7824 672
rect 1475 632 7716 633
rect 1475 562 1481 632
rect 1550 562 7716 632
rect 1475 560 7716 562
rect 7792 560 7824 633
rect 1475 556 7824 560
rect 7686 555 7770 556
use CLK_div_3_mag  CLK_div_3_mag_0
timestamp 1693072129
transform 1 0 0 0 1 1
box -34 -1 6461 3249
use CLK_div_3_mag  CLK_div_3_mag_1
timestamp 1693072129
transform -1 0 6016 0 -1 5299
box -34 -1 6461 3249
use CLK_div_3_mag  CLK_div_3_mag_2
timestamp 1693072129
transform 1 0 6247 0 1 9
box -34 -1 6461 3249
use JK_FF_mag  JK_FF_mag_0
timestamp 1692973937
transform -1 0 12003 0 -1 5389
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_1
timestamp 1692973937
transform -1 0 8828 0 -1 4272
box -390 0 2603 2148
<< labels >>
flabel via1 5850 4671 5850 4671 0 FreeSans 640 0 0 0 CLK
port 1 nsew
flabel via2 9139 4463 9139 4463 0 FreeSans 640 0 0 0 RST
port 2 nsew
flabel metal1 6093 5289 6093 5289 0 FreeSans 640 0 0 0 VSS
port 3 nsew
flabel metal1 9287 2137 9287 2137 0 FreeSans 640 0 0 0 VDD
port 4 nsew
flabel via1 6151 4466 6151 4466 0 FreeSans 640 0 0 0 Vdiv108
port 0 nsew
<< end >>
