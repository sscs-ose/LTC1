magic
tech gf180mcuC
magscale 1 10
timestamp 1694693600
<< nwell >>
rect -122 538 286 631
rect -118 526 286 538
rect -36 525 130 526
rect -32 292 31 525
<< psubdiff >>
rect -80 -95 236 -82
rect -80 -141 -67 -95
rect 223 -141 236 -95
rect -80 -154 236 -141
<< nsubdiff >>
rect -80 594 243 607
rect -80 538 -65 594
rect 229 538 243 594
rect -80 525 243 538
<< psubdiffcont >>
rect -67 -141 223 -95
<< nsubdiffcont >>
rect -65 538 229 594
<< polysilicon >>
rect -44 187 156 250
rect -44 141 31 187
rect 87 141 156 187
rect -44 103 156 141
<< polycontact >>
rect 31 141 87 187
<< metal1 >>
rect -122 594 286 631
rect -122 538 -65 594
rect 229 538 286 594
rect -122 525 286 538
rect -122 292 -59 525
rect -118 187 93 200
rect -118 141 31 187
rect 87 141 93 187
rect -118 128 93 141
rect 179 189 242 450
rect 179 131 286 189
rect -134 -69 -67 60
rect 179 14 242 131
rect -134 -95 286 -69
rect -134 -141 -67 -95
rect 223 -141 286 -95
rect -134 -175 286 -141
use nmos_3p3_MGBSF7  nmos_3p3_MGBSF7_0
timestamp 1694669839
transform 1 0 56 0 1 37
box -216 -97 216 97
use pmos_3p3_MW53B7  pmos_3p3_MW53B7_0
timestamp 1694669839
transform 1 0 56 0 1 369
box -274 -210 274 210
<< labels >>
flabel nsubdiffcont 82 566 82 566 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel psubdiffcont 80 -120 80 -120 0 FreeSans 640 0 0 0 VSS
port 1 nsew
flabel metal1 -106 158 -106 158 0 FreeSans 640 0 0 0 IN
port 2 nsew
flabel metal1 276 159 276 159 0 FreeSans 640 0 0 0 OUT
port 3 nsew
<< end >>
