magic
tech gf180mcuC
magscale 1 10
timestamp 1694669839
<< nwell >>
rect -64 708 500 863
rect -64 682 32 708
rect 33 682 500 708
rect 191 384 243 624
<< psubdiff >>
rect 13 -105 402 -91
rect 13 -151 75 -105
rect 333 -151 402 -105
rect 13 -167 402 -151
<< nsubdiff >>
rect 41 774 395 826
rect 41 728 85 774
rect 312 728 395 774
rect 41 710 395 728
<< psubdiffcont >>
rect 75 -151 333 -105
<< nsubdiffcont >>
rect 85 728 312 774
<< polysilicon >>
rect 311 421 391 427
rect 112 334 166 421
rect 63 318 166 334
rect 63 268 81 318
rect 130 268 166 318
rect 63 254 166 268
rect 112 200 166 254
rect 272 414 391 421
rect 272 366 326 414
rect 374 366 391 414
rect 272 360 391 366
rect 272 350 390 360
rect 272 200 327 350
<< polycontact >>
rect 81 268 130 318
rect 326 366 374 414
<< metal1 >>
rect -64 817 500 863
rect -64 774 499 817
rect -64 728 85 774
rect 312 728 499 774
rect -64 708 499 728
rect 33 471 89 708
rect 191 545 243 624
rect 186 470 253 545
rect 354 473 411 708
rect 63 325 144 334
rect 53 318 144 325
rect 53 278 81 318
rect 63 268 81 278
rect 130 268 144 318
rect 63 254 144 268
rect 191 314 243 470
rect 311 414 465 418
rect 311 366 326 414
rect 374 366 465 414
rect 311 361 465 366
rect 311 360 391 361
rect 191 265 406 314
rect 34 -79 88 149
rect 186 70 255 156
rect 351 80 406 265
rect -70 -105 493 -79
rect -70 -151 75 -105
rect 333 -151 493 -105
rect -70 -188 493 -151
use nmos_3p3_5QNVWA  nmos_3p3_5QNVWA_0
timestamp 1694669839
transform 1 0 140 0 1 112
box -140 -112 140 112
use nmos_3p3_5QNVWA  nmos_3p3_5QNVWA_1
timestamp 1694669839
transform 1 0 300 0 1 112
box -140 -112 140 112
use pmos_3p3_M8SWPS  pmos_3p3_M8SWPS_0
timestamp 1694669839
transform 1 0 300 0 1 545
box -202 -210 202 210
use pmos_3p3_M8SWPS  pmos_3p3_M8SWPS_1
timestamp 1694669839
transform 1 0 140 0 1 545
box -202 -210 202 210
<< labels >>
flabel nsubdiffcont 200 749 200 749 0 FreeSans 480 0 0 0 VDD
port 0 nsew
flabel polycontact 101 293 101 293 0 FreeSans 480 0 0 0 IN2
port 1 nsew
flabel metal1 425 394 425 394 0 FreeSans 480 0 0 0 IN1
port 2 nsew
flabel metal1 374 282 374 282 0 FreeSans 480 0 0 0 OUT
port 3 nsew
flabel psubdiffcont 204 -128 204 -128 0 FreeSans 480 0 0 0 VSS
port 4 nsew
<< end >>
