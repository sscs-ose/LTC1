* NGSPICE file created from mux_8x1_flat.ext - technology: gf180mcuC

.subckt mux_8x1_flat I1 I2 I3 I4 I5 I6 I7 VSS VDD OUT S0 S1 S2 I0
X0 mux_4x1_0.mux_2x1_1.I1 mux_4x1_0.mux_2x1_0.nand2_1.IN2 VDD.t42 VDD.t41 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 mux_2x1_0.nand2_1.IN2 S2.t0 a_3615_1307# VSS.t32 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X2 VDD mux_4x1_0.mux_2x1_0.nand2_2.OUT mux_4x1_0.mux_2x1_1.I1 VDD.t50 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 mux_4x1_1.mux_2x1_1.nand2_1.IN2 S1.t0 a_2490_n1395# VSS.t42 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X4 mux_4x1_1.mux_2x1_1.nand2_2.IN2 S1.t1 VDD.t79 VDD.t78 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X5 VDD mux_2x1_0.I0 mux_2x1_0.nand2_2.OUT VDD.t92 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X6 mux_2x1_0.nand2_1.IN2 mux_2x1_0.I1 VDD.t4 VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 mux_4x1_0.mux_2x1_0.nand2_2.OUT mux_4x1_0.mux_2x1_0.nand2_2.IN2 VDD.t35 VDD.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 mux_2x1_0.nand2_2.OUT mux_2x1_0.I0 a_4178_707# VSS.t4 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X9 a_1927_707# mux_4x1_0.mux_2x1_0.nand2_2.IN2 VSS.t22 VSS.t21 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X10 mux_4x1_1.mux_2x1_2.nand2_2.IN2 S0.t0 VDD.t96 VDD.t95 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X11 mux_4x1_0.mux_2x1_1.nand2_2.OUT mux_4x1_0.mux_2x1_1.nand2_2.IN2 VDD.t32 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X12 VDD S1.t2 mux_4x1_1.mux_2x1_1.nand2_1.IN2 VDD.t80 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X13 a_3053_707# mux_4x1_0.mux_2x1_1.nand2_2.IN2 VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X14 mux_4x1_1.mux_2x1_1.nand2_2.OUT mux_4x1_1.mux_2x1_1.nand2_2.IN2 VDD.t33 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 mux_4x1_1.mux_2x1_2.nand2_1.IN2 S0.t1 a_238_n1395# VSS.t57 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 a_1927_n1395# mux_4x1_1.mux_2x1_0.nand2_1.IN2 VSS.t55 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X17 mux_4x1_1.mux_2x1_2.nand2_2.OUT mux_4x1_1.mux_2x1_2.nand2_2.IN2 VDD.t40 VDD.t36 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 mux_4x1_0.mux_2x1_2.nand2_2.IN2 S0.t2 VDD.t44 VDD.t43 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 VDD mux_4x1_1.mux_2x1_1.I0 mux_4x1_1.mux_2x1_1.nand2_2.OUT VDD.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X20 VDD I4.t0 mux_4x1_0.mux_2x1_2.nand2_2.OUT VDD.t69 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X21 a_1927_1307# mux_4x1_0.mux_2x1_0.nand2_1.IN2 VSS.t28 VSS.t21 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X22 mux_4x1_0.mux_2x1_2.nand2_2.OUT I4.t1 a_801_707# VSS.t29 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X23 VDD S0.t3 mux_4x1_1.mux_2x1_2.nand2_1.IN2 VDD.t45 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X24 a_1364_n1395# I3.t0 VSS.t52 VSS.t51 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X25 mux_4x1_1.mux_2x1_1.I1 mux_4x1_1.mux_2x1_0.nand2_1.IN2 VDD.t84 VDD.t83 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X26 mux_4x1_0.mux_2x1_1.I1 mux_4x1_0.mux_2x1_0.nand2_2.OUT a_1927_1307# VSS.t14 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X27 VDD S1.t3 mux_4x1_0.mux_2x1_1.nand2_1.IN2 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X28 VDD I6.t0 mux_4x1_0.mux_2x1_0.nand2_2.OUT VDD.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X29 VDD mux_4x1_0.mux_2x1_2.nand2_2.OUT mux_4x1_0.mux_2x1_1.I0 VDD.t53 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X30 mux_4x1_1.mux_2x1_0.nand2_2.IN2 S0.t4 VDD.t65 VDD.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X31 mux_4x1_0.mux_2x1_0.nand2_2.OUT I6.t1 a_1927_707# VSS.t14 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X32 VDD mux_4x1_0.mux_2x1_1.I0 mux_4x1_0.mux_2x1_1.nand2_2.OUT VDD.t105 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 VDD S0.t5 mux_4x1_0.mux_2x1_2.nand2_1.IN2 VDD.t66 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X34 mux_4x1_0.mux_2x1_1.nand2_2.OUT mux_4x1_0.mux_2x1_1.I0 a_3053_707# VSS.t13 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X35 mux_4x1_0.mux_2x1_1.nand2_1.IN2 mux_4x1_0.mux_2x1_1.I1 VDD.t104 VDD.t103 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X36 mux_4x1_1.mux_2x1_0.nand2_1.IN2 I3.t1 VDD.t23 VDD.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 a_3615_1307# mux_2x1_0.I1 VSS.t3 VSS.t2 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X38 a_1927_n795# mux_4x1_1.mux_2x1_0.nand2_2.IN2 VSS.t46 VSS.t45 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X39 a_238_n1395# I1.t0 VSS.t49 VSS.t48 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X40 mux_4x1_1.mux_2x1_0.nand2_2.OUT I2.t0 a_1927_n795# VSS.t10 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X41 mux_4x1_1.mux_2x1_1.nand2_2.IN2 S1.t4 VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X42 mux_4x1_1.mux_2x1_2.nand2_1.IN2 I1.t1 VDD.t28 VDD.t27 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X43 mux_4x1_1.mux_2x1_2.nand2_2.IN2 S0.t6 VSS.t12 VSS.t11 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X44 mux_2x1_0.I0 mux_4x1_1.mux_2x1_1.nand2_2.OUT a_3053_n1395# VSS.t56 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X45 VDD S0.t7 mux_4x1_0.mux_2x1_0.nand2_1.IN2 VDD.t16 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X46 mux_4x1_0.mux_2x1_2.nand2_2.IN2 S0.t8 VSS.t40 VSS.t39 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X47 mux_4x1_0.mux_2x1_1.nand2_1.IN2 S1.t5 a_2490_1307# VSS.t58 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X48 mux_4x1_0.mux_2x1_1.I0 mux_4x1_0.mux_2x1_2.nand2_2.OUT a_801_1307# VSS.t29 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X49 mux_4x1_0.mux_2x1_0.nand2_1.IN2 I7.t0 VDD.t49 VDD.t48 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X50 mux_2x1_0.I1 mux_4x1_0.mux_2x1_1.nand2_1.IN2 VDD.t75 VDD.t74 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X51 mux_4x1_0.mux_2x1_1.nand2_2.IN2 S1.t6 VDD.t98 VDD.t97 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X52 a_2490_1307# mux_4x1_0.mux_2x1_1.I1 VSS.t62 VSS.t61 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X53 mux_4x1_0.mux_2x1_2.nand2_1.IN2 S0.t9 a_238_1307# VSS.t41 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X54 VDD mux_4x1_1.mux_2x1_1.nand2_2.OUT mux_2x1_0.I0 VDD.t87 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X55 mux_4x1_0.mux_2x1_0.nand2_2.IN2 S0.t10 VDD.t57 VDD.t56 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X56 mux_4x1_0.mux_2x1_1.I0 mux_4x1_0.mux_2x1_2.nand2_1.IN2 VDD.t73 VDD.t72 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X57 VDD mux_4x1_0.mux_2x1_1.nand2_2.OUT mux_2x1_0.I1 VDD.t19 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X58 mux_4x1_0.mux_2x1_2.nand2_1.IN2 I5.t0 VDD.t91 VDD.t90 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X59 a_2490_n1395# mux_4x1_1.mux_2x1_1.I1 VSS.t54 VSS.t53 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X60 mux_4x1_1.mux_2x1_0.nand2_2.IN2 S0.t11 VSS.t38 VSS.t37 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X61 mux_4x1_1.mux_2x1_0.nand2_2.OUT mux_4x1_1.mux_2x1_0.nand2_2.IN2 VDD.t58 VDD.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X62 mux_2x1_0.nand2_2.IN2 S2.t1 VDD.t30 VDD.t29 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X63 VDD mux_2x1_0.nand2_2.OUT OUT.t0 VDD.t5 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X64 mux_4x1_1.mux_2x1_2.nand2_2.OUT I0.t0 a_801_n795# VSS.t5 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X65 OUT mux_2x1_0.nand2_1.IN2 VDD.t9 VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X66 mux_4x1_1.mux_2x1_1.nand2_1.IN2 mux_4x1_1.mux_2x1_1.I1 VDD.t77 VDD.t76 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X67 VDD I2.t1 mux_4x1_1.mux_2x1_0.nand2_2.OUT VDD.t24 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X68 mux_4x1_0.mux_2x1_0.nand2_1.IN2 S0.t12 a_1364_1307# VSS.t15 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X69 mux_4x1_1.mux_2x1_0.nand2_1.IN2 S0.t13 a_1364_n1395# VSS.t16 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X70 mux_4x1_1.mux_2x1_1.I0 mux_4x1_1.mux_2x1_2.nand2_2.OUT a_801_n1395# VSS.t5 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X71 a_1364_1307# I7.t1 VSS.t44 VSS.t43 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X72 a_3053_1307# mux_4x1_0.mux_2x1_1.nand2_1.IN2 VSS.t50 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X73 VDD S0.t14 mux_4x1_1.mux_2x1_0.nand2_1.IN2 VDD.t10 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X74 VDD mux_4x1_1.mux_2x1_2.nand2_2.OUT mux_4x1_1.mux_2x1_1.I0 VDD.t59 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X75 mux_4x1_0.mux_2x1_2.nand2_2.OUT mux_4x1_0.mux_2x1_2.nand2_2.IN2 VDD.t37 VDD.t36 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X76 a_801_1307# mux_4x1_0.mux_2x1_2.nand2_1.IN2 VSS.t47 VSS.t23 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X77 a_3053_n1395# mux_4x1_1.mux_2x1_1.nand2_1.IN2 VSS.t59 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X78 a_801_707# mux_4x1_0.mux_2x1_2.nand2_2.IN2 VSS.t24 VSS.t23 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X79 mux_2x1_0.I1 mux_4x1_0.mux_2x1_1.nand2_2.OUT a_3053_1307# VSS.t13 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X80 VDD S2.t2 mux_2x1_0.nand2_1.IN2 VDD.t108 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 mux_4x1_0.mux_2x1_1.nand2_2.IN2 S1.t7 VSS.t36 VSS.t35 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X82 a_238_1307# I5.t1 VSS.t34 VSS.t33 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X83 mux_4x1_0.mux_2x1_0.nand2_2.IN2 S0.t15 VSS.t9 VSS.t8 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X84 OUT mux_2x1_0.nand2_2.OUT a_4178_1307# VSS.t4 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X85 mux_2x1_0.I0 mux_4x1_1.mux_2x1_1.nand2_1.IN2 VDD.t100 VDD.t99 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X86 mux_4x1_1.mux_2x1_1.I1 mux_4x1_1.mux_2x1_0.nand2_2.OUT a_1927_n1395# VSS.t10 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X87 a_3053_n795# mux_4x1_1.mux_2x1_1.nand2_2.IN2 VSS.t20 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X88 a_4178_1307# mux_2x1_0.nand2_1.IN2 VSS.t7 VSS.t6 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X89 VDD I0.t1 mux_4x1_1.mux_2x1_2.nand2_2.OUT VDD.t69 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X90 mux_2x1_0.nand2_2.IN2 S2.t3 VSS.t31 VSS.t30 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X91 a_801_n1395# mux_4x1_1.mux_2x1_2.nand2_1.IN2 VSS.t26 VSS.t25 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X92 a_801_n795# mux_4x1_1.mux_2x1_2.nand2_2.IN2 VSS.t27 VSS.t25 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X93 mux_4x1_1.mux_2x1_1.nand2_2.OUT mux_4x1_1.mux_2x1_1.I0 a_3053_n795# VSS.t56 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X94 mux_2x1_0.nand2_2.OUT mux_2x1_0.nand2_2.IN2 VDD.t102 VDD.t101 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X95 VDD mux_4x1_1.mux_2x1_0.nand2_2.OUT mux_4x1_1.mux_2x1_1.I1 VDD.t13 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X96 a_4178_707# mux_2x1_0.nand2_2.IN2 VSS.t60 VSS.t6 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X97 mux_4x1_1.mux_2x1_1.I0 mux_4x1_1.mux_2x1_2.nand2_1.IN2 VDD.t39 VDD.t38 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 VDD.t97 VDD.n83 40818.4
R1 VDD.n12 VDD.t43 40818.4
R2 VDD.t56 VDD.n4 40818.4
R3 VDD.t108 VDD.t8 763.259
R4 VDD.t0 VDD.t74 763.259
R5 VDD.t50 VDD.t103 763.259
R6 VDD.t16 VDD.t41 763.259
R7 VDD.t53 VDD.t48 763.259
R8 VDD.t66 VDD.t72 763.259
R9 VDD.t99 VDD.t80 763.259
R10 VDD.t13 VDD.t76 763.259
R11 VDD.t83 VDD.t10 763.259
R12 VDD.t59 VDD.t22 763.259
R13 VDD.t45 VDD.t38 763.259
R14 VDD.t19 VDD.t3 761.365
R15 VDD.n76 VDD.t101 386.348
R16 VDD.n84 VDD.t97 365.673
R17 VDD.n15 VDD.t43 365.673
R18 VDD.n5 VDD.t56 365.673
R19 VDD.n76 VDD.t29 362.409
R20 VDD.n81 VDD.t78 360.012
R21 VDD.n13 VDD.t95 360.012
R22 VDD.n3 VDD.t64 360.012
R23 VDD.n92 VDD.n84 322.221
R24 VDD.n15 VDD.n14 322.221
R25 VDD.n125 VDD.n5 322.221
R26 VDD.n77 VDD.n76 319.75
R27 VDD.n85 VDD.n84 319.733
R28 VDD.n16 VDD.n15 319.733
R29 VDD.n6 VDD.n5 319.733
R30 VDD.n33 VDD.t5 193.183
R31 VDD.n34 VDD.t108 193.183
R32 VDD.n36 VDD.t19 193.183
R33 VDD.n39 VDD.t0 193.183
R34 VDD.n41 VDD.t50 193.183
R35 VDD.n43 VDD.t16 193.183
R36 VDD.n45 VDD.t53 193.183
R37 VDD.n48 VDD.t66 193.183
R38 VDD.n75 VDD.t92 193.183
R39 VDD.n24 VDD.t87 193.183
R40 VDD.n103 VDD.t80 193.183
R41 VDD.n104 VDD.t13 193.183
R42 VDD.n112 VDD.t10 193.183
R43 VDD.n113 VDD.t59 193.183
R44 VDD.n114 VDD.t45 193.183
R45 VDD.n83 VDD.t31 192.236
R46 VDD.n12 VDD.t36 192.236
R47 VDD.n4 VDD.t34 192.236
R48 VDD.t8 VDD.n33 109.849
R49 VDD.t3 VDD.n34 109.849
R50 VDD.t74 VDD.n36 109.849
R51 VDD.t103 VDD.n39 109.849
R52 VDD.t41 VDD.n41 109.849
R53 VDD.t48 VDD.n43 109.849
R54 VDD.t72 VDD.n45 109.849
R55 VDD.n48 VDD.t90 109.849
R56 VDD.t101 VDD.n75 109.849
R57 VDD.n24 VDD.t99 109.849
R58 VDD.t76 VDD.n103 109.849
R59 VDD.n104 VDD.t83 109.849
R60 VDD.t22 VDD.n112 109.849
R61 VDD.t38 VDD.n113 109.849
R62 VDD.n114 VDD.t27 109.849
R63 VDD.n82 VDD.t105 96.5914
R64 VDD.n10 VDD.t69 96.5914
R65 VDD.n0 VDD.t24 96.5914
R66 VDD.t31 VDD.n82 54.9247
R67 VDD.t36 VDD.n10 54.9247
R68 VDD.t34 VDD.n0 54.9247
R69 VDD.n93 VDD 18.0631
R70 VDD.n73 VDD 11.7877
R71 VDD.n115 VDD.n114 6.3005
R72 VDD.n113 VDD.n18 6.3005
R73 VDD.n112 VDD.n111 6.3005
R74 VDD.n105 VDD.n104 6.3005
R75 VDD.n103 VDD.n102 6.3005
R76 VDD.n25 VDD.n24 6.3005
R77 VDD.n75 VDD.n74 6.3005
R78 VDD.n33 VDD.n31 6.3005
R79 VDD.n68 VDD.n34 6.3005
R80 VDD.n65 VDD.n36 6.3005
R81 VDD.n62 VDD.n39 6.3005
R82 VDD.n59 VDD.n41 6.3005
R83 VDD.n55 VDD.n43 6.3005
R84 VDD.n52 VDD.n45 6.3005
R85 VDD.n49 VDD.n48 6.3005
R86 VDD VDD.n23 5.23855
R87 VDD VDD.n30 5.23855
R88 VDD VDD.n29 5.23796
R89 VDD.n49 VDD.t91 5.21701
R90 VDD.n115 VDD.t28 5.21701
R91 VDD.n16 VDD.t44 5.19258
R92 VDD.n14 VDD.t96 5.19258
R93 VDD.n78 VDD.t30 5.1858
R94 VDD.n86 VDD.t98 5.14703
R95 VDD.n91 VDD.t79 5.14703
R96 VDD.n124 VDD.t65 5.14703
R97 VDD.n7 VDD.t57 5.14703
R98 VDD.n54 VDD.t49 5.13746
R99 VDD.n61 VDD.t104 5.13746
R100 VDD.n67 VDD.t4 5.13746
R101 VDD.n101 VDD.t77 5.13746
R102 VDD.n110 VDD.t23 5.13746
R103 VDD.n89 VDD.n87 5.13287
R104 VDD.n89 VDD.n88 5.13287
R105 VDD.n50 VDD.n47 5.13287
R106 VDD.n53 VDD.n44 5.13287
R107 VDD.n56 VDD.n42 5.13287
R108 VDD.n60 VDD.n40 5.13287
R109 VDD.n63 VDD.n38 5.13287
R110 VDD.n66 VDD.n35 5.13287
R111 VDD.n69 VDD.n32 5.13287
R112 VDD.n79 VDD.n27 5.13287
R113 VDD.n79 VDD.n28 5.13287
R114 VDD.n98 VDD.n22 5.13287
R115 VDD.n100 VDD.n99 5.13287
R116 VDD.n107 VDD.n20 5.13287
R117 VDD.n109 VDD.n108 5.13287
R118 VDD.n122 VDD.n8 5.13287
R119 VDD.n122 VDD.n9 5.13287
R120 VDD.n116 VDD.n19 5.13287
R121 VDD.n46 VDD.t73 3.91303
R122 VDD.n37 VDD.t75 3.91303
R123 VDD.n57 VDD.t42 3.91303
R124 VDD.n71 VDD.t9 3.91303
R125 VDD.n21 VDD.t84 3.9128
R126 VDD.n118 VDD.t39 3.9128
R127 VDD.n96 VDD.t100 3.91277
R128 VDD.n96 VDD.n95 3.87701
R129 VDD.n119 VDD.n118 3.87649
R130 VDD.n46 VDD.n11 3.87623
R131 VDD.n37 VDD.n26 3.87623
R132 VDD.n57 VDD.n1 3.87623
R133 VDD.n21 VDD.n2 3.87585
R134 VDD.n72 VDD.n71 3.87523
R135 VDD.n1 VDD.t35 3.51093
R136 VDD.n72 VDD.t102 3.51093
R137 VDD.n11 VDD.t37 3.51093
R138 VDD.n26 VDD.t32 3.51093
R139 VDD.n119 VDD.t40 3.51079
R140 VDD.n95 VDD.t33 3.51063
R141 VDD.n2 VDD.t58 3.51063
R142 VDD.n79 VDD.n78 3.45802
R143 VDD.n82 VDD.n80 3.15287
R144 VDD.n121 VDD.n10 3.1505
R145 VDD.n128 VDD.n0 3.1505
R146 VDD.n83 VDD.n81 0.939698
R147 VDD.n13 VDD.n12 0.939698
R148 VDD.n4 VDD.n3 0.939698
R149 VDD.n17 VDD 0.412255
R150 VDD.n126 VDD 0.412255
R151 VDD.n126 VDD 0.412255
R152 VDD.n93 VDD 0.411896
R153 VDD.n17 VDD 0.411255
R154 VDD.n120 VDD.n119 0.274239
R155 VDD.n95 VDD.n94 0.273886
R156 VDD.n127 VDD.n2 0.273886
R157 VDD.n120 VDD.n11 0.272927
R158 VDD.n94 VDD.n26 0.272927
R159 VDD.n73 VDD.n72 0.272927
R160 VDD.n127 VDD.n1 0.272927
R161 VDD.n51 VDD.n46 0.22389
R162 VDD.n64 VDD.n37 0.22389
R163 VDD.n71 VDD.n70 0.22389
R164 VDD.n58 VDD.n57 0.22389
R165 VDD.n106 VDD.n21 0.22353
R166 VDD.n118 VDD.n117 0.22353
R167 VDD.n97 VDD.n96 0.223424
R168 VDD.n90 VDD.n86 0.176707
R169 VDD.n91 VDD.n90 0.143461
R170 VDD.n98 VDD.n97 0.141016
R171 VDD.n101 VDD.n100 0.141016
R172 VDD.n107 VDD.n106 0.141016
R173 VDD.n110 VDD.n109 0.141016
R174 VDD.n117 VDD.n116 0.141016
R175 VDD.n70 VDD.n69 0.141016
R176 VDD.n64 VDD.n63 0.141016
R177 VDD.n61 VDD.n60 0.141016
R178 VDD.n58 VDD.n56 0.141016
R179 VDD.n54 VDD.n53 0.141016
R180 VDD.n51 VDD.n50 0.141016
R181 VDD.n67 VDD.n66 0.140435
R182 VDD.n123 VDD.n7 0.139013
R183 VDD.n124 VDD.n123 0.139013
R184 VDD VDD.n98 0.106177
R185 VDD.n100 VDD 0.106177
R186 VDD VDD.n107 0.106177
R187 VDD.n109 VDD 0.106177
R188 VDD.n116 VDD 0.106177
R189 VDD.n69 VDD 0.106177
R190 VDD.n66 VDD 0.106177
R191 VDD.n63 VDD 0.106177
R192 VDD.n60 VDD 0.106177
R193 VDD.n56 VDD 0.106177
R194 VDD.n53 VDD 0.106177
R195 VDD.n50 VDD 0.106177
R196 VDD.n97 VDD.n25 0.0800484
R197 VDD.n102 VDD.n101 0.0800484
R198 VDD.n106 VDD.n105 0.0800484
R199 VDD.n117 VDD.n18 0.0800484
R200 VDD.n74 VDD.n73 0.0800484
R201 VDD.n70 VDD.n31 0.0800484
R202 VDD.n68 VDD.n67 0.0800484
R203 VDD.n65 VDD.n64 0.0800484
R204 VDD.n62 VDD.n61 0.0800484
R205 VDD.n59 VDD.n58 0.0800484
R206 VDD.n52 VDD.n51 0.0800484
R207 VDD VDD.n110 0.0788871
R208 VDD VDD.n54 0.0788871
R209 VDD.n122 VDD 0.0530484
R210 VDD VDD.n79 0.0530484
R211 VDD.n89 VDD 0.0513065
R212 VDD.n86 VDD.n85 0.0460556
R213 VDD.n92 VDD.n91 0.0460556
R214 VDD.n7 VDD.n6 0.0460556
R215 VDD.n125 VDD.n124 0.0460556
R216 VDD.n121 VDD.n120 0.0402742
R217 VDD.n94 VDD.n80 0.0402742
R218 VDD.n128 VDD.n127 0.0402742
R219 VDD.n123 VDD.n122 0.0338871
R220 VDD.n90 VDD.n89 0.0318548
R221 VDD.n94 VDD.n93 0.0239437
R222 VDD.n120 VDD.n17 0.0225645
R223 VDD.n127 VDD.n126 0.0225645
R224 VDD.n84 VDD.n81 0.00925055
R225 VDD.n15 VDD.n13 0.00925055
R226 VDD.n5 VDD.n3 0.00925055
R227 VDD.n78 VDD.n77 0.00883333
R228 VDD.n25 VDD 0.00166129
R229 VDD.n102 VDD 0.00166129
R230 VDD.n105 VDD 0.00166129
R231 VDD.n111 VDD 0.00166129
R232 VDD.n111 VDD 0.00166129
R233 VDD VDD.n18 0.00166129
R234 VDD VDD.n115 0.00166129
R235 VDD.n74 VDD 0.00166129
R236 VDD.n31 VDD 0.00166129
R237 VDD VDD.n68 0.00166129
R238 VDD VDD.n65 0.00166129
R239 VDD VDD.n62 0.00166129
R240 VDD VDD.n59 0.00166129
R241 VDD VDD.n55 0.00166129
R242 VDD.n55 VDD 0.00166129
R243 VDD VDD.n52 0.00166129
R244 VDD VDD.n49 0.00166129
R245 VDD VDD.n121 0.00108064
R246 VDD.n80 VDD 0.00108064
R247 VDD VDD.n128 0.00108064
R248 VDD.n85 VDD 0.00105556
R249 VDD VDD.n92 0.00105556
R250 VDD.n14 VDD 0.00105556
R251 VDD VDD.n16 0.00105556
R252 VDD.n6 VDD 0.00105556
R253 VDD VDD.n125 0.00105556
R254 VDD.n77 VDD 0.00105556
R255 S2.n1 S2.t0 31.528
R256 S2.n0 S2.t1 25.7638
R257 S2.n1 S2.t2 15.3826
R258 S2.n0 S2.t3 13.2969
R259 S2.n2 S2.n1 7.62851
R260 S2.n7 S2.n4 2.2505
R261 S2.n3 S2.n2 2.2324
R262 S2.n7 S2.n0 2.11815
R263 S2.n2 S2 0.107918
R264 S2.n4 S2.n3 0.0289694
R265 S2 S2.n5 0.0124388
R266 S2.n7 S2.n6 0.00421134
R267 S2.n5 S2.n4 0.00417347
R268 S2.n6 S2 0.00235567
R269 S2 S2.n7 0.00142783
R270 VSS.n37 VSS.n36 28802.9
R271 VSS.t33 VSS.t48 23952.8
R272 VSS.t56 VSS.n25 21804.7
R273 VSS.t53 VSS.t10 1483.3
R274 VSS.t45 VSS.t16 1483.3
R275 VSS.t51 VSS.t5 1483.3
R276 VSS.t25 VSS.t57 1483.3
R277 VSS.t32 VSS.t6 1483.3
R278 VSS.t17 VSS.t58 1483.3
R279 VSS.t43 VSS.t29 1483.3
R280 VSS.t41 VSS.t23 1483.3
R281 VSS.t2 VSS.t13 1479.61
R282 VSS.t42 VSS.t19 1367.44
R283 VSS.n13 VSS.t4 353.341
R284 VSS.n36 VSS.n35 349.661
R285 VSS.n58 VSS.n57 349.661
R286 VSS.n38 VSS.n37 349.661
R287 VSS.n47 VSS.n6 349.661
R288 VSS.n25 VSS.n24 345.981
R289 VSS.n27 VSS.t56 298.279
R290 VSS.n29 VSS.t53 235.561
R291 VSS.n35 VSS.t45 235.561
R292 VSS.n59 VSS.t51 235.561
R293 VSS.n57 VSS.t25 235.561
R294 VSS.t48 VSS.n49 235.561
R295 VSS.t6 VSS.n13 235.561
R296 VSS.n15 VSS.t2 235.561
R297 VSS.n24 VSS.t17 235.561
R298 VSS.n18 VSS.t61 235.561
R299 VSS.n38 VSS.t21 235.561
R300 VSS.n43 VSS.t43 235.561
R301 VSS.t23 VSS.n47 235.561
R302 VSS.n50 VSS.t33 235.561
R303 VSS.t19 VSS.n27 198.853
R304 VSS.n54 VSS.t12 9.34566
R305 VSS.n10 VSS.t31 9.34566
R306 VSS.n21 VSS.t36 9.34566
R307 VSS.n40 VSS.t9 9.34566
R308 VSS.n4 VSS.t40 9.34566
R309 VSS.n8 VSS.t1 9.34566
R310 VSS.n32 VSS.t38 9.34566
R311 VSS.n25 VSS.t13 7.36177
R312 VSS.n3 VSS.t27 7.19156
R313 VSS.n3 VSS.t26 7.19156
R314 VSS.n12 VSS.t7 7.19156
R315 VSS.n12 VSS.t60 7.19156
R316 VSS.n17 VSS.t3 7.19156
R317 VSS.n20 VSS.t50 7.19156
R318 VSS.n20 VSS.t18 7.19156
R319 VSS.n7 VSS.t62 7.19156
R320 VSS.n39 VSS.t28 7.19156
R321 VSS.n39 VSS.t22 7.19156
R322 VSS.n45 VSS.t44 7.19156
R323 VSS.n46 VSS.t47 7.19156
R324 VSS.n46 VSS.t24 7.19156
R325 VSS.n52 VSS.t34 7.19156
R326 VSS.n53 VSS.t49 7.19156
R327 VSS.n26 VSS.t20 7.19156
R328 VSS.n26 VSS.t59 7.19156
R329 VSS.n31 VSS.t54 7.19156
R330 VSS.n34 VSS.t46 7.19156
R331 VSS.n34 VSS.t55 7.19156
R332 VSS.n0 VSS.t52 7.19156
R333 VSS.t0 VSS.t42 3.68113
R334 VSS.n36 VSS.t10 3.68113
R335 VSS.t16 VSS.t37 3.68113
R336 VSS.t5 VSS.n58 3.68113
R337 VSS.t57 VSS.t11 3.68113
R338 VSS.t30 VSS.t32 3.68113
R339 VSS.t58 VSS.t35 3.68113
R340 VSS.n37 VSS.t14 3.68113
R341 VSS.t8 VSS.t15 3.68113
R342 VSS.t29 VSS.n6 3.68113
R343 VSS.t39 VSS.t41 3.68113
R344 VSS.n60 VSS.n1 3.37613
R345 VSS.n30 VSS.n28 3.37613
R346 VSS.n16 VSS.n14 3.37613
R347 VSS.n23 VSS.n19 3.37613
R348 VSS.n44 VSS.n42 3.37613
R349 VSS.n51 VSS.n48 3.37613
R350 VSS.n56 VSS.n2 3.37613
R351 VSS.n57 VSS 2.6035
R352 VSS.n47 VSS 2.6035
R353 VSS VSS.n38 2.6035
R354 VSS.n24 VSS 2.6035
R355 VSS.n13 VSS 2.6035
R356 VSS.n35 VSS 2.6035
R357 VSS.n27 VSS 2.60269
R358 VSS.n56 VSS.n55 2.6005
R359 VSS.t11 VSS.n56 2.6005
R360 VSS VSS.n2 2.6005
R361 VSS.n49 VSS.n2 2.6005
R362 VSS VSS.n51 2.6005
R363 VSS.n51 VSS.n50 2.6005
R364 VSS VSS.n44 2.6005
R365 VSS.n44 VSS.n43 2.6005
R366 VSS VSS.n19 2.6005
R367 VSS.n19 VSS.n18 2.6005
R368 VSS VSS.n16 2.6005
R369 VSS.n16 VSS.n15 2.6005
R370 VSS.n14 VSS.n11 2.6005
R371 VSS.n14 VSS.t30 2.6005
R372 VSS.n23 VSS.n22 2.6005
R373 VSS.t35 VSS.n23 2.6005
R374 VSS.n42 VSS.n41 2.6005
R375 VSS.n42 VSS.t8 2.6005
R376 VSS.n48 VSS.n5 2.6005
R377 VSS.n48 VSS.t39 2.6005
R378 VSS.n28 VSS.n9 2.6005
R379 VSS.n28 VSS.t0 2.6005
R380 VSS VSS.n30 2.6005
R381 VSS.n30 VSS.n29 2.6005
R382 VSS.n33 VSS.n1 2.6005
R383 VSS.t37 VSS.n1 2.6005
R384 VSS VSS.n60 2.6005
R385 VSS.n60 VSS.n59 2.6005
R386 VSS.n53 VSS.n52 2.54306
R387 VSS VSS.n0 0.171522
R388 VSS VSS.n7 0.171522
R389 VSS VSS.n45 0.171522
R390 VSS VSS.n31 0.171522
R391 VSS VSS.n17 0.17111
R392 VSS VSS.n3 0.113253
R393 VSS.n12 VSS 0.113253
R394 VSS VSS.n20 0.113253
R395 VSS VSS.n39 0.113253
R396 VSS.n46 VSS 0.113253
R397 VSS.n26 VSS 0.113253
R398 VSS.n34 VSS 0.113253
R399 VSS.n3 VSS 0.0595367
R400 VSS VSS.n12 0.0595367
R401 VSS.n20 VSS 0.0595367
R402 VSS.n39 VSS 0.0595367
R403 VSS VSS.n46 0.0595367
R404 VSS VSS.n26 0.0595367
R405 VSS VSS.n34 0.0595367
R406 VSS.n17 VSS 0.0569474
R407 VSS VSS.n7 0.0569474
R408 VSS.n45 VSS 0.0569474
R409 VSS.n52 VSS 0.0569474
R410 VSS VSS.n53 0.0569474
R411 VSS.n31 VSS 0.0569474
R412 VSS VSS.n0 0.0569474
R413 VSS VSS.n10 0.0340526
R414 VSS VSS.n21 0.0340526
R415 VSS VSS.n40 0.0340526
R416 VSS VSS.n4 0.0340526
R417 VSS VSS.n54 0.0340526
R418 VSS VSS.n8 0.0340526
R419 VSS VSS.n32 0.0320789
R420 VSS VSS.n11 0.0182632
R421 VSS.n22 VSS 0.0182632
R422 VSS.n41 VSS 0.0182632
R423 VSS VSS.n5 0.0182632
R424 VSS.n55 VSS 0.0182632
R425 VSS VSS.n9 0.0182632
R426 VSS VSS.n33 0.0182632
R427 VSS VSS.n10 0.00405263
R428 VSS.n21 VSS 0.00405263
R429 VSS VSS.n4 0.00405263
R430 VSS.n54 VSS 0.00405263
R431 VSS VSS.n8 0.00405263
R432 VSS.n40 VSS 0.00247368
R433 VSS.n32 VSS 0.00247368
R434 VSS.n11 VSS 0.000894737
R435 VSS.n22 VSS 0.000894737
R436 VSS.n41 VSS 0.000894737
R437 VSS.n5 VSS 0.000894737
R438 VSS.n55 VSS 0.000894737
R439 VSS.n9 VSS 0.000894737
R440 VSS.n33 VSS 0.000894737
R441 S1.n0 S1.t5 31.528
R442 S1.n5 S1.t0 31.528
R443 S1.n16 S1.t6 25.7638
R444 S1.n3 S1.t1 25.7638
R445 S1.n0 S1.t3 15.3826
R446 S1.n5 S1.t2 15.3826
R447 S1.n16 S1.t7 13.2969
R448 S1.n3 S1.t4 13.2969
R449 S1.n21 S1.n0 7.62076
R450 S1.n6 S1.n5 7.62076
R451 S1.n14 S1.n13 6.87179
R452 S1.n8 S1.n7 4.54699
R453 S1.n20 S1.n19 4.54699
R454 S1.n15 S1.n14 4.52926
R455 S1.n13 S1.n12 4.52926
R456 S1.n18 S1 4.52833
R457 S1.n9 S1 4.52833
R458 S1.n11 S1.n10 2.2505
R459 S1.n17 S1.n1 2.2505
R460 S1.n17 S1.n16 2.11815
R461 S1.n11 S1.n3 2.11815
R462 S1.n9 S1.n8 1.33991
R463 S1.n20 S1.n18 1.33848
R464 S1.n8 S1.n6 1.12145
R465 S1.n21 S1.n20 1.12145
R466 S1.n7 S1 0.0780197
R467 S1.n19 S1 0.0780197
R468 S1.n7 S1 0.0359098
R469 S1.n19 S1 0.032959
R470 S1.n10 S1.n9 0.0289694
R471 S1.n18 S1.n1 0.0289694
R472 S1.n14 S1 0.0170306
R473 S1.n13 S1 0.0161122
R474 S1.n4 S1 0.0133571
R475 S1 S1.n2 0.0124388
R476 S1.n17 S1.n15 0.00421134
R477 S1.n2 S1.n1 0.00417347
R478 S1.n12 S1.n11 0.00328351
R479 S1.n10 S1.n4 0.0032551
R480 S1 S1.n6 0.00197541
R481 S1 S1.n21 0.00197541
R482 S1 S1.n17 0.00142783
R483 S1.n11 S1 0.00142783
R484 S0.n0 S0.t9 31.528
R485 S0.n21 S0.t1 31.528
R486 S0.n13 S0.t13 31.528
R487 S0.n2 S0.t12 31.528
R488 S0.n33 S0.t2 25.7638
R489 S0.n11 S0.t0 25.7638
R490 S0.n16 S0.t4 25.7638
R491 S0.n5 S0.t10 25.7638
R492 S0.n0 S0.t5 15.3826
R493 S0.n21 S0.t3 15.3826
R494 S0.n13 S0.t14 15.3826
R495 S0.n2 S0.t7 15.3826
R496 S0.n33 S0.t8 13.2969
R497 S0.n11 S0.t6 13.2969
R498 S0.n16 S0.t11 13.2969
R499 S0.n5 S0.t15 13.2969
R500 S0.n14 S0.n13 7.6291
R501 S0.n3 S0.n2 7.6289
R502 S0.n1 S0.n0 7.62076
R503 S0.n22 S0.n21 7.62076
R504 S0.n20 S0 4.53443
R505 S0.n39 S0 4.53443
R506 S0.n32 S0.n31 4.52926
R507 S0.n30 S0.n29 4.52926
R508 S0.n36 S0 4.52853
R509 S0.n35 S0 4.52833
R510 S0.n26 S0 4.52833
R511 S0.n18 S0 4.52833
R512 S0.n7 S0 4.52833
R513 S0.n28 S0.n27 2.2505
R514 S0.n34 S0.n9 2.2505
R515 S0.n37 S0.n8 2.19776
R516 S0.n24 S0.n19 2.19633
R517 S0.n34 S0.n33 2.11815
R518 S0.n28 S0.n11 2.11815
R519 S0.n17 S0.n16 2.11815
R520 S0.n6 S0.n5 2.11815
R521 S0.n31 S0.n30 1.84791
R522 S0.n23 S0.n22 1.5005
R523 S0.n38 S0.n1 1.5005
R524 S0.n26 S0.n25 1.31185
R525 S0.n36 S0.n35 1.31042
R526 S0.n19 S0.n18 1.2853
R527 S0.n8 S0.n7 1.28387
R528 S0.n6 S0.n4 1.1266
R529 S0.n17 S0.n15 1.12637
R530 S0.n8 S0.n3 0.948428
R531 S0.n19 S0.n14 0.948389
R532 S0.n14 S0 0.109321
R533 S0.n3 S0 0.108522
R534 S0 S0.n39 0.0780742
R535 S0.n20 S0 0.0780197
R536 S0.n22 S0.n20 0.0373852
R537 S0.n39 S0.n1 0.0373852
R538 S0.n25 S0.n24 0.0359098
R539 S0.n37 S0.n36 0.0359098
R540 S0.n7 S0.n4 0.0344967
R541 S0.n18 S0.n15 0.0342688
R542 S0.n27 S0.n26 0.0289694
R543 S0.n35 S0.n9 0.0289694
R544 S0.n31 S0 0.0170306
R545 S0.n30 S0 0.0161122
R546 S0.n12 S0 0.0133571
R547 S0.n15 S0 0.012774
R548 S0.n4 S0 0.0125466
R549 S0 S0.n10 0.0124388
R550 S0 S0.n1 0.00935246
R551 S0.n34 S0.n32 0.00421134
R552 S0.n10 S0.n9 0.00417347
R553 S0.n23 S0 0.00345082
R554 S0 S0.n38 0.00345082
R555 S0.n29 S0.n28 0.00328351
R556 S0.n27 S0.n12 0.0032551
R557 S0.n24 S0.n23 0.00197541
R558 S0.n38 S0.n37 0.00197541
R559 S0 S0.n34 0.00142783
R560 S0.n28 S0 0.00142783
R561 S0 S0.n17 0.00142783
R562 S0 S0.n6 0.00142783
R563 I4.n0 I4.t1 31.528
R564 I4.n0 I4.t0 15.3826
R565 I4 I4.n0 8.74076
R566 I3.n0 I3.t1 30.9379
R567 I3.n0 I3.t0 21.6422
R568 I3 I3.n0 4.0005
R569 I6.n0 I6.t1 31.528
R570 I6.n0 I6.t0 15.3826
R571 I6.n1 I6.n0 8.74076
R572 I6.n1 I6 0.00507627
R573 I6 I6.n1 0.00202542
R574 I1.n0 I1.t1 30.9379
R575 I1.n0 I1.t0 21.6422
R576 I1 I1.n0 4.005
R577 I2.n0 I2.t0 31.528
R578 I2.n0 I2.t1 15.3826
R579 I2.n1 I2.n0 8.74076
R580 I2.n1 I2 0.00197541
R581 I2 I2.n1 0.00197541
R582 I7.n0 I7.t0 30.9379
R583 I7.n0 I7.t1 21.6422
R584 I7 I7.n0 4.0005
R585 I5.n0 I5.t0 30.9379
R586 I5.n0 I5.t1 21.6422
R587 I5 I5.n0 4.005
R588 OUT OUT.n2 7.15141
R589 OUT.n3 OUT.n1 3.2163
R590 OUT.n1 OUT.t0 2.2755
R591 OUT.n1 OUT.n0 2.2755
R592 OUT OUT.n3 0.035398
R593 OUT.n3 OUT 0.0119545
R594 I0.n0 I0.t0 31.528
R595 I0.n0 I0.t1 15.3826
R596 I0 I0.n0 8.74076
C0 mux_4x1_0.mux_2x1_1.I0 S0 0.207f
C1 mux_4x1_1.mux_2x1_1.nand2_1.IN2 mux_4x1_1.mux_2x1_1.I0 0.00154f
C2 mux_2x1_0.I1 VDD 0.423f
C3 mux_4x1_1.mux_2x1_1.nand2_2.OUT mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.12f
C4 mux_4x1_1.mux_2x1_2.nand2_2.OUT a_801_n795# 0.0964f
C5 mux_4x1_1.mux_2x1_2.nand2_2.OUT I4 3e-19
C6 mux_4x1_1.mux_2x1_1.I1 mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.328f
C7 mux_2x1_0.nand2_2.OUT S1 1.54e-19
C8 mux_4x1_1.mux_2x1_0.nand2_1.IN2 mux_4x1_1.mux_2x1_0.nand2_2.IN2 0.00212f
C9 mux_4x1_1.mux_2x1_1.I0 a_801_n795# 1.5e-19
C10 mux_4x1_0.mux_2x1_0.nand2_2.OUT mux_4x1_0.mux_2x1_1.I1 0.328f
C11 mux_4x1_1.mux_2x1_1.I0 mux_4x1_0.mux_2x1_0.nand2_2.IN2 9.55e-20
C12 S1 mux_4x1_0.mux_2x1_0.nand2_1.IN2 4.51e-21
C13 mux_4x1_1.mux_2x1_1.I1 mux_4x1_1.mux_2x1_1.I0 0.00147f
C14 mux_4x1_0.mux_2x1_1.I1 mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.11f
C15 mux_2x1_0.I1 mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.329f
C16 mux_4x1_1.mux_2x1_2.nand2_1.IN2 I1 0.0959f
C17 I6 mux_4x1_1.mux_2x1_1.I0 1.04e-19
C18 I4 a_801_707# 0.00293f
C19 a_4178_1307# mux_2x1_0.nand2_1.IN2 0.00372f
C20 I7 S0 0.0665f
C21 mux_4x1_0.mux_2x1_2.nand2_2.IN2 I4 0.0473f
C22 S1 S2 0.0018f
C23 mux_4x1_0.mux_2x1_1.I1 S0 0.0109f
C24 VDD mux_4x1_0.mux_2x1_1.nand2_2.IN2 0.405f
C25 mux_4x1_0.mux_2x1_2.nand2_1.IN2 I5 0.0959f
C26 a_1364_n1395# VDD 3.14e-19
C27 mux_2x1_0.nand2_2.IN2 mux_2x1_0.nand2_1.IN2 0.00212f
C28 a_3053_n795# VDD 0.00444f
C29 a_801_n1395# VDD 0.00444f
C30 mux_4x1_0.mux_2x1_0.nand2_2.OUT VDD 0.665f
C31 a_1927_n795# VDD 0.00444f
C32 mux_4x1_0.mux_2x1_1.nand2_2.IN2 mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.12f
C33 a_801_1307# mux_4x1_0.mux_2x1_2.nand2_2.OUT 0.00949f
C34 a_3053_707# S2 2.16e-19
C35 mux_2x1_0.I1 a_3053_1307# 0.069f
C36 VDD mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.462f
C37 mux_2x1_0.I0 S0 6.5e-20
C38 a_801_1307# mux_4x1_0.mux_2x1_1.I0 0.069f
C39 mux_4x1_0.mux_2x1_0.nand2_2.OUT a_1927_707# 0.0964f
C40 OUT mux_2x1_0.nand2_2.OUT 0.303f
C41 I2 S1 0.00826f
C42 mux_4x1_1.mux_2x1_2.nand2_2.IN2 VDD 0.404f
C43 mux_2x1_0.nand2_1.IN2 VDD 0.461f
C44 VDD S0 3.48f
C45 mux_2x1_0.I0 mux_4x1_1.mux_2x1_1.nand2_2.OUT 0.419f
C46 a_238_1307# mux_4x1_0.mux_2x1_2.nand2_1.IN2 0.069f
C47 mux_4x1_0.mux_2x1_2.nand2_2.OUT mux_4x1_0.mux_2x1_1.I0 0.63f
C48 mux_4x1_0.mux_2x1_1.I0 mux_4x1_1.mux_2x1_1.nand2_2.IN2 9.55e-20
C49 mux_4x1_1.mux_2x1_0.nand2_2.IN2 mux_4x1_0.mux_2x1_1.I0 9.55e-20
C50 mux_4x1_0.mux_2x1_1.nand2_1.IN2 mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.053f
C51 mux_4x1_1.mux_2x1_1.nand2_2.OUT VDD 0.634f
C52 a_1927_707# S0 2.62e-19
C53 OUT S2 0.00946f
C54 mux_2x1_0.nand2_1.IN2 mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.0106f
C55 mux_4x1_1.mux_2x1_0.nand2_1.IN2 VDD 0.46f
C56 I6 mux_4x1_0.mux_2x1_1.nand2_2.IN2 0.0036f
C57 I2 mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.203f
C58 mux_4x1_0.mux_2x1_0.nand2_2.OUT mux_4x1_0.mux_2x1_0.nand2_2.IN2 0.12f
C59 a_238_n1395# VDD 3.14e-19
C60 mux_4x1_1.mux_2x1_1.nand2_1.IN2 S0 4.45e-19
C61 I2 mux_4x1_1.mux_2x1_1.I0 0.01f
C62 mux_2x1_0.I1 S2 0.0594f
C63 I7 mux_4x1_0.mux_2x1_2.nand2_2.OUT 0.0174f
C64 mux_4x1_1.mux_2x1_2.nand2_1.IN2 mux_4x1_1.mux_2x1_2.nand2_2.OUT 0.053f
C65 a_3053_707# S1 2.62e-19
C66 a_1927_1307# mux_4x1_0.mux_2x1_0.nand2_2.OUT 0.00949f
C67 I6 mux_4x1_0.mux_2x1_0.nand2_2.OUT 0.202f
C68 I3 VDD 0.153f
C69 S1 mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.113f
C70 mux_4x1_1.mux_2x1_2.nand2_2.IN2 a_801_n795# 0.00372f
C71 mux_4x1_1.mux_2x1_2.nand2_1.IN2 mux_4x1_1.mux_2x1_1.I0 0.109f
C72 a_801_n795# S0 6.89e-19
C73 a_3053_1307# mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.00372f
C74 mux_4x1_0.mux_2x1_0.nand2_2.OUT a_2490_1307# 9.43e-19
C75 I7 mux_4x1_0.mux_2x1_1.I0 0.0454f
C76 mux_4x1_0.mux_2x1_0.nand2_2.IN2 S0 0.136f
C77 mux_4x1_1.mux_2x1_1.nand2_1.IN2 mux_4x1_1.mux_2x1_1.nand2_2.OUT 0.053f
C78 I4 S0 0.00512f
C79 mux_4x1_0.mux_2x1_1.I1 mux_4x1_0.mux_2x1_1.I0 0.00147f
C80 S1 mux_4x1_1.mux_2x1_1.I0 0.0863f
C81 mux_4x1_1.mux_2x1_1.I1 S0 0.0109f
C82 a_2490_1307# mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.069f
C83 mux_2x1_0.nand2_2.IN2 mux_4x1_0.mux_2x1_1.I0 0.00494f
C84 mux_4x1_1.mux_2x1_2.nand2_2.OUT I0 0.202f
C85 a_1927_n1395# VDD 0.00444f
C86 a_801_1307# VDD 0.00444f
C87 mux_4x1_1.mux_2x1_1.I0 I0 0.0148f
C88 S2 mux_4x1_0.mux_2x1_1.nand2_2.IN2 3.66e-19
C89 mux_2x1_0.I0 mux_4x1_1.mux_2x1_1.nand2_2.IN2 3.43e-19
C90 mux_4x1_0.mux_2x1_0.nand2_1.IN2 mux_4x1_0.mux_2x1_0.nand2_2.OUT 0.053f
C91 a_1364_1307# S0 0.0151f
C92 a_3053_n1395# mux_4x1_1.mux_2x1_1.I0 2.44e-19
C93 mux_4x1_1.mux_2x1_0.nand2_1.IN2 mux_4x1_1.mux_2x1_1.I1 0.109f
C94 mux_4x1_0.mux_2x1_2.nand2_2.OUT VDD 0.664f
C95 VDD mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.405f
C96 mux_4x1_1.mux_2x1_0.nand2_2.IN2 VDD 0.405f
C97 a_3615_1307# VDD 3.14e-19
C98 I5 S0 0.0576f
C99 mux_2x1_0.I0 mux_4x1_0.mux_2x1_1.I0 0.0073f
C100 mux_4x1_1.mux_2x1_1.I0 mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.0241f
C101 mux_2x1_0.nand2_1.IN2 mux_2x1_0.nand2_2.OUT 0.053f
C102 mux_4x1_1.mux_2x1_2.nand2_2.OUT mux_4x1_1.mux_2x1_1.I0 0.63f
C103 S1 mux_2x1_0.I1 0.00946f
C104 VDD mux_4x1_0.mux_2x1_1.I0 1.41f
C105 mux_4x1_0.mux_2x1_0.nand2_1.IN2 S0 0.378f
C106 S2 mux_4x1_0.mux_2x1_1.nand2_1.IN2 4.52e-21
C107 a_3615_1307# mux_4x1_0.mux_2x1_1.nand2_2.OUT 9.46e-19
C108 mux_4x1_0.mux_2x1_2.nand2_1.IN2 mux_4x1_0.mux_2x1_2.nand2_2.IN2 0.00212f
C109 mux_2x1_0.nand2_1.IN2 S2 0.341f
C110 a_2490_n1395# VDD 3.14e-19
C111 a_1927_707# mux_4x1_0.mux_2x1_1.I0 8.2e-19
C112 I1 S0 0.0576f
C113 mux_4x1_0.mux_2x1_1.I0 mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.25f
C114 mux_4x1_1.mux_2x1_1.nand2_1.IN2 mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.00212f
C115 mux_4x1_1.mux_2x1_1.I1 a_1927_n1395# 0.069f
C116 I7 VDD 0.153f
C117 mux_2x1_0.I0 mux_2x1_0.nand2_2.IN2 0.051f
C118 S1 mux_4x1_0.mux_2x1_1.nand2_2.IN2 0.16f
C119 a_238_1307# S0 0.0144f
C120 a_4178_1307# VDD 0.00444f
C121 mux_4x1_0.mux_2x1_1.I1 VDD 0.423f
C122 a_1927_n795# I2 0.00293f
C123 mux_4x1_0.mux_2x1_2.nand2_2.IN2 a_801_707# 0.00372f
C124 mux_4x1_0.mux_2x1_2.nand2_2.OUT mux_4x1_0.mux_2x1_0.nand2_2.IN2 0.0112f
C125 mux_4x1_0.mux_2x1_2.nand2_2.OUT I4 0.202f
C126 mux_4x1_1.mux_2x1_0.nand2_2.IN2 mux_4x1_0.mux_2x1_0.nand2_2.IN2 0.00216f
C127 mux_4x1_1.mux_2x1_2.nand2_1.IN2 a_801_n1395# 0.00372f
C128 mux_2x1_0.nand2_2.IN2 VDD 0.402f
C129 a_3053_n795# S1 2.62e-19
C130 a_238_n1395# I1 0.00347f
C131 mux_4x1_0.mux_2x1_0.nand2_2.IN2 mux_4x1_0.mux_2x1_1.I0 0.0189f
C132 I4 mux_4x1_0.mux_2x1_1.I0 0.0148f
C133 S1 mux_4x1_0.mux_2x1_0.nand2_2.OUT 0.113f
C134 a_2490_n1395# mux_4x1_1.mux_2x1_1.nand2_1.IN2 0.069f
C135 a_1927_n795# S1 2.15e-19
C136 a_3053_707# mux_4x1_0.mux_2x1_1.nand2_2.IN2 0.00372f
C137 a_3053_1307# mux_4x1_0.mux_2x1_1.I0 2.44e-19
C138 S1 mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.342f
C139 mux_4x1_1.mux_2x1_2.nand2_1.IN2 mux_4x1_1.mux_2x1_2.nand2_2.IN2 0.00212f
C140 mux_2x1_0.nand2_2.IN2 mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.0113f
C141 a_1927_1307# mux_4x1_0.mux_2x1_1.I0 2.44e-19
C142 I6 mux_4x1_0.mux_2x1_1.I0 0.01f
C143 mux_4x1_1.mux_2x1_2.nand2_1.IN2 S0 0.368f
C144 mux_2x1_0.I0 VDD 1.44f
C145 a_2490_1307# mux_4x1_0.mux_2x1_1.I0 1.04e-19
C146 mux_4x1_1.mux_2x1_1.I1 a_2490_n1395# 0.00372f
C147 S1 S0 0.00413f
C148 mux_4x1_1.mux_2x1_1.I0 mux_4x1_0.mux_2x1_1.nand2_2.IN2 9.55e-20
C149 a_1364_1307# mux_4x1_0.mux_2x1_1.I0 0.00211f
C150 mux_4x1_1.mux_2x1_1.I0 a_1364_n1395# 0.00211f
C151 mux_4x1_1.mux_2x1_2.nand2_2.OUT a_801_n1395# 0.00949f
C152 mux_4x1_0.mux_2x1_2.nand2_2.OUT mux_4x1_0.mux_2x1_0.nand2_1.IN2 0.0102f
C153 a_3053_n795# mux_4x1_1.mux_2x1_1.I0 0.00375f
C154 a_1927_n795# mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.0964f
C155 mux_4x1_1.mux_2x1_2.nand2_2.IN2 I0 0.0473f
C156 mux_2x1_0.nand2_2.OUT mux_4x1_0.mux_2x1_1.I0 3.46e-19
C157 S1 mux_4x1_1.mux_2x1_1.nand2_2.OUT 0.00227f
C158 mux_4x1_1.mux_2x1_1.I0 a_801_n1395# 0.069f
C159 I0 S0 0.00507f
C160 VDD a_1927_707# 0.00444f
C161 mux_4x1_0.mux_2x1_0.nand2_1.IN2 mux_4x1_0.mux_2x1_1.I0 0.0169f
C162 a_1927_n795# mux_4x1_1.mux_2x1_1.I0 8.2e-19
C163 mux_4x1_1.mux_2x1_0.nand2_1.IN2 S1 4.51e-21
C164 mux_4x1_1.mux_2x1_2.nand2_1.IN2 a_238_n1395# 0.069f
C165 VDD mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.664f
C166 mux_2x1_0.nand2_2.IN2 a_4178_707# 0.00372f
C167 a_1927_1307# mux_4x1_0.mux_2x1_1.I1 0.069f
C168 I6 mux_4x1_0.mux_2x1_1.I1 1.36e-19
C169 a_3615_1307# S2 0.0144f
C170 mux_2x1_0.I0 mux_4x1_1.mux_2x1_1.nand2_1.IN2 0.11f
C171 mux_4x1_1.mux_2x1_2.nand2_2.OUT mux_4x1_1.mux_2x1_2.nand2_2.IN2 0.12f
C172 S0 mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.00112f
C173 mux_4x1_0.mux_2x1_2.nand2_1.IN2 S0 0.368f
C174 mux_4x1_1.mux_2x1_2.nand2_2.OUT S0 0.0532f
C175 a_2490_1307# mux_4x1_0.mux_2x1_1.I1 0.00372f
C176 I7 a_1364_1307# 0.00347f
C177 a_3053_n1395# mux_4x1_1.mux_2x1_1.nand2_2.OUT 0.00949f
C178 mux_4x1_1.mux_2x1_1.I0 mux_4x1_1.mux_2x1_2.nand2_2.IN2 0.0048f
C179 S2 mux_4x1_0.mux_2x1_1.I0 0.00519f
C180 mux_4x1_1.mux_2x1_1.nand2_1.IN2 VDD 0.461f
C181 mux_4x1_1.mux_2x1_1.I0 S0 0.207f
C182 mux_2x1_0.I0 a_4178_707# 0.00293f
C183 a_4178_1307# mux_2x1_0.nand2_2.OUT 0.00949f
C184 a_801_n795# VDD 0.00444f
C185 mux_4x1_0.mux_2x1_0.nand2_2.IN2 VDD 0.405f
C186 I4 VDD 0.258f
C187 mux_4x1_1.mux_2x1_0.nand2_1.IN2 mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.053f
C188 I7 mux_4x1_0.mux_2x1_0.nand2_1.IN2 0.0959f
C189 mux_4x1_1.mux_2x1_0.nand2_1.IN2 mux_4x1_1.mux_2x1_2.nand2_2.OUT 0.0102f
C190 mux_4x1_1.mux_2x1_1.I0 mux_4x1_1.mux_2x1_1.nand2_2.OUT 0.25f
C191 a_801_707# S0 6.89e-19
C192 mux_4x1_0.mux_2x1_0.nand2_1.IN2 mux_4x1_0.mux_2x1_1.I1 0.109f
C193 mux_2x1_0.nand2_2.IN2 mux_2x1_0.nand2_2.OUT 0.12f
C194 mux_4x1_1.mux_2x1_2.nand2_2.IN2 mux_4x1_0.mux_2x1_2.nand2_2.IN2 0.00216f
C195 a_4178_707# VDD 0.00444f
C196 mux_4x1_1.mux_2x1_1.I1 VDD 0.423f
C197 OUT mux_2x1_0.nand2_1.IN2 0.109f
C198 mux_4x1_0.mux_2x1_2.nand2_2.IN2 S0 0.162f
C199 mux_4x1_1.mux_2x1_0.nand2_1.IN2 mux_4x1_1.mux_2x1_1.I0 0.0169f
C200 a_3053_1307# VDD 0.00444f
C201 I2 mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.0036f
C202 mux_4x1_1.mux_2x1_0.nand2_2.IN2 I2 0.0473f
C203 mux_2x1_0.I1 mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.109f
C204 a_1927_1307# VDD 0.00444f
C205 I6 VDD 0.258f
C206 mux_4x1_0.mux_2x1_0.nand2_2.IN2 a_1927_707# 0.00372f
C207 a_2490_1307# VDD 3.14e-19
C208 I2 mux_4x1_0.mux_2x1_1.I0 1.04e-19
C209 I3 mux_4x1_1.mux_2x1_2.nand2_2.OUT 0.0174f
C210 a_1364_1307# VDD 3.14e-19
C211 mux_2x1_0.nand2_1.IN2 mux_2x1_0.I1 0.11f
C212 mux_2x1_0.I1 S0 6.5e-20
C213 mux_2x1_0.nand2_2.IN2 S2 0.136f
C214 mux_2x1_0.I0 mux_2x1_0.nand2_2.OUT 0.234f
C215 S1 mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.16f
C216 mux_4x1_1.mux_2x1_0.nand2_2.IN2 S1 0.00266f
C217 I3 mux_4x1_1.mux_2x1_1.I0 0.0454f
C218 a_3053_1307# mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.00949f
C219 I5 VDD 0.147f
C220 I6 a_1927_707# 0.00293f
C221 mux_2x1_0.nand2_2.OUT VDD 0.635f
C222 mux_4x1_0.mux_2x1_0.nand2_2.OUT mux_4x1_0.mux_2x1_1.nand2_2.IN2 0.0112f
C223 S1 mux_4x1_0.mux_2x1_1.I0 0.0874f
C224 mux_4x1_1.mux_2x1_1.I1 mux_4x1_1.mux_2x1_1.nand2_1.IN2 0.11f
C225 a_1927_n1395# mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.00949f
C226 mux_4x1_0.mux_2x1_0.nand2_1.IN2 VDD 0.46f
C227 mux_4x1_0.mux_2x1_2.nand2_2.OUT I0 3e-19
C228 mux_4x1_1.mux_2x1_0.nand2_2.IN2 I0 0.0036f
C229 mux_4x1_0.mux_2x1_1.nand2_2.IN2 mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.00212f
C230 a_801_1307# mux_4x1_0.mux_2x1_2.nand2_1.IN2 0.00372f
C231 mux_2x1_0.I0 S2 4.25e-19
C232 I4 mux_4x1_0.mux_2x1_0.nand2_2.IN2 0.0036f
C233 a_1927_n1395# mux_4x1_1.mux_2x1_1.I0 2.44e-19
C234 a_2490_n1395# S1 0.0144f
C235 mux_4x1_0.mux_2x1_2.nand2_1.IN2 mux_4x1_0.mux_2x1_2.nand2_2.OUT 0.053f
C236 mux_4x1_1.mux_2x1_0.nand2_2.OUT mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.0112f
C237 mux_4x1_1.mux_2x1_0.nand2_2.IN2 mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.12f
C238 S2 VDD 0.596f
C239 mux_4x1_0.mux_2x1_2.nand2_2.OUT mux_4x1_1.mux_2x1_2.nand2_2.OUT 0.00342f
C240 VDD I1 0.147f
C241 mux_4x1_1.mux_2x1_2.nand2_2.OUT mux_4x1_1.mux_2x1_0.nand2_2.IN2 0.0112f
C242 a_1364_n1395# S0 0.0151f
C243 I6 mux_4x1_0.mux_2x1_0.nand2_2.IN2 0.0473f
C244 mux_4x1_0.mux_2x1_0.nand2_2.OUT mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.0106f
C245 a_3053_707# mux_4x1_0.mux_2x1_1.I0 0.00375f
C246 mux_4x1_1.mux_2x1_1.I0 mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.0646f
C247 mux_4x1_1.mux_2x1_0.nand2_2.IN2 mux_4x1_1.mux_2x1_1.I0 0.0189f
C248 mux_4x1_0.mux_2x1_2.nand2_1.IN2 mux_4x1_0.mux_2x1_1.I0 0.109f
C249 a_801_n1395# S0 9.5e-19
C250 S1 mux_4x1_0.mux_2x1_1.I1 0.0593f
C251 a_238_1307# VDD 3.14e-19
C252 mux_4x1_0.mux_2x1_0.nand2_2.OUT S0 0.00113f
C253 a_1927_n795# S0 2.62e-19
C254 mux_4x1_1.mux_2x1_1.I0 mux_4x1_0.mux_2x1_1.I0 0.285f
C255 mux_2x1_0.nand2_2.IN2 S1 2.44e-19
C256 S2 mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.109f
C257 mux_4x1_0.mux_2x1_2.nand2_2.OUT a_801_707# 0.0964f
C258 a_3053_n795# mux_4x1_1.mux_2x1_1.nand2_2.OUT 0.0964f
C259 mux_4x1_1.mux_2x1_0.nand2_1.IN2 a_1364_n1395# 0.069f
C260 S0 mux_4x1_0.mux_2x1_1.nand2_1.IN2 4.45e-19
C261 a_2490_n1395# mux_4x1_1.mux_2x1_0.nand2_2.OUT 9.43e-19
C262 mux_4x1_0.mux_2x1_2.nand2_2.OUT mux_4x1_0.mux_2x1_2.nand2_2.IN2 0.12f
C263 mux_2x1_0.nand2_2.OUT a_4178_707# 0.0964f
C264 mux_4x1_0.mux_2x1_0.nand2_1.IN2 mux_4x1_0.mux_2x1_0.nand2_2.IN2 0.00212f
C265 a_801_707# mux_4x1_0.mux_2x1_1.I0 1.5e-19
C266 a_2490_n1395# mux_4x1_1.mux_2x1_1.I0 1.04e-19
C267 mux_4x1_1.mux_2x1_2.nand2_2.IN2 S0 0.162f
C268 I2 VDD 0.261f
C269 mux_4x1_0.mux_2x1_2.nand2_2.IN2 mux_4x1_0.mux_2x1_1.I0 0.0048f
C270 mux_2x1_0.I0 S1 0.0118f
C271 I3 a_1364_n1395# 0.00347f
C272 a_1927_1307# mux_4x1_0.mux_2x1_0.nand2_1.IN2 0.00372f
C273 a_3615_1307# mux_2x1_0.I1 0.00372f
C274 mux_4x1_1.mux_2x1_2.nand2_1.IN2 VDD 0.456f
C275 a_4178_707# S2 2.62e-19
C276 S1 VDD 1.58f
C277 a_1364_1307# mux_4x1_0.mux_2x1_0.nand2_1.IN2 0.069f
C278 mux_2x1_0.I1 mux_4x1_0.mux_2x1_1.I0 5.19e-19
C279 mux_4x1_1.mux_2x1_0.nand2_1.IN2 S0 0.378f
C280 mux_2x1_0.I0 a_3053_n1395# 0.069f
C281 a_238_n1395# S0 0.0144f
C282 I0 VDD 0.258f
C283 S1 a_1927_707# 2.15e-19
C284 OUT a_4178_1307# 0.069f
C285 a_3053_n1395# VDD 0.00444f
C286 S1 mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.00228f
C287 mux_4x1_0.mux_2x1_1.nand2_2.IN2 mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.00216f
C288 I3 S0 0.0665f
C289 a_3053_707# VDD 0.00444f
C290 mux_2x1_0.I0 mux_4x1_1.mux_2x1_1.I0 0.0449f
C291 VDD mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.665f
C292 mux_4x1_0.mux_2x1_2.nand2_1.IN2 VDD 0.456f
C293 mux_2x1_0.nand2_2.OUT S2 4.46e-19
C294 mux_4x1_1.mux_2x1_2.nand2_2.OUT VDD 0.664f
C295 a_3053_n795# mux_4x1_1.mux_2x1_1.nand2_2.IN2 0.00372f
C296 S1 mux_4x1_1.mux_2x1_1.nand2_1.IN2 0.342f
C297 mux_4x1_0.mux_2x1_1.nand2_2.IN2 mux_4x1_0.mux_2x1_1.I0 0.0646f
C298 mux_4x1_1.mux_2x1_1.I1 I2 1.36e-19
C299 mux_4x1_1.mux_2x1_1.I0 VDD 1.36f
C300 a_238_1307# I5 0.00347f
C301 mux_4x1_1.mux_2x1_0.nand2_2.IN2 a_1927_n795# 0.00372f
C302 I2 I6 0.00246f
C303 a_3053_707# mux_4x1_0.mux_2x1_1.nand2_2.OUT 0.0964f
C304 mux_4x1_1.mux_2x1_0.nand2_1.IN2 I3 0.0959f
C305 S1 mux_4x1_0.mux_2x1_0.nand2_2.IN2 0.00266f
C306 mux_2x1_0.I0 OUT 1.49e-19
C307 a_801_1307# S0 9.5e-19
C308 mux_4x1_0.mux_2x1_0.nand2_2.OUT mux_4x1_0.mux_2x1_1.I0 0.0241f
C309 mux_4x1_1.mux_2x1_1.I1 S1 0.0593f
C310 a_801_707# VDD 0.00444f
C311 a_3053_n1395# mux_4x1_1.mux_2x1_1.nand2_1.IN2 0.00372f
C312 mux_4x1_0.mux_2x1_2.nand2_2.IN2 VDD 0.404f
C313 OUT VDD 0.234f
C314 a_801_n795# I0 0.00293f
C315 mux_4x1_0.mux_2x1_2.nand2_2.OUT S0 0.0532f
C316 I6 S1 0.00831f
C317 mux_4x1_0.mux_2x1_1.I0 mux_4x1_0.mux_2x1_1.nand2_1.IN2 0.00154f
C318 a_3615_1307# mux_2x1_0.nand2_1.IN2 0.069f
C319 mux_4x1_1.mux_2x1_0.nand2_2.IN2 S0 0.136f
C320 I4 I0 0.00246f
C321 mux_4x1_1.mux_2x1_1.nand2_1.IN2 mux_4x1_1.mux_2x1_0.nand2_2.OUT 0.0106f
C322 mux_2x1_0.I0 mux_2x1_0.I1 2.74e-20
C323 S1 a_2490_1307# 0.0144f
C324 mux_4x1_1.mux_2x1_0.nand2_1.IN2 a_1927_n1395# 0.00372f
C325 a_3053_n1395# VSS 0.0676f
C326 a_2490_n1395# VSS 0.0676f
C327 a_1927_n1395# VSS 0.0676f
C328 a_1364_n1395# VSS 0.0676f
C329 a_801_n1395# VSS 0.0676f
C330 a_238_n1395# VSS 0.0678f
C331 mux_4x1_1.mux_2x1_1.nand2_1.IN2 VSS 0.412f
C332 mux_4x1_1.mux_2x1_1.I1 VSS 0.416f
C333 mux_4x1_1.mux_2x1_0.nand2_1.IN2 VSS 0.412f
C334 I3 VSS 0.257f
C335 mux_4x1_1.mux_2x1_2.nand2_1.IN2 VSS 0.435f
C336 I1 VSS 0.292f
C337 a_3053_n795# VSS 0.0676f
C338 a_1927_n795# VSS 0.0676f
C339 a_801_n795# VSS 0.0676f
C340 mux_4x1_1.mux_2x1_1.nand2_2.OUT VSS 0.598f
C341 mux_4x1_1.mux_2x1_1.I0 VSS 0.771f
C342 mux_4x1_1.mux_2x1_1.nand2_2.IN2 VSS 0.416f
C343 mux_4x1_1.mux_2x1_0.nand2_2.OUT VSS 0.489f
C344 I2 VSS 0.226f
C345 mux_4x1_1.mux_2x1_0.nand2_2.IN2 VSS 0.417f
C346 mux_4x1_1.mux_2x1_2.nand2_2.OUT VSS 0.43f
C347 I0 VSS 0.226f
C348 mux_4x1_1.mux_2x1_2.nand2_2.IN2 VSS 0.436f
C349 a_4178_707# VSS 0.0676f
C350 mux_2x1_0.I0 VSS 1.4f
C351 mux_2x1_0.nand2_2.IN2 VSS 0.422f
C352 a_3053_707# VSS 0.0676f
C353 mux_4x1_0.mux_2x1_1.nand2_2.IN2 VSS 0.417f
C354 a_1927_707# VSS 0.0676f
C355 I6 VSS 0.226f
C356 mux_4x1_0.mux_2x1_0.nand2_2.IN2 VSS 0.417f
C357 a_801_707# VSS 0.0676f
C358 I4 VSS 0.226f
C359 mux_4x1_0.mux_2x1_2.nand2_2.IN2 VSS 0.436f
C360 a_4178_1307# VSS 0.0676f
C361 a_3615_1307# VSS 0.0676f
C362 a_3053_1307# VSS 0.0676f
C363 a_2490_1307# VSS 0.0676f
C364 a_1927_1307# VSS 0.0676f
C365 a_1364_1307# VSS 0.0676f
C366 a_801_1307# VSS 0.0676f
C367 a_238_1307# VSS 0.0678f
C368 OUT VSS 0.14f
C369 mux_4x1_0.mux_2x1_1.I0 VSS 0.714f
C370 mux_2x1_0.nand2_2.OUT VSS 0.653f
C371 mux_2x1_0.nand2_1.IN2 VSS 0.412f
C372 S2 VSS 0.714f
C373 mux_2x1_0.I1 VSS 0.416f
C374 mux_4x1_0.mux_2x1_1.nand2_2.OUT VSS 0.489f
C375 mux_4x1_0.mux_2x1_1.nand2_1.IN2 VSS 0.412f
C376 S1 VSS 1.53f
C377 mux_4x1_0.mux_2x1_1.I1 VSS 0.416f
C378 mux_4x1_0.mux_2x1_0.nand2_2.OUT VSS 0.489f
C379 mux_4x1_0.mux_2x1_0.nand2_1.IN2 VSS 0.412f
C380 I7 VSS 0.257f
C381 mux_4x1_0.mux_2x1_2.nand2_2.OUT VSS 0.43f
C382 mux_4x1_0.mux_2x1_2.nand2_1.IN2 VSS 0.435f
C383 S0 VSS 3.97f
C384 I5 VSS 0.292f
C385 VDD VSS 27.7f
C386 S0.t5 VSS 0.0227f
C387 S0.t9 VSS 0.0284f
C388 S0.n0 VSS 0.0671f
C389 S0.n1 VSS 0.0171f
C390 S0.t7 VSS 0.0227f
C391 S0.t12 VSS 0.0284f
C392 S0.n2 VSS 0.0672f
C393 S0.n3 VSS 0.0353f
C394 S0.n4 VSS 0.00872f
C395 S0.t15 VSS 0.00827f
C396 S0.t10 VSS 0.0329f
C397 S0.n5 VSS 0.0535f
C398 S0.n6 VSS 0.0184f
C399 S0.n7 VSS 0.132f
C400 S0.n8 VSS 0.325f
C401 S0.n9 VSS 0.00731f
C402 S0.n10 VSS 0.00355f
C403 S0.t0 VSS 0.0329f
C404 S0.t6 VSS 0.00827f
C405 S0.n11 VSS 0.0535f
C406 S0.n12 VSS 0.00355f
C407 S0.t14 VSS 0.0227f
C408 S0.t13 VSS 0.0284f
C409 S0.n13 VSS 0.0672f
C410 S0.n14 VSS 0.0352f
C411 S0.n15 VSS 0.00871f
C412 S0.t4 VSS 0.0329f
C413 S0.t11 VSS 0.00827f
C414 S0.n16 VSS 0.0535f
C415 S0.n17 VSS 0.0184f
C416 S0.n18 VSS 0.132f
C417 S0.n19 VSS 0.325f
C418 S0.n20 VSS 0.00965f
C419 S0.t3 VSS 0.0227f
C420 S0.t1 VSS 0.0284f
C421 S0.n21 VSS 0.0671f
C422 S0.n22 VSS 0.0274f
C423 S0.n23 VSS 3.88e-19
C424 S0.n24 VSS 0.19f
C425 S0.n25 VSS 0.134f
C426 S0.n26 VSS 0.133f
C427 S0.n27 VSS 0.0071f
C428 S0.n28 VSS 8.22e-19
C429 S0.n29 VSS 0.0176f
C430 S0.n30 VSS 0.185f
C431 S0.n31 VSS 0.185f
C432 S0.n32 VSS 0.0174f
C433 S0.t8 VSS 0.00827f
C434 S0.t2 VSS 0.0329f
C435 S0.n33 VSS 0.0535f
C436 S0.n34 VSS 0.00103f
C437 S0.n35 VSS 0.133f
C438 S0.n36 VSS 0.134f
C439 S0.n37 VSS 0.19f
C440 S0.n38 VSS 3.88e-19
C441 S0.n39 VSS 0.00964f
C442 VDD.t24 VSS 0.0685f
C443 VDD.n0 VSS 0.0327f
C444 VDD.t35 VSS 0.00199f
C445 VDD.n1 VSS 0.0166f
C446 VDD.t58 VSS 0.00199f
C447 VDD.n2 VSS 0.0166f
C448 VDD.t64 VSS 0.0295f
C449 VDD.t34 VSS 0.0359f
C450 VDD.n4 VSS 0.0283f
C451 VDD.t56 VSS 0.0296f
C452 VDD.n5 VSS 0.0294f
C453 VDD.t65 VSS 0.00264f
C454 VDD.t57 VSS 0.00264f
C455 VDD.n6 VSS 0.0217f
C456 VDD.n7 VSS 0.0124f
C457 VDD.n8 VSS 0.00263f
C458 VDD.n9 VSS 0.00263f
C459 VDD.t69 VSS 0.0685f
C460 VDD.n10 VSS 0.0327f
C461 VDD.t37 VSS 0.00199f
C462 VDD.n11 VSS 0.0166f
C463 VDD.t43 VSS 0.0296f
C464 VDD.t36 VSS 0.0359f
C465 VDD.n12 VSS 0.0283f
C466 VDD.t95 VSS 0.0295f
C467 VDD.t96 VSS 0.00274f
C468 VDD.n14 VSS 0.0331f
C469 VDD.n15 VSS 0.0294f
C470 VDD.t44 VSS 0.00274f
C471 VDD.n16 VSS 0.033f
C472 VDD.n17 VSS 0.00812f
C473 VDD.t40 VSS 0.00199f
C474 VDD.n18 VSS 0.00814f
C475 VDD.n19 VSS 0.00263f
C476 VDD.t10 VSS 0.0347f
C477 VDD.n20 VSS 0.00263f
C478 VDD.t84 VSS 0.00216f
C479 VDD.n21 VSS 0.0183f
C480 VDD.t80 VSS 0.0347f
C481 VDD.n22 VSS 0.00263f
C482 VDD.n23 VSS 0.00289f
C483 VDD.t87 VSS 0.0343f
C484 VDD.t99 VSS 0.0317f
C485 VDD.n24 VSS 0.0163f
C486 VDD.n25 VSS 0.00814f
C487 VDD.t100 VSS 0.00216f
C488 VDD.t32 VSS 0.00199f
C489 VDD.n26 VSS 0.0166f
C490 VDD.n27 VSS 0.00263f
C491 VDD.n28 VSS 0.00263f
C492 VDD.t30 VSS 0.00269f
C493 VDD.t29 VSS 0.0296f
C494 VDD.t92 VSS 0.0343f
C495 VDD.n29 VSS 0.00289f
C496 VDD.t102 VSS 0.00199f
C497 VDD.t9 VSS 0.00216f
C498 VDD.n30 VSS 0.00289f
C499 VDD.n31 VSS 0.00814f
C500 VDD.n32 VSS 0.00263f
C501 VDD.t5 VSS 0.0343f
C502 VDD.n33 VSS 0.0163f
C503 VDD.t8 VSS 0.0317f
C504 VDD.t108 VSS 0.0347f
C505 VDD.n34 VSS 0.0163f
C506 VDD.t4 VSS 0.00263f
C507 VDD.n35 VSS 0.00263f
C508 VDD.t3 VSS 0.0316f
C509 VDD.t19 VSS 0.0346f
C510 VDD.n36 VSS 0.0163f
C511 VDD.t75 VSS 0.00216f
C512 VDD.n37 VSS 0.0183f
C513 VDD.n38 VSS 0.00263f
C514 VDD.t74 VSS 0.0317f
C515 VDD.t0 VSS 0.0347f
C516 VDD.n39 VSS 0.0163f
C517 VDD.t104 VSS 0.00263f
C518 VDD.n40 VSS 0.00263f
C519 VDD.t103 VSS 0.0317f
C520 VDD.t50 VSS 0.0347f
C521 VDD.n41 VSS 0.0163f
C522 VDD.n42 VSS 0.00263f
C523 VDD.t41 VSS 0.0317f
C524 VDD.t16 VSS 0.0347f
C525 VDD.n43 VSS 0.0163f
C526 VDD.t49 VSS 0.00263f
C527 VDD.n44 VSS 0.00263f
C528 VDD.t48 VSS 0.0317f
C529 VDD.t53 VSS 0.0347f
C530 VDD.n45 VSS 0.0163f
C531 VDD.t73 VSS 0.00216f
C532 VDD.n46 VSS 0.0183f
C533 VDD.n47 VSS 0.00263f
C534 VDD.t72 VSS 0.0317f
C535 VDD.t66 VSS 0.0347f
C536 VDD.t90 VSS 0.0316f
C537 VDD.n48 VSS 0.0163f
C538 VDD.t91 VSS 0.00282f
C539 VDD.n49 VSS 0.0202f
C540 VDD.n50 VSS 0.013f
C541 VDD.n51 VSS 0.00886f
C542 VDD.n52 VSS 0.00814f
C543 VDD.n53 VSS 0.013f
C544 VDD.n54 VSS 0.012f
C545 VDD.n55 VSS 0.00542f
C546 VDD.n56 VSS 0.013f
C547 VDD.t42 VSS 0.00216f
C548 VDD.n57 VSS 0.0183f
C549 VDD.n58 VSS 0.00886f
C550 VDD.n59 VSS 0.00814f
C551 VDD.n60 VSS 0.013f
C552 VDD.n61 VSS 0.0121f
C553 VDD.n62 VSS 0.00814f
C554 VDD.n63 VSS 0.013f
C555 VDD.n64 VSS 0.00886f
C556 VDD.n65 VSS 0.00814f
C557 VDD.n66 VSS 0.013f
C558 VDD.n67 VSS 0.0121f
C559 VDD.n68 VSS 0.00814f
C560 VDD.n69 VSS 0.013f
C561 VDD.n70 VSS 0.00886f
C562 VDD.n71 VSS 0.0183f
C563 VDD.n72 VSS 0.0166f
C564 VDD.n73 VSS 0.00949f
C565 VDD.n74 VSS 0.00814f
C566 VDD.n75 VSS 0.0163f
C567 VDD.t101 VSS 0.018f
C568 VDD.n76 VSS 0.0288f
C569 VDD.n77 VSS 0.0203f
C570 VDD.n78 VSS 0.0252f
C571 VDD.n79 VSS 0.0259f
C572 VDD.n80 VSS 0.0163f
C573 VDD.t78 VSS 0.0295f
C574 VDD.t105 VSS 0.0685f
C575 VDD.n82 VSS 0.0327f
C576 VDD.t31 VSS 0.0359f
C577 VDD.n83 VSS 0.0283f
C578 VDD.t97 VSS 0.0296f
C579 VDD.n84 VSS 0.0294f
C580 VDD.t79 VSS 0.00264f
C581 VDD.t98 VSS 0.00264f
C582 VDD.n85 VSS 0.0217f
C583 VDD.n86 VSS 0.0158f
C584 VDD.n87 VSS 0.00263f
C585 VDD.n88 VSS 0.00263f
C586 VDD.n89 VSS 0.0203f
C587 VDD.n90 VSS 0.026f
C588 VDD.n91 VSS 0.0126f
C589 VDD.n92 VSS 0.0217f
C590 VDD.n93 VSS 0.00773f
C591 VDD.n94 VSS 0.0114f
C592 VDD.t33 VSS 0.00199f
C593 VDD.n95 VSS 0.0166f
C594 VDD.n96 VSS 0.0183f
C595 VDD.n97 VSS 0.00886f
C596 VDD.n98 VSS 0.013f
C597 VDD.t77 VSS 0.00263f
C598 VDD.n99 VSS 0.00263f
C599 VDD.n100 VSS 0.013f
C600 VDD.n101 VSS 0.0121f
C601 VDD.n102 VSS 0.00814f
C602 VDD.n103 VSS 0.0163f
C603 VDD.t76 VSS 0.0317f
C604 VDD.t13 VSS 0.0347f
C605 VDD.t83 VSS 0.0317f
C606 VDD.n104 VSS 0.0163f
C607 VDD.n105 VSS 0.00814f
C608 VDD.n106 VSS 0.00886f
C609 VDD.n107 VSS 0.013f
C610 VDD.t23 VSS 0.00263f
C611 VDD.n108 VSS 0.00263f
C612 VDD.n109 VSS 0.013f
C613 VDD.n110 VSS 0.012f
C614 VDD.n111 VSS 0.00542f
C615 VDD.n112 VSS 0.0163f
C616 VDD.t22 VSS 0.0317f
C617 VDD.t59 VSS 0.0347f
C618 VDD.n113 VSS 0.0163f
C619 VDD.t38 VSS 0.0317f
C620 VDD.t45 VSS 0.0347f
C621 VDD.t27 VSS 0.0316f
C622 VDD.n114 VSS 0.0163f
C623 VDD.t28 VSS 0.00282f
C624 VDD.n115 VSS 0.0202f
C625 VDD.n116 VSS 0.013f
C626 VDD.n117 VSS 0.00886f
C627 VDD.t39 VSS 0.00216f
C628 VDD.n118 VSS 0.0183f
C629 VDD.n119 VSS 0.0166f
C630 VDD.n120 VSS 0.0111f
C631 VDD.n121 VSS 0.0163f
C632 VDD.n122 VSS 0.0208f
C633 VDD.n123 VSS 0.0292f
C634 VDD.n124 VSS 0.0124f
C635 VDD.n125 VSS 0.0217f
C636 VDD.n126 VSS 0.00812f
C637 VDD.n127 VSS 0.0111f
C638 VDD.n128 VSS 0.0163f
.ends

