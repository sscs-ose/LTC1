magic
tech gf180mcuC
magscale 1 10
timestamp 1694400330
<< nwell >>
rect 536 700 1360 813
<< psubdiff >>
rect 558 80 1329 95
rect 558 34 577 80
rect 1306 34 1329 80
rect 558 19 1329 34
<< nsubdiff >>
rect 564 774 1327 789
rect 564 728 593 774
rect 1305 728 1327 774
rect 564 715 1327 728
<< psubdiffcont >>
rect 577 34 1306 80
<< nsubdiffcont >>
rect 593 728 1305 774
<< polysilicon >>
rect 1412 664 1501 678
rect 1412 658 1425 664
rect 1126 606 1425 658
rect 1412 604 1425 606
rect 1488 604 1501 664
rect 1412 591 1501 604
rect 714 473 770 484
rect 703 460 792 473
rect 703 400 716 460
rect 779 400 792 460
rect 703 386 792 400
rect 413 301 502 315
rect 413 241 426 301
rect 489 241 502 301
rect 413 228 502 241
rect 451 179 496 228
rect 1414 206 1503 220
rect 1414 188 1427 206
rect 451 132 708 179
rect 1188 146 1427 188
rect 1490 146 1503 206
rect 1188 142 1503 146
rect 1414 133 1503 142
<< polycontact >>
rect 1425 604 1488 664
rect 716 400 779 460
rect 426 241 489 301
rect 1427 146 1490 206
<< metal1 >>
rect 404 774 1360 813
rect 404 728 593 774
rect 1305 728 1360 774
rect 404 700 1360 728
rect 440 614 527 632
rect 440 549 453 614
rect 518 576 527 614
rect 518 549 692 576
rect 440 547 692 549
rect 446 525 692 547
rect 790 525 861 700
rect 1035 525 1106 700
rect 1412 664 1501 678
rect 1412 604 1425 664
rect 1488 604 1501 664
rect 1412 591 1501 604
rect 1204 525 1335 574
rect 446 505 631 525
rect -23 398 74 415
rect -23 340 2 398
rect 60 340 74 398
rect 357 371 459 418
rect -23 337 74 340
rect 412 315 459 371
rect 412 301 502 315
rect 412 287 426 301
rect 413 241 426 287
rect 489 241 502 301
rect 413 228 502 241
rect 560 221 631 505
rect 703 460 792 473
rect 703 400 716 460
rect 779 400 792 460
rect 703 386 792 400
rect 1266 456 1335 525
rect 1266 397 1275 456
rect 1327 397 1335 456
rect 729 113 801 268
rect 1097 113 1167 268
rect 1266 221 1335 397
rect 1414 206 1503 220
rect 1414 146 1427 206
rect 1490 146 1503 206
rect 1414 133 1503 146
rect 404 80 1360 113
rect 404 34 577 80
rect 1306 34 1360 80
rect 404 0 1360 34
<< via1 >>
rect 453 549 518 614
rect 1425 604 1488 664
rect 2 340 60 398
rect 716 400 779 460
rect 1275 397 1327 456
rect 1427 146 1490 206
<< metal2 >>
rect 1412 672 1501 678
rect 453 664 1501 672
rect 453 632 1425 664
rect 440 614 1425 632
rect 440 549 453 614
rect 518 607 1425 614
rect 518 549 530 607
rect 1412 604 1425 607
rect 1488 604 1501 664
rect 1412 591 1501 604
rect 440 547 530 549
rect 703 460 792 473
rect -23 398 74 415
rect -23 340 2 398
rect 60 340 74 398
rect 703 400 716 460
rect 779 456 1339 460
rect 779 400 1275 456
rect 703 397 1275 400
rect 1327 397 1339 456
rect 703 393 1339 397
rect 703 386 792 393
rect -23 337 74 340
rect 2 202 60 337
rect 1414 206 1503 220
rect 1414 202 1427 206
rect 2 146 1427 202
rect 1490 146 1503 206
rect 2 144 1503 146
rect 1372 138 1503 144
rect 1414 133 1503 138
use Inverter  Inverter_0
timestamp 1693893072
transform 1 0 118 0 1 214
box -118 -214 286 599
use nmos_3p3_DDNVWA  nmos_3p3_DDNVWA_0
timestamp 1692705520
transform 1 0 680 0 1 245
box -144 -97 144 97
use nmos_3p3_DDNVWA  nmos_3p3_DDNVWA_1
timestamp 1692705520
transform 1 0 1216 0 1 245
box -144 -97 144 97
use pmos_3p3_M8LTNG  pmos_3p3_M8LTNG_0
timestamp 1692705520
transform 1 0 742 0 1 550
box -206 -159 206 159
use pmos_3p3_M8LTNG  pmos_3p3_M8LTNG_1
timestamp 1692705520
transform 1 0 1154 0 1 550
box -206 -159 206 159
<< labels >>
flabel nsubdiffcont 932 747 932 747 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel psubdiffcont 940 64 940 64 0 FreeSans 640 0 0 0 VSS
port 1 nsew
flabel via1 1447 643 1447 643 0 FreeSans 640 0 0 0 OUT
port 2 nsew
flabel via1 1299 417 1299 417 0 FreeSans 640 0 0 0 OUT_B
port 3 nsew
flabel via1 26 362 26 362 0 FreeSans 640 0 0 0 VIN
port 4 nsew
<< end >>
