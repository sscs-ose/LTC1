magic
tech gf180mcuC
magscale 1 10
timestamp 1694088395
<< nwell >>
rect -624 -1121 624 1121
<< nsubdiff >>
rect -600 1025 600 1097
rect -600 981 -528 1025
rect -600 -981 -587 981
rect -541 -981 -528 981
rect 528 981 600 1025
rect -600 -1025 -528 -981
rect 528 -981 541 981
rect 587 -981 600 981
rect 528 -1025 600 -981
rect -600 -1097 600 -1025
<< nsubdiffcont >>
rect -587 -981 -541 981
rect 541 -981 587 981
<< polysilicon >>
rect -440 924 -280 937
rect -440 878 -427 924
rect -293 878 -280 924
rect -440 834 -280 878
rect -440 -878 -280 -834
rect -440 -924 -427 -878
rect -293 -924 -280 -878
rect -440 -937 -280 -924
rect -200 924 -40 937
rect -200 878 -187 924
rect -53 878 -40 924
rect -200 834 -40 878
rect -200 -878 -40 -834
rect -200 -924 -187 -878
rect -53 -924 -40 -878
rect -200 -937 -40 -924
rect 40 924 200 937
rect 40 878 53 924
rect 187 878 200 924
rect 40 834 200 878
rect 40 -878 200 -834
rect 40 -924 53 -878
rect 187 -924 200 -878
rect 40 -937 200 -924
rect 280 924 440 937
rect 280 878 293 924
rect 427 878 440 924
rect 280 834 440 878
rect 280 -878 440 -834
rect 280 -924 293 -878
rect 427 -924 440 -878
rect 280 -937 440 -924
<< polycontact >>
rect -427 878 -293 924
rect -427 -924 -293 -878
rect -187 878 -53 924
rect -187 -924 -53 -878
rect 53 878 187 924
rect 53 -924 187 -878
rect 293 878 427 924
rect 293 -924 427 -878
<< ppolyres >>
rect -440 -834 -280 834
rect -200 -834 -40 834
rect 40 -834 200 834
rect 280 -834 440 834
<< metal1 >>
rect -587 1038 587 1084
rect -587 981 -541 1038
rect 541 981 587 1038
rect -438 878 -427 924
rect -293 878 -282 924
rect -198 878 -187 924
rect -53 878 -42 924
rect 42 878 53 924
rect 187 878 198 924
rect 282 878 293 924
rect 427 878 438 924
rect -438 -924 -427 -878
rect -293 -924 -282 -878
rect -198 -924 -187 -878
rect -53 -924 -42 -878
rect 42 -924 53 -878
rect 187 -924 198 -878
rect 282 -924 293 -878
rect 427 -924 438 -878
rect -587 -1038 -541 -981
rect 541 -1038 587 -981
rect -587 -1084 587 -1038
<< properties >>
string FIXED_BBOX -564 -1061 564 1061
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 8.343 m 1 nx 4 wmin 0.80 lmin 1.00 rho 315 val 3.6k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 1
<< end >>
