magic
tech gf180mcuD
magscale 1 5
timestamp 1713185578
<< checkpaint >>
rect -5927 -4180 5927 4180
<< mimcap >>
rect -4867 2972 -1867 3090
rect -4867 208 -4749 2972
rect -1985 208 -1867 2972
rect -4867 90 -1867 208
rect -1560 2972 1440 3090
rect -1560 208 -1442 2972
rect 1322 208 1440 2972
rect -1560 90 1440 208
rect 1747 2972 4747 3090
rect 1747 208 1865 2972
rect 4629 208 4747 2972
rect 1747 90 4747 208
rect -4867 -208 -1867 -90
rect -4867 -2972 -4749 -208
rect -1985 -2972 -1867 -208
rect -4867 -3090 -1867 -2972
rect -1560 -208 1440 -90
rect -1560 -2972 -1442 -208
rect 1322 -2972 1440 -208
rect -1560 -3090 1440 -2972
rect 1747 -208 4747 -90
rect 1747 -2972 1865 -208
rect 4629 -2972 4747 -208
rect 1747 -3090 4747 -2972
<< mimcapcontact >>
rect -4749 208 -1985 2972
rect -1442 208 1322 2972
rect 1865 208 4629 2972
rect -4749 -2972 -1985 -208
rect -1442 -2972 1322 -208
rect 1865 -2972 4629 -208
<< metal4 >>
rect -4927 3112 -1687 3150
rect -4927 3090 -1754 3112
rect -4927 90 -4867 3090
rect -1867 90 -1754 3090
rect -4927 68 -1754 90
rect -1726 68 -1687 3112
rect -4927 30 -1687 68
rect -1620 3112 1620 3150
rect -1620 3090 1553 3112
rect -1620 90 -1560 3090
rect 1440 90 1553 3090
rect -1620 68 1553 90
rect 1581 68 1620 3112
rect -1620 30 1620 68
rect 1687 3112 4927 3150
rect 1687 3090 4860 3112
rect 1687 90 1747 3090
rect 4747 90 4860 3090
rect 1687 68 4860 90
rect 4888 68 4927 3112
rect 1687 30 4927 68
rect -4927 -68 -1687 -30
rect -4927 -90 -1754 -68
rect -4927 -3090 -4867 -90
rect -1867 -3090 -1754 -90
rect -4927 -3112 -1754 -3090
rect -1726 -3112 -1687 -68
rect -4927 -3150 -1687 -3112
rect -1620 -68 1620 -30
rect -1620 -90 1553 -68
rect -1620 -3090 -1560 -90
rect 1440 -3090 1553 -90
rect -1620 -3112 1553 -3090
rect 1581 -3112 1620 -68
rect -1620 -3150 1620 -3112
rect 1687 -68 4927 -30
rect 1687 -90 4860 -68
rect 1687 -3090 1747 -90
rect 4747 -3090 4860 -90
rect 1687 -3112 4860 -3090
rect 4888 -3112 4927 -68
rect 1687 -3150 4927 -3112
<< via4 >>
rect -1754 68 -1726 3112
rect 1553 68 1581 3112
rect 4860 68 4888 3112
rect -1754 -3112 -1726 -68
rect 1553 -3112 1581 -68
rect 4860 -3112 4888 -68
<< metal5 >>
rect -3420 3050 -3314 3180
rect -1793 3112 -1687 3180
rect -4827 2972 -1907 3050
rect -4827 208 -4749 2972
rect -1985 208 -1907 2972
rect -4827 130 -1907 208
rect -3420 -130 -3314 130
rect -1793 68 -1754 3112
rect -1726 68 -1687 3112
rect -113 3050 -7 3180
rect 1514 3112 1620 3180
rect -1520 2972 1400 3050
rect -1520 208 -1442 2972
rect 1322 208 1400 2972
rect -1520 130 1400 208
rect -1793 -68 -1687 68
rect -4827 -208 -1907 -130
rect -4827 -2972 -4749 -208
rect -1985 -2972 -1907 -208
rect -4827 -3050 -1907 -2972
rect -3420 -3180 -3314 -3050
rect -1793 -3112 -1754 -68
rect -1726 -3112 -1687 -68
rect -113 -130 -7 130
rect 1514 68 1553 3112
rect 1581 68 1620 3112
rect 3194 3050 3300 3180
rect 4821 3112 4927 3180
rect 1787 2972 4707 3050
rect 1787 208 1865 2972
rect 4629 208 4707 2972
rect 1787 130 4707 208
rect 1514 -68 1620 68
rect -1520 -208 1400 -130
rect -1520 -2972 -1442 -208
rect 1322 -2972 1400 -208
rect -1520 -3050 1400 -2972
rect -1793 -3180 -1687 -3112
rect -113 -3180 -7 -3050
rect 1514 -3112 1553 -68
rect 1581 -3112 1620 -68
rect 3194 -130 3300 130
rect 4821 68 4860 3112
rect 4888 68 4927 3112
rect 4821 -68 4927 68
rect 1787 -208 4707 -130
rect 1787 -2972 1865 -208
rect 4629 -2972 4707 -208
rect 1787 -3050 4707 -2972
rect 1514 -3180 1620 -3112
rect 3194 -3180 3300 -3050
rect 4821 -3112 4860 -68
rect 4888 -3112 4927 -68
rect 4821 -3180 4927 -3112
<< properties >>
string FIXED_BBOX 1687 30 4807 3150
<< end >>
