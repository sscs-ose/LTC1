* NGSPICE file created from RES_74k_flat.ext - technology: gf180mcuC

.subckt Res_74k_pex P VDD M
X0 P.t63 P.t64 VDD.t12 ppolyf_u r_width=1.1u r_length=2.6u
X1 P.t53 P.t54 VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X2 P.t52 a_4414_3230.t0 VDD.t12 ppolyf_u r_width=1.1u r_length=2.6u
X3 a_7114_2196.t0 a_7414_1574.t0 VDD.t1 ppolyf_u r_width=1.1u r_length=2.6u
X4 a_7714_3852.t0 a_7414_3230.t0 VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X5 P.t16 P.t17 VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X6 P.t77 P.t78 VDD.t1 ppolyf_u r_width=1.1u r_length=2.6u
X7 P.t28 P.t29 VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X8 a_5914_540.t0 a_6214_n82.t1 VDD.t14 ppolyf_u r_width=1.1u r_length=2.6u
X9 a_7414_3024.t1 a_7714_2402.t1 VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X10 a_4414_3024.t0 a_4414_2196.t0 VDD.t12 ppolyf_u r_width=1.1u r_length=2.6u
X11 a_5314_540.t0 a_5014_n82.t1 VDD.t15 ppolyf_u r_width=1.1u r_length=2.6u
X12 P.t85 P.t86 VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X13 a_4414_540.t0 a_4414_n82.t0 VDD.t12 ppolyf_u r_width=1.1u r_length=2.6u
X14 a_6514_2196.t0 a_6814_1574.t1 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X15 P.t22 P.t23 VDD.t15 ppolyf_u r_width=1.1u r_length=2.6u
X16 P.t55 P.t56 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X17 P.t69 P.t70 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X18 a_5314_3852.t0 a_5014_3230.t1 VDD.t15 ppolyf_u r_width=1.1u r_length=2.6u
X19 a_8314_3852.t0 a_8614_3024.t0 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X20 a_5014_1368.t1 a_4714_746.t1 VDD.t2 ppolyf_u r_width=1.1u r_length=2.6u
X21 a_8314_2196.t1 a_8014_1574.t1 VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X22 a_4714_2196.t1 a_5014_1574.t1 VDD.t2 ppolyf_u r_width=1.1u r_length=2.6u
X23 P.t75 P.t76 VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X24 a_8314_540.t1 a_8014_n82.t1 VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X25 a_8614_3024.t1 a_8314_2402.t1 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X26 P.t81 P.t82 VDD.t2 ppolyf_u r_width=1.1u r_length=2.6u
X27 a_5014_3024.t1 a_5314_2402.t1 VDD.t15 ppolyf_u r_width=1.1u r_length=2.6u
X28 a_7114_540.t0 a_7414_n82.t1 VDD.t1 ppolyf_u r_width=1.1u r_length=2.6u
X29 a_4414_1368.t1 a_4414_540.t1 VDD.t12 ppolyf_u r_width=1.1u r_length=2.6u
X30 P.t59 P.t60 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X31 a_6514_540.t1 a_6214_n82.t0 VDD.t16 ppolyf_u r_width=1.1u r_length=2.6u
X32 a_5014_1368.t0 a_5314_746.t1 VDD.t15 ppolyf_u r_width=1.1u r_length=2.6u
X33 a_4714_3852.t1 a_4414_3230.t1 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X34 a_7714_2196.t1 a_7414_1574.t1 VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X35 a_4414_2196.t1 a_4414_1574.t1 VDD.t12 ppolyf_u r_width=1.1u r_length=2.6u
X36 P.t71 P.t72 VDD.t14 ppolyf_u r_width=1.1u r_length=2.6u
X37 P.t87 P.t88 VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X38 P.t73 P.t74 VDD.t12 ppolyf_u r_width=1.1u r_length=2.6u
X39 a_5314_540.t1 a_5614_n82.t1 VDD.t13 ppolyf_u r_width=1.1u r_length=2.6u
X40 a_4414_3024.t1 a_4714_2402.t1 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X41 a_4414_1368.t0 a_4714_746.t0 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X42 a_5914_3852.t0 a_6214_3230.t1 VDD.t14 ppolyf_u r_width=1.1u r_length=2.6u
X43 a_6214_1368.t0 a_5914_746.t1 VDD.t14 ppolyf_u r_width=1.1u r_length=2.6u
X44 a_6214_3024.t1 a_5914_2402.t0 VDD.t14 ppolyf_u r_width=1.1u r_length=2.6u
X45 a_4714_540.t1 a_4414_n82.t1 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X46 a_5614_1368.t1 a_5314_746.t0 VDD.t13 ppolyf_u r_width=1.1u r_length=2.6u
X47 a_6814_1368.t0 a_7114_746.t1 VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X48 a_8314_540.t0 M.t0 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X49 P.t38 P.t39 VDD.t13 ppolyf_u r_width=1.1u r_length=2.6u
X50 P.t30 P.t31 VDD.t11 ppolyf_u r_width=1.1u r_length=2.6u
X51 a_6214_1368.t1 a_6514_746.t1 VDD.t16 ppolyf_u r_width=1.1u r_length=2.6u
X52 a_5314_3852.t1 a_5614_3230.t1 VDD.t13 ppolyf_u r_width=1.1u r_length=2.6u
X53 a_8014_1368.t1 a_7714_746.t1 VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X54 P.t10 P.t11 VDD.t11 ppolyf_u r_width=1.1u r_length=2.6u
X55 a_8314_2196.t0 a_8614_1368.t1 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X56 a_5314_2196.t1 a_5014_1574.t0 VDD.t15 ppolyf_u r_width=1.1u r_length=2.6u
X57 P.t12 P.t13 VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X58 P.t14 P.t15 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X59 P.t46 P.t47 VDD.t15 ppolyf_u r_width=1.1u r_length=2.6u
X60 a_7714_540.t0 a_7414_n82.t0 VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X61 P.t36 P.t37 VDD.t11 ppolyf_u r_width=1.1u r_length=2.6u
X62 a_5614_3024.t0 a_5314_2402.t0 VDD.t13 ppolyf_u r_width=1.1u r_length=2.6u
X63 a_7114_3852.t0 a_6814_3230.t1 VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X64 a_5614_1368.t0 a_5914_746.t0 VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X65 a_7414_1368.t1 a_7114_746.t0 VDD.t1 ppolyf_u r_width=1.1u r_length=2.6u
X66 a_6814_3024.t1 a_7114_2402.t1 VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X67 a_6514_540.t0 a_6814_n82.t0 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X68 a_6814_1368.t1 a_6514_746.t0 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X69 a_5914_540.t1 a_5614_n82.t0 VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X70 a_8014_1368.t0 a_8314_746.t1 VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X71 a_4714_2196.t0 a_4414_1574.t0 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X72 P.t26 P.t27 VDD.t16 ppolyf_u r_width=1.1u r_length=2.6u
X73 P.t0 P.t1 VDD.t5 ppolyf_u r_width=1.1u r_length=2.6u
X74 a_7414_1368.t0 a_7714_746.t0 VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X75 a_5914_2196.t0 a_6214_1574.t0 VDD.t14 ppolyf_u r_width=1.1u r_length=2.6u
X76 a_6514_3852.t1 a_6214_3230.t0 VDD.t16 ppolyf_u r_width=1.1u r_length=2.6u
X77 P.t44 P.t45 VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X78 P.t42 P.t43 VDD.t14 ppolyf_u r_width=1.1u r_length=2.6u
X79 a_6214_3024.t0 a_6514_2402.t1 VDD.t16 ppolyf_u r_width=1.1u r_length=2.6u
X80 a_7714_3852.t1 a_8014_3230.t0 VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X81 P.t32 P.t33 VDD.t11 ppolyf_u r_width=1.1u r_length=2.6u
X82 a_8014_3024.t1 a_7714_2402.t0 VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X83 a_8614_1368.t0 a_8314_746.t0 VDD.t4 ppolyf_u r_width=1.1u r_length=2.6u
X84 P.t2 P.t3 VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X85 P.t48 P.t49 VDD.t11 ppolyf_u r_width=1.1u r_length=2.6u
X86 a_5314_2196.t0 a_5614_1574.t0 VDD.t13 ppolyf_u r_width=1.1u r_length=2.6u
X87 a_5914_3852.t1 a_5614_3230.t0 VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X88 P.t57 P.t58 VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X89 P.t50 P.t51 VDD.t1 ppolyf_u r_width=1.1u r_length=2.6u
X90 P.t61 P.t62 VDD.t11 ppolyf_u r_width=1.1u r_length=2.6u
X91 P.t40 P.t41 VDD.t13 ppolyf_u r_width=1.1u r_length=2.6u
X92 a_5614_3024.t1 a_5914_2402.t1 VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X93 P.t4 P.t5 VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X94 a_7114_3852.t1 a_7414_3230.t1 VDD.t1 ppolyf_u r_width=1.1u r_length=2.6u
X95 P.t67 P.t68 VDD.t11 ppolyf_u r_width=1.1u r_length=2.6u
X96 a_7114_2196.t1 a_6814_1574.t0 VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X97 P.t65 P.t66 VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
X98 a_7414_3024.t0 a_7114_2402.t0 VDD.t1 ppolyf_u r_width=1.1u r_length=2.6u
X99 P.t20 P.t21 VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X100 P.t83 P.t84 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X101 a_4714_540.t0 a_5014_n82.t0 VDD.t2 ppolyf_u r_width=1.1u r_length=2.6u
X102 a_6514_3852.t0 a_6814_3230.t0 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X103 a_6514_2196.t1 a_6214_1574.t1 VDD.t16 ppolyf_u r_width=1.1u r_length=2.6u
X104 P.t34 P.t35 VDD.t2 ppolyf_u r_width=1.1u r_length=2.6u
X105 P.t18 P.t19 VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X106 P.t24 P.t25 VDD.t16 ppolyf_u r_width=1.1u r_length=2.6u
X107 P.t6 P.t7 VDD.t7 ppolyf_u r_width=1.1u r_length=2.6u
X108 a_6814_3024.t0 a_6514_2402.t0 VDD.t3 ppolyf_u r_width=1.1u r_length=2.6u
X109 a_8314_3852.t1 a_8014_3230.t1 VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X110 a_4714_3852.t0 a_5014_3230.t0 VDD.t2 ppolyf_u r_width=1.1u r_length=2.6u
X111 a_7714_2196.t0 a_8014_1574.t0 VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X112 P.t8 P.t9 VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X113 a_8014_3024.t0 a_8314_2402.t0 VDD.t9 ppolyf_u r_width=1.1u r_length=2.6u
X114 a_5014_3024.t0 a_4714_2402.t0 VDD.t2 ppolyf_u r_width=1.1u r_length=2.6u
X115 a_7714_540.t1 a_8014_n82.t0 VDD.t8 ppolyf_u r_width=1.1u r_length=2.6u
X116 a_5914_2196.t1 a_5614_1574.t1 VDD.t6 ppolyf_u r_width=1.1u r_length=2.6u
X117 P.t79 P.t80 VDD.t0 ppolyf_u r_width=1.1u r_length=2.6u
X118 a_7114_540.t1 a_6814_n82.t1 VDD.t10 ppolyf_u r_width=1.1u r_length=2.6u
R0 P.n92 P.t4 6.1905
R1 P.n28 P.t31 6.1905
R2 P.n44 P.t58 6.1905
R3 P.n43 P.t64 6.1905
R4 P.n42 P.t60 6.1905
R5 P.n41 P.t35 6.1905
R6 P.n40 P.t23 6.1905
R7 P.n39 P.t39 6.1905
R8 P.n38 P.t3 6.1905
R9 P.n37 P.t72 6.1905
R10 P.n36 P.t27 6.1905
R11 P.n35 P.t84 6.1905
R12 P.n34 P.t13 6.1905
R13 P.n33 P.t51 6.1905
R14 P.n32 P.t80 6.1905
R15 P.n31 P.t45 6.1905
R16 P.n30 P.t19 6.1905
R17 P.n29 P.t56 6.1905
R18 P.n26 P.t10 6.1905
R19 P.n25 P.t11 6.1905
R20 P.n24 P.t36 6.1905
R21 P.n23 P.t37 6.1905
R22 P.n22 P.t48 6.1905
R23 P.n21 P.t49 6.1905
R24 P.n20 P.t67 6.1905
R25 P.n19 P.t68 6.1905
R26 P.n18 P.t32 6.1905
R27 P.n17 P.t33 6.1905
R28 P.n64 P.t61 6.1905
R29 P.n80 P.t28 6.1905
R30 P.n79 P.t73 6.1905
R31 P.n78 P.t0 6.1905
R32 P.n77 P.t81 6.1905
R33 P.n76 P.t46 6.1905
R34 P.n75 P.t40 6.1905
R35 P.n74 P.t53 6.1905
R36 P.n73 P.t42 6.1905
R37 P.n72 P.t24 6.1905
R38 P.n71 P.t69 6.1905
R39 P.n70 P.t65 6.1905
R40 P.n69 P.t77 6.1905
R41 P.n68 P.t87 6.1905
R42 P.n67 P.t8 6.1905
R43 P.n66 P.t75 6.1905
R44 P.n65 P.t14 6.1905
R45 P.n46 P.t62 6.1905
R46 P.n47 P.t15 6.1905
R47 P.n48 P.t76 6.1905
R48 P.n49 P.t9 6.1905
R49 P.n50 P.t88 6.1905
R50 P.n51 P.t78 6.1905
R51 P.n52 P.t66 6.1905
R52 P.n53 P.t70 6.1905
R53 P.n54 P.t25 6.1905
R54 P.n55 P.t43 6.1905
R55 P.n56 P.t54 6.1905
R56 P.n57 P.t41 6.1905
R57 P.n58 P.t47 6.1905
R58 P.n59 P.t82 6.1905
R59 P.n60 P.t1 6.1905
R60 P.n61 P.t74 6.1905
R61 P.n62 P.t29 6.1905
R62 P.n82 P.t7 6.1905
R63 P.n83 P.t6 6.1905
R64 P.n84 P.t86 6.1905
R65 P.n85 P.t85 6.1905
R66 P.n86 P.t17 6.1905
R67 P.n87 P.t16 6.1905
R68 P.n88 P.t21 6.1905
R69 P.n89 P.t20 6.1905
R70 P.n90 P.t5 6.1905
R71 P.n16 P.t57 6.1905
R72 P.n15 P.t63 6.1905
R73 P.n14 P.t59 6.1905
R74 P.n13 P.t34 6.1905
R75 P.n12 P.t22 6.1905
R76 P.n11 P.t38 6.1905
R77 P.n10 P.t2 6.1905
R78 P.n9 P.t71 6.1905
R79 P.n8 P.t26 6.1905
R80 P.n7 P.t83 6.1905
R81 P.n6 P.t12 6.1905
R82 P.n5 P.t50 6.1905
R83 P.n4 P.t79 6.1905
R84 P.n3 P.t44 6.1905
R85 P.n2 P.t18 6.1905
R86 P.n1 P.t55 6.1905
R87 P.n0 P.t30 6.1905
R88 P P.n93 4.949
R89 P.n93 P.t52 3.49604
R90 P.n81 P.n62 1.2155
R91 P.n45 P.n16 1.2155
R92 P.n89 P.n88 1.20532
R93 P.n87 P.n86 1.20532
R94 P.n85 P.n84 1.20532
R95 P.n83 P.n82 1.20532
R96 P.n18 P.n17 1.20532
R97 P.n20 P.n19 1.20532
R98 P.n22 P.n21 1.20532
R99 P.n24 P.n23 1.20532
R100 P.n26 P.n25 1.20532
R101 P.n91 P.n90 1.19574
R102 P.n47 P.n46 0.587457
R103 P.n48 P.n47 0.587457
R104 P.n49 P.n48 0.587457
R105 P.n50 P.n49 0.587457
R106 P.n51 P.n50 0.587457
R107 P.n52 P.n51 0.587457
R108 P.n53 P.n52 0.587457
R109 P.n54 P.n53 0.587457
R110 P.n55 P.n54 0.587457
R111 P.n56 P.n55 0.587457
R112 P.n57 P.n56 0.587457
R113 P.n58 P.n57 0.587457
R114 P.n59 P.n58 0.587457
R115 P.n60 P.n59 0.587457
R116 P.n61 P.n60 0.587457
R117 P.n62 P.n61 0.587457
R118 P.n65 P.n64 0.587457
R119 P.n66 P.n65 0.587457
R120 P.n67 P.n66 0.587457
R121 P.n68 P.n67 0.587457
R122 P.n69 P.n68 0.587457
R123 P.n70 P.n69 0.587457
R124 P.n71 P.n70 0.587457
R125 P.n72 P.n71 0.587457
R126 P.n73 P.n72 0.587457
R127 P.n74 P.n73 0.587457
R128 P.n75 P.n74 0.587457
R129 P.n76 P.n75 0.587457
R130 P.n77 P.n76 0.587457
R131 P.n78 P.n77 0.587457
R132 P.n79 P.n78 0.587457
R133 P.n80 P.n79 0.587457
R134 P.n1 P.n0 0.587457
R135 P.n2 P.n1 0.587457
R136 P.n3 P.n2 0.587457
R137 P.n4 P.n3 0.587457
R138 P.n5 P.n4 0.587457
R139 P.n6 P.n5 0.587457
R140 P.n7 P.n6 0.587457
R141 P.n8 P.n7 0.587457
R142 P.n9 P.n8 0.587457
R143 P.n10 P.n9 0.587457
R144 P.n11 P.n10 0.587457
R145 P.n12 P.n11 0.587457
R146 P.n13 P.n12 0.587457
R147 P.n14 P.n13 0.587457
R148 P.n15 P.n14 0.587457
R149 P.n16 P.n15 0.587457
R150 P.n29 P.n28 0.587457
R151 P.n30 P.n29 0.587457
R152 P.n31 P.n30 0.587457
R153 P.n32 P.n31 0.587457
R154 P.n33 P.n32 0.587457
R155 P.n34 P.n33 0.587457
R156 P.n35 P.n34 0.587457
R157 P.n36 P.n35 0.587457
R158 P.n37 P.n36 0.587457
R159 P.n38 P.n37 0.587457
R160 P.n39 P.n38 0.587457
R161 P.n40 P.n39 0.587457
R162 P.n41 P.n40 0.587457
R163 P.n42 P.n41 0.587457
R164 P.n43 P.n42 0.587457
R165 P.n44 P.n43 0.587457
R166 P.n93 P.n92 0.54333
R167 P.n90 P.n89 0.274015
R168 P.n88 P.n87 0.274015
R169 P.n86 P.n85 0.274015
R170 P.n84 P.n83 0.274015
R171 P.n19 P.n18 0.274015
R172 P.n21 P.n20 0.274015
R173 P.n23 P.n22 0.274015
R174 P.n25 P.n24 0.274015
R175 P.n82 P.n81 0.264431
R176 P.n27 P.n26 0.264431
R177 P.n91 P.n45 0.254848
R178 P.n81 P.n80 0.0298478
R179 P.n45 P.n44 0.0298478
R180 P.n92 P.n91 0.0298478
R181 P.n64 P.n63 0.00441304
R182 P.n28 P.n27 0.00441304
R183 VDD.t11 VDD.t4 49.5054
R184 VDD.t4 VDD.t9 49.5054
R185 VDD.t9 VDD.t8 49.5054
R186 VDD.t1 VDD.t0 49.5054
R187 VDD.t10 VDD.t1 49.5054
R188 VDD.t3 VDD.t10 49.5054
R189 VDD.t16 VDD.t3 49.5054
R190 VDD.t16 VDD.t14 49.5054
R191 VDD.t14 VDD.t6 49.5054
R192 VDD.t6 VDD.t13 49.5054
R193 VDD.t13 VDD.t15 49.5054
R194 VDD.t5 VDD.t2 49.5054
R195 VDD.t12 VDD.t5 49.5054
R196 VDD.t7 VDD.t12 49.5054
R197 VDD.n0 VDD.t11 41.7644
R198 VDD.n6 VDD.t7 41.7644
R199 VDD.n5 VDD.n1 10.573
R200 VDD VDD.n7 10.171
R201 VDD.n7 VDD.n6 3.1505
R202 VDD.n3 VDD.n2 3.1505
R203 VDD.t16 VDD.n3 3.1505
R204 VDD.n1 VDD.n0 3.1505
R205 VDD.n4 VDD.t16 3.1505
R206 VDD.n5 VDD.n4 3.1505
R207 VDD VDD.n5 0.218882
R208 a_4414_3230.t0 a_4414_3230.t1 12.9675
R209 a_7114_2196.t0 a_7114_2196.t1 12.9675
R210 a_7414_1574.t0 a_7414_1574.t1 12.9675
R211 a_7714_3852.t0 a_7714_3852.t1 12.9675
R212 a_7414_3230.t0 a_7414_3230.t1 12.9675
R213 a_5914_540.t0 a_5914_540.t1 12.9675
R214 a_6214_n82.t0 a_6214_n82.t1 12.9675
R215 a_7414_3024.t0 a_7414_3024.t1 12.9675
R216 a_7714_2402.t0 a_7714_2402.t1 12.9675
R217 a_4414_3024.t0 a_4414_3024.t1 12.9675
R218 a_4414_2196.t0 a_4414_2196.t1 10.2205
R219 a_5314_540.t0 a_5314_540.t1 12.9675
R220 a_5014_n82.t0 a_5014_n82.t1 12.9675
R221 a_4414_540.t0 a_4414_540.t1 10.2205
R222 a_4414_n82.t0 a_4414_n82.t1 12.9675
R223 a_6514_2196.t0 a_6514_2196.t1 12.9675
R224 a_6814_1574.t0 a_6814_1574.t1 12.9675
R225 a_5314_3852.t0 a_5314_3852.t1 12.9675
R226 a_5014_3230.t0 a_5014_3230.t1 12.9675
R227 a_8314_3852.t0 a_8314_3852.t1 12.9675
R228 a_8614_3024.t0 a_8614_3024.t1 10.2205
R229 a_5014_1368.t0 a_5014_1368.t1 12.9675
R230 a_4714_746.t0 a_4714_746.t1 12.9675
R231 a_8314_2196.t0 a_8314_2196.t1 12.9675
R232 a_8014_1574.t0 a_8014_1574.t1 12.9675
R233 a_4714_2196.t0 a_4714_2196.t1 12.9675
R234 a_5014_1574.t0 a_5014_1574.t1 12.9675
R235 a_8314_540.t0 a_8314_540.t1 12.9675
R236 a_8014_n82.t0 a_8014_n82.t1 12.9675
R237 a_8314_2402.t0 a_8314_2402.t1 12.9675
R238 a_5014_3024.t0 a_5014_3024.t1 12.9675
R239 a_5314_2402.t0 a_5314_2402.t1 12.9675
R240 a_7114_540.t0 a_7114_540.t1 12.9675
R241 a_7414_n82.t0 a_7414_n82.t1 12.9675
R242 a_4414_1368.t0 a_4414_1368.t1 12.9675
R243 a_6514_540.t0 a_6514_540.t1 12.9675
R244 a_5314_746.t0 a_5314_746.t1 12.9675
R245 a_4714_3852.t0 a_4714_3852.t1 12.9675
R246 a_7714_2196.t0 a_7714_2196.t1 12.9675
R247 a_4414_1574.t0 a_4414_1574.t1 12.9675
R248 a_5614_n82.t0 a_5614_n82.t1 12.9675
R249 a_4714_2402.t0 a_4714_2402.t1 12.9675
R250 a_5914_3852.t0 a_5914_3852.t1 12.9675
R251 a_6214_3230.t0 a_6214_3230.t1 12.9675
R252 a_6214_1368.t0 a_6214_1368.t1 12.9675
R253 a_5914_746.t0 a_5914_746.t1 12.9675
R254 a_6214_3024.t0 a_6214_3024.t1 12.9675
R255 a_5914_2402.t0 a_5914_2402.t1 12.9675
R256 a_4714_540.t0 a_4714_540.t1 12.9675
R257 a_5614_1368.t0 a_5614_1368.t1 12.9675
R258 a_6814_1368.t0 a_6814_1368.t1 12.9675
R259 a_7114_746.t0 a_7114_746.t1 12.9675
R260 M M.t0 8.52434
R261 a_6514_746.t0 a_6514_746.t1 12.9675
R262 a_5614_3230.t0 a_5614_3230.t1 12.9675
R263 a_8014_1368.t0 a_8014_1368.t1 12.9675
R264 a_7714_746.t0 a_7714_746.t1 12.9675
R265 a_8614_1368.t0 a_8614_1368.t1 10.2205
R266 a_5314_2196.t0 a_5314_2196.t1 12.9675
R267 a_7714_540.t0 a_7714_540.t1 12.9675
R268 a_5614_3024.t0 a_5614_3024.t1 12.9675
R269 a_7114_3852.t0 a_7114_3852.t1 12.9675
R270 a_6814_3230.t0 a_6814_3230.t1 12.9675
R271 a_7414_1368.t0 a_7414_1368.t1 12.9675
R272 a_6814_3024.t0 a_6814_3024.t1 12.9675
R273 a_7114_2402.t0 a_7114_2402.t1 12.9675
R274 a_6814_n82.t0 a_6814_n82.t1 12.9675
R275 a_8314_746.t0 a_8314_746.t1 12.9675
R276 a_5914_2196.t0 a_5914_2196.t1 12.9675
R277 a_6214_1574.t0 a_6214_1574.t1 12.9675
R278 a_6514_3852.t0 a_6514_3852.t1 12.9675
R279 a_6514_2402.t0 a_6514_2402.t1 12.9675
R280 a_8014_3230.t0 a_8014_3230.t1 12.9675
R281 a_8014_3024.t0 a_8014_3024.t1 12.9675
R282 a_5614_1574.t0 a_5614_1574.t1 12.9675
C0 M P 0.217f
C1 M VDD 0.248f
C2 P VDD 20.4f
C3 M VSUBS 0.386f
C4 P VSUBS 10.6f
C5 VDD VSUBS 0.104p
C6 VDD.t8 VSUBS 1.05f
C7 VDD.t9 VSUBS 1.05f
C8 VDD.t4 VSUBS 1.05f
C9 VDD.t11 VSUBS 0.981f
C10 VDD.n0 VSUBS 0.806f
C11 VDD.n1 VSUBS 0.147f
C12 VDD.t0 VSUBS 1.05f
C13 VDD.t1 VSUBS 1.05f
C14 VDD.t10 VSUBS 1.05f
C15 VDD.t3 VSUBS 1.05f
C16 VDD.t15 VSUBS 1.05f
C17 VDD.t13 VSUBS 1.05f
C18 VDD.t6 VSUBS 1.05f
C19 VDD.t14 VSUBS 1.05f
C20 VDD.n2 VSUBS 0.149f
C21 VDD.n3 VSUBS 0.233f
C22 VDD.t16 VSUBS 1.05f
C23 VDD.n4 VSUBS 0.233f
C24 VDD.n5 VSUBS 0.0866f
C25 VDD.t2 VSUBS 1.05f
C26 VDD.t5 VSUBS 1.05f
C27 VDD.t12 VSUBS 1.05f
C28 VDD.t7 VSUBS 0.981f
C29 VDD.n6 VSUBS 0.806f
C30 VDD.n7 VSUBS 0.144f
C31 P.t4 VSUBS 0.0952f
C32 P.t30 VSUBS 0.0952f
C33 P.n0 VSUBS 0.173f
C34 P.t55 VSUBS 0.0952f
C35 P.n1 VSUBS 0.107f
C36 P.t18 VSUBS 0.0952f
C37 P.n2 VSUBS 0.107f
C38 P.t44 VSUBS 0.0952f
C39 P.n3 VSUBS 0.107f
C40 P.t79 VSUBS 0.0952f
C41 P.n4 VSUBS 0.107f
C42 P.t50 VSUBS 0.0952f
C43 P.n5 VSUBS 0.107f
C44 P.t12 VSUBS 0.0952f
C45 P.n6 VSUBS 0.107f
C46 P.t83 VSUBS 0.0952f
C47 P.n7 VSUBS 0.107f
C48 P.t26 VSUBS 0.0952f
C49 P.n8 VSUBS 0.107f
C50 P.t71 VSUBS 0.0952f
C51 P.n9 VSUBS 0.107f
C52 P.t2 VSUBS 0.0952f
C53 P.n10 VSUBS 0.107f
C54 P.t38 VSUBS 0.0952f
C55 P.n11 VSUBS 0.107f
C56 P.t22 VSUBS 0.0952f
C57 P.n12 VSUBS 0.107f
C58 P.t34 VSUBS 0.0952f
C59 P.n13 VSUBS 0.107f
C60 P.t59 VSUBS 0.0952f
C61 P.n14 VSUBS 0.107f
C62 P.t63 VSUBS 0.0952f
C63 P.n15 VSUBS 0.107f
C64 P.t57 VSUBS 0.0952f
C65 P.n16 VSUBS 0.171f
C66 P.t10 VSUBS 0.0952f
C67 P.t11 VSUBS 0.0952f
C68 P.t36 VSUBS 0.0952f
C69 P.t37 VSUBS 0.0952f
C70 P.t48 VSUBS 0.0952f
C71 P.t49 VSUBS 0.0952f
C72 P.t67 VSUBS 0.0952f
C73 P.t68 VSUBS 0.0952f
C74 P.t32 VSUBS 0.0952f
C75 P.t33 VSUBS 0.0952f
C76 P.n17 VSUBS 0.179f
C77 P.n18 VSUBS 0.18f
C78 P.n19 VSUBS 0.18f
C79 P.n20 VSUBS 0.18f
C80 P.n21 VSUBS 0.18f
C81 P.n22 VSUBS 0.18f
C82 P.n23 VSUBS 0.18f
C83 P.n24 VSUBS 0.18f
C84 P.n25 VSUBS 0.18f
C85 P.n26 VSUBS 0.179f
C86 P.n27 VSUBS 0.123f
C87 P.t31 VSUBS 0.0952f
C88 P.n28 VSUBS 0.0687f
C89 P.t56 VSUBS 0.0952f
C90 P.n29 VSUBS 0.107f
C91 P.t19 VSUBS 0.0952f
C92 P.n30 VSUBS 0.107f
C93 P.t45 VSUBS 0.0952f
C94 P.n31 VSUBS 0.107f
C95 P.t80 VSUBS 0.0952f
C96 P.n32 VSUBS 0.107f
C97 P.t51 VSUBS 0.0952f
C98 P.n33 VSUBS 0.107f
C99 P.t13 VSUBS 0.0952f
C100 P.n34 VSUBS 0.107f
C101 P.t84 VSUBS 0.0952f
C102 P.n35 VSUBS 0.107f
C103 P.t27 VSUBS 0.0952f
C104 P.n36 VSUBS 0.107f
C105 P.t72 VSUBS 0.0952f
C106 P.n37 VSUBS 0.107f
C107 P.t3 VSUBS 0.0952f
C108 P.n38 VSUBS 0.107f
C109 P.t39 VSUBS 0.0952f
C110 P.n39 VSUBS 0.107f
C111 P.t23 VSUBS 0.0952f
C112 P.n40 VSUBS 0.107f
C113 P.t35 VSUBS 0.0952f
C114 P.n41 VSUBS 0.107f
C115 P.t60 VSUBS 0.0952f
C116 P.n42 VSUBS 0.107f
C117 P.t64 VSUBS 0.0952f
C118 P.n43 VSUBS 0.107f
C119 P.t58 VSUBS 0.0952f
C120 P.n44 VSUBS 0.0703f
C121 P.n45 VSUBS 0.123f
C122 P.t5 VSUBS 0.0952f
C123 P.t20 VSUBS 0.0952f
C124 P.t21 VSUBS 0.0952f
C125 P.t16 VSUBS 0.0952f
C126 P.t17 VSUBS 0.0952f
C127 P.t85 VSUBS 0.0952f
C128 P.t86 VSUBS 0.0952f
C129 P.t6 VSUBS 0.0952f
C130 P.t7 VSUBS 0.0952f
C131 P.t62 VSUBS 0.0952f
C132 P.n46 VSUBS 0.173f
C133 P.t15 VSUBS 0.0952f
C134 P.n47 VSUBS 0.107f
C135 P.t76 VSUBS 0.0952f
C136 P.n48 VSUBS 0.107f
C137 P.t9 VSUBS 0.0952f
C138 P.n49 VSUBS 0.107f
C139 P.t88 VSUBS 0.0952f
C140 P.n50 VSUBS 0.107f
C141 P.t78 VSUBS 0.0952f
C142 P.n51 VSUBS 0.107f
C143 P.t66 VSUBS 0.0952f
C144 P.n52 VSUBS 0.107f
C145 P.t70 VSUBS 0.0952f
C146 P.n53 VSUBS 0.107f
C147 P.t25 VSUBS 0.0952f
C148 P.n54 VSUBS 0.107f
C149 P.t43 VSUBS 0.0952f
C150 P.n55 VSUBS 0.107f
C151 P.t54 VSUBS 0.0952f
C152 P.n56 VSUBS 0.107f
C153 P.t41 VSUBS 0.0952f
C154 P.n57 VSUBS 0.107f
C155 P.t47 VSUBS 0.0952f
C156 P.n58 VSUBS 0.107f
C157 P.t82 VSUBS 0.0952f
C158 P.n59 VSUBS 0.107f
C159 P.t1 VSUBS 0.0952f
C160 P.n60 VSUBS 0.107f
C161 P.t74 VSUBS 0.0952f
C162 P.n61 VSUBS 0.107f
C163 P.t29 VSUBS 0.0952f
C164 P.n62 VSUBS 0.171f
C165 P.n63 VSUBS 0.124f
C166 P.t61 VSUBS 0.0952f
C167 P.n64 VSUBS 0.0687f
C168 P.t14 VSUBS 0.0952f
C169 P.n65 VSUBS 0.107f
C170 P.t75 VSUBS 0.0952f
C171 P.n66 VSUBS 0.107f
C172 P.t8 VSUBS 0.0952f
C173 P.n67 VSUBS 0.107f
C174 P.t87 VSUBS 0.0952f
C175 P.n68 VSUBS 0.107f
C176 P.t77 VSUBS 0.0952f
C177 P.n69 VSUBS 0.107f
C178 P.t65 VSUBS 0.0952f
C179 P.n70 VSUBS 0.107f
C180 P.t69 VSUBS 0.0952f
C181 P.n71 VSUBS 0.107f
C182 P.t24 VSUBS 0.0952f
C183 P.n72 VSUBS 0.107f
C184 P.t42 VSUBS 0.0952f
C185 P.n73 VSUBS 0.107f
C186 P.t53 VSUBS 0.0952f
C187 P.n74 VSUBS 0.107f
C188 P.t40 VSUBS 0.0952f
C189 P.n75 VSUBS 0.107f
C190 P.t46 VSUBS 0.0952f
C191 P.n76 VSUBS 0.107f
C192 P.t81 VSUBS 0.0952f
C193 P.n77 VSUBS 0.107f
C194 P.t0 VSUBS 0.0952f
C195 P.n78 VSUBS 0.107f
C196 P.t73 VSUBS 0.0952f
C197 P.n79 VSUBS 0.107f
C198 P.t28 VSUBS 0.0952f
C199 P.n80 VSUBS 0.0703f
C200 P.n81 VSUBS 0.124f
C201 P.n82 VSUBS 0.179f
C202 P.n83 VSUBS 0.18f
C203 P.n84 VSUBS 0.18f
C204 P.n85 VSUBS 0.18f
C205 P.n86 VSUBS 0.18f
C206 P.n87 VSUBS 0.18f
C207 P.n88 VSUBS 0.18f
C208 P.n89 VSUBS 0.18f
C209 P.n90 VSUBS 0.179f
C210 P.n91 VSUBS 0.121f
C211 P.n92 VSUBS 0.0679f
C212 P.t52 VSUBS 0.0721f
C213 P.n93 VSUBS 0.301f
.ends

