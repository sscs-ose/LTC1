magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2692 -2128 2692 2128
<< nwell >>
rect -692 -128 692 128
<< nsubdiff >>
rect -609 23 609 45
rect -609 -23 -587 23
rect 587 -23 609 23
rect -609 -45 609 -23
<< nsubdiffcont >>
rect -587 -23 587 23
<< metal1 >>
rect -598 23 598 34
rect -598 -23 -587 23
rect 587 -23 598 23
rect -598 -34 598 -23
<< end >>
