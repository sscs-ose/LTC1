magic
tech gf180mcuC
magscale 1 10
timestamp 1692080300
<< error_p >>
rect -162 83 -151 129
rect 54 83 65 129
rect -239 -48 -193 48
rect -23 -48 23 48
rect 193 -48 239 48
rect -162 -129 -151 -83
rect 54 -129 65 -83
<< nwell >>
rect -414 -258 414 258
<< pmos >>
rect -164 -50 -52 50
rect 52 -50 164 50
<< pdiff >>
rect -252 37 -164 50
rect -252 -37 -239 37
rect -193 -37 -164 37
rect -252 -50 -164 -37
rect -52 37 52 50
rect -52 -37 -23 37
rect 23 -37 52 37
rect -52 -50 52 -37
rect 164 37 252 50
rect 164 -37 193 37
rect 239 -37 252 37
rect 164 -50 252 -37
<< pdiffc >>
rect -239 -37 -193 37
rect -23 -37 23 37
rect 193 -37 239 37
<< nsubdiff >>
rect -390 162 390 234
rect -390 118 -318 162
rect -390 -118 -377 118
rect -331 -118 -318 118
rect 318 118 390 162
rect -390 -162 -318 -118
rect 318 -118 331 118
rect 377 -118 390 118
rect 318 -162 390 -118
rect -390 -234 390 -162
<< nsubdiffcont >>
rect -377 -118 -331 118
rect 331 -118 377 118
<< polysilicon >>
rect -164 129 -52 142
rect -164 83 -151 129
rect -65 83 -52 129
rect -164 50 -52 83
rect 52 129 164 142
rect 52 83 65 129
rect 151 83 164 129
rect 52 50 164 83
rect -164 -83 -52 -50
rect -164 -129 -151 -83
rect -65 -129 -52 -83
rect -164 -142 -52 -129
rect 52 -83 164 -50
rect 52 -129 65 -83
rect 151 -129 164 -83
rect 52 -142 164 -129
<< polycontact >>
rect -151 83 -65 129
rect 65 83 151 129
rect -151 -129 -65 -83
rect 65 -129 151 -83
<< metal1 >>
rect -377 175 377 221
rect -377 118 -331 175
rect -162 83 -151 129
rect -65 83 -54 129
rect 54 83 65 129
rect 151 83 162 129
rect 331 118 377 175
rect -239 37 -193 48
rect -239 -48 -193 -37
rect -23 37 23 48
rect -23 -48 23 -37
rect 193 37 239 48
rect 193 -48 239 -37
rect -377 -175 -331 -118
rect -162 -129 -151 -83
rect -65 -129 -54 -83
rect 54 -129 65 -83
rect 151 -129 162 -83
rect 331 -175 377 -118
rect -377 -221 377 -175
<< properties >>
string FIXED_BBOX -354 -198 354 198
string gencell pmos_3p3
string library gf180mcu
string parameters w 0.5 l 0.560 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
