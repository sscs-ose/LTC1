* NGSPICE file created from CLK_div_108_new_mag_flat.ext - technology: gf180mcuC

.subckt CLK_div_108_new_mag_flat VDD VSS RST Vdiv108 CLK
X0 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t78 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X1 a_11440_215# RST.t0 a_11280_215# VSS.t173 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2 VDD VDD.t171 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VDD.t172 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X3 a_13857_4607# VDD.t453 VSS.t115 VSS.t114 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X4 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_18289_4654# VSS.t65 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X5 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t315 VDD.t314 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X6 a_18853_4654# JK_FF_mag_0.nand2_mag_1.IN2 VSS.t239 VSS.t238 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X7 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.QB a_14017_4607# VSS.t191 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X8 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.CLK.t2 VDD.t429 VDD.t428 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X9 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.CLK.t3 VDD.t404 VDD.t403 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X10 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t360 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X11 a_17846_214# RST.t1 a_17686_214# VSS.t172 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X12 VSS CLK_div_3_mag_1.CLK.t4 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t254 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X13 a_18289_4654# JK_FF_mag_0.nand3_mag_1.IN1 VSS.t251 VSS.t250 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X14 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t61 VDD.t60 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X15 JK_FF_mag_1.QB JK_FF_mag_1.Q a_15863_3554# VSS.t269 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X16 VDD CLK_div_3_mag_2.JK_FF_mag_1.K.t2 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VDD.t107 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X17 VSS VDD.t454 a_9147_215# VSS.t111 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X18 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t329 VDD.t328 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X19 VSS CLK.t0 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VSS.t85 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X20 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK.t1 VDD.t132 VDD.t131 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X21 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 a_10674_5199# VSS.t120 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X22 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.Q0 VDD.t180 VDD.t179 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X23 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t381 VDD.t380 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X24 VDD CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t220 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD.t305 VDD.t304 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X26 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t449 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X27 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t400 VDD.t399 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X28 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_15299_3554# VSS.t54 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X29 VSS CLK_div_3_mag_1.CLK.t5 a_8705_2455# VSS.t257 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X30 a_7699_259# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t26 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X31 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 a_11398_5199# VSS.t21 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X32 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t34 VDD.t33 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X33 a_15863_3554# JK_FF_mag_1.nand2_mag_4.IN2 VSS.t43 VSS.t42 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X34 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK.t2 VDD.t229 VDD.t228 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 a_11962_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS.t137 VSS.t136 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X36 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t227 VDD.t226 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X37 VSS CLK.t3 a_15111_2454# VSS.t138 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X38 VSS VDD.t455 a_15553_214# VSS.t108 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X39 a_10674_5199# CLK_div_3_mag_0.CLK.t2 a_10514_5199# VSS.t237 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X40 VDD CLK_div_3_mag_0.CLK.t3 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t181 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X41 a_8227_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS.t41 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X42 JK_FF_mag_1.nand3_mag_2.OUT VDD.t168 VDD.t170 VDD.t169 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X43 a_17122_258# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t178 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X44 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t251 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X45 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.Q0.t0 VDD.t377 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X46 VDD RST.t2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t254 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X47 VSS CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.or_2_mag_0.IN2 VSS.t145 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X48 a_9141_1312# CLK_div_3_mag_1.CLK.t6 a_8981_1312# VSS.t260 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X49 a_12164_215# CLK_div_3_mag_1.CLK.t7 a_12004_215# VSS.t261 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X50 a_9355_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t233 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X51 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q1 a_10956_3003# VSS.t81 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X52 JK_FF_mag_0.nand3_mag_2.OUT VDD.t165 VDD.t167 VDD.t166 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X53 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 VDD.t101 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X54 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS.t189 VSS.t188 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X55 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t35 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X56 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t195 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X57 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT VDD.t204 VDD.t203 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X58 VDD CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.IN2 VDD.t371 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X59 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.Q1.t3 VDD.t82 VDD.t81 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X60 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.Q1.t0 VDD.t104 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X61 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.JK_FF_mag_1.K.t3 VDD.t111 VDD.t110 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X62 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VDD.t290 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X63 VSS CLK_div_3_mag_2.JK_FF_mag_1.K.t4 a_18564_1311# VSS.t69 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X64 JK_FF_mag_0.nand3_mag_2.OUT Vdiv108.t3 VDD.t317 VDD.t316 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X65 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VDD.t325 VDD.t324 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X66 VDD CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.CLK.t0 VDD.t441 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X67 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t327 VDD.t326 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X68 a_18570_214# CLK.t4 a_18410_214# VSS.t141 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X69 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.Q1.t4 VDD.t84 VDD.t83 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X70 a_7732_2691# CLK_div_3_mag_1.Q0.t3 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD.t432 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X71 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.Q1.t3 VDD.t116 VDD.t115 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X72 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X73 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 a_17879_3513# VSS.t249 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X74 a_14138_2690# CLK_div_3_mag_2.Q0.t3 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VDD.t348 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X75 a_7135_259# CLK_div_3_mag_1.Q0.t4 CLK_div_3_mag_1.JK_FF_mag_1.K VSS.t272 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X76 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t88 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X77 a_13541_258# CLK_div_3_mag_2.Q0.t4 CLK_div_3_mag_2.JK_FF_mag_1.K VSS.t213 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X78 a_18564_1311# CLK.t5 a_18404_1311# VSS.t142 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X79 VDD CLK_div_3_mag_0.CLK.t4 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t184 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X80 VDD VDD.t161 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t162 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 a_13851_3510# VDD.t457 VSS.t107 VSS.t106 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X82 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t223 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X83 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t4 a_10680_4102# VSS.t91 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X84 a_17879_3513# RST.t3 a_17719_3513# VSS.t171 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X85 VSS CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.CLK.t1 VSS.t281 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X86 VDD VDD.t157 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VDD.t158 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X87 a_16995_3513# VDD.t459 VSS.t105 VSS.t104 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X88 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT a_8423_215# VSS.t123 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X89 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11808_4102# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X90 a_8417_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t195 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X91 VSS CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT a_14829_214# VSS.t179 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X92 JK_FF_mag_0.nand3_mag_2.OUT Vdiv108.t4 a_17155_3513# VSS.t199 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X93 a_10680_4102# CLK_div_3_mag_0.CLK.t5 a_10520_4102# VSS.t91 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X94 JK_FF_mag_1.Q JK_FF_mag_1.nand2_mag_1.IN2 VDD.t431 VDD.t430 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X95 VSS CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_17840_1355# VSS.t219 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X96 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_11244_4102# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X97 a_16712_1355# CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.Q1.t1 VSS.t16 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X98 VDD JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t49 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X99 a_10716_259# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t198 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X100 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t311 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X101 VSS VDD.t460 a_12164_215# VSS.t101 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X102 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand3_mag_1.IN1 VDD.t393 VDD.t392 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X103 JK_FF_mag_1.CLK CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD.t402 VDD.t401 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X104 VSS CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_14105_258# VSS.t288 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X105 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t93 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X106 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t70 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X107 VSS VDD.t461 a_18570_214# VSS.t98 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X108 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VDD.t92 VDD.t91 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X109 VSS CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 a_13695_1355# VSS.t230 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X110 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t345 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X111 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_10870_1356# VSS.t150 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X112 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t289 VDD.t288 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X113 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_18443_3557# VSS.t64 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X114 VSS CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_14823_1355# VSS.t22 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X115 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0 a_12526_5199# VSS.t119 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X116 VDD CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VDD.t176 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X117 a_15299_3554# JK_FF_mag_1.nand3_mag_1.OUT VSS.t127 VSS.t54 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X118 a_8705_2455# CLK_div_3_mag_1.Q1.t5 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS.t55 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X119 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_10306_1356# VSS.t66 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X120 a_13695_1355# CLK_div_3_mag_2.JK_FF_mag_1.K.t5 CLK_div_3_mag_2.Q0.t2 VSS.t72 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X121 a_10152_259# CLK_div_3_mag_1.Q1.t6 CLK_div_3_mag_1.JK_FF_mag_1.QB VSS.t56 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X122 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VDD.t205 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X123 a_11398_5199# RST.t4 a_11238_5199# VSS.t170 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X124 VDD RST.t5 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD.t366 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X125 VDD CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VDD.t24 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X126 a_10870_1356# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t197 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X127 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K.t0 VDD.t387 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X128 a_15111_2454# CLK_div_3_mag_2.Q1.t4 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VSS.t74 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X129 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.K.t1 VDD.t374 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X130 a_10514_5199# VDD.t462 VSS.t97 VSS.t96 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X131 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11962_5199# VSS.t57 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X132 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t154 VDD.t156 VDD.t155 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X133 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t85 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X134 a_11929_2535# CLK_div_3_mag_0.or_2_mag_0.IN2 VDD.t338 VDD.t337 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X135 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_11434_1356# VSS.t0 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X136 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_4.IN2 VDD.t97 VDD.t96 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X137 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT VDD.t126 VDD.t125 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X138 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t275 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X139 VDD CLK_div_3_mag_2.Q0.t5 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VDD.t353 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X140 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT a_14581_4651# VSS.t126 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X141 JK_FF_mag_1.CLK CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t253 VSS.t252 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X142 VDD CLK_div_3_mag_2.Q1.t5 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VDD.t117 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X143 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t48 VDD.t47 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X144 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t6 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X145 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VDD.t448 VDD.t447 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X146 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT a_11440_215# VSS.t210 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X147 VDD CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t208 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X148 VDD JK_FF_mag_1.Q JK_FF_mag_0.nand3_mag_2.OUT VDD.t425 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X149 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t140 VDD.t139 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X150 VDD CLK_div_3_mag_1.JK_FF_mag_1.K.t2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VDD.t44 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X151 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.Q1.t6 VDD.t121 VDD.t120 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X152 JK_FF_mag_1.Q JK_FF_mag_1.QB a_15709_4651# VSS.t190 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X153 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT a_17725_4654# VSS.t33 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X154 VDD Vdiv108.t5 JK_FF_mag_0.QB VDD.t330 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X155 VSS CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.IN2 VSS.t224 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X156 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0 a_11929_2535# VDD.t175 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X157 VDD CLK_div_3_mag_1.CLK.t8 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t405 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X158 a_14581_4651# JK_FF_mag_1.nand3_mag_0.OUT VSS.t52 VSS.t51 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X159 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t56 VDD.t55 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X160 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t342 VDD.t341 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X161 VSS CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_17846_214# VSS.t128 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X162 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_15145_4651# VSS.t53 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X163 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK.t6 VDD.t188 VDD.t187 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X164 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t32 VDD.t31 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X165 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t52 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X166 a_18404_1311# CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VSS.t15 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X167 VDD CLK_div_3_mag_0.CLK.t7 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD.t189 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X168 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 VDD.t219 VDD.t218 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X169 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.CLK.t9 VDD.t409 VDD.t408 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X170 VDD CLK_div_3_mag_0.JK_FF_mag_1.K.t5 CLK_div_3_mag_0.Q0 VDD.t243 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X171 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD.t334 VDD.t333 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X172 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.CLK VSS.t12 VSS.t11 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X173 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB a_7663_4102# VSS.t91 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X174 a_17719_3513# JK_FF_mag_0.nand3_mag_2.OUT VSS.t79 VSS.t78 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X175 a_15393_214# CLK_div_3_mag_2.Q0.t6 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VSS.t216 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X176 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT a_7699_259# VSS.t192 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X177 VSS CLK_div_3_mag_2.Q1.t7 a_15547_1311# VSS.t75 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X178 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.or_2_mag_0.IN2 VSS.t204 VSS.t116 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X179 a_11808_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t20 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X180 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD.t344 VDD.t343 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X181 a_11998_1312# CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS.t132 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X182 VSS CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_17122_258# VSS.t59 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X183 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.CLK.t10 VDD.t411 VDD.t410 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X184 a_17155_3513# JK_FF_mag_1.Q a_16995_3513# VSS.t268 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X185 VSS CLK_div_3_mag_1.JK_FF_mag_1.K.t3 a_12158_1312# VSS.t28 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X186 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_1.Q VDD.t424 VDD.t423 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X187 a_7663_4102# CLK_div_3_mag_0.CLK.t8 a_7503_4102# VSS.t91 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X188 a_10520_4102# CLK_div_3_mag_0.Q1 VSS.t135 VSS.t91 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X189 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 a_12372_4102# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X190 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t391 VDD.t390 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X191 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VDD.t272 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X192 VSS CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_17276_1355# VSS.t48 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X193 JK_FF_mag_0.nand3_mag_0.OUT VDD.t151 VDD.t153 VDD.t152 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X194 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VDD.t3 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X195 a_17840_1355# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t58 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X196 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB VDD.t12 VDD.t11 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X197 VDD JK_FF_mag_0.QB Vdiv108.t1 VDD.t9 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X198 a_11244_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS.t201 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X199 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT VDD.t258 VDD.t257 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X200 VDD CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.CLK.t0 VDD.t264 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X201 a_12158_1312# CLK_div_3_mag_1.CLK.t11 a_11998_1312# VSS.t262 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X202 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT CLK.t6 VDD.t231 VDD.t230 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X203 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB VDD.t382 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X204 a_12372_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t207 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X205 a_17276_1355# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VSS.t177 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X206 a_17001_4610# VDD.t463 VSS.t95 VSS.t94 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X207 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK.t9 VSS.t122 VSS.t121 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X208 VDD JK_FF_mag_1.Q JK_FF_mag_0.nand3_mag_0.OUT VDD.t420 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X209 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.QB a_17161_4610# VSS.t8 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X210 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 a_7135_259# VSS.t240 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X211 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 VDD.t217 VDD.t216 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X212 VSS CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 a_13541_258# VSS.t227 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X213 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.QB VDD.t269 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X214 VDD CLK_div_3_mag_1.Q0.t5 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t281 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X215 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.Q1 a_7657_5199# VSS.t134 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X216 a_9147_215# CLK_div_3_mag_1.CLK.t12 a_8987_215# VSS.t263 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X217 a_19007_3557# JK_FF_mag_0.nand2_mag_4.IN2 VSS.t63 VSS.t62 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X218 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 a_7853_1356# VSS.t163 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X219 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_8381_5199# VSS.t215 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X220 a_8945_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS.t187 VSS.t186 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X221 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t352 VDD.t351 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X222 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t303 VDD.t302 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X223 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 a_14735_3510# VSS.t245 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X224 VSS CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.CLK.t1 VSS.t156 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X225 a_8263_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS.t162 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X226 VDD CLK_div_3_mag_2.Q1.t8 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VDD.t122 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X227 a_17161_4610# JK_FF_mag_1.Q a_17001_4610# VSS.t267 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X228 VDD CLK_div_3_mag_0.CLK.t10 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t192 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X229 a_18443_3557# JK_FF_mag_0.nand3_mag_1.OUT VSS.t32 VSS.t31 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X230 VDD CLK.t7 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t232 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X231 a_14669_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VSS.t6 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X232 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t340 VDD.t339 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X233 a_14823_1355# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VSS.t287 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X234 VSS CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_14259_1355# VSS.t3 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X235 a_7657_5199# CLK_div_3_mag_0.CLK.t11 a_7497_5199# VSS.t80 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X236 a_12526_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t223 VSS.t222 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X237 VDD CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD.t213 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X238 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD.t370 VDD.t369 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X239 a_10306_1356# CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.Q1.t2 VSS.t131 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X240 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 a_9509_5199# VSS.t133 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X241 a_11238_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS.t203 VSS.t202 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X242 VDD RST.t6 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VDD.t363 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X243 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VDD.t336 VDD.t335 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X244 a_16558_258# CLK_div_3_mag_2.Q1.t9 CLK_div_3_mag_2.JK_FF_mag_1.QB VSS.t208 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X245 a_15553_214# CLK.t8 a_15393_214# VSS.t143 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X246 a_8381_5199# RST.t7 a_8221_5199# VSS.t169 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X247 JK_FF_mag_0.QB Vdiv108.t6 a_19007_3557# VSS.t200 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X248 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t321 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X249 a_11434_1356# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t37 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X250 a_14259_1355# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t206 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X251 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_8945_5199# VSS.t196 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X252 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.Q0.t1 VDD.t133 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X253 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t41 VDD.t40 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X254 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_10716_259# VSS.t34 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X255 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK.t9 VDD.t236 VDD.t235 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X256 a_8987_215# CLK_div_3_mag_1.Q0.t6 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS.t174 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X257 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT RST.t8 VDD.t268 VDD.t267 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X258 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD.t318 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X259 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VDD.t57 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X260 VDD CLK_div_3_mag_1.JK_FF_mag_1.K.t4 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t259 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X261 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT RST.t9 VDD.t199 VDD.t198 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X262 Vdiv108 JK_FF_mag_0.QB a_18853_4654# VSS.t7 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X263 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 VDD.t263 VDD.t262 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X264 a_18410_214# CLK_div_3_mag_2.Q1.t10 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VSS.t209 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X265 a_15709_4651# JK_FF_mag_1.nand2_mag_1.IN2 VSS.t271 VSS.t270 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X266 a_17725_4654# JK_FF_mag_0.nand3_mag_0.OUT VSS.t154 VSS.t153 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X267 VDD CLK_div_3_mag_1.Q1.t7 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VDD.t293 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X268 VDD CLK_div_3_mag_1.CLK.t13 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t412 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X269 VDD CLK_div_3_mag_2.JK_FF_mag_1.K.t6 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VDD.t112 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X270 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VDD.t248 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X271 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.Q1.t2 VDD.t64 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X272 VSS CLK_div_3_mag_1.CLK.t14 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t284 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X273 a_15145_4651# JK_FF_mag_1.nand3_mag_1.IN1 VSS.t244 VSS.t243 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X274 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t299 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X275 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VDD.t350 VDD.t349 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X276 VDD CLK.t10 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t237 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X277 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK.t12 VDD.t128 VDD.t127 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X278 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VDD.t247 VDD.t246 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X279 VSS CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS.t246 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X280 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.CLK.t13 VDD.t130 VDD.t129 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X281 VDD CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 VDD.t136 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X282 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VDD.t67 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X283 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 a_8791_4102# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X284 VSS CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS.t116 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X285 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_1.Q VSS.t266 VSS.t265 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X286 VSS CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VSS.t278 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X287 VSS CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 a_10152_259# VSS.t234 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X288 a_15547_1311# CLK.t11 a_15387_1311# VSS.t144 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X289 a_8423_215# RST.t10 a_8263_215# VSS.t168 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X290 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT a_8227_4102# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X291 VDD JK_FF_mag_1.CLK JK_FF_mag_1.nand3_mag_2.OUT VDD.t19 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X292 a_8981_1312# CLK_div_3_mag_1.JK_FF_mag_1.K.t6 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS.t155 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X293 a_14829_214# RST.t11 a_14669_214# VSS.t167 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X294 a_8791_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS.t214 VSS.t19 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X295 VDD JK_FF_mag_1.Q JK_FF_mag_1.QB VDD.t417 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X296 a_10956_3003# CLK_div_3_mag_0.CLK.t14 VSS.t82 VSS.t81 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X297 VDD CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.or_2_mag_0.IN2 VDD.t240 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X298 a_7503_4102# CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS.t148 VSS.t91 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X299 VDD RST.t12 JK_FF_mag_1.nand3_mag_1.OUT VDD.t278 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X300 VSS CLK_div_3_mag_1.Q1.t8 a_9141_1312# VSS.t182 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X301 VSS CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_16558_258# VSS.t159 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X302 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t98 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X303 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.QB a_9355_4102# VSS.t19 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X304 a_11280_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS.t149 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X305 a_15387_1311# CLK_div_3_mag_2.JK_FF_mag_1.K.t7 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VSS.t73 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X306 Vdiv108 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t386 VDD.t385 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X307 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.Q0.t7 VSS.t176 VSS.t175 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X308 VDD CLK_div_3_mag_1.Q1.t9 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VDD.t296 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X309 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 VDD.t75 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X310 VDD CLK_div_3_mag_1.CLK.t15 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD.t444 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X311 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VDD.t39 VDD.t38 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X312 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.Q VDD.t416 VDD.t415 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X313 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_4.IN2 VDD.t63 VDD.t62 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X314 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.Q0.t7 VSS.t218 VSS.t217 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X315 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_2.OUT VDD.t434 VDD.t433 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X316 VDD CLK_div_3_mag_1.or_2_mag_0.IN2 a_7732_2691# VDD.t394 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X317 a_17686_214# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VSS.t47 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X318 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 VDD.t398 VDD.t397 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X319 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.CLK.t15 VSS.t84 VSS.t83 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X320 VDD CLK.t12 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VDD.t435 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X321 a_14105_258# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VSS.t205 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X322 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VDD.t287 VDD.t286 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X323 VDD CLK_div_3_mag_2.or_2_mag_0.IN2 a_14138_2690# VDD.t438 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X324 a_14011_3510# JK_FF_mag_1.CLK a_13851_3510# VSS.t10 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X325 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT RST.t13 VDD.t285 VDD.t284 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X326 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 a_7289_1356# VSS.t88 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X327 a_7853_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS.t25 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X328 a_14735_3510# RST.t14 a_14575_3510# VSS.t166 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X329 VDD JK_FF_mag_1.CLK JK_FF_mag_1.nand3_mag_0.OUT VDD.t16 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X330 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t148 VDD.t150 VDD.t149 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X331 a_12004_215# CLK_div_3_mag_1.Q1.t10 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS.t185 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X332 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT RST.t15 VDD.t359 VDD.t358 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X333 a_7497_5199# VDD.t464 VSS.t93 VSS.t92 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X334 VDD JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t200 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X335 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD.t23 VDD.t22 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X336 VSS CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT a_8417_1356# VSS.t38 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X337 VDD VDD.t144 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VDD.t145 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X338 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.Q0.t8 VDD.t43 VDD.t42 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X339 a_9509_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS.t14 VSS.t13 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X340 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.CLK VDD.t15 VDD.t14 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X341 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VDD.t30 VDD.t29 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X342 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.Q a_14011_3510# VSS.t264 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X343 a_7289_1356# CLK_div_3_mag_1.JK_FF_mag_1.K.t7 CLK_div_3_mag_1.Q0.t0 VSS.t27 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X344 VSS CLK.t13 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VSS.t275 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X345 a_8221_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS.t18 VSS.t17 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X346 JK_FF_mag_1.nand3_mag_0.OUT VDD.t141 VDD.t143 VDD.t142 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X347 a_14575_3510# JK_FF_mag_1.nand3_mag_2.OUT VSS.t274 VSS.t273 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X348 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.Q0.t8 VDD.t357 VDD.t356 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X349 VDD JK_FF_mag_1.QB JK_FF_mag_1.Q VDD.t308 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X350 a_14017_4607# JK_FF_mag_1.CLK a_13857_4607# VSS.t9 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X351 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.QB VDD.t307 VDD.t306 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X352 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT VDD.t74 VDD.t73 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X353 VSS CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 a_16712_1355# VSS.t44 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
R0 VDD.n157 VDD.t356 107239
R1 VDD.n352 VDD.t42 107239
R2 VDD.t149 VDD.n260 57397.6
R3 VDD.n350 VDD.n334 4006.3
R4 VDD.n155 VDD.n139 4006.3
R5 VDD.n157 VDD.n137 3116.02
R6 VDD.n352 VDD.n332 3116.02
R7 VDD.n156 VDD.n137 2331.49
R8 VDD.n351 VDD.n332 2331.49
R9 VDD.n156 VDD.n155 1668.51
R10 VDD.n351 VDD.n350 1668.51
R11 VDD.t290 VDD.t353 1164.27
R12 VDD.t374 VDD.t339 1164.27
R13 VDD.t195 VDD.t281 1164.27
R14 VDD.t387 VDD.t38 1164.27
R15 VDD.t449 VDD.n156 1046.11
R16 VDD.t311 VDD.n351 1046.11
R17 VDD.t321 VDD.t22 961.905
R18 VDD.t216 VDD.t29 961.905
R19 VDD.n260 VDD.t302 864.287
R20 VDD.t78 VDD.t430 765.152
R21 VDD.t392 VDD.t200 765.152
R22 VDD.t306 VDD.t73 765.152
R23 VDD.t385 VDD.t98 765.152
R24 VDD.t49 VDD.t397 765.152
R25 VDD.t257 VDD.t11 765.152
R26 VDD.t101 VDD.t96 765.152
R27 VDD.t399 VDD.t47 765.152
R28 VDD.t316 VDD.t125 765.152
R29 VDD.t360 VDD.t24 765.152
R30 VDD.t70 VDD.t91 765.152
R31 VDD.t64 VDD.t288 765.152
R32 VDD.t345 VDD.t296 765.152
R33 VDD.t52 VDD.t248 765.152
R34 VDD.t382 VDD.t328 765.152
R35 VDD.t0 VDD.t208 765.152
R36 VDD.t55 VDD.t251 765.152
R37 VDD.t104 VDD.t326 765.152
R38 VDD.t318 VDD.t380 765.152
R39 VDD.t299 VDD.t349 765.152
R40 VDD.t139 VDD.t60 765.152
R41 VDD.t259 VDD.t57 765.152
R42 VDD.t275 VDD.t314 765.152
R43 VDD.t133 VDD.t40 765.152
R44 VDD.t88 VDD.t343 765.152
R45 VDD.t31 VDD.t223 765.152
R46 VDD.t324 VDD.t333 765.152
R47 VDD.t85 VDD.t369 765.152
R48 VDD.t33 VDD.t226 765.152
R49 VDD.t179 VDD.t335 765.152
R50 VDD.t112 VDD.t35 765.152
R51 VDD.t447 VDD.t6 765.152
R52 VDD.t341 VDD.t377 765.152
R53 VDD.t205 VDD.t122 765.152
R54 VDD.t67 VDD.t93 765.152
R55 VDD.t269 VDD.t286 765.152
R56 VDD.t75 VDD.t62 765.152
R57 VDD.t390 VDD.t203 765.152
R58 VDD.t415 VDD.t433 765.152
R59 VDD.t230 VDD.t172 461.096
R60 VDD.t353 VDD.t230 461.096
R61 VDD.t198 VDD.t290 461.096
R62 VDD.t3 VDD.t198 461.096
R63 VDD.t339 VDD.t449 461.096
R64 VDD.t356 VDD.t374 461.096
R65 VDD.t410 VDD.t145 461.096
R66 VDD.t281 VDD.t410 461.096
R67 VDD.t267 VDD.t195 461.096
R68 VDD.t272 VDD.t267 461.096
R69 VDD.t38 VDD.t311 461.096
R70 VDD.t42 VDD.t387 461.096
R71 VDD VDD.n196 429.187
R72 VDD.n325 VDD 429.187
R73 VDD VDD.n108 429.187
R74 VDD VDD.n64 429.187
R75 VDD VDD.n442 429.187
R76 VDD VDD.n462 429.187
R77 VDD VDD.n301 427.092
R78 VDD VDD.n119 427.092
R79 VDD VDD.n303 426.699
R80 VDD VDD.n373 426.699
R81 VDD VDD.n192 424.618
R82 VDD VDD.n292 420.935
R83 VDD VDD.n115 420.935
R84 VDD.n208 VDD 418.495
R85 VDD.n442 VDD.t152 386.365
R86 VDD.t107 VDD.n64 386.365
R87 VDD.n196 VDD.t44 386.365
R88 VDD.n303 VDD.t246 386.365
R89 VDD.t293 VDD.n325 386.365
R90 VDD.n373 VDD.t218 386.365
R91 VDD.t117 VDD.n108 386.365
R92 VDD.t351 VDD.t363 380.952
R93 VDD.t192 VDD.t216 380.952
R94 VDD.t220 VDD.n208 378.788
R95 VDD.n292 VDD.t81 378.788
R96 VDD.n115 VDD.t115 378.788
R97 VDD.n208 VDD.t337 322.223
R98 VDD.t394 VDD.n292 322.223
R99 VDD.t438 VDD.n115 322.223
R100 VDD.n192 VDD.t175 320.635
R101 VDD.n301 VDD.t432 320.635
R102 VDD.n119 VDD.t348 320.635
R103 VDD.t16 VDD.t306 303.031
R104 VDD.t11 VDD.t420 303.031
R105 VDD.t254 VDD.t399 303.031
R106 VDD.t425 VDD.t316 303.031
R107 VDD.t24 VDD.t228 303.031
R108 VDD.t296 VDD.t403 303.031
R109 VDD.t248 VDD.t284 303.031
R110 VDD.t208 VDD.t408 303.031
R111 VDD.t189 VDD.t139 303.031
R112 VDD.t428 VDD.t259 303.031
R113 VDD.t184 VDD.t324 303.031
R114 VDD.t366 VDD.t33 303.031
R115 VDD.t181 VDD.t179 303.031
R116 VDD.t235 VDD.t112 303.031
R117 VDD.t122 VDD.t131 303.031
R118 VDD.t358 VDD.t67 303.031
R119 VDD.t278 VDD.t390 303.031
R120 VDD.t19 VDD.t415 303.031
R121 VDD.n252 VDD.t213 242.857
R122 VDD.n254 VDD.t321 242.857
R123 VDD.t363 VDD.n257 242.857
R124 VDD.n261 VDD.t192 242.857
R125 VDD.n447 VDD.t308 193.183
R126 VDD.n448 VDD.t78 193.183
R127 VDD.n457 VDD.t200 193.183
R128 VDD.n458 VDD.t16 193.183
R129 VDD.n428 VDD.t9 193.183
R130 VDD.n434 VDD.t98 193.183
R131 VDD.n435 VDD.t49 193.183
R132 VDD.n441 VDD.t420 193.183
R133 VDD.n38 VDD.t330 193.183
R134 VDD.n40 VDD.t101 193.183
R135 VDD.n43 VDD.t254 193.183
R136 VDD.n46 VDD.t425 193.183
R137 VDD.n209 VDD.t220 193.183
R138 VDD.n286 VDD.t136 193.183
R139 VDD.n289 VDD.t318 193.183
R140 VDD.n294 VDD.t299 193.183
R141 VDD.n299 VDD.t189 193.183
R142 VDD.n242 VDD.t243 193.183
R143 VDD.n243 VDD.t88 193.183
R144 VDD.n249 VDD.t223 193.183
R145 VDD.n250 VDD.t184 193.183
R146 VDD.n219 VDD.t176 193.183
R147 VDD.n221 VDD.t85 193.183
R148 VDD.n224 VDD.t366 193.183
R149 VDD.n227 VDD.t181 193.183
R150 VDD.n5 VDD.t417 193.183
R151 VDD.n7 VDD.t75 193.183
R152 VDD.n10 VDD.t278 193.183
R153 VDD.n13 VDD.t19 193.183
R154 VDD.t228 VDD.n66 191.288
R155 VDD.t91 VDD.n70 191.288
R156 VDD.t288 VDD.n72 191.288
R157 VDD.n74 VDD.t27 191.288
R158 VDD.t403 VDD.n170 191.288
R159 VDD.t284 VDD.n174 191.288
R160 VDD.t328 VDD.n178 191.288
R161 VDD.n180 VDD.t83 191.288
R162 VDD.t408 VDD.n200 191.288
R163 VDD.n201 VDD.t55 191.288
R164 VDD.t326 VDD.n383 191.288
R165 VDD.n384 VDD.t211 191.288
R166 VDD.t81 VDD.n290 191.288
R167 VDD.n364 VDD.t428 191.288
R168 VDD.n363 VDD.t314 191.288
R169 VDD.t40 VDD.n329 191.288
R170 VDD.n331 VDD.t262 191.288
R171 VDD.n406 VDD.t235 191.288
R172 VDD.n405 VDD.t447 191.288
R173 VDD.n404 VDD.t341 191.288
R174 VDD.n403 VDD.t110 191.288
R175 VDD.t115 VDD.n113 191.288
R176 VDD.t131 VDD.n94 191.288
R177 VDD.n95 VDD.t358 191.288
R178 VDD.t286 VDD.n103 191.288
R179 VDD.n104 VDD.t120 191.288
R180 VDD.n207 VDD.t175 142.857
R181 VDD.t432 VDD.n296 142.857
R182 VDD.t348 VDD.n117 142.857
R183 VDD.t22 VDD.n252 138.095
R184 VDD.t302 VDD.n254 138.095
R185 VDD.t29 VDD.n257 138.095
R186 VDD.n261 VDD.t149 138.095
R187 VDD.n156 VDD.t3 118.156
R188 VDD.n351 VDD.t272 118.156
R189 VDD.n66 VDD.t107 111.743
R190 VDD.n70 VDD.t360 111.743
R191 VDD.n72 VDD.t70 111.743
R192 VDD.n74 VDD.t64 111.743
R193 VDD.n170 VDD.t162 111.743
R194 VDD.n174 VDD.t345 111.743
R195 VDD.n178 VDD.t52 111.743
R196 VDD.n180 VDD.t382 111.743
R197 VDD.n200 VDD.t44 111.743
R198 VDD.n201 VDD.t0 111.743
R199 VDD.n383 VDD.t251 111.743
R200 VDD.n384 VDD.t104 111.743
R201 VDD.n290 VDD.t444 111.743
R202 VDD.n364 VDD.t293 111.743
R203 VDD.t57 VDD.n363 111.743
R204 VDD.n329 VDD.t275 111.743
R205 VDD.n331 VDD.t133 111.743
R206 VDD.n406 VDD.t117 111.743
R207 VDD.t35 VDD.n405 111.743
R208 VDD.t6 VDD.n404 111.743
R209 VDD.t377 VDD.n403 111.743
R210 VDD.n113 VDD.t435 111.743
R211 VDD.n94 VDD.t158 111.743
R212 VDD.n95 VDD.t205 111.743
R213 VDD.n103 VDD.t93 111.743
R214 VDD.n104 VDD.t269 111.743
R215 VDD.t337 VDD.n207 111.112
R216 VDD.n296 VDD.t394 111.112
R217 VDD.n117 VDD.t438 111.112
R218 VDD.t430 VDD.n447 109.849
R219 VDD.n448 VDD.t392 109.849
R220 VDD.t73 VDD.n457 109.849
R221 VDD.n458 VDD.t142 109.849
R222 VDD.n428 VDD.t385 109.849
R223 VDD.t397 VDD.n434 109.849
R224 VDD.n435 VDD.t257 109.849
R225 VDD.t152 VDD.n441 109.849
R226 VDD.t96 VDD.n38 109.849
R227 VDD.t47 VDD.n40 109.849
R228 VDD.t125 VDD.n43 109.849
R229 VDD.n46 VDD.t166 109.849
R230 VDD.n209 VDD.t129 109.849
R231 VDD.t380 VDD.n286 109.849
R232 VDD.t349 VDD.n289 109.849
R233 VDD.t60 VDD.n294 109.849
R234 VDD.t246 VDD.n299 109.849
R235 VDD.t343 VDD.n242 109.849
R236 VDD.n243 VDD.t31 109.849
R237 VDD.t333 VDD.n249 109.849
R238 VDD.t218 VDD.n250 109.849
R239 VDD.t369 VDD.n219 109.849
R240 VDD.t226 VDD.n221 109.849
R241 VDD.t335 VDD.n224 109.849
R242 VDD.n227 VDD.t155 109.849
R243 VDD.t62 VDD.n5 109.849
R244 VDD.t203 VDD.n7 109.849
R245 VDD.t433 VDD.n10 109.849
R246 VDD.n13 VDD.t169 109.849
R247 VDD.n260 VDD.t351 97.6195
R248 VDD.n303 VDD.t127 62.1896
R249 VDD.n373 VDD.t187 62.1896
R250 VDD.n192 VDD.t401 61.8817
R251 VDD.n208 VDD.t304 60.9761
R252 VDD.n462 VDD.t14 59.702
R253 VDD.n442 VDD.t423 59.702
R254 VDD.n64 VDD.t232 59.702
R255 VDD.n196 VDD.t405 59.702
R256 VDD.n325 VDD.t412 59.702
R257 VDD.n108 VDD.t237 59.702
R258 VDD.n301 VDD.t441 59.4064
R259 VDD.n119 VDD.t264 59.4064
R260 VDD.n292 VDD.t371 58.5371
R261 VDD.n115 VDD.t240 58.5371
R262 VDD.n49 VDD.t165 30.9379
R263 VDD.n47 VDD.t151 30.9379
R264 VDD.n264 VDD.t154 30.9379
R265 VDD.n162 VDD.t144 30.9379
R266 VDD.n82 VDD.t171 30.9379
R267 VDD.n14 VDD.t141 30.9379
R268 VDD.n15 VDD.t168 30.9379
R269 VDD.n165 VDD.t161 30.3459
R270 VDD.n85 VDD.t157 30.3459
R271 VDD.n263 VDD.t148 29.9642
R272 VDD.n49 VDD.t459 24.5101
R273 VDD.n47 VDD.t463 24.5101
R274 VDD.n269 VDD.t464 24.5101
R275 VDD.n264 VDD.t462 24.5101
R276 VDD.n162 VDD.t454 24.5101
R277 VDD.n82 VDD.t455 24.5101
R278 VDD.n14 VDD.t453 24.5101
R279 VDD.n15 VDD.t457 24.5101
R280 VDD.n166 VDD.t460 24.4392
R281 VDD.n86 VDD.t461 24.4392
R282 VDD.n164 VDD.n163 8.14079
R283 VDD.n84 VDD.n83 8.14079
R284 VDD.n270 VDD.n269 8.0005
R285 VDD.n167 VDD.n166 8.0005
R286 VDD.n87 VDD.n86 8.0005
R287 VDD.n266 VDD.n265 6.99025
R288 VDD.n52 VDD.n46 6.3005
R289 VDD.n55 VDD.n43 6.3005
R290 VDD.n58 VDD.n40 6.3005
R291 VDD.n61 VDD.n38 6.3005
R292 VDD.n207 VDD.n206 6.3005
R293 VDD.n210 VDD.n209 6.3005
R294 VDD.n383 VDD.n382 6.3005
R295 VDD.n203 VDD.n201 6.3005
R296 VDD.n200 VDD.n199 6.3005
R297 VDD.n308 VDD.n296 6.3005
R298 VDD.n317 VDD.n289 6.3005
R299 VDD.n311 VDD.n294 6.3005
R300 VDD.n306 VDD.n299 6.3005
R301 VDD.n316 VDD.n290 6.3005
R302 VDD.n353 VDD.n352 6.3005
R303 VDD.n346 VDD.n332 6.3005
R304 VDD.n350 VDD.n349 6.3005
R305 VDD.n363 VDD.n362 6.3005
R306 VDD.n359 VDD.n329 6.3005
R307 VDD.n356 VDD.n331 6.3005
R308 VDD.n365 VDD.n364 6.3005
R309 VDD.n369 VDD.n286 6.3005
R310 VDD.n283 VDD.n252 6.3005
R311 VDD.n280 VDD.n254 6.3005
R312 VDD.n277 VDD.n257 6.3005
R313 VDD.n274 VDD.n261 6.3005
R314 VDD.n237 VDD.n219 6.3005
R315 VDD.n234 VDD.n221 6.3005
R316 VDD.n231 VDD.n224 6.3005
R317 VDD.n228 VDD.n227 6.3005
R318 VDD.n242 VDD.n241 6.3005
R319 VDD.n244 VDD.n243 6.3005
R320 VDD.n249 VDD.n248 6.3005
R321 VDD.n375 VDD.n250 6.3005
R322 VDD.n385 VDD.n384 6.3005
R323 VDD.n398 VDD.n170 6.3005
R324 VDD.n395 VDD.n174 6.3005
R325 VDD.n392 VDD.n178 6.3005
R326 VDD.n389 VDD.n180 6.3005
R327 VDD.n158 VDD.n157 6.3005
R328 VDD.n151 VDD.n137 6.3005
R329 VDD.n155 VDD.n154 6.3005
R330 VDD.n403 VDD.n402 6.3005
R331 VDD.n404 VDD.n133 6.3005
R332 VDD.n405 VDD.n129 6.3005
R333 VDD.n121 VDD.n117 6.3005
R334 VDD.n125 VDD.n113 6.3005
R335 VDD.n407 VDD.n406 6.3005
R336 VDD.n105 VDD.n104 6.3005
R337 VDD.n103 VDD.n102 6.3005
R338 VDD.n96 VDD.n95 6.3005
R339 VDD.n94 VDD.n93 6.3005
R340 VDD.n414 VDD.n74 6.3005
R341 VDD.n417 VDD.n72 6.3005
R342 VDD.n420 VDD.n70 6.3005
R343 VDD.n423 VDD.n66 6.3005
R344 VDD.n429 VDD.n428 6.3005
R345 VDD.n434 VDD.n433 6.3005
R346 VDD.n436 VDD.n435 6.3005
R347 VDD.n441 VDD.n440 6.3005
R348 VDD.n19 VDD.n13 6.3005
R349 VDD.n22 VDD.n10 6.3005
R350 VDD.n25 VDD.n7 6.3005
R351 VDD.n28 VDD.n5 6.3005
R352 VDD.n447 VDD.n446 6.3005
R353 VDD.n449 VDD.n448 6.3005
R354 VDD.n457 VDD.n456 6.3005
R355 VDD.n459 VDD.n458 6.3005
R356 VDD.n30 VDD.t424 5.85907
R357 VDD.n202 VDD.t305 5.85907
R358 VDD.n461 VDD.t15 5.85907
R359 VDD.n312 VDD.n293 5.85007
R360 VDD.n304 VDD.t247 5.22601
R361 VDD.n410 VDD.n409 5.21771
R362 VDD.n334 VDD.n333 5.213
R363 VDD.n228 VDD.t156 5.213
R364 VDD.n139 VDD.n138 5.213
R365 VDD.n368 VDD.t381 5.18919
R366 VDD VDD.n195 5.16369
R367 VDD.n197 VDD.n194 5.13761
R368 VDD.n439 VDD.t153 5.13287
R369 VDD.n437 VDD.t258 5.13287
R370 VDD.n34 VDD.n33 5.13287
R371 VDD.n432 VDD.t398 5.13287
R372 VDD.n431 VDD.n35 5.13287
R373 VDD.n430 VDD.t386 5.13287
R374 VDD.n427 VDD.n36 5.13287
R375 VDD.n51 VDD.t167 5.13287
R376 VDD.n54 VDD.t126 5.13287
R377 VDD.n57 VDD.t48 5.13287
R378 VDD.n59 VDD.n39 5.13287
R379 VDD.n60 VDD.t97 5.13287
R380 VDD.n62 VDD.n37 5.13287
R381 VDD.n386 VDD.t212 5.13287
R382 VDD.n186 VDD.n185 5.13287
R383 VDD.n381 VDD.t130 5.13287
R384 VDD.n380 VDD.t327 5.13287
R385 VDD.n184 VDD.n183 5.13287
R386 VDD.n187 VDD.t56 5.13287
R387 VDD.n204 VDD.n191 5.13287
R388 VDD.n370 VDD.n285 5.13287
R389 VDD.n319 VDD.n287 5.13287
R390 VDD.n315 VDD.t350 5.13287
R391 VDD.n313 VDD.n291 5.13287
R392 VDD.n310 VDD.t61 5.13287
R393 VDD.n314 VDD.t82 5.13287
R394 VDD.n318 VDD.n288 5.13287
R395 VDD.n324 VDD.n323 5.13287
R396 VDD.n354 VDD.t43 5.13287
R397 VDD.n344 VDD.n343 5.13287
R398 VDD.n345 VDD.t39 5.13287
R399 VDD.n347 VDD.n342 5.13287
R400 VDD.n339 VDD.n335 5.13287
R401 VDD.n355 VDD.t263 5.13287
R402 VDD.n357 VDD.n330 5.13287
R403 VDD.n358 VDD.t41 5.13287
R404 VDD.n360 VDD.n328 5.13287
R405 VDD.n361 VDD.t315 5.13287
R406 VDD.n327 VDD.n326 5.13287
R407 VDD.n284 VDD.n251 5.13287
R408 VDD.n282 VDD.t23 5.13287
R409 VDD.n281 VDD.n253 5.13287
R410 VDD.n279 VDD.t303 5.13287
R411 VDD.n276 VDD.t30 5.13287
R412 VDD.n238 VDD.n218 5.13287
R413 VDD.n236 VDD.t370 5.13287
R414 VDD.n235 VDD.n220 5.13287
R415 VDD.n233 VDD.t227 5.13287
R416 VDD.n230 VDD.t336 5.13287
R417 VDD.n239 VDD.n217 5.13287
R418 VDD.n240 VDD.t344 5.13287
R419 VDD.n216 VDD.n215 5.13287
R420 VDD.n245 VDD.t32 5.13287
R421 VDD.n246 VDD.n214 5.13287
R422 VDD.n247 VDD.t334 5.13287
R423 VDD.n374 VDD.t219 5.13287
R424 VDD.n388 VDD.t84 5.13287
R425 VDD.n390 VDD.n179 5.13287
R426 VDD.n391 VDD.t329 5.13287
R427 VDD.n393 VDD.n177 5.13287
R428 VDD.n396 VDD.n173 5.13287
R429 VDD.n159 VDD.t357 5.13287
R430 VDD.n149 VDD.n148 5.13287
R431 VDD.n150 VDD.t340 5.13287
R432 VDD.n152 VDD.n147 5.13287
R433 VDD.n144 VDD.n140 5.13287
R434 VDD.n401 VDD.t111 5.13287
R435 VDD.n136 VDD.n134 5.13287
R436 VDD.n135 VDD.t342 5.13287
R437 VDD.n132 VDD.n130 5.13287
R438 VDD.n131 VDD.t448 5.13287
R439 VDD.n128 VDD.n127 5.13287
R440 VDD.n124 VDD.t116 5.13287
R441 VDD.n126 VDD.n112 5.13287
R442 VDD.n106 VDD.t121 5.13287
R443 VDD.n100 VDD.n99 5.13287
R444 VDD.n101 VDD.t287 5.13287
R445 VDD.n98 VDD.n75 5.13287
R446 VDD.n79 VDD.n78 5.13287
R447 VDD.n460 VDD.t143 5.13287
R448 VDD.n455 VDD.t74 5.13287
R449 VDD.n451 VDD.n0 5.13287
R450 VDD.n450 VDD.t393 5.13287
R451 VDD.n2 VDD.n1 5.13287
R452 VDD.n445 VDD.t431 5.13287
R453 VDD.n444 VDD.n3 5.13287
R454 VDD.n18 VDD.t170 5.13287
R455 VDD.n21 VDD.t434 5.13287
R456 VDD.n24 VDD.t204 5.13287
R457 VDD.n26 VDD.n6 5.13287
R458 VDD.n27 VDD.t63 5.13287
R459 VDD.n29 VDD.n4 5.13287
R460 VDD.n413 VDD.t28 5.12655
R461 VDD.n415 VDD.n73 5.12655
R462 VDD.n416 VDD.t289 5.12655
R463 VDD.n418 VDD.n71 5.12655
R464 VDD.n419 VDD.t92 5.12655
R465 VDD.n421 VDD.n69 5.12655
R466 VDD.n424 VDD.n65 5.12655
R467 VDD VDD.t128 5.11529
R468 VDD.n193 VDD.t402 5.09407
R469 VDD.n302 VDD.n300 5.09407
R470 VDD.n182 VDD.n181 5.09407
R471 VDD.n372 VDD.t188 5.09407
R472 VDD.n120 VDD.n118 5.09407
R473 VDD.n123 VDD.n114 5.09407
R474 VDD.n411 VDD.n107 5.09407
R475 VDD.n425 VDD.n63 5.09407
R476 VDD.n400 VDD.n399 5.08521
R477 VDD.n378 VDD.n377 4.99361
R478 VDD.n273 VDD.t150 4.8755
R479 VDD.n169 VDD.n160 4.8755
R480 VDD.n89 VDD.n80 4.8755
R481 VDD.n266 VDD.n262 4.51272
R482 VDD.n269 VDD.n268 4.5005
R483 VDD VDD.n14 4.35564
R484 VDD.n205 VDD.t338 4.12326
R485 VDD.n309 VDD.n295 4.12326
R486 VDD.n122 VDD.n116 4.12326
R487 VDD VDD.n49 4.09565
R488 VDD.n48 VDD.n47 4.08504
R489 VDD VDD.n15 4.00785
R490 VDD.n267 VDD.n263 3.6022
R491 VDD.n17 VDD 3.06902
R492 VDD.n50 VDD.n48 2.93012
R493 VDD.n17 VDD.n16 2.86671
R494 VDD.n438 VDD.n32 2.85787
R495 VDD.n53 VDD.n45 2.85787
R496 VDD.n56 VDD.n42 2.85787
R497 VDD.n190 VDD.n189 2.85787
R498 VDD.n307 VDD.n298 2.85787
R499 VDD.n348 VDD.n341 2.85787
R500 VDD.n338 VDD.n337 2.85787
R501 VDD.n322 VDD.n321 2.85787
R502 VDD.n278 VDD.n256 2.85787
R503 VDD.n275 VDD.n259 2.85787
R504 VDD.n232 VDD.n223 2.85787
R505 VDD.n229 VDD.n226 2.85787
R506 VDD.n213 VDD.n212 2.85787
R507 VDD.n394 VDD.n176 2.85787
R508 VDD.n397 VDD.n172 2.85787
R509 VDD.n153 VDD.n146 2.85787
R510 VDD.n143 VDD.n142 2.85787
R511 VDD.n111 VDD.n110 2.85787
R512 VDD.n97 VDD.n77 2.85787
R513 VDD.n92 VDD.n91 2.85787
R514 VDD.n454 VDD.n453 2.85787
R515 VDD.n20 VDD.n12 2.85787
R516 VDD.n23 VDD.n9 2.85787
R517 VDD.n422 VDD.n68 2.85155
R518 VDD.n50 VDD 2.83528
R519 VDD.n18 VDD.n17 2.28244
R520 VDD.n32 VDD.t12 2.2755
R521 VDD.n32 VDD.n31 2.2755
R522 VDD.n45 VDD.t317 2.2755
R523 VDD.n45 VDD.n44 2.2755
R524 VDD.n42 VDD.t400 2.2755
R525 VDD.n42 VDD.n41 2.2755
R526 VDD.n189 VDD.t409 2.2755
R527 VDD.n189 VDD.n188 2.2755
R528 VDD.n298 VDD.t140 2.2755
R529 VDD.n298 VDD.n297 2.2755
R530 VDD.n341 VDD.t268 2.2755
R531 VDD.n341 VDD.n340 2.2755
R532 VDD.n337 VDD.t411 2.2755
R533 VDD.n337 VDD.n336 2.2755
R534 VDD.n321 VDD.t429 2.2755
R535 VDD.n321 VDD.n320 2.2755
R536 VDD.n256 VDD.t352 2.2755
R537 VDD.n256 VDD.n255 2.2755
R538 VDD.n259 VDD.t217 2.2755
R539 VDD.n259 VDD.n258 2.2755
R540 VDD.n223 VDD.t34 2.2755
R541 VDD.n223 VDD.n222 2.2755
R542 VDD.n226 VDD.t180 2.2755
R543 VDD.n226 VDD.n225 2.2755
R544 VDD.n212 VDD.t325 2.2755
R545 VDD.n212 VDD.n211 2.2755
R546 VDD.n176 VDD.t285 2.2755
R547 VDD.n176 VDD.n175 2.2755
R548 VDD.n172 VDD.t404 2.2755
R549 VDD.n172 VDD.n171 2.2755
R550 VDD.n146 VDD.t199 2.2755
R551 VDD.n146 VDD.n145 2.2755
R552 VDD.n142 VDD.t231 2.2755
R553 VDD.n142 VDD.n141 2.2755
R554 VDD.n110 VDD.t236 2.2755
R555 VDD.n110 VDD.n109 2.2755
R556 VDD.n77 VDD.t359 2.2755
R557 VDD.n77 VDD.n76 2.2755
R558 VDD.n91 VDD.t132 2.2755
R559 VDD.n91 VDD.n90 2.2755
R560 VDD.n68 VDD.t229 2.2755
R561 VDD.n68 VDD.n67 2.2755
R562 VDD.n453 VDD.t307 2.2755
R563 VDD.n453 VDD.n452 2.2755
R564 VDD.n12 VDD.t416 2.2755
R565 VDD.n12 VDD.n11 2.2755
R566 VDD.n9 VDD.t391 2.2755
R567 VDD.n9 VDD.n8 2.2755
R568 VDD.n51 VDD.n50 2.27489
R569 VDD.n163 VDD.n162 2.11346
R570 VDD.n83 VDD.n82 2.11346
R571 VDD.n265 VDD.n264 2.11318
R572 VDD.n165 VDD.n164 1.81921
R573 VDD.n85 VDD.n84 1.81921
R574 VDD.n426 VDD.n425 1.78842
R575 VDD.n197 VDD 1.77385
R576 VDD VDD.n324 1.77343
R577 VDD.n268 VDD.n266 1.54696
R578 VDD.n239 VDD.n238 1.16167
R579 VDD.n355 VDD.n354 1.16051
R580 VDD.n401 VDD.n400 1.12915
R581 VDD.n388 VDD.n387 1.0737
R582 VDD.n426 VDD.n62 1.02928
R583 VDD.n443 VDD.n29 1.02928
R584 VDD.n371 VDD.n284 1.01882
R585 VDD.n412 VDD.n106 1.01824
R586 VDD.n269 VDD.n263 0.798596
R587 VDD.n378 VDD 0.59265
R588 VDD VDD.n366 0.468962
R589 VDD.n408 VDD 0.468962
R590 VDD.n166 VDD.n165 0.423118
R591 VDD.n86 VDD.n85 0.423118
R592 VDD.n121 VDD.n120 0.389068
R593 VDD.n379 VDD.n378 0.346452
R594 VDD.n274 VDD.n273 0.337997
R595 VDD.n93 VDD.n89 0.337997
R596 VDD.n273 VDD.n272 0.328132
R597 VDD.n169 VDD.n168 0.328132
R598 VDD.n89 VDD.n88 0.328132
R599 VDD VDD.n376 0.316077
R600 VDD VDD.n126 0.274338
R601 VDD VDD.n122 0.269908
R602 VDD.n399 VDD.n169 0.257868
R603 VDD.n57 VDD.n56 0.233919
R604 VDD.n54 VDD.n53 0.233919
R605 VDD.n339 VDD.n338 0.233919
R606 VDD.n348 VDD.n347 0.233919
R607 VDD.n279 VDD.n278 0.233919
R608 VDD.n276 VDD.n275 0.233919
R609 VDD.n233 VDD.n232 0.233919
R610 VDD.n230 VDD.n229 0.233919
R611 VDD.n397 VDD.n396 0.233919
R612 VDD.n394 VDD.n393 0.233919
R613 VDD.n144 VDD.n143 0.233919
R614 VDD.n153 VDD.n152 0.233919
R615 VDD.n92 VDD.n79 0.233919
R616 VDD.n98 VDD.n97 0.233919
R617 VDD.n24 VDD.n23 0.233919
R618 VDD.n21 VDD.n20 0.233919
R619 VDD.n367 VDD 0.216814
R620 VDD.n379 VDD 0.216814
R621 VDD.n124 VDD.n123 0.170499
R622 VDD VDD.n424 0.166121
R623 VDD.n387 VDD.n386 0.14292
R624 VDD.n60 VDD.n59 0.141016
R625 VDD.n345 VDD.n344 0.141016
R626 VDD.n361 VDD.n360 0.141016
R627 VDD.n358 VDD.n357 0.141016
R628 VDD.n282 VDD.n281 0.141016
R629 VDD.n236 VDD.n235 0.141016
R630 VDD.n240 VDD.n216 0.141016
R631 VDD.n246 VDD.n245 0.141016
R632 VDD.n391 VDD.n390 0.141016
R633 VDD.n150 VDD.n149 0.141016
R634 VDD.n132 VDD.n131 0.141016
R635 VDD.n136 VDD.n135 0.141016
R636 VDD.n101 VDD.n100 0.141016
R637 VDD.n27 VDD.n26 0.141016
R638 VDD VDD.n410 0.140259
R639 VDD.n387 VDD.n182 0.139745
R640 VDD.n305 VDD.n302 0.137219
R641 VDD.n198 VDD.n193 0.13637
R642 VDD.n419 VDD.n418 0.125672
R643 VDD.n416 VDD.n415 0.125672
R644 VDD.n327 VDD 0.123016
R645 VDD.n128 VDD 0.123016
R646 VDD.n247 VDD 0.122435
R647 VDD.n413 VDD.n412 0.117172
R648 VDD VDD.n213 0.111984
R649 VDD VDD.n322 0.111403
R650 VDD VDD.n111 0.111403
R651 VDD VDD.n421 0.109638
R652 VDD.n122 VDD 0.109408
R653 VDD.n163 VDD 0.107393
R654 VDD.n83 VDD 0.107393
R655 VDD.n62 VDD.n61 0.107339
R656 VDD.n59 VDD.n58 0.107339
R657 VDD.n346 VDD.n345 0.107339
R658 VDD.n354 VDD.n353 0.107339
R659 VDD.n362 VDD.n361 0.107339
R660 VDD.n359 VDD.n358 0.107339
R661 VDD.n356 VDD.n355 0.107339
R662 VDD.n284 VDD.n283 0.107339
R663 VDD.n281 VDD.n280 0.107339
R664 VDD.n238 VDD.n237 0.107339
R665 VDD.n235 VDD.n234 0.107339
R666 VDD.n241 VDD.n239 0.107339
R667 VDD.n244 VDD.n216 0.107339
R668 VDD.n248 VDD.n246 0.107339
R669 VDD.n386 VDD.n385 0.107339
R670 VDD.n392 VDD.n391 0.107339
R671 VDD.n389 VDD.n388 0.107339
R672 VDD.n151 VDD.n150 0.107339
R673 VDD.n159 VDD.n158 0.107339
R674 VDD.n131 VDD.n129 0.107339
R675 VDD.n135 VDD.n133 0.107339
R676 VDD.n402 VDD.n401 0.107339
R677 VDD.n125 VDD.n124 0.107339
R678 VDD.n102 VDD.n101 0.107339
R679 VDD.n106 VDD.n105 0.107339
R680 VDD.n29 VDD.n28 0.107339
R681 VDD.n26 VDD.n25 0.107339
R682 VDD.n265 VDD 0.106795
R683 VDD.n338 VDD 0.106758
R684 VDD VDD.n348 0.106758
R685 VDD VDD.n397 0.106758
R686 VDD VDD.n394 0.106758
R687 VDD.n143 VDD 0.106758
R688 VDD VDD.n153 0.106758
R689 VDD VDD.n92 0.106758
R690 VDD.n97 VDD 0.106758
R691 VDD.n56 VDD 0.106177
R692 VDD.n53 VDD 0.106177
R693 VDD.n278 VDD 0.106177
R694 VDD.n275 VDD 0.106177
R695 VDD.n232 VDD 0.106177
R696 VDD.n229 VDD 0.106177
R697 VDD.n23 VDD 0.106177
R698 VDD.n20 VDD 0.106177
R699 VDD.n412 VDD.n411 0.104
R700 VDD.n422 VDD 0.0992931
R701 VDD.n420 VDD.n419 0.0956724
R702 VDD.n417 VDD.n416 0.0956724
R703 VDD.n414 VDD.n413 0.0956724
R704 VDD VDD.n422 0.0951552
R705 VDD.n374 VDD 0.0847644
R706 VDD.n55 VDD.n54 0.080629
R707 VDD.n52 VDD.n51 0.080629
R708 VDD.n349 VDD.n339 0.080629
R709 VDD.n277 VDD.n276 0.080629
R710 VDD.n231 VDD.n230 0.080629
R711 VDD.n399 VDD.n398 0.080629
R712 VDD.n396 VDD.n395 0.080629
R713 VDD.n154 VDD.n144 0.080629
R714 VDD.n96 VDD.n79 0.080629
R715 VDD.n22 VDD.n21 0.080629
R716 VDD.n19 VDD.n18 0.080629
R717 VDD VDD.n60 0.0794677
R718 VDD VDD.n57 0.0794677
R719 VDD VDD.n282 0.0794677
R720 VDD VDD.n279 0.0794677
R721 VDD VDD.n236 0.0794677
R722 VDD VDD.n233 0.0794677
R723 VDD VDD.n240 0.0794677
R724 VDD.n245 VDD 0.0794677
R725 VDD VDD.n247 0.0794677
R726 VDD VDD.n27 0.0794677
R727 VDD VDD.n24 0.0794677
R728 VDD.n347 VDD 0.0788871
R729 VDD.n344 VDD 0.0788871
R730 VDD VDD.n327 0.0788871
R731 VDD.n360 VDD 0.0788871
R732 VDD.n357 VDD 0.0788871
R733 VDD.n393 VDD 0.0788871
R734 VDD.n390 VDD 0.0788871
R735 VDD.n152 VDD 0.0788871
R736 VDD.n149 VDD 0.0788871
R737 VDD VDD.n128 0.0788871
R738 VDD VDD.n132 0.0788871
R739 VDD VDD.n136 0.0788871
R740 VDD VDD.n98 0.0788871
R741 VDD.n100 VDD 0.0788871
R742 VDD.n126 VDD 0.0754032
R743 VDD.n161 VDD 0.0733571
R744 VDD.n81 VDD 0.0733571
R745 VDD.n424 VDD.n423 0.0718793
R746 VDD.n193 VDD 0.0709717
R747 VDD.n421 VDD 0.0703276
R748 VDD.n418 VDD 0.0703276
R749 VDD.n415 VDD 0.0703276
R750 VDD.n302 VDD 0.0701226
R751 VDD VDD.n182 0.0701226
R752 VDD.n120 VDD 0.0701226
R753 VDD.n123 VDD 0.0701226
R754 VDD.n271 VDD 0.0690714
R755 VDD.n376 VDD.n213 0.0616715
R756 VDD.n371 VDD.n370 0.0601785
R757 VDD.n366 VDD.n324 0.0556613
R758 VDD.n304 VDD 0.0531999
R759 VDD.n372 VDD.n371 0.0531705
R760 VDD.n370 VDD.n369 0.0489211
R761 VDD.n272 VDD.n271 0.0471071
R762 VDD.n168 VDD.n161 0.0471071
R763 VDD.n88 VDD.n81 0.0471071
R764 VDD.n366 VDD.n322 0.0417258
R765 VDD.n408 VDD.n111 0.0417258
R766 VDD.n410 VDD.n408 0.0417109
R767 VDD.n411 VDD 0.0415
R768 VDD.n425 VDD 0.0415
R769 VDD.n167 VDD.n164 0.0387491
R770 VDD.n87 VDD.n84 0.0387491
R771 VDD.n439 VDD.n30 0.037789
R772 VDD.n461 VDD.n460 0.0376465
R773 VDD.n375 VDD.n374 0.0368158
R774 VDD VDD.n190 0.0366978
R775 VDD.n307 VDD 0.0365
R776 VDD.n270 VDD.n262 0.0358571
R777 VDD.n168 VDD.n167 0.0358571
R778 VDD.n88 VDD.n87 0.0358571
R779 VDD.n205 VDD.n204 0.0349176
R780 VDD.n310 VDD.n309 0.0349176
R781 VDD.n272 VDD.n270 0.03425
R782 VDD VDD.n187 0.033533
R783 VDD.n313 VDD 0.0333352
R784 VDD VDD.n368 0.033241
R785 VDD.n400 VDD.n159 0.0318548
R786 VDD.n187 VDD.n186 0.0307637
R787 VDD.n314 VDD.n313 0.0307637
R788 VDD.n431 VDD.n430 0.0283517
R789 VDD.n432 VDD.n34 0.0283517
R790 VDD.n445 VDD.n2 0.0282452
R791 VDD.n451 VDD.n450 0.0282452
R792 VDD VDD.n310 0.0274011
R793 VDD.n204 VDD 0.0272033
R794 VDD.n427 VDD.n426 0.0267404
R795 VDD.n444 VDD.n443 0.0266401
R796 VDD.n368 VDD.n367 0.0252441
R797 VDD VDD.n437 0.0246688
R798 VDD.n455 VDD 0.0245764
R799 VDD.n198 VDD.n197 0.0230424
R800 VDD.n438 VDD 0.0225972
R801 VDD VDD.n454 0.0225127
R802 VDD VDD.n372 0.0217216
R803 VDD.n429 VDD.n427 0.0216765
R804 VDD.n433 VDD.n431 0.0216765
R805 VDD.n436 VDD.n34 0.0216765
R806 VDD.n446 VDD.n444 0.0215955
R807 VDD.n449 VDD.n2 0.0215955
R808 VDD.n456 VDD.n451 0.0215955
R809 VDD VDD.n438 0.0214463
R810 VDD.n454 VDD 0.0213662
R811 VDD.n366 VDD.n365 0.0201154
R812 VDD.n408 VDD.n407 0.0201154
R813 VDD.n210 VDD.n184 0.0192912
R814 VDD.n382 VDD.n381 0.0192912
R815 VDD.n318 VDD.n317 0.0192912
R816 VDD.n316 VDD.n315 0.0192912
R817 VDD.n186 VDD.n184 0.0181044
R818 VDD.n381 VDD.n380 0.0181044
R819 VDD.n319 VDD.n318 0.0181044
R820 VDD.n315 VDD.n314 0.0181044
R821 VDD.n440 VDD.n439 0.0163824
R822 VDD.n460 VDD.n459 0.0163217
R823 VDD.n430 VDD 0.0161522
R824 VDD VDD.n432 0.0161522
R825 VDD.n437 VDD 0.0161522
R826 VDD VDD.n445 0.0160924
R827 VDD.n450 VDD 0.0160924
R828 VDD VDD.n455 0.0160924
R829 VDD.n308 VDD.n307 0.0157308
R830 VDD.n206 VDD.n190 0.015533
R831 VDD.n199 VDD.n198 0.0149396
R832 VDD.n306 VDD.n305 0.0147418
R833 VDD.n16 VDD 0.0113333
R834 VDD.n376 VDD 0.00944737
R835 VDD.n271 VDD 0.00907143
R836 VDD.n305 VDD.n304 0.00906907
R837 VDD VDD.n205 0.00781868
R838 VDD.n367 VDD.n319 0.00762088
R839 VDD.n309 VDD 0.00762088
R840 VDD.n380 VDD.n379 0.00742308
R841 VDD VDD.n121 0.00579412
R842 VDD VDD.n125 0.00572581
R843 VDD.n48 VDD 0.00564286
R844 VDD.n443 VDD 0.00508599
R845 VDD.n161 VDD 0.00478571
R846 VDD.n81 VDD 0.00478571
R847 VDD.n16 VDD 0.00466667
R848 VDD.n267 VDD.n262 0.00371429
R849 VDD.n312 VDD.n311 0.00366484
R850 VDD.n203 VDD.n202 0.00346703
R851 VDD VDD.n316 0.00228022
R852 VDD VDD.n346 0.00224194
R853 VDD.n353 VDD 0.00224194
R854 VDD.n362 VDD 0.00224194
R855 VDD VDD.n359 0.00224194
R856 VDD VDD.n356 0.00224194
R857 VDD.n385 VDD 0.00224194
R858 VDD VDD.n392 0.00224194
R859 VDD VDD.n389 0.00224194
R860 VDD VDD.n151 0.00224194
R861 VDD.n158 VDD 0.00224194
R862 VDD.n129 VDD 0.00224194
R863 VDD.n133 VDD 0.00224194
R864 VDD.n402 VDD 0.00224194
R865 VDD.n102 VDD 0.00224194
R866 VDD.n105 VDD 0.00224194
R867 VDD.n268 VDD.n267 0.00210714
R868 VDD VDD.n210 0.00208242
R869 VDD VDD.n420 0.00205172
R870 VDD VDD.n417 0.00205172
R871 VDD VDD.n414 0.00205172
R872 VDD.n206 VDD 0.00188462
R873 VDD VDD.n308 0.00188462
R874 VDD.n61 VDD 0.00166129
R875 VDD.n58 VDD 0.00166129
R876 VDD VDD.n55 0.00166129
R877 VDD VDD.n52 0.00166129
R878 VDD.n283 VDD 0.00166129
R879 VDD.n280 VDD 0.00166129
R880 VDD VDD.n277 0.00166129
R881 VDD VDD.n274 0.00166129
R882 VDD.n237 VDD 0.00166129
R883 VDD.n234 VDD 0.00166129
R884 VDD VDD.n231 0.00166129
R885 VDD VDD.n228 0.00166129
R886 VDD.n241 VDD 0.00166129
R887 VDD VDD.n244 0.00166129
R888 VDD.n248 VDD 0.00166129
R889 VDD.n28 VDD 0.00166129
R890 VDD.n25 VDD 0.00166129
R891 VDD VDD.n22 0.00166129
R892 VDD VDD.n19 0.00166129
R893 VDD VDD.n203 0.00109341
R894 VDD.n382 VDD 0.00109341
R895 VDD VDD.n334 0.00108064
R896 VDD.n349 VDD 0.00108064
R897 VDD.n398 VDD 0.00108064
R898 VDD.n395 VDD 0.00108064
R899 VDD VDD.n139 0.00108064
R900 VDD.n154 VDD 0.00108064
R901 VDD.n93 VDD 0.00108064
R902 VDD VDD.n96 0.00108064
R903 VDD.n365 VDD 0.00107692
R904 VDD.n407 VDD 0.00107692
R905 VDD.n369 VDD 0.00102632
R906 VDD VDD.n375 0.00102632
R907 VDD.n423 VDD 0.00101724
R908 VDD.n202 VDD 0.000895604
R909 VDD.n317 VDD 0.000895604
R910 VDD VDD.n312 0.000895604
R911 VDD.n311 VDD 0.000895604
R912 VDD VDD.n306 0.000895604
R913 VDD VDD.n429 0.000730179
R914 VDD.n433 VDD 0.000730179
R915 VDD VDD.n436 0.000730179
R916 VDD.n440 VDD 0.000730179
R917 VDD VDD.n30 0.000730179
R918 VDD.n446 VDD 0.000729299
R919 VDD VDD.n449 0.000729299
R920 VDD.n456 VDD 0.000729299
R921 VDD.n459 VDD 0.000729299
R922 VDD VDD.n461 0.000729299
R923 VDD.n199 VDD 0.000697802
R924 RST.n2 RST.t4 37.2595
R925 RST.n49 RST.t10 37.1988
R926 RST.n34 RST.t11 37.1988
R927 RST.n42 RST.t0 36.935
R928 RST.n15 RST.t1 36.935
R929 RST.n24 RST.t14 36.935
R930 RST.n19 RST.t3 36.935
R931 RST.n8 RST.t7 36.935
R932 RST.n42 RST.t13 18.1962
R933 RST.n15 RST.t15 18.1962
R934 RST.n24 RST.t12 18.1962
R935 RST.n19 RST.t2 18.1962
R936 RST.n8 RST.t6 18.1962
R937 RST.n49 RST.t8 17.6613
R938 RST.n34 RST.t9 17.6613
R939 RST.n2 RST.t5 17.5939
R940 RST.n46 RST.n39 7.32578
R941 RST.n47 RST.n12 7.18787
R942 RST.n12 RST.n5 4.99277
R943 RST.n32 RST.n18 4.86625
R944 RST RST.n56 4.54717
R945 RST.n45 RST.n44 4.5005
R946 RST.n18 RST.n17 4.5005
R947 RST.n11 RST.n10 4.5005
R948 RST.n32 RST.n31 4.46212
R949 RST.n12 RST.n11 4.4249
R950 RST.n31 RST.n20 3.94094
R951 RST.n46 RST.n45 3.78663
R952 RST.n55 RST.n54 3.31947
R953 RST.n54 RST.n53 2.8446
R954 RST.n39 RST.n38 2.8446
R955 RST.n43 RST.n41 2.25022
R956 RST.n16 RST.n14 2.25022
R957 RST.n5 RST.n4 2.24196
R958 RST.n53 RST.n52 2.24157
R959 RST.n38 RST.n37 2.24157
R960 RST.n20 RST.n19 2.15477
R961 RST.n43 RST.n42 2.12393
R962 RST.n16 RST.n15 2.12393
R963 RST.n25 RST.n24 2.12188
R964 RST.n9 RST.n8 2.12075
R965 RST.n31 RST.n30 1.78745
R966 RST.n54 RST.n47 1.66471
R967 RST.n39 RST.n32 1.57395
R968 RST.n27 RST.n26 1.5005
R969 RST.n29 RST.n28 1.5005
R970 RST.n7 RST.n6 1.49653
R971 RST.n3 RST.n2 1.42098
R972 RST.n50 RST.n49 1.41601
R973 RST.n35 RST.n34 1.41601
R974 RST.n47 RST.n46 1.12471
R975 RST.n56 RST.n55 0.90484
R976 RST.n7 RST 0.0658428
R977 RST.n40 RST 0.0584663
R978 RST.n13 RST 0.0584663
R979 RST.n20 RST 0.0476942
R980 RST.n1 RST 0.0410354
R981 RST.n51 RST 0.0394837
R982 RST.n36 RST 0.0394837
R983 RST.n52 RST.n51 0.0377414
R984 RST.n37 RST.n36 0.0377414
R985 RST.n26 RST.n23 0.0361897
R986 RST.n4 RST.n1 0.0361897
R987 RST.n30 RST.n29 0.0358571
R988 RST.n23 RST 0.031725
R989 RST.n45 RST 0.0293
R990 RST.n18 RST 0.0293
R991 RST.n11 RST 0.0293
R992 RST.n5 RST.n0 0.0238218
R993 RST.n53 RST.n48 0.0230258
R994 RST.n38 RST.n33 0.0230258
R995 RST.n28 RST.n21 0.0219286
R996 RST.n44 RST.n40 0.0196058
R997 RST.n17 RST.n13 0.0196058
R998 RST RST.n55 0.0145998
R999 RST.n10 RST.n7 0.0131921
R1000 RST.n26 RST.n25 0.0129138
R1001 RST.n27 RST.n22 0.0052523
R1002 RST.n10 RST.n9 0.00515517
R1003 RST.n4 RST.n3 0.00515517
R1004 RST.n28 RST.n27 0.00371429
R1005 RST.n52 RST.n50 0.00360345
R1006 RST.n37 RST.n35 0.00360345
R1007 RST.n44 RST.n43 0.00255119
R1008 RST.n17 RST.n16 0.00255119
R1009 RST.n41 RST 0.0017
R1010 RST.n14 RST 0.0017
R1011 RST.n6 RST 0.0017
R1012 VSS.n100 VSS.n99 71260
R1013 VSS.n101 VSS.n100 39263.5
R1014 VSS.n260 VSS.n40 19564.1
R1015 VSS.n97 VSS.n95 18801.2
R1016 VSS.n188 VSS.t275 14048.5
R1017 VSS.n85 VSS.t272 7280.79
R1018 VSS.n85 VSS.n84 5639.46
R1019 VSS.t265 VSS.n140 5265.51
R1020 VSS.n132 VSS.n131 5147.52
R1021 VSS.n188 VSS.n164 4818.58
R1022 VSS.n84 VSS.n83 4659.38
R1023 VSS.n202 VSS.n201 4287.32
R1024 VSS.n130 VSS.t284 4107.43
R1025 VSS.n234 VSS.n41 3956.92
R1026 VSS.n94 VSS.n54 3893.61
R1027 VSS.n290 VSS.n288 3893.61
R1028 VSS.n134 VSS.n133 3355.98
R1029 VSS.n304 VSS.n281 3063.89
R1030 VSS.n133 VSS.n132 3017.86
R1031 VSS.t278 VSS.t145 2781.65
R1032 VSS.t246 VSS.t224 2781.65
R1033 VSS.n281 VSS.t213 2426.54
R1034 VSS.n281 VSS.t101 2421.57
R1035 VSS.t132 VSS.t0 2307.56
R1036 VSS.t37 VSS.t150 2307.56
R1037 VSS.t197 VSS.t66 2307.56
R1038 VSS.t254 VSS.t182 2307.56
R1039 VSS.t155 VSS.t38 2307.56
R1040 VSS.t195 VSS.t163 2307.56
R1041 VSS.t53 VSS.t270 2307.56
R1042 VSS.t126 VSS.t243 2307.56
R1043 VSS.t191 VSS.t51 2307.56
R1044 VSS.t238 VSS.t65 2307.56
R1045 VSS.t250 VSS.t33 2307.56
R1046 VSS.t15 VSS.t219 2307.56
R1047 VSS.t58 VSS.t48 2307.56
R1048 VSS.t177 VSS.t44 2307.56
R1049 VSS.t75 VSS.t85 2307.56
R1050 VSS.t73 VSS.t22 2307.56
R1051 VSS.t3 VSS.t287 2307.56
R1052 VSS.t264 VSS.t273 2159.54
R1053 VSS.n99 VSS.n98 1925.44
R1054 VSS.n97 VSS.n96 1922.83
R1055 VSS.n288 VSS.t208 1686.81
R1056 VSS.n54 VSS.t56 1684.74
R1057 VSS.n288 VSS.t108 1682.82
R1058 VSS.n54 VSS.t111 1680.76
R1059 VSS.t128 VSS.t209 1611.04
R1060 VSS.t159 VSS.t178 1611.04
R1061 VSS.t179 VSS.t216 1611.04
R1062 VSS.t227 VSS.t205 1611.04
R1063 VSS.t185 VSS.t210 1609.07
R1064 VSS.t234 VSS.t198 1609.07
R1065 VSS.t123 VSS.t174 1609.07
R1066 VSS.t240 VSS.t26 1609.07
R1067 VSS.n131 VSS.t156 1601.22
R1068 VSS.n84 VSS.t281 1601.22
R1069 VSS.n95 VSS.n94 1565.03
R1070 VSS.n290 VSS.n289 1565.03
R1071 VSS.t11 VSS.n112 1544.05
R1072 VSS.n234 VSS.t96 1301.85
R1073 VSS.t133 VSS.n234 1298.77
R1074 VSS.t57 VSS.t222 1243.37
R1075 VSS.t202 VSS.t120 1243.37
R1076 VSS.t196 VSS.t13 1243.37
R1077 VSS.t134 VSS.t17 1243.37
R1078 VSS.t28 VSS.n305 1199.47
R1079 VSS.t94 VSS.n203 1199.47
R1080 VSS.n186 VSS.t69 1199.47
R1081 VSS.n112 VSS.t119 1178.74
R1082 VSS.t27 VSS.n85 1153.78
R1083 VSS.n202 VSS.t190 1153.78
R1084 VSS.n164 VSS.t7 1153.78
R1085 VSS.n304 VSS.t72 1153.78
R1086 VSS.n218 VSS.n217 1041.81
R1087 VSS.n131 VSS.n130 1034.55
R1088 VSS.n213 VSS.n212 1025.15
R1089 VSS.n201 VSS.t104 943.548
R1090 VSS.t262 VSS.t132 913.885
R1091 VSS.t260 VSS.t155 913.885
R1092 VSS.t9 VSS.t191 913.885
R1093 VSS.t267 VSS.t8 913.885
R1094 VSS.t142 VSS.t15 913.885
R1095 VSS.t144 VSS.t73 913.885
R1096 VSS.t245 VSS.t166 855.264
R1097 VSS.t10 VSS.t264 855.264
R1098 VSS.t64 VSS.t62 784.35
R1099 VSS.t78 VSS.t199 784.35
R1100 VSS.n134 VSS.t11 782.221
R1101 VSS.n124 VSS.t217 776.83
R1102 VSS.n77 VSS.t175 776.83
R1103 VSS.n219 VSS.n218 763.912
R1104 VSS.n212 VSS.t42 754.639
R1105 VSS.n142 VSS.t265 699.654
R1106 VSS.n217 VSS.t106 668.119
R1107 VSS.n200 VSS.t269 650.643
R1108 VSS.n261 VSS.t83 641.721
R1109 VSS.t209 VSS.t141 638.038
R1110 VSS.t172 VSS.t47 638.038
R1111 VSS.t216 VSS.t143 638.038
R1112 VSS.t167 VSS.t6 638.038
R1113 VSS.t261 VSS.t185 637.255
R1114 VSS.t173 VSS.t149 637.255
R1115 VSS.t174 VSS.t263 637.255
R1116 VSS.t168 VSS.t162 637.255
R1117 VSS.n124 VSS.t278 554.879
R1118 VSS.n77 VSS.t246 554.879
R1119 VSS.n98 VSS.n97 548.634
R1120 VSS.n318 VSS.t262 548.331
R1121 VSS.n317 VSS.t37 548.331
R1122 VSS.n316 VSS.t197 548.331
R1123 VSS.n315 VSS.t131 548.331
R1124 VSS.n92 VSS.t260 548.331
R1125 VSS.n91 VSS.t195 548.331
R1126 VSS.n90 VSS.t25 548.331
R1127 VSS.n86 VSS.t27 548.331
R1128 VSS.t190 VSS.n154 548.331
R1129 VSS.n143 VSS.t53 548.331
R1130 VSS.n144 VSS.t126 548.331
R1131 VSS.n145 VSS.t9 548.331
R1132 VSS.t7 VSS.n163 548.331
R1133 VSS.t65 VSS.n162 548.331
R1134 VSS.t33 VSS.n161 548.331
R1135 VSS.n204 VSS.t267 548.331
R1136 VSS.n185 VSS.t142 548.331
R1137 VSS.n184 VSS.t58 548.331
R1138 VSS.n183 VSS.t177 548.331
R1139 VSS.n182 VSS.t16 548.331
R1140 VSS.n294 VSS.t144 548.331
R1141 VSS.t287 VSS.n298 548.331
R1142 VSS.n299 VSS.t206 548.331
R1143 VSS.t72 VSS.n303 548.331
R1144 VSS.n69 VSS.t55 546.41
R1145 VSS.n116 VSS.t74 546.41
R1146 VSS.t284 VSS.n23 522.021
R1147 VSS.t275 VSS.n187 508.839
R1148 VSS.t200 VSS.n188 502.839
R1149 VSS.t170 VSS.t21 492.425
R1150 VSS.t120 VSS.t237 492.425
R1151 VSS.t169 VSS.t215 492.425
R1152 VSS.t80 VSS.t134 492.425
R1153 VSS.n217 VSS.t10 400.906
R1154 VSS.t141 VSS.n2 382.822
R1155 VSS.n4 VSS.t172 382.822
R1156 VSS.t178 VSS.n6 382.822
R1157 VSS.t208 VSS.n8 382.822
R1158 VSS.t143 VSS.n11 382.822
R1159 VSS.n13 VSS.t167 382.822
R1160 VSS.t205 VSS.n15 382.822
R1161 VSS.t213 VSS.n17 382.822
R1162 VSS.n280 VSS.t261 382.353
R1163 VSS.n279 VSS.t173 382.353
R1164 VSS.t198 VSS.n28 382.353
R1165 VSS.t56 VSS.n30 382.353
R1166 VSS.t263 VSS.n33 382.353
R1167 VSS.n35 VSS.t168 382.353
R1168 VSS.t26 VSS.n37 382.353
R1169 VSS.t272 VSS.n39 382.353
R1170 VSS.n318 VSS.t28 365.555
R1171 VSS.t0 VSS.n317 365.555
R1172 VSS.t150 VSS.n316 365.555
R1173 VSS.t66 VSS.n315 365.555
R1174 VSS.t182 VSS.n92 365.555
R1175 VSS.t38 VSS.n91 365.555
R1176 VSS.t163 VSS.n90 365.555
R1177 VSS.n86 VSS.t88 365.555
R1178 VSS.n154 VSS.t270 365.555
R1179 VSS.t243 VSS.n143 365.555
R1180 VSS.t51 VSS.n144 365.555
R1181 VSS.n145 VSS.t114 365.555
R1182 VSS.n163 VSS.t238 365.555
R1183 VSS.n162 VSS.t250 365.555
R1184 VSS.n161 VSS.t153 365.555
R1185 VSS.n204 VSS.t94 365.555
R1186 VSS.t69 VSS.n185 365.555
R1187 VSS.t219 VSS.n184 365.555
R1188 VSS.t48 VSS.n183 365.555
R1189 VSS.t44 VSS.n182 365.555
R1190 VSS.n294 VSS.t75 365.555
R1191 VSS.n298 VSS.t22 365.555
R1192 VSS.n299 VSS.t3 365.555
R1193 VSS.n303 VSS.t230 365.555
R1194 VSS.n69 VSS.t257 364.274
R1195 VSS.n116 VSS.t138 364.274
R1196 VSS.t273 VSS.n216 342.106
R1197 VSS.t81 VSS.t188 327.675
R1198 VSS.t171 VSS.t249 310.634
R1199 VSS.t199 VSS.t268 310.634
R1200 VSS.n225 VSS.t119 295.455
R1201 VSS.n226 VSS.t57 295.455
R1202 VSS.n229 VSS.t170 295.455
R1203 VSS.n233 VSS.t237 295.455
R1204 VSS.n235 VSS.t133 295.455
R1205 VSS.n236 VSS.t196 295.455
R1206 VSS.n237 VSS.t169 295.455
R1207 VSS.n238 VSS.t80 295.455
R1208 VSS.n201 VSS.n200 273.747
R1209 VSS.n102 VSS.n101 270.834
R1210 VSS.n2 VSS.t98 255.215
R1211 VSS.n4 VSS.t128 255.215
R1212 VSS.n6 VSS.t59 255.215
R1213 VSS.n8 VSS.t159 255.215
R1214 VSS.t108 VSS.n11 255.215
R1215 VSS.n13 VSS.t179 255.215
R1216 VSS.n15 VSS.t288 255.215
R1217 VSS.n17 VSS.t227 255.215
R1218 VSS.t101 VSS.n280 254.903
R1219 VSS.t210 VSS.n279 254.903
R1220 VSS.n28 VSS.t34 254.903
R1221 VSS.n30 VSS.t234 254.903
R1222 VSS.t111 VSS.n33 254.903
R1223 VSS.n35 VSS.t123 254.903
R1224 VSS.n37 VSS.t192 254.903
R1225 VSS.n39 VSS.t240 254.903
R1226 VSS.n101 VSS.n51 251.548
R1227 VSS.t222 VSS.n225 196.97
R1228 VSS.n226 VSS.t136 196.97
R1229 VSS.n229 VSS.t202 196.97
R1230 VSS.t96 VSS.n233 196.97
R1231 VSS.t13 VSS.n235 196.97
R1232 VSS.n236 VSS.t186 196.97
R1233 VSS.t17 VSS.n237 196.97
R1234 VSS.n238 VSS.t92 196.97
R1235 VSS.n103 VSS.t81 190.587
R1236 VSS.n211 VSS.t269 186.715
R1237 VSS.n191 VSS.t200 186.381
R1238 VSS.n192 VSS.t64 186.381
R1239 VSS.n195 VSS.t171 186.381
R1240 VSS.n199 VSS.t268 186.381
R1241 VSS.n101 VSS.t116 174.407
R1242 VSS.t42 VSS.n211 124.477
R1243 VSS.t62 VSS.n191 124.254
R1244 VSS.n192 VSS.t31 124.254
R1245 VSS.n195 VSS.t78 124.254
R1246 VSS.t104 VSS.n199 124.254
R1247 VSS.n94 VSS.n93 114.236
R1248 VSS.n293 VSS.n290 114.236
R1249 VSS.n260 VSS.n41 106.921
R1250 VSS.t116 VSS.t252 93.9117
R1251 VSS.t19 VSS.t121 58.5375
R1252 VSS.t156 VSS.n129 47.5615
R1253 VSS.t281 VSS.n82 47.5615
R1254 VSS.n138 VSS.t245 36.0732
R1255 VSS.n93 VSS.t254 34.2711
R1256 VSS.t85 VSS.n293 34.2711
R1257 VSS.t224 VSS.n76 34.1511
R1258 VSS.t145 VSS.n123 34.1511
R1259 VSS.n203 VSS.n142 22.5699
R1260 VSS.n259 VSS.t91 20.9066
R1261 VSS.n138 VSS.t54 17.8773
R1262 VSS.n305 VSS.n23 16.8399
R1263 VSS.n103 VSS.n102 16.7186
R1264 VSS.n261 VSS.n260 16.561
R1265 VSS.n187 VSS.n186 16.4146
R1266 VSS.n203 VSS.n202 13.5422
R1267 VSS.t91 VSS.t19 13.1415
R1268 VSS.n141 VSS.t266 9.3736
R1269 VSS.n135 VSS.t12 9.3736
R1270 VSS.n258 VSS.t122 9.3736
R1271 VSS.n292 VSS.n291 9.37275
R1272 VSS.n22 VSS.n21 9.37275
R1273 VSS.n56 VSS.n55 9.37275
R1274 VSS.n105 VSS.t189 9.364
R1275 VSS.n72 VSS.n71 9.3221
R1276 VSS.n79 VSS.t176 9.3221
R1277 VSS.n107 VSS.t204 9.3221
R1278 VSS.n109 VSS.n52 9.3221
R1279 VSS.n119 VSS.n118 9.3221
R1280 VSS.n126 VSS.t218 9.3221
R1281 VSS.n168 VSS.n167 9.30652
R1282 VSS.n74 VSS.n67 9.30652
R1283 VSS.n80 VSS.n66 9.30652
R1284 VSS.n110 VSS.t253 9.30652
R1285 VSS.n263 VSS.t84 9.30652
R1286 VSS.n121 VSS.n114 9.30652
R1287 VSS.n127 VSS.n113 9.30652
R1288 VSS.n212 VSS.n138 8.85568
R1289 VSS VSS.n115 7.30633
R1290 VSS VSS.n68 7.30633
R1291 VSS VSS.t82 7.30633
R1292 VSS.n336 VSS.n5 7.19156
R1293 VSS.n334 VSS.n7 7.19156
R1294 VSS.n327 VSS.n14 7.19156
R1295 VSS.n325 VSS.n16 7.19156
R1296 VSS.n296 VSS.n285 7.19156
R1297 VSS.n284 VSS.n283 7.19156
R1298 VSS.n301 VSS.n282 7.19156
R1299 VSS.n174 VSS.n173 7.19156
R1300 VSS.n177 VSS.n176 7.19156
R1301 VSS.n180 VSS.n179 7.19156
R1302 VSS.n277 VSS.n27 7.19156
R1303 VSS.n275 VSS.n29 7.19156
R1304 VSS.n61 VSS.n60 7.19156
R1305 VSS.n64 VSS.n63 7.19156
R1306 VSS.n88 VSS.n65 7.19156
R1307 VSS.n268 VSS.n36 7.19156
R1308 VSS.n266 VSS.n38 7.19156
R1309 VSS.n244 VSS.t41 7.19156
R1310 VSS.n242 VSS.t214 7.19156
R1311 VSS.n240 VSS.t233 7.19156
R1312 VSS.n252 VSS.t187 7.19156
R1313 VSS.n254 VSS.t14 7.19156
R1314 VSS.n47 VSS.t201 7.19156
R1315 VSS.n45 VSS.t20 7.19156
R1316 VSS.n43 VSS.t207 7.19156
R1317 VSS.n228 VSS.t137 7.19156
R1318 VSS.n223 VSS.t223 7.19156
R1319 VSS.n307 VSS.n306 7.19156
R1320 VSS.n310 VSS.n309 7.19156
R1321 VSS.n313 VSS.n312 7.19156
R1322 VSS.n152 VSS.t271 7.19156
R1323 VSS.n150 VSS.t244 7.19156
R1324 VSS.n148 VSS.t52 7.19156
R1325 VSS.n156 VSS.t239 7.19156
R1326 VSS.n158 VSS.t251 7.19156
R1327 VSS.n159 VSS.t154 7.19156
R1328 VSS.n189 VSS.t63 7.13823
R1329 VSS.n194 VSS.t32 7.13823
R1330 VSS.n209 VSS.t43 7.13323
R1331 VSS.n214 VSS.t127 7.13323
R1332 VSS.n1 VSS.n0 5.91399
R1333 VSS.n338 VSS.n3 5.91399
R1334 VSS.n331 VSS.n10 5.91399
R1335 VSS.n329 VSS.n12 5.91399
R1336 VSS.n287 VSS.n286 5.91399
R1337 VSS.n171 VSS.n166 5.91399
R1338 VSS.n19 VSS.n18 5.91399
R1339 VSS.n26 VSS.n25 5.91399
R1340 VSS.n58 VSS.n57 5.91399
R1341 VSS.n272 VSS.n32 5.91399
R1342 VSS.n270 VSS.n34 5.91399
R1343 VSS.n246 VSS.t148 5.91399
R1344 VSS.n248 VSS.t93 5.91399
R1345 VSS.n250 VSS.t18 5.91399
R1346 VSS.n49 VSS.t135 5.91399
R1347 VSS.n50 VSS.t97 5.91399
R1348 VSS.n231 VSS.t203 5.91399
R1349 VSS.n320 VSS.n20 5.91399
R1350 VSS.n146 VSS.t115 5.91399
R1351 VSS.n206 VSS.t95 5.91399
R1352 VSS.n197 VSS.t79 5.86065
R1353 VSS.n139 VSS.t105 5.86065
R1354 VSS.n137 VSS.t274 5.85565
R1355 VSS.n220 VSS.t107 5.85565
R1356 VSS.n70 VSS.n69 5.2005
R1357 VSS.n76 VSS.n75 5.2005
R1358 VSS.n78 VSS.n77 5.2005
R1359 VSS.n82 VSS.n81 5.2005
R1360 VSS.n104 VSS.n103 5.2005
R1361 VSS.n111 VSS.n51 5.2005
R1362 VSS.n319 VSS.n318 5.2005
R1363 VSS.n317 VSS.n308 5.2005
R1364 VSS.n316 VSS.n311 5.2005
R1365 VSS.n315 VSS.n314 5.2005
R1366 VSS.n92 VSS.n59 5.2005
R1367 VSS.n91 VSS.n62 5.2005
R1368 VSS.n90 VSS.n89 5.2005
R1369 VSS.n87 VSS.n86 5.2005
R1370 VSS.n93 VSS.n56 5.2005
R1371 VSS.n245 VSS.n41 5.2005
R1372 VSS.n243 VSS.n41 5.2005
R1373 VSS.n241 VSS.n41 5.2005
R1374 VSS.n239 VSS.n41 5.2005
R1375 VSS.n48 VSS.n41 5.2005
R1376 VSS.n46 VSS.n41 5.2005
R1377 VSS.n44 VSS.n41 5.2005
R1378 VSS.n42 VSS.n41 5.2005
R1379 VSS.n259 VSS.n258 5.2005
R1380 VSS.n225 VSS.n224 5.2005
R1381 VSS.n227 VSS.n226 5.2005
R1382 VSS.n230 VSS.n229 5.2005
R1383 VSS.n233 VSS.n232 5.2005
R1384 VSS.n255 VSS.n235 5.2005
R1385 VSS.n253 VSS.n236 5.2005
R1386 VSS.n251 VSS.n237 5.2005
R1387 VSS.n249 VSS.n238 5.2005
R1388 VSS.n262 VSS.n261 5.2005
R1389 VSS.n265 VSS.n39 5.2005
R1390 VSS.n267 VSS.n37 5.2005
R1391 VSS.n269 VSS.n35 5.2005
R1392 VSS.n271 VSS.n33 5.2005
R1393 VSS.n274 VSS.n30 5.2005
R1394 VSS.n276 VSS.n28 5.2005
R1395 VSS.n279 VSS.n278 5.2005
R1396 VSS.n280 VSS.n24 5.2005
R1397 VSS.n23 VSS.n22 5.2005
R1398 VSS.n135 VSS.n134 5.2005
R1399 VSS.n154 VSS.n153 5.2005
R1400 VSS.n151 VSS.n143 5.2005
R1401 VSS.n149 VSS.n144 5.2005
R1402 VSS.n147 VSS.n145 5.2005
R1403 VSS.n216 VSS.n215 5.2005
R1404 VSS.n163 VSS.n155 5.2005
R1405 VSS.n162 VSS.n157 5.2005
R1406 VSS.n161 VSS.n160 5.2005
R1407 VSS.n205 VSS.n204 5.2005
R1408 VSS.n142 VSS.n141 5.2005
R1409 VSS.n199 VSS.n198 5.2005
R1410 VSS.n196 VSS.n195 5.2005
R1411 VSS.n193 VSS.n192 5.2005
R1412 VSS.n191 VSS.n190 5.2005
R1413 VSS.n187 VSS.n165 5.2005
R1414 VSS.n185 VSS.n172 5.2005
R1415 VSS.n184 VSS.n175 5.2005
R1416 VSS.n183 VSS.n178 5.2005
R1417 VSS.n182 VSS.n181 5.2005
R1418 VSS.n295 VSS.n294 5.2005
R1419 VSS.n298 VSS.n297 5.2005
R1420 VSS.n300 VSS.n299 5.2005
R1421 VSS.n303 VSS.n302 5.2005
R1422 VSS.n293 VSS.n292 5.2005
R1423 VSS.n211 VSS.n210 5.2005
R1424 VSS.n117 VSS.n116 5.2005
R1425 VSS.n123 VSS.n122 5.2005
R1426 VSS.n125 VSS.n124 5.2005
R1427 VSS.n129 VSS.n128 5.2005
R1428 VSS.n339 VSS.n2 5.2005
R1429 VSS.n337 VSS.n4 5.2005
R1430 VSS.n335 VSS.n6 5.2005
R1431 VSS.n333 VSS.n8 5.2005
R1432 VSS.n330 VSS.n11 5.2005
R1433 VSS.n328 VSS.n13 5.2005
R1434 VSS.n326 VSS.n15 5.2005
R1435 VSS.n324 VSS.n17 5.2005
R1436 VSS.n305 VSS.n304 3.36838
R1437 VSS.n260 VSS.n259 2.38977
R1438 VSS.n323 VSS 2.24014
R1439 VSS.n264 VSS.n263 2.2128
R1440 VSS VSS.n222 2.14127
R1441 VSS VSS.n264 1.91938
R1442 VSS.n169 VSS.n168 1.36907
R1443 VSS.n248 VSS.n247 1.03389
R1444 VSS.n257 VSS.n256 0.846463
R1445 VSS.n332 VSS.n9 0.845914
R1446 VSS.n170 VSS.n169 0.845914
R1447 VSS.n273 VSS.n31 0.845914
R1448 VSS.n322 VSS.n321 0.845914
R1449 VSS.n208 VSS.n207 0.819492
R1450 VSS.n221 VSS.n136 0.817015
R1451 VSS.n230 VSS.n228 0.480225
R1452 VSS.n232 VSS.n231 0.480225
R1453 VSS.n252 VSS.n251 0.480225
R1454 VSS.n250 VSS.n249 0.480225
R1455 VSS VSS.n208 0.473
R1456 VSS.n222 VSS 0.438387
R1457 VSS.n264 VSS 0.413056
R1458 VSS.n196 VSS.n194 0.363625
R1459 VSS.n198 VSS.n197 0.363625
R1460 VSS.n215 VSS.n214 0.363625
R1461 VSS.n219 VSS.n137 0.363625
R1462 VSS VSS.n284 0.343161
R1463 VSS.n301 VSS 0.343161
R1464 VSS.n177 VSS 0.343161
R1465 VSS.n180 VSS 0.343161
R1466 VSS.n64 VSS 0.343161
R1467 VSS VSS.n88 0.343161
R1468 VSS VSS.n240 0.343161
R1469 VSS VSS.n242 0.343161
R1470 VSS VSS.n43 0.343161
R1471 VSS VSS.n45 0.343161
R1472 VSS.n223 VSS 0.343161
R1473 VSS.n254 VSS 0.343161
R1474 VSS.n310 VSS 0.343161
R1475 VSS.n313 VSS 0.343161
R1476 VSS.n152 VSS 0.343161
R1477 VSS.n150 VSS 0.343161
R1478 VSS VSS.n156 0.343161
R1479 VSS VSS.n158 0.343161
R1480 VSS.n73 VSS.n72 0.310174
R1481 VSS.n120 VSS.n119 0.310174
R1482 VSS.n107 VSS.n106 0.309418
R1483 VSS.n222 VSS.n221 0.3055
R1484 VSS VSS.n295 0.289491
R1485 VSS VSS.n172 0.289491
R1486 VSS VSS.n59 0.289491
R1487 VSS.n245 VSS 0.289491
R1488 VSS.n48 VSS 0.289491
R1489 VSS.n319 VSS 0.289491
R1490 VSS VSS.n147 0.289491
R1491 VSS.n205 VSS 0.289491
R1492 VSS.n189 VSS 0.259875
R1493 VSS.n209 VSS 0.259875
R1494 VSS.n120 VSS.n117 0.255008
R1495 VSS.n73 VSS.n70 0.255008
R1496 VSS.n106 VSS.n53 0.254245
R1497 VSS.n296 VSS 0.191234
R1498 VSS.n174 VSS 0.191234
R1499 VSS.n61 VSS 0.191234
R1500 VSS VSS.n244 0.191234
R1501 VSS VSS.n47 0.191234
R1502 VSS.n307 VSS 0.191234
R1503 VSS.n148 VSS 0.191234
R1504 VSS.n159 VSS 0.191234
R1505 VSS.n256 VSS.n50 0.187931
R1506 VSS.n256 VSS 0.183803
R1507 VSS.n110 VSS.n109 0.168119
R1508 VSS.n80 VSS.n79 0.168072
R1509 VSS.n127 VSS.n126 0.168072
R1510 VSS.n74 VSS.n73 0.142796
R1511 VSS.n121 VSS.n120 0.142796
R1512 VSS.n208 VSS.n139 0.142375
R1513 VSS.n221 VSS.n220 0.142375
R1514 VSS.n106 VSS.n105 0.141455
R1515 VSS VSS.n9 0.137685
R1516 VSS.n170 VSS 0.137685
R1517 VSS.n207 VSS 0.137685
R1518 VSS.n136 VSS 0.137685
R1519 VSS.n321 VSS 0.137685
R1520 VSS VSS.n31 0.137685
R1521 VSS.n79 VSS.n78 0.137391
R1522 VSS.n126 VSS.n125 0.137391
R1523 VSS VSS.n257 0.137136
R1524 VSS.n247 VSS 0.137136
R1525 VSS.n109 VSS.n108 0.136634
R1526 VSS.n339 VSS.n338 0.130899
R1527 VSS.n337 VSS.n336 0.130899
R1528 VSS.n330 VSS.n329 0.130899
R1529 VSS.n328 VSS.n327 0.130899
R1530 VSS.n26 VSS.n24 0.130575
R1531 VSS.n278 VSS.n277 0.130575
R1532 VSS.n271 VSS.n270 0.130575
R1533 VSS.n269 VSS.n268 0.130575
R1534 VSS.n297 VSS.n296 0.118573
R1535 VSS.n300 VSS.n284 0.118573
R1536 VSS.n302 VSS.n301 0.118573
R1537 VSS.n175 VSS.n174 0.118573
R1538 VSS.n178 VSS.n177 0.118573
R1539 VSS.n181 VSS.n180 0.118573
R1540 VSS.n62 VSS.n61 0.118573
R1541 VSS.n89 VSS.n64 0.118573
R1542 VSS.n88 VSS.n87 0.118573
R1543 VSS.n240 VSS.n239 0.118573
R1544 VSS.n242 VSS.n241 0.118573
R1545 VSS.n244 VSS.n243 0.118573
R1546 VSS.n43 VSS.n42 0.118573
R1547 VSS.n45 VSS.n44 0.118573
R1548 VSS.n47 VSS.n46 0.118573
R1549 VSS.n224 VSS.n223 0.118573
R1550 VSS.n228 VSS.n227 0.118573
R1551 VSS.n255 VSS.n254 0.118573
R1552 VSS.n253 VSS.n252 0.118573
R1553 VSS.n308 VSS.n307 0.118573
R1554 VSS.n311 VSS.n310 0.118573
R1555 VSS.n314 VSS.n313 0.118573
R1556 VSS.n153 VSS.n152 0.118573
R1557 VSS.n151 VSS.n150 0.118573
R1558 VSS.n149 VSS.n148 0.118573
R1559 VSS.n156 VSS.n155 0.118573
R1560 VSS.n158 VSS.n157 0.118573
R1561 VSS.n160 VSS.n159 0.118573
R1562 VSS.n323 VSS 0.116501
R1563 VSS VSS.n107 0.115458
R1564 VSS VSS.n287 0.115271
R1565 VSS VSS.n171 0.115271
R1566 VSS VSS.n58 0.115271
R1567 VSS.n246 VSS 0.115271
R1568 VSS.n49 VSS 0.115271
R1569 VSS.n231 VSS 0.115271
R1570 VSS VSS.n50 0.115271
R1571 VSS VSS.n250 0.115271
R1572 VSS VSS.n248 0.115271
R1573 VSS.n320 VSS 0.115271
R1574 VSS VSS.n146 0.115271
R1575 VSS.n206 VSS 0.115271
R1576 VSS.n72 VSS 0.114702
R1577 VSS.n119 VSS 0.114702
R1578 VSS.n287 VSS.n9 0.10206
R1579 VSS.n171 VSS.n170 0.10206
R1580 VSS.n58 VSS.n31 0.10206
R1581 VSS.n247 VSS.n246 0.10206
R1582 VSS.n257 VSS.n49 0.10206
R1583 VSS.n321 VSS.n320 0.10206
R1584 VSS.n146 VSS.n136 0.10206
R1585 VSS.n207 VSS.n206 0.10206
R1586 VSS VSS.n334 0.0936421
R1587 VSS VSS.n325 0.0936421
R1588 VSS VSS.n275 0.0934104
R1589 VSS VSS.n266 0.0934104
R1590 VSS VSS.n323 0.09252
R1591 VSS.n190 VSS.n189 0.089875
R1592 VSS.n194 VSS.n193 0.089875
R1593 VSS.n210 VSS.n209 0.089875
R1594 VSS.n214 VSS.n213 0.089875
R1595 VSS.n197 VSS 0.087375
R1596 VSS VSS.n139 0.087375
R1597 VSS VSS.n137 0.087375
R1598 VSS.n220 VSS 0.087375
R1599 VSS.n263 VSS.n262 0.0675755
R1600 VSS.n168 VSS.n165 0.0667264
R1601 VSS.n75 VSS.n74 0.0667264
R1602 VSS.n122 VSS.n121 0.0667264
R1603 VSS.n105 VSS.n104 0.0589403
R1604 VSS.n111 VSS.n110 0.0564843
R1605 VSS.n81 VSS.n80 0.0557756
R1606 VSS.n128 VSS.n127 0.0557756
R1607 VSS VSS.n322 0.0526154
R1608 VSS.n169 VSS.n1 0.0512232
R1609 VSS.n332 VSS.n331 0.0512232
R1610 VSS.n322 VSS.n19 0.051097
R1611 VSS.n273 VSS.n272 0.051097
R1612 VSS VSS.n332 0.0505499
R1613 VSS VSS.n273 0.0504254
R1614 VSS.n336 VSS.n335 0.0325948
R1615 VSS.n334 VSS.n333 0.0325948
R1616 VSS.n327 VSS.n326 0.0325948
R1617 VSS.n325 VSS.n324 0.0325948
R1618 VSS.n277 VSS.n276 0.0325149
R1619 VSS.n275 VSS.n274 0.0325149
R1620 VSS.n268 VSS.n267 0.0325149
R1621 VSS.n266 VSS.n265 0.0325149
R1622 VSS VSS.n1 0.031697
R1623 VSS.n338 VSS 0.031697
R1624 VSS.n331 VSS 0.031697
R1625 VSS.n329 VSS 0.031697
R1626 VSS VSS.n19 0.0316194
R1627 VSS VSS.n26 0.0316194
R1628 VSS.n272 VSS 0.0316194
R1629 VSS.n270 VSS 0.0316194
R1630 VSS.n297 VSS 0.00545413
R1631 VSS VSS.n300 0.00545413
R1632 VSS.n302 VSS 0.00545413
R1633 VSS VSS.n175 0.00545413
R1634 VSS VSS.n178 0.00545413
R1635 VSS.n181 VSS 0.00545413
R1636 VSS VSS.n62 0.00545413
R1637 VSS.n89 VSS 0.00545413
R1638 VSS.n87 VSS 0.00545413
R1639 VSS.n239 VSS 0.00545413
R1640 VSS.n241 VSS 0.00545413
R1641 VSS.n243 VSS 0.00545413
R1642 VSS.n42 VSS 0.00545413
R1643 VSS.n44 VSS 0.00545413
R1644 VSS.n46 VSS 0.00545413
R1645 VSS.n224 VSS 0.00545413
R1646 VSS.n227 VSS 0.00545413
R1647 VSS VSS.n255 0.00545413
R1648 VSS VSS.n253 0.00545413
R1649 VSS VSS.n308 0.00545413
R1650 VSS VSS.n311 0.00545413
R1651 VSS.n314 VSS 0.00545413
R1652 VSS.n153 VSS 0.00545413
R1653 VSS VSS.n151 0.00545413
R1654 VSS VSS.n149 0.00545413
R1655 VSS.n155 VSS 0.00545413
R1656 VSS.n157 VSS 0.00545413
R1657 VSS.n160 VSS 0.00545413
R1658 VSS.n190 VSS 0.00425
R1659 VSS.n193 VSS 0.00425
R1660 VSS.n210 VSS 0.00425
R1661 VSS.n213 VSS 0.00425
R1662 VSS.n117 VSS 0.00380275
R1663 VSS.n295 VSS 0.00380275
R1664 VSS.n172 VSS 0.00380275
R1665 VSS.n59 VSS 0.00380275
R1666 VSS.n70 VSS 0.00380275
R1667 VSS VSS.n245 0.00380275
R1668 VSS.n53 VSS 0.00380275
R1669 VSS VSS.n48 0.00380275
R1670 VSS VSS.n230 0.00380275
R1671 VSS.n232 VSS 0.00380275
R1672 VSS.n251 VSS 0.00380275
R1673 VSS.n249 VSS 0.00380275
R1674 VSS VSS.n319 0.00380275
R1675 VSS.n147 VSS 0.00380275
R1676 VSS VSS.n205 0.00380275
R1677 VSS.n78 VSS 0.00352521
R1678 VSS.n108 VSS 0.00352521
R1679 VSS.n125 VSS 0.00352521
R1680 VSS VSS.n196 0.003
R1681 VSS.n198 VSS 0.003
R1682 VSS.n215 VSS 0.003
R1683 VSS VSS.n219 0.003
R1684 VSS.n292 VSS 0.00219811
R1685 VSS VSS.n165 0.00219811
R1686 VSS.n141 VSS 0.00219811
R1687 VSS VSS.n135 0.00219811
R1688 VSS.n22 VSS 0.00219811
R1689 VSS.n56 VSS 0.00219811
R1690 VSS.n75 VSS 0.00219811
R1691 VSS.n104 VSS 0.00219811
R1692 VSS.n258 VSS 0.00219811
R1693 VSS.n262 VSS 0.00219811
R1694 VSS.n122 VSS 0.00219811
R1695 VSS.n81 VSS 0.00191732
R1696 VSS VSS.n111 0.00191732
R1697 VSS.n128 VSS 0.00191732
R1698 VSS.n335 VSS 0.00184663
R1699 VSS.n333 VSS 0.00184663
R1700 VSS.n326 VSS 0.00184663
R1701 VSS.n324 VSS 0.00184663
R1702 VSS.n276 VSS 0.00184328
R1703 VSS.n274 VSS 0.00184328
R1704 VSS.n267 VSS 0.00184328
R1705 VSS.n265 VSS 0.00184328
R1706 VSS VSS.n339 0.00139776
R1707 VSS VSS.n337 0.00139776
R1708 VSS VSS.n330 0.00139776
R1709 VSS VSS.n328 0.00139776
R1710 VSS.n24 VSS 0.00139552
R1711 VSS.n278 VSS 0.00139552
R1712 VSS VSS.n271 0.00139552
R1713 VSS VSS.n269 0.00139552
R1714 CLK_div_3_mag_1.CLK.n7 CLK_div_3_mag_1.CLK.t11 36.935
R1715 CLK_div_3_mag_1.CLK.n6 CLK_div_3_mag_1.CLK.t7 36.935
R1716 CLK_div_3_mag_1.CLK.n11 CLK_div_3_mag_1.CLK.t6 36.935
R1717 CLK_div_3_mag_1.CLK.n10 CLK_div_3_mag_1.CLK.t12 36.935
R1718 CLK_div_3_mag_1.CLK.n8 CLK_div_3_mag_1.CLK.t15 30.6315
R1719 CLK_div_3_mag_1.CLK.n15 CLK_div_3_mag_1.CLK.t8 25.5361
R1720 CLK_div_3_mag_1.CLK.n12 CLK_div_3_mag_1.CLK.t13 25.5361
R1721 CLK_div_3_mag_1.CLK.n8 CLK_div_3_mag_1.CLK.t5 21.7275
R1722 CLK_div_3_mag_1.CLK.n7 CLK_div_3_mag_1.CLK.t9 18.1962
R1723 CLK_div_3_mag_1.CLK.n6 CLK_div_3_mag_1.CLK.t3 18.1962
R1724 CLK_div_3_mag_1.CLK.n11 CLK_div_3_mag_1.CLK.t2 18.1962
R1725 CLK_div_3_mag_1.CLK.n10 CLK_div_3_mag_1.CLK.t10 18.1962
R1726 CLK_div_3_mag_1.CLK.n15 CLK_div_3_mag_1.CLK.t14 14.0734
R1727 CLK_div_3_mag_1.CLK.n12 CLK_div_3_mag_1.CLK.t4 14.0734
R1728 CLK_div_3_mag_1.CLK.n5 CLK_div_3_mag_1.CLK.t1 9.33985
R1729 CLK_div_3_mag_1.CLK.n0 CLK_div_3_mag_1.CLK.n9 7.41366
R1730 CLK_div_3_mag_1.CLK.n14 CLK_div_3_mag_1.CLK.n13 5.37352
R1731 CLK_div_3_mag_1.CLK.n5 CLK_div_3_mag_1.CLK.t0 5.17836
R1732 CLK_div_3_mag_1.CLK.n7 CLK_div_3_mag_1.CLK 2.13258
R1733 CLK_div_3_mag_1.CLK.n2 CLK_div_3_mag_1.CLK.n0 1.11745
R1734 CLK_div_3_mag_1.CLK.n2 CLK_div_3_mag_1.CLK.n11 2.13258
R1735 CLK_div_3_mag_1.CLK.n9 CLK_div_3_mag_1.CLK.n8 1.80525
R1736 CLK_div_3_mag_1.CLK.n1 CLK_div_3_mag_1.CLK 2.63808
R1737 CLK_div_3_mag_1.CLK.n0 CLK_div_3_mag_1.CLK 2.51975
R1738 CLK_div_3_mag_1.CLK CLK_div_3_mag_1.CLK.n10 2.13055
R1739 CLK_div_3_mag_1.CLK CLK_div_3_mag_1.CLK.n6 2.13055
R1740 CLK_div_3_mag_1.CLK.n3 CLK_div_3_mag_1.CLK.n12 1.43653
R1741 CLK_div_3_mag_1.CLK.n4 CLK_div_3_mag_1.CLK.n15 1.43653
R1742 CLK_div_3_mag_1.CLK.n3 CLK_div_3_mag_1.CLK 0.196042
R1743 CLK_div_3_mag_1.CLK CLK_div_3_mag_1.CLK.n4 0.196042
R1744 CLK_div_3_mag_1.CLK CLK_div_3_mag_1.CLK.n5 0.115328
R1745 CLK_div_3_mag_1.CLK.n9 CLK_div_3_mag_1.CLK 0.108371
R1746 CLK_div_3_mag_1.CLK.n2 CLK_div_3_mag_1.CLK 0.0763652
R1747 CLK_div_3_mag_1.CLK.n13 CLK_div_3_mag_1.CLK.n3 1.19546
R1748 CLK_div_3_mag_1.CLK.n4 CLK_div_3_mag_1.CLK.n14 1.19546
R1749 CLK_div_3_mag_1.CLK CLK_div_3_mag_1.CLK.n1 1.11745
R1750 CLK_div_3_mag_1.CLK.n13 CLK_div_3_mag_1.CLK.n0 1.01362
R1751 CLK_div_3_mag_1.CLK.n14 CLK_div_3_mag_1.CLK.n1 0.895294
R1752 CLK_div_3_mag_2.Q1.n5 CLK_div_3_mag_2.Q1.t10 36.935
R1753 CLK_div_3_mag_2.Q1.n4 CLK_div_3_mag_2.Q1.t4 31.4332
R1754 CLK_div_3_mag_2.Q1.n6 CLK_div_3_mag_2.Q1.t9 31.4332
R1755 CLK_div_3_mag_2.Q1.n3 CLK_div_3_mag_2.Q1.t5 30.5184
R1756 CLK_div_3_mag_2.Q1.n3 CLK_div_3_mag_2.Q1.t7 24.7029
R1757 CLK_div_3_mag_2.Q1.n5 CLK_div_3_mag_2.Q1.t8 18.1962
R1758 CLK_div_3_mag_2.Q1.n4 CLK_div_3_mag_2.Q1.t3 15.3826
R1759 CLK_div_3_mag_2.Q1.n6 CLK_div_3_mag_2.Q1.t6 15.3826
R1760 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.Q1.t1 7.09905
R1761 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.Q1.n6 6.86134
R1762 CLK_div_3_mag_2.Q1.n7 CLK_div_3_mag_2.Q1 5.0096
R1763 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.Q1.n0 8.55639
R1764 CLK_div_3_mag_2.Q1.n4 CLK_div_3_mag_2.Q1 5.69501
R1765 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.Q1.n2 3.25226
R1766 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.Q1.n8 2.43532
R1767 CLK_div_3_mag_2.Q1.n2 CLK_div_3_mag_2.Q1.t2 2.2755
R1768 CLK_div_3_mag_2.Q1.n2 CLK_div_3_mag_2.Q1.n1 2.2755
R1769 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.Q1.n5 2.13479
R1770 CLK_div_3_mag_2.Q1 CLK_div_3_mag_2.Q1.n3 1.81225
R1771 CLK_div_3_mag_2.Q1.n8 CLK_div_3_mag_2.Q1.n7 1.45511
R1772 CLK_div_3_mag_2.Q1.n8 CLK_div_3_mag_2.Q1.n0 1.23718
R1773 CLK_div_3_mag_2.Q1.n7 CLK_div_3_mag_2.Q1 1.12056
R1774 CLK_div_3_mag_2.Q1.n0 CLK_div_3_mag_2.Q1 0.976034
R1775 CLK_div_3_mag_2.JK_FF_mag_1.K.n5 CLK_div_3_mag_2.JK_FF_mag_1.K.t7 37.1984
R1776 CLK_div_3_mag_2.JK_FF_mag_1.K.n4 CLK_div_3_mag_2.JK_FF_mag_1.K.t5 31.4332
R1777 CLK_div_3_mag_2.JK_FF_mag_1.K.n3 CLK_div_3_mag_2.JK_FF_mag_1.K.t2 30.5184
R1778 CLK_div_3_mag_2.JK_FF_mag_1.K.n3 CLK_div_3_mag_2.JK_FF_mag_1.K.t4 24.7029
R1779 CLK_div_3_mag_2.JK_FF_mag_1.K.n5 CLK_div_3_mag_2.JK_FF_mag_1.K.t6 17.6618
R1780 CLK_div_3_mag_2.JK_FF_mag_1.K.n4 CLK_div_3_mag_2.JK_FF_mag_1.K.t3 15.3826
R1781 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_3_mag_2.JK_FF_mag_1.K 12.0839
R1782 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_3_mag_2.JK_FF_mag_1.K.n4 9.86691
R1783 CLK_div_3_mag_2.JK_FF_mag_1.K.n6 CLK_div_3_mag_2.JK_FF_mag_1.K 6.09789
R1784 CLK_div_3_mag_2.JK_FF_mag_1.K.n7 CLK_div_3_mag_2.JK_FF_mag_1.K.n2 2.99416
R1785 CLK_div_3_mag_2.JK_FF_mag_1.K.n2 CLK_div_3_mag_2.JK_FF_mag_1.K.t1 2.2755
R1786 CLK_div_3_mag_2.JK_FF_mag_1.K.n2 CLK_div_3_mag_2.JK_FF_mag_1.K.n1 2.2755
R1787 CLK_div_3_mag_2.JK_FF_mag_1.K.n7 CLK_div_3_mag_2.JK_FF_mag_1.K.n6 2.2505
R1788 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 CLK_div_3_mag_2.JK_FF_mag_1.K 2.24134
R1789 CLK_div_3_mag_2.JK_FF_mag_1.K.n6 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 1.93723
R1790 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.K.n3 1.81224
R1791 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.K.n5 1.43718
R1792 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.K.n7 0.4325
R1793 CLK.n8 CLK.t5 36.935
R1794 CLK.n1 CLK.t4 36.935
R1795 CLK.n23 CLK.t11 36.935
R1796 CLK.n15 CLK.t8 36.935
R1797 CLK.n13 CLK.t12 30.6315
R1798 CLK.n37 CLK.t7 25.5361
R1799 CLK.n30 CLK.t10 25.5361
R1800 CLK.n13 CLK.t3 21.7275
R1801 CLK.n8 CLK.t2 18.1962
R1802 CLK.n1 CLK.t1 18.1962
R1803 CLK.n23 CLK.t9 18.1962
R1804 CLK.n15 CLK.t6 18.1962
R1805 CLK.n37 CLK.t13 14.0734
R1806 CLK.n30 CLK.t0 14.0734
R1807 CLK.n21 CLK.n14 7.41366
R1808 CLK.n35 CLK.n34 5.37352
R1809 CLK.n12 CLK.n11 2.25107
R1810 CLK.n27 CLK.n26 2.25107
R1811 CLK.n33 CLK.n32 2.24385
R1812 CLK.n39 CLK.n36 2.24385
R1813 CLK.n9 CLK.n8 2.12207
R1814 CLK.n24 CLK.n23 2.12207
R1815 CLK.n2 CLK.n1 2.12188
R1816 CLK.n16 CLK.n15 2.12188
R1817 CLK.n14 CLK.n13 1.80525
R1818 CLK.n7 CLK.n6 1.74297
R1819 CLK.n21 CLK.n20 1.62464
R1820 CLK.n6 CLK.n4 1.49778
R1821 CLK.n20 CLK.n18 1.49778
R1822 CLK.n31 CLK.n30 1.42775
R1823 CLK.n38 CLK.n37 1.42775
R1824 CLK.n35 CLK.n12 0.882596
R1825 CLK.n34 CLK.n27 0.882596
R1826 CLK.n29 CLK 0.1605
R1827 CLK.n22 CLK.n21 0.118826
R1828 CLK.n14 CLK 0.108371
R1829 CLK.n34 CLK.n33 0.0726935
R1830 CLK.n36 CLK.n35 0.0726935
R1831 CLK CLK.n40 0.05925
R1832 CLK.n10 CLK 0.0457995
R1833 CLK.n3 CLK 0.0457995
R1834 CLK.n25 CLK 0.0457995
R1835 CLK.n17 CLK 0.0457995
R1836 CLK.n11 CLK.n10 0.0377414
R1837 CLK.n4 CLK.n3 0.0377414
R1838 CLK.n26 CLK.n25 0.0377414
R1839 CLK.n18 CLK.n17 0.0377414
R1840 CLK.n32 CLK.n29 0.03175
R1841 CLK.n40 CLK.n39 0.03175
R1842 CLK.n33 CLK.n28 0.0205196
R1843 CLK.n36 CLK.n0 0.0205196
R1844 CLK.n6 CLK.n5 0.0131772
R1845 CLK.n20 CLK.n19 0.0131772
R1846 CLK.n12 CLK.n7 0.0122182
R1847 CLK.n27 CLK.n22 0.0122182
R1848 CLK.n11 CLK.n9 0.00360345
R1849 CLK.n4 CLK.n2 0.00360345
R1850 CLK.n26 CLK.n24 0.00360345
R1851 CLK.n18 CLK.n16 0.00360345
R1852 CLK.n32 CLK.n31 0.00175
R1853 CLK.n39 CLK.n38 0.00175
R1854 CLK_div_3_mag_0.CLK.n10 CLK_div_3_mag_0.CLK.t8 36.935
R1855 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.t11 36.935
R1856 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.t5 36.935
R1857 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK.t2 36.935
R1858 CLK_div_3_mag_0.CLK.n12 CLK_div_3_mag_0.CLK.t13 30.5752
R1859 CLK_div_3_mag_0.CLK.n18 CLK_div_3_mag_0.CLK.t12 25.4742
R1860 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK.t6 25.4742
R1861 CLK_div_3_mag_0.CLK.n12 CLK_div_3_mag_0.CLK.t14 21.7814
R1862 CLK_div_3_mag_0.CLK.n10 CLK_div_3_mag_0.CLK.t7 18.1962
R1863 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.t10 18.1962
R1864 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.t4 18.1962
R1865 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK.t3 18.1962
R1866 CLK_div_3_mag_0.CLK.n18 CLK_div_3_mag_0.CLK.t15 14.142
R1867 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK.t9 14.142
R1868 CLK_div_3_mag_0.CLK.n8 CLK_div_3_mag_0.CLK.t1 9.33985
R1869 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n13 7.41653
R1870 CLK_div_3_mag_0.CLK.n17 CLK_div_3_mag_0.CLK.n16 5.37091
R1871 CLK_div_3_mag_0.CLK.n8 CLK_div_3_mag_0.CLK.t0 5.17836
R1872 CLK_div_3_mag_0.CLK.n9 CLK_div_3_mag_0.CLK.n4 2.13175
R1873 CLK_div_3_mag_0.CLK.n3 CLK_div_3_mag_0.CLK.n2 1.11873
R1874 CLK_div_3_mag_0.CLK.n11 CLK_div_3_mag_0.CLK.n5 2.13275
R1875 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n1 0.0786548
R1876 CLK_div_3_mag_0.CLK.n14 CLK_div_3_mag_0.CLK.n1 2.13252
R1877 CLK_div_3_mag_0.CLK.n15 CLK_div_3_mag_0.CLK.n6 1.42979
R1878 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK.n18 1.42979
R1879 CLK_div_3_mag_0.CLK.n7 CLK_div_3_mag_0.CLK.n17 1.19668
R1880 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n1 1.11863
R1881 CLK_div_3_mag_0.CLK.n3 CLK_div_3_mag_0.CLK.n10 2.13252
R1882 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK.n12 1.80834
R1883 CLK_div_3_mag_0.CLK.n2 CLK_div_3_mag_0.CLK.n4 2.63066
R1884 CLK_div_3_mag_0.CLK.n0 CLK_div_3_mag_0.CLK.n5 2.51833
R1885 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n5 0.0794261
R1886 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n8 0.115328
R1887 CLK_div_3_mag_0.CLK.n13 CLK_div_3_mag_0.CLK 0.105738
R1888 CLK_div_3_mag_0.CLK.n4 CLK_div_3_mag_0.CLK 0.0794261
R1889 CLK_div_3_mag_0.CLK.n3 CLK_div_3_mag_0.CLK 0.0786538
R1890 CLK_div_3_mag_0.CLK CLK_div_3_mag_0.CLK.n7 0.19529
R1891 CLK_div_3_mag_0.CLK.n6 CLK_div_3_mag_0.CLK 0.19529
R1892 CLK_div_3_mag_0.CLK.n16 CLK_div_3_mag_0.CLK.n6 1.19668
R1893 CLK_div_3_mag_0.CLK.n16 CLK_div_3_mag_0.CLK.n0 1.01264
R1894 CLK_div_3_mag_0.CLK.n17 CLK_div_3_mag_0.CLK.n2 0.890034
R1895 CLK_div_3_mag_2.Q0.n3 CLK_div_3_mag_2.Q0.t6 36.935
R1896 CLK_div_3_mag_2.Q0.n4 CLK_div_3_mag_2.Q0.t4 31.4332
R1897 CLK_div_3_mag_2.Q0.n2 CLK_div_3_mag_2.Q0.t3 29.8635
R1898 CLK_div_3_mag_2.Q0.n2 CLK_div_3_mag_2.Q0.t7 27.7543
R1899 CLK_div_3_mag_2.Q0.n3 CLK_div_3_mag_2.Q0.t5 18.1962
R1900 CLK_div_3_mag_2.Q0.n4 CLK_div_3_mag_2.Q0.t8 15.3826
R1901 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.Q0.t2 7.09905
R1902 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.Q0.n4 6.86134
R1903 CLK_div_3_mag_2.Q0.n5 CLK_div_3_mag_2.Q0 5.0096
R1904 CLK_div_3_mag_2.Q0.n6 CLK_div_3_mag_2.Q0 3.41823
R1905 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.Q0.n1 3.25226
R1906 CLK_div_3_mag_2.Q0.n1 CLK_div_3_mag_2.Q0.t0 2.2755
R1907 CLK_div_3_mag_2.Q0.n1 CLK_div_3_mag_2.Q0.n0 2.2755
R1908 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.Q0.n6 2.2505
R1909 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.Q0.n3 2.13479
R1910 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.Q0.n2 1.7371
R1911 CLK_div_3_mag_2.Q0.n6 CLK_div_3_mag_2.Q0.n5 1.50498
R1912 CLK_div_3_mag_2.Q0.n5 CLK_div_3_mag_2.Q0 1.12056
R1913 CLK_div_3_mag_1.Q1.n5 CLK_div_3_mag_1.Q1.t10 36.935
R1914 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1.t5 31.4332
R1915 CLK_div_3_mag_1.Q1.n6 CLK_div_3_mag_1.Q1.t6 31.4332
R1916 CLK_div_3_mag_1.Q1.n3 CLK_div_3_mag_1.Q1.t7 30.5184
R1917 CLK_div_3_mag_1.Q1.n3 CLK_div_3_mag_1.Q1.t8 24.7029
R1918 CLK_div_3_mag_1.Q1.n5 CLK_div_3_mag_1.Q1.t9 18.1962
R1919 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1.t3 15.3826
R1920 CLK_div_3_mag_1.Q1.n6 CLK_div_3_mag_1.Q1.t4 15.3826
R1921 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.t2 7.09905
R1922 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n6 6.86134
R1923 CLK_div_3_mag_1.Q1.n7 CLK_div_3_mag_1.Q1 5.0096
R1924 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n0 8.55639
R1925 CLK_div_3_mag_1.Q1.n4 CLK_div_3_mag_1.Q1 5.69501
R1926 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n2 3.25226
R1927 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n8 2.43532
R1928 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1.t0 2.2755
R1929 CLK_div_3_mag_1.Q1.n2 CLK_div_3_mag_1.Q1.n1 2.2755
R1930 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n5 2.13479
R1931 CLK_div_3_mag_1.Q1 CLK_div_3_mag_1.Q1.n3 1.81225
R1932 CLK_div_3_mag_1.Q1.n8 CLK_div_3_mag_1.Q1.n7 1.45511
R1933 CLK_div_3_mag_1.Q1.n8 CLK_div_3_mag_1.Q1.n0 1.23718
R1934 CLK_div_3_mag_1.Q1.n7 CLK_div_3_mag_1.Q1 1.12056
R1935 CLK_div_3_mag_1.Q1.n0 CLK_div_3_mag_1.Q1 0.976034
R1936 Vdiv108.n8 Vdiv108.t4 36.935
R1937 Vdiv108.n6 Vdiv108.t6 31.528
R1938 Vdiv108.n8 Vdiv108.t3 18.1962
R1939 Vdiv108.n6 Vdiv108.t5 15.3826
R1940 Vdiv108.n4 Vdiv108.n1 7.09905
R1941 Vdiv108.n7 Vdiv108.n6 6.86134
R1942 Vdiv108.n10 Vdiv108.n9 5.01109
R1943 Vdiv108.n4 Vdiv108.n3 3.25085
R1944 Vdiv108.n11 Vdiv108.n5 2.36461
R1945 Vdiv108 Vdiv108.n0 2.27595
R1946 Vdiv108.n3 Vdiv108.t1 2.2755
R1947 Vdiv108.n3 Vdiv108.n2 2.2755
R1948 Vdiv108.n9 Vdiv108.n8 2.13398
R1949 Vdiv108.n11 Vdiv108.n10 1.47724
R1950 Vdiv108.n10 Vdiv108.n7 1.12725
R1951 Vdiv108 Vdiv108.n11 1.02714
R1952 Vdiv108.n5 Vdiv108.n4 0.0919062
R1953 Vdiv108.n7 Vdiv108 0.0857632
R1954 Vdiv108.n9 Vdiv108 0.0810725
R1955 Vdiv108.n5 Vdiv108 0.073625
R1956 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 37.1981
R1957 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 31.528
R1958 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 30.4613
R1959 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 24.7562
R1960 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 17.6611
R1961 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 15.3826
R1962 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 12.0856
R1963 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 9.86714
R1964 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K 6.09789
R1965 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 2.99416
R1966 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 2.2755
R1967 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 2.2755
R1968 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 2.2505
R1969 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 CLK_div_3_mag_0.JK_FF_mag_1.K 2.24173
R1970 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 1.93771
R1971 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n3 1.81589
R1972 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n2 1.43706
R1973 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.K.n1 0.281955
R1974 CLK_div_3_mag_1.Q0.n3 CLK_div_3_mag_1.Q0.t6 36.935
R1975 CLK_div_3_mag_1.Q0.n4 CLK_div_3_mag_1.Q0.t4 31.4332
R1976 CLK_div_3_mag_1.Q0.n2 CLK_div_3_mag_1.Q0.t3 29.8635
R1977 CLK_div_3_mag_1.Q0.n2 CLK_div_3_mag_1.Q0.t7 27.7543
R1978 CLK_div_3_mag_1.Q0.n3 CLK_div_3_mag_1.Q0.t5 18.1962
R1979 CLK_div_3_mag_1.Q0.n4 CLK_div_3_mag_1.Q0.t8 15.3826
R1980 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.t0 7.09905
R1981 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n4 6.86134
R1982 CLK_div_3_mag_1.Q0.n5 CLK_div_3_mag_1.Q0 5.0096
R1983 CLK_div_3_mag_1.Q0.n6 CLK_div_3_mag_1.Q0 3.41823
R1984 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n1 3.25226
R1985 CLK_div_3_mag_1.Q0.n1 CLK_div_3_mag_1.Q0.t1 2.2755
R1986 CLK_div_3_mag_1.Q0.n1 CLK_div_3_mag_1.Q0.n0 2.2755
R1987 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n6 2.2505
R1988 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n3 2.13479
R1989 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.Q0.n2 1.7371
R1990 CLK_div_3_mag_1.Q0.n6 CLK_div_3_mag_1.Q0.n5 1.50498
R1991 CLK_div_3_mag_1.Q0.n5 CLK_div_3_mag_1.Q0 1.12056
R1992 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 37.1984
R1993 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_3_mag_1.JK_FF_mag_1.K.t7 31.4332
R1994 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_3_mag_1.JK_FF_mag_1.K.t2 30.5184
R1995 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 CLK_div_3_mag_1.JK_FF_mag_1.K.t3 24.7029
R1996 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 17.6618
R1997 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 15.3826
R1998 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K 12.0839
R1999 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 9.86691
R2000 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_3_mag_1.JK_FF_mag_1.K 6.09789
R2001 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 2.99416
R2002 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_3_mag_1.JK_FF_mag_1.K.t0 2.2755
R2003 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 CLK_div_3_mag_1.JK_FF_mag_1.K.n1 2.2755
R2004 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 2.2505
R2005 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 CLK_div_3_mag_1.JK_FF_mag_1.K 2.24134
R2006 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 1.93723
R2007 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n3 1.81224
R2008 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n5 1.43718
R2009 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K.n7 0.4325
C0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q0 7.24e-19
C1 CLK_div_3_mag_2.JK_FF_mag_1.QB a_16712_1355# 0.0112f
C2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_14259_1355# 0.011f
C3 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C4 a_12004_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0731f
C5 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_18564_1311# 0.0203f
C6 a_18853_4654# JK_FF_mag_0.QB 0.0114f
C7 JK_FF_mag_1.Q JK_FF_mag_0.nand3_mag_1.OUT 6.64e-19
C8 CLK_div_3_mag_0.JK_FF_mag_1.K a_11929_2535# 0.00168f
C9 JK_FF_mag_1.Q CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00528f
C10 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C11 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VDD 0.996f
C12 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C13 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_1.K 0.00205f
C14 a_7853_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C15 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C16 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C17 a_19007_3557# JK_FF_mag_0.QB 0.0811f
C18 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1f
C19 a_18410_214# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C20 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C21 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.312f
C22 a_9355_4102# CLK_div_3_mag_0.Q1 0.069f
C23 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.QB 0.198f
C24 VDD a_13541_258# 3.14e-19
C25 a_7732_2691# CLK_div_3_mag_0.JK_FF_mag_1.QB 2.51e-19
C26 RST a_14829_214# 0.00212f
C27 a_12372_4102# VDD 3.73e-19
C28 CLK_div_3_mag_0.Q1 a_8221_5199# 0.0102f
C29 a_10680_4102# CLK_div_3_mag_0.Q0 2.79e-20
C30 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 9.52e-19
C31 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.Q0 7.24e-19
C32 CLK_div_3_mag_2.JK_FF_mag_1.QB a_15547_1311# 1.86e-20
C33 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C34 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_13695_1355# 0.00118f
C35 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C36 a_11440_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 9.1e-19
C37 a_15299_3554# VDD 3.14e-19
C38 a_18289_4654# JK_FF_mag_0.QB 2.96e-19
C39 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_18404_1311# 0.0732f
C40 JK_FF_mag_1.CLK VDD 1.42f
C41 CLK_div_3_mag_0.JK_FF_mag_1.K a_8705_2455# 3.16e-19
C42 a_8417_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C43 CLK_div_3_mag_2.JK_FF_mag_1.K a_18564_1311# 8.64e-19
C44 a_7289_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C45 RST CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.166f
C46 a_18443_3557# JK_FF_mag_0.QB 0.00964f
C47 JK_FF_mag_0.QB Vdiv108 1.94f
C48 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_3.IN1 5.32e-21
C49 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_7732_2691# 0.132f
C50 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_17840_1355# 0.0202f
C51 a_12158_1312# CLK_div_3_mag_1.JK_FF_mag_1.K 8.64e-19
C52 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.Q0 0.0635f
C53 VDD a_12164_215# 0.0132f
C54 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT a_8227_4102# 0.00378f
C55 a_15393_214# a_15553_214# 0.0504f
C56 a_11808_4102# VDD 3.14e-19
C57 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.Q1 0.0636f
C58 JK_FF_mag_1.CLK JK_FF_mag_1.nand3_mag_0.OUT 0.267f
C59 CLK_div_3_mag_0.Q1 a_7657_5199# 0.00789f
C60 RST a_14669_214# 0.00203f
C61 CLK_div_3_mag_2.JK_FF_mag_1.QB a_15387_1311# 1.41e-20
C62 VDD CLK_div_3_mag_2.Q0 1.34f
C63 a_11280_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C64 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK 5.57e-19
C65 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT a_17840_1355# 0.00378f
C66 a_11238_5199# VDD 2.21e-19
C67 a_7853_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C68 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C69 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C70 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C71 JK_FF_mag_0.nand3_mag_2.OUT VDD 0.748f
C72 a_17879_3513# JK_FF_mag_0.QB 0.00696f
C73 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_11434_1356# 0.0697f
C74 RST CLK_div_3_mag_2.or_2_mag_0.IN2 9.19e-19
C75 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C76 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C77 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT a_17276_1355# 4.52e-20
C78 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK 0.471f
C79 VDD a_12004_215# 0.00888f
C80 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C81 a_11244_4102# VDD 3.14e-19
C82 RST a_14105_258# 0.00121f
C83 CLK_div_3_mag_0.Q1 a_7497_5199# 0.00335f
C84 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_11434_1356# 5.01e-20
C85 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C86 JK_FF_mag_1.nand3_mag_2.OUT RST 0.0498f
C87 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C88 a_14575_3510# VDD 2.21e-19
C89 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.352f
C90 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 7.02e-21
C91 JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.399f
C92 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C93 RST a_8263_215# 0.00204f
C94 CLK a_15111_2454# 0.0103f
C95 a_10674_5199# VDD 0.00305f
C96 a_13695_1355# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C97 VDD a_8987_215# 0.00305f
C98 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT RST 0.277f
C99 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 a_10870_1356# 0.0059f
C100 a_17719_3513# JK_FF_mag_0.QB 0.00695f
C101 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.231f
C102 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 1.99e-19
C103 a_14017_4607# CLK_div_3_mag_0.Q0 1.07e-20
C104 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.656f
C105 a_17122_258# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C106 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 7.02e-21
C107 VDD a_11440_215# 0.0012f
C108 RST CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.135f
C109 JK_FF_mag_1.Q JK_FF_mag_0.nand3_mag_1.IN1 9.71e-20
C110 RST a_13541_258# 0.00114f
C111 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C112 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VDD 0.469f
C113 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C114 a_10680_4102# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00392f
C115 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 0.321f
C116 a_15863_3554# JK_FF_mag_1.QB 0.0811f
C117 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C118 a_15299_3554# RST 0.00137f
C119 a_10514_5199# VDD 0.00743f
C120 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C121 JK_FF_mag_1.CLK RST 7.64e-19
C122 a_11398_5199# RST 0.00103f
C123 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C124 a_13857_4607# CLK_div_3_mag_0.Q0 1.37e-20
C125 a_17879_3513# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 1.8e-21
C126 VDD a_11280_215# 9.82e-19
C127 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C128 RST a_12164_215# 0.00218f
C129 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.198f
C130 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.K 0.0613f
C131 VDD CLK_div_3_mag_1.JK_FF_mag_1.K 2.53f
C132 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 8.58e-20
C133 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C134 a_10956_3003# VDD 5.92e-19
C135 a_17719_3513# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 1.8e-21
C136 a_13851_3510# VDD 0.00108f
C137 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 8.16e-20
C138 RST CLK_div_3_mag_2.Q0 0.129f
C139 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.002f
C140 JK_FF_mag_1.CLK JK_FF_mag_1.nand2_mag_1.IN2 1.48e-20
C141 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN a_14138_2690# 0.132f
C142 a_14735_3510# RST 0.00206f
C143 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C144 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 8.58e-20
C145 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C146 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C147 a_11238_5199# RST 0.00119f
C148 JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 1.08e-20
C149 a_8263_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C150 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 2.81e-20
C151 JK_FF_mag_0.nand3_mag_2.OUT RST 0.082f
C152 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C153 VDD a_10716_259# 0.00149f
C154 a_14669_214# a_14829_214# 0.0504f
C155 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_12526_5199# 0.00372f
C156 RST a_12004_215# 0.00218f
C157 VDD a_15111_2454# 5.92e-19
C158 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 4.44e-20
C159 a_11244_4102# RST 2.95e-19
C160 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C161 a_7732_2691# VDD 0.165f
C162 a_14575_3510# RST 0.00103f
C163 JK_FF_mag_1.QB CLK 9.53e-20
C164 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_12372_4102# 4.94e-20
C165 a_14669_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C166 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.768f
C167 JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_0.Q0 0.00444f
C168 a_10674_5199# RST 0.00218f
C169 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.Q 0.0635f
C170 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.Q1 0.104f
C171 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C172 a_10680_4102# CLK_div_3_mag_0.JK_FF_mag_1.QB 1.41e-20
C173 RST a_8987_215# 0.00218f
C174 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK 0.362f
C175 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN JK_FF_mag_1.CLK 0.131f
C176 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C177 VDD a_10152_259# 0.00149f
C178 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.213f
C179 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 a_11962_5199# 0.069f
C180 RST a_11440_215# 0.00187f
C181 VDD a_14138_2690# 0.165f
C182 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.or_2_mag_0.IN2 1.82e-19
C183 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C184 a_8263_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C185 a_15553_214# CLK_div_3_mag_2.Q0 0.00335f
C186 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN RST 0.00146f
C187 a_9355_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C188 a_11398_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C189 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C190 CLK_div_3_mag_2.JK_FF_mag_1.K a_15387_1311# 0.00392f
C191 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.175f
C192 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.Q0 3.09e-19
C193 a_10514_5199# RST 0.00218f
C194 JK_FF_mag_1.Q JK_FF_mag_0.nand2_mag_3.IN1 0.421f
C195 a_10520_4102# CLK_div_3_mag_0.JK_FF_mag_1.QB 1.86e-20
C196 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C197 CLK_div_3_mag_0.JK_FF_mag_1.QB a_8381_5199# 0.00696f
C198 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.657f
C199 a_8981_1312# CLK_div_3_mag_1.JK_FF_mag_1.K 0.00392f
C200 a_7699_259# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C201 a_17155_3513# CLK_div_3_mag_2.JK_FF_mag_1.K 2.59e-19
C202 RST a_11280_215# 0.00228f
C203 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_17122_258# 0.069f
C204 a_11808_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C205 RST CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 0.0581f
C206 VDD a_11929_2535# 0.165f
C207 RST CLK_div_3_mag_1.JK_FF_mag_1.K 0.445f
C208 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C209 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C210 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C211 a_15393_214# CLK_div_3_mag_2.Q0 0.00789f
C212 a_10956_3003# RST 3.11e-19
C213 a_8791_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C214 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_1.QB 2.81e-20
C215 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C216 a_8987_215# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C217 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C218 RST CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.0547f
C219 CLK_div_3_mag_2.JK_FF_mag_1.K a_14823_1355# 1.75e-19
C220 a_7657_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C221 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_11998_1312# 0.00119f
C222 a_18289_4654# JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C223 a_9355_4102# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0112f
C224 JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.or_2_mag_0.IN2 9.24e-19
C225 a_17725_4654# VDD 3.14e-19
C226 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C227 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.Q0 0.0175f
C228 a_8945_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C229 CLK_div_3_mag_0.JK_FF_mag_1.QB a_8221_5199# 0.00695f
C230 a_8417_1356# CLK_div_3_mag_1.JK_FF_mag_1.K 1.75e-19
C231 a_18443_3557# JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C232 JK_FF_mag_0.nand3_mag_1.OUT Vdiv108 0.0343f
C233 a_8987_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C234 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C235 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_16558_258# 0.00372f
C236 RST a_10716_259# 0.00164f
C237 JK_FF_mag_1.QB VDD 0.916f
C238 a_16995_3513# CLK_div_3_mag_2.JK_FF_mag_1.K 2.59e-19
C239 a_11244_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C240 VDD a_8705_2455# 5.92e-19
C241 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C242 RST a_15111_2454# 7.58e-19
C243 a_14829_214# CLK_div_3_mag_2.Q0 0.0102f
C244 VDD CLK_div_3_mag_2.JK_FF_mag_1.QB 0.876f
C245 a_8227_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.43e-19
C246 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.0948f
C247 CLK_div_3_mag_2.JK_FF_mag_1.K a_14259_1355# 2.96e-19
C248 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 7.35e-19
C249 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_11434_1356# 1.43e-19
C250 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C251 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C252 CLK_div_3_mag_0.JK_FF_mag_1.K JK_FF_mag_1.nand2_mag_3.IN1 2.06e-19
C253 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C254 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.Q0 0.00335f
C255 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.175f
C256 a_7853_1356# CLK_div_3_mag_1.JK_FF_mag_1.K 2.96e-19
C257 a_17879_3513# JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C258 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_1.K 0.00384f
C259 JK_FF_mag_1.Q Vdiv108 0.158f
C260 RST a_10152_259# 0.00114f
C261 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C262 JK_FF_mag_1.CLK CLK_div_3_mag_2.or_2_mag_0.IN2 4.26e-19
C263 a_14669_214# CLK_div_3_mag_2.Q0 0.0101f
C264 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C265 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C266 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK 0.00481f
C267 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 0.0881f
C268 a_17846_214# CLK_div_3_mag_2.JK_FF_mag_1.QB 0.00695f
C269 CLK_div_3_mag_1.Q0 a_7699_259# 0.00859f
C270 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_1.K 0.00542f
C271 a_8987_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C272 CLK_div_3_mag_2.JK_FF_mag_1.K a_13695_1355# 0.012f
C273 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.CLK 0.235f
C274 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_10870_1356# 0.011f
C275 a_17001_4610# VDD 0.00514f
C276 a_8227_4102# CLK_div_3_mag_0.JK_FF_mag_1.QB 3.33e-19
C277 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C278 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 7.24e-19
C279 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.or_2_mag_0.IN2 0.0655f
C280 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_9509_5199# 0.00372f
C281 a_7289_1356# CLK_div_3_mag_1.JK_FF_mag_1.K 0.012f
C282 a_17719_3513# JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C283 RST CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.0232f
C284 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT CLK 0.298f
C285 a_7663_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0732f
C286 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VDD 0.647f
C287 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C288 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.198f
C289 a_11398_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C290 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.Q1 0.0138f
C291 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_7732_2691# 3.25e-19
C292 a_7732_2691# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C293 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.359f
C294 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C295 a_14105_258# CLK_div_3_mag_2.Q0 0.00859f
C296 a_7135_259# CLK_div_3_mag_1.JK_FF_mag_1.K 0.0811f
C297 JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.Q0 1.22e-19
C298 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C299 JK_FF_mag_0.QB VDD 0.982f
C300 JK_FF_mag_1.nand3_mag_2.OUT a_14735_3510# 2.88e-20
C301 a_17686_214# CLK_div_3_mag_2.JK_FF_mag_1.QB 0.00696f
C302 a_15393_214# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C303 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_14823_1355# 0.0202f
C304 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.107f
C305 JK_FF_mag_0.nand3_mag_0.OUT a_17725_4654# 0.00378f
C306 CLK_div_3_mag_2.JK_FF_mag_1.K a_12158_1312# 1.01e-20
C307 a_11808_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C308 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 a_10306_1356# 0.00118f
C309 a_15709_4651# VDD 3.56e-19
C310 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 a_8945_5199# 0.069f
C311 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.or_2_mag_0.IN2 0.0655f
C312 a_17725_4654# RST 2.59e-19
C313 a_7663_4102# CLK_div_3_mag_0.Q1 2.79e-20
C314 a_17155_3513# JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C315 a_7503_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C316 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C317 JK_FF_mag_1.QB JK_FF_mag_0.nand3_mag_0.OUT 2.4e-20
C318 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0635f
C319 CLK_div_3_mag_0.JK_FF_mag_1.K JK_FF_mag_1.Q 3.16e-21
C320 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_1.K 0.69f
C321 a_11238_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C322 a_18570_214# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C323 CLK_div_3_mag_2.JK_FF_mag_1.K CLK 2.11f
C324 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1f
C325 JK_FF_mag_1.QB RST 0.162f
C326 RST a_8705_2455# 4.71e-19
C327 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT 2.29e-20
C328 a_13541_258# CLK_div_3_mag_2.Q0 0.0157f
C329 a_18289_4654# JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C330 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C331 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C332 JK_FF_mag_1.nand3_mag_2.OUT a_14575_3510# 9.1e-19
C333 a_17122_258# CLK_div_3_mag_2.JK_FF_mag_1.QB 0.00964f
C334 a_18404_1311# a_18564_1311# 0.0504f
C335 RST CLK_div_3_mag_2.JK_FF_mag_1.QB 0.596f
C336 CLK_div_3_mag_2.JK_FF_mag_1.K a_11998_1312# 6.09e-21
C337 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT a_14259_1355# 4.52e-20
C338 JK_FF_mag_0.nand3_mag_0.OUT a_17161_4610# 0.0732f
C339 JK_FF_mag_0.nand3_mag_1.IN1 Vdiv108 0.00335f
C340 a_11244_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C341 a_15145_4651# VDD 3.14e-19
C342 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.392f
C343 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 7.3e-19
C344 a_17161_4610# RST 7.58e-19
C345 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C346 JK_FF_mag_1.CLK CLK_div_3_mag_2.Q0 9.37e-19
C347 a_16995_3513# JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C348 a_17155_3513# JK_FF_mag_1.Q 0.00208f
C349 a_7503_4102# a_7663_4102# 0.0504f
C350 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_1.IN2 0.0592f
C351 a_10520_4102# VDD 2.21e-19
C352 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 1f
C353 a_10674_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C354 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.00205f
C355 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C356 a_18410_214# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C357 a_11238_5199# a_11398_5199# 0.0504f
C358 VDD a_8381_5199# 9.82e-19
C359 a_12164_215# CLK_div_3_mag_2.Q0 1.27e-20
C360 CLK_div_3_mag_1.Q0 a_7663_4102# 3.49e-20
C361 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.Q0 0.0655f
C362 a_16558_258# CLK_div_3_mag_2.JK_FF_mag_1.QB 0.0811f
C363 JK_FF_mag_1.nand3_mag_2.OUT a_14011_3510# 0.0731f
C364 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C365 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN a_11929_2535# 0.132f
C366 a_17879_3513# JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C367 JK_FF_mag_0.nand3_mag_0.OUT a_17001_4610# 0.0203f
C368 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.653f
C369 a_14581_4651# VDD 3.14e-19
C370 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C371 JK_FF_mag_1.nand3_mag_1.OUT CLK 0.00156f
C372 JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.657f
C373 CLK_div_3_mag_1.Q0 a_8423_215# 0.0102f
C374 a_17001_4610# RST 9.1e-19
C375 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C376 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C377 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_8705_2455# 0.069f
C378 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C379 a_12004_215# a_12164_215# 0.0504f
C380 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.161f
C381 a_16995_3513# JK_FF_mag_1.Q 0.00174f
C382 a_9355_4102# VDD 3.56e-19
C383 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.Q0 0.0285f
C384 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11962_5199# 0.0036f
C385 a_17846_214# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C386 a_10514_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C387 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT RST 0.00494f
C388 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.or_2_mag_0.IN2 5.32e-19
C389 VDD a_8221_5199# 0.0012f
C390 a_12004_215# CLK_div_3_mag_2.Q0 1.01e-20
C391 JK_FF_mag_1.nand3_mag_0.OUT a_14581_4651# 0.00378f
C392 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C393 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_0.OUT 0.343f
C394 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C395 JK_FF_mag_1.nand3_mag_2.OUT a_13851_3510# 0.0202f
C396 JK_FF_mag_0.QB RST 0.0999f
C397 a_8263_215# CLK_div_3_mag_1.JK_FF_mag_1.K 0.00696f
C398 a_14105_258# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C399 JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 7.72e-21
C400 CLK_div_3_mag_2.or_2_mag_0.IN2 a_15111_2454# 7.48e-20
C401 JK_FF_mag_1.nand2_mag_3.IN1 CLK 7.92e-20
C402 a_14575_3510# a_14735_3510# 0.0504f
C403 a_15709_4651# RST 5.97e-19
C404 VDD CLK_div_3_mag_2.JK_FF_mag_1.K 2.32f
C405 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_1.CLK 1e-19
C406 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C407 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.313f
C408 a_14011_3510# JK_FF_mag_1.CLK 0.00233f
C409 a_18853_4654# JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C410 a_15863_3554# JK_FF_mag_1.Q 0.0157f
C411 a_8791_4102# VDD 3.14e-19
C412 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C413 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK 0.00302f
C414 a_17686_214# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C415 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.395f
C416 a_10680_4102# RST 0.0012f
C417 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C418 VDD a_7657_5199# 0.00888f
C419 JK_FF_mag_1.nand3_mag_0.OUT a_14017_4607# 0.0732f
C420 RST CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.316f
C421 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 1.11e-20
C422 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C423 JK_FF_mag_1.nand2_mag_1.IN2 a_15709_4651# 0.00372f
C424 a_14011_3510# CLK_div_3_mag_2.Q0 4.06e-19
C425 JK_FF_mag_1.CLK CLK_div_3_mag_1.JK_FF_mag_1.K 0.00195f
C426 a_13857_4607# VDD 0.00484f
C427 CLK_div_3_mag_2.or_2_mag_0.IN2 a_14138_2690# 8.64e-19
C428 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.394f
C429 a_15145_4651# RST 5.97e-19
C430 a_13851_3510# JK_FF_mag_1.CLK 0.00211f
C431 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 RST 0.00239f
C432 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.00586f
C433 a_18289_4654# JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C434 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_1.QB 4.28e-19
C435 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C436 a_8227_4102# VDD 3.14e-19
C437 JK_FF_mag_0.nand3_mag_1.OUT CLK 3.92e-21
C438 a_17122_258# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C439 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK 0.0983f
C440 a_10520_4102# RST 0.00163f
C441 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C442 RST CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.313f
C443 VDD a_7497_5199# 0.0132f
C444 a_18443_3557# JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C445 JK_FF_mag_0.nand2_mag_3.IN1 Vdiv108 0.0168f
C446 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 6.62e-20
C447 JK_FF_mag_1.nand3_mag_0.OUT a_13857_4607# 0.0203f
C448 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C449 RST a_8381_5199# 0.00135f
C450 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.0948f
C451 JK_FF_mag_1.nand3_mag_1.OUT VDD 1f
C452 CLK_div_3_mag_2.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K 0.0437f
C453 a_18853_4654# JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C454 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C455 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.00761f
C456 a_10306_1356# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C457 JK_FF_mag_1.nand2_mag_1.IN2 a_15145_4651# 0.069f
C458 a_13851_3510# CLK_div_3_mag_2.Q0 2.99e-19
C459 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 3.81e-19
C460 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C461 a_19007_3557# JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C462 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.Q0 0.0175f
C463 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0881f
C464 a_14105_258# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C465 JK_FF_mag_1.nand3_mag_1.IN1 RST 0.189f
C466 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C467 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C468 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 3.76e-19
C469 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.53e-20
C470 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C471 JK_FF_mag_1.Q CLK 0.014f
C472 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C473 CLK_div_3_mag_1.Q0 a_9147_215# 0.00335f
C474 a_10514_5199# a_10674_5199# 0.0504f
C475 a_9355_4102# RST 0.00208f
C476 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q1 0.362f
C477 a_18853_4654# Vdiv108 0.069f
C478 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 7.3e-19
C479 RST a_8221_5199# 8.64e-19
C480 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C481 JK_FF_mag_1.nand2_mag_3.IN1 VDD 1.3f
C482 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1 1.12e-19
C483 a_19007_3557# Vdiv108 0.0157f
C484 JK_FF_mag_1.CLK a_14138_2690# 3.27e-19
C485 JK_FF_mag_1.QB CLK_div_3_mag_2.or_2_mag_0.IN2 9.3e-20
C486 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C487 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C488 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C489 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 8.58e-20
C490 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 2.34e-19
C491 a_18443_3557# JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C492 JK_FF_mag_0.nand2_mag_4.IN2 Vdiv108 0.0635f
C493 a_13541_258# CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C494 RST CLK_div_3_mag_2.JK_FF_mag_1.K 0.442f
C495 a_11280_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C496 a_11280_215# a_11440_215# 0.0504f
C497 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand2_mag_3.IN1 0.0893f
C498 JK_FF_mag_1.Q CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 3.37e-19
C499 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 8.58e-20
C500 a_8791_4102# RST 8.99e-19
C501 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 a_17276_1355# 0.069f
C502 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C503 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.QB 0.103f
C504 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 RST 0.0592f
C505 a_10956_3003# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 4.98e-20
C506 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0169f
C507 a_7503_4102# CLK_div_3_mag_0.JK_FF_mag_1.K 8.64e-19
C508 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 4.28e-19
C509 a_7663_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.00119f
C510 CLK_div_3_mag_2.Q0 a_14138_2690# 0.0134f
C511 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_1.K 0.00559f
C512 a_18443_3557# Vdiv108 0.00859f
C513 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.K 0.027f
C514 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 1.8e-21
C515 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.QB 0.343f
C516 a_10956_3003# CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN 0.069f
C517 JK_FF_mag_0.nand3_mag_1.OUT VDD 0.997f
C518 JK_FF_mag_1.Q CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 9.01e-22
C519 VDD CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.465f
C520 a_13851_3510# a_14011_3510# 0.0504f
C521 a_9141_1312# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C522 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C523 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.0625f
C524 CLK_div_3_mag_0.Q0 CLK_div_3_mag_1.JK_FF_mag_1.QB 4.1e-21
C525 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C526 a_8227_4102# RST 1.21e-19
C527 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 a_16712_1355# 0.00372f
C528 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_2.Q0 0.0635f
C529 a_17155_3513# JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C530 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C531 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C532 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.Q0 2.37f
C533 a_10956_3003# CLK_div_3_mag_1.JK_FF_mag_1.K 3.16e-19
C534 a_15299_3554# JK_FF_mag_1.QB 0.00964f
C535 JK_FF_mag_1.nand3_mag_1.OUT RST 0.262f
C536 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_9355_4102# 0.00372f
C537 a_17879_3513# Vdiv108 0.0101f
C538 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.Q1 1.94f
C539 JK_FF_mag_1.CLK JK_FF_mag_1.QB 0.307f
C540 JK_FF_mag_0.nand3_mag_1.IN1 CLK 7.07e-21
C541 a_7663_4102# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00392f
C542 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.99e-20
C543 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.08f
C544 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.Q0 0.107f
C545 JK_FF_mag_1.Q VDD 2.25f
C546 a_8981_1312# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C547 a_15863_3554# JK_FF_mag_1.nand2_mag_4.IN2 0.00372f
C548 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00698f
C549 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C550 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.Q 7.24e-19
C551 a_12526_5199# CLK_div_3_mag_0.Q0 0.0157f
C552 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C553 a_14735_3510# JK_FF_mag_1.QB 0.00696f
C554 a_7732_2691# CLK_div_3_mag_1.JK_FF_mag_1.K 0.00168f
C555 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 a_8791_4102# 0.069f
C556 JK_FF_mag_1.nand2_mag_3.IN1 RST 0.0611f
C557 a_17719_3513# Vdiv108 0.0102f
C558 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C559 a_9509_5199# CLK_div_3_mag_0.Q1 0.0157f
C560 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C561 a_8417_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C562 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN a_8227_4102# 5.01e-20
C563 RST CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.311f
C564 CLK_div_3_mag_1.Q0 CLK_div_3_mag_0.JK_FF_mag_1.QB 4.1e-21
C565 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.36f
C566 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 8.31e-21
C567 a_17719_3513# a_17879_3513# 0.0504f
C568 a_14575_3510# JK_FF_mag_1.QB 0.00695f
C569 a_11962_5199# CLK_div_3_mag_0.Q0 0.00859f
C570 a_17155_3513# Vdiv108 0.00789f
C571 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN a_11929_2535# 3.25e-19
C572 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT 0.803f
C573 a_8945_5199# CLK_div_3_mag_0.Q1 0.00859f
C574 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C575 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_14138_2690# 1.4e-19
C576 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 0.209f
C577 a_14829_214# CLK_div_3_mag_2.JK_FF_mag_1.K 0.00695f
C578 JK_FF_mag_0.nand3_mag_1.OUT RST 0.254f
C579 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C580 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK 0.235f
C581 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_11434_1356# 0.0202f
C582 RST CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00746f
C583 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C584 a_18564_1311# CLK 0.0101f
C585 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.Q0 5.76e-20
C586 VDD a_7699_259# 3.14e-19
C587 JK_FF_mag_1.nand2_mag_4.IN2 CLK 2.59e-19
C588 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C589 JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.653f
C590 a_11929_2535# CLK_div_3_mag_1.JK_FF_mag_1.K 0.00263f
C591 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C592 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C593 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C594 a_16995_3513# Vdiv108 0.00335f
C595 a_15387_1311# a_15547_1311# 0.0504f
C596 JK_FF_mag_1.Q JK_FF_mag_0.nand3_mag_0.OUT 0.267f
C597 a_15553_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C598 JK_FF_mag_1.Q RST 0.164f
C599 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 RST 0.0143f
C600 a_14669_214# CLK_div_3_mag_2.JK_FF_mag_1.K 0.00696f
C601 a_12372_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C602 a_12004_215# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C603 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand3_mag_1.IN1 0.00163f
C604 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT a_10870_1356# 4.52e-20
C605 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 0.0725f
C606 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C607 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1f
C608 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT a_11244_4102# 0.00378f
C609 a_18404_1311# CLK 0.00939f
C610 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.QB 0.103f
C611 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_1.CLK 5.6e-20
C612 JK_FF_mag_0.nand2_mag_3.IN1 CLK 1.29e-19
C613 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.398f
C614 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.or_2_mag_0.IN2 0.00761f
C615 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00975f
C616 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0854f
C617 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.QB 0.175f
C618 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_18570_214# 0.0202f
C619 CLK_div_3_mag_1.or_2_mag_0.IN2 VDD 0.493f
C620 a_12526_5199# CLK_div_3_mag_0.JK_FF_mag_1.K 0.0811f
C621 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.Q 0.107f
C622 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C623 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.391f
C624 a_15393_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C625 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.231f
C626 a_14105_258# CLK_div_3_mag_2.JK_FF_mag_1.K 0.00964f
C627 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.0622f
C628 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_1.IN2 0.0592f
C629 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VDD 0.65f
C630 JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.K 6.21e-20
C631 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.QB 7.08e-20
C632 a_17840_1355# CLK 6.43e-21
C633 CLK_div_3_mag_0.or_2_mag_0.IN2 VDD 0.493f
C634 JK_FF_mag_1.CLK a_14581_4651# 6.43e-21
C635 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.35e-20
C636 JK_FF_mag_1.CLK JK_FF_mag_1.nand3_mag_1.IN1 9.71e-20
C637 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C638 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.74f
C639 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C640 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_18410_214# 0.0731f
C641 a_11962_5199# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00964f
C642 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT RST 0.0551f
C643 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.0718f
C644 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT CLK 0.235f
C645 VDD a_18564_1311# 6.01e-19
C646 a_14829_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C647 a_13541_258# CLK_div_3_mag_2.JK_FF_mag_1.K 0.0811f
C648 JK_FF_mag_0.nand2_mag_4.IN2 CLK 1.05e-20
C649 VDD CLK_div_3_mag_0.Q1 2.52f
C650 JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.391f
C651 CLK_div_3_mag_0.Q0 a_11998_1312# 3.49e-20
C652 a_7663_4102# VDD 2.65e-19
C653 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.K 3.28e-19
C654 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.K 0.0718f
C655 a_17276_1355# CLK 6.06e-21
C656 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C657 a_14735_3510# JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C658 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.122f
C659 JK_FF_mag_1.CLK a_14017_4607# 0.00939f
C660 CLK_div_3_mag_0.Q1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 1.45e-19
C661 RST a_7699_259# 0.00122f
C662 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C663 a_16995_3513# a_17155_3513# 0.0504f
C664 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C665 JK_FF_mag_0.nand3_mag_1.IN1 RST 0.157f
C666 CLK_div_3_mag_0.Q0 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 3.09e-19
C667 VDD a_8423_215# 2.21e-19
C668 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_17846_214# 9.1e-19
C669 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.653f
C670 Vdiv108 CLK 1.56e-19
C671 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK 0.0215f
C672 VDD a_18404_1311# 2.65e-19
C673 a_14669_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C674 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C675 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00542f
C676 a_10716_259# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C677 a_14017_4607# CLK_div_3_mag_2.Q0 1.98e-21
C678 a_7503_4102# VDD 5.99e-19
C679 JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.31f
C680 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.Q0 2.37f
C681 CLK_div_3_mag_0.JK_FF_mag_1.QB CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C682 a_16712_1355# CLK 9.45e-19
C683 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_8705_2455# 4.98e-20
C684 JK_FF_mag_1.CLK a_13857_4607# 0.0101f
C685 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.337f
C686 CLK_div_3_mag_1.Q0 VDD 1.27f
C687 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 6.02e-20
C688 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C689 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.or_2_mag_0.IN2 4.52e-20
C690 RST CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00355f
C691 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C692 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT a_17686_214# 2.88e-20
C693 JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.K 6.19e-20
C694 CLK_div_3_mag_1.or_2_mag_0.IN2 RST 8.93e-19
C695 VDD a_17840_1355# 3.16e-19
C696 a_15299_3554# JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C697 a_14105_258# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C698 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 6.62e-20
C699 RST CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.0239f
C700 JK_FF_mag_1.CLK JK_FF_mag_1.nand3_mag_1.OUT 6.64e-19
C701 a_18853_4654# VDD 3.56e-19
C702 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT RST 9.38e-19
C703 a_7699_259# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C704 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C705 VDD CLK_div_3_mag_0.Q0 1.33f
C706 a_15547_1311# CLK 0.0101f
C707 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C708 a_19007_3557# VDD 3.48e-19
C709 JK_FF_mag_1.Q CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 1.4e-20
C710 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C711 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C712 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C713 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.00166f
C714 JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.392f
C715 CLK_div_3_mag_1.JK_FF_mag_1.QB a_11998_1312# 0.00392f
C716 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.101f
C717 RST CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT 0.0545f
C718 JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.Q0 6.96e-19
C719 a_14735_3510# JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C720 VDD a_17276_1355# 3.16e-19
C721 a_15299_3554# JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C722 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 a_14259_1355# 0.069f
C723 JK_FF_mag_1.QB a_17161_4610# 1.08e-20
C724 JK_FF_mag_1.CLK JK_FF_mag_1.nand2_mag_3.IN1 0.419f
C725 a_18289_4654# VDD 3.14e-19
C726 CLK_div_3_mag_0.Q1 RST 0.273f
C727 JK_FF_mag_1.nand2_mag_4.IN2 RST 0.0235f
C728 a_8945_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C729 a_15387_1311# CLK 0.00939f
C730 a_7853_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C731 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.QB 4.75e-20
C732 a_18443_3557# VDD 3.14e-19
C733 Vdiv108 VDD 1.15f
C734 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C735 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.399f
C736 CLK_div_3_mag_1.or_2_mag_0.IN2 a_7853_1356# 4.9e-20
C737 JK_FF_mag_1.Q CLK_div_3_mag_2.or_2_mag_0.IN2 0.00549f
C738 a_9509_5199# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0811f
C739 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 0.124f
C740 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 7.35e-19
C741 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C742 CLK_div_3_mag_1.JK_FF_mag_1.QB a_11434_1356# 3.33e-19
C743 RST a_8423_215# 0.00212f
C744 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C745 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_15547_1311# 0.0203f
C746 VDD a_16712_1355# 3.57e-19
C747 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.166f
C748 a_14575_3510# JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C749 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 a_13695_1355# 0.00372f
C750 JK_FF_mag_1.nand3_mag_2.OUT JK_FF_mag_1.Q 0.338f
C751 JK_FF_mag_1.QB a_17001_4610# 1.38e-20
C752 VDD a_9147_215# 0.00743f
C753 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_1.IN2 8.16e-20
C754 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C755 CLK_div_3_mag_1.Q0 a_8981_1312# 2.79e-20
C756 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K 8.05e-19
C757 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.Q0 0.0343f
C758 a_7699_259# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C759 a_7289_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.00372f
C760 JK_FF_mag_0.nand2_mag_3.IN1 RST 0.00475f
C761 a_14823_1355# CLK 6.43e-21
C762 a_14735_3510# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 8.31e-21
C763 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C764 JK_FF_mag_0.QB a_17725_4654# 3.33e-19
C765 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.16f
C766 JK_FF_mag_1.CLK CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 1.73e-19
C767 CLK_div_3_mag_1.Q0 RST 0.139f
C768 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 0.69f
C769 a_8945_5199# CLK_div_3_mag_0.JK_FF_mag_1.QB 0.00964f
C770 a_8417_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C771 a_17001_4610# a_17161_4610# 0.0504f
C772 JK_FF_mag_1.QB JK_FF_mag_0.QB 4.17e-22
C773 a_7289_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 4.52e-20
C774 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C775 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_17840_1355# 0.0697f
C776 a_14011_3510# JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C777 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_15387_1311# 0.0732f
C778 VDD CLK_div_3_mag_1.JK_FF_mag_1.QB 0.878f
C779 VDD a_15547_1311# 2.21e-19
C780 a_12372_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C781 JK_FF_mag_1.QB a_15709_4651# 0.0114f
C782 a_7135_259# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 0.00372f
C783 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 1.76e-19
C784 a_15299_3554# JK_FF_mag_1.Q 0.00859f
C785 CLK_div_3_mag_2.Q0 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C786 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C787 JK_FF_mag_0.QB a_17161_4610# 0.00392f
C788 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C789 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 a_8381_5199# 8.64e-19
C790 a_17719_3513# VDD 2.21e-19
C791 RST CLK_div_3_mag_0.Q0 0.0457f
C792 JK_FF_mag_1.CLK JK_FF_mag_1.Q 0.161f
C793 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C794 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q1 0.0014f
C795 CLK_div_3_mag_0.JK_FF_mag_1.K VDD 2.66f
C796 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_1.CLK 2.14e-20
C797 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK 7.81e-19
C798 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.Q1 0.107f
C799 a_7853_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C800 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C801 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C802 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C803 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00169f
C804 RST CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.107f
C805 CLK_div_3_mag_1.JK_FF_mag_1.QB a_10306_1356# 0.0112f
C806 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.233f
C807 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C808 JK_FF_mag_0.nand2_mag_4.IN2 RST 3.69e-19
C809 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C810 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 a_17276_1355# 0.0059f
C811 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT a_14823_1355# 0.00378f
C812 a_13851_3510# JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C813 a_14011_3510# JK_FF_mag_1.nand2_mag_3.IN1 1.46e-19
C814 a_8423_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C815 JK_FF_mag_1.QB a_15145_4651# 2.96e-19
C816 a_10716_259# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.069f
C817 a_11808_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C818 RST a_17276_1355# 7.1e-19
C819 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 6.7e-19
C820 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.00169f
C821 JK_FF_mag_1.Q CLK_div_3_mag_2.Q0 0.00335f
C822 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C823 CLK_div_3_mag_2.JK_FF_mag_1.K a_14138_2690# 0.00168f
C824 a_14735_3510# JK_FF_mag_1.Q 0.0101f
C825 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C826 JK_FF_mag_0.nand3_mag_0.OUT Vdiv108 7.24e-19
C827 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand2_mag_1.IN2 0.00975f
C828 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 4.81e-22
C829 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C830 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.109f
C831 a_12526_5199# VDD 3.14e-19
C832 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 1.53e-19
C833 Vdiv108 RST 0.0434f
C834 VDD CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.01f
C835 RST CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.00536f
C836 CLK_div_3_mag_0.Q0 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 2.29e-20
C837 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_1.Q 0.235f
C838 CLK_div_3_mag_1.JK_FF_mag_1.QB a_9141_1312# 1.86e-20
C839 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C840 JK_FF_mag_1.nand3_mag_1.OUT a_15111_2454# 1.82e-21
C841 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.215f
C842 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.198f
C843 VDD a_14823_1355# 3.14e-19
C844 JK_FF_mag_1.QB a_14581_4651# 3.33e-19
C845 a_11244_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C846 a_10152_259# CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.00372f
C847 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_1.IN1 0.0383f
C848 RST a_16712_1355# 0.00154f
C849 RST a_9147_215# 0.00218f
C850 a_8791_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C851 CLK_div_3_mag_1.Q0 a_7289_1356# 0.069f
C852 a_10680_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C853 a_13695_1355# CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 4.94e-20
C854 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C855 a_14575_3510# JK_FF_mag_1.Q 0.0102f
C856 JK_FF_mag_1.Q JK_FF_mag_0.nand2_mag_1.IN2 1.48e-20
C857 a_16995_3513# VDD 0.00108f
C858 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C859 a_10674_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C860 a_11962_5199# VDD 3.14e-19
C861 CLK_div_3_mag_1.Q0 a_7135_259# 0.0157f
C862 a_17879_3513# RST 0.00154f
C863 a_8423_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C864 a_15553_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C865 a_11998_1312# a_12158_1312# 0.0504f
C866 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C867 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.Q0 0.209f
C868 CLK_div_3_mag_1.JK_FF_mag_1.QB a_8981_1312# 1.41e-20
C869 CLK_div_3_mag_0.JK_FF_mag_1.QB VDD 0.88f
C870 VDD a_14259_1355# 3.14e-19
C871 JK_FF_mag_1.QB a_14017_4607# 0.00392f
C872 RST CLK_div_3_mag_1.JK_FF_mag_1.QB 0.696f
C873 RST a_15547_1311# 0.00214f
C874 JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.K 5.25e-20
C875 a_8227_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.0697f
C876 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.399f
C877 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C878 a_10520_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C879 a_14011_3510# JK_FF_mag_1.Q 0.00789f
C880 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C881 CLK_div_3_mag_0.Q0 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C882 a_15863_3554# VDD 3.14e-19
C883 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.QB 3.28e-19
C884 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 3.67e-20
C885 a_17719_3513# RST 0.00177f
C886 a_15393_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C887 CLK_div_3_mag_0.JK_FF_mag_1.K RST 0.292f
C888 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VDD 0.415f
C889 CLK CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 6.28e-21
C890 a_9509_5199# VDD 0.00149f
C891 VDD a_13695_1355# 3.56e-19
C892 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C893 RST a_15387_1311# 0.00154f
C894 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN a_15111_2454# 0.069f
C895 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.121f
C896 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.IN1 0.00158f
C897 a_10520_4102# a_10680_4102# 0.0504f
C898 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C899 a_13851_3510# JK_FF_mag_1.Q 0.00335f
C900 a_9147_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C901 a_12164_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C902 JK_FF_mag_1.Q CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 6.27e-22
C903 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT CLK 0.272f
C904 a_17155_3513# RST 0.00251f
C905 a_18570_214# CLK 0.00117f
C906 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C907 a_14829_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C908 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.Q1 4.33e-19
C909 a_8381_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C910 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_1.OUT 0.25f
C911 RST CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.139f
C912 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 7.08e-20
C913 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 0.122f
C914 a_8945_5199# VDD 0.00149f
C915 VDD a_12158_1312# 5.99e-19
C916 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_1.K 3.03e-20
C917 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.109f
C918 RST a_14823_1355# 5.61e-19
C919 a_8263_215# a_8423_215# 0.0504f
C920 JK_FF_mag_1.Q a_15111_2454# 2.99e-19
C921 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN a_14138_2690# 3.25e-19
C922 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C923 a_11398_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C924 a_8263_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C925 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00559f
C926 a_12004_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C927 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_1.QB 4.75e-20
C928 CLK_div_3_mag_0.or_2_mag_0.IN2 a_11808_4102# 4.9e-20
C929 JK_FF_mag_1.nand2_mag_4.IN2 a_15299_3554# 0.069f
C930 JK_FF_mag_0.QB CLK_div_3_mag_2.JK_FF_mag_1.K 5.16e-20
C931 VDD CLK 2.42f
C932 a_16995_3513# RST 0.00266f
C933 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.802f
C934 a_18410_214# CLK 0.00164f
C935 a_14669_214# CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C936 a_8221_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C937 JK_FF_mag_1.CLK CLK_div_3_mag_0.Q1 2.53e-19
C938 JK_FF_mag_1.nand3_mag_1.IN1 a_15145_4651# 0.0059f
C939 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_3.IN1 0.28f
C940 CLK_div_3_mag_1.Q0 a_8263_215# 0.0101f
C941 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_18404_1311# 0.00119f
C942 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00205f
C943 a_9147_215# CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C944 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C945 VDD a_11998_1312# 2.65e-19
C946 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C947 CLK_div_3_mag_0.JK_FF_mag_1.QB RST 0.625f
C948 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.K 8.58e-20
C949 RST a_14259_1355# 5.02e-19
C950 JK_FF_mag_1.Q a_14138_2690# 0.00263f
C951 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C952 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.765f
C953 a_11238_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C954 a_11440_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0203f
C955 RST CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 0.00356f
C956 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 1.35e-20
C957 a_8791_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C958 VDD CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.416f
C959 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C960 a_15863_3554# RST 0.00203f
C961 a_7699_259# CLK_div_3_mag_1.JK_FF_mag_1.K 0.00964f
C962 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.122f
C963 JK_FF_mag_0.nand3_mag_1.OUT a_17725_4654# 0.0202f
C964 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 3.76e-19
C965 a_7657_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.5e-20
C966 a_11238_5199# CLK_div_3_mag_0.Q1 3.6e-22
C967 a_8221_5199# a_8381_5199# 0.0504f
C968 JK_FF_mag_1.nand3_mag_1.IN1 a_14581_4651# 0.0697f
C969 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C970 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_17840_1355# 1.43e-19
C971 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.Q0 0.0343f
C972 VDD a_11434_1356# 3.14e-19
C973 a_9509_5199# RST 0.00114f
C974 RST a_13695_1355# 5.02e-19
C975 JK_FF_mag_1.QB CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 4.37e-20
C976 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 a_11929_2535# 1.4e-19
C977 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C978 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 0.359f
C979 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 9.62e-20
C980 VDD a_18570_214# 0.0132f
C981 a_10674_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C982 a_18410_214# a_18570_214# 0.0504f
C983 a_11280_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C984 JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.QB 1.22e-19
C985 a_12372_4102# CLK_div_3_mag_0.Q0 0.069f
C986 a_8227_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0202f
C987 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_1.JK_FF_mag_1.K 9.62e-20
C988 JK_FF_mag_1.Q a_17725_4654# 6.43e-21
C989 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.0948f
C990 a_7497_5199# CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C991 a_10674_5199# CLK_div_3_mag_0.Q1 1.86e-20
C992 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 0.0725f
C993 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.or_2_mag_0.IN2 0.124f
C994 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_17276_1355# 0.011f
C995 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.K 6.15e-20
C996 JK_FF_mag_1.CLK CLK_div_3_mag_0.Q0 0.209f
C997 a_11398_5199# CLK_div_3_mag_0.Q0 0.0101f
C998 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand2_mag_3.IN1 0.00118f
C999 VDD a_10870_1356# 3.14e-19
C1000 CLK_div_3_mag_1.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 0.00761f
C1001 a_8945_5199# RST 5.68e-19
C1002 CLK_div_3_mag_0.Q1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 3.17e-19
C1003 JK_FF_mag_1.QB JK_FF_mag_1.Q 1.96f
C1004 RST a_12158_1312# 7.78e-19
C1005 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 0.198f
C1006 VDD a_18410_214# 0.00888f
C1007 a_10514_5199# CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C1008 JK_FF_mag_1.nand3_mag_1.OUT a_15145_4651# 4.52e-20
C1009 a_10716_259# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C1010 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_10870_1356# 0.069f
C1011 JK_FF_mag_1.nand2_mag_3.IN1 a_15709_4651# 0.00118f
C1012 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1.26e-19
C1013 a_9355_4102# CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C1014 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q1 0.305f
C1015 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 0.359f
C1016 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_1.QB 0.0576f
C1017 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 CLK 0.013f
C1018 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN 3.34e-19
C1019 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_1.K 0.00586f
C1020 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C1021 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.397f
C1022 a_10514_5199# CLK_div_3_mag_0.Q1 2.55e-20
C1023 JK_FF_mag_1.Q a_17161_4610# 0.00939f
C1024 RST CLK 0.132f
C1025 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 0.36f
C1026 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0843f
C1027 a_10956_3003# CLK_div_3_mag_0.or_2_mag_0.IN2 7.48e-20
C1028 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00166f
C1029 JK_FF_mag_1.nand3_mag_0.OUT VDD 0.742f
C1030 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 a_16712_1355# 0.00118f
C1031 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT CLK_div_3_mag_2.Q0 0.338f
C1032 a_11238_5199# CLK_div_3_mag_0.Q0 0.0102f
C1033 VDD a_10306_1356# 3.56e-19
C1034 RST a_11998_1312# 6.43e-19
C1035 CLK_div_3_mag_1.or_2_mag_0.IN2 a_7732_2691# 8.64e-19
C1036 CLK_div_3_mag_1.Q0 a_8987_215# 0.00789f
C1037 VDD a_17846_214# 0.0012f
C1038 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_12158_1312# 0.0203f
C1039 JK_FF_mag_1.nand3_mag_1.OUT a_14581_4651# 0.0202f
C1040 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 a_10306_1356# 0.00372f
C1041 CLK_div_3_mag_0.Q1 CLK_div_3_mag_1.JK_FF_mag_1.K 0.0209f
C1042 JK_FF_mag_1.nand2_mag_3.IN1 a_15145_4651# 0.011f
C1043 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_1.OUT 0.25f
C1044 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 0.768f
C1045 a_10956_3003# CLK_div_3_mag_0.Q1 0.01f
C1046 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN a_7289_1356# 4.94e-20
C1047 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_14823_1355# 0.0697f
C1048 JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 4.95e-20
C1049 a_13857_4607# a_14017_4607# 0.0504f
C1050 a_18853_4654# JK_FF_mag_0.nand2_mag_1.IN2 0.00372f
C1051 JK_FF_mag_1.Q a_17001_4610# 0.0101f
C1052 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C1053 a_10674_5199# CLK_div_3_mag_0.Q0 0.00789f
C1054 a_8423_215# CLK_div_3_mag_1.JK_FF_mag_1.K 0.00695f
C1055 VDD a_9141_1312# 2.21e-19
C1056 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.0894f
C1057 CLK_div_3_mag_1.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 0.0435f
C1058 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_0.JK_FF_mag_1.K 0.23f
C1059 RST a_11434_1356# 2.23e-19
C1060 VDD a_17686_214# 9.82e-19
C1061 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C1062 JK_FF_mag_0.nand3_mag_2.OUT Vdiv108 0.338f
C1063 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_11998_1312# 0.0732f
C1064 JK_FF_mag_0.nand3_mag_1.IN1 a_17725_4654# 0.0697f
C1065 RST CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.00702f
C1066 JK_FF_mag_1.nand2_mag_3.IN1 a_14581_4651# 1.43e-19
C1067 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C1068 JK_FF_mag_1.Q JK_FF_mag_0.QB 0.307f
C1069 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.K 1.22e-23
C1070 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_3.IN1 0.233f
C1071 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 a_14259_1355# 0.0059f
C1072 a_15553_214# CLK 0.00117f
C1073 a_12372_4102# CLK_div_3_mag_0.JK_FF_mag_1.K 0.012f
C1074 a_7497_5199# a_7657_5199# 0.0504f
C1075 a_18289_4654# JK_FF_mag_0.nand2_mag_1.IN2 0.069f
C1076 CLK_div_3_mag_1.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K 2.37f
C1077 JK_FF_mag_1.Q a_15709_4651# 0.069f
C1078 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.Q0 8.04e-19
C1079 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C1080 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_12372_4102# 0.00372f
C1081 a_10514_5199# CLK_div_3_mag_0.Q0 0.00335f
C1082 JK_FF_mag_0.nand2_mag_1.IN2 Vdiv108 0.107f
C1083 a_10680_4102# CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 0.00119f
C1084 RST a_10870_1356# 0.00121f
C1085 CLK_div_3_mag_0.JK_FF_mag_1.K JK_FF_mag_1.CLK 0.00199f
C1086 a_11398_5199# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00696f
C1087 VDD CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.654f
C1088 JK_FF_mag_0.nand3_mag_0.OUT VDD 0.742f
C1089 a_17879_3513# JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C1090 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.122f
C1091 VDD a_17122_258# 0.00149f
C1092 a_17686_214# a_17846_214# 0.0504f
C1093 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT a_11434_1356# 0.00378f
C1094 VDD RST 3.29f
C1095 a_17155_3513# CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 1.8e-21
C1096 JK_FF_mag_1.nand2_mag_3.IN1 a_14017_4607# 0.00119f
C1097 CLK_div_3_mag_0.or_2_mag_0.IN2 a_11929_2535# 8.64e-19
C1098 a_15393_214# CLK 0.00164f
C1099 CLK_div_3_mag_0.Q0 CLK_div_3_mag_1.JK_FF_mag_1.K 0.027f
C1100 a_11808_4102# CLK_div_3_mag_0.JK_FF_mag_1.K 2.96e-19
C1101 a_14259_1355# CLK_div_3_mag_2.or_2_mag_0.IN2 4.9e-20
C1102 JK_FF_mag_1.Q a_15145_4651# 3.74e-21
C1103 RST CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 0.00721f
C1104 a_14581_4651# CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 1.46e-22
C1105 a_8987_215# a_9147_215# 0.0504f
C1106 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 0.321f
C1107 CLK_div_3_mag_1.Q0 a_7732_2691# 0.0134f
C1108 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.or_2_mag_0.IN2 3.81e-19
C1109 JK_FF_mag_1.nand3_mag_1.IN1 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 1.22e-19
C1110 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C1111 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 a_11808_4102# 0.069f
C1112 VDD a_8417_1356# 3.14e-19
C1113 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 7.89e-19
C1114 CLK_div_3_mag_1.or_2_mag_0.IN2 a_8705_2455# 7.48e-20
C1115 a_12526_5199# JK_FF_mag_1.CLK 4.77e-20
C1116 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 0.00335f
C1117 RST a_10306_1356# 0.00154f
C1118 JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.399f
C1119 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT a_11962_5199# 0.00378f
C1120 a_11238_5199# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00695f
C1121 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C1122 VDD a_16558_258# 0.00149f
C1123 a_17719_3513# JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C1124 a_15387_1311# CLK_div_3_mag_2.Q0 2.79e-20
C1125 CLK_div_3_mag_0.Q1 a_11929_2535# 6.83e-19
C1126 RST a_17846_214# 8.64e-19
C1127 VDD CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.65f
C1128 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 8.59e-20
C1129 a_11244_4102# CLK_div_3_mag_0.JK_FF_mag_1.K 1.75e-19
C1130 a_8981_1312# a_9141_1312# 0.0504f
C1131 JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.JK_FF_mag_1.K 6.19e-22
C1132 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.Q 0.00335f
C1133 CLK_div_3_mag_2.JK_FF_mag_1.K CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 0.00384f
C1134 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 0.0147f
C1135 VDD a_7853_1356# 3.14e-19
C1136 a_11440_215# CLK_div_3_mag_1.JK_FF_mag_1.QB 0.00695f
C1137 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VDD 0.469f
C1138 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 a_16712_1355# 4.52e-20
C1139 JK_FF_mag_0.QB JK_FF_mag_0.nand3_mag_1.IN1 0.0378f
C1140 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C1141 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_3.IN1 0.16f
C1142 a_11962_5199# JK_FF_mag_1.CLK 1.73e-20
C1143 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.08f
C1144 RST a_9141_1312# 0.00211f
C1145 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK 0.00254f
C1146 a_17686_214# CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C1147 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT 0.159f
C1148 a_17155_3513# JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C1149 VDD a_15553_214# 0.00743f
C1150 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.QB 0.103f
C1151 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.QB 0.198f
C1152 RST a_17686_214# 0.00135f
C1153 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.739f
C1154 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VDD 0.415f
C1155 JK_FF_mag_1.Q a_14017_4607# 2.79e-20
C1156 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.399f
C1157 JK_FF_mag_1.Q CLK_div_3_mag_2.JK_FF_mag_1.K 0.0372f
C1158 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN CLK_div_3_mag_0.JK_FF_mag_1.K 0.00384f
C1159 a_14011_3510# CLK_div_3_mag_0.JK_FF_mag_1.K 9.44e-21
C1160 JK_FF_mag_0.nand2_mag_3.IN1 a_17725_4654# 1.43e-19
C1161 VDD a_7289_1356# 3.56e-19
C1162 a_11280_215# CLK_div_3_mag_1.JK_FF_mag_1.QB 0.00696f
C1163 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_8381_5199# 2.88e-20
C1164 RST a_8981_1312# 0.00152f
C1165 a_16995_3513# JK_FF_mag_0.nand3_mag_2.OUT 0.0202f
C1166 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK 6.62e-20
C1167 CLK_div_3_mag_1.JK_FF_mag_1.QB CLK_div_3_mag_1.JK_FF_mag_1.K 3.28e-19
C1168 VDD a_15393_214# 0.00305f
C1169 VDD CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.654f
C1170 RST CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 0.196f
C1171 JK_FF_mag_0.nand3_mag_0.OUT RST 0.00523f
C1172 VDD a_7135_259# 3.14e-19
C1173 RST a_17122_258# 5.68e-19
C1174 JK_FF_mag_1.QB JK_FF_mag_0.nand2_mag_3.IN1 2.72e-19
C1175 CLK_div_3_mag_0.or_2_mag_0.IN2 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.53e-20
C1176 JK_FF_mag_1.nand3_mag_1.OUT CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 5.14e-20
C1177 CLK_div_3_mag_2.JK_FF_mag_1.QB a_18404_1311# 0.00392f
C1178 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 CLK_div_3_mag_2.Q0 0.107f
C1179 CLK_div_3_mag_0.Q0 a_11929_2535# 0.0134f
C1180 CLK_div_3_mag_0.JK_FF_mag_1.K CLK_div_3_mag_1.JK_FF_mag_1.K 0.089f
C1181 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C1182 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT 0.00183f
C1183 JK_FF_mag_0.nand2_mag_3.IN1 a_17161_4610# 0.00119f
C1184 a_13851_3510# CLK_div_3_mag_0.JK_FF_mag_1.K 1.17e-20
C1185 a_10716_259# CLK_div_3_mag_1.JK_FF_mag_1.QB 0.00964f
C1186 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_8221_5199# 9.1e-19
C1187 CLK_div_3_mag_0.Q1 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 5.95e-20
C1188 VDD CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C1189 RST a_8417_1356# 5.58e-19
C1190 CLK_div_3_mag_2.or_2_mag_0.IN2 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.0445f
C1191 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT CLK_div_3_mag_0.Q1 0.101f
C1192 VDD a_14829_214# 2.21e-19
C1193 JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 1.26e-19
C1194 JK_FF_mag_1.nand2_mag_1.IN2 RST 0.00422f
C1195 a_13695_1355# CLK_div_3_mag_2.Q0 0.069f
C1196 RST a_16558_258# 0.00114f
C1197 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.Q 0.0343f
C1198 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 CLK 1.31f
C1199 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0622f
C1200 CLK_div_3_mag_2.JK_FF_mag_1.QB a_17840_1355# 3.33e-19
C1201 JK_FF_mag_1.QB CLK_div_3_mag_0.Q0 2.61e-19
C1202 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_15387_1311# 0.00119f
C1203 RST CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT 0.0042f
C1204 VDD CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 0.652f
C1205 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN 6.11e-19
C1206 JK_FF_mag_1.nand2_mag_4.IN2 a_15709_4651# 4.52e-20
C1207 a_7732_2691# CLK_div_3_mag_0.JK_FF_mag_1.K 0.00263f
C1208 a_8981_1312# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.00119f
C1209 a_15299_3554# CLK 3.54e-21
C1210 a_10152_259# CLK_div_3_mag_1.JK_FF_mag_1.QB 0.0811f
C1211 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_7657_5199# 0.0731f
C1212 RST a_7853_1356# 5.01e-19
C1213 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN RST 0.00333f
C1214 RST CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 0.0541f
C1215 a_12158_1312# CLK_div_3_mag_2.Q0 3.51e-19
C1216 CLK_div_3_mag_0.Q1 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT 0.0343f
C1217 RST a_15553_214# 0.00218f
C1218 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.Q 0.0179f
C1219 JK_FF_mag_0.nand3_mag_1.IN1 CLK_div_3_mag_2.JK_FF_mag_1.K 6.13e-20
C1220 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 a_14823_1355# 1.43e-19
C1221 a_12164_215# CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C1222 RST CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT 0.107f
C1223 JK_FF_mag_1.QB Vdiv108 1.43e-19
C1224 JK_FF_mag_0.QB JK_FF_mag_0.nand2_mag_3.IN1 0.28f
C1225 JK_FF_mag_1.Q CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT 4.18e-21
C1226 VDD CLK_div_3_mag_2.or_2_mag_0.IN2 0.49f
C1227 a_8417_1356# CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C1228 CLK_div_3_mag_2.Q0 CLK 0.149f
C1229 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.Q0 5.26e-19
C1230 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 RST 0.00797f
C1231 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT 0.121f
C1232 Vdiv108 CLK_div_3_mag_2.JK_FF_mag_1.QB 5.82e-21
C1233 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT a_7497_5199# 0.0202f
C1234 JK_FF_mag_1.CLK CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN 0.00121f
C1235 CLK_div_3_mag_2.JK_FF_mag_1.QB CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C1236 RST a_7289_1356# 5.01e-19
C1237 CLK_div_3_mag_1.JK_FF_mag_1.QB a_11929_2535# 2.51e-19
C1238 a_10520_4102# CLK_div_3_mag_0.Q1 0.00149f
C1239 VDD a_14105_258# 3.14e-19
C1240 Vdiv108 a_17161_4610# 2.79e-20
C1241 CLK_div_3_mag_0.Q0 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 1.99e-20
C1242 JK_FF_mag_0.nand3_mag_2.OUT CLK 1.17e-20
C1243 JK_FF_mag_1.nand3_mag_2.OUT VDD 0.756f
C1244 CLK_div_3_mag_0.Q1 a_8381_5199# 0.0101f
C1245 RST a_15393_214# 0.00218f
C1246 RST CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 0.143f
C1247 RST a_7135_259# 0.00114f
C1248 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT 0.00183f
C1249 JK_FF_mag_1.nand3_mag_0.OUT CLK_div_3_mag_2.or_2_mag_0.IN2 1.19e-20
C1250 a_18570_214# VSS 0.0881f
C1251 a_18410_214# VSS 0.0343f
C1252 a_17846_214# VSS 0.0881f
C1253 a_17686_214# VSS 0.0343f
C1254 a_17122_258# VSS 0.0676f
C1255 a_16558_258# VSS 0.0675f
C1256 a_15553_214# VSS 0.0881f
C1257 a_15393_214# VSS 0.0343f
C1258 a_14829_214# VSS 0.0881f
C1259 a_14669_214# VSS 0.0343f
C1260 a_14105_258# VSS 0.0676f
C1261 a_13541_258# VSS 0.0675f
C1262 a_12164_215# VSS 0.0881f
C1263 a_12004_215# VSS 0.0343f
C1264 a_11440_215# VSS 0.0881f
C1265 a_11280_215# VSS 0.0343f
C1266 a_10716_259# VSS 0.0676f
C1267 a_10152_259# VSS 0.0675f
C1268 a_9147_215# VSS 0.0881f
C1269 a_8987_215# VSS 0.0343f
C1270 a_8423_215# VSS 0.0881f
C1271 a_8263_215# VSS 0.0343f
C1272 a_7699_259# VSS 0.0676f
C1273 a_7135_259# VSS 0.0675f
C1274 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C1275 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C1276 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.541f
C1277 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C1278 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.521f
C1279 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.417f
C1280 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.541f
C1281 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.417f
C1282 a_18564_1311# VSS 0.0881f
C1283 a_18404_1311# VSS 0.0343f
C1284 a_17840_1355# VSS 0.0676f
C1285 a_17276_1355# VSS 0.0676f
C1286 a_16712_1355# VSS 0.0676f
C1287 a_15547_1311# VSS 0.0881f
C1288 a_15387_1311# VSS 0.0343f
C1289 a_14823_1355# VSS 0.0676f
C1290 a_14259_1355# VSS 0.0676f
C1291 a_13695_1355# VSS 0.0676f
C1292 a_12158_1312# VSS 0.0881f
C1293 a_11998_1312# VSS 0.0343f
C1294 a_11434_1356# VSS 0.0676f
C1295 a_10870_1356# VSS 0.0676f
C1296 a_10306_1356# VSS 0.0676f
C1297 a_9141_1312# VSS 0.0881f
C1298 a_8981_1312# VSS 0.0343f
C1299 a_8417_1356# VSS 0.0676f
C1300 a_7853_1356# VSS 0.0676f
C1301 a_7289_1356# VSS 0.0676f
C1302 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C1303 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.811f
C1304 CLK_div_3_mag_2.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.726f
C1305 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.699f
C1306 CLK_div_3_mag_2.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1307 CLK_div_3_mag_2.JK_FF_mag_1.QB VSS 0.859f
C1308 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1309 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C1310 CLK_div_3_mag_2.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C1311 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.692f
C1312 CLK_div_3_mag_2.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.414f
C1313 CLK_div_3_mag_2.JK_FF_mag_1.K VSS 4.43f
C1314 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C1315 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.809f
C1316 CLK_div_3_mag_1.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.724f
C1317 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.698f
C1318 CLK_div_3_mag_1.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1319 CLK_div_3_mag_1.JK_FF_mag_1.QB VSS 0.857f
C1320 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1321 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.811f
C1322 CLK_div_3_mag_1.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.726f
C1323 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.692f
C1324 CLK_div_3_mag_1.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1325 CLK_div_3_mag_1.JK_FF_mag_1.K VSS 4.19f
C1326 a_15111_2454# VSS 0.0676f
C1327 a_14138_2690# VSS 0.0247f
C1328 a_11929_2535# VSS 0.0247f
C1329 a_8705_2455# VSS 0.0676f
C1330 CLK_div_3_mag_2.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.598f
C1331 CLK VSS 2.77f
C1332 CLK_div_3_mag_2.and2_mag_0.GF_INV_MAG_0.IN VSS 0.434f
C1333 CLK_div_3_mag_2.or_2_mag_0.IN2 VSS 0.419f
C1334 CLK_div_3_mag_2.Q0 VSS 2.65f
C1335 CLK_div_3_mag_0.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.597f
C1336 CLK_div_3_mag_0.or_2_mag_0.IN2 VSS 0.416f
C1337 CLK_div_3_mag_0.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C1338 a_10956_3003# VSS 0.0676f
C1339 a_7732_2691# VSS 0.0247f
C1340 CLK_div_3_mag_1.or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C1341 CLK_div_3_mag_1.and2_mag_0.GF_INV_MAG_0.IN VSS 0.433f
C1342 CLK_div_3_mag_1.or_2_mag_0.IN2 VSS 0.416f
C1343 CLK_div_3_mag_1.Q0 VSS 2.76f
C1344 a_19007_3557# VSS 0.0729f
C1345 a_18443_3557# VSS 0.073f
C1346 a_17879_3513# VSS 0.0439f
C1347 a_17719_3513# VSS 0.0977f
C1348 a_17155_3513# VSS 0.0439f
C1349 a_16995_3513# VSS 0.0978f
C1350 a_15863_3554# VSS 0.0736f
C1351 a_15299_3554# VSS 0.0737f
C1352 a_14735_3510# VSS 0.0454f
C1353 a_14575_3510# VSS 0.0992f
C1354 a_14011_3510# VSS 0.0454f
C1355 a_13851_3510# VSS 0.0992f
C1356 JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.423f
C1357 JK_FF_mag_0.nand3_mag_2.OUT VSS 0.57f
C1358 JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.424f
C1359 JK_FF_mag_1.nand3_mag_2.OUT VSS 0.57f
C1360 a_12372_4102# VSS 0.0676f
C1361 a_11808_4102# VSS 0.0676f
C1362 a_11244_4102# VSS 0.0676f
C1363 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1364 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1365 a_10680_4102# VSS 0.0343f
C1366 a_10520_4102# VSS 0.0881f
C1367 a_9355_4102# VSS 0.0676f
C1368 a_8791_4102# VSS 0.0676f
C1369 a_8227_4102# VSS 0.0676f
C1370 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1371 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_0.OUT VSS 0.508f
C1372 a_7663_4102# VSS 0.0343f
C1373 a_7503_4102# VSS 0.0881f
C1374 a_18853_4654# VSS 0.0676f
C1375 a_18289_4654# VSS 0.0676f
C1376 a_17725_4654# VSS 0.0676f
C1377 a_17161_4610# VSS 0.0343f
C1378 a_17001_4610# VSS 0.0881f
C1379 a_15709_4651# VSS 0.0676f
C1380 a_15145_4651# VSS 0.0676f
C1381 a_14581_4651# VSS 0.0676f
C1382 a_14017_4607# VSS 0.0343f
C1383 a_13857_4607# VSS 0.0881f
C1384 Vdiv108 VSS 1.5f
C1385 JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C1386 JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.835f
C1387 JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.725f
C1388 JK_FF_mag_0.nand3_mag_1.OUT VSS 0.84f
C1389 JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C1390 JK_FF_mag_0.QB VSS 0.88f
C1391 JK_FF_mag_1.Q VSS 2.1f
C1392 JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C1393 JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.84f
C1394 JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.723f
C1395 JK_FF_mag_1.nand3_mag_1.OUT VSS 0.84f
C1396 JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C1397 JK_FF_mag_1.QB VSS 0.906f
C1398 JK_FF_mag_1.CLK VSS 2.12f
C1399 CLK_div_3_mag_0.JK_FF_mag_1.K VSS 4.4f
C1400 a_12526_5199# VSS 0.0675f
C1401 a_11962_5199# VSS 0.0676f
C1402 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C1403 CLK_div_3_mag_0.JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.69f
C1404 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.OUT VSS 0.809f
C1405 a_11398_5199# VSS 0.0343f
C1406 a_11238_5199# VSS 0.0881f
C1407 a_10674_5199# VSS 0.0343f
C1408 a_10514_5199# VSS 0.0881f
C1409 CLK_div_3_mag_0.JK_FF_mag_1.QB VSS 0.857f
C1410 a_9509_5199# VSS 0.0675f
C1411 a_8945_5199# VSS 0.0676f
C1412 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.416f
C1413 CLK_div_3_mag_0.JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.697f
C1414 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.OUT VSS 0.808f
C1415 a_8381_5199# VSS 0.0343f
C1416 a_8221_5199# VSS 0.0881f
C1417 a_7657_5199# VSS 0.0343f
C1418 a_7497_5199# VSS 0.0881f
C1419 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C1420 CLK_div_3_mag_0.JK_FF_mag_0.nand3_mag_2.OUT VSS 0.539f
C1421 CLK_div_3_mag_0.Q0 VSS 1.64f
C1422 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.722f
C1423 RST VSS 7.24f
C1424 CLK_div_3_mag_0.JK_FF_mag_1.nand3_mag_2.OUT VSS 0.519f
C1425 CLK_div_3_mag_0.Q1 VSS 1.7f
C1426 VDD VSS 0.138p
C1427 CLK_div_3_mag_1.JK_FF_mag_1.K.n0 VSS 2.12f
C1428 CLK_div_3_mag_1.JK_FF_mag_1.K.t0 VSS 0.0346f
C1429 CLK_div_3_mag_1.JK_FF_mag_1.K.n1 VSS 0.0346f
C1430 CLK_div_3_mag_1.JK_FF_mag_1.K.n2 VSS 0.0817f
C1431 CLK_div_3_mag_1.JK_FF_mag_1.K.t3 VSS 0.0554f
C1432 CLK_div_3_mag_1.JK_FF_mag_1.K.t2 VSS 0.0714f
C1433 CLK_div_3_mag_1.JK_FF_mag_1.K.n3 VSS 0.141f
C1434 CLK_div_3_mag_1.JK_FF_mag_1.K.t5 VSS 0.0443f
C1435 CLK_div_3_mag_1.JK_FF_mag_1.K.t7 VSS 0.0553f
C1436 CLK_div_3_mag_1.JK_FF_mag_1.K.n4 VSS 0.143f
C1437 CLK_div_3_mag_1.JK_FF_mag_1.K.t6 VSS 0.0779f
C1438 CLK_div_3_mag_1.JK_FF_mag_1.K.t4 VSS 0.0496f
C1439 CLK_div_3_mag_1.JK_FF_mag_1.K.n5 VSS 0.138f
C1440 CLK_div_3_mag_1.JK_FF_mag_1.K.n6 VSS 1.18f
C1441 CLK_div_3_mag_1.JK_FF_mag_1.K.n7 VSS 0.268f
C1442 CLK_div_3_mag_1.Q0.t0 VSS 0.0246f
C1443 CLK_div_3_mag_1.Q0.t1 VSS 0.0203f
C1444 CLK_div_3_mag_1.Q0.n0 VSS 0.0203f
C1445 CLK_div_3_mag_1.Q0.n1 VSS 0.0557f
C1446 CLK_div_3_mag_1.Q0.t3 VSS 0.0632f
C1447 CLK_div_3_mag_1.Q0.t7 VSS 0.0195f
C1448 CLK_div_3_mag_1.Q0.n2 VSS 0.0665f
C1449 CLK_div_3_mag_1.Q0.t5 VSS 0.0298f
C1450 CLK_div_3_mag_1.Q0.t6 VSS 0.0452f
C1451 CLK_div_3_mag_1.Q0.n3 VSS 0.0802f
C1452 CLK_div_3_mag_1.Q0.t8 VSS 0.0259f
C1453 CLK_div_3_mag_1.Q0.t4 VSS 0.0324f
C1454 CLK_div_3_mag_1.Q0.n4 VSS 0.0753f
C1455 CLK_div_3_mag_1.Q0.n5 VSS 0.597f
C1456 CLK_div_3_mag_1.Q0.n6 VSS 0.441f
C1457 CLK_div_3_mag_0.JK_FF_mag_1.K.n0 VSS 2.2f
C1458 CLK_div_3_mag_0.JK_FF_mag_1.K.n1 VSS 0.159f
C1459 CLK_div_3_mag_0.JK_FF_mag_1.K.t3 VSS 0.0515f
C1460 CLK_div_3_mag_0.JK_FF_mag_1.K.t4 VSS 0.0808f
C1461 CLK_div_3_mag_0.JK_FF_mag_1.K.n2 VSS 0.143f
C1462 CLK_div_3_mag_0.JK_FF_mag_1.K.t7 VSS 0.0739f
C1463 CLK_div_3_mag_0.JK_FF_mag_1.K.t8 VSS 0.0576f
C1464 CLK_div_3_mag_0.JK_FF_mag_1.K.n3 VSS 0.147f
C1465 CLK_div_3_mag_0.JK_FF_mag_1.K.t5 VSS 0.046f
C1466 CLK_div_3_mag_0.JK_FF_mag_1.K.t6 VSS 0.0576f
C1467 CLK_div_3_mag_0.JK_FF_mag_1.K.n4 VSS 0.148f
C1468 CLK_div_3_mag_0.JK_FF_mag_1.K.n5 VSS 1.23f
C1469 CLK_div_3_mag_0.JK_FF_mag_1.K.t0 VSS 0.0359f
C1470 CLK_div_3_mag_0.JK_FF_mag_1.K.n6 VSS 0.0359f
C1471 CLK_div_3_mag_0.JK_FF_mag_1.K.n7 VSS 0.0766f
C1472 CLK_div_3_mag_1.Q1.n0 VSS 0.317f
C1473 CLK_div_3_mag_1.Q1.t2 VSS 0.0207f
C1474 CLK_div_3_mag_1.Q1.t0 VSS 0.0171f
C1475 CLK_div_3_mag_1.Q1.n1 VSS 0.0171f
C1476 CLK_div_3_mag_1.Q1.n2 VSS 0.047f
C1477 CLK_div_3_mag_1.Q1.t8 VSS 0.0273f
C1478 CLK_div_3_mag_1.Q1.t7 VSS 0.0352f
C1479 CLK_div_3_mag_1.Q1.n3 VSS 0.0697f
C1480 CLK_div_3_mag_1.Q1.t3 VSS 0.0218f
C1481 CLK_div_3_mag_1.Q1.t5 VSS 0.0273f
C1482 CLK_div_3_mag_1.Q1.n4 VSS 0.0618f
C1483 CLK_div_3_mag_1.Q1.t9 VSS 0.0251f
C1484 CLK_div_3_mag_1.Q1.t10 VSS 0.0381f
C1485 CLK_div_3_mag_1.Q1.n5 VSS 0.0676f
C1486 CLK_div_3_mag_1.Q1.t4 VSS 0.0218f
C1487 CLK_div_3_mag_1.Q1.t6 VSS 0.0273f
C1488 CLK_div_3_mag_1.Q1.n6 VSS 0.0634f
C1489 CLK_div_3_mag_1.Q1.n7 VSS 0.499f
C1490 CLK_div_3_mag_1.Q1.n8 VSS 0.207f
C1491 CLK_div_3_mag_2.Q0.t2 VSS 0.0246f
C1492 CLK_div_3_mag_2.Q0.t0 VSS 0.0203f
C1493 CLK_div_3_mag_2.Q0.n0 VSS 0.0203f
C1494 CLK_div_3_mag_2.Q0.n1 VSS 0.0557f
C1495 CLK_div_3_mag_2.Q0.t3 VSS 0.0632f
C1496 CLK_div_3_mag_2.Q0.t7 VSS 0.0195f
C1497 CLK_div_3_mag_2.Q0.n2 VSS 0.0665f
C1498 CLK_div_3_mag_2.Q0.t5 VSS 0.0298f
C1499 CLK_div_3_mag_2.Q0.t6 VSS 0.0452f
C1500 CLK_div_3_mag_2.Q0.n3 VSS 0.0802f
C1501 CLK_div_3_mag_2.Q0.t8 VSS 0.0259f
C1502 CLK_div_3_mag_2.Q0.t4 VSS 0.0324f
C1503 CLK_div_3_mag_2.Q0.n4 VSS 0.0753f
C1504 CLK_div_3_mag_2.Q0.n5 VSS 0.597f
C1505 CLK_div_3_mag_2.Q0.n6 VSS 0.441f
C1506 CLK_div_3_mag_0.CLK.n0 VSS 0.521f
C1507 CLK_div_3_mag_0.CLK.n1 VSS 0.0208f
C1508 CLK_div_3_mag_0.CLK.n2 VSS 0.337f
C1509 CLK_div_3_mag_0.CLK.n3 VSS 0.0208f
C1510 CLK_div_3_mag_0.CLK.n4 VSS 0.141f
C1511 CLK_div_3_mag_0.CLK.n5 VSS 0.131f
C1512 CLK_div_3_mag_0.CLK.n6 VSS 0.0495f
C1513 CLK_div_3_mag_0.CLK.n7 VSS 0.0495f
C1514 CLK_div_3_mag_0.CLK.t0 VSS 0.0571f
C1515 CLK_div_3_mag_0.CLK.t1 VSS 0.0172f
C1516 CLK_div_3_mag_0.CLK.n8 VSS 0.198f
C1517 CLK_div_3_mag_0.CLK.t11 VSS 0.0509f
C1518 CLK_div_3_mag_0.CLK.t10 VSS 0.0335f
C1519 CLK_div_3_mag_0.CLK.n9 VSS 0.09f
C1520 CLK_div_3_mag_0.CLK.t8 VSS 0.0509f
C1521 CLK_div_3_mag_0.CLK.t7 VSS 0.0335f
C1522 CLK_div_3_mag_0.CLK.n10 VSS 0.09f
C1523 CLK_div_3_mag_0.CLK.t2 VSS 0.0509f
C1524 CLK_div_3_mag_0.CLK.t3 VSS 0.0335f
C1525 CLK_div_3_mag_0.CLK.n11 VSS 0.09f
C1526 CLK_div_3_mag_0.CLK.t13 VSS 0.0472f
C1527 CLK_div_3_mag_0.CLK.t14 VSS 0.0264f
C1528 CLK_div_3_mag_0.CLK.n12 VSS 0.0899f
C1529 CLK_div_3_mag_0.CLK.n13 VSS 0.288f
C1530 CLK_div_3_mag_0.CLK.t5 VSS 0.0509f
C1531 CLK_div_3_mag_0.CLK.t4 VSS 0.0335f
C1532 CLK_div_3_mag_0.CLK.n14 VSS 0.09f
C1533 CLK_div_3_mag_0.CLK.t6 VSS 0.042f
C1534 CLK_div_3_mag_0.CLK.t9 VSS 0.0109f
C1535 CLK_div_3_mag_0.CLK.n15 VSS 0.0697f
C1536 CLK_div_3_mag_0.CLK.n16 VSS 0.671f
C1537 CLK_div_3_mag_0.CLK.n17 VSS 0.67f
C1538 CLK_div_3_mag_0.CLK.t12 VSS 0.042f
C1539 CLK_div_3_mag_0.CLK.t15 VSS 0.0109f
C1540 CLK_div_3_mag_0.CLK.n18 VSS 0.0697f
C1541 CLK.n0 VSS 0.0183f
C1542 CLK.t1 VSS 0.0348f
C1543 CLK.t4 VSS 0.0528f
C1544 CLK.n1 VSS 0.0933f
C1545 CLK.n2 VSS 0.0122f
C1546 CLK.n3 VSS 0.00876f
C1547 CLK.n4 VSS 0.00438f
C1548 CLK.n5 VSS 0.0171f
C1549 CLK.n6 VSS 0.173f
C1550 CLK.n7 VSS 0.175f
C1551 CLK.t2 VSS 0.0348f
C1552 CLK.t5 VSS 0.0528f
C1553 CLK.n8 VSS 0.0933f
C1554 CLK.n9 VSS 0.0122f
C1555 CLK.n10 VSS 0.00876f
C1556 CLK.n11 VSS 0.00433f
C1557 CLK.n12 VSS 0.101f
C1558 CLK.t12 VSS 0.049f
C1559 CLK.t3 VSS 0.0273f
C1560 CLK.n13 VSS 0.0932f
C1561 CLK.n14 VSS 0.299f
C1562 CLK.t6 VSS 0.0348f
C1563 CLK.t8 VSS 0.0528f
C1564 CLK.n15 VSS 0.0933f
C1565 CLK.n16 VSS 0.0122f
C1566 CLK.n17 VSS 0.00876f
C1567 CLK.n18 VSS 0.00438f
C1568 CLK.n19 VSS 0.0171f
C1569 CLK.n20 VSS 0.161f
C1570 CLK.n21 VSS 0.362f
C1571 CLK.n22 VSS 0.0135f
C1572 CLK.t9 VSS 0.0348f
C1573 CLK.t11 VSS 0.0528f
C1574 CLK.n23 VSS 0.0933f
C1575 CLK.n24 VSS 0.0122f
C1576 CLK.n25 VSS 0.00876f
C1577 CLK.n26 VSS 0.00433f
C1578 CLK.n27 VSS 0.101f
C1579 CLK.n28 VSS 0.0183f
C1580 CLK.n29 VSS 0.0314f
C1581 CLK.t10 VSS 0.0436f
C1582 CLK.t0 VSS 0.0111f
C1583 CLK.n30 VSS 0.0722f
C1584 CLK.n31 VSS 0.0153f
C1585 CLK.n32 VSS 0.00533f
C1586 CLK.n33 VSS 0.0116f
C1587 CLK.n34 VSS 0.667f
C1588 CLK.n35 VSS 0.668f
C1589 CLK.n36 VSS 0.0116f
C1590 CLK.t7 VSS 0.0436f
C1591 CLK.t13 VSS 0.0111f
C1592 CLK.n37 VSS 0.0722f
C1593 CLK.n38 VSS 0.0153f
C1594 CLK.n39 VSS 0.00533f
C1595 CLK.n40 VSS 0.0148f
C1596 CLK_div_3_mag_2.JK_FF_mag_1.K.n0 VSS 2.06f
C1597 CLK_div_3_mag_2.JK_FF_mag_1.K.t1 VSS 0.0336f
C1598 CLK_div_3_mag_2.JK_FF_mag_1.K.n1 VSS 0.0336f
C1599 CLK_div_3_mag_2.JK_FF_mag_1.K.n2 VSS 0.0793f
C1600 CLK_div_3_mag_2.JK_FF_mag_1.K.t4 VSS 0.0538f
C1601 CLK_div_3_mag_2.JK_FF_mag_1.K.t2 VSS 0.0693f
C1602 CLK_div_3_mag_2.JK_FF_mag_1.K.n3 VSS 0.137f
C1603 CLK_div_3_mag_2.JK_FF_mag_1.K.t3 VSS 0.043f
C1604 CLK_div_3_mag_2.JK_FF_mag_1.K.t5 VSS 0.0537f
C1605 CLK_div_3_mag_2.JK_FF_mag_1.K.n4 VSS 0.139f
C1606 CLK_div_3_mag_2.JK_FF_mag_1.K.t7 VSS 0.0756f
C1607 CLK_div_3_mag_2.JK_FF_mag_1.K.t6 VSS 0.0482f
C1608 CLK_div_3_mag_2.JK_FF_mag_1.K.n5 VSS 0.134f
C1609 CLK_div_3_mag_2.JK_FF_mag_1.K.n6 VSS 1.15f
C1610 CLK_div_3_mag_2.JK_FF_mag_1.K.n7 VSS 0.261f
C1611 CLK_div_3_mag_2.Q1.n0 VSS 0.317f
C1612 CLK_div_3_mag_2.Q1.t1 VSS 0.0207f
C1613 CLK_div_3_mag_2.Q1.t2 VSS 0.0171f
C1614 CLK_div_3_mag_2.Q1.n1 VSS 0.0171f
C1615 CLK_div_3_mag_2.Q1.n2 VSS 0.047f
C1616 CLK_div_3_mag_2.Q1.t7 VSS 0.0273f
C1617 CLK_div_3_mag_2.Q1.t5 VSS 0.0352f
C1618 CLK_div_3_mag_2.Q1.n3 VSS 0.0697f
C1619 CLK_div_3_mag_2.Q1.t3 VSS 0.0218f
C1620 CLK_div_3_mag_2.Q1.t4 VSS 0.0273f
C1621 CLK_div_3_mag_2.Q1.n4 VSS 0.0618f
C1622 CLK_div_3_mag_2.Q1.t8 VSS 0.0251f
C1623 CLK_div_3_mag_2.Q1.t10 VSS 0.0381f
C1624 CLK_div_3_mag_2.Q1.n5 VSS 0.0676f
C1625 CLK_div_3_mag_2.Q1.t6 VSS 0.0218f
C1626 CLK_div_3_mag_2.Q1.t9 VSS 0.0273f
C1627 CLK_div_3_mag_2.Q1.n6 VSS 0.0634f
C1628 CLK_div_3_mag_2.Q1.n7 VSS 0.499f
C1629 CLK_div_3_mag_2.Q1.n8 VSS 0.207f
C1630 CLK_div_3_mag_1.CLK.n0 VSS 0.511f
C1631 CLK_div_3_mag_1.CLK.n1 VSS 0.322f
C1632 CLK_div_3_mag_1.CLK.n2 VSS 0.0205f
C1633 CLK_div_3_mag_1.CLK.n3 VSS 0.0485f
C1634 CLK_div_3_mag_1.CLK.n4 VSS 0.0485f
C1635 CLK_div_3_mag_1.CLK.t0 VSS 0.0562f
C1636 CLK_div_3_mag_1.CLK.t1 VSS 0.0169f
C1637 CLK_div_3_mag_1.CLK.n5 VSS 0.194f
C1638 CLK_div_3_mag_1.CLK.t3 VSS 0.033f
C1639 CLK_div_3_mag_1.CLK.t7 VSS 0.0501f
C1640 CLK_div_3_mag_1.CLK.n6 VSS 0.0885f
C1641 CLK_div_3_mag_1.CLK.t9 VSS 0.033f
C1642 CLK_div_3_mag_1.CLK.t11 VSS 0.0501f
C1643 CLK_div_3_mag_1.CLK.n7 VSS 0.0885f
C1644 CLK_div_3_mag_1.CLK.t15 VSS 0.0465f
C1645 CLK_div_3_mag_1.CLK.t5 VSS 0.0259f
C1646 CLK_div_3_mag_1.CLK.n8 VSS 0.0884f
C1647 CLK_div_3_mag_1.CLK.n9 VSS 0.283f
C1648 CLK_div_3_mag_1.CLK.t10 VSS 0.033f
C1649 CLK_div_3_mag_1.CLK.t12 VSS 0.0501f
C1650 CLK_div_3_mag_1.CLK.n10 VSS 0.0885f
C1651 CLK_div_3_mag_1.CLK.t2 VSS 0.033f
C1652 CLK_div_3_mag_1.CLK.t6 VSS 0.0501f
C1653 CLK_div_3_mag_1.CLK.n11 VSS 0.0885f
C1654 CLK_div_3_mag_1.CLK.t13 VSS 0.0414f
C1655 CLK_div_3_mag_1.CLK.t4 VSS 0.0106f
C1656 CLK_div_3_mag_1.CLK.n12 VSS 0.0686f
C1657 CLK_div_3_mag_1.CLK.n13 VSS 0.66f
C1658 CLK_div_3_mag_1.CLK.n14 VSS 0.66f
C1659 CLK_div_3_mag_1.CLK.t8 VSS 0.0414f
C1660 CLK_div_3_mag_1.CLK.t14 VSS 0.0106f
C1661 CLK_div_3_mag_1.CLK.n15 VSS 0.0686f
C1662 RST.n0 VSS 0.00428f
C1663 RST.n1 VSS 0.00228f
C1664 RST.t5 VSS 0.00953f
C1665 RST.t4 VSS 0.015f
C1666 RST.n2 VSS 0.0264f
C1667 RST.n3 VSS 0.00339f
C1668 RST.n4 VSS 0.00121f
C1669 RST.n5 VSS 0.0665f
C1670 RST.n6 VSS 0.00461f
C1671 RST.n7 VSS 0.00142f
C1672 RST.t7 VSS 0.0149f
C1673 RST.t6 VSS 0.0098f
C1674 RST.n8 VSS 0.0263f
C1675 RST.n9 VSS 0.00339f
C1676 RST.n10 VSS 0.00123f
C1677 RST.n11 VSS 0.0919f
C1678 RST.n12 VSS 0.367f
C1679 RST.n13 VSS 0.00154f
C1680 RST.n14 VSS 0.00461f
C1681 RST.t15 VSS 0.0098f
C1682 RST.t1 VSS 0.0149f
C1683 RST.n15 VSS 0.0263f
C1684 RST.n16 VSS 0.00343f
C1685 RST.n17 VSS 0.00123f
C1686 RST.n18 VSS 0.0982f
C1687 RST.t2 VSS 0.0098f
C1688 RST.t3 VSS 0.0149f
C1689 RST.n19 VSS 0.0264f
C1690 RST.n20 VSS 0.0794f
C1691 RST.n21 VSS 0.00458f
C1692 RST.n22 VSS 0.00568f
C1693 RST.n23 VSS 0.002f
C1694 RST.t12 VSS 0.0098f
C1695 RST.t14 VSS 0.0149f
C1696 RST.n24 VSS 0.0263f
C1697 RST.n25 VSS 0.00372f
C1698 RST.n26 VSS 0.00144f
C1699 RST.n27 VSS 7.41e-19
C1700 RST.n28 VSS 0.00155f
C1701 RST.n29 VSS 0.00881f
C1702 RST.n30 VSS 0.0766f
C1703 RST.n31 VSS 0.399f
C1704 RST.n32 VSS 0.311f
C1705 RST.n33 VSS 0.00441f
C1706 RST.t11 VSS 0.015f
C1707 RST.t9 VSS 0.00956f
C1708 RST.n34 VSS 0.0264f
C1709 RST.n35 VSS 0.00343f
C1710 RST.n36 VSS 0.00228f
C1711 RST.n37 VSS 0.00121f
C1712 RST.n38 VSS 0.0362f
C1713 RST.n39 VSS 0.264f
C1714 RST.n40 VSS 0.00154f
C1715 RST.n41 VSS 0.00461f
C1716 RST.t13 VSS 0.0098f
C1717 RST.t0 VSS 0.0149f
C1718 RST.n42 VSS 0.0263f
C1719 RST.n43 VSS 0.00343f
C1720 RST.n44 VSS 0.00123f
C1721 RST.n45 VSS 0.0854f
C1722 RST.n46 VSS 0.267f
C1723 RST.n47 VSS 0.289f
C1724 RST.n48 VSS 0.00441f
C1725 RST.t10 VSS 0.015f
C1726 RST.t8 VSS 0.00956f
C1727 RST.n49 VSS 0.0264f
C1728 RST.n50 VSS 0.00343f
C1729 RST.n51 VSS 0.00228f
C1730 RST.n52 VSS 0.00121f
C1731 RST.n53 VSS 0.0362f
C1732 RST.n54 VSS 0.149f
C1733 RST.n55 VSS 0.103f
C1734 RST.n56 VSS 0.0416f
C1735 VDD.t15 VSS 0.00772f
C1736 VDD.t143 VSS 0.00614f
C1737 VDD.t200 VSS 0.0811f
C1738 VDD.n0 VSS 0.00613f
C1739 VDD.t393 VSS 0.00614f
C1740 VDD.n1 VSS 0.00613f
C1741 VDD.n2 VSS 0.112f
C1742 VDD.t308 VSS 0.0799f
C1743 VDD.n3 VSS 0.00613f
C1744 VDD.n4 VSS 0.00613f
C1745 VDD.t417 VSS 0.0799f
C1746 VDD.n5 VSS 0.0381f
C1747 VDD.t63 VSS 0.00614f
C1748 VDD.n6 VSS 0.00613f
C1749 VDD.t62 VSS 0.074f
C1750 VDD.t75 VSS 0.0811f
C1751 VDD.n7 VSS 0.0381f
C1752 VDD.t204 VSS 0.00614f
C1753 VDD.t391 VSS 0.00252f
C1754 VDD.n8 VSS 0.00252f
C1755 VDD.n9 VSS 0.00551f
C1756 VDD.t203 VSS 0.074f
C1757 VDD.t390 VSS 0.0904f
C1758 VDD.t278 VSS 0.042f
C1759 VDD.n10 VSS 0.0381f
C1760 VDD.t434 VSS 0.00614f
C1761 VDD.t416 VSS 0.00252f
C1762 VDD.n11 VSS 0.00252f
C1763 VDD.n12 VSS 0.00551f
C1764 VDD.t433 VSS 0.074f
C1765 VDD.t415 VSS 0.0904f
C1766 VDD.t19 VSS 0.042f
C1767 VDD.t169 VSS 0.0738f
C1768 VDD.n13 VSS 0.0381f
C1769 VDD.t170 VSS 0.00614f
C1770 VDD.t141 VSS 0.00527f
C1771 VDD.t453 VSS 0.00399f
C1772 VDD.n14 VSS 0.0106f
C1773 VDD.t168 VSS 0.00527f
C1774 VDD.t457 VSS 0.00399f
C1775 VDD.n15 VSS 0.0103f
C1776 VDD.n16 VSS 0.00356f
C1777 VDD.n17 VSS 0.043f
C1778 VDD.n18 VSS 0.0285f
C1779 VDD.n19 VSS 0.019f
C1780 VDD.n20 VSS 0.035f
C1781 VDD.n21 VSS 0.0359f
C1782 VDD.n22 VSS 0.019f
C1783 VDD.n23 VSS 0.035f
C1784 VDD.n24 VSS 0.0358f
C1785 VDD.n25 VSS 0.0212f
C1786 VDD.n26 VSS 0.0304f
C1787 VDD.n27 VSS 0.0283f
C1788 VDD.n28 VSS 0.0212f
C1789 VDD.n29 VSS 0.0533f
C1790 VDD.t424 VSS 0.00772f
C1791 VDD.n30 VSS 0.0895f
C1792 VDD.t420 VSS 0.042f
C1793 VDD.t12 VSS 0.00252f
C1794 VDD.n31 VSS 0.00252f
C1795 VDD.n32 VSS 0.00551f
C1796 VDD.t258 VSS 0.00614f
C1797 VDD.n33 VSS 0.00613f
C1798 VDD.n34 VSS 0.111f
C1799 VDD.t98 VSS 0.0811f
C1800 VDD.n35 VSS 0.00613f
C1801 VDD.t386 VSS 0.00614f
C1802 VDD.n36 VSS 0.00613f
C1803 VDD.n37 VSS 0.00613f
C1804 VDD.t330 VSS 0.0799f
C1805 VDD.n38 VSS 0.0381f
C1806 VDD.t97 VSS 0.00614f
C1807 VDD.n39 VSS 0.00613f
C1808 VDD.t96 VSS 0.074f
C1809 VDD.t101 VSS 0.0811f
C1810 VDD.n40 VSS 0.0381f
C1811 VDD.t48 VSS 0.00614f
C1812 VDD.t400 VSS 0.00252f
C1813 VDD.n41 VSS 0.00252f
C1814 VDD.n42 VSS 0.00551f
C1815 VDD.t47 VSS 0.074f
C1816 VDD.t399 VSS 0.0904f
C1817 VDD.t254 VSS 0.042f
C1818 VDD.n43 VSS 0.0381f
C1819 VDD.t126 VSS 0.00614f
C1820 VDD.t317 VSS 0.00252f
C1821 VDD.n44 VSS 0.00252f
C1822 VDD.n45 VSS 0.00551f
C1823 VDD.t125 VSS 0.074f
C1824 VDD.t316 VSS 0.0904f
C1825 VDD.t425 VSS 0.042f
C1826 VDD.t166 VSS 0.0738f
C1827 VDD.n46 VSS 0.0381f
C1828 VDD.t167 VSS 0.00614f
C1829 VDD.t151 VSS 0.00527f
C1830 VDD.t463 VSS 0.00399f
C1831 VDD.n47 VSS 0.0104f
C1832 VDD.n48 VSS 0.00848f
C1833 VDD.t165 VSS 0.00527f
C1834 VDD.t459 VSS 0.00399f
C1835 VDD.n49 VSS 0.0104f
C1836 VDD.n50 VSS 0.0473f
C1837 VDD.n51 VSS 0.0285f
C1838 VDD.n52 VSS 0.019f
C1839 VDD.n53 VSS 0.035f
C1840 VDD.n54 VSS 0.0359f
C1841 VDD.n55 VSS 0.019f
C1842 VDD.n56 VSS 0.035f
C1843 VDD.n57 VSS 0.0358f
C1844 VDD.n58 VSS 0.0212f
C1845 VDD.n59 VSS 0.0304f
C1846 VDD.n60 VSS 0.0283f
C1847 VDD.n61 VSS 0.0212f
C1848 VDD.n62 VSS 0.0533f
C1849 VDD.n63 VSS 0.00611f
C1850 VDD.t232 VSS 0.0542f
C1851 VDD.n64 VSS 0.057f
C1852 VDD.n65 VSS 0.00613f
C1853 VDD.t107 VSS 0.0421f
C1854 VDD.n66 VSS 0.0381f
C1855 VDD.t229 VSS 0.00252f
C1856 VDD.n67 VSS 0.00252f
C1857 VDD.n68 VSS 0.0055f
C1858 VDD.n69 VSS 0.00613f
C1859 VDD.t228 VSS 0.0418f
C1860 VDD.t24 VSS 0.0904f
C1861 VDD.t360 VSS 0.0742f
C1862 VDD.n70 VSS 0.0381f
C1863 VDD.t92 VSS 0.00612f
C1864 VDD.n71 VSS 0.00613f
C1865 VDD.t91 VSS 0.0809f
C1866 VDD.t70 VSS 0.0742f
C1867 VDD.n72 VSS 0.0381f
C1868 VDD.t289 VSS 0.00612f
C1869 VDD.n73 VSS 0.00613f
C1870 VDD.t288 VSS 0.0809f
C1871 VDD.t64 VSS 0.0742f
C1872 VDD.t27 VSS 0.0798f
C1873 VDD.n74 VSS 0.0381f
C1874 VDD.t28 VSS 0.00612f
C1875 VDD.t121 VSS 0.00613f
C1876 VDD.t93 VSS 0.0742f
C1877 VDD.n75 VSS 0.00614f
C1878 VDD.t359 VSS 0.00252f
C1879 VDD.n76 VSS 0.00252f
C1880 VDD.n77 VSS 0.00551f
C1881 VDD.n78 VSS 0.00614f
C1882 VDD.n79 VSS 0.0359f
C1883 VDD.t158 VSS 0.074f
C1884 VDD.n80 VSS 0.00574f
C1885 VDD.n81 VSS 6.07e-19
C1886 VDD.t171 VSS 0.00527f
C1887 VDD.t455 VSS 0.00399f
C1888 VDD.n82 VSS 0.0103f
C1889 VDD.n83 VSS 0.0684f
C1890 VDD.n84 VSS 0.0676f
C1891 VDD.t461 VSS 0.00398f
C1892 VDD.t157 VSS 0.00517f
C1893 VDD.n85 VSS 0.005f
C1894 VDD.n86 VSS 0.0054f
C1895 VDD.n87 VSS 8.68e-19
C1896 VDD.n88 VSS 0.00458f
C1897 VDD.n89 VSS 0.0143f
C1898 VDD.t132 VSS 0.00252f
C1899 VDD.n90 VSS 0.00252f
C1900 VDD.n91 VSS 0.00551f
C1901 VDD.n92 VSS 0.035f
C1902 VDD.n93 VSS 0.0351f
C1903 VDD.n94 VSS 0.0381f
C1904 VDD.t131 VSS 0.0418f
C1905 VDD.t122 VSS 0.0904f
C1906 VDD.t205 VSS 0.0742f
C1907 VDD.t67 VSS 0.0904f
C1908 VDD.t358 VSS 0.0418f
C1909 VDD.n95 VSS 0.0381f
C1910 VDD.n96 VSS 0.019f
C1911 VDD.n97 VSS 0.035f
C1912 VDD.n98 VSS 0.0358f
C1913 VDD.t287 VSS 0.00613f
C1914 VDD.n99 VSS 0.00614f
C1915 VDD.n100 VSS 0.0282f
C1916 VDD.n101 VSS 0.0304f
C1917 VDD.n102 VSS 0.0213f
C1918 VDD.n103 VSS 0.0381f
C1919 VDD.t286 VSS 0.0809f
C1920 VDD.t269 VSS 0.0742f
C1921 VDD.t120 VSS 0.0798f
C1922 VDD.n104 VSS 0.0381f
C1923 VDD.n105 VSS 0.0213f
C1924 VDD.n106 VSS 0.0529f
C1925 VDD.n107 VSS 0.00611f
C1926 VDD.t237 VSS 0.0542f
C1927 VDD.n108 VSS 0.057f
C1928 VDD.t236 VSS 0.00252f
C1929 VDD.n109 VSS 0.00252f
C1930 VDD.n110 VSS 0.00551f
C1931 VDD.n111 VSS 0.0198f
C1932 VDD.n112 VSS 0.00614f
C1933 VDD.t435 VSS 0.074f
C1934 VDD.n113 VSS 0.0381f
C1935 VDD.t116 VSS 0.00613f
C1936 VDD.n114 VSS 0.00611f
C1937 VDD.t115 VSS 0.0482f
C1938 VDD.t240 VSS 0.0552f
C1939 VDD.n115 VSS 0.0957f
C1940 VDD.n116 VSS 0.0147f
C1941 VDD.t438 VSS 0.0522f
C1942 VDD.n117 VSS 0.0371f
C1943 VDD.n118 VSS 0.00611f
C1944 VDD.t348 VSS 0.055f
C1945 VDD.t264 VSS 0.0544f
C1946 VDD.n119 VSS 0.0631f
C1947 VDD.n120 VSS 0.0328f
C1948 VDD.n121 VSS 0.0327f
C1949 VDD.n122 VSS 0.0333f
C1950 VDD.n123 VSS 0.0216f
C1951 VDD.n124 VSS 0.0301f
C1952 VDD.n125 VSS 0.0215f
C1953 VDD.n126 VSS 0.0422f
C1954 VDD.t117 VSS 0.0421f
C1955 VDD.n127 VSS 0.00614f
C1956 VDD.n128 VSS 0.0268f
C1957 VDD.n129 VSS 0.0213f
C1958 VDD.n130 VSS 0.00614f
C1959 VDD.t448 VSS 0.00613f
C1960 VDD.n131 VSS 0.0304f
C1961 VDD.n132 VSS 0.0282f
C1962 VDD.n133 VSS 0.0213f
C1963 VDD.n134 VSS 0.00614f
C1964 VDD.t342 VSS 0.00613f
C1965 VDD.n135 VSS 0.0304f
C1966 VDD.n136 VSS 0.0282f
C1967 VDD.t111 VSS 0.00613f
C1968 VDD.t357 VSS 0.00613f
C1969 VDD.n137 VSS 0.0666f
C1970 VDD.t172 VSS 0.0594f
C1971 VDD.t230 VSS 0.0337f
C1972 VDD.t353 VSS 0.0594f
C1973 VDD.t290 VSS 0.0594f
C1974 VDD.t198 VSS 0.0337f
C1975 VDD.t3 VSS 0.0212f
C1976 VDD.n138 VSS 0.00658f
C1977 VDD.n139 VSS 0.128f
C1978 VDD.n140 VSS 0.00614f
C1979 VDD.t231 VSS 0.00252f
C1980 VDD.n141 VSS 0.00252f
C1981 VDD.n142 VSS 0.00551f
C1982 VDD.n143 VSS 0.035f
C1983 VDD.n144 VSS 0.0359f
C1984 VDD.t199 VSS 0.00252f
C1985 VDD.n145 VSS 0.00252f
C1986 VDD.n146 VSS 0.00551f
C1987 VDD.n147 VSS 0.00614f
C1988 VDD.t340 VSS 0.00613f
C1989 VDD.n148 VSS 0.00614f
C1990 VDD.n149 VSS 0.0282f
C1991 VDD.n150 VSS 0.0304f
C1992 VDD.n151 VSS 0.0213f
C1993 VDD.n152 VSS 0.0358f
C1994 VDD.n153 VSS 0.035f
C1995 VDD.n154 VSS 0.019f
C1996 VDD.n155 VSS 0.0689f
C1997 VDD.n156 VSS 0.0823f
C1998 VDD.t449 VSS 0.0551f
C1999 VDD.t339 VSS 0.0594f
C2000 VDD.t374 VSS 0.0594f
C2001 VDD.t356 VSS 0.0595f
C2002 VDD.n157 VSS 0.0765f
C2003 VDD.n158 VSS 0.0213f
C2004 VDD.n159 VSS 0.0216f
C2005 VDD.n160 VSS 0.00574f
C2006 VDD.n161 VSS 6.07e-19
C2007 VDD.t144 VSS 0.00527f
C2008 VDD.t454 VSS 0.00399f
C2009 VDD.n162 VSS 0.0103f
C2010 VDD.n163 VSS 0.0684f
C2011 VDD.n164 VSS 0.0676f
C2012 VDD.t460 VSS 0.00398f
C2013 VDD.t161 VSS 0.00517f
C2014 VDD.n165 VSS 0.005f
C2015 VDD.n166 VSS 0.0054f
C2016 VDD.n167 VSS 8.68e-19
C2017 VDD.n168 VSS 0.00458f
C2018 VDD.n169 VSS 0.00934f
C2019 VDD.t162 VSS 0.074f
C2020 VDD.n170 VSS 0.0381f
C2021 VDD.t404 VSS 0.00252f
C2022 VDD.n171 VSS 0.00252f
C2023 VDD.n172 VSS 0.00551f
C2024 VDD.n173 VSS 0.00614f
C2025 VDD.t403 VSS 0.0418f
C2026 VDD.t296 VSS 0.0904f
C2027 VDD.t345 VSS 0.0742f
C2028 VDD.n174 VSS 0.0381f
C2029 VDD.t285 VSS 0.00252f
C2030 VDD.n175 VSS 0.00252f
C2031 VDD.n176 VSS 0.00551f
C2032 VDD.n177 VSS 0.00614f
C2033 VDD.t284 VSS 0.0418f
C2034 VDD.t248 VSS 0.0904f
C2035 VDD.t52 VSS 0.0742f
C2036 VDD.n178 VSS 0.0381f
C2037 VDD.t329 VSS 0.00613f
C2038 VDD.n179 VSS 0.00614f
C2039 VDD.t328 VSS 0.0809f
C2040 VDD.t382 VSS 0.0742f
C2041 VDD.t83 VSS 0.0798f
C2042 VDD.n180 VSS 0.0381f
C2043 VDD.t84 VSS 0.00613f
C2044 VDD.n181 VSS 0.00611f
C2045 VDD.n182 VSS 0.0193f
C2046 VDD.t212 VSS 0.00613f
C2047 VDD.t251 VSS 0.0742f
C2048 VDD.n183 VSS 0.00614f
C2049 VDD.n184 VSS 0.0359f
C2050 VDD.t304 VSS 0.0554f
C2051 VDD.t56 VSS 0.00613f
C2052 VDD.n185 VSS 0.00613f
C2053 VDD.n186 VSS 0.0438f
C2054 VDD.n187 VSS 0.0546f
C2055 VDD.t175 VSS 0.055f
C2056 VDD.t409 VSS 0.00252f
C2057 VDD.n188 VSS 0.00252f
C2058 VDD.n189 VSS 0.00551f
C2059 VDD.n190 VSS 0.0433f
C2060 VDD.t338 VSS 0.0147f
C2061 VDD.n191 VSS 0.00614f
C2062 VDD.t44 VSS 0.0421f
C2063 VDD.t402 VSS 0.00611f
C2064 VDD.t401 VSS 0.0546f
C2065 VDD.n192 VSS 0.0631f
C2066 VDD.n193 VSS 0.02f
C2067 VDD.n194 VSS 0.00614f
C2068 VDD.n195 VSS 0.0064f
C2069 VDD.t405 VSS 0.0542f
C2070 VDD.n196 VSS 0.057f
C2071 VDD.n197 VSS 0.026f
C2072 VDD.n198 VSS 0.025f
C2073 VDD.n199 VSS 0.0227f
C2074 VDD.n200 VSS 0.0381f
C2075 VDD.t408 VSS 0.0418f
C2076 VDD.t208 VSS 0.0904f
C2077 VDD.t0 VSS 0.0742f
C2078 VDD.t55 VSS 0.0809f
C2079 VDD.n201 VSS 0.0381f
C2080 VDD.t305 VSS 0.00772f
C2081 VDD.n202 VSS 0.0145f
C2082 VDD.n203 VSS 0.0149f
C2083 VDD.n204 VSS 0.0532f
C2084 VDD.n205 VSS 0.0455f
C2085 VDD.n206 VSS 0.0249f
C2086 VDD.n207 VSS 0.0371f
C2087 VDD.t337 VSS 0.0522f
C2088 VDD.n208 VSS 0.0957f
C2089 VDD.t220 VSS 0.0484f
C2090 VDD.t129 VSS 0.0738f
C2091 VDD.n209 VSS 0.0381f
C2092 VDD.n210 VSS 0.0267f
C2093 VDD.t130 VSS 0.00614f
C2094 VDD.t327 VSS 0.00613f
C2095 VDD.t325 VSS 0.00252f
C2096 VDD.n211 VSS 0.00252f
C2097 VDD.n212 VSS 0.00551f
C2098 VDD.n213 VSS 0.0236f
C2099 VDD.t223 VSS 0.0811f
C2100 VDD.n214 VSS 0.00613f
C2101 VDD.t32 VSS 0.00614f
C2102 VDD.n215 VSS 0.00613f
C2103 VDD.n216 VSS 0.0304f
C2104 VDD.t243 VSS 0.0799f
C2105 VDD.n217 VSS 0.00613f
C2106 VDD.n218 VSS 0.00613f
C2107 VDD.t176 VSS 0.0799f
C2108 VDD.n219 VSS 0.0381f
C2109 VDD.t370 VSS 0.00614f
C2110 VDD.n220 VSS 0.00613f
C2111 VDD.t369 VSS 0.074f
C2112 VDD.t85 VSS 0.0811f
C2113 VDD.n221 VSS 0.0381f
C2114 VDD.t227 VSS 0.00614f
C2115 VDD.t34 VSS 0.00252f
C2116 VDD.n222 VSS 0.00252f
C2117 VDD.n223 VSS 0.00551f
C2118 VDD.t226 VSS 0.074f
C2119 VDD.t33 VSS 0.0904f
C2120 VDD.t366 VSS 0.042f
C2121 VDD.n224 VSS 0.0381f
C2122 VDD.t336 VSS 0.00614f
C2123 VDD.t180 VSS 0.00252f
C2124 VDD.n225 VSS 0.00252f
C2125 VDD.n226 VSS 0.00551f
C2126 VDD.t335 VSS 0.074f
C2127 VDD.t179 VSS 0.0904f
C2128 VDD.t181 VSS 0.042f
C2129 VDD.t155 VSS 0.0738f
C2130 VDD.n227 VSS 0.0381f
C2131 VDD.t156 VSS 0.00658f
C2132 VDD.n228 VSS 0.0473f
C2133 VDD.n229 VSS 0.035f
C2134 VDD.n230 VSS 0.0359f
C2135 VDD.n231 VSS 0.019f
C2136 VDD.n232 VSS 0.035f
C2137 VDD.n233 VSS 0.0358f
C2138 VDD.n234 VSS 0.0212f
C2139 VDD.n235 VSS 0.0304f
C2140 VDD.n236 VSS 0.0283f
C2141 VDD.n237 VSS 0.0212f
C2142 VDD.n238 VSS 0.0579f
C2143 VDD.n239 VSS 0.0658f
C2144 VDD.t344 VSS 0.00614f
C2145 VDD.n240 VSS 0.0283f
C2146 VDD.n241 VSS 0.0212f
C2147 VDD.n242 VSS 0.0381f
C2148 VDD.t343 VSS 0.074f
C2149 VDD.t88 VSS 0.0811f
C2150 VDD.t31 VSS 0.074f
C2151 VDD.n243 VSS 0.0381f
C2152 VDD.n244 VSS 0.0212f
C2153 VDD.n245 VSS 0.0283f
C2154 VDD.n246 VSS 0.0304f
C2155 VDD.t334 VSS 0.00614f
C2156 VDD.n247 VSS 0.0268f
C2157 VDD.n248 VSS 0.0212f
C2158 VDD.n249 VSS 0.0381f
C2159 VDD.t333 VSS 0.074f
C2160 VDD.t324 VSS 0.0904f
C2161 VDD.t184 VSS 0.042f
C2162 VDD.n250 VSS 0.0381f
C2163 VDD.t219 VSS 0.00614f
C2164 VDD.t188 VSS 0.00611f
C2165 VDD.n251 VSS 0.00613f
C2166 VDD.t213 VSS 0.0645f
C2167 VDD.n252 VSS 0.0329f
C2168 VDD.t23 VSS 0.00614f
C2169 VDD.n253 VSS 0.00613f
C2170 VDD.t22 VSS 0.0589f
C2171 VDD.t321 VSS 0.0645f
C2172 VDD.n254 VSS 0.0329f
C2173 VDD.t303 VSS 0.00614f
C2174 VDD.t352 VSS 0.00252f
C2175 VDD.n255 VSS 0.00252f
C2176 VDD.n256 VSS 0.00551f
C2177 VDD.n257 VSS 0.0329f
C2178 VDD.t30 VSS 0.00614f
C2179 VDD.t217 VSS 0.00252f
C2180 VDD.n258 VSS 0.00252f
C2181 VDD.n259 VSS 0.00551f
C2182 VDD.t29 VSS 0.0589f
C2183 VDD.t216 VSS 0.0719f
C2184 VDD.t192 VSS 0.0334f
C2185 VDD.t302 VSS 0.0537f
C2186 VDD.t363 VSS 0.0334f
C2187 VDD.t351 VSS 0.0256f
C2188 VDD.n260 VSS 0.212f
C2189 VDD.t149 VSS 0.0676f
C2190 VDD.n261 VSS 0.0329f
C2191 VDD.n262 VSS 0.00158f
C2192 VDD.t464 VSS 0.00399f
C2193 VDD.t148 VSS 0.00511f
C2194 VDD.n263 VSS 0.00496f
C2195 VDD.t462 VSS 0.00399f
C2196 VDD.t154 VSS 0.00527f
C2197 VDD.n264 VSS 0.0103f
C2198 VDD.n265 VSS 0.0577f
C2199 VDD.n266 VSS 0.0754f
C2200 VDD.n267 VSS 5.1e-20
C2201 VDD.n268 VSS 0.00134f
C2202 VDD.n269 VSS 0.00548f
C2203 VDD.n270 VSS 7.31e-19
C2204 VDD.n271 VSS 6.08e-19
C2205 VDD.n272 VSS 0.00457f
C2206 VDD.t150 VSS 0.00574f
C2207 VDD.n273 VSS 0.0143f
C2208 VDD.n274 VSS 0.035f
C2209 VDD.n275 VSS 0.035f
C2210 VDD.n276 VSS 0.0359f
C2211 VDD.n277 VSS 0.019f
C2212 VDD.n278 VSS 0.035f
C2213 VDD.n279 VSS 0.0358f
C2214 VDD.n280 VSS 0.0212f
C2215 VDD.n281 VSS 0.0304f
C2216 VDD.n282 VSS 0.0283f
C2217 VDD.n283 VSS 0.0212f
C2218 VDD.n284 VSS 0.053f
C2219 VDD.n285 VSS 0.00613f
C2220 VDD.t136 VSS 0.0799f
C2221 VDD.n286 VSS 0.0381f
C2222 VDD.n287 VSS 0.00613f
C2223 VDD.n288 VSS 0.00614f
C2224 VDD.t380 VSS 0.074f
C2225 VDD.t318 VSS 0.0811f
C2226 VDD.n289 VSS 0.0381f
C2227 VDD.t444 VSS 0.074f
C2228 VDD.n290 VSS 0.0381f
C2229 VDD.t350 VSS 0.00614f
C2230 VDD.t82 VSS 0.00613f
C2231 VDD.n291 VSS 0.00613f
C2232 VDD.t81 VSS 0.0482f
C2233 VDD.t371 VSS 0.0552f
C2234 VDD.n292 VSS 0.0957f
C2235 VDD.n293 VSS 0.0077f
C2236 VDD.t349 VSS 0.074f
C2237 VDD.t299 VSS 0.0811f
C2238 VDD.n294 VSS 0.0381f
C2239 VDD.t61 VSS 0.00614f
C2240 VDD.n295 VSS 0.0147f
C2241 VDD.t394 VSS 0.0522f
C2242 VDD.n296 VSS 0.0371f
C2243 VDD.t140 VSS 0.00252f
C2244 VDD.n297 VSS 0.00252f
C2245 VDD.n298 VSS 0.00551f
C2246 VDD.t60 VSS 0.074f
C2247 VDD.t139 VSS 0.0904f
C2248 VDD.t189 VSS 0.042f
C2249 VDD.n299 VSS 0.0381f
C2250 VDD.n300 VSS 0.00611f
C2251 VDD.t432 VSS 0.055f
C2252 VDD.t441 VSS 0.0544f
C2253 VDD.n301 VSS 0.0631f
C2254 VDD.n302 VSS 0.02f
C2255 VDD.t247 VSS 0.00646f
C2256 VDD.t246 VSS 0.042f
C2257 VDD.t127 VSS 0.0543f
C2258 VDD.n303 VSS 0.057f
C2259 VDD.t128 VSS 0.0063f
C2260 VDD.n304 VSS 0.0673f
C2261 VDD.n305 VSS 0.0207f
C2262 VDD.n306 VSS 0.0227f
C2263 VDD.n307 VSS 0.0433f
C2264 VDD.n308 VSS 0.0251f
C2265 VDD.n309 VSS 0.0454f
C2266 VDD.n310 VSS 0.0533f
C2267 VDD.n311 VSS 0.0149f
C2268 VDD.n312 VSS 0.0147f
C2269 VDD.n313 VSS 0.0544f
C2270 VDD.n314 VSS 0.0438f
C2271 VDD.n315 VSS 0.0359f
C2272 VDD.n316 VSS 0.0268f
C2273 VDD.n317 VSS 0.0259f
C2274 VDD.n318 VSS 0.0359f
C2275 VDD.n319 VSS 0.0276f
C2276 VDD.t429 VSS 0.00252f
C2277 VDD.n320 VSS 0.00252f
C2278 VDD.n321 VSS 0.00551f
C2279 VDD.n322 VSS 0.0198f
C2280 VDD.n323 VSS 0.00614f
C2281 VDD.n324 VSS 0.027f
C2282 VDD.t412 VSS 0.0542f
C2283 VDD.n325 VSS 0.057f
C2284 VDD.t293 VSS 0.0421f
C2285 VDD.t314 VSS 0.0809f
C2286 VDD.n326 VSS 0.00614f
C2287 VDD.n327 VSS 0.0268f
C2288 VDD.t315 VSS 0.00613f
C2289 VDD.n328 VSS 0.00614f
C2290 VDD.t275 VSS 0.0742f
C2291 VDD.n329 VSS 0.0381f
C2292 VDD.t41 VSS 0.00613f
C2293 VDD.n330 VSS 0.00614f
C2294 VDD.t40 VSS 0.0809f
C2295 VDD.t133 VSS 0.0742f
C2296 VDD.t262 VSS 0.0798f
C2297 VDD.n331 VSS 0.0381f
C2298 VDD.t263 VSS 0.00613f
C2299 VDD.t43 VSS 0.00613f
C2300 VDD.n332 VSS 0.0666f
C2301 VDD.t145 VSS 0.0594f
C2302 VDD.t410 VSS 0.0337f
C2303 VDD.t281 VSS 0.0594f
C2304 VDD.t195 VSS 0.0594f
C2305 VDD.t267 VSS 0.0337f
C2306 VDD.t272 VSS 0.0212f
C2307 VDD.n333 VSS 0.00658f
C2308 VDD.n334 VSS 0.128f
C2309 VDD.n335 VSS 0.00614f
C2310 VDD.t411 VSS 0.00252f
C2311 VDD.n336 VSS 0.00252f
C2312 VDD.n337 VSS 0.00551f
C2313 VDD.n338 VSS 0.035f
C2314 VDD.n339 VSS 0.0359f
C2315 VDD.t268 VSS 0.00252f
C2316 VDD.n340 VSS 0.00252f
C2317 VDD.n341 VSS 0.00551f
C2318 VDD.n342 VSS 0.00614f
C2319 VDD.t39 VSS 0.00613f
C2320 VDD.n343 VSS 0.00614f
C2321 VDD.n344 VSS 0.0282f
C2322 VDD.n345 VSS 0.0304f
C2323 VDD.n346 VSS 0.0213f
C2324 VDD.n347 VSS 0.0358f
C2325 VDD.n348 VSS 0.035f
C2326 VDD.n349 VSS 0.019f
C2327 VDD.n350 VSS 0.0689f
C2328 VDD.n351 VSS 0.0823f
C2329 VDD.t311 VSS 0.0551f
C2330 VDD.t38 VSS 0.0594f
C2331 VDD.t387 VSS 0.0594f
C2332 VDD.t42 VSS 0.0595f
C2333 VDD.n352 VSS 0.0765f
C2334 VDD.n353 VSS 0.0213f
C2335 VDD.n354 VSS 0.0578f
C2336 VDD.n355 VSS 0.0657f
C2337 VDD.n356 VSS 0.0213f
C2338 VDD.n357 VSS 0.0282f
C2339 VDD.n358 VSS 0.0304f
C2340 VDD.n359 VSS 0.0213f
C2341 VDD.n360 VSS 0.0282f
C2342 VDD.n361 VSS 0.0304f
C2343 VDD.n362 VSS 0.0213f
C2344 VDD.n363 VSS 0.0381f
C2345 VDD.t57 VSS 0.0742f
C2346 VDD.t259 VSS 0.0904f
C2347 VDD.t428 VSS 0.0418f
C2348 VDD.n364 VSS 0.0381f
C2349 VDD.n365 VSS 0.0141f
C2350 VDD.n366 VSS 0.0479f
C2351 VDD.n367 VSS 0.039f
C2352 VDD.t381 VSS 0.00632f
C2353 VDD.n368 VSS 0.0483f
C2354 VDD.n369 VSS 0.0318f
C2355 VDD.n370 VSS 0.0531f
C2356 VDD.n371 VSS 0.0717f
C2357 VDD.n372 VSS 0.0422f
C2358 VDD.t187 VSS 0.0543f
C2359 VDD.t218 VSS 0.042f
C2360 VDD.n373 VSS 0.057f
C2361 VDD.n374 VSS 0.0588f
C2362 VDD.n375 VSS 0.027f
C2363 VDD.n376 VSS 0.0451f
C2364 VDD.n377 VSS 0.00589f
C2365 VDD.n378 VSS 0.0139f
C2366 VDD.n379 VSS 0.0608f
C2367 VDD.n380 VSS 0.0275f
C2368 VDD.n381 VSS 0.0359f
C2369 VDD.n382 VSS 0.026f
C2370 VDD.n383 VSS 0.0381f
C2371 VDD.t326 VSS 0.0809f
C2372 VDD.t104 VSS 0.0742f
C2373 VDD.t211 VSS 0.0798f
C2374 VDD.n384 VSS 0.0381f
C2375 VDD.n385 VSS 0.0213f
C2376 VDD.n386 VSS 0.0311f
C2377 VDD.n387 VSS 0.0434f
C2378 VDD.n388 VSS 0.0543f
C2379 VDD.n389 VSS 0.0213f
C2380 VDD.n390 VSS 0.0282f
C2381 VDD.n391 VSS 0.0304f
C2382 VDD.n392 VSS 0.0213f
C2383 VDD.n393 VSS 0.0358f
C2384 VDD.n394 VSS 0.035f
C2385 VDD.n395 VSS 0.019f
C2386 VDD.n396 VSS 0.0359f
C2387 VDD.n397 VSS 0.035f
C2388 VDD.n398 VSS 0.019f
C2389 VDD.n399 VSS 0.0684f
C2390 VDD.n400 VSS 0.0855f
C2391 VDD.n401 VSS 0.0647f
C2392 VDD.n402 VSS 0.0213f
C2393 VDD.t110 VSS 0.0798f
C2394 VDD.n403 VSS 0.0381f
C2395 VDD.t377 VSS 0.0742f
C2396 VDD.t341 VSS 0.0809f
C2397 VDD.n404 VSS 0.0381f
C2398 VDD.t6 VSS 0.0742f
C2399 VDD.t447 VSS 0.0809f
C2400 VDD.n405 VSS 0.0381f
C2401 VDD.t35 VSS 0.0742f
C2402 VDD.t112 VSS 0.0904f
C2403 VDD.t235 VSS 0.0418f
C2404 VDD.n406 VSS 0.0381f
C2405 VDD.n407 VSS 0.0141f
C2406 VDD.n408 VSS 0.0469f
C2407 VDD.n409 VSS 0.00634f
C2408 VDD.n410 VSS 0.0352f
C2409 VDD.n411 VSS 0.0271f
C2410 VDD.n412 VSS 0.0491f
C2411 VDD.n413 VSS 0.0319f
C2412 VDD.n414 VSS 0.0223f
C2413 VDD.n415 VSS 0.0303f
C2414 VDD.n416 VSS 0.0327f
C2415 VDD.n417 VSS 0.0223f
C2416 VDD.n418 VSS 0.0303f
C2417 VDD.n419 VSS 0.0327f
C2418 VDD.n420 VSS 0.0223f
C2419 VDD.n421 VSS 0.0286f
C2420 VDD.n422 VSS 0.0271f
C2421 VDD.n423 VSS 0.0198f
C2422 VDD.n424 VSS 0.035f
C2423 VDD.n425 VSS 0.224f
C2424 VDD.n426 VSS 0.548f
C2425 VDD.n427 VSS 0.108f
C2426 VDD.t9 VSS 0.0799f
C2427 VDD.t385 VSS 0.074f
C2428 VDD.n428 VSS 0.0381f
C2429 VDD.n429 VSS 0.0566f
C2430 VDD.n430 VSS 0.1f
C2431 VDD.n431 VSS 0.111f
C2432 VDD.t398 VSS 0.00614f
C2433 VDD.n432 VSS 0.1f
C2434 VDD.n433 VSS 0.0566f
C2435 VDD.n434 VSS 0.0381f
C2436 VDD.t397 VSS 0.074f
C2437 VDD.t49 VSS 0.0811f
C2438 VDD.t11 VSS 0.0904f
C2439 VDD.t257 VSS 0.074f
C2440 VDD.n435 VSS 0.0381f
C2441 VDD.n436 VSS 0.0566f
C2442 VDD.n437 VSS 0.0926f
C2443 VDD.n438 VSS 0.0963f
C2444 VDD.t153 VSS 0.00614f
C2445 VDD.n439 VSS 0.12f
C2446 VDD.n440 VSS 0.0457f
C2447 VDD.n441 VSS 0.0381f
C2448 VDD.t152 VSS 0.042f
C2449 VDD.t423 VSS 0.0542f
C2450 VDD.n442 VSS 0.057f
C2451 VDD.n443 VSS 0.0898f
C2452 VDD.n444 VSS 0.109f
C2453 VDD.t431 VSS 0.00614f
C2454 VDD.n445 VSS 0.101f
C2455 VDD.n446 VSS 0.0568f
C2456 VDD.n447 VSS 0.0381f
C2457 VDD.t430 VSS 0.074f
C2458 VDD.t78 VSS 0.0811f
C2459 VDD.t392 VSS 0.074f
C2460 VDD.n448 VSS 0.0381f
C2461 VDD.n449 VSS 0.0568f
C2462 VDD.n450 VSS 0.101f
C2463 VDD.n451 VSS 0.112f
C2464 VDD.t74 VSS 0.00614f
C2465 VDD.t307 VSS 0.00252f
C2466 VDD.n452 VSS 0.00252f
C2467 VDD.n453 VSS 0.00551f
C2468 VDD.n454 VSS 0.0966f
C2469 VDD.n455 VSS 0.0929f
C2470 VDD.n456 VSS 0.0568f
C2471 VDD.n457 VSS 0.0381f
C2472 VDD.t73 VSS 0.074f
C2473 VDD.t306 VSS 0.0904f
C2474 VDD.t16 VSS 0.042f
C2475 VDD.t142 VSS 0.042f
C2476 VDD.n458 VSS 0.0381f
C2477 VDD.n459 VSS 0.0458f
C2478 VDD.n460 VSS 0.121f
C2479 VDD.n461 VSS 0.0898f
C2480 VDD.t14 VSS 0.0542f
C2481 VDD.n462 VSS 0.057f
.ends

