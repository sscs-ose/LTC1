magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2208 -2120 2348 2720
<< nwell >>
rect -208 -120 348 720
<< mvpmos >>
rect 0 0 140 600
<< mvpdiff >>
rect -88 587 0 600
rect -88 541 -75 587
rect -29 541 0 587
rect -88 482 0 541
rect -88 436 -75 482
rect -29 436 0 482
rect -88 377 0 436
rect -88 331 -75 377
rect -29 331 0 377
rect -88 271 0 331
rect -88 225 -75 271
rect -29 225 0 271
rect -88 165 0 225
rect -88 119 -75 165
rect -29 119 0 165
rect -88 59 0 119
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 587 228 600
rect 140 541 169 587
rect 215 541 228 587
rect 140 482 228 541
rect 140 436 169 482
rect 215 436 228 482
rect 140 377 228 436
rect 140 331 169 377
rect 215 331 228 377
rect 140 271 228 331
rect 140 225 169 271
rect 215 225 228 271
rect 140 165 228 225
rect 140 119 169 165
rect 215 119 228 165
rect 140 59 228 119
rect 140 13 169 59
rect 215 13 228 59
rect 140 0 228 13
<< mvpdiffc >>
rect -75 541 -29 587
rect -75 436 -29 482
rect -75 331 -29 377
rect -75 225 -29 271
rect -75 119 -29 165
rect -75 13 -29 59
rect 169 541 215 587
rect 169 436 215 482
rect 169 331 215 377
rect 169 225 215 271
rect 169 119 215 165
rect 169 13 215 59
<< polysilicon >>
rect 0 600 140 644
rect 0 -44 140 0
<< metal1 >>
rect -75 587 -29 600
rect -75 482 -29 541
rect -75 377 -29 436
rect -75 271 -29 331
rect -75 165 -29 225
rect -75 59 -29 119
rect -75 0 -29 13
rect 169 587 215 600
rect 169 482 215 541
rect 169 377 215 436
rect 169 271 215 331
rect 169 165 215 225
rect 169 59 215 119
rect 169 0 215 13
<< labels >>
rlabel metal1 192 300 192 300 4 D
rlabel metal1 -52 300 -52 300 4 S
<< end >>
