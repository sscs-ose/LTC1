magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7545 -2245 7545 2245
<< psubdiff >>
rect -5545 223 5545 245
rect -5545 -223 -5523 223
rect 5523 -223 5545 223
rect -5545 -245 5545 -223
<< psubdiffcont >>
rect -5523 -223 5523 223
<< metal1 >>
rect -5534 223 5534 234
rect -5534 -223 -5523 223
rect 5523 -223 5534 223
rect -5534 -234 5534 -223
<< end >>
