magic
tech gf180mcuC
magscale 1 10
timestamp 1699882188
<< nwell >>
rect -284 -1136 284 1136
<< nsubdiff >>
rect -260 1040 260 1112
rect -260 -1040 -188 1040
rect 188 -1040 260 1040
rect -260 -1112 260 -1040
<< polysilicon >>
rect -100 939 100 952
rect -100 893 -87 939
rect 87 893 100 939
rect -100 850 100 893
rect -100 -893 100 -850
rect -100 -939 -87 -893
rect 87 -939 100 -893
rect -100 -952 100 -939
<< polycontact >>
rect -87 893 87 939
rect -87 -939 87 -893
<< ppolyres >>
rect -100 -850 100 850
<< metal1 >>
rect -98 893 -87 939
rect 87 893 98 939
rect -98 -939 -87 -893
rect 87 -939 98 -893
<< properties >>
string FIXED_BBOX -224 -1076 224 1076
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 8.5 m 1 nx 1 wmin 0.80 lmin 1.00 rho 315 val 2.879k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
