** sch_path: /home/shahid/GF180Projects/GF_INV/Xschem/nmos_char_dc.sch
**.subckt nmos_char_dc
XM1 d g GND GND nfet_03v3 L=.28u W=.3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
VGS g GND DC{vgs}
.save i(vgs)
VDS d GND DC{vds}
.save i(vds)
**** begin user architecture code



*Parameters
.param vds = 200m
.param vgs = 1.2

.options TEMP = 50.0

*Models

*Data to save
.save all  @M.xm1.m0[id]  @M.xm1.m0[vds]  @M.xm1.m0[vgs]  @M.xm1.m0[vth]  @M.xm1.m0[cgg]  @M.xm1.m0[cgs]  @M.xm1.m0[gds]  @M.xm1.m0[gm]  @M.xm1.m0[vdsat]

*Simulation
.control

dc VDS 0 3.3 0.01
setplot dc1
plot @M.xm1.m0[id] ylabel Id xlabel Vds
set filetype = binary
write nmos_char_dc_1.raw

reset
dc VGS 0 3.3 0.01
setplot dc2
plot @M.xm1.m0[id] ylabel Id xlabel Vgs
set filetype = binary
write nmos_char_dc_2.raw

reset
op
save all
set filetype = binary
write nmos_char_dc.raw

.endc
.end



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
