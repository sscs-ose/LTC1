* NGSPICE file created from NOR_Layout.ext - technology: gf180mcuC

.subckt pmos_3p3_MEVUAR a_n196_n100# a_n52_n100# w_n282_n230# a_108_n100# a_52_n144#
+ a_n108_n144#
X0 a_n52_n100# a_n108_n144# a_n196_n100# w_n282_n230# pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1 a_108_n100# a_52_n144# a_n52_n100# w_n282_n230# pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
.ends

.subckt nmos_3p3_GGGST2 a_n28_n94# a_n116_n50# a_28_n50# VSUBS
X0 a_28_n50# a_n28_n94# a_n116_n50# VSUBS nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
.ends

.subckt NOR_Layout A B OUT VDD VSS
Xpmos_3p3_MEVUAR_0 m1_99_317# OUT VDD m1_99_317# B B pmos_3p3_MEVUAR
Xpmos_3p3_MEVUAR_1 m1_99_317# VDD VDD m1_99_317# A A pmos_3p3_MEVUAR
Xnmos_3p3_GGGST2_0 B OUT VSS VSS nmos_3p3_GGGST2
Xnmos_3p3_GGGST2_1 A VSS OUT VSS nmos_3p3_GGGST2
.ends

