magic
tech gf180mcuC
magscale 1 10
timestamp 1691396512
<< pwell >>
rect -460 -872 460 872
<< nmos >>
rect -348 504 -292 804
rect -188 504 -132 804
rect -28 504 28 804
rect 132 504 188 804
rect 292 504 348 804
rect -348 68 -292 368
rect -188 68 -132 368
rect -28 68 28 368
rect 132 68 188 368
rect 292 68 348 368
rect -348 -368 -292 -68
rect -188 -368 -132 -68
rect -28 -368 28 -68
rect 132 -368 188 -68
rect 292 -368 348 -68
rect -348 -804 -292 -504
rect -188 -804 -132 -504
rect -28 -804 28 -504
rect 132 -804 188 -504
rect 292 -804 348 -504
<< ndiff >>
rect -436 791 -348 804
rect -436 517 -423 791
rect -377 517 -348 791
rect -436 504 -348 517
rect -292 791 -188 804
rect -292 517 -263 791
rect -217 517 -188 791
rect -292 504 -188 517
rect -132 791 -28 804
rect -132 517 -103 791
rect -57 517 -28 791
rect -132 504 -28 517
rect 28 791 132 804
rect 28 517 57 791
rect 103 517 132 791
rect 28 504 132 517
rect 188 791 292 804
rect 188 517 217 791
rect 263 517 292 791
rect 188 504 292 517
rect 348 791 436 804
rect 348 517 377 791
rect 423 517 436 791
rect 348 504 436 517
rect -436 355 -348 368
rect -436 81 -423 355
rect -377 81 -348 355
rect -436 68 -348 81
rect -292 355 -188 368
rect -292 81 -263 355
rect -217 81 -188 355
rect -292 68 -188 81
rect -132 355 -28 368
rect -132 81 -103 355
rect -57 81 -28 355
rect -132 68 -28 81
rect 28 355 132 368
rect 28 81 57 355
rect 103 81 132 355
rect 28 68 132 81
rect 188 355 292 368
rect 188 81 217 355
rect 263 81 292 355
rect 188 68 292 81
rect 348 355 436 368
rect 348 81 377 355
rect 423 81 436 355
rect 348 68 436 81
rect -436 -81 -348 -68
rect -436 -355 -423 -81
rect -377 -355 -348 -81
rect -436 -368 -348 -355
rect -292 -81 -188 -68
rect -292 -355 -263 -81
rect -217 -355 -188 -81
rect -292 -368 -188 -355
rect -132 -81 -28 -68
rect -132 -355 -103 -81
rect -57 -355 -28 -81
rect -132 -368 -28 -355
rect 28 -81 132 -68
rect 28 -355 57 -81
rect 103 -355 132 -81
rect 28 -368 132 -355
rect 188 -81 292 -68
rect 188 -355 217 -81
rect 263 -355 292 -81
rect 188 -368 292 -355
rect 348 -81 436 -68
rect 348 -355 377 -81
rect 423 -355 436 -81
rect 348 -368 436 -355
rect -436 -517 -348 -504
rect -436 -791 -423 -517
rect -377 -791 -348 -517
rect -436 -804 -348 -791
rect -292 -517 -188 -504
rect -292 -791 -263 -517
rect -217 -791 -188 -517
rect -292 -804 -188 -791
rect -132 -517 -28 -504
rect -132 -791 -103 -517
rect -57 -791 -28 -517
rect -132 -804 -28 -791
rect 28 -517 132 -504
rect 28 -791 57 -517
rect 103 -791 132 -517
rect 28 -804 132 -791
rect 188 -517 292 -504
rect 188 -791 217 -517
rect 263 -791 292 -517
rect 188 -804 292 -791
rect 348 -517 436 -504
rect 348 -791 377 -517
rect 423 -791 436 -517
rect 348 -804 436 -791
<< ndiffc >>
rect -423 517 -377 791
rect -263 517 -217 791
rect -103 517 -57 791
rect 57 517 103 791
rect 217 517 263 791
rect 377 517 423 791
rect -423 81 -377 355
rect -263 81 -217 355
rect -103 81 -57 355
rect 57 81 103 355
rect 217 81 263 355
rect 377 81 423 355
rect -423 -355 -377 -81
rect -263 -355 -217 -81
rect -103 -355 -57 -81
rect 57 -355 103 -81
rect 217 -355 263 -81
rect 377 -355 423 -81
rect -423 -791 -377 -517
rect -263 -791 -217 -517
rect -103 -791 -57 -517
rect 57 -791 103 -517
rect 217 -791 263 -517
rect 377 -791 423 -517
<< polysilicon >>
rect -348 804 -292 848
rect -188 804 -132 848
rect -28 804 28 848
rect 132 804 188 848
rect 292 804 348 848
rect -348 460 -292 504
rect -188 460 -132 504
rect -28 460 28 504
rect 132 460 188 504
rect 292 460 348 504
rect -348 368 -292 412
rect -188 368 -132 412
rect -28 368 28 412
rect 132 368 188 412
rect 292 368 348 412
rect -348 24 -292 68
rect -188 24 -132 68
rect -28 24 28 68
rect 132 24 188 68
rect 292 24 348 68
rect -348 -68 -292 -24
rect -188 -68 -132 -24
rect -28 -68 28 -24
rect 132 -68 188 -24
rect 292 -68 348 -24
rect -348 -412 -292 -368
rect -188 -412 -132 -368
rect -28 -412 28 -368
rect 132 -412 188 -368
rect 292 -412 348 -368
rect -348 -504 -292 -460
rect -188 -504 -132 -460
rect -28 -504 28 -460
rect 132 -504 188 -460
rect 292 -504 348 -460
rect -348 -848 -292 -804
rect -188 -848 -132 -804
rect -28 -848 28 -804
rect 132 -848 188 -804
rect 292 -848 348 -804
<< metal1 >>
rect -423 791 -377 802
rect -423 506 -377 517
rect -263 791 -217 802
rect -263 506 -217 517
rect -103 791 -57 802
rect -103 506 -57 517
rect 57 791 103 802
rect 57 506 103 517
rect 217 791 263 802
rect 217 506 263 517
rect 377 791 423 802
rect 377 506 423 517
rect -423 355 -377 366
rect -423 70 -377 81
rect -263 355 -217 366
rect -263 70 -217 81
rect -103 355 -57 366
rect -103 70 -57 81
rect 57 355 103 366
rect 57 70 103 81
rect 217 355 263 366
rect 217 70 263 81
rect 377 355 423 366
rect 377 70 423 81
rect -423 -81 -377 -70
rect -423 -366 -377 -355
rect -263 -81 -217 -70
rect -263 -366 -217 -355
rect -103 -81 -57 -70
rect -103 -366 -57 -355
rect 57 -81 103 -70
rect 57 -366 103 -355
rect 217 -81 263 -70
rect 217 -366 263 -355
rect 377 -81 423 -70
rect 377 -366 423 -355
rect -423 -517 -377 -506
rect -423 -802 -377 -791
rect -263 -517 -217 -506
rect -263 -802 -217 -791
rect -103 -517 -57 -506
rect -103 -802 -57 -791
rect 57 -517 103 -506
rect 57 -802 103 -791
rect 217 -517 263 -506
rect 217 -802 263 -791
rect 377 -517 423 -506
rect 377 -802 423 -791
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 1.5 l 0.280 m 4 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
