magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2038 -2535 2038 2535
<< metal2 >>
rect -38 525 38 535
rect -38 469 -28 525
rect 28 469 38 525
rect -38 383 38 469
rect -38 327 -28 383
rect 28 327 38 383
rect -38 241 38 327
rect -38 185 -28 241
rect 28 185 38 241
rect -38 99 38 185
rect -38 43 -28 99
rect 28 43 38 99
rect -38 -43 38 43
rect -38 -99 -28 -43
rect 28 -99 38 -43
rect -38 -185 38 -99
rect -38 -241 -28 -185
rect 28 -241 38 -185
rect -38 -327 38 -241
rect -38 -383 -28 -327
rect 28 -383 38 -327
rect -38 -469 38 -383
rect -38 -525 -28 -469
rect 28 -525 38 -469
rect -38 -535 38 -525
<< via2 >>
rect -28 469 28 525
rect -28 327 28 383
rect -28 185 28 241
rect -28 43 28 99
rect -28 -99 28 -43
rect -28 -241 28 -185
rect -28 -383 28 -327
rect -28 -525 28 -469
<< metal3 >>
rect -38 525 38 535
rect -38 469 -28 525
rect 28 469 38 525
rect -38 383 38 469
rect -38 327 -28 383
rect 28 327 38 383
rect -38 241 38 327
rect -38 185 -28 241
rect 28 185 38 241
rect -38 99 38 185
rect -38 43 -28 99
rect 28 43 38 99
rect -38 -43 38 43
rect -38 -99 -28 -43
rect 28 -99 38 -43
rect -38 -185 38 -99
rect -38 -241 -28 -185
rect 28 -241 38 -185
rect -38 -327 38 -241
rect -38 -383 -28 -327
rect 28 -383 38 -327
rect -38 -469 38 -383
rect -38 -525 -28 -469
rect 28 -525 38 -469
rect -38 -535 38 -525
<< end >>
