magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1127 -1073 1127 1073
<< metal1 >>
rect -127 67 127 73
rect -127 41 -121 67
rect -95 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 95 67
rect 121 41 127 67
rect -127 13 127 41
rect -127 -13 -121 13
rect -95 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 95 13
rect 121 -13 127 13
rect -127 -41 127 -13
rect -127 -67 -121 -41
rect -95 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 95 -41
rect 121 -67 127 -41
rect -127 -73 127 -67
<< via1 >>
rect -121 41 -95 67
rect -67 41 -41 67
rect -13 41 13 67
rect 41 41 67 67
rect 95 41 121 67
rect -121 -13 -95 13
rect -67 -13 -41 13
rect -13 -13 13 13
rect 41 -13 67 13
rect 95 -13 121 13
rect -121 -67 -95 -41
rect -67 -67 -41 -41
rect -13 -67 13 -41
rect 41 -67 67 -41
rect 95 -67 121 -41
<< metal2 >>
rect -127 67 127 73
rect -127 41 -121 67
rect -95 41 -67 67
rect -41 41 -13 67
rect 13 41 41 67
rect 67 41 95 67
rect 121 41 127 67
rect -127 13 127 41
rect -127 -13 -121 13
rect -95 -13 -67 13
rect -41 -13 -13 13
rect 13 -13 41 13
rect 67 -13 95 13
rect 121 -13 127 13
rect -127 -41 127 -13
rect -127 -67 -121 -41
rect -95 -67 -67 -41
rect -41 -67 -13 -41
rect 13 -67 41 -41
rect 67 -67 95 -41
rect 121 -67 127 -41
rect -127 -73 127 -67
<< end >>
