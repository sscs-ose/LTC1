magic
tech gf180mcuC
magscale 1 10
timestamp 1698649173
<< nwell >>
rect -367 1688 1644 1873
rect 405 267 482 345
<< psubdiff >>
rect -337 -767 1614 -737
rect -337 -821 -124 -767
rect 37 -821 97 -767
rect 258 -821 318 -767
rect 479 -821 539 -767
rect 700 -821 760 -767
rect 921 -821 981 -767
rect 1142 -821 1202 -767
rect 1363 -821 1423 -767
rect 1584 -821 1614 -767
rect -337 -851 1614 -821
<< nsubdiff >>
rect -343 1813 1614 1843
rect -343 1759 -124 1813
rect 37 1759 97 1813
rect 258 1759 318 1813
rect 479 1759 539 1813
rect 700 1759 760 1813
rect 921 1759 981 1813
rect 1142 1759 1202 1813
rect 1363 1759 1423 1813
rect 1584 1759 1614 1813
rect -343 1729 1614 1759
<< psubdiffcont >>
rect -124 -821 37 -767
rect 97 -821 258 -767
rect 318 -821 479 -767
rect 539 -821 700 -767
rect 760 -821 921 -767
rect 981 -821 1142 -767
rect 1202 -821 1363 -767
rect 1423 -821 1584 -767
<< nsubdiffcont >>
rect -124 1759 37 1813
rect 97 1759 258 1813
rect 318 1759 479 1813
rect 539 1759 700 1813
rect 760 1759 921 1813
rect 981 1759 1142 1813
rect 1202 1759 1363 1813
rect 1423 1759 1584 1813
<< polysilicon >>
rect -193 1266 -137 1316
rect 406 1314 481 1326
rect 211 1266 267 1314
rect 406 1313 1470 1314
rect 406 1267 421 1313
rect 467 1267 1470 1313
rect 406 1266 1470 1267
rect 406 1252 481 1266
rect -193 930 -137 980
rect 406 978 481 990
rect 211 930 267 978
rect 406 977 1470 978
rect 406 931 421 977
rect 467 931 1470 977
rect 406 930 1470 931
rect 406 916 481 930
rect -193 594 -137 644
rect 406 642 481 654
rect 211 594 267 642
rect 406 641 1470 642
rect 406 595 421 641
rect 467 595 1470 641
rect 406 594 1470 595
rect 406 580 481 594
rect -193 107 -137 350
rect -437 90 -137 107
rect -437 44 -416 90
rect -370 44 -318 90
rect -272 44 -220 90
rect -174 44 -137 90
rect 211 89 267 336
rect 614 279 670 309
rect 774 279 830 309
rect 934 279 990 309
rect 1094 279 1150 310
rect 1254 279 1310 309
rect 1414 279 1470 310
rect 614 229 1471 279
rect -437 27 -137 44
rect -193 -11 -137 27
rect 42 76 267 89
rect 42 68 163 76
rect 42 22 56 68
rect 104 30 163 68
rect 209 30 267 76
rect 104 22 267 30
rect 42 17 267 22
rect 42 9 118 17
rect 211 12 267 17
rect -193 -325 -137 -275
rect 240 -276 670 -272
rect 211 -324 1470 -276
rect 240 -328 670 -324
rect 211 -644 1469 -588
<< polycontact >>
rect 421 1267 467 1313
rect 421 931 467 977
rect 421 595 467 641
rect -416 44 -370 90
rect -318 44 -272 90
rect -220 44 -174 90
rect 56 22 104 68
rect 163 30 209 76
<< metal1 >>
rect -367 1813 1644 1873
rect -367 1759 -124 1813
rect 37 1759 97 1813
rect 258 1759 318 1813
rect 479 1759 539 1813
rect 700 1759 760 1813
rect 921 1759 981 1813
rect 1142 1759 1202 1813
rect 1363 1759 1423 1813
rect 1584 1759 1644 1813
rect -367 1699 1644 1759
rect -268 352 -222 1699
rect -439 90 -163 107
rect -439 44 -416 90
rect -370 44 -318 90
rect -272 44 -220 90
rect -174 44 -163 90
rect -439 27 -163 44
rect -108 86 -62 1556
rect 136 1545 182 1699
rect 539 1602 1545 1650
rect 539 1544 585 1602
rect 859 1545 905 1602
rect 1179 1545 1225 1602
rect 1499 1545 1545 1602
rect 136 537 182 1371
rect 296 1312 342 1371
rect 406 1313 481 1326
rect 406 1312 421 1313
rect 296 1267 421 1312
rect 467 1267 481 1313
rect 296 1266 481 1267
rect 296 976 342 1266
rect 406 1252 481 1266
rect 406 977 481 990
rect 406 976 421 977
rect 296 931 421 976
rect 467 931 481 977
rect 296 930 481 931
rect 296 640 342 930
rect 406 916 481 930
rect 406 641 481 654
rect 406 640 421 641
rect 296 595 421 640
rect 467 595 481 641
rect 296 594 481 595
rect 296 537 342 594
rect 406 580 481 594
rect 539 537 585 1371
rect 699 1370 744 1371
rect 699 1191 745 1370
rect 699 884 745 1064
rect 699 565 745 700
rect 698 519 745 565
rect 859 519 905 1372
rect 1019 526 1065 1379
rect 1179 533 1225 1386
rect 1339 530 1385 1383
rect 1499 530 1545 1383
rect 42 86 236 89
rect -108 76 236 86
rect -108 68 163 76
rect -108 23 56 68
rect -268 -707 -222 -34
rect -108 -566 -62 23
rect 42 22 56 23
rect 104 30 163 68
rect 209 30 236 76
rect 104 22 236 30
rect 42 17 236 22
rect 42 9 118 17
rect 296 -45 342 363
rect 405 333 482 345
rect 405 279 419 333
rect 473 329 482 333
rect 539 329 585 363
rect 473 279 585 329
rect 405 221 585 279
rect 699 306 745 363
rect 1018 306 1065 363
rect 1338 306 1385 363
rect 699 304 1385 306
rect 699 229 1724 304
rect 699 227 1385 229
rect 405 162 415 221
rect 474 162 585 221
rect 405 149 585 162
rect 539 -45 585 149
rect 1289 122 1385 227
rect 699 13 1385 122
rect 699 -45 745 13
rect 1019 -46 1065 13
rect 1339 -45 1385 13
rect 136 -381 182 -219
rect 296 -381 342 -219
rect 539 -381 585 -219
rect 699 -370 745 -219
rect 859 -381 905 -219
rect 1019 -381 1065 -219
rect 1179 -381 1225 -219
rect 1339 -381 1385 -219
rect 1499 -381 1545 -219
rect 136 -707 182 -555
rect 539 -613 585 -554
rect 859 -613 905 -555
rect 1179 -613 1225 -555
rect 1499 -613 1545 -555
rect 539 -661 1545 -613
rect -367 -767 1644 -707
rect -367 -821 -124 -767
rect 37 -821 97 -767
rect 258 -821 318 -767
rect 479 -821 539 -767
rect 700 -821 760 -767
rect 921 -821 981 -767
rect 1142 -821 1202 -767
rect 1363 -821 1423 -767
rect 1584 -821 1644 -767
rect -367 -881 1644 -821
<< via1 >>
rect 419 279 473 333
rect 415 162 474 221
<< metal2 >>
rect 405 334 482 345
rect -432 333 482 334
rect -432 279 419 333
rect 473 279 482 333
rect -432 221 482 279
rect -432 162 415 221
rect 474 162 482 221
rect -432 158 482 162
rect 405 149 482 158
use nmos_3p3_CU6RT2  nmos_3p3_CU6RT2_0
timestamp 1690971400
transform 1 0 1042 0 1 -300
box -540 -336 540 336
use nmos_3p3_K66RT2  nmos_3p3_K66RT2_1
timestamp 1690971400
transform 1 0 239 0 1 -300
box -140 -336 140 336
use nmos_3p3_K66RT2  nmos_3p3_K66RT2_2
timestamp 1690971400
transform 1 0 -165 0 1 -300
box -140 -336 140 336
use pmos_3p3_MENMAR  pmos_3p3_MENMAR_0
timestamp 1690971400
transform 1 0 1042 0 1 954
box -602 -734 602 734
use pmos_3p3_MNHNAR  pmos_3p3_MNHNAR_0
timestamp 1690971400
transform 1 0 -165 0 1 954
box -202 -734 202 734
use pmos_3p3_MNHNAR  pmos_3p3_MNHNAR_1
timestamp 1690971400
transform 1 0 239 0 1 954
box -202 -734 202 734
<< labels >>
flabel metal1 1624 282 1624 282 0 FreeSans 800 0 0 0 B
port 12 nsew
flabel nsubdiffcont 842 1781 842 1781 0 FreeSans 800 0 0 0 VDD
port 13 nsew
flabel psubdiffcont 833 -798 833 -798 0 FreeSans 800 0 0 0 VSS
port 14 nsew
flabel metal2 -409 257 -409 257 0 FreeSans 1600 0 0 0 A
port 16 nsew
flabel metal1 -438 84 -438 84 0 FreeSans 1600 0 0 0 CLK
port 18 nsew
<< end >>
