magic
tech gf180mcuC
magscale 1 10
timestamp 1694669839
<< error_s >>
rect 38878 5623 38890 5635
rect 38998 5623 39010 5635
rect 39259 5623 39271 5635
rect 39381 5623 39393 5635
rect 38866 5611 38878 5623
rect 39010 5611 39022 5623
rect 39247 5611 39259 5623
rect 39393 5611 39405 5623
rect 38866 5565 38878 5577
rect 39010 5565 39022 5577
rect 38878 5553 38890 5565
rect 38998 5553 39010 5565
rect 39247 5563 39259 5575
rect 39393 5563 39405 5575
rect 39259 5551 39271 5563
rect 39381 5551 39393 5563
<< nwell >>
rect 43378 2071 43473 2203
<< metal1 >>
rect 41644 12213 42163 12279
rect 34910 12114 35109 12141
rect 34910 11960 34943 12114
rect 35080 11960 35109 12114
rect 34910 11930 35109 11960
rect 35173 12121 35372 12144
rect 35173 11965 35195 12121
rect 35347 11965 35372 12121
rect 35173 11931 35372 11965
rect 35500 12114 35699 12142
rect 35500 11961 35531 12114
rect 35675 11961 35699 12114
rect 35500 11929 35699 11961
rect 41644 11933 41698 12213
rect 42092 11933 42163 12213
rect 41644 11850 42163 11933
rect 17816 11251 18569 11314
rect 17816 10801 17869 11251
rect 18491 10801 18569 11251
rect 17816 10741 18569 10801
rect 18869 11248 19620 11309
rect 18869 10845 18958 11248
rect 19533 10845 19620 11248
rect 18869 10739 19620 10845
rect 34570 10370 43150 11600
rect 34320 9992 34529 10022
rect 34320 9825 34351 9992
rect 34507 9825 34529 9992
rect 34320 9810 34529 9825
rect 33844 8358 34045 8418
rect 33844 8183 33891 8358
rect 34002 8183 34045 8358
rect 33844 8137 34045 8183
rect 36903 7505 37080 10370
rect 37400 7520 37577 10370
rect 37870 7540 38047 10370
rect 38380 7570 38557 10370
rect 38810 7580 38987 10370
rect 39230 7580 39407 10370
rect 39670 7570 39847 10370
rect 40120 7580 40297 10370
rect 34933 7155 35087 7167
rect 34933 7068 34948 7155
rect 35070 7149 35087 7155
rect 35070 7068 35528 7149
rect 34933 7058 35087 7068
rect 33840 6681 35792 6705
rect 33840 6557 35864 6681
rect 33840 6547 35792 6557
rect 43492 6498 43650 6606
rect 35202 6148 35347 6164
rect 38189 6156 38265 6164
rect 35202 6147 35524 6148
rect 35202 6036 35217 6147
rect 35329 6067 35524 6147
rect 38189 6099 38201 6156
rect 38257 6099 38265 6156
rect 38189 6087 38265 6099
rect 35329 6036 35347 6067
rect 35202 6019 35347 6036
rect 57209 5698 57574 5773
rect 41704 5484 42114 5519
rect 39707 5464 39887 5470
rect 41704 5464 41778 5484
rect 39707 5451 41778 5464
rect 39707 5348 39733 5451
rect 39863 5348 41778 5451
rect 39707 5338 41778 5348
rect 42037 5338 42114 5484
rect 39707 5316 42114 5338
rect 39707 5309 39887 5316
rect 41704 5307 42114 5316
rect 57209 5367 57270 5698
rect 57533 5367 57574 5698
rect 34940 5268 38740 5280
rect 57209 5279 57574 5367
rect 34940 5158 34958 5268
rect 35071 5260 38740 5268
rect 35071 5170 38620 5260
rect 38730 5170 38740 5260
rect 35071 5158 38740 5170
rect 34940 5150 38740 5158
rect 41708 5090 42113 5094
rect 41702 5053 42113 5090
rect 41702 5009 41757 5053
rect 33758 4795 41757 5009
rect 42024 5009 42113 5053
rect 42024 4795 45064 5009
rect 33758 4728 45064 4795
rect 41702 4717 42113 4728
rect 41708 4689 42113 4717
rect 42708 4265 43121 4516
rect 32588 3449 33088 3505
rect 37815 3449 38032 3471
rect 32588 3415 38032 3449
rect 32588 3397 37856 3415
rect 32588 3159 32655 3397
rect 32948 3247 37856 3397
rect 38001 3247 38032 3415
rect 32948 3202 38032 3247
rect 32948 3159 33088 3202
rect 37815 3171 38032 3202
rect 32588 3048 33088 3159
rect 19154 2873 19426 2933
rect 19154 2716 19196 2873
rect 19360 2716 19426 2873
rect 42201 2792 42374 2793
rect 42199 2782 42377 2792
rect 42199 2780 42213 2782
rect 19154 2679 19426 2716
rect 34551 2763 42213 2780
rect 34551 2622 34562 2763
rect 34665 2622 42213 2763
rect 34551 2603 42213 2622
rect 42369 2603 42377 2782
rect 34551 2601 42377 2603
rect 42199 2591 42377 2601
rect 34731 2456 34935 2492
rect 38108 2456 38302 2470
rect 34731 2455 38302 2456
rect 33824 2330 34082 2367
rect 30436 2124 33880 2330
rect 34068 2124 34082 2330
rect 34731 2297 34759 2455
rect 34905 2450 38302 2455
rect 34905 2299 38140 2450
rect 38281 2299 38302 2450
rect 34905 2297 38302 2299
rect 34731 2272 38302 2297
rect 34731 2262 34935 2272
rect 38108 2267 38302 2272
rect 30436 2093 34082 2124
rect 33824 2062 34082 2093
rect 43378 2178 43473 2203
rect 43378 2098 43396 2178
rect 43457 2098 43473 2178
rect 43378 2071 43473 2098
rect 35185 2027 35372 2044
rect 37477 2027 37606 2030
rect 35185 2024 37606 2027
rect 35185 1899 35214 2024
rect 35346 2008 37606 2024
rect 35346 1902 37502 2008
rect 37585 1902 37606 2008
rect 35346 1899 37606 1902
rect 35185 1895 37606 1899
rect 35185 1872 35372 1895
rect 37477 1881 37606 1895
rect 28028 1821 28258 1856
rect 28028 1665 28065 1821
rect 28228 1665 28258 1821
rect 28028 1630 28258 1665
rect 33883 1660 34022 1666
rect 30611 1647 34022 1660
rect 30611 1630 33894 1647
rect 30605 1572 33894 1630
rect 30611 1541 33894 1572
rect 34008 1541 34022 1647
rect 30611 1532 34022 1541
rect 33883 1531 34022 1532
rect 34550 1175 34672 1193
rect 34550 1088 34564 1175
rect 34662 1137 34672 1175
rect 39734 1167 39882 1185
rect 39734 1157 39754 1167
rect 34662 1090 35116 1137
rect 36204 1134 36286 1146
rect 34662 1088 34672 1090
rect 34550 1068 34672 1088
rect 36204 1075 36213 1134
rect 36273 1075 36286 1134
rect 39485 1123 39754 1157
rect 36204 1066 36286 1075
rect 39307 1068 39754 1123
rect 39485 1051 39754 1068
rect 39734 1037 39754 1051
rect 39872 1037 39882 1167
rect 39734 1018 39882 1037
rect 41742 797 42116 892
rect 41742 758 41837 797
rect 39320 675 41837 758
rect 39289 515 41837 675
rect 41742 480 41837 515
rect 42106 480 42116 797
rect 43366 544 43458 551
rect 43366 488 43380 544
rect 43440 488 43458 544
rect 43366 482 43458 488
rect 41742 417 42116 480
rect 37238 271 37329 284
rect 37238 213 37251 271
rect 37308 213 37329 271
rect 37238 197 37329 213
rect 37252 75 37309 197
rect 37113 18 37309 75
rect 34767 -1892 34909 -1880
rect 34767 -2000 34780 -1892
rect 34897 -1912 34909 -1892
rect 34897 -1996 35159 -1912
rect 36196 -1929 36287 -1916
rect 36196 -1992 36210 -1929
rect 36276 -1992 36287 -1929
rect 34897 -2000 34909 -1996
rect 34767 -2017 34909 -2000
rect 36196 -2004 36287 -1992
rect 41701 -2990 42314 -2932
rect 41701 -3053 41771 -2990
rect 30721 -3242 41771 -3053
rect 42236 -3053 42314 -2990
rect 45023 -3053 45212 -2394
rect 42236 -3242 45212 -3053
rect 41701 -3316 42314 -3242
rect 18971 -4176 19435 -3950
rect 18971 -4572 19061 -4176
rect 19310 -4572 19435 -4176
rect 57240 -4138 57627 -3991
rect 18971 -4719 19435 -4572
rect 42454 -4299 42680 -4298
rect 42454 -4352 43394 -4299
rect 42454 -4605 42485 -4352
rect 42645 -4605 43394 -4352
rect 42454 -4632 43394 -4605
rect 57240 -4593 57314 -4138
rect 57541 -4593 57627 -4138
rect 42454 -4656 42680 -4632
rect 57240 -4718 57627 -4593
rect 34226 -4954 34596 -4895
rect 34226 -5168 34281 -4954
rect 34547 -5168 34596 -4954
rect 34226 -5220 34596 -5168
rect 34768 -5556 34931 -5539
rect 42328 -5549 42544 -5529
rect 42328 -5556 42348 -5549
rect 34768 -5560 42348 -5556
rect 34768 -5708 34788 -5560
rect 34910 -5708 42348 -5560
rect 34768 -5722 42348 -5708
rect 42526 -5722 42544 -5549
rect 34768 -5732 42544 -5722
rect 42328 -5756 42544 -5732
rect 42326 -7564 42560 -7540
rect 42326 -7604 42354 -7564
rect 19088 -7739 19417 -7703
rect 41311 -7728 42354 -7604
rect 42530 -7728 42560 -7564
rect 41311 -7734 42560 -7728
rect 19088 -8019 19119 -7739
rect 19368 -8019 19417 -7739
rect 42326 -7750 42560 -7734
rect 19088 -8079 19417 -8019
rect 55478 -8641 55756 -8589
rect 55478 -8825 55513 -8641
rect 55696 -8825 55756 -8641
rect 55478 -8880 55756 -8825
rect 57244 -9679 57490 -9673
rect 57211 -9746 57563 -9679
rect 57211 -10038 57251 -9746
rect 57457 -10038 57563 -9746
rect 57211 -10104 57563 -10038
rect 41438 -10171 42929 -10127
rect 41438 -10421 41745 -10171
rect 42266 -10421 42929 -10171
rect 41438 -10472 42929 -10421
rect 19826 -12000 21571 -11979
rect 19804 -12058 21571 -12000
rect 19804 -12310 19869 -12058
rect 20071 -12310 21571 -12058
rect 19804 -12397 21571 -12310
rect 19826 -12404 21571 -12397
rect 41273 -12235 41674 -12161
rect 41273 -12413 41335 -12235
rect 41604 -12413 41674 -12235
rect 41273 -12454 41674 -12413
rect 35138 -12875 35375 -12834
rect 35138 -12881 35169 -12875
rect 34924 -13041 35169 -12881
rect 35138 -13044 35169 -13041
rect 35348 -13044 35375 -12875
rect 35138 -13077 35375 -13044
rect 37211 -14965 40395 -14903
rect 37211 -15247 38672 -14965
rect 39016 -15247 40395 -14965
rect 37211 -15309 40395 -15247
rect 57220 -16173 57646 -16072
rect 57220 -16547 57289 -16173
rect 57564 -16547 57646 -16173
rect 57220 -16623 57646 -16547
rect 19108 -17013 19454 -16917
rect 19108 -17206 19180 -17013
rect 19363 -17206 19454 -17013
rect 19108 -17290 19454 -17206
rect 36001 -18806 36246 -18777
rect 36001 -19007 36043 -18806
rect 36207 -19007 36246 -18806
rect 36001 -19062 36246 -19007
rect 56390 -19738 56703 -19713
rect 56390 -19819 56421 -19738
rect 55676 -19888 56421 -19819
rect 56390 -19908 56421 -19888
rect 56676 -19908 56703 -19738
rect 56390 -19946 56703 -19908
rect 21421 -23059 56289 -22738
rect 21421 -23526 38572 -23059
rect 39145 -23526 56289 -23059
rect 21421 -23960 56289 -23526
<< via1 >>
rect 34943 11960 35080 12114
rect 35195 11965 35347 12121
rect 35531 11961 35675 12114
rect 41698 11933 42092 12213
rect 17869 10801 18491 11251
rect 18958 10845 19533 11248
rect 34351 9825 34507 9992
rect 33891 8183 34002 8358
rect 43502 8412 43573 8494
rect 43521 7768 43575 7831
rect 33707 7359 33780 7419
rect 34948 7068 35070 7155
rect 35217 6036 35329 6147
rect 38201 6099 38257 6156
rect 38878 5565 39010 5623
rect 39259 5563 39393 5623
rect 39733 5348 39863 5451
rect 41778 5338 42037 5484
rect 57270 5367 57533 5698
rect 34958 5158 35071 5268
rect 38620 5170 38730 5260
rect 41757 4795 42024 5053
rect 32655 3159 32948 3397
rect 37856 3247 38001 3415
rect 19196 2716 19360 2873
rect 34562 2622 34665 2763
rect 42213 2603 42369 2782
rect 33880 2124 34068 2330
rect 34759 2297 34905 2455
rect 38140 2299 38281 2450
rect 43396 2098 43457 2178
rect 35214 1899 35346 2024
rect 37502 1902 37585 2008
rect 28065 1665 28228 1821
rect 33894 1541 34008 1647
rect 38890 1560 39000 1650
rect 39270 1590 39390 1660
rect 34564 1088 34662 1175
rect 36213 1075 36273 1134
rect 39754 1037 39872 1167
rect 41837 480 42106 797
rect 43380 488 43440 544
rect 37251 213 37308 271
rect 35903 19 35972 73
rect 35902 -926 35975 -873
rect 37032 -927 37108 -874
rect 34780 -2000 34897 -1892
rect 36210 -1992 36276 -1929
rect 41771 -3242 42236 -2990
rect 19061 -4572 19310 -4176
rect 42485 -4605 42645 -4352
rect 57314 -4593 57541 -4138
rect 34281 -5168 34547 -4954
rect 34788 -5708 34910 -5560
rect 42348 -5722 42526 -5549
rect 42354 -7728 42530 -7564
rect 19119 -8019 19368 -7739
rect 55513 -8825 55696 -8641
rect 57251 -10038 57457 -9746
rect 38709 -10438 38970 -10288
rect 41745 -10421 42266 -10171
rect 19869 -12310 20071 -12058
rect 41335 -12413 41604 -12235
rect 35169 -13044 35348 -12875
rect 38672 -15247 39016 -14965
rect 57289 -16547 57564 -16173
rect 19180 -17206 19363 -17013
rect 36043 -19007 36207 -18806
rect 56421 -19908 56676 -19738
rect 38572 -23526 39145 -23059
<< metal2 >>
rect 41644 12213 42163 12279
rect 34910 12114 35109 12141
rect 34910 11960 34943 12114
rect 35080 11960 35109 12114
rect 34910 11930 35109 11960
rect 35173 12121 35372 12144
rect 35173 11965 35195 12121
rect 35347 11965 35372 12121
rect 35173 11931 35372 11965
rect 35500 12114 35699 12142
rect 35500 11961 35531 12114
rect 35675 11961 35699 12114
rect 17817 11314 18567 11315
rect 17816 11251 18569 11314
rect 17816 10801 17869 11251
rect 18491 10801 18569 11251
rect 17816 10741 18569 10801
rect 18869 11273 19620 11309
rect 18869 11248 19621 11273
rect 18869 10845 18958 11248
rect 19533 10845 19621 11248
rect 17817 4646 18567 10741
rect 18869 10739 19621 10845
rect 17817 4174 18015 4646
rect 18361 4174 18567 4646
rect 17817 -5667 18567 4174
rect 17817 -6036 18068 -5667
rect 18326 -6036 18567 -5667
rect 17817 -21293 18567 -6036
rect 18871 2897 19621 10739
rect 34320 10022 34527 10023
rect 34320 9992 34529 10022
rect 34320 9825 34351 9992
rect 34507 9825 34529 9992
rect 34320 9810 34529 9825
rect 33844 8387 34045 8418
rect 33844 8160 33865 8387
rect 34022 8160 34045 8387
rect 33844 8137 34045 8160
rect 33855 8000 34077 8002
rect 33855 7980 34083 8000
rect 33855 7836 33877 7980
rect 34060 7836 34083 7980
rect 33855 7820 34083 7836
rect 33699 7436 33786 7447
rect 33699 7347 33707 7436
rect 33778 7419 33786 7436
rect 33780 7359 33786 7419
rect 33778 7347 33786 7359
rect 33699 7333 33786 7347
rect 27990 4485 28310 4525
rect 27990 4259 28023 4485
rect 28259 4259 28310 4485
rect 27990 4223 28310 4259
rect 20027 3416 20444 3462
rect 20027 3193 20069 3416
rect 20374 3193 20444 3416
rect 20027 3126 20444 3193
rect 18871 2703 19172 2897
rect 19390 2703 19621 2897
rect 18871 -4097 19621 2703
rect 18871 -4640 19016 -4097
rect 19333 -4640 19621 -4097
rect 18871 -7733 19621 -4640
rect 20070 -4934 20353 3126
rect 28027 1821 28261 4223
rect 32588 3464 33088 3505
rect 32588 3090 32613 3464
rect 33033 3090 33088 3464
rect 32588 3048 33088 3090
rect 33863 2387 34083 7820
rect 34140 7446 34252 7465
rect 34140 7338 34151 7446
rect 34237 7338 34252 7446
rect 34140 7321 34252 7338
rect 33863 2367 34082 2387
rect 33824 2330 34082 2367
rect 33824 2124 33880 2330
rect 34068 2124 34082 2330
rect 33824 2062 34082 2124
rect 28027 1665 28065 1821
rect 28228 1665 28261 1821
rect 28027 1626 28261 1665
rect 33883 1647 34022 1666
rect 33883 1541 33894 1647
rect 34008 1541 34022 1647
rect 33883 1531 34022 1541
rect 33883 -1051 34020 1531
rect 34149 -820 34229 7321
rect 34320 4580 34527 9810
rect 34703 7749 34882 7784
rect 34703 7639 34728 7749
rect 34864 7639 34882 7749
rect 34703 7594 34882 7639
rect 34289 4511 34610 4580
rect 34289 4239 34321 4511
rect 34580 4239 34610 4511
rect 34289 4173 34610 4239
rect 34704 3019 34846 7594
rect 34940 7167 35085 11930
rect 34933 7155 35087 7167
rect 34933 7068 34948 7155
rect 35070 7068 35087 7155
rect 34933 7058 35087 7068
rect 34940 5268 35085 7058
rect 34940 5158 34958 5268
rect 35071 5158 35085 5268
rect 34940 5150 35085 5158
rect 35201 6164 35346 11931
rect 35500 11929 35699 11961
rect 41644 11933 41698 12213
rect 42092 11933 42163 12213
rect 35540 8631 35681 11929
rect 41644 11850 42163 11933
rect 35519 8606 35699 8631
rect 35519 8475 35551 8606
rect 35675 8475 35699 8606
rect 35519 8454 35699 8475
rect 36673 8308 36811 8325
rect 36673 8211 36696 8308
rect 36795 8211 36811 8308
rect 36673 8187 36811 8211
rect 36723 7772 36810 8187
rect 36723 7756 36831 7772
rect 36723 7691 36743 7756
rect 36814 7691 36831 7756
rect 36723 7679 36831 7691
rect 36723 7676 36810 7679
rect 38190 6170 38259 6329
rect 35201 6147 35347 6164
rect 35201 6036 35217 6147
rect 35329 6036 35347 6147
rect 38184 6159 38271 6170
rect 38184 6091 38193 6159
rect 38261 6091 38271 6159
rect 38184 6080 38271 6091
rect 35201 6019 35347 6036
rect 34318 2877 34846 3019
rect 34108 -839 34251 -820
rect 34108 -969 34119 -839
rect 34237 -969 34251 -839
rect 34108 -982 34251 -969
rect 33879 -1061 34025 -1051
rect 33879 -1160 33893 -1061
rect 34011 -1160 34025 -1061
rect 33879 -1165 34025 -1160
rect 34318 -4895 34460 2877
rect 34551 2763 34680 2780
rect 34551 2622 34562 2763
rect 34665 2622 34680 2763
rect 34551 2601 34680 2622
rect 34558 1193 34663 2601
rect 34731 2455 34935 2492
rect 34731 2297 34759 2455
rect 34905 2297 34935 2455
rect 34731 2262 34935 2297
rect 34755 1225 34902 2262
rect 35201 2044 35346 6019
rect 38862 5623 39024 5630
rect 38862 5565 38878 5623
rect 39010 5565 39024 5623
rect 38862 5558 39024 5565
rect 39242 5623 39408 5635
rect 39242 5563 39259 5623
rect 39393 5563 39408 5623
rect 39242 5558 39408 5563
rect 37887 5487 38018 5511
rect 37887 5388 37904 5487
rect 37999 5388 38018 5487
rect 38124 5485 38290 5515
rect 38124 5463 38153 5485
rect 37887 5372 38018 5388
rect 38123 5389 38153 5463
rect 38269 5389 38290 5485
rect 37894 3471 38016 5372
rect 37815 3415 38032 3471
rect 37815 3247 37856 3415
rect 38001 3247 38032 3415
rect 37815 3171 38032 3247
rect 38123 2470 38290 5389
rect 38610 5260 38740 5280
rect 38610 5170 38620 5260
rect 38730 5170 38740 5260
rect 38610 5150 38740 5170
rect 38108 2450 38302 2470
rect 38108 2299 38140 2450
rect 38281 2299 38302 2450
rect 38108 2267 38302 2299
rect 35185 2024 35372 2044
rect 35185 1899 35214 2024
rect 35346 1899 35372 2024
rect 35185 1872 35372 1899
rect 37477 2008 37606 2030
rect 37477 1902 37502 2008
rect 37585 1902 37606 2008
rect 37477 1881 37606 1902
rect 34550 1175 34672 1193
rect 34550 1088 34564 1175
rect 34662 1088 34672 1175
rect 34755 1162 35323 1225
rect 34550 1068 34672 1088
rect 36204 1139 36286 1146
rect 36204 1075 36211 1139
rect 36279 1075 36286 1139
rect 37512 1126 37575 1881
rect 38637 1170 38700 5150
rect 38870 1650 39020 5558
rect 38870 1560 38890 1650
rect 39000 1560 39020 1650
rect 39250 1660 39400 5558
rect 41708 5519 42114 11850
rect 43491 8498 43585 8505
rect 43491 8407 43499 8498
rect 43577 8407 43585 8498
rect 43491 8394 43585 8407
rect 43136 8029 43257 8056
rect 43136 7945 43149 8029
rect 43238 7945 43257 8029
rect 43136 7932 43257 7945
rect 42436 7793 42610 7811
rect 42436 7690 42458 7793
rect 42589 7690 42610 7793
rect 42436 7676 42610 7690
rect 42204 7564 42373 7576
rect 42204 7438 42218 7564
rect 42355 7438 42373 7564
rect 42204 7419 42373 7438
rect 41704 5484 42114 5519
rect 39707 5451 39887 5470
rect 39707 5348 39733 5451
rect 39863 5348 39887 5451
rect 39707 5309 39887 5348
rect 41140 5395 41368 5415
rect 39250 1590 39270 1660
rect 39390 1590 39400 1660
rect 39250 1580 39400 1590
rect 38870 1550 39020 1560
rect 39736 1185 39881 5309
rect 41140 5288 41168 5395
rect 41335 5288 41368 5395
rect 41704 5338 41778 5484
rect 42037 5338 42114 5484
rect 41704 5307 42114 5338
rect 41140 5244 41368 5288
rect 40772 3478 40932 3492
rect 40772 3333 40784 3478
rect 40913 3333 40932 3478
rect 40772 3318 40932 3333
rect 40783 1850 40929 3318
rect 40758 1825 40961 1850
rect 40758 1710 40793 1825
rect 40930 1710 40961 1825
rect 40758 1684 40961 1710
rect 39734 1167 39882 1185
rect 36204 1066 36286 1075
rect 39734 1037 39754 1167
rect 39872 1037 39882 1167
rect 39734 1018 39882 1037
rect 39736 1016 39881 1018
rect 37238 272 37329 284
rect 40844 283 40979 302
rect 40844 277 40858 283
rect 37238 204 37249 272
rect 37317 204 37329 272
rect 37238 197 37329 204
rect 40843 200 40858 277
rect 40964 200 40979 283
rect 40843 182 40979 200
rect 35883 84 35985 94
rect 35883 7 35893 84
rect 35976 7 35985 84
rect 35883 -5 35985 7
rect 35889 -859 35982 -848
rect 35889 -938 35895 -859
rect 35978 -938 35982 -859
rect 35889 -949 35982 -938
rect 37013 -855 37113 -846
rect 37013 -933 37022 -855
rect 37101 -874 37113 -855
rect 37108 -927 37113 -874
rect 37101 -933 37113 -927
rect 37013 -940 37113 -933
rect 34767 -1892 34909 -1880
rect 34767 -2000 34780 -1892
rect 34897 -2000 34909 -1892
rect 34767 -2017 34909 -2000
rect 36196 -1924 36287 -1916
rect 36196 -1996 36205 -1924
rect 36279 -1996 36287 -1924
rect 36196 -2004 36287 -1996
rect 18871 -8031 19101 -7733
rect 19398 -8031 19621 -7733
rect 18871 -16979 19621 -8031
rect 19806 -5217 20353 -4934
rect 34226 -4954 34596 -4895
rect 34226 -5168 34281 -4954
rect 34547 -5168 34596 -4954
rect 19806 -10256 20089 -5217
rect 34226 -5220 34596 -5168
rect 34790 -5539 34904 -2017
rect 35155 -2569 35392 -2546
rect 40843 -2569 40971 182
rect 35155 -2707 35175 -2569
rect 35355 -2707 35392 -2569
rect 35155 -2732 35392 -2707
rect 40834 -2590 41014 -2569
rect 34768 -5560 34931 -5539
rect 34768 -5708 34788 -5560
rect 34910 -5708 34931 -5560
rect 34768 -5732 34931 -5708
rect 35189 -8000 35353 -2732
rect 40834 -2791 40849 -2590
rect 40987 -2791 41014 -2590
rect 40834 -2804 41014 -2791
rect 41169 -5943 41328 5244
rect 41708 5090 42114 5094
rect 41702 5053 42114 5090
rect 41702 4795 41757 5053
rect 42024 4795 42114 5053
rect 41702 4717 42114 4795
rect 41708 915 42114 4717
rect 42208 2793 42365 7419
rect 42201 2792 42374 2793
rect 42199 2782 42377 2792
rect 42199 2603 42213 2782
rect 42369 2603 42377 2782
rect 42199 2591 42377 2603
rect 41708 797 42116 915
rect 41708 480 41837 797
rect 42106 480 42116 797
rect 41708 317 42116 480
rect 41708 81 42118 317
rect 41708 -2854 42116 81
rect 41708 -2932 42316 -2854
rect 41701 -2990 42316 -2932
rect 41701 -3242 41771 -2990
rect 42236 -3242 42316 -2990
rect 41701 -3316 42316 -3242
rect 41708 -4991 42316 -3316
rect 42455 -4298 42603 7676
rect 42819 6613 42993 6614
rect 42818 6600 42993 6613
rect 42818 6474 42834 6600
rect 42970 6474 42993 6600
rect 42818 4516 42993 6474
rect 43151 6161 43255 7932
rect 43500 7836 43586 7846
rect 43500 7759 43510 7836
rect 43575 7759 43586 7836
rect 43500 7749 43586 7759
rect 43489 6590 43651 6606
rect 43489 6512 43530 6590
rect 43610 6512 43651 6590
rect 43489 6494 43651 6512
rect 43151 6057 43329 6161
rect 42708 4471 43121 4516
rect 42708 4310 42782 4471
rect 43061 4310 43121 4471
rect 42708 4265 43121 4310
rect 42890 -734 42947 4265
rect 43225 3483 43329 6057
rect 57001 5739 57751 8305
rect 57001 5320 57242 5739
rect 57547 5320 57751 5739
rect 43060 3379 43329 3483
rect 56354 3492 56692 3519
rect 43060 2187 43164 3379
rect 56354 3260 56384 3492
rect 56662 3260 56692 3492
rect 56354 3217 56692 3260
rect 43378 2187 43473 2203
rect 43060 2178 43473 2187
rect 43060 2098 43396 2178
rect 43457 2098 43473 2178
rect 43060 2083 43473 2098
rect 43378 2071 43473 2083
rect 43034 549 43146 560
rect 43034 473 43051 549
rect 43135 473 43146 549
rect 43366 547 43458 551
rect 43366 485 43376 547
rect 43448 485 43458 547
rect 43366 482 43458 485
rect 43034 458 43146 473
rect 43046 103 43140 458
rect 43040 87 43152 103
rect 43040 11 43056 87
rect 43140 11 43152 87
rect 43040 -1 43152 11
rect 42890 -791 43679 -734
rect 55980 -2585 56278 -2546
rect 55980 -2807 56003 -2585
rect 56241 -2807 56278 -2585
rect 55980 -2852 56278 -2807
rect 42454 -4352 42680 -4298
rect 42454 -4605 42485 -4352
rect 42645 -4605 42680 -4352
rect 42454 -4656 42680 -4605
rect 41169 -6102 41567 -5943
rect 35189 -8971 35271 -8000
rect 35189 -8972 35336 -8971
rect 19807 -12000 20087 -10256
rect 19804 -12058 20143 -12000
rect 19804 -12310 19869 -12058
rect 20071 -12310 20143 -12058
rect 19804 -12397 20143 -12310
rect 35186 -12834 35336 -8972
rect 38608 -10288 39073 -10254
rect 38608 -10438 38709 -10288
rect 38970 -10438 39073 -10288
rect 35138 -12875 35375 -12834
rect 35138 -13044 35169 -12875
rect 35348 -13044 35375 -12875
rect 35138 -13077 35375 -13044
rect 18871 -17246 19155 -16979
rect 19388 -17246 19621 -16979
rect 18871 -21147 19621 -17246
rect 38608 -14965 39073 -10438
rect 41408 -12161 41567 -6102
rect 41708 -9877 42116 -4991
rect 42328 -5549 42544 -5529
rect 56008 -5530 56265 -2852
rect 42328 -5722 42348 -5549
rect 42526 -5722 42544 -5549
rect 55770 -5666 56265 -5530
rect 42328 -5756 42544 -5722
rect 42350 -7540 42529 -5756
rect 42326 -7564 42560 -7540
rect 42326 -7728 42354 -7564
rect 42530 -7728 42560 -7564
rect 42326 -7750 42560 -7728
rect 55478 -8618 55756 -8589
rect 55478 -8866 55495 -8618
rect 55721 -8866 55756 -8618
rect 55478 -8880 55756 -8866
rect 41708 -10171 42316 -9877
rect 41708 -10421 41745 -10171
rect 42266 -10421 42316 -10171
rect 41708 -10469 42316 -10421
rect 41273 -12235 41674 -12161
rect 41273 -12413 41335 -12235
rect 41604 -12413 41674 -12235
rect 41273 -12454 41674 -12413
rect 38608 -15247 38672 -14965
rect 39016 -15247 39073 -14965
rect 35977 -18806 36310 -18773
rect 35977 -19007 36043 -18806
rect 36207 -19007 36310 -18806
rect 17794 -21374 18567 -21293
rect 17794 -21836 17929 -21374
rect 18465 -21836 18567 -21374
rect 35977 -21412 36310 -19007
rect 17794 -21924 18567 -21836
rect 35823 -21527 36450 -21412
rect 35823 -21809 35912 -21527
rect 36348 -21809 36450 -21527
rect 35823 -21873 36450 -21809
rect 17794 -21951 18560 -21924
rect 38608 -22941 39073 -15247
rect 41992 -16829 42276 -16807
rect 41992 -17003 42022 -16829
rect 42239 -17003 42276 -16829
rect 41992 -17041 42276 -17003
rect 42891 -16856 43179 -16830
rect 42891 -16990 42947 -16856
rect 43146 -16990 43179 -16856
rect 42891 -17026 43179 -16990
rect 42019 -21404 42241 -17041
rect 56404 -19713 56685 3217
rect 57001 -1680 57751 5320
rect 57001 -2071 57206 -1680
rect 57480 -2071 57751 -1680
rect 57001 -4082 57751 -2071
rect 57001 -4667 57286 -4082
rect 57576 -4667 57751 -4082
rect 57001 -9726 57751 -4667
rect 57001 -10051 57237 -9726
rect 57490 -10051 57751 -9726
rect 57001 -16141 57751 -10051
rect 57001 -16560 57269 -16141
rect 57584 -16560 57751 -16141
rect 56390 -19738 56703 -19713
rect 56390 -19908 56421 -19738
rect 56676 -19908 56703 -19738
rect 56390 -19946 56703 -19908
rect 57001 -21282 57751 -16560
rect 58223 4673 58973 8277
rect 58223 4114 58446 4673
rect 58860 4114 58973 4673
rect 58223 -8539 58973 4114
rect 58223 -8967 58398 -8539
rect 58813 -8967 58973 -8539
rect 58223 -21286 58973 -8967
rect 58202 -21340 58979 -21286
rect 41930 -21483 42382 -21404
rect 41930 -21764 41995 -21483
rect 42303 -21764 42382 -21483
rect 41930 -21823 42382 -21764
rect 58202 -21871 58283 -21340
rect 58922 -21871 58979 -21340
rect 58202 -21942 58979 -21871
rect 38465 -23059 39241 -22941
rect 38465 -23526 38572 -23059
rect 39145 -23526 39241 -23059
rect 38465 -23610 39241 -23526
<< via2 >>
rect 19179 10964 19388 11180
rect 18015 4174 18361 4646
rect 18068 -6036 18326 -5667
rect 33865 8358 34022 8387
rect 33865 8183 33891 8358
rect 33891 8183 34002 8358
rect 34002 8183 34022 8358
rect 33865 8160 34022 8183
rect 33877 7836 34060 7980
rect 33707 7419 33778 7436
rect 33707 7359 33778 7419
rect 33707 7347 33778 7359
rect 28023 4259 28259 4485
rect 20069 3193 20374 3416
rect 19172 2873 19390 2897
rect 19172 2716 19196 2873
rect 19196 2716 19360 2873
rect 19360 2716 19390 2873
rect 19172 2703 19390 2716
rect 19016 -4176 19333 -4097
rect 19016 -4572 19061 -4176
rect 19061 -4572 19310 -4176
rect 19310 -4572 19333 -4176
rect 19016 -4640 19333 -4572
rect 32613 3397 33033 3464
rect 32613 3159 32655 3397
rect 32655 3159 32948 3397
rect 32948 3159 33033 3397
rect 32613 3090 33033 3159
rect 34151 7338 34237 7446
rect 34728 7639 34864 7749
rect 34321 4239 34580 4511
rect 35551 8475 35675 8606
rect 36696 8211 36795 8308
rect 36743 7691 36814 7756
rect 38193 6156 38261 6159
rect 38193 6099 38201 6156
rect 38201 6099 38257 6156
rect 38257 6099 38261 6156
rect 38193 6091 38261 6099
rect 34119 -969 34237 -839
rect 33893 -1160 34011 -1061
rect 37904 5388 37999 5487
rect 38153 5389 38269 5485
rect 36211 1134 36279 1139
rect 36211 1075 36213 1134
rect 36213 1075 36273 1134
rect 36273 1075 36279 1134
rect 43499 8494 43577 8498
rect 43499 8412 43502 8494
rect 43502 8412 43573 8494
rect 43573 8412 43577 8494
rect 43499 8407 43577 8412
rect 43149 7945 43238 8029
rect 42458 7690 42589 7793
rect 42218 7438 42355 7564
rect 41168 5288 41335 5395
rect 40784 3333 40913 3478
rect 40793 1710 40930 1825
rect 37249 271 37317 272
rect 37249 213 37251 271
rect 37251 213 37308 271
rect 37308 213 37317 271
rect 37249 204 37317 213
rect 40858 200 40964 283
rect 35893 73 35976 84
rect 35893 19 35903 73
rect 35903 19 35972 73
rect 35972 19 35976 73
rect 35893 7 35976 19
rect 35895 -873 35978 -859
rect 35895 -926 35902 -873
rect 35902 -926 35975 -873
rect 35975 -926 35978 -873
rect 35895 -938 35978 -926
rect 37022 -874 37101 -855
rect 37022 -927 37032 -874
rect 37032 -927 37101 -874
rect 37022 -933 37101 -927
rect 36205 -1929 36279 -1924
rect 36205 -1992 36210 -1929
rect 36210 -1992 36276 -1929
rect 36276 -1992 36279 -1929
rect 36205 -1996 36279 -1992
rect 19101 -7739 19398 -7733
rect 19101 -8019 19119 -7739
rect 19119 -8019 19368 -7739
rect 19368 -8019 19398 -7739
rect 19101 -8031 19398 -8019
rect 35175 -2707 35355 -2569
rect 40849 -2791 40987 -2590
rect 42834 6474 42970 6600
rect 43510 7831 43575 7836
rect 43510 7768 43521 7831
rect 43521 7768 43575 7831
rect 43510 7759 43575 7768
rect 43530 6512 43610 6590
rect 42782 4310 43061 4471
rect 57242 5698 57547 5739
rect 57242 5367 57270 5698
rect 57270 5367 57533 5698
rect 57533 5367 57547 5698
rect 57242 5320 57547 5367
rect 56384 3260 56662 3492
rect 43051 473 43135 549
rect 43376 544 43448 547
rect 43376 488 43380 544
rect 43380 488 43440 544
rect 43440 488 43448 544
rect 43376 485 43448 488
rect 43056 11 43140 87
rect 56003 -2807 56241 -2585
rect 19155 -17013 19388 -16979
rect 19155 -17206 19180 -17013
rect 19180 -17206 19363 -17013
rect 19363 -17206 19388 -17013
rect 19155 -17246 19388 -17206
rect 55495 -8641 55721 -8618
rect 55495 -8825 55513 -8641
rect 55513 -8825 55696 -8641
rect 55696 -8825 55721 -8641
rect 55495 -8866 55721 -8825
rect 17929 -21836 18465 -21374
rect 35912 -21809 36348 -21527
rect 42022 -17003 42239 -16829
rect 42947 -16990 43146 -16856
rect 57206 -2071 57480 -1680
rect 57286 -4138 57576 -4082
rect 57286 -4593 57314 -4138
rect 57314 -4593 57541 -4138
rect 57541 -4593 57576 -4138
rect 57286 -4667 57576 -4593
rect 57237 -9746 57490 -9726
rect 57237 -10038 57251 -9746
rect 57251 -10038 57457 -9746
rect 57457 -10038 57490 -9746
rect 57237 -10051 57490 -10038
rect 57269 -16173 57584 -16141
rect 57269 -16547 57289 -16173
rect 57289 -16547 57564 -16173
rect 57564 -16547 57584 -16173
rect 57269 -16560 57584 -16547
rect 58446 4114 58860 4673
rect 58398 -8967 58813 -8539
rect 41995 -21764 42303 -21483
rect 58283 -21871 58922 -21340
<< metal3 >>
rect 19158 11180 19415 11195
rect 19158 10964 19179 11180
rect 19388 11103 19415 11180
rect 19388 11026 21798 11103
rect 19388 10964 19415 11026
rect 19158 10929 19415 10964
rect 35519 8606 35699 8631
rect 35519 8475 35551 8606
rect 35675 8574 35699 8606
rect 35675 8475 38320 8574
rect 43491 8498 43585 8505
rect 43491 8493 43499 8498
rect 35519 8470 38320 8475
rect 35519 8454 35699 8470
rect 33844 8387 34045 8418
rect 33844 8160 33865 8387
rect 34022 8322 34045 8387
rect 36673 8322 36811 8325
rect 34022 8308 36811 8322
rect 34022 8211 36696 8308
rect 36795 8211 36811 8308
rect 34022 8187 36811 8211
rect 34022 8184 36808 8187
rect 34022 8160 34045 8184
rect 33844 8137 34045 8160
rect 33855 7998 34077 8002
rect 33855 7980 38123 7998
rect 33855 7836 33877 7980
rect 34060 7911 38123 7980
rect 34060 7910 37811 7911
rect 34060 7836 34077 7910
rect 33855 7820 34077 7836
rect 34703 7766 34882 7784
rect 34703 7749 36674 7766
rect 34703 7639 34728 7749
rect 34864 7700 36674 7749
rect 34864 7639 34882 7700
rect 34703 7594 34882 7639
rect 33699 7446 33786 7447
rect 34140 7446 34252 7465
rect 33699 7436 34151 7446
rect 33699 7347 33707 7436
rect 33778 7347 34151 7436
rect 33699 7338 34151 7347
rect 34237 7338 34253 7446
rect 36608 7427 36674 7700
rect 36731 7756 36831 7772
rect 36731 7691 36743 7756
rect 36814 7691 36831 7756
rect 36731 7679 36831 7691
rect 36731 7460 36802 7679
rect 38036 7440 38123 7911
rect 33699 7333 34253 7338
rect 34140 7321 34252 7333
rect 37916 5511 38002 6591
rect 38216 6378 38320 8470
rect 38828 8407 43499 8493
rect 43577 8407 43585 8498
rect 38828 7424 38914 8407
rect 43491 8394 43585 8407
rect 43136 8029 43257 8056
rect 43136 8016 43149 8029
rect 39048 7958 43149 8016
rect 39048 7441 39106 7958
rect 43136 7945 43149 7958
rect 43238 7945 43257 8029
rect 43136 7932 43257 7945
rect 43500 7839 43586 7846
rect 42859 7836 43586 7839
rect 42436 7793 42610 7811
rect 42436 7761 42458 7793
rect 39886 7409 39972 7759
rect 40148 7701 42458 7761
rect 40148 7444 40208 7701
rect 42436 7690 42458 7701
rect 42589 7690 42610 7793
rect 42436 7676 42610 7690
rect 42859 7759 43510 7836
rect 43575 7759 43586 7836
rect 42859 7758 43586 7759
rect 42204 7564 42373 7576
rect 42859 7564 42957 7758
rect 43500 7749 43586 7758
rect 42204 7438 42218 7564
rect 42355 7438 42957 7564
rect 42204 7423 42957 7438
rect 42204 7419 42373 7423
rect 42819 6607 42993 6614
rect 42819 6606 43602 6607
rect 42819 6600 43651 6606
rect 42819 6474 42834 6600
rect 42970 6590 43651 6600
rect 42970 6512 43530 6590
rect 43610 6512 43651 6590
rect 42970 6494 43651 6512
rect 42970 6474 42993 6494
rect 42819 6454 42993 6474
rect 38161 6274 38320 6378
rect 38161 6170 38265 6274
rect 38161 6159 38271 6170
rect 38161 6091 38193 6159
rect 38261 6091 38271 6159
rect 38161 6080 38271 6091
rect 38161 5515 38265 6080
rect 37887 5487 38018 5511
rect 37887 5388 37904 5487
rect 37999 5388 38018 5487
rect 37887 5372 38018 5388
rect 38124 5485 38290 5515
rect 38124 5389 38153 5485
rect 38269 5389 38290 5485
rect 38124 5368 38290 5389
rect 39886 5359 39972 6312
rect 57209 5739 57574 5773
rect 57209 5557 57242 5739
rect 53733 5480 57242 5557
rect 41140 5395 41368 5415
rect 41140 5359 41168 5395
rect 39886 5288 41168 5359
rect 41335 5288 41368 5395
rect 39886 5273 41368 5288
rect 57209 5320 57242 5480
rect 57547 5320 57574 5739
rect 57209 5279 57574 5320
rect 41140 5244 41368 5273
rect 17918 4646 18476 4749
rect 17918 4174 18015 4646
rect 18361 4578 18476 4646
rect 58325 4673 58921 4807
rect 34257 4578 34638 4580
rect 58325 4578 58446 4673
rect 18361 4511 58446 4578
rect 18361 4485 34321 4511
rect 18361 4259 28023 4485
rect 28259 4259 34321 4485
rect 18361 4239 34321 4259
rect 34580 4471 58446 4511
rect 34580 4310 42782 4471
rect 43061 4310 58446 4471
rect 34580 4239 58446 4310
rect 18361 4174 58446 4239
rect 17918 4083 18476 4174
rect 34257 4173 34638 4174
rect 58325 4114 58446 4174
rect 58860 4114 58921 4673
rect 58325 4004 58921 4114
rect 32588 3464 33088 3505
rect 56354 3492 56692 3519
rect 20027 3416 20444 3462
rect 20027 3193 20069 3416
rect 20374 3413 20444 3416
rect 32588 3413 32613 3464
rect 20374 3193 32613 3413
rect 20027 3176 32613 3193
rect 20027 3126 20444 3176
rect 32588 3090 32613 3176
rect 33033 3090 33088 3464
rect 40772 3478 56384 3492
rect 40772 3333 40784 3478
rect 40913 3333 56384 3478
rect 40772 3318 56384 3333
rect 56354 3260 56384 3318
rect 56662 3260 56692 3492
rect 56354 3217 56692 3260
rect 32588 3048 33088 3090
rect 19154 2897 19426 2933
rect 19154 2703 19172 2897
rect 19390 2848 19426 2897
rect 19390 2752 24487 2848
rect 19390 2703 19426 2752
rect 19154 2679 19426 2703
rect 40758 1825 40961 1850
rect 40758 1786 40793 1825
rect 36204 1710 40793 1786
rect 40930 1710 40961 1825
rect 36204 1704 40961 1710
rect 36204 1139 36286 1704
rect 40758 1684 40961 1704
rect 36204 1075 36211 1139
rect 36279 1075 36286 1139
rect 36204 1066 36286 1075
rect 43034 551 43146 560
rect 43034 549 43458 551
rect 43034 473 43051 549
rect 43135 547 43458 549
rect 43135 485 43376 547
rect 43448 485 43458 547
rect 43135 481 43458 485
rect 43135 473 43146 481
rect 43034 458 43146 473
rect 37238 278 37329 284
rect 40844 283 40979 302
rect 40844 278 40858 283
rect 37238 272 40858 278
rect 37238 204 37249 272
rect 37317 204 40858 272
rect 37238 200 40858 204
rect 40964 200 40979 283
rect 37238 199 40979 200
rect 37238 197 37329 199
rect 40844 182 40979 199
rect 35883 89 35985 94
rect 43040 89 43152 103
rect 35883 87 43152 89
rect 35883 84 43056 87
rect 35883 7 35893 84
rect 35976 11 43056 84
rect 43140 11 43152 87
rect 35976 7 43152 11
rect 35883 2 43152 7
rect 35883 -5 35985 2
rect 43040 -1 43152 2
rect 34108 -839 34251 -820
rect 34108 -969 34119 -839
rect 34237 -850 34251 -839
rect 35889 -850 35982 -848
rect 34237 -859 35982 -850
rect 34237 -938 35895 -859
rect 35978 -938 35982 -859
rect 34237 -946 35982 -938
rect 34237 -969 34251 -946
rect 35889 -949 35982 -946
rect 37013 -855 37113 -846
rect 37013 -933 37022 -855
rect 37101 -933 37113 -855
rect 34108 -982 34251 -969
rect 33879 -1059 34025 -1051
rect 37013 -1059 37113 -933
rect 33879 -1061 37113 -1059
rect 33879 -1160 33893 -1061
rect 34011 -1159 37113 -1061
rect 34011 -1160 34025 -1159
rect 33879 -1165 34025 -1160
rect 57144 -1680 57542 -1584
rect 57144 -1829 57206 -1680
rect 52444 -1906 57206 -1829
rect 36196 -1924 36287 -1916
rect 36196 -1996 36205 -1924
rect 36279 -1996 36287 -1924
rect 36196 -2004 36287 -1996
rect 35155 -2569 35392 -2546
rect 35155 -2707 35175 -2569
rect 35355 -2586 35392 -2569
rect 36196 -2586 36284 -2004
rect 57144 -2071 57206 -1906
rect 57480 -2071 57542 -1680
rect 57144 -2201 57542 -2071
rect 35355 -2674 36284 -2586
rect 40834 -2571 41014 -2569
rect 55980 -2571 56278 -2546
rect 40834 -2585 56278 -2571
rect 40834 -2590 56003 -2585
rect 35355 -2707 35392 -2674
rect 35155 -2732 35392 -2707
rect 40834 -2791 40849 -2590
rect 40987 -2791 56003 -2590
rect 40834 -2804 56003 -2791
rect 55980 -2807 56003 -2804
rect 56241 -2807 56278 -2585
rect 55980 -2852 56278 -2807
rect 18971 -4097 19435 -3950
rect 18971 -4640 19016 -4097
rect 19333 -4165 19435 -4097
rect 57240 -4082 57627 -3991
rect 57240 -4165 57286 -4082
rect 19333 -4569 57286 -4165
rect 19333 -4640 19435 -4569
rect 18971 -4719 19435 -4640
rect 57240 -4667 57286 -4569
rect 57576 -4667 57627 -4082
rect 57240 -4718 57627 -4667
rect 18018 -5667 18388 -5581
rect 18018 -6036 18068 -5667
rect 18326 -5855 18388 -5667
rect 18326 -5944 20728 -5855
rect 18326 -6036 18388 -5944
rect 18018 -6110 18388 -6036
rect 19088 -7733 19417 -7703
rect 19088 -8031 19101 -7733
rect 19398 -7844 19417 -7733
rect 19398 -7961 21052 -7844
rect 19398 -8031 19417 -7961
rect 19088 -8079 19417 -8031
rect 58352 -8539 58873 -8459
rect 58352 -8586 58398 -8539
rect 55478 -8618 58398 -8586
rect 55478 -8866 55495 -8618
rect 55721 -8866 58398 -8618
rect 55478 -8880 58398 -8866
rect 58352 -8967 58398 -8880
rect 58813 -8967 58873 -8539
rect 58352 -9020 58873 -8967
rect 57244 -9679 57490 -9673
rect 57211 -9726 57563 -9679
rect 57211 -9879 57237 -9726
rect 52242 -9936 57237 -9879
rect 57211 -10051 57237 -9936
rect 57490 -10051 57563 -9726
rect 57211 -10104 57563 -10051
rect 20882 -11188 55877 -10784
rect 57220 -16141 57646 -16072
rect 57220 -16311 57269 -16141
rect 53784 -16459 57269 -16311
rect 57220 -16560 57269 -16459
rect 57584 -16560 57646 -16141
rect 57220 -16623 57646 -16560
rect 41992 -16829 42276 -16807
rect 19108 -16979 19454 -16917
rect 19108 -17246 19155 -16979
rect 19388 -17066 19454 -16979
rect 41992 -17003 42022 -16829
rect 42239 -16856 43193 -16829
rect 42239 -16990 42947 -16856
rect 43146 -16990 43193 -16856
rect 42239 -17003 43193 -16990
rect 41992 -17032 43193 -17003
rect 41992 -17041 42276 -17032
rect 19388 -17147 23318 -17066
rect 19388 -17246 19454 -17147
rect 19108 -17290 19454 -17246
rect 58202 -21289 58979 -21286
rect 17773 -21340 58979 -21289
rect 17773 -21374 58283 -21340
rect 17773 -21836 17929 -21374
rect 18465 -21483 58283 -21374
rect 18465 -21527 41995 -21483
rect 18465 -21809 35912 -21527
rect 36348 -21764 41995 -21527
rect 42303 -21764 58283 -21483
rect 36348 -21809 58283 -21764
rect 18465 -21836 58283 -21809
rect 17773 -21871 58283 -21836
rect 58922 -21871 58979 -21340
rect 17773 -21942 58979 -21871
rect 17773 -21947 58961 -21942
rect 17794 -21951 18560 -21947
use CLK_div_90_mag  CLK_div_90_mag_0
timestamp 1694669839
transform 1 0 18281 0 1 301
box 3140 4330 16201 11389
use CLK_div_93_mag  CLK_div_93_mag_0
timestamp 1694669839
transform 1 0 20761 0 1 -10236
box -502 -242 21015 5340
use CLK_div_96_mag  CLK_div_96_mag_0
timestamp 1694669839
transform 1 0 21556 0 1 -3347
box 52 105 9646 6783
use CLK_div_99_mag  CLK_div_99_mag_0
timestamp 1694669839
transform 1 0 19954 0 1 -28521
box 1317 7658 17710 16746
use CLK_div_100_mag  CLK_div_100_mag_0
timestamp 1694669839
transform 1 0 43329 0 1 -2455
box -125 0 12197 5567
use CLK_div_100_mag  CLK_div_100_mag_1
timestamp 1694669839
transform 1 0 43441 0 1 4931
box -125 0 12197 5567
use CLK_div_108_new_mag  CLK_div_108_new_mag_0
timestamp 1694669839
transform 1 0 36094 0 1 -10375
box 6435 -290 19896 6076
use CLK_div_110_mag  CLK_div_110_mag_0
timestamp 1694669839
transform 1 0 42879 0 1 -18358
box -2562 -2430 13288 6270
use mux_8x1_ibr  mux_8x1_ibr_0
timestamp 1694669839
transform 1 0 34946 0 1 -427
box 0 -2102 4512 2102
<< labels >>
flabel metal1 30140 -23490 30140 -23490 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal1 37488 10946 37488 10946 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel via1 35001 12031 35001 12031 0 FreeSans 1600 0 0 0 F2
port 2 nsew
flabel via1 35267 12049 35267 12049 0 FreeSans 1440 0 0 0 F1
port 3 nsew
flabel via1 35596 12043 35596 12043 0 FreeSans 1440 0 0 0 F0
port 4 nsew
flabel via1 18121 11047 18121 11047 0 FreeSans 1440 0 0 0 CLK
port 5 nsew
flabel via1 19095 11035 19095 11035 0 FreeSans 1440 0 0 0 RST
port 6 nsew
flabel via1 41870 12076 41870 12076 0 FreeSans 1440 0 0 0 Vdiv
port 7 nsew
<< end >>
