magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1539 1045 1539
<< metal2 >>
rect -45 534 45 539
rect -45 -534 -40 534
rect 40 -534 45 534
rect -45 -539 45 -534
<< via2 >>
rect -40 -534 40 534
<< metal3 >>
rect -45 534 45 539
rect -45 -534 -40 534
rect 40 -534 45 534
rect -45 -539 45 -534
<< end >>
