* NGSPICE file created from INV_2_flat.ext - technology: gf180mcuC

.subckt INV_2_flat VDD VSS IN OUT
X0 OUT IN.t0 VSS.t9 VSS.t8 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X1 OUT IN.t1 VSS.t7 VSS.t6 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X2 OUT IN.t2 VDD.t15 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
X3 OUT IN.t3 VDD.t14 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X4 VDD IN.t4 OUT.t4 VDD.t9 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X5 VDD IN.t5 OUT.t3 VDD.t9 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X6 VDD IN.t6 OUT.t2 VDD.t2 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X7 OUT IN.t7 VDD.t6 VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X8 VSS IN.t8 OUT.t8 VSS.t3 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.5u
X9 VSS IN.t9 OUT.t7 VSS.t0 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X10 VDD IN.t10 OUT.t1 VDD.t2 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.5u
X11 OUT IN.t11 VDD.t1 VDD.t0 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.5u
R0 IN.n4 IN.t9 28.3986
R1 IN.n5 IN.n4 23.7519
R2 IN.n6 IN.n5 19.7846
R3 IN.n1 IN.n0 12.2457
R4 IN.n2 IN.n1 12.2457
R5 IN.n3 IN.n2 12.2457
R6 IN.n7 IN.t11 11.6285
R7 IN.n0 IN.t10 8.9065
R8 IN.n1 IN.t7 8.9065
R9 IN.n2 IN.t4 8.9065
R10 IN.n3 IN.t2 8.9065
R11 IN.n6 IN.t0 8.59715
R12 IN.n0 IN.t6 8.3225
R13 IN.n1 IN.t3 8.3225
R14 IN.n2 IN.t5 8.3225
R15 IN.t11 IN.n3 8.3225
R16 IN IN.n7 4.223
R17 IN.n4 IN.t1 3.6505
R18 IN.n5 IN.t8 3.6505
R19 IN.n7 IN.n6 3.1807
R20 VSS.n17 VSS.n16 759.951
R21 VSS.n8 VSS.t0 250.623
R22 VSS.n23 VSS.t8 137.439
R23 VSS.n16 VSS.t6 121.269
R24 VSS.n18 VSS.n15 9.13939
R25 VSS.n30 VSS.n18 9.13939
R26 VSS.n29 VSS.t3 8.08508
R27 VSS.n4 VSS.n3 6.65541
R28 VSS.n19 VSS.t9 6.65541
R29 VSS VSS.n18 5.2005
R30 VSS VSS.n18 5.2005
R31 VSS.n2 VSS.n1 3.37941
R32 VSS.n1 VSS.t7 3.2765
R33 VSS.n1 VSS.n0 3.2765
R34 VSS.n7 VSS.n6 2.6005
R35 VSS.n10 VSS.n9 2.6005
R36 VSS.n9 VSS.n8 2.6005
R37 VSS.n13 VSS.n12 2.6005
R38 VSS.n12 VSS.n11 2.6005
R39 VSS.n15 VSS.n14 2.6005
R40 VSS.n16 VSS.n15 2.6005
R41 VSS.n18 VSS.n17 2.6005
R42 VSS.n31 VSS.n30 2.6005
R43 VSS.n30 VSS.n29 2.6005
R44 VSS.n28 VSS.n27 2.6005
R45 VSS.n27 VSS.n26 2.6005
R46 VSS.n25 VSS.n24 2.6005
R47 VSS.n24 VSS.n23 2.6005
R48 VSS.n22 VSS.n21 2.6005
R49 VSS.n10 VSS.n7 0.0596608
R50 VSS.n13 VSS.n10 0.0596608
R51 VSS.n14 VSS.n13 0.0596608
R52 VSS VSS.n31 0.0596608
R53 VSS.n31 VSS.n28 0.0596608
R54 VSS.n28 VSS.n25 0.0596608
R55 VSS.n25 VSS.n22 0.0596608
R56 VSS.n14 VSS.n2 0.0552552
R57 VSS.n21 VSS.n20 0.0316876
R58 VSS.n6 VSS.n5 0.0316876
R59 VSS.n7 VSS.n4 0.0250455
R60 VSS.n22 VSS.n19 0.0162343
R61 VSS VSS.n2 0.00490559
R62 OUT.n3 OUT.t2 3.6405
R63 OUT.n3 OUT.n2 3.6405
R64 OUT.n1 OUT.t1 3.6405
R65 OUT.n1 OUT.n0 3.6405
R66 OUT.n10 OUT.t3 3.6405
R67 OUT.n10 OUT.n9 3.6405
R68 OUT.n8 OUT.t4 3.6405
R69 OUT.n8 OUT.n7 3.6405
R70 OUT.n15 OUT.n6 3.50463
R71 OUT.n14 OUT.n13 3.50463
R72 OUT.n6 OUT.t7 3.2765
R73 OUT.n6 OUT.n5 3.2765
R74 OUT.n13 OUT.t8 3.2765
R75 OUT.n13 OUT.n12 3.2765
R76 OUT.n4 OUT.n1 3.06224
R77 OUT.n11 OUT.n8 3.05425
R78 OUT.n4 OUT.n3 2.6005
R79 OUT.n11 OUT.n10 2.6005
R80 OUT.n15 OUT.n14 0.798761
R81 OUT OUT.n15 0.562022
R82 OUT.n15 OUT.n4 0.18637
R83 OUT.n14 OUT.n11 0.18637
R84 VDD.n32 VDD.n31 128.591
R85 VDD.n25 VDD.t0 39.6722
R86 VDD.n32 VDD.t9 21.8883
R87 VDD.n5 VDD.t2 13.6804
R88 VDD.n14 VDD.n13 8.488
R89 VDD.n33 VDD.n14 8.2255
R90 VDD.n20 VDD.t1 6.70224
R91 VDD.n2 VDD.n1 6.70224
R92 VDD VDD.n14 6.3005
R93 VDD VDD.n14 6.3005
R94 VDD.n20 VDD.t15 6.2405
R95 VDD.n2 VDD.n0 6.2405
R96 VDD.n12 VDD.t5 4.10447
R97 VDD.n16 VDD.t6 3.6405
R98 VDD.n16 VDD.n15 3.6405
R99 VDD.n18 VDD.t14 3.6405
R100 VDD.n18 VDD.n17 3.6405
R101 VDD.n4 VDD.n3 3.1505
R102 VDD.n7 VDD.n6 3.1505
R103 VDD.n6 VDD.n5 3.1505
R104 VDD.n10 VDD.n9 3.1505
R105 VDD.n9 VDD.n8 3.1505
R106 VDD.n13 VDD.n11 3.1505
R107 VDD.n13 VDD.n12 3.1505
R108 VDD.n31 VDD.n14 3.1505
R109 VDD.n34 VDD.n33 3.1505
R110 VDD.n33 VDD.n32 3.1505
R111 VDD.n30 VDD.n29 3.1505
R112 VDD.n29 VDD.n28 3.1505
R113 VDD.n27 VDD.n26 3.1505
R114 VDD.n26 VDD.n25 3.1505
R115 VDD.n24 VDD.n23 3.1505
R116 VDD.n19 VDD.n18 3.06224
R117 VDD.n19 VDD.n16 2.6005
R118 VDD.n4 VDD.n2 0.352424
R119 VDD.n21 VDD.n20 0.340935
R120 VDD.n35 VDD.n19 0.340935
R121 VDD.n23 VDD.n22 0.182033
R122 VDD.n10 VDD.n7 0.0624149
R123 VDD VDD.n11 0.0624149
R124 VDD.n34 VDD.n30 0.0624149
R125 VDD.n27 VDD.n24 0.0624149
R126 VDD.n7 VDD.n4 0.0605
R127 VDD.n11 VDD.n10 0.0605
R128 VDD.n30 VDD.n27 0.0605
R129 VDD.n35 VDD.n34 0.0553936
R130 VDD.n24 VDD.n21 0.0222021
R131 VDD VDD.n35 0.00560638
C0 OUT VDD 0.665f
C1 IN OUT 0.328f
C2 IN VDD 1.14f
.ends

