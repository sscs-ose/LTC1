magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1227 1019 1227
<< metal1 >>
rect -19 221 19 227
rect -19 -221 -13 221
rect 13 -221 19 221
rect -19 -227 19 -221
<< via1 >>
rect -13 -221 13 221
<< metal2 >>
rect -19 221 19 227
rect -19 -221 -13 221
rect 13 -221 19 221
rect -19 -227 19 -221
<< end >>
