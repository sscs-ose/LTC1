magic
tech gf180mcuC
magscale 1 10
timestamp 1714559806
<< nwell >>
rect 236 1820 2544 1837
rect 236 1789 2546 1820
rect 239 1686 2546 1789
rect 239 1665 314 1686
rect 524 1665 2546 1686
rect 239 1638 2546 1665
rect 1190 1279 2173 1638
rect 2180 1637 2546 1638
rect 1322 1217 1499 1279
<< pwell >>
rect 531 1064 693 1122
rect 294 1002 717 1064
rect 1364 856 1497 950
rect 1698 922 2038 1110
<< psubdiff >>
rect 276 771 601 961
rect 276 704 412 771
rect 558 704 601 771
rect 276 684 601 704
rect 879 766 1103 784
rect 879 704 911 766
rect 1066 704 1103 766
rect 879 688 1103 704
rect 1491 763 1715 779
rect 1491 701 1525 763
rect 1680 701 1715 763
rect 1491 683 1715 701
rect 1981 763 2205 781
rect 1981 701 2005 763
rect 2160 701 2205 763
rect 1981 685 2205 701
<< nsubdiff >>
rect 314 1740 524 1760
<< psubdiffcont >>
rect 412 704 558 771
rect 911 704 1066 766
rect 1525 701 1680 763
rect 2005 701 2160 763
<< polysilicon >>
rect 1030 1365 1574 1366
rect 814 1314 1574 1365
rect 814 1265 955 1314
rect 1002 1265 1574 1314
rect 814 1216 1574 1265
rect 2046 1283 2374 1364
rect 2046 1237 2307 1283
rect 2359 1237 2374 1283
rect 2046 1219 2374 1237
rect 898 951 1048 964
rect 805 950 1141 951
rect 805 943 1589 950
rect 805 882 942 943
rect 1011 882 1589 943
rect 805 856 1589 882
rect 2049 917 2385 941
rect 2049 871 2299 917
rect 2346 871 2385 917
rect 2049 828 2385 871
<< polycontact >>
rect 955 1265 1002 1314
rect 2307 1237 2359 1283
rect 942 882 1011 943
rect 2299 871 2346 917
<< metal1 >>
rect 239 1820 2544 1837
rect 239 1656 2546 1820
rect 76 1488 175 1507
rect 76 1433 99 1488
rect 164 1433 175 1488
rect 76 1413 175 1433
rect 730 1414 795 1656
rect 929 1497 1010 1507
rect 929 1423 942 1497
rect 1001 1423 1010 1497
rect 929 1413 1010 1423
rect 1160 1413 1225 1656
rect 78 1299 181 1329
rect 597 1304 671 1319
rect 78 1249 317 1299
rect 78 1229 181 1249
rect 597 1238 603 1304
rect 664 1238 671 1304
rect 945 1314 1010 1413
rect 945 1265 955 1314
rect 1002 1265 1010 1314
rect 1376 1326 1440 1511
rect 1592 1416 1657 1656
rect 1966 1553 2454 1602
rect 1595 1415 1654 1416
rect 1966 1413 2024 1553
rect 1967 1326 2024 1413
rect 1376 1265 2024 1326
rect 2177 1429 2242 1506
rect 2177 1368 2183 1429
rect 2236 1368 2242 1429
rect 2396 1419 2454 1553
rect 2540 1428 2629 1436
rect 945 1249 1010 1265
rect 597 1224 671 1238
rect 1946 1159 2025 1160
rect 1391 1153 2025 1159
rect 1391 1110 1959 1153
rect 77 1085 176 1094
rect 77 1008 87 1085
rect 162 1008 176 1085
rect 929 1066 1025 1082
rect 77 997 176 1008
rect 79 918 179 929
rect 79 845 90 918
rect 169 845 179 918
rect 276 862 601 961
rect 79 834 179 845
rect 234 809 640 862
rect 716 809 781 1055
rect 929 1012 941 1066
rect 1003 1012 1025 1066
rect 929 943 1025 1012
rect 929 882 942 943
rect 1011 882 1025 943
rect 929 873 1025 882
rect 1164 809 1229 1053
rect 1391 990 1453 1110
rect 1946 1100 1959 1110
rect 2012 1100 2025 1153
rect 1946 1089 2025 1100
rect 1612 809 1677 1052
rect 1971 995 2025 1089
rect 2177 980 2242 1368
rect 2540 1373 2552 1428
rect 2617 1373 2629 1428
rect 2540 1364 2629 1373
rect 2294 1305 2373 1306
rect 2293 1286 2373 1305
rect 2293 1232 2304 1286
rect 2362 1232 2373 1286
rect 2293 1220 2373 1232
rect 2294 1219 2373 1220
rect 2408 1161 2492 1170
rect 2408 1100 2420 1161
rect 2480 1100 2492 1161
rect 2408 1093 2492 1100
rect 2410 1038 2464 1093
rect 2410 983 2465 1038
rect 2410 981 2464 983
rect 2281 919 2366 926
rect 2281 864 2293 919
rect 2353 864 2366 919
rect 2281 855 2366 864
rect 234 771 2546 809
rect 234 704 412 771
rect 558 766 2546 771
rect 558 704 911 766
rect 1066 763 2546 766
rect 1066 704 1525 763
rect 234 701 1525 704
rect 1680 701 2005 763
rect 2160 701 2546 763
rect 234 665 2546 701
<< via1 >>
rect 99 1433 164 1488
rect 942 1423 1001 1497
rect 603 1238 664 1304
rect 2183 1368 2236 1429
rect 87 1008 162 1085
rect 90 845 169 918
rect 941 1012 1003 1066
rect 1959 1100 2012 1153
rect 2552 1373 2617 1428
rect 2304 1283 2362 1286
rect 2304 1237 2307 1283
rect 2307 1237 2359 1283
rect 2359 1237 2362 1283
rect 2304 1232 2362 1237
rect 2420 1100 2480 1161
rect 2293 917 2353 919
rect 2293 871 2299 917
rect 2299 871 2346 917
rect 2346 871 2353 917
rect 2293 864 2353 871
<< metal2 >>
rect 76 1497 1010 1507
rect 76 1488 942 1497
rect 76 1433 99 1488
rect 164 1433 942 1488
rect 76 1423 942 1433
rect 1001 1423 1010 1497
rect 76 1413 1010 1423
rect 2163 1436 2254 1449
rect 2163 1429 2629 1436
rect 2163 1368 2183 1429
rect 2236 1428 2629 1429
rect 2236 1373 2552 1428
rect 2617 1373 2629 1428
rect 2236 1368 2629 1373
rect 2163 1364 2629 1368
rect 2163 1356 2254 1364
rect 597 1304 671 1319
rect 597 1238 603 1304
rect 664 1298 671 1304
rect 2294 1298 2373 1306
rect 664 1286 2373 1298
rect 664 1238 2304 1286
rect 597 1232 2304 1238
rect 2362 1232 2373 1286
rect 597 1226 2373 1232
rect 597 1224 671 1226
rect 2294 1219 2373 1226
rect 2408 1161 2492 1170
rect 1946 1157 2025 1160
rect 2408 1157 2420 1161
rect 1946 1153 2420 1157
rect 1946 1100 1959 1153
rect 2012 1101 2420 1153
rect 2012 1100 2025 1101
rect 77 1085 176 1094
rect 1946 1089 2025 1100
rect 2408 1100 2420 1101
rect 2480 1100 2492 1161
rect 2408 1093 2492 1100
rect 77 1008 87 1085
rect 162 1081 176 1085
rect 162 1066 1014 1081
rect 162 1012 941 1066
rect 1003 1012 1014 1066
rect 162 1008 1014 1012
rect 77 1001 1014 1008
rect 77 997 176 1001
rect 937 986 1014 1001
rect 79 926 179 929
rect 79 919 2366 926
rect 79 918 2293 919
rect 79 845 90 918
rect 169 864 2293 918
rect 2353 864 2366 919
rect 169 845 2366 864
rect 79 842 2366 845
rect 79 834 179 842
use inv  inv_0
timestamp 1714553867
transform 1 0 296 0 1 804
box -61 58 345 1035
use nmos_3p3_GYTGVN  nmos_3p3_GYTGVN_0
timestamp 1714126980
transform 1 0 2217 0 1 1010
box -284 -100 284 100
use nmos_3p3_GYTGVN  nmos_3p3_GYTGVN_1
timestamp 1714126980
transform 1 0 973 0 1 1022
box -284 -100 284 100
use nmos_3p3_GYTGVN  nmos_3p3_GYTGVN_2
timestamp 1714126980
transform 1 0 1421 0 1 1022
box -284 -100 284 100
use pmos_3p3_HVHFD7  pmos_3p3_HVHFD7_0
timestamp 1714126980
transform -1 0 1410 0 1 1459
box -338 -180 338 180
use pmos_3p3_HVHFD7  pmos_3p3_HVHFD7_1
timestamp 1714126980
transform 1 0 2210 0 1 1458
box -338 -180 338 180
use pmos_3p3_HVHFD7  pmos_3p3_HVHFD7_2
timestamp 1714126980
transform 1 0 978 0 1 1459
box -338 -180 338 180
<< labels >>
flabel metal1 1323 728 1323 728 0 FreeSans 480 0 0 0 VSS
port 1 nsew
flabel via1 2582 1398 2582 1398 0 FreeSans 480 0 0 0 VCNTL
port 2 nsew
flabel metal1 112 1276 112 1276 0 FreeSans 480 0 0 0 PU
port 3 nsew
flabel via1 112 874 112 874 0 FreeSans 480 0 0 0 PD
port 4 nsew
flabel via1 124 1462 124 1462 0 FreeSans 480 0 0 0 IPD_
port 5 nsew
flabel via1 100 1043 100 1043 0 FreeSans 480 0 0 0 IPD+
port 6 nsew
<< end >>
