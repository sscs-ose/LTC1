magic
tech gf180mcuD
magscale 1 10
timestamp 1713349043
<< checkpaint >>
rect -2184 -3564 3665 2536
<< nwell >>
rect 936 535 1450 536
rect 0 430 1450 535
rect 281 426 1450 430
rect 888 420 1450 426
rect 936 240 1450 420
rect 936 214 1065 240
rect 936 187 1060 214
rect 997 186 1060 187
rect 611 -68 708 0
<< pwell >>
rect 1046 -1225 1055 -505
<< psubdiff >>
rect 502 -1491 641 -1454
rect 502 -1537 545 -1491
rect 591 -1537 641 -1491
rect 502 -1564 641 -1537
<< nsubdiff >>
rect 281 487 888 506
rect 281 441 306 487
rect 822 441 888 487
rect 281 426 888 441
<< psubdiffcont >>
rect 545 -1537 591 -1491
<< nsubdiffcont >>
rect 306 441 822 487
<< polysilicon >>
rect 1166 81 1278 88
rect 174 37 286 39
rect 1166 35 1200 81
rect 1246 35 1278 81
rect 174 -86 286 32
rect 390 -86 502 32
rect 606 -6 718 33
rect 606 -52 637 -6
rect 683 -52 718 -6
rect 606 -86 718 -52
rect 822 -86 934 33
rect 1166 19 1278 35
rect 174 -529 286 -376
rect 390 -447 502 -376
rect 390 -493 407 -447
rect 453 -493 502 -447
rect 390 -529 502 -493
rect 606 -529 718 -376
rect 1165 -388 1278 -375
rect 822 -435 934 -397
rect 820 -450 934 -435
rect 1165 -434 1201 -388
rect 1247 -434 1278 -388
rect 1165 -448 1278 -434
rect 820 -496 834 -450
rect 880 -496 934 -450
rect 820 -529 934 -496
rect 174 -889 286 -841
rect 390 -889 502 -841
rect 1167 -889 1279 -840
rect 174 -1239 286 -1168
rect -87 -1276 286 -1239
rect 388 -1240 718 -1196
rect -87 -1322 -58 -1276
rect -12 -1290 286 -1276
rect 822 -1290 934 -1201
rect 1167 -1224 1279 -1198
rect -12 -1322 934 -1290
rect 1162 -1245 1279 -1224
rect 1162 -1291 1181 -1245
rect 1227 -1291 1279 -1245
rect 1162 -1307 1279 -1291
rect -87 -1351 934 -1322
rect 174 -1385 934 -1351
<< polycontact >>
rect 1200 35 1246 81
rect 637 -52 683 -6
rect 407 -493 453 -447
rect 1201 -434 1247 -388
rect 834 -496 880 -450
rect -58 -1322 -12 -1276
rect 1181 -1291 1227 -1245
<< metal1 >>
rect 88 487 1386 505
rect 88 441 306 487
rect 822 441 1386 487
rect 88 426 1386 441
rect 99 25 145 298
rect 299 206 374 219
rect 299 154 311 206
rect 363 154 374 206
rect 299 140 374 154
rect 531 25 577 298
rect 747 220 793 426
rect 1091 350 1137 426
rect 731 207 807 220
rect 731 155 743 207
rect 795 155 807 207
rect 731 142 807 155
rect -47 4 35 17
rect -89 3 35 4
rect -89 -49 -34 3
rect 18 -49 35 3
rect -89 -52 35 -49
rect -47 -62 35 -52
rect 99 -22 577 25
rect -46 -445 47 -429
rect -112 -446 47 -445
rect -112 -498 -24 -446
rect 28 -498 47 -446
rect -112 -499 47 -498
rect -46 -510 47 -499
rect -81 -1266 15 -1248
rect -184 -1276 15 -1266
rect -184 -1322 -58 -1276
rect -12 -1322 15 -1276
rect -184 -1335 15 -1322
rect -81 -1348 15 -1335
rect 99 -1346 145 -22
rect 300 -232 377 -217
rect 300 -284 312 -232
rect 364 -284 377 -232
rect 300 -297 377 -284
rect 382 -444 479 -422
rect 382 -496 404 -444
rect 456 -496 479 -444
rect 531 -448 577 -22
rect 623 -4 700 13
rect 623 -56 634 -4
rect 686 -56 700 -4
rect 623 -76 700 -56
rect 747 -217 793 142
rect 963 -39 1009 298
rect 1091 130 1135 350
rect 1308 339 1354 426
rect 1308 182 1352 339
rect 1305 93 1354 182
rect 1188 81 1354 93
rect 1188 35 1200 81
rect 1246 35 1354 81
rect 1188 26 1354 35
rect 1188 19 1261 26
rect 963 -86 1665 -39
rect 731 -231 807 -217
rect 731 -283 743 -231
rect 795 -283 807 -231
rect 731 -296 807 -283
rect 747 -352 793 -296
rect 822 -446 892 -435
rect 789 -448 892 -446
rect 531 -450 892 -448
rect 531 -494 834 -450
rect 382 -517 479 -496
rect 789 -496 834 -494
rect 880 -496 892 -450
rect 789 -499 892 -496
rect 822 -510 892 -499
rect 315 -1214 361 -575
rect 531 -842 577 -575
rect 732 -664 808 -650
rect 732 -716 744 -664
rect 796 -716 808 -664
rect 732 -729 808 -716
rect 963 -795 1009 -86
rect 1092 -89 1665 -86
rect 1092 -338 1138 -89
rect 1089 -376 1138 -338
rect 1307 -376 1353 -89
rect 1441 -169 1518 -152
rect 1441 -221 1452 -169
rect 1504 -221 1518 -169
rect 1441 -237 1518 -221
rect 1089 -388 1353 -376
rect 1089 -434 1201 -388
rect 1247 -434 1353 -388
rect 1089 -438 1353 -434
rect 1185 -439 1353 -438
rect 1185 -445 1262 -439
rect 1092 -842 1138 -575
rect 1308 -638 1354 -575
rect 1295 -655 1372 -638
rect 1295 -707 1305 -655
rect 1357 -707 1372 -655
rect 1295 -725 1372 -707
rect 531 -889 1138 -842
rect 531 -1155 577 -889
rect 748 -1214 794 -1114
rect 315 -1260 794 -1214
rect 966 -1346 1012 -1069
rect 1092 -1155 1138 -889
rect 1160 -1243 1250 -1228
rect 1160 -1295 1178 -1243
rect 1230 -1295 1250 -1243
rect 1160 -1311 1250 -1295
rect 99 -1392 1012 -1346
rect 1308 -1442 1354 -725
rect 1446 -1223 1509 -237
rect 1438 -1234 1520 -1223
rect 1438 -1286 1452 -1234
rect 1504 -1286 1520 -1234
rect 1438 -1304 1520 -1286
rect -51 -1491 1427 -1442
rect -51 -1537 545 -1491
rect 591 -1537 1427 -1491
rect -51 -1563 1427 -1537
<< via1 >>
rect 311 154 363 206
rect 743 155 795 207
rect -34 -49 18 3
rect -24 -498 28 -446
rect 312 -284 364 -232
rect 404 -447 456 -444
rect 404 -493 407 -447
rect 407 -493 453 -447
rect 453 -493 456 -447
rect 404 -496 456 -493
rect 634 -6 686 -4
rect 634 -52 637 -6
rect 637 -52 683 -6
rect 683 -52 686 -6
rect 634 -56 686 -52
rect 743 -283 795 -231
rect 744 -716 796 -664
rect 1452 -221 1504 -169
rect 1305 -707 1357 -655
rect 1178 -1245 1230 -1243
rect 1178 -1291 1181 -1245
rect 1181 -1291 1227 -1245
rect 1227 -1291 1230 -1245
rect 1178 -1295 1230 -1291
rect 1452 -1286 1504 -1234
<< metal2 >>
rect 299 212 374 219
rect 731 212 807 220
rect 299 207 807 212
rect 299 206 743 207
rect 299 154 311 206
rect 363 155 743 206
rect 795 155 807 207
rect 363 154 807 155
rect 299 147 807 154
rect 299 140 374 147
rect 731 142 807 147
rect -47 13 35 17
rect -47 4 718 13
rect 1441 4 1511 5
rect -47 3 1511 4
rect -47 -49 -34 3
rect 18 -4 1511 3
rect 18 -49 634 -4
rect -47 -56 634 -49
rect 686 -56 1511 -4
rect -47 -62 35 -56
rect 597 -61 1511 -56
rect 597 -76 718 -61
rect 1441 -152 1511 -61
rect 1441 -169 1518 -152
rect 300 -224 377 -217
rect 731 -224 807 -217
rect 300 -231 807 -224
rect 300 -232 743 -231
rect 300 -284 312 -232
rect 364 -283 743 -232
rect 795 -283 807 -231
rect 1441 -221 1452 -169
rect 1504 -221 1518 -169
rect 1441 -237 1518 -221
rect 364 -284 807 -283
rect 300 -292 807 -284
rect 300 -297 377 -292
rect 731 -296 807 -292
rect 382 -429 479 -422
rect -46 -444 479 -429
rect -46 -446 404 -444
rect -46 -498 -24 -446
rect 28 -496 404 -446
rect 456 -496 479 -444
rect 28 -498 479 -496
rect -46 -510 479 -498
rect 382 -517 479 -510
rect 732 -651 808 -650
rect 1295 -651 1372 -638
rect 732 -655 1372 -651
rect 732 -664 1305 -655
rect 732 -716 744 -664
rect 796 -707 1305 -664
rect 1357 -707 1372 -655
rect 796 -716 1372 -707
rect 732 -721 1372 -716
rect 732 -729 808 -721
rect 1295 -725 1372 -721
rect 1152 -1234 1250 -1224
rect 1438 -1234 1520 -1223
rect 1152 -1243 1452 -1234
rect 1152 -1295 1178 -1243
rect 1230 -1286 1452 -1243
rect 1504 -1286 1520 -1234
rect 1230 -1295 1520 -1286
rect 1152 -1299 1520 -1295
rect 1152 -1309 1250 -1299
rect 1438 -1304 1520 -1299
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_0
timestamp 1713185578
transform 1 0 446 0 1 -685
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_1
timestamp 1713185578
transform 1 0 230 0 1 -685
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_2
timestamp 1713185578
transform 1 0 662 0 1 -685
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_3
timestamp 1713185578
transform 1 0 878 0 1 -685
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_4
timestamp 1713185578
transform 1 0 1223 0 1 -1045
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_5
timestamp 1713185578
transform 1 0 1223 0 1 -685
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_9
timestamp 1713185578
transform 1 0 878 0 1 -1045
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_10
timestamp 1713185578
transform 1 0 662 0 1 -1045
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_11
timestamp 1713185578
transform 1 0 446 0 1 -1045
box -168 -180 168 180
use nmos_3p3_A2UGVV  nmos_3p3_A2UGVV_12
timestamp 1713185578
transform 1 0 230 0 1 -1045
box -168 -180 168 180
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_0
timestamp 1713185578
transform 1 0 878 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_1
timestamp 1713185578
transform 1 0 230 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_2
timestamp 1713185578
transform 1 0 446 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_3
timestamp 1713185578
transform 1 0 662 0 1 -242
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_4
timestamp 1713185578
transform 1 0 878 0 1 188
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_5
timestamp 1713185578
transform 1 0 662 0 1 188
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_6
timestamp 1713185578
transform 1 0 446 0 1 188
box -230 -242 230 242
use pmos_3p3_V9Y6F7  pmos_3p3_V9Y6F7_7
timestamp 1713185578
transform 1 0 230 0 1 188
box -230 -242 230 242
use pmos_3p3_Z9Y6F7  pmos_3p3_Z9Y6F7_0
timestamp 1713185578
transform 1 0 1222 0 1 -242
box -230 -242 230 242
use pmos_3p3_Z9Y6F7  pmos_3p3_Z9Y6F7_1
timestamp 1713185578
transform 1 0 1222 0 1 240
box -230 -242 230 242
<< labels >>
flabel psubdiffcont 567 -1517 567 -1517 0 FreeSans 750 0 0 0 VSS
flabel metal1 s -137 -1305 -137 -1305 0 FreeSans 750 0 0 0 A
port 1 nsew
flabel metal1 s -87 -476 -87 -476 0 FreeSans 750 0 0 0 B
port 2 nsew
flabel metal1 s -72 -29 -72 -29 0 FreeSans 750 0 0 0 C
port 3 nsew
flabel metal1 s 1615 -68 1615 -68 0 FreeSans 750 0 0 0 VOUT
port 4 nsew
flabel metal1 s 653 465 653 465 0 FreeSans 750 0 0 0 VDD
port 5 nsew
<< end >>
