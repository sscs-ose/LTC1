magic
tech gf180mcuC
magscale 1 10
timestamp 1692250459
<< nwell >>
rect -1464 -1307 1464 1307
<< nsubdiff >>
rect -1440 1211 1440 1283
rect -1440 -1211 -1368 1211
rect 1368 -1211 1440 1211
rect -1440 -1283 1440 -1211
<< polysilicon >>
rect -1280 1110 -1120 1123
rect -1280 1064 -1267 1110
rect -1133 1064 -1120 1110
rect -1280 1020 -1120 1064
rect -1280 -1064 -1120 -1020
rect -1280 -1110 -1267 -1064
rect -1133 -1110 -1120 -1064
rect -1280 -1123 -1120 -1110
rect -1040 1110 -880 1123
rect -1040 1064 -1027 1110
rect -893 1064 -880 1110
rect -1040 1020 -880 1064
rect -1040 -1064 -880 -1020
rect -1040 -1110 -1027 -1064
rect -893 -1110 -880 -1064
rect -1040 -1123 -880 -1110
rect -800 1110 -640 1123
rect -800 1064 -787 1110
rect -653 1064 -640 1110
rect -800 1020 -640 1064
rect -800 -1064 -640 -1020
rect -800 -1110 -787 -1064
rect -653 -1110 -640 -1064
rect -800 -1123 -640 -1110
rect -560 1110 -400 1123
rect -560 1064 -547 1110
rect -413 1064 -400 1110
rect -560 1020 -400 1064
rect -560 -1064 -400 -1020
rect -560 -1110 -547 -1064
rect -413 -1110 -400 -1064
rect -560 -1123 -400 -1110
rect -320 1110 -160 1123
rect -320 1064 -307 1110
rect -173 1064 -160 1110
rect -320 1020 -160 1064
rect -320 -1064 -160 -1020
rect -320 -1110 -307 -1064
rect -173 -1110 -160 -1064
rect -320 -1123 -160 -1110
rect -80 1110 80 1123
rect -80 1064 -67 1110
rect 67 1064 80 1110
rect -80 1020 80 1064
rect -80 -1064 80 -1020
rect -80 -1110 -67 -1064
rect 67 -1110 80 -1064
rect -80 -1123 80 -1110
rect 160 1110 320 1123
rect 160 1064 173 1110
rect 307 1064 320 1110
rect 160 1020 320 1064
rect 160 -1064 320 -1020
rect 160 -1110 173 -1064
rect 307 -1110 320 -1064
rect 160 -1123 320 -1110
rect 400 1110 560 1123
rect 400 1064 413 1110
rect 547 1064 560 1110
rect 400 1020 560 1064
rect 400 -1064 560 -1020
rect 400 -1110 413 -1064
rect 547 -1110 560 -1064
rect 400 -1123 560 -1110
rect 640 1110 800 1123
rect 640 1064 653 1110
rect 787 1064 800 1110
rect 640 1020 800 1064
rect 640 -1064 800 -1020
rect 640 -1110 653 -1064
rect 787 -1110 800 -1064
rect 640 -1123 800 -1110
rect 880 1110 1040 1123
rect 880 1064 893 1110
rect 1027 1064 1040 1110
rect 880 1020 1040 1064
rect 880 -1064 1040 -1020
rect 880 -1110 893 -1064
rect 1027 -1110 1040 -1064
rect 880 -1123 1040 -1110
rect 1120 1110 1280 1123
rect 1120 1064 1133 1110
rect 1267 1064 1280 1110
rect 1120 1020 1280 1064
rect 1120 -1064 1280 -1020
rect 1120 -1110 1133 -1064
rect 1267 -1110 1280 -1064
rect 1120 -1123 1280 -1110
<< polycontact >>
rect -1267 1064 -1133 1110
rect -1267 -1110 -1133 -1064
rect -1027 1064 -893 1110
rect -1027 -1110 -893 -1064
rect -787 1064 -653 1110
rect -787 -1110 -653 -1064
rect -547 1064 -413 1110
rect -547 -1110 -413 -1064
rect -307 1064 -173 1110
rect -307 -1110 -173 -1064
rect -67 1064 67 1110
rect -67 -1110 67 -1064
rect 173 1064 307 1110
rect 173 -1110 307 -1064
rect 413 1064 547 1110
rect 413 -1110 547 -1064
rect 653 1064 787 1110
rect 653 -1110 787 -1064
rect 893 1064 1027 1110
rect 893 -1110 1027 -1064
rect 1133 1064 1267 1110
rect 1133 -1110 1267 -1064
<< ppolyres >>
rect -1280 -1020 -1120 1020
rect -1040 -1020 -880 1020
rect -800 -1020 -640 1020
rect -560 -1020 -400 1020
rect -320 -1020 -160 1020
rect -80 -1020 80 1020
rect 160 -1020 320 1020
rect 400 -1020 560 1020
rect 640 -1020 800 1020
rect 880 -1020 1040 1020
rect 1120 -1020 1280 1020
<< metal1 >>
rect -1278 1064 -1267 1110
rect -1133 1064 -1122 1110
rect -1038 1064 -1027 1110
rect -893 1064 -882 1110
rect -798 1064 -787 1110
rect -653 1064 -642 1110
rect -558 1064 -547 1110
rect -413 1064 -402 1110
rect -318 1064 -307 1110
rect -173 1064 -162 1110
rect -78 1064 -67 1110
rect 67 1064 78 1110
rect 162 1064 173 1110
rect 307 1064 318 1110
rect 402 1064 413 1110
rect 547 1064 558 1110
rect 642 1064 653 1110
rect 787 1064 798 1110
rect 882 1064 893 1110
rect 1027 1064 1038 1110
rect 1122 1064 1133 1110
rect 1267 1064 1278 1110
rect -1278 -1110 -1267 -1064
rect -1133 -1110 -1122 -1064
rect -1038 -1110 -1027 -1064
rect -893 -1110 -882 -1064
rect -798 -1110 -787 -1064
rect -653 -1110 -642 -1064
rect -558 -1110 -547 -1064
rect -413 -1110 -402 -1064
rect -318 -1110 -307 -1064
rect -173 -1110 -162 -1064
rect -78 -1110 -67 -1064
rect 67 -1110 78 -1064
rect 162 -1110 173 -1064
rect 307 -1110 318 -1064
rect 402 -1110 413 -1064
rect 547 -1110 558 -1064
rect 642 -1110 653 -1064
rect 787 -1110 798 -1064
rect 882 -1110 893 -1064
rect 1027 -1110 1038 -1064
rect 1122 -1110 1133 -1064
rect 1267 -1110 1278 -1064
<< properties >>
string FIXED_BBOX -1404 -1247 1404 1247
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 10.2 m 1 nx 11 wmin 0.80 lmin 1.00 rho 315 val 4.401k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
