** sch_path: /home/shahid/GF180Projects/Top_test/Decoder_muxes/Xschem/decoder_2x4_PEX_TB_ibr.sym
**.subckt decoder_2x4_PEX_TB_ibr
V1 VDD VSS 3.3
.save i(v1)
V2 VSS GND 0
.save i(v2)
V3 IN1 VSS pulse(3.3 0 0 100p 100p 50n 100n)
.save i(v3)
V4 IN2 VSS pulse(3.3 0 0 100p 100p 100n 200n)
.save i(v4)
x1 IN1 VSS VDD D0 D1 D2 D3 IN2 pex_dec_2x4_ibr_mag
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_dec_2x4_ibr_mag.spice
.control
save all
tran 50p 500n
plot v(IN1) V(IN2)+4 v(D0)+8 v(D1)+12 v(D2)+16 v(D3)+20


*write test_nfet_03v3.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
