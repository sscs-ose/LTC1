magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1075 -1299 1075 1299
<< metal2 >>
rect -75 294 75 299
rect -75 266 -70 294
rect -42 266 -14 294
rect 14 266 42 294
rect 70 266 75 294
rect -75 238 75 266
rect -75 210 -70 238
rect -42 210 -14 238
rect 14 210 42 238
rect 70 210 75 238
rect -75 182 75 210
rect -75 154 -70 182
rect -42 154 -14 182
rect 14 154 42 182
rect 70 154 75 182
rect -75 126 75 154
rect -75 98 -70 126
rect -42 98 -14 126
rect 14 98 42 126
rect 70 98 75 126
rect -75 70 75 98
rect -75 42 -70 70
rect -42 42 -14 70
rect 14 42 42 70
rect 70 42 75 70
rect -75 14 75 42
rect -75 -14 -70 14
rect -42 -14 -14 14
rect 14 -14 42 14
rect 70 -14 75 14
rect -75 -42 75 -14
rect -75 -70 -70 -42
rect -42 -70 -14 -42
rect 14 -70 42 -42
rect 70 -70 75 -42
rect -75 -98 75 -70
rect -75 -126 -70 -98
rect -42 -126 -14 -98
rect 14 -126 42 -98
rect 70 -126 75 -98
rect -75 -154 75 -126
rect -75 -182 -70 -154
rect -42 -182 -14 -154
rect 14 -182 42 -154
rect 70 -182 75 -154
rect -75 -210 75 -182
rect -75 -238 -70 -210
rect -42 -238 -14 -210
rect 14 -238 42 -210
rect 70 -238 75 -210
rect -75 -266 75 -238
rect -75 -294 -70 -266
rect -42 -294 -14 -266
rect 14 -294 42 -266
rect 70 -294 75 -266
rect -75 -299 75 -294
<< via2 >>
rect -70 266 -42 294
rect -14 266 14 294
rect 42 266 70 294
rect -70 210 -42 238
rect -14 210 14 238
rect 42 210 70 238
rect -70 154 -42 182
rect -14 154 14 182
rect 42 154 70 182
rect -70 98 -42 126
rect -14 98 14 126
rect 42 98 70 126
rect -70 42 -42 70
rect -14 42 14 70
rect 42 42 70 70
rect -70 -14 -42 14
rect -14 -14 14 14
rect 42 -14 70 14
rect -70 -70 -42 -42
rect -14 -70 14 -42
rect 42 -70 70 -42
rect -70 -126 -42 -98
rect -14 -126 14 -98
rect 42 -126 70 -98
rect -70 -182 -42 -154
rect -14 -182 14 -154
rect 42 -182 70 -154
rect -70 -238 -42 -210
rect -14 -238 14 -210
rect 42 -238 70 -210
rect -70 -294 -42 -266
rect -14 -294 14 -266
rect 42 -294 70 -266
<< metal3 >>
rect -75 294 75 299
rect -75 266 -70 294
rect -42 266 -14 294
rect 14 266 42 294
rect 70 266 75 294
rect -75 238 75 266
rect -75 210 -70 238
rect -42 210 -14 238
rect 14 210 42 238
rect 70 210 75 238
rect -75 182 75 210
rect -75 154 -70 182
rect -42 154 -14 182
rect 14 154 42 182
rect 70 154 75 182
rect -75 126 75 154
rect -75 98 -70 126
rect -42 98 -14 126
rect 14 98 42 126
rect 70 98 75 126
rect -75 70 75 98
rect -75 42 -70 70
rect -42 42 -14 70
rect 14 42 42 70
rect 70 42 75 70
rect -75 14 75 42
rect -75 -14 -70 14
rect -42 -14 -14 14
rect 14 -14 42 14
rect 70 -14 75 14
rect -75 -42 75 -14
rect -75 -70 -70 -42
rect -42 -70 -14 -42
rect 14 -70 42 -42
rect 70 -70 75 -42
rect -75 -98 75 -70
rect -75 -126 -70 -98
rect -42 -126 -14 -98
rect 14 -126 42 -98
rect 70 -126 75 -98
rect -75 -154 75 -126
rect -75 -182 -70 -154
rect -42 -182 -14 -154
rect 14 -182 42 -154
rect 70 -182 75 -154
rect -75 -210 75 -182
rect -75 -238 -70 -210
rect -42 -238 -14 -210
rect 14 -238 42 -210
rect 70 -238 75 -210
rect -75 -266 75 -238
rect -75 -294 -70 -266
rect -42 -294 -14 -266
rect 14 -294 42 -266
rect 70 -294 75 -266
rect -75 -299 75 -294
<< end >>
