magic
tech gf180mcuC
magscale 1 10
timestamp 1714534647
<< nwell >>
rect 36 631 330 669
rect -122 579 330 631
rect 36 502 330 579
<< psubdiff >>
rect -80 -95 236 -82
rect -80 -141 -67 -95
rect 223 -141 236 -95
rect -80 -154 236 -141
<< nsubdiff >>
rect 69 622 306 636
rect 69 576 231 622
rect 277 576 306 622
rect 69 559 306 576
<< psubdiffcont >>
rect -67 -141 223 -95
<< nsubdiffcont >>
rect 231 576 277 622
<< polysilicon >>
rect -44 187 156 250
rect -44 141 31 187
rect 87 141 156 187
rect -44 103 156 141
<< polycontact >>
rect 31 141 87 187
<< metal1 >>
rect 69 631 306 636
rect -122 622 330 631
rect -122 576 231 622
rect 277 576 330 622
rect -122 522 330 576
rect -122 292 -59 522
rect -118 187 93 200
rect -118 141 31 187
rect 87 141 93 187
rect -118 128 93 141
rect 179 189 242 450
rect 179 131 286 189
rect -134 -69 -67 60
rect 179 14 242 131
rect -134 -95 286 -69
rect -134 -141 -67 -95
rect 223 -141 286 -95
rect -134 -175 286 -141
use nmos_3p3_MGBSF7  nmos_3p3_MGBSF7_0
timestamp 1714126980
transform 1 0 56 0 1 37
box -216 -97 216 97
use pmos_3p3_MW53B7  pmos_3p3_MW53B7_0
timestamp 1714126980
transform 1 0 56 0 1 369
box -274 -210 274 210
<< labels >>
flabel psubdiffcont 80 -120 80 -120 0 FreeSans 640 0 0 0 VSS
port 1 nsew
flabel metal1 -106 158 -106 158 0 FreeSans 640 0 0 0 IN
port 2 nsew
flabel metal1 276 159 276 159 0 FreeSans 640 0 0 0 OUT
port 3 nsew
flabel nsubdiffcont 251 601 251 601 0 FreeSans 640 0 0 0 VDD
port 4 nsew
<< end >>
