magic
tech gf180mcuC
magscale 1 10
timestamp 1692949218
<< error_p >>
rect -3306 -3722 -3267 -3716
rect -3221 -3722 -3182 -3716
rect -3306 -3740 -3182 -3722
rect -1330 -3722 -1291 -3716
rect -1245 -3722 -1206 -3716
rect -1330 -3740 -1206 -3722
rect -3282 -3764 -3206 -3740
rect -1306 -3764 -1230 -3740
rect -2438 -4035 -2370 -3968
rect -3282 -4250 -3206 -4226
rect -1306 -4250 -1230 -4226
rect -3306 -4274 -3182 -4250
rect -1330 -4274 -1206 -4250
<< nwell >>
rect -3327 -4250 -1192 -3740
<< pdiff >>
rect -2438 -4035 -2370 -3968
<< nsubdiff >>
rect -3282 -3768 -3267 -3740
rect -3221 -3768 -3206 -3740
rect -3282 -3816 -3206 -3768
rect -3282 -3862 -3267 -3816
rect -3221 -3862 -3206 -3816
rect -3282 -3910 -3206 -3862
rect -3282 -3956 -3267 -3910
rect -3221 -3956 -3206 -3910
rect -3282 -4004 -3206 -3956
rect -1306 -3768 -1291 -3740
rect -1245 -3768 -1230 -3740
rect -1306 -3816 -1230 -3768
rect -1306 -3862 -1291 -3816
rect -1245 -3862 -1230 -3816
rect -1306 -3910 -1230 -3862
rect -1306 -3956 -1291 -3910
rect -1245 -3956 -1230 -3910
rect -3282 -4050 -3267 -4004
rect -3221 -4050 -3206 -4004
rect -1306 -4004 -1230 -3956
rect -3282 -4098 -3206 -4050
rect -3282 -4144 -3267 -4098
rect -3221 -4144 -3206 -4098
rect -3282 -4192 -3206 -4144
rect -3282 -4238 -3267 -4192
rect -3221 -4238 -3206 -4192
rect -3282 -4250 -3206 -4238
rect -1306 -4050 -1291 -4004
rect -1245 -4050 -1230 -4004
rect -1306 -4098 -1230 -4050
rect -1306 -4144 -1291 -4098
rect -1245 -4144 -1230 -4098
rect -1306 -4192 -1230 -4144
rect -1306 -4238 -1291 -4192
rect -1245 -4238 -1230 -4192
rect -1306 -4250 -1230 -4238
<< nsubdiffcont >>
rect -3267 -3768 -3221 -3740
rect -3267 -3862 -3221 -3816
rect -3267 -3956 -3221 -3910
rect -1291 -3768 -1245 -3740
rect -1291 -3862 -1245 -3816
rect -1291 -3956 -1245 -3910
rect -3267 -4050 -3221 -4004
rect -3267 -4144 -3221 -4098
rect -3267 -4238 -3221 -4192
rect -1291 -4050 -1245 -4004
rect -1291 -4144 -1245 -4098
rect -1291 -4238 -1245 -4192
<< metal1 >>
rect -3293 -3768 -3267 -3740
rect -3221 -3768 -3195 -3740
rect -3293 -3816 -3195 -3768
rect -1317 -3768 -1291 -3740
rect -1245 -3768 -1219 -3740
rect -3293 -3862 -3267 -3816
rect -3221 -3862 -3195 -3816
rect -3293 -3910 -3195 -3862
rect -2607 -3822 -2524 -3808
rect -2607 -3878 -2593 -3822
rect -2537 -3878 -2524 -3822
rect -2607 -3890 -2524 -3878
rect -1965 -3822 -1882 -3809
rect -1965 -3878 -1952 -3822
rect -1896 -3878 -1882 -3822
rect -1965 -3891 -1882 -3878
rect -1317 -3816 -1219 -3768
rect -1317 -3862 -1291 -3816
rect -1245 -3862 -1219 -3816
rect -3293 -3956 -3267 -3910
rect -3221 -3956 -3195 -3910
rect -1317 -3910 -1219 -3862
rect -3293 -4004 -3195 -3956
rect -3293 -4050 -3267 -4004
rect -3221 -4050 -3195 -4004
rect -2767 -3975 -2684 -3961
rect -2767 -4031 -2753 -3975
rect -2697 -4031 -2684 -3975
rect -2767 -4043 -2684 -4031
rect -2453 -3968 -2354 -3953
rect -1317 -3956 -1291 -3910
rect -1245 -3956 -1219 -3910
rect -2453 -4035 -2438 -3968
rect -2370 -4035 -2354 -3968
rect -2453 -4046 -2354 -4035
rect -2126 -3974 -2043 -3960
rect -2126 -4030 -2112 -3974
rect -2056 -4030 -2043 -3974
rect -2126 -4042 -2043 -4030
rect -1806 -3975 -1723 -3961
rect -1806 -4031 -1792 -3975
rect -1736 -4031 -1723 -3975
rect -1806 -4043 -1723 -4031
rect -1317 -4004 -1219 -3956
rect -3293 -4098 -3195 -4050
rect -3293 -4144 -3267 -4098
rect -3221 -4144 -3195 -4098
rect -1317 -4050 -1291 -4004
rect -1245 -4050 -1219 -4004
rect -1317 -4098 -1219 -4050
rect -3293 -4192 -3195 -4144
rect -3293 -4238 -3267 -4192
rect -3221 -4238 -3195 -4192
rect -3088 -4134 -3004 -4120
rect -3088 -4190 -3074 -4134
rect -3018 -4190 -3004 -4134
rect -3088 -4204 -3004 -4190
rect -2927 -4134 -2843 -4119
rect -2927 -4190 -2913 -4134
rect -2857 -4190 -2843 -4134
rect -2927 -4203 -2843 -4190
rect -2288 -4134 -2202 -4120
rect -2288 -4190 -2274 -4134
rect -2216 -4190 -2202 -4134
rect -2288 -4204 -2202 -4190
rect -1647 -4134 -1563 -4119
rect -1647 -4190 -1633 -4134
rect -1577 -4190 -1563 -4134
rect -1647 -4203 -1563 -4190
rect -1487 -4134 -1403 -4120
rect -1487 -4190 -1473 -4134
rect -1417 -4190 -1403 -4134
rect -1487 -4204 -1403 -4190
rect -1317 -4144 -1291 -4098
rect -1245 -4121 -1219 -4098
rect -1245 -4144 -1120 -4121
rect -1317 -4192 -1120 -4144
rect -3293 -4250 -3195 -4238
rect -1317 -4238 -1291 -4192
rect -1245 -4238 -1120 -4192
rect -1317 -4250 -1120 -4238
<< via1 >>
rect -2593 -3878 -2537 -3822
rect -1952 -3878 -1896 -3822
rect -2753 -4031 -2697 -3975
rect -2438 -4035 -2370 -3968
rect -2112 -4030 -2056 -3974
rect -1792 -4031 -1736 -3975
rect -3074 -4190 -3018 -4134
rect -2913 -4190 -2857 -4134
rect -2274 -4190 -2216 -4134
rect -1633 -4190 -1577 -4134
rect -1473 -4190 -1417 -4134
<< metal2 >>
rect -3472 -3973 -3352 -3740
rect -2524 -3808 -2332 -3806
rect -2607 -3819 -2332 -3808
rect -2607 -3822 -2510 -3819
rect -2607 -3878 -2593 -3822
rect -2537 -3875 -2510 -3822
rect -2454 -3875 -2400 -3819
rect -2344 -3820 -2332 -3819
rect -1965 -3820 -1882 -3809
rect -2344 -3822 -1882 -3820
rect -2344 -3875 -1952 -3822
rect -2537 -3878 -1952 -3875
rect -1896 -3878 -1882 -3822
rect -2607 -3880 -1882 -3878
rect -2607 -3890 -2332 -3880
rect -1965 -3891 -1882 -3880
rect -2767 -3973 -2684 -3961
rect -2453 -3968 -2354 -3953
rect -2453 -3973 -2438 -3968
rect -3472 -3975 -2438 -3973
rect -3472 -4031 -2753 -3975
rect -2697 -4031 -2438 -3975
rect -3472 -4034 -2438 -4031
rect -3472 -4250 -3352 -4034
rect -2767 -4043 -2684 -4034
rect -2453 -4035 -2438 -4034
rect -2370 -3973 -2354 -3968
rect -2126 -3973 -2043 -3960
rect -1806 -3973 -1723 -3961
rect -2370 -3974 -1723 -3973
rect -2370 -4030 -2112 -3974
rect -2056 -3975 -1723 -3974
rect -2056 -4030 -1792 -3975
rect -2370 -4031 -1792 -4030
rect -1736 -4031 -1723 -3975
rect -2370 -4034 -1723 -4031
rect -2370 -4035 -2354 -4034
rect -2453 -4046 -2354 -4035
rect -2126 -4042 -2043 -4034
rect -1806 -4043 -1723 -4034
rect -3088 -4132 -3004 -4120
rect -2927 -4132 -2843 -4119
rect -2288 -4132 -2202 -4120
rect -2121 -4131 -1929 -4118
rect -2121 -4132 -2107 -4131
rect -3088 -4134 -2107 -4132
rect -3088 -4190 -3074 -4134
rect -3018 -4190 -2913 -4134
rect -2857 -4190 -2274 -4134
rect -2216 -4187 -2107 -4134
rect -2051 -4187 -1997 -4131
rect -1941 -4132 -1929 -4131
rect -1647 -4132 -1563 -4119
rect -1487 -4132 -1403 -4120
rect -1941 -4134 -1403 -4132
rect -1941 -4187 -1633 -4134
rect -2216 -4190 -1633 -4187
rect -1577 -4190 -1473 -4134
rect -1417 -4190 -1403 -4134
rect -3088 -4192 -1403 -4190
rect -3088 -4204 -3004 -4192
rect -2927 -4203 -2843 -4192
rect -2288 -4204 -2202 -4192
rect -2121 -4202 -1929 -4192
rect -1647 -4203 -1563 -4192
rect -1487 -4204 -1403 -4192
<< via2 >>
rect -2510 -3875 -2454 -3819
rect -2400 -3875 -2344 -3819
rect -2107 -4187 -2051 -4131
rect -1997 -4187 -1941 -4131
<< metal3 >>
rect -2833 -4250 -2767 -3740
rect -2458 -3806 -2392 -3740
rect -2524 -3819 -2332 -3806
rect -2524 -3875 -2510 -3819
rect -2454 -3875 -2400 -3819
rect -2344 -3875 -2332 -3819
rect -2524 -3890 -2332 -3875
rect -2458 -4250 -2392 -3890
rect -2097 -4118 -2031 -3740
rect -2121 -4131 -1929 -4118
rect -2121 -4187 -2107 -4131
rect -2051 -4187 -1997 -4131
rect -1941 -4187 -1929 -4131
rect -2121 -4202 -1929 -4187
rect -2097 -4250 -2031 -4202
rect -1726 -4250 -1660 -3740
<< end >>
