magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2195 -6145 2195 6145
<< psubdiff >>
rect -195 4123 195 4145
rect -195 -4123 -173 4123
rect 173 -4123 195 4123
rect -195 -4145 195 -4123
<< psubdiffcont >>
rect -173 -4123 173 4123
<< metal1 >>
rect -184 4123 184 4134
rect -184 -4123 -173 4123
rect 173 -4123 184 4123
rect -184 -4134 184 -4123
<< end >>
