magic
tech gf180mcuC
magscale 1 10
timestamp 1693543231
<< pwell >>
rect 0 1734 4200 2070
rect 0 1283 4200 1619
rect 0 519 4200 855
rect 0 71 4200 407
<< nmos >>
rect 112 1802 212 2002
rect 316 1802 416 2002
rect 520 1802 620 2002
rect 724 1802 824 2002
rect 928 1802 1028 2002
rect 1132 1802 1232 2002
rect 1336 1802 1436 2002
rect 1540 1802 1640 2002
rect 1744 1802 1844 2002
rect 1948 1802 2048 2002
rect 2152 1802 2252 2002
rect 2356 1802 2456 2002
rect 2560 1802 2660 2002
rect 2764 1802 2864 2002
rect 2968 1802 3068 2002
rect 3172 1802 3272 2002
rect 3376 1802 3476 2002
rect 3580 1802 3680 2002
rect 3784 1802 3884 2002
rect 3988 1802 4088 2002
rect 112 1351 212 1551
rect 316 1351 416 1551
rect 520 1351 620 1551
rect 724 1351 824 1551
rect 928 1351 1028 1551
rect 1132 1351 1232 1551
rect 1336 1351 1436 1551
rect 1540 1351 1640 1551
rect 1744 1351 1844 1551
rect 1948 1351 2048 1551
rect 2152 1351 2252 1551
rect 2356 1351 2456 1551
rect 2560 1351 2660 1551
rect 2764 1351 2864 1551
rect 2968 1351 3068 1551
rect 3172 1351 3272 1551
rect 3376 1351 3476 1551
rect 3580 1351 3680 1551
rect 3784 1351 3884 1551
rect 3988 1351 4088 1551
rect 112 587 212 787
rect 316 587 416 787
rect 520 587 620 787
rect 724 587 824 787
rect 928 587 1028 787
rect 1132 587 1232 787
rect 1336 587 1436 787
rect 1540 587 1640 787
rect 1744 587 1844 787
rect 1948 587 2048 787
rect 2152 587 2252 787
rect 2356 587 2456 787
rect 2560 587 2660 787
rect 2764 587 2864 787
rect 2968 587 3068 787
rect 3172 587 3272 787
rect 3376 587 3476 787
rect 3580 587 3680 787
rect 3784 587 3884 787
rect 3988 587 4088 787
rect 112 139 212 339
rect 316 139 416 339
rect 520 139 620 339
rect 724 139 824 339
rect 928 139 1028 339
rect 1132 139 1232 339
rect 1336 139 1436 339
rect 1540 139 1640 339
rect 1744 139 1844 339
rect 1948 139 2048 339
rect 2152 139 2252 339
rect 2356 139 2456 339
rect 2560 139 2660 339
rect 2764 139 2864 339
rect 2968 139 3068 339
rect 3172 139 3272 339
rect 3376 139 3476 339
rect 3580 139 3680 339
rect 3784 139 3884 339
rect 3988 139 4088 339
<< ndiff >>
rect 24 1989 112 2002
rect 24 1815 37 1989
rect 83 1815 112 1989
rect 24 1802 112 1815
rect 212 1989 316 2002
rect 212 1815 241 1989
rect 287 1815 316 1989
rect 212 1802 316 1815
rect 416 1989 520 2002
rect 416 1815 445 1989
rect 491 1815 520 1989
rect 416 1802 520 1815
rect 620 1989 724 2002
rect 620 1815 649 1989
rect 695 1815 724 1989
rect 620 1802 724 1815
rect 824 1989 928 2002
rect 824 1815 853 1989
rect 899 1815 928 1989
rect 824 1802 928 1815
rect 1028 1989 1132 2002
rect 1028 1815 1057 1989
rect 1103 1815 1132 1989
rect 1028 1802 1132 1815
rect 1232 1989 1336 2002
rect 1232 1815 1261 1989
rect 1307 1815 1336 1989
rect 1232 1802 1336 1815
rect 1436 1989 1540 2002
rect 1436 1815 1465 1989
rect 1511 1815 1540 1989
rect 1436 1802 1540 1815
rect 1640 1989 1744 2002
rect 1640 1815 1669 1989
rect 1715 1815 1744 1989
rect 1640 1802 1744 1815
rect 1844 1989 1948 2002
rect 1844 1815 1873 1989
rect 1919 1815 1948 1989
rect 1844 1802 1948 1815
rect 2048 1989 2152 2002
rect 2048 1815 2077 1989
rect 2123 1815 2152 1989
rect 2048 1802 2152 1815
rect 2252 1989 2356 2002
rect 2252 1815 2281 1989
rect 2327 1815 2356 1989
rect 2252 1802 2356 1815
rect 2456 1989 2560 2002
rect 2456 1815 2485 1989
rect 2531 1815 2560 1989
rect 2456 1802 2560 1815
rect 2660 1989 2764 2002
rect 2660 1815 2689 1989
rect 2735 1815 2764 1989
rect 2660 1802 2764 1815
rect 2864 1989 2968 2002
rect 2864 1815 2893 1989
rect 2939 1815 2968 1989
rect 2864 1802 2968 1815
rect 3068 1989 3172 2002
rect 3068 1815 3097 1989
rect 3143 1815 3172 1989
rect 3068 1802 3172 1815
rect 3272 1989 3376 2002
rect 3272 1815 3301 1989
rect 3347 1815 3376 1989
rect 3272 1802 3376 1815
rect 3476 1989 3580 2002
rect 3476 1815 3505 1989
rect 3551 1815 3580 1989
rect 3476 1802 3580 1815
rect 3680 1989 3784 2002
rect 3680 1815 3709 1989
rect 3755 1815 3784 1989
rect 3680 1802 3784 1815
rect 3884 1989 3988 2002
rect 3884 1815 3913 1989
rect 3959 1815 3988 1989
rect 3884 1802 3988 1815
rect 4088 1989 4176 2002
rect 4088 1815 4117 1989
rect 4163 1815 4176 1989
rect 4088 1802 4176 1815
rect 24 1538 112 1551
rect 24 1364 37 1538
rect 83 1364 112 1538
rect 24 1351 112 1364
rect 212 1538 316 1551
rect 212 1364 241 1538
rect 287 1364 316 1538
rect 212 1351 316 1364
rect 416 1538 520 1551
rect 416 1364 445 1538
rect 491 1364 520 1538
rect 416 1351 520 1364
rect 620 1538 724 1551
rect 620 1364 649 1538
rect 695 1364 724 1538
rect 620 1351 724 1364
rect 824 1538 928 1551
rect 824 1364 853 1538
rect 899 1364 928 1538
rect 824 1351 928 1364
rect 1028 1538 1132 1551
rect 1028 1364 1057 1538
rect 1103 1364 1132 1538
rect 1028 1351 1132 1364
rect 1232 1538 1336 1551
rect 1232 1364 1261 1538
rect 1307 1364 1336 1538
rect 1232 1351 1336 1364
rect 1436 1538 1540 1551
rect 1436 1364 1465 1538
rect 1511 1364 1540 1538
rect 1436 1351 1540 1364
rect 1640 1538 1744 1551
rect 1640 1364 1669 1538
rect 1715 1364 1744 1538
rect 1640 1351 1744 1364
rect 1844 1538 1948 1551
rect 1844 1364 1873 1538
rect 1919 1364 1948 1538
rect 1844 1351 1948 1364
rect 2048 1538 2152 1551
rect 2048 1364 2077 1538
rect 2123 1364 2152 1538
rect 2048 1351 2152 1364
rect 2252 1538 2356 1551
rect 2252 1364 2281 1538
rect 2327 1364 2356 1538
rect 2252 1351 2356 1364
rect 2456 1538 2560 1551
rect 2456 1364 2485 1538
rect 2531 1364 2560 1538
rect 2456 1351 2560 1364
rect 2660 1538 2764 1551
rect 2660 1364 2689 1538
rect 2735 1364 2764 1538
rect 2660 1351 2764 1364
rect 2864 1538 2968 1551
rect 2864 1364 2893 1538
rect 2939 1364 2968 1538
rect 2864 1351 2968 1364
rect 3068 1538 3172 1551
rect 3068 1364 3097 1538
rect 3143 1364 3172 1538
rect 3068 1351 3172 1364
rect 3272 1538 3376 1551
rect 3272 1364 3301 1538
rect 3347 1364 3376 1538
rect 3272 1351 3376 1364
rect 3476 1538 3580 1551
rect 3476 1364 3505 1538
rect 3551 1364 3580 1538
rect 3476 1351 3580 1364
rect 3680 1538 3784 1551
rect 3680 1364 3709 1538
rect 3755 1364 3784 1538
rect 3680 1351 3784 1364
rect 3884 1538 3988 1551
rect 3884 1364 3913 1538
rect 3959 1364 3988 1538
rect 3884 1351 3988 1364
rect 4088 1538 4176 1551
rect 4088 1364 4117 1538
rect 4163 1364 4176 1538
rect 4088 1351 4176 1364
rect 24 774 112 787
rect 24 600 37 774
rect 83 600 112 774
rect 24 587 112 600
rect 212 774 316 787
rect 212 600 241 774
rect 287 600 316 774
rect 212 587 316 600
rect 416 774 520 787
rect 416 600 445 774
rect 491 600 520 774
rect 416 587 520 600
rect 620 774 724 787
rect 620 600 649 774
rect 695 600 724 774
rect 620 587 724 600
rect 824 774 928 787
rect 824 600 853 774
rect 899 600 928 774
rect 824 587 928 600
rect 1028 774 1132 787
rect 1028 600 1057 774
rect 1103 600 1132 774
rect 1028 587 1132 600
rect 1232 774 1336 787
rect 1232 600 1261 774
rect 1307 600 1336 774
rect 1232 587 1336 600
rect 1436 774 1540 787
rect 1436 600 1465 774
rect 1511 600 1540 774
rect 1436 587 1540 600
rect 1640 774 1744 787
rect 1640 600 1669 774
rect 1715 600 1744 774
rect 1640 587 1744 600
rect 1844 774 1948 787
rect 1844 600 1873 774
rect 1919 600 1948 774
rect 1844 587 1948 600
rect 2048 774 2152 787
rect 2048 600 2077 774
rect 2123 600 2152 774
rect 2048 587 2152 600
rect 2252 774 2356 787
rect 2252 600 2281 774
rect 2327 600 2356 774
rect 2252 587 2356 600
rect 2456 774 2560 787
rect 2456 600 2485 774
rect 2531 600 2560 774
rect 2456 587 2560 600
rect 2660 774 2764 787
rect 2660 600 2689 774
rect 2735 600 2764 774
rect 2660 587 2764 600
rect 2864 774 2968 787
rect 2864 600 2893 774
rect 2939 600 2968 774
rect 2864 587 2968 600
rect 3068 774 3172 787
rect 3068 600 3097 774
rect 3143 600 3172 774
rect 3068 587 3172 600
rect 3272 774 3376 787
rect 3272 600 3301 774
rect 3347 600 3376 774
rect 3272 587 3376 600
rect 3476 774 3580 787
rect 3476 600 3505 774
rect 3551 600 3580 774
rect 3476 587 3580 600
rect 3680 774 3784 787
rect 3680 600 3709 774
rect 3755 600 3784 774
rect 3680 587 3784 600
rect 3884 774 3988 787
rect 3884 600 3913 774
rect 3959 600 3988 774
rect 3884 587 3988 600
rect 4088 774 4176 787
rect 4088 600 4117 774
rect 4163 600 4176 774
rect 4088 587 4176 600
rect 24 326 112 339
rect 24 152 37 326
rect 83 152 112 326
rect 24 139 112 152
rect 212 326 316 339
rect 212 152 241 326
rect 287 152 316 326
rect 212 139 316 152
rect 416 326 520 339
rect 416 152 445 326
rect 491 152 520 326
rect 416 139 520 152
rect 620 326 724 339
rect 620 152 649 326
rect 695 152 724 326
rect 620 139 724 152
rect 824 326 928 339
rect 824 152 853 326
rect 899 152 928 326
rect 824 139 928 152
rect 1028 326 1132 339
rect 1028 152 1057 326
rect 1103 152 1132 326
rect 1028 139 1132 152
rect 1232 326 1336 339
rect 1232 152 1261 326
rect 1307 152 1336 326
rect 1232 139 1336 152
rect 1436 326 1540 339
rect 1436 152 1465 326
rect 1511 152 1540 326
rect 1436 139 1540 152
rect 1640 326 1744 339
rect 1640 152 1669 326
rect 1715 152 1744 326
rect 1640 139 1744 152
rect 1844 326 1948 339
rect 1844 152 1873 326
rect 1919 152 1948 326
rect 1844 139 1948 152
rect 2048 326 2152 339
rect 2048 152 2077 326
rect 2123 152 2152 326
rect 2048 139 2152 152
rect 2252 326 2356 339
rect 2252 152 2281 326
rect 2327 152 2356 326
rect 2252 139 2356 152
rect 2456 326 2560 339
rect 2456 152 2485 326
rect 2531 152 2560 326
rect 2456 139 2560 152
rect 2660 326 2764 339
rect 2660 152 2689 326
rect 2735 152 2764 326
rect 2660 139 2764 152
rect 2864 326 2968 339
rect 2864 152 2893 326
rect 2939 152 2968 326
rect 2864 139 2968 152
rect 3068 326 3172 339
rect 3068 152 3097 326
rect 3143 152 3172 326
rect 3068 139 3172 152
rect 3272 326 3376 339
rect 3272 152 3301 326
rect 3347 152 3376 326
rect 3272 139 3376 152
rect 3476 326 3580 339
rect 3476 152 3505 326
rect 3551 152 3580 326
rect 3476 139 3580 152
rect 3680 326 3784 339
rect 3680 152 3709 326
rect 3755 152 3784 326
rect 3680 139 3784 152
rect 3884 326 3988 339
rect 3884 152 3913 326
rect 3959 152 3988 326
rect 3884 139 3988 152
rect 4088 326 4176 339
rect 4088 152 4117 326
rect 4163 152 4176 326
rect 4088 139 4176 152
<< ndiffc >>
rect 37 1815 83 1989
rect 241 1815 287 1989
rect 445 1815 491 1989
rect 649 1815 695 1989
rect 853 1815 899 1989
rect 1057 1815 1103 1989
rect 1261 1815 1307 1989
rect 1465 1815 1511 1989
rect 1669 1815 1715 1989
rect 1873 1815 1919 1989
rect 2077 1815 2123 1989
rect 2281 1815 2327 1989
rect 2485 1815 2531 1989
rect 2689 1815 2735 1989
rect 2893 1815 2939 1989
rect 3097 1815 3143 1989
rect 3301 1815 3347 1989
rect 3505 1815 3551 1989
rect 3709 1815 3755 1989
rect 3913 1815 3959 1989
rect 4117 1815 4163 1989
rect 37 1364 83 1538
rect 241 1364 287 1538
rect 445 1364 491 1538
rect 649 1364 695 1538
rect 853 1364 899 1538
rect 1057 1364 1103 1538
rect 1261 1364 1307 1538
rect 1465 1364 1511 1538
rect 1669 1364 1715 1538
rect 1873 1364 1919 1538
rect 2077 1364 2123 1538
rect 2281 1364 2327 1538
rect 2485 1364 2531 1538
rect 2689 1364 2735 1538
rect 2893 1364 2939 1538
rect 3097 1364 3143 1538
rect 3301 1364 3347 1538
rect 3505 1364 3551 1538
rect 3709 1364 3755 1538
rect 3913 1364 3959 1538
rect 4117 1364 4163 1538
rect 37 600 83 774
rect 241 600 287 774
rect 445 600 491 774
rect 649 600 695 774
rect 853 600 899 774
rect 1057 600 1103 774
rect 1261 600 1307 774
rect 1465 600 1511 774
rect 1669 600 1715 774
rect 1873 600 1919 774
rect 2077 600 2123 774
rect 2281 600 2327 774
rect 2485 600 2531 774
rect 2689 600 2735 774
rect 2893 600 2939 774
rect 3097 600 3143 774
rect 3301 600 3347 774
rect 3505 600 3551 774
rect 3709 600 3755 774
rect 3913 600 3959 774
rect 4117 600 4163 774
rect 37 152 83 326
rect 241 152 287 326
rect 445 152 491 326
rect 649 152 695 326
rect 853 152 899 326
rect 1057 152 1103 326
rect 1261 152 1307 326
rect 1465 152 1511 326
rect 1669 152 1715 326
rect 1873 152 1919 326
rect 2077 152 2123 326
rect 2281 152 2327 326
rect 2485 152 2531 326
rect 2689 152 2735 326
rect 2893 152 2939 326
rect 3097 152 3143 326
rect 3301 152 3347 326
rect 3505 152 3551 326
rect 3709 152 3755 326
rect 3913 152 3959 326
rect 4117 152 4163 326
<< psubdiff >>
rect 0 2341 128 2357
rect 0 2230 17 2341
rect 111 2230 128 2341
rect 0 2211 128 2230
rect 210 2341 338 2357
rect 210 2230 227 2341
rect 321 2230 338 2341
rect 210 2211 338 2230
rect 420 2341 548 2357
rect 420 2230 437 2341
rect 531 2230 548 2341
rect 420 2211 548 2230
rect 630 2341 758 2357
rect 630 2230 647 2341
rect 741 2230 758 2341
rect 630 2211 758 2230
rect 840 2341 968 2357
rect 840 2230 857 2341
rect 951 2230 968 2341
rect 840 2211 968 2230
rect 1050 2341 1178 2357
rect 1050 2230 1067 2341
rect 1161 2230 1178 2341
rect 1050 2211 1178 2230
rect 1260 2341 1388 2357
rect 1260 2230 1277 2341
rect 1371 2230 1388 2341
rect 1260 2211 1388 2230
rect 1470 2341 1598 2357
rect 1470 2230 1487 2341
rect 1581 2230 1598 2341
rect 1470 2211 1598 2230
rect 1680 2341 1808 2357
rect 1680 2230 1697 2341
rect 1791 2230 1808 2341
rect 1680 2211 1808 2230
rect 1890 2341 2018 2357
rect 1890 2230 1907 2341
rect 2001 2230 2018 2341
rect 1890 2211 2018 2230
rect 2100 2341 2228 2357
rect 2100 2230 2117 2341
rect 2211 2230 2228 2341
rect 2100 2211 2228 2230
rect 2310 2341 2438 2357
rect 2310 2230 2327 2341
rect 2421 2230 2438 2341
rect 2310 2211 2438 2230
rect 2520 2341 2648 2357
rect 2520 2230 2537 2341
rect 2631 2230 2648 2341
rect 2520 2211 2648 2230
rect 2730 2341 2858 2357
rect 2730 2230 2747 2341
rect 2841 2230 2858 2341
rect 2730 2211 2858 2230
rect 2940 2341 3068 2357
rect 2940 2230 2957 2341
rect 3051 2230 3068 2341
rect 2940 2211 3068 2230
rect 3150 2341 3278 2357
rect 3150 2230 3167 2341
rect 3261 2230 3278 2341
rect 3150 2211 3278 2230
rect 3360 2341 3488 2357
rect 3360 2230 3377 2341
rect 3471 2230 3488 2341
rect 3360 2211 3488 2230
rect 3570 2341 3698 2357
rect 3570 2230 3587 2341
rect 3681 2230 3698 2341
rect 3570 2211 3698 2230
rect 3780 2341 3908 2357
rect 3780 2230 3797 2341
rect 3891 2230 3908 2341
rect 3780 2211 3908 2230
rect 3990 2341 4118 2357
rect 3990 2230 4007 2341
rect 4101 2230 4118 2341
rect 3990 2211 4118 2230
rect 0 1126 128 1142
rect 0 1015 17 1126
rect 111 1015 128 1126
rect 0 996 128 1015
rect 210 1126 338 1142
rect 210 1015 227 1126
rect 321 1015 338 1126
rect 210 996 338 1015
rect 420 1126 548 1142
rect 420 1015 437 1126
rect 531 1015 548 1126
rect 420 996 548 1015
rect 630 1126 758 1142
rect 630 1015 647 1126
rect 741 1015 758 1126
rect 630 996 758 1015
rect 840 1126 968 1142
rect 840 1015 857 1126
rect 951 1015 968 1126
rect 840 996 968 1015
rect 1050 1126 1178 1142
rect 1050 1015 1067 1126
rect 1161 1015 1178 1126
rect 1050 996 1178 1015
rect 1260 1126 1388 1142
rect 1260 1015 1277 1126
rect 1371 1015 1388 1126
rect 1260 996 1388 1015
rect 1470 1126 1598 1142
rect 1470 1015 1487 1126
rect 1581 1015 1598 1126
rect 1470 996 1598 1015
rect 1680 1126 1808 1142
rect 1680 1015 1697 1126
rect 1791 1015 1808 1126
rect 1680 996 1808 1015
rect 1890 1126 2018 1142
rect 1890 1015 1907 1126
rect 2001 1015 2018 1126
rect 1890 996 2018 1015
rect 2100 1126 2228 1142
rect 2100 1015 2117 1126
rect 2211 1015 2228 1126
rect 2100 996 2228 1015
rect 2310 1126 2438 1142
rect 2310 1015 2327 1126
rect 2421 1015 2438 1126
rect 2310 996 2438 1015
rect 2520 1126 2648 1142
rect 2520 1015 2537 1126
rect 2631 1015 2648 1126
rect 2520 996 2648 1015
rect 2730 1126 2858 1142
rect 2730 1015 2747 1126
rect 2841 1015 2858 1126
rect 2730 996 2858 1015
rect 2940 1126 3068 1142
rect 2940 1015 2957 1126
rect 3051 1015 3068 1126
rect 2940 996 3068 1015
rect 3150 1126 3278 1142
rect 3150 1015 3167 1126
rect 3261 1015 3278 1126
rect 3150 996 3278 1015
rect 3360 1126 3488 1142
rect 3360 1015 3377 1126
rect 3471 1015 3488 1126
rect 3360 996 3488 1015
rect 3570 1126 3698 1142
rect 3570 1015 3587 1126
rect 3681 1015 3698 1126
rect 3570 996 3698 1015
rect 3780 1126 3908 1142
rect 3780 1015 3797 1126
rect 3891 1015 3908 1126
rect 3780 996 3908 1015
rect 3990 1126 4118 1142
rect 3990 1015 4007 1126
rect 4101 1015 4118 1126
rect 3990 996 4118 1015
rect 0 -79 128 -63
rect 0 -190 17 -79
rect 111 -190 128 -79
rect 0 -209 128 -190
rect 210 -79 338 -63
rect 210 -190 227 -79
rect 321 -190 338 -79
rect 210 -209 338 -190
rect 420 -79 548 -63
rect 420 -190 437 -79
rect 531 -190 548 -79
rect 420 -209 548 -190
rect 630 -79 758 -63
rect 630 -190 647 -79
rect 741 -190 758 -79
rect 630 -209 758 -190
rect 840 -79 968 -63
rect 840 -190 857 -79
rect 951 -190 968 -79
rect 840 -209 968 -190
rect 1050 -79 1178 -63
rect 1050 -190 1067 -79
rect 1161 -190 1178 -79
rect 1050 -209 1178 -190
rect 1260 -79 1388 -63
rect 1260 -190 1277 -79
rect 1371 -190 1388 -79
rect 1260 -209 1388 -190
rect 1470 -79 1598 -63
rect 1470 -190 1487 -79
rect 1581 -190 1598 -79
rect 1470 -209 1598 -190
rect 1680 -79 1808 -63
rect 1680 -190 1697 -79
rect 1791 -190 1808 -79
rect 1680 -209 1808 -190
rect 1890 -79 2018 -63
rect 1890 -190 1907 -79
rect 2001 -190 2018 -79
rect 1890 -209 2018 -190
rect 2100 -79 2228 -63
rect 2100 -190 2117 -79
rect 2211 -190 2228 -79
rect 2100 -209 2228 -190
rect 2310 -79 2438 -63
rect 2310 -190 2327 -79
rect 2421 -190 2438 -79
rect 2310 -209 2438 -190
rect 2520 -79 2648 -63
rect 2520 -190 2537 -79
rect 2631 -190 2648 -79
rect 2520 -209 2648 -190
rect 2730 -79 2858 -63
rect 2730 -190 2747 -79
rect 2841 -190 2858 -79
rect 2730 -209 2858 -190
rect 2940 -79 3068 -63
rect 2940 -190 2957 -79
rect 3051 -190 3068 -79
rect 2940 -209 3068 -190
rect 3150 -79 3278 -63
rect 3150 -190 3167 -79
rect 3261 -190 3278 -79
rect 3150 -209 3278 -190
rect 3360 -79 3488 -63
rect 3360 -190 3377 -79
rect 3471 -190 3488 -79
rect 3360 -209 3488 -190
rect 3570 -79 3698 -63
rect 3570 -190 3587 -79
rect 3681 -190 3698 -79
rect 3570 -209 3698 -190
rect 3780 -79 3908 -63
rect 3780 -190 3797 -79
rect 3891 -190 3908 -79
rect 3780 -209 3908 -190
rect 3990 -79 4118 -63
rect 3990 -190 4007 -79
rect 4101 -190 4118 -79
rect 3990 -209 4118 -190
<< psubdiffcont >>
rect 17 2230 111 2341
rect 227 2230 321 2341
rect 437 2230 531 2341
rect 647 2230 741 2341
rect 857 2230 951 2341
rect 1067 2230 1161 2341
rect 1277 2230 1371 2341
rect 1487 2230 1581 2341
rect 1697 2230 1791 2341
rect 1907 2230 2001 2341
rect 2117 2230 2211 2341
rect 2327 2230 2421 2341
rect 2537 2230 2631 2341
rect 2747 2230 2841 2341
rect 2957 2230 3051 2341
rect 3167 2230 3261 2341
rect 3377 2230 3471 2341
rect 3587 2230 3681 2341
rect 3797 2230 3891 2341
rect 4007 2230 4101 2341
rect 17 1015 111 1126
rect 227 1015 321 1126
rect 437 1015 531 1126
rect 647 1015 741 1126
rect 857 1015 951 1126
rect 1067 1015 1161 1126
rect 1277 1015 1371 1126
rect 1487 1015 1581 1126
rect 1697 1015 1791 1126
rect 1907 1015 2001 1126
rect 2117 1015 2211 1126
rect 2327 1015 2421 1126
rect 2537 1015 2631 1126
rect 2747 1015 2841 1126
rect 2957 1015 3051 1126
rect 3167 1015 3261 1126
rect 3377 1015 3471 1126
rect 3587 1015 3681 1126
rect 3797 1015 3891 1126
rect 4007 1015 4101 1126
rect 17 -190 111 -79
rect 227 -190 321 -79
rect 437 -190 531 -79
rect 647 -190 741 -79
rect 857 -190 951 -79
rect 1067 -190 1161 -79
rect 1277 -190 1371 -79
rect 1487 -190 1581 -79
rect 1697 -190 1791 -79
rect 1907 -190 2001 -79
rect 2117 -190 2211 -79
rect 2327 -190 2421 -79
rect 2537 -190 2631 -79
rect 2747 -190 2841 -79
rect 2957 -190 3051 -79
rect 3167 -190 3261 -79
rect 3377 -190 3471 -79
rect 3587 -190 3681 -79
rect 3797 -190 3891 -79
rect 4007 -190 4101 -79
<< polysilicon >>
rect 112 2130 4088 2144
rect 112 2108 1758 2130
rect 112 2002 212 2108
rect 316 2002 416 2046
rect 520 2002 620 2046
rect 724 2002 824 2108
rect 928 2002 1028 2108
rect 1132 2002 1232 2046
rect 1336 2002 1436 2046
rect 1540 2002 1640 2108
rect 1744 2058 1758 2108
rect 1830 2128 4088 2130
rect 1830 2108 2370 2128
rect 1830 2058 1844 2108
rect 1744 2002 1844 2058
rect 2356 2056 2370 2108
rect 2442 2108 4088 2128
rect 2442 2056 2456 2108
rect 1948 2002 2048 2046
rect 2152 2002 2252 2046
rect 2356 2002 2456 2056
rect 2560 2002 2660 2108
rect 2764 2002 2864 2046
rect 2968 2002 3068 2046
rect 3172 2002 3272 2108
rect 3376 2002 3476 2108
rect 3580 2002 3680 2046
rect 3784 2002 3884 2046
rect 3988 2002 4088 2108
rect 112 1758 212 1802
rect 316 1693 416 1802
rect 520 1693 620 1802
rect 724 1758 824 1802
rect 928 1758 1028 1802
rect 1132 1693 1232 1802
rect 1336 1693 1436 1802
rect 1540 1758 1640 1802
rect 1744 1758 1844 1802
rect 1948 1693 2048 1802
rect 2152 1693 2252 1802
rect 2356 1758 2456 1802
rect 2560 1758 2660 1802
rect 2764 1693 2864 1802
rect 2968 1693 3068 1802
rect 3172 1758 3272 1802
rect 3376 1758 3476 1802
rect 3580 1693 3680 1802
rect 3784 1693 3884 1802
rect 3988 1758 4088 1802
rect -151 1657 4354 1693
rect -151 1579 -115 1657
rect -181 1564 -92 1579
rect -181 1513 -165 1564
rect -111 1513 -92 1564
rect 112 1551 212 1657
rect 316 1551 416 1595
rect 520 1551 620 1595
rect 724 1551 824 1657
rect 928 1551 1028 1657
rect 1132 1551 1232 1595
rect 1336 1551 1436 1595
rect 1540 1551 1640 1657
rect 1744 1551 1844 1657
rect 1948 1551 2048 1595
rect 2152 1551 2252 1595
rect 2356 1551 2456 1657
rect 2560 1551 2660 1657
rect 2764 1551 2864 1595
rect 2968 1551 3068 1595
rect 3172 1551 3272 1657
rect 3376 1551 3476 1657
rect 3580 1551 3680 1595
rect 3784 1551 3884 1595
rect 3988 1551 4088 1657
rect 4318 1598 4354 1657
rect 4296 1582 4385 1598
rect -181 1498 -92 1513
rect 4296 1528 4312 1582
rect 4368 1528 4385 1582
rect 4296 1515 4385 1528
rect 112 1307 212 1351
rect 316 1248 416 1351
rect 520 1248 620 1351
rect 724 1307 824 1351
rect 928 1307 1028 1351
rect 1132 1248 1232 1351
rect 1336 1298 1436 1351
rect 1540 1307 1640 1351
rect 1744 1307 1844 1351
rect 1336 1248 1350 1298
rect 316 1226 1350 1248
rect 1422 1248 1436 1298
rect 1948 1248 2048 1351
rect 2152 1298 2252 1351
rect 2356 1307 2456 1351
rect 2560 1307 2660 1351
rect 2152 1248 2166 1298
rect 1422 1226 2166 1248
rect 2238 1248 2252 1298
rect 2764 1298 2864 1351
rect 2764 1248 2778 1298
rect 2238 1226 2778 1248
rect 2850 1248 2864 1298
rect 2968 1248 3068 1351
rect 3172 1307 3272 1351
rect 3376 1307 3476 1351
rect 3580 1248 3680 1351
rect 3784 1248 3884 1351
rect 3988 1307 4088 1351
rect 2850 1226 3884 1248
rect 316 1212 3884 1226
rect 112 915 4088 929
rect 112 843 126 915
rect 198 914 942 915
rect 198 893 738 914
rect 198 843 212 893
rect 112 787 212 843
rect 724 842 738 893
rect 810 893 942 914
rect 810 842 824 893
rect 316 787 416 831
rect 520 787 620 831
rect 724 787 824 842
rect 928 843 942 893
rect 1014 893 1554 915
rect 1014 843 1028 893
rect 928 787 1028 843
rect 1540 843 1554 893
rect 1626 893 1758 915
rect 1626 843 1640 893
rect 1132 787 1232 831
rect 1336 787 1436 831
rect 1540 787 1640 843
rect 1744 843 1758 893
rect 1830 893 2370 915
rect 1830 843 1844 893
rect 1744 787 1844 843
rect 2356 843 2370 893
rect 2442 893 2574 915
rect 2442 843 2456 893
rect 1948 787 2048 831
rect 2152 787 2252 831
rect 2356 787 2456 843
rect 2560 843 2574 893
rect 2646 893 3186 915
rect 2646 843 2660 893
rect 2560 787 2660 843
rect 3172 843 3186 893
rect 3258 893 3390 915
rect 3258 843 3272 893
rect 2764 787 2864 831
rect 2968 787 3068 831
rect 3172 787 3272 843
rect 3376 843 3390 893
rect 3462 893 4002 915
rect 3462 843 3476 893
rect 3376 787 3476 843
rect 3988 843 4002 893
rect 4074 843 4088 915
rect 3580 787 3680 831
rect 3784 787 3884 831
rect 3988 787 4088 843
rect 112 543 212 587
rect 316 531 416 587
rect 316 481 330 531
rect 112 459 330 481
rect 402 481 416 531
rect 520 531 620 587
rect 724 543 824 587
rect 928 543 1028 587
rect 520 481 534 531
rect 402 459 534 481
rect 606 481 620 531
rect 1132 531 1232 587
rect 1132 481 1146 531
rect 606 467 1146 481
rect 606 459 738 467
rect 112 445 738 459
rect 112 339 212 445
rect 724 395 738 445
rect 810 445 942 467
rect 810 395 824 445
rect 316 339 416 383
rect 520 339 620 383
rect 724 339 824 395
rect 928 395 942 445
rect 1014 459 1146 467
rect 1218 481 1232 531
rect 1336 531 1436 587
rect 1540 543 1640 587
rect 1744 543 1844 587
rect 1336 481 1350 531
rect 1218 459 1350 481
rect 1422 481 1436 531
rect 1948 531 2048 587
rect 1948 481 1962 531
rect 1422 467 1962 481
rect 1422 459 1554 467
rect 1014 445 1554 459
rect 1014 395 1028 445
rect 928 339 1028 395
rect 1540 395 1554 445
rect 1626 445 1758 467
rect 1626 395 1640 445
rect 1132 339 1232 383
rect 1336 339 1436 383
rect 1540 339 1640 395
rect 1744 395 1758 445
rect 1830 459 1962 467
rect 2034 481 2048 531
rect 2152 531 2252 587
rect 2356 543 2456 587
rect 2560 543 2660 587
rect 2152 481 2166 531
rect 2034 459 2166 481
rect 2238 481 2252 531
rect 2764 531 2864 587
rect 2764 481 2778 531
rect 2238 467 2778 481
rect 2238 459 2370 467
rect 1830 445 2370 459
rect 1830 395 1844 445
rect 1744 339 1844 395
rect 2356 395 2370 445
rect 2442 445 2574 467
rect 2442 395 2456 445
rect 1948 339 2048 383
rect 2152 339 2252 383
rect 2356 339 2456 395
rect 2560 395 2574 445
rect 2646 459 2778 467
rect 2850 481 2864 531
rect 2968 531 3068 587
rect 3172 543 3272 587
rect 3376 543 3476 587
rect 2968 481 2982 531
rect 2850 459 2982 481
rect 3054 481 3068 531
rect 3580 531 3680 587
rect 3580 481 3594 531
rect 3054 467 3594 481
rect 3054 459 3186 467
rect 2646 445 3186 459
rect 2646 395 2660 445
rect 2560 339 2660 395
rect 3172 395 3186 445
rect 3258 445 3390 467
rect 3258 395 3272 445
rect 2764 339 2864 383
rect 2968 339 3068 383
rect 3172 339 3272 395
rect 3376 395 3390 445
rect 3462 459 3594 467
rect 3666 481 3680 531
rect 3784 531 3884 587
rect 3988 543 4088 587
rect 3784 481 3798 531
rect 3666 459 3798 481
rect 3870 481 3884 531
rect 3870 459 4088 481
rect 3462 445 4088 459
rect 3462 395 3476 445
rect 3376 339 3476 395
rect 3580 339 3680 383
rect 3784 339 3884 383
rect 3988 339 4088 445
rect 112 95 212 139
rect 316 86 416 139
rect 316 14 330 86
rect 402 36 416 86
rect 520 86 620 139
rect 724 95 824 139
rect 928 95 1028 139
rect 520 36 534 86
rect 402 14 534 36
rect 606 36 620 86
rect 1132 86 1232 139
rect 1132 36 1146 86
rect 606 14 1146 36
rect 1218 36 1232 86
rect 1336 86 1436 139
rect 1540 95 1640 139
rect 1744 95 1844 139
rect 1336 36 1350 86
rect 1218 14 1350 36
rect 1422 36 1436 86
rect 1948 86 2048 139
rect 1948 36 1962 86
rect 1422 14 1962 36
rect 2034 36 2048 86
rect 2152 86 2252 139
rect 2356 95 2456 139
rect 2560 95 2660 139
rect 2152 36 2166 86
rect 2034 14 2166 36
rect 2238 36 2252 86
rect 2764 86 2864 139
rect 2764 36 2778 86
rect 2238 14 2778 36
rect 2850 36 2864 86
rect 2968 86 3068 139
rect 3172 95 3272 139
rect 3376 95 3476 139
rect 2968 36 2982 86
rect 2850 14 2982 36
rect 3054 36 3068 86
rect 3580 86 3680 139
rect 3580 36 3594 86
rect 3054 14 3594 36
rect 3666 36 3680 86
rect 3784 86 3884 139
rect 3988 95 4088 139
rect 3784 36 3798 86
rect 3666 14 3798 36
rect 3870 14 3884 86
rect 316 0 3884 14
<< polycontact >>
rect 1758 2058 1830 2130
rect 2370 2056 2442 2128
rect -165 1513 -111 1564
rect 4312 1528 4368 1582
rect 1350 1226 1422 1298
rect 2166 1226 2238 1298
rect 2778 1226 2850 1298
rect 126 843 198 915
rect 738 842 810 914
rect 942 843 1014 915
rect 1554 843 1626 915
rect 1758 843 1830 915
rect 2370 843 2442 915
rect 2574 843 2646 915
rect 3186 843 3258 915
rect 3390 843 3462 915
rect 4002 843 4074 915
rect 330 459 402 531
rect 534 459 606 531
rect 738 395 810 467
rect 942 395 1014 467
rect 1146 459 1218 531
rect 1350 459 1422 531
rect 1554 395 1626 467
rect 1758 395 1830 467
rect 1962 459 2034 531
rect 2166 459 2238 531
rect 2370 395 2442 467
rect 2574 395 2646 467
rect 2778 459 2850 531
rect 2982 459 3054 531
rect 3186 395 3258 467
rect 3390 395 3462 467
rect 3594 459 3666 531
rect 3798 459 3870 531
rect 330 14 402 86
rect 534 14 606 86
rect 1146 14 1218 86
rect 1350 14 1422 86
rect 1962 14 2034 86
rect 2166 14 2238 86
rect 2778 14 2850 86
rect 2982 14 3054 86
rect 3594 14 3666 86
rect 3798 14 3870 86
<< metal1 >>
rect -442 2840 -369 2850
rect -442 2782 -433 2840
rect -379 2782 -369 2840
rect -442 2771 -369 2782
rect 0 2341 4200 2357
rect 0 2230 17 2341
rect 111 2230 227 2341
rect 321 2230 437 2341
rect 531 2230 647 2341
rect 741 2230 857 2341
rect 951 2230 1067 2341
rect 1161 2230 1277 2341
rect 1371 2230 1487 2341
rect 1581 2230 1697 2341
rect 1791 2230 1907 2341
rect 2001 2230 2117 2341
rect 2211 2230 2327 2341
rect 2421 2230 2537 2341
rect 2631 2230 2747 2341
rect 2841 2230 2957 2341
rect 3051 2230 3167 2341
rect 3261 2230 3377 2341
rect 3471 2230 3587 2341
rect 3681 2230 3797 2341
rect 3891 2230 4007 2341
rect 4101 2230 4200 2341
rect 0 2211 4200 2230
rect 37 1989 83 2000
rect 241 1989 287 2000
rect 220 1926 241 1936
rect 445 1989 491 2211
rect 220 1868 229 1926
rect 220 1857 241 1868
rect 37 1718 83 1815
rect 287 1857 293 1936
rect 241 1804 287 1815
rect 649 1989 695 2000
rect 631 1934 649 1944
rect 853 1989 899 2000
rect 631 1876 640 1934
rect 631 1865 649 1876
rect 445 1804 491 1815
rect 695 1865 704 1944
rect 649 1804 695 1815
rect 1057 1989 1103 2000
rect 1038 1933 1057 1943
rect 1261 1989 1307 2211
rect 1749 2130 1839 2139
rect 1749 2058 1758 2130
rect 1830 2058 1839 2130
rect 1749 2049 1839 2058
rect 1038 1875 1047 1933
rect 1038 1864 1057 1875
rect 853 1718 899 1815
rect 1103 1864 1111 1943
rect 1057 1804 1103 1815
rect 1465 1989 1511 2000
rect 1448 1933 1465 1943
rect 1669 1989 1715 2000
rect 1448 1875 1457 1933
rect 1448 1864 1465 1875
rect 1261 1804 1307 1815
rect 1511 1864 1521 1943
rect 1465 1804 1511 1815
rect 1873 1989 1919 2000
rect 1854 1933 1873 1943
rect 2077 1989 2123 2211
rect 2361 2128 2451 2137
rect 2361 2056 2370 2128
rect 2442 2056 2451 2128
rect 2361 2047 2451 2056
rect 1854 1875 1863 1933
rect 1854 1864 1873 1875
rect 1669 1718 1715 1815
rect 1919 1864 1927 1943
rect 1873 1804 1919 1815
rect 2281 1989 2327 2000
rect 2264 1933 2281 1943
rect 2485 1989 2531 2000
rect 2264 1875 2273 1933
rect 2264 1864 2281 1875
rect 2077 1804 2123 1815
rect 2327 1864 2337 1943
rect 2281 1804 2327 1815
rect 2689 1989 2735 2000
rect 2671 1933 2689 1943
rect 2893 1989 2939 2211
rect 2671 1875 2680 1933
rect 2671 1864 2689 1875
rect 2485 1718 2531 1815
rect 2735 1864 2744 1943
rect 2689 1804 2735 1815
rect 3097 1989 3143 2000
rect 3076 1933 3097 1943
rect 3301 1989 3347 2000
rect 3076 1875 3085 1933
rect 3076 1864 3097 1875
rect 2893 1804 2939 1815
rect 3143 1864 3149 1943
rect 3097 1804 3143 1815
rect 3505 1989 3551 2000
rect 3486 1933 3505 1943
rect 3709 1989 3755 2211
rect 3486 1875 3495 1933
rect 3486 1864 3505 1875
rect 3301 1718 3347 1815
rect 3551 1864 3559 1943
rect 3505 1804 3551 1815
rect 3913 1989 3959 2000
rect 3897 1937 3913 1947
rect 4117 1989 4163 2000
rect 3959 1937 3970 1947
rect 3897 1879 3906 1937
rect 3960 1879 3970 1937
rect 3897 1868 3913 1879
rect 3709 1804 3755 1815
rect 3959 1868 3970 1879
rect 3913 1804 3959 1815
rect 4117 1718 4163 1815
rect 37 1653 4163 1718
rect -181 1564 -92 1579
rect -181 1513 -165 1564
rect -111 1513 -92 1564
rect -181 530 -92 1513
rect 37 1538 83 1549
rect 241 1538 287 1549
rect 224 1482 241 1492
rect 445 1538 491 1653
rect 224 1424 233 1482
rect 224 1413 241 1424
rect 37 1142 83 1364
rect 287 1413 297 1492
rect 241 1353 287 1364
rect 649 1538 695 1549
rect 634 1481 649 1491
rect 853 1538 899 1549
rect 695 1481 707 1491
rect 634 1423 643 1481
rect 697 1423 707 1481
rect 634 1412 649 1423
rect 445 1353 491 1364
rect 695 1412 707 1423
rect 649 1353 695 1364
rect 1057 1538 1103 1549
rect 1043 1480 1057 1490
rect 1261 1538 1307 1653
rect 1103 1480 1116 1490
rect 1043 1422 1052 1480
rect 1106 1422 1116 1480
rect 1043 1411 1057 1422
rect 853 1142 899 1364
rect 1103 1411 1116 1422
rect 1057 1353 1103 1364
rect 1465 1538 1511 1549
rect 1452 1479 1465 1489
rect 1669 1538 1715 1549
rect 1511 1479 1525 1489
rect 1452 1421 1461 1479
rect 1515 1421 1525 1479
rect 1452 1410 1465 1421
rect 1261 1353 1307 1364
rect 1511 1410 1525 1421
rect 1465 1353 1511 1364
rect 1873 1538 1919 1549
rect 1861 1479 1873 1489
rect 2077 1538 2123 1603
rect 1919 1479 1934 1489
rect 1861 1421 1870 1479
rect 1924 1421 1934 1479
rect 1861 1410 1873 1421
rect 1341 1298 1431 1307
rect 1341 1226 1350 1298
rect 1422 1226 1431 1298
rect 1341 1217 1431 1226
rect 1669 1142 1715 1364
rect 1919 1410 1934 1421
rect 1873 1353 1919 1364
rect 2281 1538 2327 1549
rect 2267 1479 2281 1489
rect 2485 1538 2531 1549
rect 2327 1479 2340 1489
rect 2267 1421 2276 1479
rect 2330 1421 2340 1479
rect 2267 1410 2281 1421
rect 2077 1353 2123 1364
rect 2327 1410 2340 1421
rect 2281 1353 2327 1364
rect 2689 1538 2735 1549
rect 2674 1479 2689 1489
rect 2893 1538 2939 1653
rect 2735 1479 2747 1489
rect 2674 1421 2683 1479
rect 2737 1421 2747 1479
rect 2674 1410 2689 1421
rect 2157 1298 2247 1307
rect 2157 1226 2166 1298
rect 2238 1226 2247 1298
rect 2157 1217 2247 1226
rect 2485 1142 2531 1364
rect 2735 1410 2747 1421
rect 2689 1353 2735 1364
rect 3097 1538 3143 1549
rect 3082 1478 3097 1488
rect 3301 1538 3347 1549
rect 3143 1478 3155 1488
rect 3082 1420 3091 1478
rect 3145 1420 3155 1478
rect 3082 1409 3097 1420
rect 2893 1353 2939 1364
rect 3143 1409 3155 1420
rect 3097 1353 3143 1364
rect 3505 1538 3551 1549
rect 3490 1480 3505 1490
rect 3709 1538 3755 1653
rect 4296 1582 4385 1598
rect 3551 1480 3563 1490
rect 3490 1422 3499 1480
rect 3553 1422 3563 1480
rect 3490 1411 3505 1422
rect 2769 1298 2859 1307
rect 2769 1226 2778 1298
rect 2850 1226 2859 1298
rect 2769 1217 2859 1226
rect 3301 1142 3347 1364
rect 3551 1411 3563 1422
rect 3505 1353 3551 1364
rect 3913 1538 3959 1549
rect 3898 1479 3913 1489
rect 4117 1538 4163 1549
rect 3959 1479 3971 1489
rect 3898 1421 3907 1479
rect 3961 1421 3971 1479
rect 3898 1410 3913 1421
rect 3709 1353 3755 1364
rect 3959 1410 3971 1421
rect 3913 1353 3959 1364
rect 4117 1142 4163 1364
rect 4296 1528 4312 1582
rect 4368 1528 4385 1582
rect 0 1126 4200 1142
rect 0 1015 17 1126
rect 111 1015 227 1126
rect 321 1015 437 1126
rect 531 1015 647 1126
rect 741 1015 857 1126
rect 951 1015 1067 1126
rect 1161 1015 1277 1126
rect 1371 1015 1487 1126
rect 1581 1015 1697 1126
rect 1791 1015 1907 1126
rect 2001 1015 2117 1126
rect 2211 1015 2327 1126
rect 2421 1015 2537 1126
rect 2631 1015 2747 1126
rect 2841 1015 2957 1126
rect 3051 1015 3167 1126
rect 3261 1015 3377 1126
rect 3471 1015 3587 1126
rect 3681 1015 3797 1126
rect 3891 1015 4007 1126
rect 4101 1015 4200 1126
rect 0 996 4200 1015
rect 117 915 207 924
rect 117 880 126 915
rect 37 843 126 880
rect 198 843 207 915
rect 37 834 207 843
rect 37 774 83 834
rect 37 589 83 600
rect 241 774 287 785
rect 241 548 287 600
rect 445 774 491 996
rect 729 914 819 923
rect 729 842 738 914
rect 810 880 819 914
rect 933 915 1023 924
rect 933 880 942 915
rect 810 843 942 880
rect 1014 843 1023 915
rect 810 842 1023 843
rect 729 834 1023 842
rect 729 833 933 834
rect 445 589 491 600
rect 649 774 695 785
rect 241 540 359 548
rect 649 547 695 600
rect 853 774 899 833
rect 853 589 899 600
rect 1057 774 1103 785
rect 601 540 695 547
rect 241 531 411 540
rect 241 530 330 531
rect -181 459 330 530
rect 402 530 411 531
rect 525 531 695 540
rect 525 530 534 531
rect 402 459 534 530
rect 606 530 695 531
rect 1057 543 1103 600
rect 1261 774 1307 996
rect 1545 915 1635 924
rect 1545 843 1554 915
rect 1626 881 1635 915
rect 1749 915 1839 924
rect 1749 881 1758 915
rect 1626 843 1758 881
rect 1830 843 1839 915
rect 1545 834 1839 843
rect 1261 589 1307 600
rect 1465 774 1511 785
rect 1465 554 1511 600
rect 1669 774 1715 834
rect 1669 589 1715 600
rect 1873 774 1919 785
rect 1057 540 1169 543
rect 1405 540 1511 554
rect 1057 531 1227 540
rect 1057 530 1146 531
rect 606 467 1146 530
rect 606 459 738 467
rect -181 441 738 459
rect 241 430 358 441
rect 37 326 83 337
rect 37 -63 83 152
rect 241 326 287 430
rect 649 395 738 441
rect 810 441 942 467
rect 810 395 819 441
rect 649 386 819 395
rect 933 395 942 441
rect 1014 459 1146 467
rect 1218 530 1227 531
rect 1341 531 1511 540
rect 1341 530 1350 531
rect 1218 459 1350 530
rect 1422 530 1511 531
rect 1873 543 1919 600
rect 2077 774 2123 996
rect 2361 915 2451 924
rect 2361 843 2370 915
rect 2442 881 2451 915
rect 2565 915 2655 924
rect 2565 881 2574 915
rect 2442 843 2574 881
rect 2646 843 2655 915
rect 2361 834 2655 843
rect 2077 589 2123 600
rect 2281 774 2327 785
rect 2281 560 2327 600
rect 2485 774 2531 834
rect 2485 589 2531 600
rect 2689 774 2735 785
rect 1873 540 1974 543
rect 2224 540 2327 560
rect 1873 531 2043 540
rect 1873 530 1962 531
rect 1422 467 1962 530
rect 1422 459 1554 467
rect 1014 441 1554 459
rect 1014 395 1103 441
rect 933 386 1103 395
rect 241 141 287 152
rect 445 326 491 337
rect 445 95 491 152
rect 649 326 695 386
rect 987 379 1103 386
rect 649 141 695 152
rect 853 326 899 337
rect 321 86 615 95
rect 321 14 330 86
rect 402 48 534 86
rect 402 14 411 48
rect 321 5 411 14
rect 525 14 534 48
rect 606 14 615 86
rect 525 5 615 14
rect 853 -63 899 152
rect 1057 326 1103 379
rect 1465 395 1554 441
rect 1626 441 1758 467
rect 1626 395 1635 441
rect 1465 386 1635 395
rect 1749 395 1758 441
rect 1830 459 1962 467
rect 2034 530 2043 531
rect 2157 531 2327 540
rect 2157 530 2166 531
rect 2034 459 2166 530
rect 2238 530 2327 531
rect 2689 556 2735 600
rect 2893 774 2939 996
rect 3177 915 3267 924
rect 3177 843 3186 915
rect 3258 881 3267 915
rect 3381 915 3471 924
rect 3381 881 3390 915
rect 3258 843 3390 881
rect 3462 843 3471 915
rect 3177 834 3471 843
rect 2893 589 2939 600
rect 3097 774 3143 785
rect 3097 564 3143 600
rect 3301 774 3347 834
rect 3301 589 3347 600
rect 3505 774 3551 785
rect 2689 540 2785 556
rect 3031 540 3143 564
rect 2689 531 2859 540
rect 2689 530 2778 531
rect 2238 467 2778 530
rect 2238 459 2370 467
rect 1830 441 2370 459
rect 1830 395 1919 441
rect 1749 386 1919 395
rect 1465 383 1610 386
rect 1057 141 1103 152
rect 1261 326 1307 337
rect 1261 95 1307 152
rect 1465 326 1511 383
rect 1781 377 1919 386
rect 1465 141 1511 152
rect 1669 326 1715 337
rect 1137 86 1431 95
rect 1137 14 1146 86
rect 1218 48 1350 86
rect 1218 14 1227 48
rect 1137 5 1227 14
rect 1341 14 1350 48
rect 1422 14 1431 86
rect 1341 5 1431 14
rect 1669 -63 1715 152
rect 1873 326 1919 377
rect 2281 395 2370 441
rect 2442 441 2574 467
rect 2442 395 2451 441
rect 2281 386 2451 395
rect 2565 395 2574 441
rect 2646 459 2778 467
rect 2850 530 2859 531
rect 2973 531 3143 540
rect 2973 530 2982 531
rect 2850 459 2982 530
rect 3054 530 3143 531
rect 3505 567 3551 600
rect 3709 774 3755 996
rect 3993 915 4083 924
rect 3993 843 4002 915
rect 4074 880 4083 915
rect 4074 843 4163 880
rect 3993 834 4163 843
rect 3709 589 3755 600
rect 3913 774 3959 785
rect 3505 540 3625 567
rect 3913 566 3959 600
rect 4117 774 4163 834
rect 4117 589 4163 600
rect 3858 540 3959 566
rect 3505 531 3675 540
rect 3505 530 3594 531
rect 3054 467 3594 530
rect 3054 459 3186 467
rect 2646 441 3186 459
rect 2646 395 2735 441
rect 2565 386 2735 395
rect 2281 367 2389 386
rect 2622 372 2735 386
rect 1873 141 1919 152
rect 2077 326 2123 337
rect 2077 95 2123 152
rect 2281 326 2327 367
rect 2281 141 2327 152
rect 2485 326 2531 337
rect 1953 86 2247 95
rect 1953 14 1962 86
rect 2034 48 2166 86
rect 2034 14 2043 48
rect 1953 5 2043 14
rect 2157 14 2166 48
rect 2238 14 2247 86
rect 2157 5 2247 14
rect 2485 -63 2531 152
rect 2689 326 2735 372
rect 3097 395 3186 441
rect 3258 441 3390 467
rect 3258 395 3267 441
rect 3097 386 3267 395
rect 3381 395 3390 441
rect 3462 459 3594 467
rect 3666 530 3675 531
rect 3789 531 3959 540
rect 3789 530 3798 531
rect 3666 459 3798 530
rect 3870 530 3959 531
rect 4296 530 4385 1528
rect 3870 459 4385 530
rect 3462 441 4385 459
rect 3462 395 3551 441
rect 3381 386 3551 395
rect 3097 378 3229 386
rect 2689 141 2735 152
rect 2893 326 2939 337
rect 2893 95 2939 152
rect 3097 326 3143 378
rect 3439 368 3551 386
rect 3097 141 3143 152
rect 3301 326 3347 337
rect 2769 86 3063 95
rect 2769 14 2778 86
rect 2850 48 2982 86
rect 2850 14 2859 48
rect 2769 5 2859 14
rect 2973 14 2982 48
rect 3054 14 3063 86
rect 2973 5 3063 14
rect 3301 -63 3347 152
rect 3505 326 3551 368
rect 3505 141 3551 152
rect 3709 326 3755 337
rect 3709 95 3755 152
rect 3913 326 3959 441
rect 3913 141 3959 152
rect 4117 326 4163 337
rect 3585 86 3879 95
rect 3585 14 3594 86
rect 3666 48 3798 86
rect 3666 14 3675 48
rect 3585 5 3675 14
rect 3789 14 3798 48
rect 3870 14 3879 86
rect 3789 5 3879 14
rect 4117 -63 4163 152
rect 0 -79 4200 -63
rect 0 -190 17 -79
rect 111 -190 227 -79
rect 321 -190 437 -79
rect 531 -190 647 -79
rect 741 -190 857 -79
rect 951 -190 1067 -79
rect 1161 -190 1277 -79
rect 1371 -190 1487 -79
rect 1581 -190 1697 -79
rect 1791 -190 1907 -79
rect 2001 -190 2117 -79
rect 2211 -190 2327 -79
rect 2421 -190 2537 -79
rect 2631 -190 2747 -79
rect 2841 -190 2957 -79
rect 3051 -190 3167 -79
rect 3261 -190 3377 -79
rect 3471 -190 3587 -79
rect 3681 -190 3797 -79
rect 3891 -190 4007 -79
rect 4101 -190 4200 -79
rect 0 -209 4200 -190
<< via1 >>
rect -433 2782 -379 2840
rect 34 2268 89 2321
rect 4022 2256 4077 2309
rect 229 1868 241 1926
rect 241 1868 283 1926
rect 640 1876 649 1934
rect 649 1876 694 1934
rect 1764 2064 1819 2120
rect 1047 1875 1057 1933
rect 1057 1875 1101 1933
rect 1457 1875 1465 1933
rect 1465 1875 1511 1933
rect 2379 2065 2434 2121
rect 1863 1875 1873 1933
rect 1873 1875 1917 1933
rect 2273 1875 2281 1933
rect 2281 1875 2327 1933
rect 2680 1875 2689 1933
rect 2689 1875 2734 1933
rect 3085 1875 3097 1933
rect 3097 1875 3139 1933
rect 3495 1875 3505 1933
rect 3505 1875 3549 1933
rect 3906 1879 3913 1937
rect 3913 1879 3959 1937
rect 3959 1879 3960 1937
rect 233 1424 241 1482
rect 241 1424 287 1482
rect 643 1423 649 1481
rect 649 1423 695 1481
rect 695 1423 697 1481
rect 1052 1422 1057 1480
rect 1057 1422 1103 1480
rect 1103 1422 1106 1480
rect 1461 1421 1465 1479
rect 1465 1421 1511 1479
rect 1511 1421 1515 1479
rect 1870 1421 1873 1479
rect 1873 1421 1919 1479
rect 1919 1421 1924 1479
rect 1357 1234 1414 1289
rect 2276 1421 2281 1479
rect 2281 1421 2327 1479
rect 2327 1421 2330 1479
rect 2683 1421 2689 1479
rect 2689 1421 2735 1479
rect 2735 1421 2737 1479
rect 2173 1235 2230 1290
rect 3091 1420 3097 1478
rect 3097 1420 3143 1478
rect 3143 1420 3145 1478
rect 3499 1422 3505 1480
rect 3505 1422 3551 1480
rect 3551 1422 3553 1480
rect 2782 1231 2842 1291
rect 3907 1421 3913 1479
rect 3913 1421 3959 1479
rect 3959 1421 3961 1479
rect 34 1053 89 1106
rect 4022 1041 4077 1094
rect 1561 851 1616 906
rect 2380 854 2432 906
rect 1154 21 1207 77
rect 1974 21 2029 79
rect 2785 21 2842 80
rect 34 -162 89 -109
rect 4025 -165 4080 -112
<< metal2 >>
rect -442 2840 -369 2850
rect -442 2782 -433 2840
rect -379 2782 -369 2840
rect -442 2771 -369 2782
rect 24 2321 101 2332
rect 24 2268 34 2321
rect 89 2268 101 2321
rect 24 2256 101 2268
rect 4012 2309 4089 2320
rect 4012 2256 4022 2309
rect 4077 2256 4089 2309
rect 33 1117 89 2256
rect 4012 2244 4089 2256
rect 1749 2126 1839 2139
rect 1749 2063 1762 2126
rect 1826 2063 1839 2126
rect 1749 2049 1839 2063
rect 2361 2123 2451 2137
rect 2361 2061 2375 2123
rect 2437 2061 2451 2123
rect 2361 2047 2451 2061
rect 220 1926 293 1936
rect 220 1868 229 1926
rect 283 1919 293 1926
rect 631 1934 704 1944
rect 631 1919 640 1934
rect 283 1876 640 1919
rect 694 1919 704 1934
rect 1038 1933 1111 1943
rect 1038 1919 1047 1933
rect 694 1876 1047 1919
rect 283 1875 1047 1876
rect 1101 1919 1111 1933
rect 1448 1933 1521 1943
rect 1448 1919 1457 1933
rect 1101 1875 1457 1919
rect 1511 1919 1521 1933
rect 1854 1933 1927 1943
rect 1854 1919 1863 1933
rect 1511 1875 1863 1919
rect 1917 1919 1927 1933
rect 2264 1933 2337 1943
rect 2264 1919 2273 1933
rect 1917 1875 2273 1919
rect 2327 1919 2337 1933
rect 2671 1933 2744 1943
rect 2671 1919 2680 1933
rect 2327 1875 2680 1919
rect 2734 1919 2744 1933
rect 3076 1933 3149 1943
rect 3076 1919 3085 1933
rect 2734 1875 3085 1919
rect 3139 1919 3149 1933
rect 3486 1933 3559 1943
rect 3486 1919 3495 1933
rect 3139 1875 3495 1919
rect 3549 1919 3559 1933
rect 3897 1937 3970 1947
rect 3897 1919 3906 1937
rect 3549 1879 3906 1919
rect 3960 1879 3970 1937
rect 3549 1875 3970 1879
rect 283 1868 3970 1875
rect 220 1863 3966 1868
rect 220 1857 293 1863
rect 229 1492 285 1857
rect 224 1482 297 1492
rect 638 1491 694 1863
rect 224 1424 233 1482
rect 287 1424 297 1482
rect 224 1413 297 1424
rect 634 1481 707 1491
rect 1047 1490 1103 1863
rect 634 1423 643 1481
rect 697 1423 707 1481
rect 634 1412 707 1423
rect 1043 1480 1116 1490
rect 1458 1489 1514 1863
rect 1865 1489 1921 1863
rect 2280 1489 2336 1863
rect 2677 1489 2733 1863
rect 1043 1422 1052 1480
rect 1106 1422 1116 1480
rect 1043 1411 1116 1422
rect 1452 1479 1525 1489
rect 1452 1421 1461 1479
rect 1515 1421 1525 1479
rect 1452 1410 1525 1421
rect 1861 1479 1934 1489
rect 1861 1421 1870 1479
rect 1924 1421 1934 1479
rect 1861 1410 1934 1421
rect 2267 1479 2340 1489
rect 2267 1421 2276 1479
rect 2330 1421 2340 1479
rect 2267 1410 2340 1421
rect 2674 1479 2747 1489
rect 3088 1488 3144 1863
rect 3504 1490 3560 1863
rect 2674 1421 2683 1479
rect 2737 1421 2747 1479
rect 2674 1410 2747 1421
rect 3082 1478 3155 1488
rect 3082 1420 3091 1478
rect 3145 1420 3155 1478
rect 3082 1409 3155 1420
rect 3490 1480 3563 1490
rect 3910 1489 3966 1863
rect 3490 1422 3499 1480
rect 3553 1422 3563 1480
rect 3490 1411 3563 1422
rect 3898 1479 3971 1489
rect 3898 1421 3907 1479
rect 3961 1421 3971 1479
rect 3898 1410 3971 1421
rect 1341 1293 1431 1307
rect 1341 1230 1353 1293
rect 1417 1290 1431 1293
rect 2157 1293 2246 1307
rect 2157 1290 2171 1293
rect 2232 1290 2246 1293
rect 2769 1292 2859 1307
rect 2769 1290 2782 1292
rect 1417 1234 2171 1290
rect 1417 1230 1431 1234
rect 1341 1217 1431 1230
rect 2157 1231 2171 1234
rect 2232 1234 2782 1290
rect 2232 1231 2263 1234
rect 2157 1217 2263 1231
rect 2769 1230 2782 1234
rect 2843 1230 2859 1292
rect 2769 1217 2859 1230
rect 24 1106 101 1117
rect 24 1053 34 1106
rect 89 1053 101 1106
rect 24 1041 101 1053
rect 33 -98 89 1041
rect 1367 904 1423 1217
rect 1548 906 1630 921
rect 1548 904 1561 906
rect 1367 851 1561 904
rect 1616 904 1630 906
rect 2207 904 2263 1217
rect 2366 906 2447 920
rect 2366 904 2380 906
rect 1616 854 2380 904
rect 2432 904 2447 906
rect 2799 904 2855 1217
rect 4029 1105 4085 2244
rect 4012 1094 4089 1105
rect 4012 1041 4022 1094
rect 4077 1041 4089 1094
rect 4012 1029 4089 1041
rect 2432 854 2855 904
rect 1616 851 2855 854
rect 1367 848 2855 851
rect 1548 837 1630 848
rect 2363 840 2447 848
rect 1139 77 1222 91
rect 1139 21 1154 77
rect 1207 75 1222 77
rect 1554 75 1610 837
rect 1961 79 2044 91
rect 1961 75 1974 79
rect 1207 21 1974 75
rect 2029 75 2044 79
rect 2363 75 2419 840
rect 2772 80 2855 92
rect 2772 75 2785 80
rect 2029 21 2785 75
rect 2842 21 2855 80
rect 1139 19 2855 21
rect 1139 8 1222 19
rect 1961 8 2044 19
rect 2772 8 2855 19
rect 24 -109 101 -98
rect 4029 -101 4085 1029
rect 24 -162 34 -109
rect 89 -162 101 -109
rect 24 -174 101 -162
rect 4015 -112 4092 -101
rect 4015 -165 4025 -112
rect 4080 -165 4092 -112
rect 4015 -177 4092 -165
<< via2 >>
rect 1762 2120 1826 2126
rect 1762 2064 1764 2120
rect 1764 2064 1819 2120
rect 1819 2064 1826 2120
rect 1762 2063 1826 2064
rect 2375 2121 2437 2123
rect 2375 2065 2379 2121
rect 2379 2065 2434 2121
rect 2434 2065 2437 2121
rect 2375 2061 2437 2065
rect 1353 1289 1417 1293
rect 2171 1290 2232 1293
rect 2782 1291 2843 1292
rect 1353 1234 1357 1289
rect 1357 1234 1414 1289
rect 1414 1234 1417 1289
rect 2171 1235 2173 1290
rect 2173 1235 2230 1290
rect 2230 1235 2232 1290
rect 1353 1230 1417 1234
rect 2171 1231 2232 1235
rect 2782 1231 2842 1291
rect 2842 1231 2843 1291
rect 2782 1230 2843 1231
<< metal3 >>
rect 1749 2128 1839 2139
rect 2361 2128 2451 2137
rect 1749 2126 2451 2128
rect 1749 2063 1762 2126
rect 1826 2123 2451 2126
rect 1826 2067 2375 2123
rect 1826 2063 1839 2067
rect 1749 2049 1839 2063
rect 2361 2061 2375 2067
rect 2437 2061 2451 2123
rect 1341 1293 1431 1307
rect 1341 1230 1353 1293
rect 1417 1291 1431 1293
rect 1417 1290 1478 1291
rect 1769 1290 1830 2049
rect 2361 2047 2451 2061
rect 2157 1293 2247 1307
rect 2157 1290 2171 1293
rect 1417 1231 2171 1290
rect 2232 1290 2247 1293
rect 2375 1290 2436 2047
rect 2769 1292 2859 1307
rect 2769 1290 2782 1292
rect 2232 1231 2782 1290
rect 1417 1230 2782 1231
rect 2843 1230 2859 1292
rect 1341 1229 2859 1230
rect 1341 1217 1431 1229
rect 2157 1217 2247 1229
rect 2769 1217 2859 1229
<< end >>
