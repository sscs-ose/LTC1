magic
tech gf180mcuC
magscale 1 10
timestamp 1694501647
<< nwell >>
rect -304 -386 304 386
<< nsubdiff >>
rect -280 290 280 362
rect -280 -290 -208 290
rect 208 -290 280 290
rect -280 -362 280 -290
<< polysilicon >>
rect -120 189 120 202
rect -120 143 -107 189
rect 107 143 120 189
rect -120 100 120 143
rect -120 -143 120 -100
rect -120 -189 -107 -143
rect 107 -189 120 -143
rect -120 -202 120 -189
<< polycontact >>
rect -107 143 107 189
rect -107 -189 107 -143
<< ppolyres >>
rect -120 -100 120 100
<< metal1 >>
rect -118 143 -107 189
rect 107 143 118 189
rect -118 -189 -107 -143
rect 107 -189 118 -143
<< properties >>
string FIXED_BBOX -244 -326 244 326
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.2 l 1.0 m 1 nx 1 wmin 0.80 lmin 1.00 rho 315 val 278.761 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
