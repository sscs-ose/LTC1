magic
tech gf180mcuC
magscale 1 10
timestamp 1693141036
<< nwell >>
rect 21 513 1081 648
rect 21 507 166 513
rect 168 507 525 508
rect 528 507 1081 513
rect 371 470 907 483
rect 321 180 324 242
<< psubdiff >>
rect 38 -385 1061 -372
rect 38 -431 51 -385
rect 97 -431 145 -385
rect 191 -431 239 -385
rect 285 -431 333 -385
rect 379 -431 427 -385
rect 473 -431 521 -385
rect 567 -431 615 -385
rect 661 -431 709 -385
rect 755 -431 803 -385
rect 849 -431 897 -385
rect 943 -431 991 -385
rect 1037 -431 1061 -385
rect 38 -444 1061 -431
<< nsubdiff >>
rect 47 604 1002 617
rect 47 558 60 604
rect 106 558 154 604
rect 200 558 251 604
rect 297 558 345 604
rect 391 558 442 604
rect 488 558 536 604
rect 582 558 633 604
rect 679 558 727 604
rect 773 558 824 604
rect 870 558 918 604
rect 964 558 1002 604
rect 47 545 1002 558
<< psubdiffcont >>
rect 51 -431 97 -385
rect 145 -431 191 -385
rect 239 -431 285 -385
rect 333 -431 379 -385
rect 427 -431 473 -385
rect 521 -431 567 -385
rect 615 -431 661 -385
rect 709 -431 755 -385
rect 803 -431 849 -385
rect 897 -431 943 -385
rect 991 -431 1037 -385
<< nsubdiffcont >>
rect 60 558 106 604
rect 154 558 200 604
rect 251 558 297 604
rect 345 558 391 604
rect 442 558 488 604
rect 536 558 582 604
rect 633 558 679 604
rect 727 558 773 604
rect 824 558 870 604
rect 918 558 964 604
<< polysilicon >>
rect 195 417 907 483
rect 195 180 907 242
rect 194 -39 295 9
rect 194 -87 207 -39
rect 255 -83 295 -39
rect 399 -83 499 3
rect 603 -83 703 3
rect 807 -83 907 3
rect 255 -87 907 -83
rect 194 -131 907 -87
<< polycontact >>
rect 207 -87 255 -39
<< metal1 >>
rect 21 604 1081 648
rect 21 558 60 604
rect 106 558 154 604
rect 200 558 251 604
rect 297 558 345 604
rect 391 558 442 604
rect 488 558 536 604
rect 582 558 633 604
rect 679 558 727 604
rect 773 558 824 604
rect 870 558 918 604
rect 964 558 1081 604
rect 21 525 1081 558
rect 21 524 574 525
rect 40 381 106 524
rect 40 295 166 381
rect 120 135 166 295
rect 324 141 370 381
rect 528 372 574 524
rect 936 372 982 525
rect 528 140 574 302
rect 732 142 778 290
rect 936 134 982 298
rect 324 2 370 53
rect 732 2 778 50
rect 35 -39 266 -27
rect 35 -87 207 -39
rect 255 -87 266 -39
rect 35 -99 266 -87
rect 324 -44 1071 2
rect 324 -189 370 -44
rect 732 -182 778 -44
rect 120 -342 166 -256
rect 528 -342 574 -253
rect 936 -342 982 -252
rect 22 -385 1080 -342
rect 22 -431 51 -385
rect 97 -431 145 -385
rect 191 -431 239 -385
rect 285 -431 333 -385
rect 379 -431 427 -385
rect 473 -431 521 -385
rect 567 -431 615 -385
rect 661 -431 709 -385
rect 755 -431 803 -385
rect 849 -431 897 -385
rect 943 -431 991 -385
rect 1037 -431 1080 -385
rect 22 -485 1080 -431
use nmos_3p3_6FEA4B  nmos_3p3_6FEA4B_0
timestamp 1692505534
transform 1 0 551 0 1 -225
box -468 -118 468 118
use pmos_3p3_KYEELV  pmos_3p3_KYEELV_0
timestamp 1692985371
transform 1 0 551 0 1 215
box -530 -298 530 298
<< labels >>
flabel nsubdiffcont 559 581 559 581 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel psubdiffcont 544 -408 544 -408 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal1 53 -64 53 -64 0 FreeSans 800 0 0 0 IN
port 2 nsew
flabel metal1 1042 -23 1042 -23 0 FreeSans 800 0 0 0 OUT
port 3 nsew
<< end >>
