magic
tech gf180mcuC
magscale 1 10
timestamp 1695104611
<< nwell >>
rect -260 -1592 3252 1626
<< nsubdiff >>
rect -210 1559 3202 1576
rect -210 1513 -193 1559
rect -147 1513 -95 1559
rect -49 1513 3 1559
rect 49 1513 101 1559
rect 147 1513 199 1559
rect 245 1513 297 1559
rect 343 1513 395 1559
rect 441 1513 493 1559
rect 539 1513 591 1559
rect 637 1513 689 1559
rect 735 1513 787 1559
rect 833 1513 885 1559
rect 931 1513 983 1559
rect 1029 1513 1081 1559
rect 1127 1513 1179 1559
rect 1225 1513 1277 1559
rect 1323 1513 1375 1559
rect 1421 1513 1473 1559
rect 1519 1513 1571 1559
rect 1617 1513 1669 1559
rect 1715 1513 1767 1559
rect 1813 1513 1865 1559
rect 1911 1513 1963 1559
rect 2009 1513 2061 1559
rect 2107 1513 2159 1559
rect 2205 1513 2257 1559
rect 2303 1513 2355 1559
rect 2401 1513 2453 1559
rect 2499 1513 2551 1559
rect 2597 1513 2649 1559
rect 2695 1513 2747 1559
rect 2793 1513 2845 1559
rect 2891 1513 2943 1559
rect 2989 1513 3041 1559
rect 3087 1513 3139 1559
rect 3185 1513 3202 1559
rect -210 1496 3202 1513
rect -210 1461 -130 1496
rect -210 1415 -193 1461
rect -147 1415 -130 1461
rect -210 1363 -130 1415
rect -210 1317 -193 1363
rect -147 1317 -130 1363
rect -210 1265 -130 1317
rect 3122 1461 3202 1496
rect 3122 1415 3139 1461
rect 3185 1415 3202 1461
rect 3122 1363 3202 1415
rect 3122 1317 3139 1363
rect 3185 1317 3202 1363
rect -210 1219 -193 1265
rect -147 1219 -130 1265
rect -210 1167 -130 1219
rect -210 1121 -193 1167
rect -147 1121 -130 1167
rect -210 1069 -130 1121
rect -210 1023 -193 1069
rect -147 1023 -130 1069
rect -210 971 -130 1023
rect -210 925 -193 971
rect -147 925 -130 971
rect -210 873 -130 925
rect -210 827 -193 873
rect -147 827 -130 873
rect -210 775 -130 827
rect -210 729 -193 775
rect -147 729 -130 775
rect -210 677 -130 729
rect -210 631 -193 677
rect -147 631 -130 677
rect -210 579 -130 631
rect -210 533 -193 579
rect -147 533 -130 579
rect -210 481 -130 533
rect -210 435 -193 481
rect -147 435 -130 481
rect -210 383 -130 435
rect -210 337 -193 383
rect -147 337 -130 383
rect -210 285 -130 337
rect -210 239 -193 285
rect -147 239 -130 285
rect -210 187 -130 239
rect -210 141 -193 187
rect -147 141 -130 187
rect -210 89 -130 141
rect -210 43 -193 89
rect -147 43 -130 89
rect -210 -9 -130 43
rect -210 -55 -193 -9
rect -147 -55 -130 -9
rect -210 -107 -130 -55
rect -210 -153 -193 -107
rect -147 -153 -130 -107
rect -210 -205 -130 -153
rect -210 -251 -193 -205
rect -147 -251 -130 -205
rect -210 -303 -130 -251
rect -210 -349 -193 -303
rect -147 -349 -130 -303
rect -210 -401 -130 -349
rect -210 -447 -193 -401
rect -147 -447 -130 -401
rect -210 -499 -130 -447
rect -210 -545 -193 -499
rect -147 -545 -130 -499
rect -210 -597 -130 -545
rect -210 -643 -193 -597
rect -147 -643 -130 -597
rect -210 -695 -130 -643
rect -210 -741 -193 -695
rect -147 -741 -130 -695
rect -210 -793 -130 -741
rect -210 -839 -193 -793
rect -147 -839 -130 -793
rect -210 -891 -130 -839
rect -210 -937 -193 -891
rect -147 -937 -130 -891
rect -210 -989 -130 -937
rect -210 -1035 -193 -989
rect -147 -1035 -130 -989
rect -210 -1087 -130 -1035
rect -210 -1133 -193 -1087
rect -147 -1133 -130 -1087
rect -210 -1185 -130 -1133
rect -210 -1231 -193 -1185
rect -147 -1231 -130 -1185
rect -210 -1283 -130 -1231
rect -36 1196 3004 1268
rect -36 36 36 1196
rect 2932 36 3004 1196
rect -36 -36 3004 36
rect -36 -1196 36 -36
rect 2932 -1196 3004 -36
rect -36 -1268 3004 -1196
rect 3122 1265 3202 1317
rect 3122 1219 3139 1265
rect 3185 1219 3202 1265
rect 3122 1167 3202 1219
rect 3122 1121 3139 1167
rect 3185 1121 3202 1167
rect 3122 1069 3202 1121
rect 3122 1023 3139 1069
rect 3185 1023 3202 1069
rect 3122 971 3202 1023
rect 3122 925 3139 971
rect 3185 925 3202 971
rect 3122 873 3202 925
rect 3122 827 3139 873
rect 3185 827 3202 873
rect 3122 775 3202 827
rect 3122 729 3139 775
rect 3185 729 3202 775
rect 3122 677 3202 729
rect 3122 631 3139 677
rect 3185 631 3202 677
rect 3122 579 3202 631
rect 3122 533 3139 579
rect 3185 533 3202 579
rect 3122 481 3202 533
rect 3122 435 3139 481
rect 3185 435 3202 481
rect 3122 383 3202 435
rect 3122 337 3139 383
rect 3185 337 3202 383
rect 3122 285 3202 337
rect 3122 239 3139 285
rect 3185 239 3202 285
rect 3122 187 3202 239
rect 3122 141 3139 187
rect 3185 141 3202 187
rect 3122 89 3202 141
rect 3122 43 3139 89
rect 3185 43 3202 89
rect 3122 -9 3202 43
rect 3122 -55 3139 -9
rect 3185 -55 3202 -9
rect 3122 -107 3202 -55
rect 3122 -153 3139 -107
rect 3185 -153 3202 -107
rect 3122 -205 3202 -153
rect 3122 -251 3139 -205
rect 3185 -251 3202 -205
rect 3122 -303 3202 -251
rect 3122 -349 3139 -303
rect 3185 -349 3202 -303
rect 3122 -401 3202 -349
rect 3122 -447 3139 -401
rect 3185 -447 3202 -401
rect 3122 -499 3202 -447
rect 3122 -545 3139 -499
rect 3185 -545 3202 -499
rect 3122 -597 3202 -545
rect 3122 -643 3139 -597
rect 3185 -643 3202 -597
rect 3122 -695 3202 -643
rect 3122 -741 3139 -695
rect 3185 -741 3202 -695
rect 3122 -793 3202 -741
rect 3122 -839 3139 -793
rect 3185 -839 3202 -793
rect 3122 -891 3202 -839
rect 3122 -937 3139 -891
rect 3185 -937 3202 -891
rect 3122 -989 3202 -937
rect 3122 -1035 3139 -989
rect 3185 -1035 3202 -989
rect 3122 -1087 3202 -1035
rect 3122 -1133 3139 -1087
rect 3185 -1133 3202 -1087
rect 3122 -1185 3202 -1133
rect 3122 -1231 3139 -1185
rect 3185 -1231 3202 -1185
rect -210 -1329 -193 -1283
rect -147 -1329 -130 -1283
rect -210 -1381 -130 -1329
rect -210 -1427 -193 -1381
rect -147 -1427 -130 -1381
rect -210 -1462 -130 -1427
rect 3122 -1283 3202 -1231
rect 3122 -1329 3139 -1283
rect 3185 -1329 3202 -1283
rect 3122 -1381 3202 -1329
rect 3122 -1427 3139 -1381
rect 3185 -1427 3202 -1381
rect 3122 -1462 3202 -1427
rect -210 -1479 3202 -1462
rect -210 -1525 -193 -1479
rect -147 -1525 -95 -1479
rect -49 -1525 3 -1479
rect 49 -1525 101 -1479
rect 147 -1525 199 -1479
rect 245 -1525 297 -1479
rect 343 -1525 395 -1479
rect 441 -1525 493 -1479
rect 539 -1525 591 -1479
rect 637 -1525 689 -1479
rect 735 -1525 787 -1479
rect 833 -1525 885 -1479
rect 931 -1525 983 -1479
rect 1029 -1525 1081 -1479
rect 1127 -1525 1179 -1479
rect 1225 -1525 1277 -1479
rect 1323 -1525 1375 -1479
rect 1421 -1525 1473 -1479
rect 1519 -1525 1571 -1479
rect 1617 -1525 1669 -1479
rect 1715 -1525 1767 -1479
rect 1813 -1525 1865 -1479
rect 1911 -1525 1963 -1479
rect 2009 -1525 2061 -1479
rect 2107 -1525 2159 -1479
rect 2205 -1525 2257 -1479
rect 2303 -1525 2355 -1479
rect 2401 -1525 2453 -1479
rect 2499 -1525 2551 -1479
rect 2597 -1525 2649 -1479
rect 2695 -1525 2747 -1479
rect 2793 -1525 2845 -1479
rect 2891 -1525 2943 -1479
rect 2989 -1525 3041 -1479
rect 3087 -1525 3139 -1479
rect 3185 -1525 3202 -1479
rect -210 -1542 3202 -1525
<< nsubdiffcont >>
rect -193 1513 -147 1559
rect -95 1513 -49 1559
rect 3 1513 49 1559
rect 101 1513 147 1559
rect 199 1513 245 1559
rect 297 1513 343 1559
rect 395 1513 441 1559
rect 493 1513 539 1559
rect 591 1513 637 1559
rect 689 1513 735 1559
rect 787 1513 833 1559
rect 885 1513 931 1559
rect 983 1513 1029 1559
rect 1081 1513 1127 1559
rect 1179 1513 1225 1559
rect 1277 1513 1323 1559
rect 1375 1513 1421 1559
rect 1473 1513 1519 1559
rect 1571 1513 1617 1559
rect 1669 1513 1715 1559
rect 1767 1513 1813 1559
rect 1865 1513 1911 1559
rect 1963 1513 2009 1559
rect 2061 1513 2107 1559
rect 2159 1513 2205 1559
rect 2257 1513 2303 1559
rect 2355 1513 2401 1559
rect 2453 1513 2499 1559
rect 2551 1513 2597 1559
rect 2649 1513 2695 1559
rect 2747 1513 2793 1559
rect 2845 1513 2891 1559
rect 2943 1513 2989 1559
rect 3041 1513 3087 1559
rect 3139 1513 3185 1559
rect -193 1415 -147 1461
rect -193 1317 -147 1363
rect 3139 1415 3185 1461
rect 3139 1317 3185 1363
rect -193 1219 -147 1265
rect -193 1121 -147 1167
rect -193 1023 -147 1069
rect -193 925 -147 971
rect -193 827 -147 873
rect -193 729 -147 775
rect -193 631 -147 677
rect -193 533 -147 579
rect -193 435 -147 481
rect -193 337 -147 383
rect -193 239 -147 285
rect -193 141 -147 187
rect -193 43 -147 89
rect -193 -55 -147 -9
rect -193 -153 -147 -107
rect -193 -251 -147 -205
rect -193 -349 -147 -303
rect -193 -447 -147 -401
rect -193 -545 -147 -499
rect -193 -643 -147 -597
rect -193 -741 -147 -695
rect -193 -839 -147 -793
rect -193 -937 -147 -891
rect -193 -1035 -147 -989
rect -193 -1133 -147 -1087
rect -193 -1231 -147 -1185
rect 3139 1219 3185 1265
rect 3139 1121 3185 1167
rect 3139 1023 3185 1069
rect 3139 925 3185 971
rect 3139 827 3185 873
rect 3139 729 3185 775
rect 3139 631 3185 677
rect 3139 533 3185 579
rect 3139 435 3185 481
rect 3139 337 3185 383
rect 3139 239 3185 285
rect 3139 141 3185 187
rect 3139 43 3185 89
rect 3139 -55 3185 -9
rect 3139 -153 3185 -107
rect 3139 -251 3185 -205
rect 3139 -349 3185 -303
rect 3139 -447 3185 -401
rect 3139 -545 3185 -499
rect 3139 -643 3185 -597
rect 3139 -741 3185 -695
rect 3139 -839 3185 -793
rect 3139 -937 3185 -891
rect 3139 -1035 3185 -989
rect 3139 -1133 3185 -1087
rect 3139 -1231 3185 -1185
rect -193 -1329 -147 -1283
rect -193 -1427 -147 -1381
rect 3139 -1329 3185 -1283
rect 3139 -1427 3185 -1381
rect -193 -1525 -147 -1479
rect -95 -1525 -49 -1479
rect 3 -1525 49 -1479
rect 101 -1525 147 -1479
rect 199 -1525 245 -1479
rect 297 -1525 343 -1479
rect 395 -1525 441 -1479
rect 493 -1525 539 -1479
rect 591 -1525 637 -1479
rect 689 -1525 735 -1479
rect 787 -1525 833 -1479
rect 885 -1525 931 -1479
rect 983 -1525 1029 -1479
rect 1081 -1525 1127 -1479
rect 1179 -1525 1225 -1479
rect 1277 -1525 1323 -1479
rect 1375 -1525 1421 -1479
rect 1473 -1525 1519 -1479
rect 1571 -1525 1617 -1479
rect 1669 -1525 1715 -1479
rect 1767 -1525 1813 -1479
rect 1865 -1525 1911 -1479
rect 1963 -1525 2009 -1479
rect 2061 -1525 2107 -1479
rect 2159 -1525 2205 -1479
rect 2257 -1525 2303 -1479
rect 2355 -1525 2401 -1479
rect 2453 -1525 2499 -1479
rect 2551 -1525 2597 -1479
rect 2649 -1525 2695 -1479
rect 2747 -1525 2793 -1479
rect 2845 -1525 2891 -1479
rect 2943 -1525 2989 -1479
rect 3041 -1525 3087 -1479
rect 3139 -1525 3185 -1479
<< polysilicon >>
rect 124 1095 324 1108
rect 124 1049 137 1095
rect 311 1049 324 1095
rect 124 1006 324 1049
rect 124 183 324 226
rect 124 137 137 183
rect 311 137 324 183
rect 124 124 324 137
rect 404 1095 604 1108
rect 404 1049 417 1095
rect 591 1049 604 1095
rect 404 1006 604 1049
rect 404 183 604 226
rect 404 137 417 183
rect 591 137 604 183
rect 404 124 604 137
rect 684 1095 884 1108
rect 684 1049 697 1095
rect 871 1049 884 1095
rect 684 1006 884 1049
rect 684 183 884 226
rect 684 137 697 183
rect 871 137 884 183
rect 684 124 884 137
rect 964 1095 1164 1108
rect 964 1049 977 1095
rect 1151 1049 1164 1095
rect 964 1006 1164 1049
rect 964 183 1164 226
rect 964 137 977 183
rect 1151 137 1164 183
rect 964 124 1164 137
rect 1244 1095 1444 1108
rect 1244 1049 1257 1095
rect 1431 1049 1444 1095
rect 1244 1006 1444 1049
rect 1244 183 1444 226
rect 1244 137 1257 183
rect 1431 137 1444 183
rect 1244 124 1444 137
rect 1524 1095 1724 1108
rect 1524 1049 1537 1095
rect 1711 1049 1724 1095
rect 1524 1006 1724 1049
rect 1524 183 1724 226
rect 1524 137 1537 183
rect 1711 137 1724 183
rect 1524 124 1724 137
rect 1804 1095 2004 1108
rect 1804 1049 1817 1095
rect 1991 1049 2004 1095
rect 1804 1006 2004 1049
rect 1804 183 2004 226
rect 1804 137 1817 183
rect 1991 137 2004 183
rect 1804 124 2004 137
rect 2084 1095 2284 1108
rect 2084 1049 2097 1095
rect 2271 1049 2284 1095
rect 2084 1006 2284 1049
rect 2084 183 2284 226
rect 2084 137 2097 183
rect 2271 137 2284 183
rect 2084 124 2284 137
rect 2364 1095 2564 1108
rect 2364 1049 2377 1095
rect 2551 1049 2564 1095
rect 2364 1006 2564 1049
rect 2364 183 2564 226
rect 2364 137 2377 183
rect 2551 137 2564 183
rect 2364 124 2564 137
rect 2644 1095 2844 1108
rect 2644 1049 2657 1095
rect 2831 1049 2844 1095
rect 2644 1006 2844 1049
rect 2644 183 2844 226
rect 2644 137 2657 183
rect 2831 137 2844 183
rect 2644 124 2844 137
rect 124 -137 324 -124
rect 124 -183 137 -137
rect 311 -183 324 -137
rect 124 -226 324 -183
rect 124 -1049 324 -1006
rect 124 -1095 137 -1049
rect 311 -1095 324 -1049
rect 124 -1108 324 -1095
rect 404 -137 604 -124
rect 404 -183 417 -137
rect 591 -183 604 -137
rect 404 -226 604 -183
rect 404 -1049 604 -1006
rect 404 -1095 417 -1049
rect 591 -1095 604 -1049
rect 404 -1108 604 -1095
rect 684 -137 884 -124
rect 684 -183 697 -137
rect 871 -183 884 -137
rect 684 -226 884 -183
rect 684 -1049 884 -1006
rect 684 -1095 697 -1049
rect 871 -1095 884 -1049
rect 684 -1108 884 -1095
rect 964 -137 1164 -124
rect 964 -183 977 -137
rect 1151 -183 1164 -137
rect 964 -226 1164 -183
rect 964 -1049 1164 -1006
rect 964 -1095 977 -1049
rect 1151 -1095 1164 -1049
rect 964 -1108 1164 -1095
rect 1244 -137 1444 -124
rect 1244 -183 1257 -137
rect 1431 -183 1444 -137
rect 1244 -226 1444 -183
rect 1244 -1049 1444 -1006
rect 1244 -1095 1257 -1049
rect 1431 -1095 1444 -1049
rect 1244 -1108 1444 -1095
rect 1524 -137 1724 -124
rect 1524 -183 1537 -137
rect 1711 -183 1724 -137
rect 1524 -226 1724 -183
rect 1524 -1049 1724 -1006
rect 1524 -1095 1537 -1049
rect 1711 -1095 1724 -1049
rect 1524 -1108 1724 -1095
rect 1804 -137 2004 -124
rect 1804 -183 1817 -137
rect 1991 -183 2004 -137
rect 1804 -226 2004 -183
rect 1804 -1049 2004 -1006
rect 1804 -1095 1817 -1049
rect 1991 -1095 2004 -1049
rect 1804 -1108 2004 -1095
rect 2084 -137 2284 -124
rect 2084 -183 2097 -137
rect 2271 -183 2284 -137
rect 2084 -226 2284 -183
rect 2084 -1049 2284 -1006
rect 2084 -1095 2097 -1049
rect 2271 -1095 2284 -1049
rect 2084 -1108 2284 -1095
rect 2364 -137 2564 -124
rect 2364 -183 2377 -137
rect 2551 -183 2564 -137
rect 2364 -226 2564 -183
rect 2364 -1049 2564 -1006
rect 2364 -1095 2377 -1049
rect 2551 -1095 2564 -1049
rect 2364 -1108 2564 -1095
rect 2644 -137 2844 -124
rect 2644 -183 2657 -137
rect 2831 -183 2844 -137
rect 2644 -226 2844 -183
rect 2644 -1049 2844 -1006
rect 2644 -1095 2657 -1049
rect 2831 -1095 2844 -1049
rect 2644 -1108 2844 -1095
<< polycontact >>
rect 137 1049 311 1095
rect 137 137 311 183
rect 417 1049 591 1095
rect 417 137 591 183
rect 697 1049 871 1095
rect 697 137 871 183
rect 977 1049 1151 1095
rect 977 137 1151 183
rect 1257 1049 1431 1095
rect 1257 137 1431 183
rect 1537 1049 1711 1095
rect 1537 137 1711 183
rect 1817 1049 1991 1095
rect 1817 137 1991 183
rect 2097 1049 2271 1095
rect 2097 137 2271 183
rect 2377 1049 2551 1095
rect 2377 137 2551 183
rect 2657 1049 2831 1095
rect 2657 137 2831 183
rect 137 -183 311 -137
rect 137 -1095 311 -1049
rect 417 -183 591 -137
rect 417 -1095 591 -1049
rect 697 -183 871 -137
rect 697 -1095 871 -1049
rect 977 -183 1151 -137
rect 977 -1095 1151 -1049
rect 1257 -183 1431 -137
rect 1257 -1095 1431 -1049
rect 1537 -183 1711 -137
rect 1537 -1095 1711 -1049
rect 1817 -183 1991 -137
rect 1817 -1095 1991 -1049
rect 2097 -183 2271 -137
rect 2097 -1095 2271 -1049
rect 2377 -183 2551 -137
rect 2377 -1095 2551 -1049
rect 2657 -183 2831 -137
rect 2657 -1095 2831 -1049
<< ppolyres >>
rect 124 226 324 1006
rect 404 226 604 1006
rect 684 226 884 1006
rect 964 226 1164 1006
rect 1244 226 1444 1006
rect 1524 226 1724 1006
rect 1804 226 2004 1006
rect 2084 226 2284 1006
rect 2364 226 2564 1006
rect 2644 226 2844 1006
rect 124 -1006 324 -226
rect 404 -1006 604 -226
rect 684 -1006 884 -226
rect 964 -1006 1164 -226
rect 1244 -1006 1444 -226
rect 1524 -1006 1724 -226
rect 1804 -1006 2004 -226
rect 2084 -1006 2284 -226
rect 2364 -1006 2564 -226
rect 2644 -1006 2844 -226
<< metal1 >>
rect -210 1559 3202 1576
rect -210 1513 -193 1559
rect -147 1513 -95 1559
rect -49 1513 3 1559
rect 49 1513 101 1559
rect 147 1513 199 1559
rect 245 1513 297 1559
rect 343 1513 395 1559
rect 441 1513 493 1559
rect 539 1513 591 1559
rect 637 1513 689 1559
rect 735 1513 787 1559
rect 833 1513 885 1559
rect 931 1513 983 1559
rect 1029 1513 1081 1559
rect 1127 1513 1179 1559
rect 1225 1513 1277 1559
rect 1323 1513 1375 1559
rect 1421 1513 1473 1559
rect 1519 1513 1571 1559
rect 1617 1513 1669 1559
rect 1715 1513 1767 1559
rect 1813 1513 1865 1559
rect 1911 1513 1963 1559
rect 2009 1513 2061 1559
rect 2107 1513 2159 1559
rect 2205 1513 2257 1559
rect 2303 1513 2355 1559
rect 2401 1513 2453 1559
rect 2499 1513 2551 1559
rect 2597 1513 2649 1559
rect 2695 1513 2747 1559
rect 2793 1513 2845 1559
rect 2891 1513 2943 1559
rect 2989 1513 3041 1559
rect 3087 1513 3139 1559
rect 3185 1513 3202 1559
rect -210 1496 3202 1513
rect -210 1461 -130 1496
rect -210 1415 -193 1461
rect -147 1415 -130 1461
rect -210 1363 -130 1415
rect 3122 1461 3202 1496
rect 3122 1415 3139 1461
rect 3185 1415 3202 1461
rect -210 1317 -193 1363
rect -147 1317 -130 1363
rect -210 1265 -130 1317
rect -210 1219 -193 1265
rect -147 1219 -130 1265
rect -210 1167 -130 1219
rect -210 1121 -193 1167
rect -147 1121 -130 1167
rect -210 1103 -130 1121
rect 406 1357 2282 1382
rect 406 1301 709 1357
rect 765 1301 819 1357
rect 875 1301 929 1357
rect 985 1301 1039 1357
rect 1095 1301 1149 1357
rect 1205 1301 2282 1357
rect 406 1247 2282 1301
rect 406 1191 709 1247
rect 765 1191 819 1247
rect 875 1191 929 1247
rect 985 1191 1039 1247
rect 1095 1191 1149 1247
rect 1205 1191 2282 1247
rect 406 1155 2282 1191
rect -210 1095 240 1103
rect 406 1095 602 1155
rect 966 1095 1162 1155
rect 1526 1095 1722 1155
rect 2086 1095 2282 1155
rect 3122 1363 3202 1415
rect 3122 1317 3139 1363
rect 3185 1317 3202 1363
rect 3122 1265 3202 1317
rect 3122 1219 3139 1265
rect 3185 1219 3202 1265
rect 3122 1167 3202 1219
rect 3122 1121 3139 1167
rect 3185 1121 3202 1167
rect 3122 1101 3202 1121
rect -210 1069 137 1095
rect -210 1023 -193 1069
rect -147 1049 137 1069
rect 311 1049 322 1095
rect 406 1049 417 1095
rect 591 1049 602 1095
rect 686 1049 697 1095
rect 871 1049 882 1095
rect 966 1049 977 1095
rect 1151 1049 1162 1095
rect 1246 1049 1257 1095
rect 1431 1049 1442 1095
rect 1526 1049 1537 1095
rect 1711 1049 1722 1095
rect 1806 1049 1817 1095
rect 1991 1049 2002 1095
rect 2086 1049 2097 1095
rect 2271 1049 2282 1095
rect 2366 1095 2561 1096
rect 2773 1095 3202 1101
rect 2366 1049 2377 1095
rect 2551 1049 2562 1095
rect 2646 1049 2657 1095
rect 2831 1069 3202 1095
rect 2831 1049 3139 1069
rect -147 1032 240 1049
rect -147 1023 -130 1032
rect -210 971 -130 1023
rect -210 925 -193 971
rect -147 925 -130 971
rect -210 873 -130 925
rect -210 827 -193 873
rect -147 827 -130 873
rect -210 775 -130 827
rect -210 729 -193 775
rect -147 729 -130 775
rect 686 989 882 1049
rect 1246 989 1441 1049
rect 1806 989 2001 1049
rect 2366 989 2561 1049
rect 2773 1030 3139 1049
rect 686 943 2561 989
rect 686 887 1771 943
rect 1827 887 1881 943
rect 1937 887 1991 943
rect 2047 887 2101 943
rect 2157 887 2211 943
rect 2267 887 2561 943
rect 686 833 2561 887
rect 686 777 1771 833
rect 1827 777 1881 833
rect 1937 777 1991 833
rect 2047 777 2101 833
rect 2157 777 2211 833
rect 2267 777 2561 833
rect 686 762 2561 777
rect 3122 1023 3139 1030
rect 3185 1023 3202 1069
rect 3122 971 3202 1023
rect 3122 925 3139 971
rect 3185 925 3202 971
rect 3122 873 3202 925
rect 3122 827 3139 873
rect 3185 827 3202 873
rect 3122 775 3202 827
rect -210 677 -130 729
rect -210 631 -193 677
rect -147 631 -130 677
rect -210 579 -130 631
rect -210 533 -193 579
rect -147 533 -130 579
rect -210 481 -130 533
rect -210 435 -193 481
rect -147 435 -130 481
rect -210 383 -130 435
rect -210 337 -193 383
rect -147 337 -130 383
rect -210 285 -130 337
rect -210 239 -193 285
rect -147 239 -130 285
rect -210 197 -130 239
rect 3122 729 3139 775
rect 3185 729 3202 775
rect 3122 677 3202 729
rect 3122 631 3139 677
rect 3185 631 3202 677
rect 3122 579 3202 631
rect 3122 533 3139 579
rect 3185 533 3202 579
rect 3122 481 3202 533
rect 3122 435 3139 481
rect 3185 435 3202 481
rect 3122 383 3202 435
rect 3122 337 3139 383
rect 3185 337 3202 383
rect 3122 285 3202 337
rect 3122 239 3139 285
rect 3185 239 3202 285
rect 3122 198 3202 239
rect -210 187 229 197
rect -210 141 -193 187
rect -147 183 229 187
rect 2764 187 3202 198
rect 2764 183 3139 187
rect -147 141 137 183
rect -210 137 137 141
rect 311 137 322 183
rect -210 126 229 137
rect -210 89 -130 126
rect -210 43 -193 89
rect -147 43 -130 89
rect -210 -9 -130 43
rect -210 -55 -193 -9
rect -147 -55 -130 -9
rect -210 -107 -130 -55
rect -210 -153 -193 -107
rect -147 -129 -130 -107
rect 406 119 417 183
rect 591 137 602 183
rect 473 119 527 137
rect 583 119 602 137
rect 406 82 602 119
rect 686 137 697 183
rect 871 137 882 183
rect 686 82 882 137
rect 966 137 977 183
rect 1151 137 1162 183
rect 966 82 1162 137
rect 1246 137 1257 183
rect 1431 137 1442 183
rect 1246 82 1442 137
rect 1526 137 1537 183
rect 1711 138 1722 183
rect 1711 137 1723 138
rect 1526 82 1723 137
rect 1806 137 1817 183
rect 1991 137 2002 183
rect 1806 82 2002 137
rect 2086 137 2097 183
rect 2271 137 2282 183
rect 2086 82 2282 137
rect 2366 137 2377 183
rect 2551 137 2562 183
rect 2646 137 2657 183
rect 2831 141 3139 183
rect 3185 141 3202 187
rect 2831 137 3202 141
rect 2366 82 2562 137
rect 2764 127 3202 137
rect 406 65 2562 82
rect 406 9 417 65
rect 473 9 527 65
rect 583 9 2562 65
rect 406 -45 2562 9
rect 406 -101 417 -45
rect 473 -101 527 -45
rect 583 -82 2562 -45
rect 583 -101 602 -82
rect -147 -137 238 -129
rect 406 -137 602 -101
rect -147 -153 137 -137
rect -210 -183 137 -153
rect 311 -183 322 -137
rect -210 -200 238 -183
rect -210 -205 -130 -200
rect -210 -251 -193 -205
rect -147 -251 -130 -205
rect 406 -211 417 -137
rect 591 -183 602 -137
rect 686 -137 882 -82
rect 686 -183 697 -137
rect 871 -183 882 -137
rect 966 -137 1162 -82
rect 966 -183 977 -137
rect 1151 -183 1162 -137
rect 1246 -137 1442 -82
rect 1246 -183 1257 -137
rect 1431 -183 1442 -137
rect 1526 -137 1723 -82
rect 1806 -137 2002 -82
rect 1526 -183 1537 -137
rect 1711 -183 1722 -137
rect 1806 -183 1817 -137
rect 1991 -183 2002 -137
rect 2086 -137 2282 -82
rect 2086 -183 2097 -137
rect 2271 -183 2282 -137
rect 2366 -137 2562 -82
rect 3122 89 3202 127
rect 3122 43 3139 89
rect 3185 43 3202 89
rect 3122 -9 3202 43
rect 3122 -55 3139 -9
rect 3185 -55 3202 -9
rect 3122 -107 3202 -55
rect 3122 -130 3139 -107
rect 2771 -137 3139 -130
rect 2366 -183 2377 -137
rect 2551 -183 2562 -137
rect 2646 -183 2657 -137
rect 2831 -153 3139 -137
rect 3185 -153 3202 -107
rect 2831 -183 3202 -153
rect 473 -211 527 -183
rect 583 -211 602 -183
rect 2771 -201 3202 -183
rect 406 -228 602 -211
rect 3122 -205 3202 -201
rect -210 -303 -130 -251
rect -210 -349 -193 -303
rect -147 -349 -130 -303
rect -210 -401 -130 -349
rect -210 -447 -193 -401
rect -147 -447 -130 -401
rect -210 -499 -130 -447
rect -210 -545 -193 -499
rect -147 -545 -130 -499
rect -210 -597 -130 -545
rect -210 -643 -193 -597
rect -147 -643 -130 -597
rect -210 -695 -130 -643
rect -210 -741 -193 -695
rect -147 -741 -130 -695
rect -210 -793 -130 -741
rect 3122 -251 3139 -205
rect 3185 -251 3202 -205
rect 3122 -303 3202 -251
rect 3122 -349 3139 -303
rect 3185 -349 3202 -303
rect 3122 -401 3202 -349
rect 3122 -447 3139 -401
rect 3185 -447 3202 -401
rect 3122 -499 3202 -447
rect 3122 -545 3139 -499
rect 3185 -545 3202 -499
rect 3122 -597 3202 -545
rect 3122 -643 3139 -597
rect 3185 -643 3202 -597
rect 3122 -695 3202 -643
rect 3122 -741 3139 -695
rect 3185 -741 3202 -695
rect -210 -839 -193 -793
rect -147 -839 -130 -793
rect -210 -891 -130 -839
rect -210 -937 -193 -891
rect -147 -937 -130 -891
rect -210 -989 -130 -937
rect -210 -1035 -193 -989
rect -147 -1035 -130 -989
rect 686 -799 2562 -762
rect 686 -855 702 -799
rect 758 -855 812 -799
rect 868 -855 922 -799
rect 978 -855 1032 -799
rect 1088 -855 1142 -799
rect 1198 -855 2562 -799
rect 686 -909 2562 -855
rect 686 -965 702 -909
rect 758 -965 812 -909
rect 868 -965 922 -909
rect 978 -965 1032 -909
rect 1088 -965 1142 -909
rect 1198 -965 2562 -909
rect 686 -989 2562 -965
rect -210 -1049 234 -1035
rect 686 -1049 882 -989
rect 1246 -1049 1442 -989
rect 1806 -1049 2002 -989
rect 2366 -1049 2562 -989
rect 3122 -793 3202 -741
rect 3122 -839 3139 -793
rect 3185 -839 3202 -793
rect 3122 -891 3202 -839
rect 3122 -937 3139 -891
rect 3185 -937 3202 -891
rect 3122 -989 3202 -937
rect 3122 -1032 3139 -989
rect 2747 -1035 3139 -1032
rect 3185 -1035 3202 -989
rect 2747 -1049 3202 -1035
rect -210 -1087 137 -1049
rect -210 -1133 -193 -1087
rect -147 -1095 137 -1087
rect 311 -1095 322 -1049
rect 406 -1095 417 -1049
rect 591 -1095 602 -1049
rect 686 -1095 697 -1049
rect 871 -1095 882 -1049
rect 966 -1095 977 -1049
rect 1151 -1095 1162 -1049
rect 1246 -1095 1257 -1049
rect 1431 -1095 1442 -1049
rect 1526 -1095 1537 -1049
rect 1711 -1095 1722 -1049
rect 1806 -1095 1817 -1049
rect 1991 -1095 2002 -1049
rect 2086 -1095 2097 -1049
rect 2271 -1095 2282 -1049
rect 2366 -1095 2377 -1049
rect 2551 -1095 2562 -1049
rect 2646 -1095 2657 -1049
rect 2831 -1087 3202 -1049
rect 2831 -1095 3139 -1087
rect -147 -1106 234 -1095
rect -147 -1133 -130 -1106
rect -210 -1185 -130 -1133
rect -210 -1231 -193 -1185
rect -147 -1231 -130 -1185
rect -210 -1283 -130 -1231
rect -210 -1329 -193 -1283
rect -147 -1329 -130 -1283
rect -210 -1381 -130 -1329
rect -210 -1427 -193 -1381
rect -147 -1427 -130 -1381
rect 406 -1155 602 -1095
rect 966 -1155 1162 -1095
rect 1526 -1155 1722 -1095
rect 2086 -1155 2282 -1095
rect 2747 -1103 3139 -1095
rect 406 -1183 2282 -1155
rect 406 -1239 1730 -1183
rect 1786 -1239 1840 -1183
rect 1896 -1239 1950 -1183
rect 2006 -1239 2060 -1183
rect 2116 -1239 2170 -1183
rect 2226 -1239 2282 -1183
rect 406 -1293 2282 -1239
rect 406 -1349 1730 -1293
rect 1786 -1349 1840 -1293
rect 1896 -1349 1950 -1293
rect 2006 -1349 2060 -1293
rect 2116 -1349 2170 -1293
rect 2226 -1349 2282 -1293
rect 406 -1382 2282 -1349
rect 3122 -1133 3139 -1103
rect 3185 -1133 3202 -1087
rect 3122 -1185 3202 -1133
rect 3122 -1231 3139 -1185
rect 3185 -1231 3202 -1185
rect 3122 -1283 3202 -1231
rect 3122 -1329 3139 -1283
rect 3185 -1329 3202 -1283
rect 3122 -1381 3202 -1329
rect -210 -1462 -130 -1427
rect 3122 -1427 3139 -1381
rect 3185 -1427 3202 -1381
rect 3122 -1462 3202 -1427
rect -210 -1479 3202 -1462
rect -210 -1525 -193 -1479
rect -147 -1525 -95 -1479
rect -49 -1525 3 -1479
rect 49 -1525 101 -1479
rect 147 -1525 199 -1479
rect 245 -1525 297 -1479
rect 343 -1525 395 -1479
rect 441 -1525 493 -1479
rect 539 -1525 591 -1479
rect 637 -1525 689 -1479
rect 735 -1525 787 -1479
rect 833 -1525 885 -1479
rect 931 -1525 983 -1479
rect 1029 -1525 1081 -1479
rect 1127 -1525 1179 -1479
rect 1225 -1525 1277 -1479
rect 1323 -1525 1375 -1479
rect 1421 -1525 1473 -1479
rect 1519 -1525 1571 -1479
rect 1617 -1525 1669 -1479
rect 1715 -1525 1767 -1479
rect 1813 -1525 1865 -1479
rect 1911 -1525 1963 -1479
rect 2009 -1525 2061 -1479
rect 2107 -1525 2159 -1479
rect 2205 -1525 2257 -1479
rect 2303 -1525 2355 -1479
rect 2401 -1525 2453 -1479
rect 2499 -1525 2551 -1479
rect 2597 -1525 2649 -1479
rect 2695 -1525 2747 -1479
rect 2793 -1525 2845 -1479
rect 2891 -1525 2943 -1479
rect 2989 -1525 3041 -1479
rect 3087 -1525 3139 -1479
rect 3185 -1525 3202 -1479
rect -210 -1542 3202 -1525
<< via1 >>
rect 709 1301 765 1357
rect 819 1301 875 1357
rect 929 1301 985 1357
rect 1039 1301 1095 1357
rect 1149 1301 1205 1357
rect 709 1191 765 1247
rect 819 1191 875 1247
rect 929 1191 985 1247
rect 1039 1191 1095 1247
rect 1149 1191 1205 1247
rect 1771 887 1827 943
rect 1881 887 1937 943
rect 1991 887 2047 943
rect 2101 887 2157 943
rect 2211 887 2267 943
rect 1771 777 1827 833
rect 1881 777 1937 833
rect 1991 777 2047 833
rect 2101 777 2157 833
rect 2211 777 2267 833
rect 417 137 473 175
rect 527 137 583 175
rect 417 119 473 137
rect 527 119 583 137
rect 417 9 473 65
rect 527 9 583 65
rect 417 -101 473 -45
rect 527 -101 583 -45
rect 417 -183 473 -155
rect 527 -183 583 -155
rect 417 -211 473 -183
rect 527 -211 583 -183
rect 702 -855 758 -799
rect 812 -855 868 -799
rect 922 -855 978 -799
rect 1032 -855 1088 -799
rect 1142 -855 1198 -799
rect 702 -965 758 -909
rect 812 -965 868 -909
rect 922 -965 978 -909
rect 1032 -965 1088 -909
rect 1142 -965 1198 -909
rect 1730 -1239 1786 -1183
rect 1840 -1239 1896 -1183
rect 1950 -1239 2006 -1183
rect 2060 -1239 2116 -1183
rect 2170 -1239 2226 -1183
rect 1730 -1349 1786 -1293
rect 1840 -1349 1896 -1293
rect 1950 -1349 2006 -1293
rect 2060 -1349 2116 -1293
rect 2170 -1349 2226 -1293
<< metal2 >>
rect 686 1357 1280 1382
rect 686 1301 709 1357
rect 765 1301 819 1357
rect 875 1301 929 1357
rect 985 1301 1039 1357
rect 1095 1301 1149 1357
rect 1205 1301 1280 1357
rect 686 1247 1280 1301
rect 686 1191 709 1247
rect 765 1191 819 1247
rect 875 1191 929 1247
rect 985 1191 1039 1247
rect 1095 1191 1149 1247
rect 1205 1191 1280 1247
rect 686 1155 1280 1191
rect 406 175 602 183
rect 406 119 417 175
rect 473 119 527 175
rect 583 119 602 175
rect 406 65 602 119
rect 406 9 417 65
rect 473 9 527 65
rect 583 9 602 65
rect 406 -45 602 9
rect 406 -101 417 -45
rect 473 -101 527 -45
rect 583 -101 602 -45
rect 406 -155 602 -101
rect 406 -211 417 -155
rect 473 -211 527 -155
rect 583 -211 602 -155
rect 406 -228 602 -211
rect 686 -762 913 1155
rect 1754 943 2282 989
rect 1754 887 1771 943
rect 1827 887 1881 943
rect 1937 887 1991 943
rect 2047 887 2101 943
rect 2157 887 2211 943
rect 2267 887 2282 943
rect 1754 833 2282 887
rect 1754 777 1771 833
rect 1827 777 1881 833
rect 1937 777 1991 833
rect 2047 777 2101 833
rect 2157 777 2211 833
rect 2267 777 2282 833
rect 1754 762 2282 777
rect 686 -799 1211 -762
rect 686 -855 702 -799
rect 758 -855 812 -799
rect 868 -855 922 -799
rect 978 -855 1032 -799
rect 1088 -855 1142 -799
rect 1198 -855 1211 -799
rect 686 -909 1211 -855
rect 686 -965 702 -909
rect 758 -965 812 -909
rect 868 -965 922 -909
rect 978 -965 1032 -909
rect 1088 -965 1142 -909
rect 1198 -965 1211 -909
rect 686 -989 1211 -965
rect 2055 -1155 2282 762
rect 1688 -1183 2282 -1155
rect 1688 -1239 1730 -1183
rect 1786 -1239 1840 -1183
rect 1896 -1239 1950 -1183
rect 2006 -1239 2060 -1183
rect 2116 -1239 2170 -1183
rect 2226 -1239 2282 -1183
rect 1688 -1293 2282 -1239
rect 1688 -1349 1730 -1293
rect 1786 -1349 1840 -1293
rect 1896 -1349 1950 -1293
rect 2006 -1349 2060 -1293
rect 2116 -1349 2170 -1293
rect 2226 -1349 2282 -1293
rect 1688 -1382 2282 -1349
<< labels >>
flabel metal1 533 1310 533 1310 0 FreeSans 800 0 0 0 R1_IN
port 0 nsew
flabel metal1 459 -1284 459 -1284 0 FreeSans 800 0 0 0 R2_IN
port 1 nsew
flabel metal2 491 -27 491 -27 0 FreeSans 800 0 0 0 COMMON
port 2 nsew
flabel metal1 1424 1537 1424 1537 0 FreeSans 800 0 0 0 VDD
port 3 nsew
<< end >>
