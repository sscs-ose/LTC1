magic
tech gf180mcuC
magscale 1 10
timestamp 1693477706
<< nwell >>
rect -15 428 577 524
<< psubdiff >>
rect -146 636 701 650
rect -146 583 -124 636
rect -72 583 1 636
rect 53 583 126 636
rect 178 583 251 636
rect 303 583 376 636
rect 428 583 501 636
rect 553 583 626 636
rect 678 583 701 636
rect -146 560 701 583
rect -146 501 -54 560
rect -146 448 -124 501
rect -72 448 -54 501
rect 611 535 701 560
rect -146 366 -54 448
rect 611 482 625 535
rect 677 482 701 535
rect -146 313 -124 366
rect -72 313 -54 366
rect -146 231 -54 313
rect -146 178 -124 231
rect -72 178 -54 231
rect -146 96 -54 178
rect -146 43 -124 96
rect -72 43 -54 96
rect -146 -39 -54 43
rect 611 400 701 482
rect 611 347 625 400
rect 677 347 701 400
rect 611 265 701 347
rect 611 212 625 265
rect 677 212 701 265
rect 611 130 701 212
rect 611 77 625 130
rect 677 77 701 130
rect -146 -92 -124 -39
rect -72 -92 -54 -39
rect -146 -174 -54 -92
rect 611 -5 701 77
rect 611 -58 625 -5
rect 677 -58 701 -5
rect -146 -227 -124 -174
rect -72 -227 -54 -174
rect -146 -309 -54 -227
rect -146 -362 -124 -309
rect -72 -362 -54 -309
rect -146 -391 -54 -362
rect 611 -140 701 -58
rect 611 -193 625 -140
rect 677 -193 701 -140
rect 611 -275 701 -193
rect 611 -328 625 -275
rect 677 -328 701 -275
rect 611 -391 701 -328
rect -146 -410 701 -391
rect -146 -463 -125 -410
rect -73 -463 0 -410
rect 52 -463 125 -410
rect 177 -463 250 -410
rect 302 -463 375 -410
rect 427 -463 500 -410
rect 552 -463 625 -410
rect 677 -463 701 -410
rect -146 -481 701 -463
<< nsubdiff >>
rect 27 479 534 499
rect 27 432 49 479
rect 95 432 149 479
rect 195 432 249 479
rect 295 432 349 479
rect 395 432 449 479
rect 495 432 534 479
rect 27 411 534 432
<< psubdiffcont >>
rect -124 583 -72 636
rect 1 583 53 636
rect 126 583 178 636
rect 251 583 303 636
rect 376 583 428 636
rect 501 583 553 636
rect 626 583 678 636
rect -124 448 -72 501
rect 625 482 677 535
rect -124 313 -72 366
rect -124 178 -72 231
rect -124 43 -72 96
rect 625 347 677 400
rect 625 212 677 265
rect 625 77 677 130
rect -124 -92 -72 -39
rect 625 -58 677 -5
rect -124 -227 -72 -174
rect -124 -362 -72 -309
rect 625 -193 677 -140
rect 625 -328 677 -275
rect -125 -463 -73 -410
rect 0 -463 52 -410
rect 125 -463 177 -410
rect 250 -463 302 -410
rect 375 -463 427 -410
rect 500 -463 552 -410
rect 625 -463 677 -410
<< nsubdiffcont >>
rect 49 432 95 479
rect 149 432 195 479
rect 249 432 295 479
rect 349 432 395 479
rect 449 432 495 479
<< polysilicon >>
rect 159 0 229 16
rect 79 -13 229 0
rect 333 -13 403 17
rect 79 -82 94 -13
rect 162 -82 403 -13
rect 79 -86 403 -82
rect 79 -95 229 -86
rect 159 -117 229 -95
rect 333 -116 403 -86
<< polycontact >>
rect 94 -82 162 -13
<< metal1 >>
rect -146 636 701 650
rect -146 583 -124 636
rect -72 583 1 636
rect 53 583 126 636
rect 178 583 251 636
rect 303 583 376 636
rect 428 583 501 636
rect 553 583 626 636
rect 678 583 701 636
rect -146 560 701 583
rect -146 501 -54 560
rect -146 448 -124 501
rect -72 448 -54 501
rect 611 535 701 560
rect -146 366 -54 448
rect 27 479 534 499
rect 27 432 49 479
rect 95 432 149 479
rect 195 432 249 479
rect 295 432 349 479
rect 395 432 449 479
rect 495 432 534 479
rect 27 411 534 432
rect 611 482 625 535
rect 677 482 701 535
rect -146 313 -124 366
rect -72 313 -54 366
rect 84 333 130 411
rect 432 334 478 411
rect 611 400 701 482
rect 611 347 625 400
rect 677 347 701 400
rect -146 231 -54 313
rect -146 178 -124 231
rect -72 178 -54 231
rect -146 96 -54 178
rect -146 43 -124 96
rect -72 43 -54 96
rect 611 265 701 347
rect 611 212 625 265
rect 677 212 701 265
rect 611 130 701 212
rect 611 77 625 130
rect 677 77 701 130
rect -146 -39 -54 43
rect 79 -13 173 0
rect 79 -22 94 -13
rect -146 -92 -124 -39
rect -72 -92 -54 -39
rect 10 -74 94 -22
rect -146 -174 -54 -92
rect 79 -82 94 -74
rect 162 -82 173 -13
rect 79 -95 173 -82
rect 258 -35 304 77
rect 611 -5 701 77
rect 258 -81 502 -35
rect 611 -58 625 -5
rect 677 -58 701 -5
rect -146 -227 -124 -174
rect -72 -227 -54 -174
rect 258 -175 304 -81
rect 611 -140 701 -58
rect -146 -309 -54 -227
rect 611 -193 625 -140
rect 677 -193 701 -140
rect -146 -362 -124 -309
rect -72 -362 -54 -309
rect -146 -391 -54 -362
rect 84 -391 131 -263
rect 431 -391 478 -262
rect 611 -275 701 -193
rect 611 -328 625 -275
rect 677 -328 701 -275
rect 611 -391 701 -328
rect -146 -410 701 -391
rect -146 -463 -125 -410
rect -73 -463 0 -410
rect 52 -463 125 -410
rect 177 -463 250 -410
rect 302 -463 375 -410
rect 427 -463 500 -410
rect 552 -463 625 -410
rect 677 -463 701 -410
rect -146 -481 701 -463
use nmos_3p3_9MTZEK  nmos_3p3_9MTZEK_0
timestamp 1693477706
transform 1 0 281 0 1 -229
box -234 -138 234 138
use pmos_3p3_585UPK  pmos_3p3_585UPK_0
timestamp 1693477706
transform 1 0 281 0 1 197
box -296 -270 296 270
<< labels >>
flabel metal1 121 454 121 454 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal1 25 -53 25 -53 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 452 -60 452 -60 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 216 -425 216 -425 0 FreeSans 320 0 0 0 VSS
port 3 nsew
<< end >>
