magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2554 -2242 2554 2242
<< nwell >>
rect -554 -242 554 242
<< pmos >>
rect -380 -112 -268 112
rect -164 -112 -52 112
rect 52 -112 164 112
rect 268 -112 380 112
<< pdiff >>
rect -468 70 -380 112
rect -468 -70 -455 70
rect -409 -70 -380 70
rect -468 -112 -380 -70
rect -268 70 -164 112
rect -268 -70 -239 70
rect -193 -70 -164 70
rect -268 -112 -164 -70
rect -52 70 52 112
rect -52 -70 -23 70
rect 23 -70 52 70
rect -52 -112 52 -70
rect 164 70 268 112
rect 164 -70 193 70
rect 239 -70 268 70
rect 164 -112 268 -70
rect 380 70 468 112
rect 380 -70 409 70
rect 455 -70 468 70
rect 380 -112 468 -70
<< pdiffc >>
rect -455 -70 -409 70
rect -239 -70 -193 70
rect -23 -70 23 70
rect 193 -70 239 70
rect 409 -70 455 70
<< polysilicon >>
rect -380 112 -268 156
rect -164 112 -52 156
rect 52 112 164 156
rect 268 112 380 156
rect -380 -156 -268 -112
rect -164 -156 -52 -112
rect 52 -156 164 -112
rect 268 -156 380 -112
<< metal1 >>
rect -455 70 -409 110
rect -455 -110 -409 -70
rect -239 70 -193 110
rect -239 -110 -193 -70
rect -23 70 23 110
rect -23 -110 23 -70
rect 193 70 239 110
rect 193 -110 239 -70
rect 409 70 455 110
rect 409 -110 455 -70
<< end >>
