* NGSPICE file created from cap_240p_flat.ext - technology: gf180mcuC

.subckt cap_240p_pex P M
X0 P.t0 M.t131 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X1 P.t1 M.t130 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X2 P.t2 M.t129 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X3 P.t3 M.t128 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X4 P.t4 M.t127 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X5 P.t5 M.t126 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X6 P.t6 M.t125 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X7 P.t7 M.t124 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X8 P.t8 M.t123 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X9 P.t9 M.t122 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X10 P.t10 M.t121 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X11 P.t11 M.t120 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X12 P.t12 M.t119 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X13 P.t13 M.t118 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X14 P.t14 M.t117 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X15 P.t15 M.t116 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X16 P.t16 M.t115 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X17 P.t17 M.t114 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X18 P.t18 M.t113 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X19 P.t19 M.t112 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X20 P.t20 M.t111 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X21 P.t21 M.t110 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X22 P.t22 M.t109 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X23 P.t23 M.t108 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X24 P.t24 M.t107 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X25 P.t25 M.t106 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X26 P.t26 M.t105 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X27 P.t27 M.t104 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X28 P.t28 M.t103 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X29 P.t29 M.t102 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X30 P.t30 M.t101 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X31 P.t31 M.t100 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X32 P.t32 M.t99 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X33 P.t33 M.t98 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X34 P.t34 M.t97 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X35 P.t35 M.t96 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X36 P.t36 M.t95 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X37 P.t37 M.t94 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X38 P.t38 M.t93 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X39 P.t39 M.t92 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X40 P.t40 M.t91 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X41 P.t41 M.t90 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X42 P.t42 M.t89 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X43 P.t43 M.t88 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X44 P.t44 M.t87 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X45 P.t45 M.t86 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X46 P.t46 M.t85 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X47 P.t47 M.t84 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X48 P.t48 M.t83 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X49 P.t49 M.t82 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X50 P.t50 M.t81 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X51 P.t51 M.t80 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X52 P.t52 M.t79 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X53 P.t53 M.t78 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X54 P.t54 M.t77 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X55 P.t55 M.t76 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X56 P.t56 M.t75 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X57 P.t57 M.t74 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X58 P.t58 M.t73 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X59 P.t59 M.t72 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X60 P.t60 M.t71 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X61 P.t61 M.t70 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X62 P.t62 M.t69 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X63 P.t63 M.t68 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X64 P.t64 M.t67 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X65 P.t65 M.t66 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X66 P.t66 M.t65 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X67 P.t67 M.t64 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X68 P.t68 M.t63 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X69 P.t69 M.t62 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X70 P.t70 M.t61 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X71 P.t71 M.t60 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X72 P.t72 M.t59 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X73 P.t73 M.t58 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X74 P.t74 M.t57 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X75 P.t75 M.t56 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X76 P.t76 M.t55 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X77 P.t77 M.t54 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X78 P.t78 M.t53 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X79 P.t79 M.t52 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X80 P.t80 M.t51 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X81 P.t81 M.t50 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X82 P.t82 M.t49 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X83 P.t83 M.t48 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X84 P.t84 M.t47 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X85 P.t85 M.t46 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X86 P.t86 M.t45 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X87 P.t87 M.t44 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X88 P.t88 M.t43 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X89 P.t89 M.t42 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X90 P.t90 M.t41 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X91 P.t91 M.t40 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X92 P.t92 M.t39 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X93 P.t93 M.t38 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X94 P.t94 M.t37 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X95 P.t95 M.t36 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X96 P.t96 M.t35 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X97 P.t97 M.t34 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X98 P.t98 M.t33 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X99 P.t99 M.t32 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X100 P.t100 M.t31 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X101 P.t101 M.t30 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X102 P.t102 M.t29 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X103 P.t103 M.t28 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X104 P.t104 M.t27 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X105 P.t105 M.t26 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X106 P.t106 M.t25 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X107 P.t107 M.t24 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X108 P.t108 M.t23 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X109 P.t109 M.t22 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X110 P.t110 M.t21 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X111 P.t111 M.t20 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X112 P.t112 M.t19 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X113 P.t113 M.t18 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X114 P.t114 M.t17 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X115 P.t115 M.t16 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X116 P.t116 M.t15 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X117 P.t117 M.t14 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X118 P.t118 M.t13 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X119 P.t119 M.t12 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X120 P.t120 M.t11 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X121 P.t121 M.t10 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X122 P.t122 M.t9 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X123 P.t123 M.t8 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X124 P.t124 M.t7 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X125 P.t125 M.t6 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X126 P.t126 M.t5 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X127 P.t127 M.t4 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X128 P.t128 M.t3 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X129 P.t129 M.t2 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X130 P.t130 M.t1 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
X131 P.t131 M.t0 cap_mim_2f0_m4m5_noshield c_width=31u c_length=29u
R0 P.n2017 P.t64 2.38596
R1 P.n3106 P.t74 2.38596
R2 P.n2782 P.t18 2.38596
R3 P.n2511 P.t36 2.38596
R4 P.n2192 P.t119 2.38596
R5 P.n0 P.t24 2.38596
R6 P.n11 P.t82 2.38596
R7 P.n22 P.t27 2.38596
R8 P.n33 P.t112 2.38596
R9 P.n44 P.t129 2.38596
R10 P.n62 P.t14 2.38596
R11 P.n720 P.n719 2.25096
R12 P.n636 P.n635 2.25096
R13 P.n329 P.n328 2.25096
R14 P.n190 P.n189 2.25096
R15 P.n93 P.n92 2.25096
R16 P.n346 P.n345 2.25096
R17 P.n354 P.n353 2.25096
R18 P.n900 P.n899 2.25096
R19 P.n1340 P.n1316 2.25096
R20 P.n1400 P.n1399 2.25096
R21 P.n1682 P.n1681 2.25096
R22 P.n876 P.n875 2.25096
R23 P.n754 P.n753 2.25096
R24 P.n512 P.n511 2.25096
R25 P.n1089 P.n1084 2.25096
R26 P.n1355 P.n1347 2.25096
R27 P.n368 P.n367 2.25096
R28 P.n293 P.n292 2.25096
R29 P.n385 P.n384 2.25096
R30 P.n101 P.n100 2.25096
R31 P.n395 P.n394 2.25096
R32 P.n781 P.n780 2.25096
R33 P.n1047 P.n1046 2.25096
R34 P.n1014 P.n1013 2.25096
R35 P.n713 P.n712 2.25096
R36 P.n1089 P.n1088 2.25096
R37 P.n1038 P.n1037 2.25096
R38 P.n1355 P.n1354 2.25096
R39 P.n1294 P.n1207 2.25096
R40 P.n1547 P.n1546 2.25096
R41 P.n1340 P.n1339 2.25096
R42 P.n1674 P.n1673 2.25096
R43 P.n1738 P.n1737 2.25096
R44 P.n1979 P.n1978 2.25096
R45 P.n1642 P.n1641 2.25096
R46 P.n1294 P.n1293 2.25096
R47 P.n1666 P.n1665 2.25096
R48 P.n1719 P.n1718 2.25096
R49 P.n1971 P.n1970 2.25096
R50 P.n2003 P.n2002 2.25096
R51 P.n2010 P.n2009 2.25096
R52 P.n1745 P.n1744 2.25096
R53 P.n1729 P.n1728 2.25096
R54 P.n1523 P.n1522 2.25096
R55 P.n1841 P.n1840 2.25096
R56 P.n1865 P.n1864 2.25096
R57 P.n1076 P.n1075 2.25096
R58 P.n1393 P.n1392 2.25096
R59 P.n766 P.n765 2.25096
R60 P.n774 P.n773 2.25096
R61 P.n908 P.n907 2.25096
R62 P.n309 P.n308 2.25096
R63 P.n523 P.n522 2.25096
R64 P.n626 P.n625 2.25096
R65 P.n697 P.n696 2.25096
R66 P.n677 P.n676 2.25096
R67 P.n654 P.n653 2.25096
R68 P.n670 P.n669 2.25096
R69 P.n302 P.n301 2.25096
R70 P.n3439 P.n2732 2.25095
R71 P.n3436 P.n2743 2.25095
R72 P.n3694 P.n2170 2.25095
R73 P.n3701 P.n2146 2.25095
R74 P.n3516 P.n2446 2.25095
R75 P.n3533 P.n2245 2.25095
R76 P.n3706 P.n2121 2.25095
R77 P.n3704 P.n2132 2.25095
R78 P.n3699 P.n2160 2.25095
R79 P.n3535 P.n2232 2.25095
R80 P.n3504 P.n2451 2.25095
R81 P.n3575 P.n3574 2.25095
R82 P.n3501 P.n2457 2.25095
R83 P.n3485 P.n2467 2.25095
R84 P.n3471 P.n2510 2.25095
R85 P.n3305 P.n2919 2.25095
R86 P.n3292 P.n2924 2.25095
R87 P.n3402 P.n2781 2.25095
R88 P.n3476 P.n2484 2.25095
R89 P.n3397 P.n3396 2.25095
R90 P.n3397 P.n2913 2.25095
R91 P.n3540 P.n2211 2.25095
R92 P.n3473 P.n2497 2.25095
R93 P.n3305 P.n3304 2.25095
R94 P.n3292 P.n3291 2.25095
R95 P.n3478 P.n2476 2.25095
R96 P.n3465 P.n3464 2.25095
R97 P.n3453 P.n2722 2.25095
R98 P.n3453 P.n2711 2.25095
R99 P.n3465 P.n2625 2.25095
R100 P.n3397 P.n2811 2.25095
R101 P.n3490 P.n2462 2.25095
R102 P.n3528 P.n3527 2.25095
R103 P.n3528 P.n2349 2.25095
R104 P.n3402 P.n2767 2.25095
R105 P.n3416 P.n3415 2.25095
R106 P.n3516 P.n2435 2.25095
R107 P.n3693 P.n3692 2.25095
R108 P.n3577 P.n2191 2.25095
R109 P.n3693 P.n2180 2.25095
R110 P.n3538 P.n2219 2.25095
R111 P.n3417 P.n2753 2.25079
R112 P.n3398 P.n2801 2.25079
R113 P.n413 P.n61 2.25079
R114 P.n426 P.n425 2.25078
R115 P.n2017 P.t12 2.2505
R116 P.n2018 P.t123 2.2505
R117 P.n2019 P.t130 2.2505
R118 P.n2020 P.t77 2.2505
R119 P.n2021 P.t46 2.2505
R120 P.n2022 P.t128 2.2505
R121 P.n2023 P.t109 2.2505
R122 P.n2024 P.t116 2.2505
R123 P.n2025 P.t62 2.2505
R124 P.n2026 P.t121 2.2505
R125 P.n2027 P.t13 2.2505
R126 P.n3106 P.t20 2.2505
R127 P.n3107 P.t126 2.2505
R128 P.n3108 P.t4 2.2505
R129 P.n3109 P.t84 2.2505
R130 P.n3110 P.t50 2.2505
R131 P.n3111 P.t3 2.2505
R132 P.n3112 P.t114 2.2505
R133 P.n3113 P.t122 2.2505
R134 P.n3114 P.t73 2.2505
R135 P.n3115 P.t30 2.2505
R136 P.n3116 P.t51 2.2505
R137 P.n2782 P.t103 2.2505
R138 P.n2783 P.t80 2.2505
R139 P.n2784 P.t92 2.2505
R140 P.n2785 P.t29 2.2505
R141 P.n2786 P.t1 2.2505
R142 P.n2787 P.t90 2.2505
R143 P.n2788 P.t56 2.2505
R144 P.n2789 P.t72 2.2505
R145 P.n2790 P.t16 2.2505
R146 P.n2791 P.t87 2.2505
R147 P.n2792 P.t9 2.2505
R148 P.n2511 P.t113 2.2505
R149 P.n2512 P.t97 2.2505
R150 P.n2513 P.t104 2.2505
R151 P.n2514 P.t40 2.2505
R152 P.n2515 P.t17 2.2505
R153 P.n2516 P.t102 2.2505
R154 P.n2517 P.t78 2.2505
R155 P.n2518 P.t91 2.2505
R156 P.n2519 P.t34 2.2505
R157 P.n2520 P.t37 2.2505
R158 P.n2521 P.t15 2.2505
R159 P.n2192 P.t71 2.2505
R160 P.n2193 P.t43 2.2505
R161 P.n2194 P.t49 2.2505
R162 P.n2195 P.t124 2.2505
R163 P.n2196 P.t107 2.2505
R164 P.n2197 P.t48 2.2505
R165 P.n2198 P.t32 2.2505
R166 P.n2199 P.t39 2.2505
R167 P.n2200 P.t117 2.2505
R168 P.n2201 P.t67 2.2505
R169 P.n2202 P.t60 2.2505
R170 P.n0 P.t105 2.2505
R171 P.n1 P.t83 2.2505
R172 P.n2 P.t95 2.2505
R173 P.n3 P.t31 2.2505
R174 P.n4 P.t5 2.2505
R175 P.n5 P.t94 2.2505
R176 P.n6 P.t61 2.2505
R177 P.n7 P.t75 2.2505
R178 P.n8 P.t19 2.2505
R179 P.n9 P.t21 2.2505
R180 P.n10 P.t57 2.2505
R181 P.n11 P.t28 2.2505
R182 P.n12 P.t0 2.2505
R183 P.n13 P.t10 2.2505
R184 P.n14 P.t93 2.2505
R185 P.n15 P.t59 2.2505
R186 P.n16 P.t8 2.2505
R187 P.n17 P.t120 2.2505
R188 P.n18 P.t125 2.2505
R189 P.n19 P.t81 2.2505
R190 P.n20 P.t2 2.2505
R191 P.n21 P.t70 2.2505
R192 P.n22 P.t106 2.2505
R193 P.n23 P.t88 2.2505
R194 P.n24 P.t98 2.2505
R195 P.n25 P.t35 2.2505
R196 P.n26 P.t7 2.2505
R197 P.n27 P.t96 2.2505
R198 P.n28 P.t65 2.2505
R199 P.n29 P.t79 2.2505
R200 P.n30 P.t25 2.2505
R201 P.n31 P.t54 2.2505
R202 P.n32 P.t23 2.2505
R203 P.n33 P.t55 2.2505
R204 P.n34 P.t38 2.2505
R205 P.n35 P.t44 2.2505
R206 P.n36 P.t118 2.2505
R207 P.n37 P.t101 2.2505
R208 P.n38 P.t42 2.2505
R209 P.n39 P.t22 2.2505
R210 P.n40 P.t33 2.2505
R211 P.n41 P.t110 2.2505
R212 P.n42 P.t99 2.2505
R213 P.n43 P.t66 2.2505
R214 P.n44 P.t85 2.2505
R215 P.n45 P.t52 2.2505
R216 P.n46 P.t68 2.2505
R217 P.n47 P.t6 2.2505
R218 P.n48 P.t115 2.2505
R219 P.n49 P.t63 2.2505
R220 P.n50 P.t41 2.2505
R221 P.n51 P.t47 2.2505
R222 P.n52 P.t127 2.2505
R223 P.n53 P.t45 2.2505
R224 P.n54 P.t111 2.2505
R225 P.n62 P.t100 2.2505
R226 P.n63 P.t76 2.2505
R227 P.n64 P.t89 2.2505
R228 P.n65 P.t26 2.2505
R229 P.n66 P.t131 2.2505
R230 P.n67 P.t86 2.2505
R231 P.n68 P.t53 2.2505
R232 P.n69 P.t69 2.2505
R233 P.n70 P.t11 2.2505
R234 P.n71 P.t58 2.2505
R235 P.n72 P.t108 2.2505
R236 P.n2857 P.n2856 1.13834
R237 P.n2291 P.n2290 1.13834
R238 P.n3628 P.n3627 1.13834
R239 P.n2570 P.n2569 1.13834
R240 P.n2999 P.n2998 1.13834
R241 P.n1903 P.n1902 1.13792
R242 P.n1465 P.n1464 1.13792
R243 P.n1150 P.n1149 1.13792
R244 P.n946 P.n945 1.13792
R245 P.n230 P.n229 1.13792
R246 P.n570 P.n569 1.13792
R247 P.n3084 P.n3083 1.1255
R248 P.n3266 P.n3265 1.1255
R249 P.n2884 P.n2883 0.9005
R250 P.n3368 P.n3367 0.9005
R251 P.n2408 P.n2407 0.9005
R252 P.n2318 P.n2317 0.9005
R253 P.n2083 P.n2082 0.9005
R254 P.n3655 P.n3654 0.9005
R255 P.n1930 P.n1929 0.9005
R256 P.n1802 P.n1801 0.9005
R257 P.n1492 P.n1491 0.9005
R258 P.n1603 P.n1602 0.9005
R259 P.n1177 P.n1176 0.9005
R260 P.n1255 P.n1254 0.9005
R261 P.n973 P.n972 0.9005
R262 P.n846 P.n845 0.9005
R263 P.n162 P.n161 0.9005
R264 P.n257 P.n256 0.9005
R265 P.n597 P.n596 0.9005
R266 P.n477 P.n476 0.9005
R267 P.n2597 P.n2596 0.9005
R268 P.n2681 P.n2680 0.9005
R269 P.n3026 P.n3025 0.9005
R270 P.n3210 P.n3209 0.9005
R271 P.n3248 P.n3235 0.9005
R272 P.n3066 P.n3052 0.9005
R273 P.n188 P.n187 0.9005
R274 P.n872 P.n871 0.9005
R275 P.n1204 P.n1203 0.9005
R276 P.n2109 P.n2108 0.9005
R277 P.n1519 P.n1518 0.9005
R278 P.n1629 P.n1628 0.9005
R279 P.n2707 P.n2706 0.9005
R280 P.n2911 P.n2910 0.9005
R281 P.n2345 P.n2344 0.9005
R282 P.n2624 P.n2623 0.9005
R283 P.n2434 P.n2433 0.9005
R284 P.n3394 P.n3393 0.9005
R285 P.n3690 P.n3681 0.9005
R286 P.n1957 P.n1956 0.9005
R287 P.n1828 P.n1827 0.9005
R288 P.n1281 P.n1280 0.9005
R289 P.n1000 P.n999 0.9005
R290 P.n284 P.n283 0.9005
R291 P.n624 P.n623 0.9005
R292 P.n503 P.n502 0.9005
R293 P.n724 P.n723 0.143661
R294 P.n2018 P.n2017 0.135964
R295 P.n2019 P.n2018 0.135964
R296 P.n2020 P.n2019 0.135964
R297 P.n2021 P.n2020 0.135964
R298 P.n2022 P.n2021 0.135964
R299 P.n2023 P.n2022 0.135964
R300 P.n2024 P.n2023 0.135964
R301 P.n2025 P.n2024 0.135964
R302 P.n2026 P.n2025 0.135964
R303 P.n2027 P.n2026 0.135964
R304 P.n3107 P.n3106 0.135964
R305 P.n3108 P.n3107 0.135964
R306 P.n3109 P.n3108 0.135964
R307 P.n3110 P.n3109 0.135964
R308 P.n3111 P.n3110 0.135964
R309 P.n3112 P.n3111 0.135964
R310 P.n3113 P.n3112 0.135964
R311 P.n3114 P.n3113 0.135964
R312 P.n3115 P.n3114 0.135964
R313 P.n3116 P.n3115 0.135964
R314 P.n2783 P.n2782 0.135964
R315 P.n2784 P.n2783 0.135964
R316 P.n2785 P.n2784 0.135964
R317 P.n2786 P.n2785 0.135964
R318 P.n2787 P.n2786 0.135964
R319 P.n2788 P.n2787 0.135964
R320 P.n2789 P.n2788 0.135964
R321 P.n2790 P.n2789 0.135964
R322 P.n2791 P.n2790 0.135964
R323 P.n2792 P.n2791 0.135964
R324 P.n2512 P.n2511 0.135964
R325 P.n2513 P.n2512 0.135964
R326 P.n2514 P.n2513 0.135964
R327 P.n2515 P.n2514 0.135964
R328 P.n2516 P.n2515 0.135964
R329 P.n2517 P.n2516 0.135964
R330 P.n2518 P.n2517 0.135964
R331 P.n2519 P.n2518 0.135964
R332 P.n2520 P.n2519 0.135964
R333 P.n2521 P.n2520 0.135964
R334 P.n2193 P.n2192 0.135964
R335 P.n2194 P.n2193 0.135964
R336 P.n2195 P.n2194 0.135964
R337 P.n2196 P.n2195 0.135964
R338 P.n2197 P.n2196 0.135964
R339 P.n2198 P.n2197 0.135964
R340 P.n2199 P.n2198 0.135964
R341 P.n2200 P.n2199 0.135964
R342 P.n2201 P.n2200 0.135964
R343 P.n2202 P.n2201 0.135964
R344 P.n1 P.n0 0.135964
R345 P.n2 P.n1 0.135964
R346 P.n3 P.n2 0.135964
R347 P.n4 P.n3 0.135964
R348 P.n5 P.n4 0.135964
R349 P.n6 P.n5 0.135964
R350 P.n7 P.n6 0.135964
R351 P.n8 P.n7 0.135964
R352 P.n9 P.n8 0.135964
R353 P.n10 P.n9 0.135964
R354 P.n12 P.n11 0.135964
R355 P.n13 P.n12 0.135964
R356 P.n14 P.n13 0.135964
R357 P.n15 P.n14 0.135964
R358 P.n16 P.n15 0.135964
R359 P.n17 P.n16 0.135964
R360 P.n18 P.n17 0.135964
R361 P.n19 P.n18 0.135964
R362 P.n20 P.n19 0.135964
R363 P.n21 P.n20 0.135964
R364 P.n23 P.n22 0.135964
R365 P.n24 P.n23 0.135964
R366 P.n25 P.n24 0.135964
R367 P.n26 P.n25 0.135964
R368 P.n27 P.n26 0.135964
R369 P.n28 P.n27 0.135964
R370 P.n29 P.n28 0.135964
R371 P.n30 P.n29 0.135964
R372 P.n31 P.n30 0.135964
R373 P.n32 P.n31 0.135964
R374 P.n34 P.n33 0.135964
R375 P.n35 P.n34 0.135964
R376 P.n36 P.n35 0.135964
R377 P.n37 P.n36 0.135964
R378 P.n38 P.n37 0.135964
R379 P.n39 P.n38 0.135964
R380 P.n40 P.n39 0.135964
R381 P.n41 P.n40 0.135964
R382 P.n42 P.n41 0.135964
R383 P.n43 P.n42 0.135964
R384 P.n45 P.n44 0.135964
R385 P.n46 P.n45 0.135964
R386 P.n47 P.n46 0.135964
R387 P.n48 P.n47 0.135964
R388 P.n49 P.n48 0.135964
R389 P.n50 P.n49 0.135964
R390 P.n51 P.n50 0.135964
R391 P.n52 P.n51 0.135964
R392 P.n53 P.n52 0.135964
R393 P.n54 P.n53 0.135964
R394 P.n63 P.n62 0.135964
R395 P.n64 P.n63 0.135964
R396 P.n65 P.n64 0.135964
R397 P.n66 P.n65 0.135964
R398 P.n67 P.n66 0.135964
R399 P.n68 P.n67 0.135964
R400 P.n69 P.n68 0.135964
R401 P.n70 P.n69 0.135964
R402 P.n71 P.n70 0.135964
R403 P.n72 P.n71 0.135964
R404 P.n3419 P.n3418 0.135597
R405 P.n1053 P.n1052 0.134522
R406 P.n1359 P.n1358 0.131145
R407 P.n1689 P.n1688 0.130758
R408 P.n3544 P.n3543 0.128242
R409 P.n3481 P.n3480 0.124113
R410 P.n400 P.n399 0.106366
R411 P.n3284 P.n3283 0.0959839
R412 P P.n2016 0.0776398
R413 P P.n3708 0.0578978
R414 P.n222 P.n221 0.0558778
R415 P.n938 P.n937 0.0523449
R416 P.n562 P.n561 0.0512851
R417 P.n2283 P.n2282 0.0492919
R418 P.n2849 P.n2848 0.0445406
R419 P.n1895 P.n1894 0.044131
R420 P.n2562 P.n2561 0.0432614
R421 P.n1142 P.n1141 0.0410397
R422 P.n3620 P.n3619 0.0407944
R423 P.n1457 P.n1456 0.03892
R424 P.n2991 P.n2990 0.0388756
R425 P.n3117 P.n3116 0.0376056
R426 P.n3468 P.n2521 0.0354299
R427 P.n3707 P.n2027 0.0340142
R428 P.n3401 P.n2792 0.0340142
R429 P.n3543 P.n2202 0.0340142
R430 P.n1689 P.n10 0.0340142
R431 P.n1365 P.n21 0.0340142
R432 P.n1060 P.n32 0.0340142
R433 P.n741 P.n43 0.0340142
R434 P.n417 P.n54 0.0340142
R435 P.n104 P.n72 0.0340142
R436 P.n2853 P.n2852 0.0140228
R437 P.n2843 P.n2842 0.0140228
R438 P.n2287 P.n2286 0.0140228
R439 P.n2277 P.n2276 0.0140228
R440 P.n3624 P.n3623 0.0140228
R441 P.n3614 P.n3613 0.0140228
R442 P.n2566 P.n2565 0.0140228
R443 P.n2556 P.n2555 0.0140228
R444 P.n2995 P.n2994 0.0140228
R445 P.n2985 P.n2984 0.0140228
R446 P.n1899 P.n1898 0.0135716
R447 P.n1889 P.n1888 0.0135716
R448 P.n1461 P.n1460 0.0135716
R449 P.n1451 P.n1450 0.0135716
R450 P.n1146 P.n1145 0.0135716
R451 P.n1136 P.n1135 0.0135716
R452 P.n942 P.n941 0.0135716
R453 P.n932 P.n931 0.0135716
R454 P.n226 P.n225 0.0135716
R455 P.n216 P.n215 0.0135716
R456 P.n566 P.n565 0.0135716
R457 P.n556 P.n555 0.0135716
R458 P.n2847 P.n2846 0.012835
R459 P.n2281 P.n2280 0.012835
R460 P.n3618 P.n3617 0.012835
R461 P.n2560 P.n2559 0.012835
R462 P.n2989 P.n2988 0.012835
R463 P.n1893 P.n1892 0.0124235
R464 P.n1455 P.n1454 0.0124235
R465 P.n1140 P.n1139 0.0124235
R466 P.n936 P.n935 0.0124235
R467 P.n220 P.n219 0.0124235
R468 P.n560 P.n559 0.0124235
R469 P.n2878 P.n2877 0.00790102
R470 P.n3362 P.n3361 0.00790102
R471 P.n2312 P.n2311 0.00790102
R472 P.n2402 P.n2401 0.00790102
R473 P.n3649 P.n3648 0.00790102
R474 P.n2077 P.n2076 0.00790102
R475 P.n2591 P.n2590 0.00790102
R476 P.n2675 P.n2674 0.00790102
R477 P.n3020 P.n3019 0.00790102
R478 P.n3204 P.n3203 0.00790102
R479 P.n1924 P.n1923 0.00765407
R480 P.n1796 P.n1795 0.00765407
R481 P.n1486 P.n1485 0.00765407
R482 P.n1597 P.n1596 0.00765407
R483 P.n1171 P.n1170 0.00765407
R484 P.n1249 P.n1248 0.00765407
R485 P.n967 P.n966 0.00765407
R486 P.n840 P.n839 0.00765407
R487 P.n251 P.n250 0.00765407
R488 P.n156 P.n155 0.00765407
R489 P.n591 P.n590 0.00765407
R490 P.n471 P.n470 0.00765407
R491 P.n2894 P.n2893 0.00717005
R492 P.n3378 P.n3377 0.00717005
R493 P.n2328 P.n2327 0.00717005
R494 P.n2418 P.n2417 0.00717005
R495 P.n3665 P.n3664 0.00717005
R496 P.n2093 P.n2092 0.00717005
R497 P.n2607 P.n2606 0.00717005
R498 P.n2691 P.n2690 0.00717005
R499 P.n3036 P.n3035 0.00717005
R500 P.n3220 P.n3219 0.00717005
R501 P.n1940 P.n1939 0.0069475
R502 P.n1812 P.n1811 0.0069475
R503 P.n1502 P.n1501 0.0069475
R504 P.n1613 P.n1612 0.0069475
R505 P.n1187 P.n1186 0.0069475
R506 P.n1265 P.n1264 0.0069475
R507 P.n983 P.n982 0.0069475
R508 P.n856 P.n855 0.0069475
R509 P.n267 P.n266 0.0069475
R510 P.n172 P.n171 0.0069475
R511 P.n607 P.n606 0.0069475
R512 P.n487 P.n486 0.0069475
R513 P.n2861 P.n2860 0.0067132
R514 P.n3346 P.n3345 0.0067132
R515 P.n2295 P.n2294 0.0067132
R516 P.n2386 P.n2385 0.0067132
R517 P.n3632 P.n3631 0.0067132
R518 P.n2061 P.n2060 0.0067132
R519 P.n2574 P.n2573 0.0067132
R520 P.n2659 P.n2658 0.0067132
R521 P.n3003 P.n3002 0.0067132
R522 P.n3188 P.n3187 0.0067132
R523 P.n1907 P.n1906 0.00650589
R524 P.n1780 P.n1779 0.00650589
R525 P.n1469 P.n1468 0.00650589
R526 P.n1581 P.n1580 0.00650589
R527 P.n1154 P.n1153 0.00650589
R528 P.n1233 P.n1232 0.00650589
R529 P.n950 P.n949 0.00650589
R530 P.n824 P.n823 0.00650589
R531 P.n234 P.n233 0.00650589
R532 P.n140 P.n139 0.00650589
R533 P.n574 P.n573 0.00650589
R534 P.n455 P.n454 0.00650589
R535 P.n3283 P.n3282 0.0065
R536 P.n3075 P.n3074 0.00616497
R537 P.n3257 P.n3256 0.00616497
R538 P.n2829 P.n2828 0.00598223
R539 P.n3331 P.n3330 0.00598223
R540 P.n2263 P.n2262 0.00598223
R541 P.n2371 P.n2370 0.00598223
R542 P.n3600 P.n3599 0.00598223
R543 P.n2046 P.n2045 0.00598223
R544 P.n2542 P.n2541 0.00598223
R545 P.n2644 P.n2643 0.00598223
R546 P.n2971 P.n2970 0.00598223
R547 P.n3173 P.n3172 0.00598223
R548 P.n1875 P.n1874 0.00579931
R549 P.n1765 P.n1764 0.00579931
R550 P.n1437 P.n1436 0.00579931
R551 P.n1566 P.n1565 0.00579931
R552 P.n1122 P.n1121 0.00579931
R553 P.n1218 P.n1217 0.00579931
R554 P.n918 P.n917 0.00579931
R555 P.n809 P.n808 0.00579931
R556 P.n202 P.n201 0.00579931
R557 P.n125 P.n124 0.00579931
R558 P.n542 P.n541 0.00579931
R559 P.n440 P.n439 0.00579931
R560 P.n2806 P.n2805 0.00497716
R561 P.n2794 P.n2793 0.00497716
R562 P.n3522 P.n3521 0.00497716
R563 P.n2437 P.n2436 0.00497716
R564 P.n2172 P.n2171 0.00497716
R565 P.n2165 P.n2164 0.00497716
R566 P.n3455 P.n3454 0.00497716
R567 P.n2717 P.n2716 0.00497716
R568 P.n2949 P.n2948 0.00497716
R569 P.n3150 P.n3149 0.00497716
R570 P.n2856 P.n2855 0.0036066
R571 P.n2846 P.n2845 0.0036066
R572 P.n2290 P.n2289 0.0036066
R573 P.n2280 P.n2279 0.0036066
R574 P.n3627 P.n3626 0.0036066
R575 P.n3617 P.n3616 0.0036066
R576 P.n2569 P.n2568 0.0036066
R577 P.n2559 P.n2558 0.0036066
R578 P.n2998 P.n2997 0.0036066
R579 P.n2988 P.n2987 0.0036066
R580 P.n2862 P.n2861 0.00351523
R581 P.n3347 P.n3346 0.00351523
R582 P.n2296 P.n2295 0.00351523
R583 P.n2387 P.n2386 0.00351523
R584 P.n3633 P.n3632 0.00351523
R585 P.n2062 P.n2061 0.00351523
R586 P.n2575 P.n2574 0.00351523
R587 P.n2660 P.n2659 0.00351523
R588 P.n3004 P.n3003 0.00351523
R589 P.n3189 P.n3188 0.00351523
R590 P.n1902 P.n1901 0.00350294
R591 P.n1892 P.n1891 0.00350294
R592 P.n1464 P.n1463 0.00350294
R593 P.n1454 P.n1453 0.00350294
R594 P.n1149 P.n1148 0.00350294
R595 P.n1139 P.n1138 0.00350294
R596 P.n945 P.n944 0.00350294
R597 P.n935 P.n934 0.00350294
R598 P.n229 P.n228 0.00350294
R599 P.n219 P.n218 0.00350294
R600 P.n569 P.n568 0.00350294
R601 P.n559 P.n558 0.00350294
R602 P.n1066 P.n1065 0.00346774
R603 P.n3312 P.n3311 0.00346774
R604 P.n1908 P.n1907 0.00341462
R605 P.n1781 P.n1780 0.00341462
R606 P.n1470 P.n1469 0.00341462
R607 P.n1582 P.n1581 0.00341462
R608 P.n1155 P.n1154 0.00341462
R609 P.n1234 P.n1233 0.00341462
R610 P.n951 P.n950 0.00341462
R611 P.n825 P.n824 0.00341462
R612 P.n235 P.n234 0.00341462
R613 P.n141 P.n140 0.00341462
R614 P.n575 P.n574 0.00341462
R615 P.n456 P.n455 0.00341462
R616 P.n2831 P.n2830 0.00324112
R617 P.n3333 P.n3332 0.00324112
R618 P.n2265 P.n2264 0.00324112
R619 P.n2373 P.n2372 0.00324112
R620 P.n3602 P.n3601 0.00324112
R621 P.n2048 P.n2047 0.00324112
R622 P.n2544 P.n2543 0.00324112
R623 P.n2646 P.n2645 0.00324112
R624 P.n2973 P.n2972 0.00324112
R625 P.n3175 P.n3174 0.00324112
R626 P.n1378 P.n1377 0.00323118
R627 P.n3589 P.n3588 0.00323118
R628 P.n1877 P.n1876 0.00314966
R629 P.n1767 P.n1766 0.00314966
R630 P.n1439 P.n1438 0.00314966
R631 P.n1568 P.n1567 0.00314966
R632 P.n1124 P.n1123 0.00314966
R633 P.n1220 P.n1219 0.00314966
R634 P.n920 P.n919 0.00314966
R635 P.n811 P.n810 0.00314966
R636 P.n204 P.n203 0.00314966
R637 P.n127 P.n126 0.00314966
R638 P.n544 P.n543 0.00314966
R639 P.n442 P.n441 0.00314966
R640 P.n1708 P.n1707 0.00310215
R641 P.n3415 P.n3414 0.00310152
R642 P.n2132 P.n2123 0.00310152
R643 P.n2121 P.n2113 0.00310152
R644 P.n3451 P.n3450 0.00303763
R645 P.n1969 P.n1968 0.0030314
R646 P.n1839 P.n1838 0.0030314
R647 P.n1419 P.n1418 0.0030314
R648 P.n1640 P.n1639 0.0030314
R649 P.n1292 P.n1291 0.0030314
R650 P.n1012 P.n1011 0.0030314
R651 P.n798 P.n797 0.0030314
R652 P.n366 P.n365 0.0030314
R653 P.n693 P.n692 0.0030314
R654 P.n743 P.n742 0.00297312
R655 P.n2808 P.n2807 0.00296701
R656 P.n2796 P.n2795 0.00296701
R657 P.n3524 P.n3523 0.00296701
R658 P.n2439 P.n2438 0.00296701
R659 P.n2174 P.n2173 0.00296701
R660 P.n2167 P.n2166 0.00296701
R661 P.n3457 P.n3456 0.00296701
R662 P.n2719 P.n2718 0.00296701
R663 P.n2951 P.n2950 0.00296701
R664 P.n3152 P.n3151 0.00296701
R665 P.n1982 P.n1981 0.00288469
R666 P.n1853 P.n1852 0.00288469
R667 P.n1535 P.n1534 0.00288469
R668 P.n1654 P.n1653 0.00288469
R669 P.n1319 P.n1318 0.00288469
R670 P.n1306 P.n1305 0.00288469
R671 P.n1026 P.n1025 0.00288469
R672 P.n888 P.n887 0.00288469
R673 P.n96 P.n95 0.00288469
R674 P.n88 P.n87 0.00288469
R675 P.n421 P.n420 0.00288469
R676 P.n57 P.n56 0.00288469
R677 P.n3514 P.n3513 0.00284409
R678 P.n3304 P.n3302 0.00282741
R679 P.n2919 P.n2917 0.00282741
R680 P.n2451 P.n2450 0.00282741
R681 P.n2457 P.n2455 0.00282741
R682 P.n3574 P.n3567 0.00282741
R683 P.n2191 P.n2184 0.00282741
R684 P.n2732 P.n2731 0.00282741
R685 P.n2743 P.n2742 0.00282741
R686 P.n3400 P.n3399 0.00282258
R687 P.n1744 P.n1742 0.00276644
R688 P.n1737 P.n1736 0.00276644
R689 P.n1392 P.n1391 0.00276644
R690 P.n1399 P.n1398 0.00276644
R691 P.n1088 P.n1087 0.00276644
R692 P.n1084 P.n1083 0.00276644
R693 P.n780 P.n779 0.00276644
R694 P.n773 P.n772 0.00276644
R695 P.n308 P.n307 0.00276644
R696 P.n301 P.n300 0.00276644
R697 P.n635 P.n633 0.00276644
R698 P.n522 P.n520 0.00276644
R699 P.n2767 P.n2766 0.00273604
R700 P.n2781 P.n2780 0.00273604
R701 P.n2232 P.n2231 0.00273604
R702 P.n2245 P.n2244 0.00273604
R703 P.n2160 P.n2152 0.00273604
R704 P.n2146 P.n2138 0.00273604
R705 P.n2497 P.n2489 0.00273604
R706 P.n2510 P.n2502 0.00273604
R707 P.n2850 P.n2849 0.00269289
R708 P.n2867 P.n2866 0.00269289
R709 P.n2284 P.n2283 0.00269289
R710 P.n2301 P.n2300 0.00269289
R711 P.n3621 P.n3620 0.00269289
R712 P.n3638 P.n3637 0.00269289
R713 P.n2563 P.n2562 0.00269289
R714 P.n2580 P.n2579 0.00269289
R715 P.n2992 P.n2991 0.00269289
R716 P.n3009 P.n3008 0.00269289
R717 P.n2001 P.n2000 0.00267811
R718 P.n1850 P.n1849 0.00267811
R719 P.n1532 P.n1531 0.00267811
R720 P.n1651 P.n1650 0.00267811
R721 P.n1338 P.n1337 0.00267811
R722 P.n1303 P.n1302 0.00267811
R723 P.n1023 P.n1022 0.00267811
R724 P.n885 P.n884 0.00267811
R725 P.n383 P.n382 0.00267811
R726 P.n338 P.n337 0.00267811
R727 P.n663 P.n662 0.00267811
R728 P.n1896 P.n1895 0.00261973
R729 P.n1913 P.n1912 0.00261973
R730 P.n1458 P.n1457 0.00261973
R731 P.n1475 P.n1474 0.00261973
R732 P.n1143 P.n1142 0.00261973
R733 P.n1160 P.n1159 0.00261973
R734 P.n939 P.n938 0.00261973
R735 P.n956 P.n955 0.00261973
R736 P.n223 P.n222 0.00261973
R737 P.n240 P.n239 0.00261973
R738 P.n563 P.n562 0.00261973
R739 P.n580 P.n579 0.00261973
R740 P.n1372 P.n1371 0.00258602
R741 P.n3697 P.n3696 0.00258602
R742 P.n3290 P.n3289 0.00251015
R743 P.n2923 P.n2922 0.00251015
R744 P.n2746 P.n2745 0.00251015
R745 P.n2461 P.n2460 0.00251015
R746 P.n2466 P.n2465 0.00251015
R747 P.n3571 P.n3570 0.00251015
R748 P.n2188 P.n2187 0.00251015
R749 P.n2726 P.n2725 0.00251015
R750 P.n2736 P.n2735 0.00251015
R751 P.n2945 P.n2944 0.00251015
R752 P.n3062 P.n3061 0.00251015
R753 P.n3146 P.n3145 0.00251015
R754 P.n3244 P.n3243 0.00251015
R755 P.n1702 P.n1701 0.00245699
R756 P.n2008 P.n2007 0.00244308
R757 P.n1977 P.n1976 0.00244308
R758 P.n1672 P.n1671 0.00244308
R759 P.n1680 P.n1679 0.00244308
R760 P.n1353 P.n1352 0.00244308
R761 P.n1104 P.n1103 0.00244308
R762 P.n1346 P.n1345 0.00244308
R763 P.n1045 P.n1044 0.00244308
R764 P.n905 P.n904 0.00244308
R765 P.n392 P.n391 0.00244308
R766 P.n352 P.n351 0.00244308
R767 P.n327 P.n326 0.00244308
R768 P.n718 P.n717 0.00244308
R769 P.n675 P.n674 0.00244308
R770 P.n652 P.n651 0.00244308
R771 P.n2871 P.n2870 0.00241878
R772 P.n3355 P.n3354 0.00241878
R773 P.n2907 P.n2906 0.00241878
R774 P.n3390 P.n3389 0.00241878
R775 P.n2305 P.n2304 0.00241878
R776 P.n2395 P.n2394 0.00241878
R777 P.n2341 P.n2340 0.00241878
R778 P.n2430 P.n2429 0.00241878
R779 P.n3642 P.n3641 0.00241878
R780 P.n2070 P.n2069 0.00241878
R781 P.n3678 P.n3677 0.00241878
R782 P.n2105 P.n2104 0.00241878
R783 P.n2584 P.n2583 0.00241878
R784 P.n2668 P.n2667 0.00241878
R785 P.n2620 P.n2619 0.00241878
R786 P.n2703 P.n2702 0.00241878
R787 P.n3013 P.n3012 0.00241878
R788 P.n3197 P.n3196 0.00241878
R789 P.n3049 P.n3048 0.00241878
R790 P.n3232 P.n3231 0.00241878
R791 P.n1092 P.n1091 0.00241398
R792 P.n3298 P.n3297 0.00241398
R793 P.n3573 P.n3572 0.00237056
R794 P.n2190 P.n2189 0.00237056
R795 P.n2728 P.n2727 0.00237056
R796 P.n2738 P.n2737 0.00237056
R797 P.n1917 P.n1916 0.00235476
R798 P.n1789 P.n1788 0.00235476
R799 P.n1953 P.n1952 0.00235476
R800 P.n1824 P.n1823 0.00235476
R801 P.n1479 P.n1478 0.00235476
R802 P.n1590 P.n1589 0.00235476
R803 P.n1515 P.n1514 0.00235476
R804 P.n1625 P.n1624 0.00235476
R805 P.n1164 P.n1163 0.00235476
R806 P.n1242 P.n1241 0.00235476
R807 P.n1200 P.n1199 0.00235476
R808 P.n1277 P.n1276 0.00235476
R809 P.n960 P.n959 0.00235476
R810 P.n833 P.n832 0.00235476
R811 P.n996 P.n995 0.00235476
R812 P.n868 P.n867 0.00235476
R813 P.n244 P.n243 0.00235476
R814 P.n149 P.n148 0.00235476
R815 P.n280 P.n279 0.00235476
R816 P.n184 P.n183 0.00235476
R817 P.n584 P.n583 0.00235476
R818 P.n464 P.n463 0.00235476
R819 P.n620 P.n619 0.00235476
R820 P.n499 P.n498 0.00235476
R821 P.n736 P.n735 0.00232796
R822 P.n2854 P.n2853 0.00232741
R823 P.n2844 P.n2843 0.00232741
R824 P.n2865 P.n2864 0.00232741
R825 P.n2882 P.n2881 0.00232741
R826 P.n2879 P.n2878 0.00232741
R827 P.n2875 P.n2874 0.00232741
R828 P.n3350 P.n3349 0.00232741
R829 P.n3366 P.n3365 0.00232741
R830 P.n3363 P.n3362 0.00232741
R831 P.n3359 P.n3358 0.00232741
R832 P.n2887 P.n2886 0.00232741
R833 P.n2910 P.n2898 0.00232741
R834 P.n2901 P.n2900 0.00232741
R835 P.n3371 P.n3370 0.00232741
R836 P.n3393 P.n3382 0.00232741
R837 P.n3384 P.n3383 0.00232741
R838 P.n3407 P.n3406 0.00232741
R839 P.n2748 P.n2747 0.00232741
R840 P.n2288 P.n2287 0.00232741
R841 P.n2278 P.n2277 0.00232741
R842 P.n2299 P.n2298 0.00232741
R843 P.n2316 P.n2315 0.00232741
R844 P.n2313 P.n2312 0.00232741
R845 P.n2309 P.n2308 0.00232741
R846 P.n2390 P.n2389 0.00232741
R847 P.n2406 P.n2405 0.00232741
R848 P.n2403 P.n2402 0.00232741
R849 P.n2399 P.n2398 0.00232741
R850 P.n2321 P.n2320 0.00232741
R851 P.n2344 P.n2332 0.00232741
R852 P.n2335 P.n2334 0.00232741
R853 P.n2411 P.n2410 0.00232741
R854 P.n2433 P.n2422 0.00232741
R855 P.n2424 P.n2423 0.00232741
R856 P.n2205 P.n2204 0.00232741
R857 P.n2213 P.n2212 0.00232741
R858 P.n3625 P.n3624 0.00232741
R859 P.n3615 P.n3614 0.00232741
R860 P.n3636 P.n3635 0.00232741
R861 P.n3653 P.n3652 0.00232741
R862 P.n3650 P.n3649 0.00232741
R863 P.n3646 P.n3645 0.00232741
R864 P.n2065 P.n2064 0.00232741
R865 P.n2081 P.n2080 0.00232741
R866 P.n2078 P.n2077 0.00232741
R867 P.n2074 P.n2073 0.00232741
R868 P.n3658 P.n3657 0.00232741
R869 P.n3681 P.n3669 0.00232741
R870 P.n3672 P.n3671 0.00232741
R871 P.n2086 P.n2085 0.00232741
R872 P.n2108 P.n2097 0.00232741
R873 P.n2099 P.n2098 0.00232741
R874 P.n2126 P.n2125 0.00232741
R875 P.n2115 P.n2114 0.00232741
R876 P.n2567 P.n2566 0.00232741
R877 P.n2557 P.n2556 0.00232741
R878 P.n2578 P.n2577 0.00232741
R879 P.n2595 P.n2594 0.00232741
R880 P.n2592 P.n2591 0.00232741
R881 P.n2588 P.n2587 0.00232741
R882 P.n2663 P.n2662 0.00232741
R883 P.n2679 P.n2678 0.00232741
R884 P.n2676 P.n2675 0.00232741
R885 P.n2672 P.n2671 0.00232741
R886 P.n2600 P.n2599 0.00232741
R887 P.n2623 P.n2611 0.00232741
R888 P.n2614 P.n2613 0.00232741
R889 P.n2684 P.n2683 0.00232741
R890 P.n2706 P.n2695 0.00232741
R891 P.n2697 P.n2696 0.00232741
R892 P.n2470 P.n2469 0.00232741
R893 P.n2478 P.n2477 0.00232741
R894 P.n2996 P.n2995 0.00232741
R895 P.n2986 P.n2985 0.00232741
R896 P.n3007 P.n3006 0.00232741
R897 P.n3024 P.n3023 0.00232741
R898 P.n3021 P.n3020 0.00232741
R899 P.n3017 P.n3016 0.00232741
R900 P.n3192 P.n3191 0.00232741
R901 P.n3208 P.n3207 0.00232741
R902 P.n3205 P.n3204 0.00232741
R903 P.n3201 P.n3200 0.00232741
R904 P.n3029 P.n3028 0.00232741
R905 P.n3052 P.n3040 0.00232741
R906 P.n3043 P.n3042 0.00232741
R907 P.n3213 P.n3212 0.00232741
R908 P.n3235 P.n3224 0.00232741
R909 P.n3226 P.n3225 0.00232741
R910 P.n3055 P.n3054 0.00232741
R911 P.n3237 P.n3236 0.00232741
R912 P.n1978 P.n1972 0.00232483
R913 P.n1673 P.n1667 0.00232483
R914 P.n1681 P.n1675 0.00232483
R915 P.n1354 P.n1348 0.00232483
R916 P.n1347 P.n1341 0.00232483
R917 P.n1046 P.n1040 0.00232483
R918 P.n907 P.n906 0.00232483
R919 P.n394 P.n393 0.00232483
R920 P.n1900 P.n1899 0.00226644
R921 P.n1890 P.n1889 0.00226644
R922 P.n1911 P.n1910 0.00226644
R923 P.n1928 P.n1927 0.00226644
R924 P.n1925 P.n1924 0.00226644
R925 P.n1921 P.n1920 0.00226644
R926 P.n1784 P.n1783 0.00226644
R927 P.n1800 P.n1799 0.00226644
R928 P.n1797 P.n1796 0.00226644
R929 P.n1793 P.n1792 0.00226644
R930 P.n1933 P.n1932 0.00226644
R931 P.n1956 P.n1944 0.00226644
R932 P.n1947 P.n1946 0.00226644
R933 P.n1805 P.n1804 0.00226644
R934 P.n1827 P.n1816 0.00226644
R935 P.n1818 P.n1817 0.00226644
R936 P.n1962 P.n1961 0.00226644
R937 P.n1832 P.n1831 0.00226644
R938 P.n1462 P.n1461 0.00226644
R939 P.n1452 P.n1451 0.00226644
R940 P.n1473 P.n1472 0.00226644
R941 P.n1490 P.n1489 0.00226644
R942 P.n1487 P.n1486 0.00226644
R943 P.n1483 P.n1482 0.00226644
R944 P.n1585 P.n1584 0.00226644
R945 P.n1601 P.n1600 0.00226644
R946 P.n1598 P.n1597 0.00226644
R947 P.n1594 P.n1593 0.00226644
R948 P.n1495 P.n1494 0.00226644
R949 P.n1518 P.n1506 0.00226644
R950 P.n1509 P.n1508 0.00226644
R951 P.n1606 P.n1605 0.00226644
R952 P.n1628 P.n1617 0.00226644
R953 P.n1619 P.n1618 0.00226644
R954 P.n1412 P.n1411 0.00226644
R955 P.n1633 P.n1632 0.00226644
R956 P.n1147 P.n1146 0.00226644
R957 P.n1137 P.n1136 0.00226644
R958 P.n1158 P.n1157 0.00226644
R959 P.n1175 P.n1174 0.00226644
R960 P.n1172 P.n1171 0.00226644
R961 P.n1168 P.n1167 0.00226644
R962 P.n1237 P.n1236 0.00226644
R963 P.n1253 P.n1252 0.00226644
R964 P.n1250 P.n1249 0.00226644
R965 P.n1246 P.n1245 0.00226644
R966 P.n1180 P.n1179 0.00226644
R967 P.n1203 P.n1191 0.00226644
R968 P.n1194 P.n1193 0.00226644
R969 P.n1258 P.n1257 0.00226644
R970 P.n1280 P.n1269 0.00226644
R971 P.n1271 P.n1270 0.00226644
R972 P.n1097 P.n1096 0.00226644
R973 P.n1285 P.n1284 0.00226644
R974 P.n943 P.n942 0.00226644
R975 P.n933 P.n932 0.00226644
R976 P.n954 P.n953 0.00226644
R977 P.n971 P.n970 0.00226644
R978 P.n968 P.n967 0.00226644
R979 P.n964 P.n963 0.00226644
R980 P.n828 P.n827 0.00226644
R981 P.n844 P.n843 0.00226644
R982 P.n841 P.n840 0.00226644
R983 P.n837 P.n836 0.00226644
R984 P.n976 P.n975 0.00226644
R985 P.n999 P.n987 0.00226644
R986 P.n990 P.n989 0.00226644
R987 P.n849 P.n848 0.00226644
R988 P.n871 P.n860 0.00226644
R989 P.n862 P.n861 0.00226644
R990 P.n1005 P.n1004 0.00226644
R991 P.n791 P.n790 0.00226644
R992 P.n227 P.n226 0.00226644
R993 P.n217 P.n216 0.00226644
R994 P.n238 P.n237 0.00226644
R995 P.n255 P.n254 0.00226644
R996 P.n252 P.n251 0.00226644
R997 P.n248 P.n247 0.00226644
R998 P.n144 P.n143 0.00226644
R999 P.n160 P.n159 0.00226644
R1000 P.n157 P.n156 0.00226644
R1001 P.n153 P.n152 0.00226644
R1002 P.n260 P.n259 0.00226644
R1003 P.n283 P.n271 0.00226644
R1004 P.n274 P.n273 0.00226644
R1005 P.n165 P.n164 0.00226644
R1006 P.n187 P.n176 0.00226644
R1007 P.n178 P.n177 0.00226644
R1008 P.n359 P.n358 0.00226644
R1009 P.n320 P.n319 0.00226644
R1010 P.n567 P.n566 0.00226644
R1011 P.n557 P.n556 0.00226644
R1012 P.n578 P.n577 0.00226644
R1013 P.n595 P.n594 0.00226644
R1014 P.n592 P.n591 0.00226644
R1015 P.n588 P.n587 0.00226644
R1016 P.n459 P.n458 0.00226644
R1017 P.n475 P.n474 0.00226644
R1018 P.n472 P.n471 0.00226644
R1019 P.n468 P.n467 0.00226644
R1020 P.n600 P.n599 0.00226644
R1021 P.n623 P.n611 0.00226644
R1022 P.n614 P.n613 0.00226644
R1023 P.n480 P.n479 0.00226644
R1024 P.n502 P.n491 0.00226644
R1025 P.n493 P.n492 0.00226644
R1026 P.n686 P.n685 0.00226644
R1027 P.n645 P.n644 0.00226644
R1028 P.n412 P.n411 0.00224727
R1029 P.n2941 P.n2940 0.00223604
R1030 P.n3142 P.n3141 0.00223604
R1031 P.n84 P.n83 0.00219892
R1032 P.n3531 P.n3530 0.00219892
R1033 P.n1404 P.n1403 0.00217742
R1034 P.n3562 P.n3561 0.00217742
R1035 P.n2859 P.n2858 0.00214467
R1036 P.n3344 P.n3343 0.00214467
R1037 P.n2825 P.n2824 0.00214467
R1038 P.n3327 P.n3326 0.00214467
R1039 P.n2293 P.n2292 0.00214467
R1040 P.n2384 P.n2383 0.00214467
R1041 P.n2259 P.n2258 0.00214467
R1042 P.n2367 P.n2366 0.00214467
R1043 P.n3630 P.n3629 0.00214467
R1044 P.n2059 P.n2058 0.00214467
R1045 P.n3596 P.n3595 0.00214467
R1046 P.n2042 P.n2041 0.00214467
R1047 P.n2572 P.n2571 0.00214467
R1048 P.n2657 P.n2656 0.00214467
R1049 P.n2538 P.n2537 0.00214467
R1050 P.n2640 P.n2639 0.00214467
R1051 P.n3001 P.n3000 0.00214467
R1052 P.n3186 P.n3185 0.00214467
R1053 P.n2967 P.n2966 0.00214467
R1054 P.n3169 P.n3168 0.00214467
R1055 P.n3083 P.n3082 0.00214467
R1056 P.n3265 P.n3264 0.00214467
R1057 P.n1905 P.n1904 0.00208979
R1058 P.n1778 P.n1777 0.00208979
R1059 P.n1871 P.n1870 0.00208979
R1060 P.n1761 P.n1760 0.00208979
R1061 P.n1467 P.n1466 0.00208979
R1062 P.n1579 P.n1578 0.00208979
R1063 P.n1433 P.n1432 0.00208979
R1064 P.n1562 P.n1561 0.00208979
R1065 P.n1152 P.n1151 0.00208979
R1066 P.n1231 P.n1230 0.00208979
R1067 P.n1118 P.n1117 0.00208979
R1068 P.n1214 P.n1213 0.00208979
R1069 P.n948 P.n947 0.00208979
R1070 P.n822 P.n821 0.00208979
R1071 P.n914 P.n913 0.00208979
R1072 P.n805 P.n804 0.00208979
R1073 P.n232 P.n231 0.00208979
R1074 P.n138 P.n137 0.00208979
R1075 P.n198 P.n197 0.00208979
R1076 P.n121 P.n120 0.00208979
R1077 P.n572 P.n571 0.00208979
R1078 P.n453 P.n452 0.00208979
R1079 P.n538 P.n537 0.00208979
R1080 P.n436 P.n435 0.00208979
R1081 P.n711 P.n710 0.00208979
R1082 P.n2839 P.n2838 0.0020533
R1083 P.n3342 P.n3341 0.0020533
R1084 P.n2823 P.n2822 0.0020533
R1085 P.n3325 P.n3324 0.0020533
R1086 P.n2818 P.n2817 0.0020533
R1087 P.n3319 P.n3318 0.0020533
R1088 P.n2273 P.n2272 0.0020533
R1089 P.n2382 P.n2381 0.0020533
R1090 P.n2257 P.n2256 0.0020533
R1091 P.n2365 P.n2364 0.0020533
R1092 P.n2252 P.n2251 0.0020533
R1093 P.n2359 P.n2358 0.0020533
R1094 P.n3610 P.n3609 0.0020533
R1095 P.n2057 P.n2056 0.0020533
R1096 P.n3594 P.n3593 0.0020533
R1097 P.n2040 P.n2039 0.0020533
R1098 P.n3688 P.n3687 0.0020533
R1099 P.n2034 P.n2033 0.0020533
R1100 P.n2552 P.n2551 0.0020533
R1101 P.n2655 P.n2654 0.0020533
R1102 P.n2536 P.n2535 0.0020533
R1103 P.n2638 P.n2637 0.0020533
R1104 P.n2531 P.n2530 0.0020533
R1105 P.n2632 P.n2631 0.0020533
R1106 P.n2981 P.n2980 0.0020533
R1107 P.n3184 P.n3183 0.0020533
R1108 P.n2965 P.n2964 0.0020533
R1109 P.n3167 P.n3166 0.0020533
R1110 P.n3069 P.n3068 0.0020533
R1111 P.n3251 P.n3250 0.0020533
R1112 P.n2940 P.n2939 0.00205068
R1113 P.n1749 P.n1748 0.00204839
R1114 P.n3469 P.n3468 0.00200538
R1115 P.n1885 P.n1884 0.00200147
R1116 P.n1776 P.n1775 0.00200147
R1117 P.n1869 P.n1868 0.00200147
R1118 P.n1759 P.n1758 0.00200147
R1119 P.n1727 P.n1726 0.00200147
R1120 P.n1717 P.n1716 0.00200147
R1121 P.n1447 P.n1446 0.00200147
R1122 P.n1577 P.n1576 0.00200147
R1123 P.n1431 P.n1430 0.00200147
R1124 P.n1560 P.n1559 0.00200147
R1125 P.n1426 P.n1425 0.00200147
R1126 P.n1554 P.n1553 0.00200147
R1127 P.n1132 P.n1131 0.00200147
R1128 P.n1229 P.n1228 0.00200147
R1129 P.n1116 P.n1115 0.00200147
R1130 P.n1212 P.n1211 0.00200147
R1131 P.n1111 P.n1110 0.00200147
R1132 P.n1074 P.n1073 0.00200147
R1133 P.n928 P.n927 0.00200147
R1134 P.n820 P.n819 0.00200147
R1135 P.n912 P.n911 0.00200147
R1136 P.n803 P.n802 0.00200147
R1137 P.n764 P.n763 0.00200147
R1138 P.n752 P.n751 0.00200147
R1139 P.n212 P.n211 0.00200147
R1140 P.n136 P.n135 0.00200147
R1141 P.n196 P.n195 0.00200147
R1142 P.n119 P.n118 0.00200147
R1143 P.n291 P.n290 0.00200147
R1144 P.n114 P.n113 0.00200147
R1145 P.n552 P.n551 0.00200147
R1146 P.n451 P.n450 0.00200147
R1147 P.n536 P.n535 0.00200147
R1148 P.n434 P.n433 0.00200147
R1149 P.n532 P.n531 0.00200147
R1150 P.n510 P.n509 0.00200147
R1151 P.n3433 P.n3432 0.00198387
R1152 P.n428 P.n427 0.00196237
R1153 P.n2848 P.n2847 0.00196193
R1154 P.n2860 P.n2859 0.00196193
R1155 P.n3341 P.n3340 0.00196193
R1156 P.n3343 P.n3342 0.00196193
R1157 P.n3345 P.n3344 0.00196193
R1158 P.n2824 P.n2823 0.00196193
R1159 P.n2836 P.n2835 0.00196193
R1160 P.n2892 P.n2891 0.00196193
R1161 P.n3326 P.n3325 0.00196193
R1162 P.n3338 P.n3337 0.00196193
R1163 P.n3376 P.n3375 0.00196193
R1164 P.n2756 P.n2755 0.00196193
R1165 P.n2770 P.n2769 0.00196193
R1166 P.n2282 P.n2281 0.00196193
R1167 P.n2294 P.n2293 0.00196193
R1168 P.n2381 P.n2380 0.00196193
R1169 P.n2383 P.n2382 0.00196193
R1170 P.n2385 P.n2384 0.00196193
R1171 P.n2258 P.n2257 0.00196193
R1172 P.n2270 P.n2269 0.00196193
R1173 P.n2326 P.n2325 0.00196193
R1174 P.n2366 P.n2365 0.00196193
R1175 P.n2378 P.n2377 0.00196193
R1176 P.n2416 P.n2415 0.00196193
R1177 P.n2222 P.n2221 0.00196193
R1178 P.n2235 P.n2234 0.00196193
R1179 P.n3619 P.n3618 0.00196193
R1180 P.n3631 P.n3630 0.00196193
R1181 P.n2056 P.n2055 0.00196193
R1182 P.n2058 P.n2057 0.00196193
R1183 P.n2060 P.n2059 0.00196193
R1184 P.n3595 P.n3594 0.00196193
R1185 P.n3607 P.n3606 0.00196193
R1186 P.n3663 P.n3662 0.00196193
R1187 P.n2041 P.n2040 0.00196193
R1188 P.n2053 P.n2052 0.00196193
R1189 P.n2091 P.n2090 0.00196193
R1190 P.n2155 P.n2154 0.00196193
R1191 P.n2141 P.n2140 0.00196193
R1192 P.n2561 P.n2560 0.00196193
R1193 P.n2573 P.n2572 0.00196193
R1194 P.n2654 P.n2653 0.00196193
R1195 P.n2656 P.n2655 0.00196193
R1196 P.n2658 P.n2657 0.00196193
R1197 P.n2537 P.n2536 0.00196193
R1198 P.n2549 P.n2548 0.00196193
R1199 P.n2605 P.n2604 0.00196193
R1200 P.n2639 P.n2638 0.00196193
R1201 P.n2651 P.n2650 0.00196193
R1202 P.n2689 P.n2688 0.00196193
R1203 P.n2492 P.n2491 0.00196193
R1204 P.n2505 P.n2504 0.00196193
R1205 P.n2990 P.n2989 0.00196193
R1206 P.n3002 P.n3001 0.00196193
R1207 P.n3183 P.n3182 0.00196193
R1208 P.n3185 P.n3184 0.00196193
R1209 P.n3187 P.n3186 0.00196193
R1210 P.n2966 P.n2965 0.00196193
R1211 P.n2978 P.n2977 0.00196193
R1212 P.n3034 P.n3033 0.00196193
R1213 P.n3168 P.n3167 0.00196193
R1214 P.n3180 P.n3179 0.00196193
R1215 P.n3218 P.n3217 0.00196193
R1216 P.n3077 P.n3076 0.00196193
R1217 P.n3259 P.n3258 0.00196193
R1218 P.n1061 P.n1060 0.00194086
R1219 P.n104 P.n103 0.00191935
R1220 P.n785 P.n784 0.00191935
R1221 P.n1894 P.n1893 0.00191315
R1222 P.n1906 P.n1905 0.00191315
R1223 P.n1775 P.n1774 0.00191315
R1224 P.n1777 P.n1776 0.00191315
R1225 P.n1779 P.n1778 0.00191315
R1226 P.n1870 P.n1869 0.00191315
R1227 P.n1882 P.n1881 0.00191315
R1228 P.n1938 P.n1937 0.00191315
R1229 P.n1760 P.n1759 0.00191315
R1230 P.n1772 P.n1771 0.00191315
R1231 P.n1810 P.n1809 0.00191315
R1232 P.n1995 P.n1994 0.00191315
R1233 P.n1844 P.n1843 0.00191315
R1234 P.n1456 P.n1455 0.00191315
R1235 P.n1468 P.n1467 0.00191315
R1236 P.n1576 P.n1575 0.00191315
R1237 P.n1578 P.n1577 0.00191315
R1238 P.n1580 P.n1579 0.00191315
R1239 P.n1432 P.n1431 0.00191315
R1240 P.n1444 P.n1443 0.00191315
R1241 P.n1500 P.n1499 0.00191315
R1242 P.n1561 P.n1560 0.00191315
R1243 P.n1573 P.n1572 0.00191315
R1244 P.n1611 P.n1610 0.00191315
R1245 P.n1526 P.n1525 0.00191315
R1246 P.n1645 P.n1644 0.00191315
R1247 P.n1141 P.n1140 0.00191315
R1248 P.n1153 P.n1152 0.00191315
R1249 P.n1228 P.n1227 0.00191315
R1250 P.n1230 P.n1229 0.00191315
R1251 P.n1232 P.n1231 0.00191315
R1252 P.n1117 P.n1116 0.00191315
R1253 P.n1129 P.n1128 0.00191315
R1254 P.n1185 P.n1184 0.00191315
R1255 P.n1213 P.n1212 0.00191315
R1256 P.n1225 P.n1224 0.00191315
R1257 P.n1263 P.n1262 0.00191315
R1258 P.n1332 P.n1331 0.00191315
R1259 P.n1297 P.n1296 0.00191315
R1260 P.n937 P.n936 0.00191315
R1261 P.n949 P.n948 0.00191315
R1262 P.n819 P.n818 0.00191315
R1263 P.n821 P.n820 0.00191315
R1264 P.n823 P.n822 0.00191315
R1265 P.n913 P.n912 0.00191315
R1266 P.n925 P.n924 0.00191315
R1267 P.n981 P.n980 0.00191315
R1268 P.n804 P.n803 0.00191315
R1269 P.n816 P.n815 0.00191315
R1270 P.n854 P.n853 0.00191315
R1271 P.n1017 P.n1016 0.00191315
R1272 P.n879 P.n878 0.00191315
R1273 P.n221 P.n220 0.00191315
R1274 P.n233 P.n232 0.00191315
R1275 P.n135 P.n134 0.00191315
R1276 P.n137 P.n136 0.00191315
R1277 P.n139 P.n138 0.00191315
R1278 P.n197 P.n196 0.00191315
R1279 P.n209 P.n208 0.00191315
R1280 P.n265 P.n264 0.00191315
R1281 P.n120 P.n119 0.00191315
R1282 P.n132 P.n131 0.00191315
R1283 P.n170 P.n169 0.00191315
R1284 P.n377 P.n376 0.00191315
R1285 P.n332 P.n331 0.00191315
R1286 P.n561 P.n560 0.00191315
R1287 P.n573 P.n572 0.00191315
R1288 P.n450 P.n449 0.00191315
R1289 P.n452 P.n451 0.00191315
R1290 P.n454 P.n453 0.00191315
R1291 P.n537 P.n536 0.00191315
R1292 P.n549 P.n548 0.00191315
R1293 P.n605 P.n604 0.00191315
R1294 P.n435 P.n434 0.00191315
R1295 P.n447 P.n446 0.00191315
R1296 P.n485 P.n484 0.00191315
R1297 P.n705 P.n704 0.00191315
R1298 P.n657 P.n656 0.00191315
R1299 P.n3090 P.n3089 0.00183333
R1300 P.n3133 P.n3132 0.00183333
R1301 P.n312 P.n311 0.00179032
R1302 P.n3499 P.n3498 0.00179032
R1303 P.n2943 P.n2942 0.00177919
R1304 P.n3144 P.n3143 0.00177919
R1305 P.n2857 P.n2839 0.00173096
R1306 P.n2291 P.n2273 0.00173096
R1307 P.n3628 P.n3610 0.00173096
R1308 P.n2570 P.n2552 0.00173096
R1309 P.n2999 P.n2981 0.00173096
R1310 P.n2762 P.n2761 0.00173096
R1311 P.n2913 P.n2911 0.00173096
R1312 P.n2776 P.n2775 0.00173096
R1313 P.n3396 P.n3394 0.00173096
R1314 P.n2349 P.n2345 0.00173096
R1315 P.n2435 P.n2434 0.00173096
R1316 P.n2148 P.n2147 0.00173096
R1317 P.n3692 P.n3690 0.00173096
R1318 P.n2134 P.n2133 0.00173096
R1319 P.n2110 P.n2109 0.00173096
R1320 P.n2625 P.n2624 0.00173096
R1321 P.n2711 P.n2707 0.00173096
R1322 P.n2858 P.n2857 0.00173049
R1323 P.n2292 P.n2291 0.00173049
R1324 P.n3629 P.n3628 0.00173049
R1325 P.n2571 P.n2570 0.00173049
R1326 P.n3000 P.n2999 0.00173049
R1327 P.n1903 P.n1885 0.00170658
R1328 P.n1465 P.n1447 0.00170658
R1329 P.n1150 P.n1132 0.00170658
R1330 P.n946 P.n928 0.00170658
R1331 P.n230 P.n212 0.00170658
R1332 P.n570 P.n552 0.00170658
R1333 P.n1990 P.n1989 0.00170657
R1334 P.n1958 P.n1957 0.00170657
R1335 P.n1861 P.n1860 0.00170657
R1336 P.n1829 P.n1828 0.00170657
R1337 P.n1543 P.n1542 0.00170657
R1338 P.n1520 P.n1519 0.00170657
R1339 P.n1662 P.n1661 0.00170657
R1340 P.n1630 P.n1629 0.00170657
R1341 P.n1327 P.n1326 0.00170657
R1342 P.n1313 P.n1312 0.00170657
R1343 P.n1282 P.n1281 0.00170657
R1344 P.n1034 P.n1033 0.00170657
R1345 P.n1001 P.n1000 0.00170657
R1346 P.n896 P.n895 0.00170657
R1347 P.n873 P.n872 0.00170657
R1348 P.n372 P.n371 0.00170657
R1349 P.n342 P.n341 0.00170657
R1350 P.n700 P.n699 0.00170657
R1351 P.n666 P.n665 0.00170657
R1352 P.n1904 P.n1903 0.00170613
R1353 P.n1466 P.n1465 0.00170613
R1354 P.n1151 P.n1150 0.00170613
R1355 P.n947 P.n946 0.00170613
R1356 P.n231 P.n230 0.00170613
R1357 P.n571 P.n570 0.00170613
R1358 P.n2803 P.n2802 0.00168782
R1359 P.n2800 P.n2799 0.00168782
R1360 P.n3519 P.n3518 0.00168782
R1361 P.n2444 P.n2443 0.00168782
R1362 P.n2178 P.n2177 0.00168782
R1363 P.n2162 P.n2161 0.00168782
R1364 P.n3462 P.n3461 0.00168782
R1365 P.n2714 P.n2713 0.00168782
R1366 P.n2956 P.n2955 0.00168782
R1367 P.n3157 P.n3156 0.00168782
R1368 P.n3283 P.n3105 0.0016828
R1369 P.n1988 P.n1987 0.00164818
R1370 P.n1859 P.n1858 0.00164818
R1371 P.n1541 P.n1540 0.00164818
R1372 P.n1660 P.n1659 0.00164818
R1373 P.n1325 P.n1324 0.00164818
R1374 P.n1311 P.n1310 0.00164818
R1375 P.n1032 P.n1031 0.00164818
R1376 P.n894 P.n893 0.00164818
R1377 P.n370 P.n369 0.00164818
R1378 P.n340 P.n339 0.00164818
R1379 P.n2821 P.n2820 0.00159645
R1380 P.n2827 P.n2826 0.00159645
R1381 P.n3323 P.n3322 0.00159645
R1382 P.n3329 P.n3328 0.00159645
R1383 P.n3288 P.n3287 0.00159645
R1384 P.n2921 P.n2920 0.00159645
R1385 P.n2255 P.n2254 0.00159645
R1386 P.n2261 P.n2260 0.00159645
R1387 P.n2363 P.n2362 0.00159645
R1388 P.n2369 P.n2368 0.00159645
R1389 P.n2459 P.n2458 0.00159645
R1390 P.n2464 P.n2463 0.00159645
R1391 P.n3592 P.n3591 0.00159645
R1392 P.n3598 P.n3597 0.00159645
R1393 P.n2038 P.n2037 0.00159645
R1394 P.n2044 P.n2043 0.00159645
R1395 P.n3569 P.n3568 0.00159645
R1396 P.n2186 P.n2185 0.00159645
R1397 P.n2534 P.n2533 0.00159645
R1398 P.n2540 P.n2539 0.00159645
R1399 P.n2636 P.n2635 0.00159645
R1400 P.n2642 P.n2641 0.00159645
R1401 P.n2724 P.n2723 0.00159645
R1402 P.n2734 P.n2733 0.00159645
R1403 P.n2963 P.n2962 0.00159645
R1404 P.n2969 P.n2968 0.00159645
R1405 P.n3165 P.n3164 0.00159645
R1406 P.n3171 P.n3170 0.00159645
R1407 P.n2947 P.n2946 0.00159645
R1408 P.n3148 P.n3147 0.00159645
R1409 P.n1867 P.n1866 0.00155986
R1410 P.n1873 P.n1872 0.00155986
R1411 P.n1757 P.n1756 0.00155986
R1412 P.n1763 P.n1762 0.00155986
R1413 P.n2006 P.n2005 0.00155986
R1414 P.n1975 P.n1974 0.00155986
R1415 P.n1429 P.n1428 0.00155986
R1416 P.n1435 P.n1434 0.00155986
R1417 P.n1558 P.n1557 0.00155986
R1418 P.n1564 P.n1563 0.00155986
R1419 P.n1670 P.n1669 0.00155986
R1420 P.n1678 P.n1677 0.00155986
R1421 P.n1114 P.n1113 0.00155986
R1422 P.n1120 P.n1119 0.00155986
R1423 P.n1210 P.n1209 0.00155986
R1424 P.n1216 P.n1215 0.00155986
R1425 P.n1351 P.n1350 0.00155986
R1426 P.n1344 P.n1343 0.00155986
R1427 P.n910 P.n909 0.00155986
R1428 P.n916 P.n915 0.00155986
R1429 P.n801 P.n800 0.00155986
R1430 P.n807 P.n806 0.00155986
R1431 P.n1043 P.n1042 0.00155986
R1432 P.n903 P.n902 0.00155986
R1433 P.n194 P.n193 0.00155986
R1434 P.n200 P.n199 0.00155986
R1435 P.n117 P.n116 0.00155986
R1436 P.n123 P.n122 0.00155986
R1437 P.n390 P.n389 0.00155986
R1438 P.n350 P.n349 0.00155986
R1439 P.n534 P.n533 0.00155986
R1440 P.n540 P.n539 0.00155986
R1441 P.n432 P.n431 0.00155986
R1442 P.n438 P.n437 0.00155986
R1443 P.n716 P.n715 0.00155986
R1444 P.n673 P.n672 0.00155986
R1445 P.n2931 P.n2930 0.00155376
R1446 P.n3275 P.n3274 0.00155376
R1447 P.n2819 P.n2818 0.00154822
R1448 P.n3320 P.n3319 0.00154822
R1449 P.n2253 P.n2252 0.00154822
R1450 P.n2360 P.n2359 0.00154822
R1451 P.n3689 P.n3688 0.00154822
R1452 P.n2035 P.n2034 0.00154822
R1453 P.n2532 P.n2531 0.00154822
R1454 P.n2633 P.n2632 0.00154822
R1455 P.n1728 P.n1727 0.00152993
R1456 P.n1718 P.n1717 0.00152993
R1457 P.n1427 P.n1426 0.00152993
R1458 P.n1555 P.n1554 0.00152993
R1459 P.n1112 P.n1111 0.00152993
R1460 P.n1075 P.n1074 0.00152993
R1461 P.n765 P.n764 0.00152993
R1462 P.n753 P.n752 0.00152993
R1463 P.n292 P.n291 0.00152993
R1464 P.n189 P.n114 0.00152993
R1465 P.n625 P.n532 0.00152993
R1466 P.n511 P.n510 0.00152993
R1467 P.n427 P.n426 0.00143007
R1468 P.n1065 P.n1064 0.00143007
R1469 P.n1064 P.n1063 0.00143007
R1470 P.n426 P.n418 0.00143007
R1471 P.n411 P.n410 0.00143007
R1472 P.n105 P.n104 0.00142473
R1473 P.n414 P.n413 0.00141932
R1474 P.n1055 P.n1054 0.00141932
R1475 P.n1063 P.n1062 0.00141932
R1476 P.n3417 P.n3416 0.00141932
R1477 P.n3398 P.n3397 0.00141932
R1478 P.n413 P.n412 0.00141932
R1479 P.n401 P.n400 0.00141932
R1480 P.n1062 P.n1061 0.00141932
R1481 P.n1054 P.n1053 0.00141932
R1482 P.n3399 P.n3398 0.00141932
R1483 P.n3418 P.n3417 0.00141932
R1484 P.n2760 P.n2759 0.00141371
R1485 P.n2774 P.n2773 0.00141371
R1486 P.n2226 P.n2225 0.00141371
R1487 P.n2239 P.n2238 0.00141371
R1488 P.n2159 P.n2158 0.00141371
R1489 P.n2145 P.n2144 0.00141371
R1490 P.n2496 P.n2495 0.00141371
R1491 P.n2509 P.n2508 0.00141371
R1492 P.n3081 P.n3080 0.00141371
R1493 P.n3263 P.n3262 0.00141371
R1494 P.n1999 P.n1998 0.00138322
R1495 P.n1848 P.n1847 0.00138322
R1496 P.n1530 P.n1529 0.00138322
R1497 P.n1649 P.n1648 0.00138322
R1498 P.n1336 P.n1335 0.00138322
R1499 P.n1301 P.n1300 0.00138322
R1500 P.n1021 P.n1020 0.00138322
R1501 P.n883 P.n882 0.00138322
R1502 P.n381 P.n380 0.00138322
R1503 P.n336 P.n335 0.00138322
R1504 P.n709 P.n708 0.00138322
R1505 P.n661 P.n660 0.00138322
R1506 P.n1060 P.n1059 0.00138172
R1507 P.n1059 P.n1058 0.00136021
R1508 P.n3397 P.n3312 0.00136021
R1509 P.n2852 P.n2851 0.00132234
R1510 P.n2842 P.n2841 0.00132234
R1511 P.n2877 P.n2876 0.00132234
R1512 P.n3361 P.n3360 0.00132234
R1513 P.n3301 P.n3300 0.00132234
R1514 P.n2916 P.n2915 0.00132234
R1515 P.n2286 P.n2285 0.00132234
R1516 P.n2276 P.n2275 0.00132234
R1517 P.n2311 P.n2310 0.00132234
R1518 P.n2401 P.n2400 0.00132234
R1519 P.n2449 P.n2448 0.00132234
R1520 P.n2454 P.n2453 0.00132234
R1521 P.n3623 P.n3622 0.00132234
R1522 P.n3613 P.n3612 0.00132234
R1523 P.n3648 P.n3647 0.00132234
R1524 P.n2076 P.n2075 0.00132234
R1525 P.n3566 P.n3565 0.00132234
R1526 P.n2183 P.n2182 0.00132234
R1527 P.n2565 P.n2564 0.00132234
R1528 P.n2555 P.n2554 0.00132234
R1529 P.n2590 P.n2589 0.00132234
R1530 P.n2674 P.n2673 0.00132234
R1531 P.n2730 P.n2729 0.00132234
R1532 P.n2741 P.n2740 0.00132234
R1533 P.n2994 P.n2993 0.00132234
R1534 P.n2984 P.n2983 0.00132234
R1535 P.n3019 P.n3018 0.00132234
R1536 P.n3203 P.n3202 0.00132234
R1537 P.n3140 P.n3139 0.00132234
R1538 P.n1898 P.n1897 0.0012949
R1539 P.n1888 P.n1887 0.0012949
R1540 P.n1923 P.n1922 0.0012949
R1541 P.n1795 P.n1794 0.0012949
R1542 P.n1741 P.n1740 0.0012949
R1543 P.n1735 P.n1734 0.0012949
R1544 P.n1460 P.n1459 0.0012949
R1545 P.n1450 P.n1449 0.0012949
R1546 P.n1485 P.n1484 0.0012949
R1547 P.n1596 P.n1595 0.0012949
R1548 P.n1390 P.n1389 0.0012949
R1549 P.n1397 P.n1396 0.0012949
R1550 P.n1145 P.n1144 0.0012949
R1551 P.n1135 P.n1134 0.0012949
R1552 P.n1170 P.n1169 0.0012949
R1553 P.n1248 P.n1247 0.0012949
R1554 P.n1086 P.n1085 0.0012949
R1555 P.n1082 P.n1081 0.0012949
R1556 P.n941 P.n940 0.0012949
R1557 P.n931 P.n930 0.0012949
R1558 P.n966 P.n965 0.0012949
R1559 P.n839 P.n838 0.0012949
R1560 P.n778 P.n777 0.0012949
R1561 P.n771 P.n770 0.0012949
R1562 P.n225 P.n224 0.0012949
R1563 P.n215 P.n214 0.0012949
R1564 P.n250 P.n249 0.0012949
R1565 P.n155 P.n154 0.0012949
R1566 P.n306 P.n305 0.0012949
R1567 P.n299 P.n298 0.0012949
R1568 P.n565 P.n564 0.0012949
R1569 P.n555 P.n554 0.0012949
R1570 P.n590 P.n589 0.0012949
R1571 P.n470 P.n469 0.0012949
R1572 P.n632 P.n631 0.0012949
R1573 P.n519 P.n518 0.0012949
R1574 P.n1057 P.n1056 0.00127419
R1575 P.n3404 P.n3403 0.00127419
R1576 P.n2765 P.n2764 0.00127411
R1577 P.n2779 P.n2778 0.00127411
R1578 P.n2230 P.n2229 0.00127411
R1579 P.n2348 P.n2347 0.00127411
R1580 P.n2243 P.n2242 0.00127411
R1581 P.n2352 P.n2351 0.00127411
R1582 P.n2151 P.n2150 0.00127411
R1583 P.n2137 P.n2136 0.00127411
R1584 P.n2112 P.n2111 0.00127411
R1585 P.n2488 P.n2487 0.00127411
R1586 P.n2524 P.n2523 0.00127411
R1587 P.n2501 P.n2500 0.00127411
R1588 P.n2710 P.n2709 0.00127411
R1589 P.n2002 P.n1992 0.00126496
R1590 P.n1970 P.n1959 0.00126496
R1591 P.n1864 P.n1863 0.00126496
R1592 P.n1840 P.n1830 0.00126496
R1593 P.n1546 P.n1545 0.00126496
R1594 P.n1522 P.n1521 0.00126496
R1595 P.n1665 P.n1664 0.00126496
R1596 P.n1641 P.n1631 0.00126496
R1597 P.n1339 P.n1329 0.00126496
R1598 P.n1207 P.n1206 0.00126496
R1599 P.n1316 P.n1315 0.00126496
R1600 P.n1293 P.n1283 0.00126496
R1601 P.n1037 P.n1036 0.00126496
R1602 P.n1013 P.n1002 0.00126496
R1603 P.n899 P.n898 0.00126496
R1604 P.n875 P.n874 0.00126496
R1605 P.n384 P.n374 0.00126496
R1606 P.n367 P.n356 0.00126496
R1607 P.n345 P.n344 0.00126496
R1608 P.n328 P.n318 0.00126496
R1609 P.n712 P.n702 0.00126496
R1610 P.n696 P.n695 0.00126496
R1611 P.n669 P.n668 0.00126496
R1612 P.n653 P.n643 0.00126496
R1613 P.n2932 P.n2931 0.00123118
R1614 P.n3274 P.n3273 0.00123118
R1615 P.n2855 P.n2854 0.00123096
R1616 P.n2845 P.n2844 0.00123096
R1617 P.n2864 P.n2863 0.00123096
R1618 P.n2883 P.n2882 0.00123096
R1619 P.n2880 P.n2879 0.00123096
R1620 P.n3349 P.n3348 0.00123096
R1621 P.n3367 P.n3366 0.00123096
R1622 P.n3364 P.n3363 0.00123096
R1623 P.n2289 P.n2288 0.00123096
R1624 P.n2279 P.n2278 0.00123096
R1625 P.n2298 P.n2297 0.00123096
R1626 P.n2317 P.n2316 0.00123096
R1627 P.n2314 P.n2313 0.00123096
R1628 P.n2389 P.n2388 0.00123096
R1629 P.n2407 P.n2406 0.00123096
R1630 P.n2404 P.n2403 0.00123096
R1631 P.n3626 P.n3625 0.00123096
R1632 P.n3616 P.n3615 0.00123096
R1633 P.n3635 P.n3634 0.00123096
R1634 P.n3654 P.n3653 0.00123096
R1635 P.n3651 P.n3650 0.00123096
R1636 P.n2064 P.n2063 0.00123096
R1637 P.n2082 P.n2081 0.00123096
R1638 P.n2079 P.n2078 0.00123096
R1639 P.n2568 P.n2567 0.00123096
R1640 P.n2558 P.n2557 0.00123096
R1641 P.n2577 P.n2576 0.00123096
R1642 P.n2596 P.n2595 0.00123096
R1643 P.n2593 P.n2592 0.00123096
R1644 P.n2662 P.n2661 0.00123096
R1645 P.n2680 P.n2679 0.00123096
R1646 P.n2677 P.n2676 0.00123096
R1647 P.n2997 P.n2996 0.00123096
R1648 P.n2987 P.n2986 0.00123096
R1649 P.n3006 P.n3005 0.00123096
R1650 P.n3025 P.n3024 0.00123096
R1651 P.n3022 P.n3021 0.00123096
R1652 P.n3191 P.n3190 0.00123096
R1653 P.n3209 P.n3208 0.00123096
R1654 P.n3206 P.n3205 0.00123096
R1655 P.n1901 P.n1900 0.00120658
R1656 P.n1891 P.n1890 0.00120658
R1657 P.n1910 P.n1909 0.00120658
R1658 P.n1929 P.n1928 0.00120658
R1659 P.n1926 P.n1925 0.00120658
R1660 P.n1783 P.n1782 0.00120658
R1661 P.n1801 P.n1800 0.00120658
R1662 P.n1798 P.n1797 0.00120658
R1663 P.n1463 P.n1462 0.00120658
R1664 P.n1453 P.n1452 0.00120658
R1665 P.n1472 P.n1471 0.00120658
R1666 P.n1491 P.n1490 0.00120658
R1667 P.n1488 P.n1487 0.00120658
R1668 P.n1584 P.n1583 0.00120658
R1669 P.n1602 P.n1601 0.00120658
R1670 P.n1599 P.n1598 0.00120658
R1671 P.n1148 P.n1147 0.00120658
R1672 P.n1138 P.n1137 0.00120658
R1673 P.n1157 P.n1156 0.00120658
R1674 P.n1176 P.n1175 0.00120658
R1675 P.n1173 P.n1172 0.00120658
R1676 P.n1236 P.n1235 0.00120658
R1677 P.n1254 P.n1253 0.00120658
R1678 P.n1251 P.n1250 0.00120658
R1679 P.n944 P.n943 0.00120658
R1680 P.n934 P.n933 0.00120658
R1681 P.n953 P.n952 0.00120658
R1682 P.n972 P.n971 0.00120658
R1683 P.n969 P.n968 0.00120658
R1684 P.n827 P.n826 0.00120658
R1685 P.n845 P.n844 0.00120658
R1686 P.n842 P.n841 0.00120658
R1687 P.n228 P.n227 0.00120658
R1688 P.n218 P.n217 0.00120658
R1689 P.n237 P.n236 0.00120658
R1690 P.n256 P.n255 0.00120658
R1691 P.n253 P.n252 0.00120658
R1692 P.n143 P.n142 0.00120658
R1693 P.n161 P.n160 0.00120658
R1694 P.n158 P.n157 0.00120658
R1695 P.n568 P.n567 0.00120658
R1696 P.n558 P.n557 0.00120658
R1697 P.n577 P.n576 0.00120658
R1698 P.n596 P.n595 0.00120658
R1699 P.n593 P.n592 0.00120658
R1700 P.n458 P.n457 0.00120658
R1701 P.n476 P.n475 0.00120658
R1702 P.n473 P.n472 0.00120658
R1703 P.n3401 P.n3400 0.00118817
R1704 P.n415 P.n414 0.00116667
R1705 P.n3302 P.n3301 0.00113959
R1706 P.n2807 P.n2806 0.00113959
R1707 P.n2809 P.n2808 0.00113959
R1708 P.n2813 P.n2812 0.00113959
R1709 P.n2915 P.n2914 0.00113959
R1710 P.n2917 P.n2916 0.00113959
R1711 P.n2795 P.n2794 0.00113959
R1712 P.n2797 P.n2796 0.00113959
R1713 P.n3314 P.n3313 0.00113959
R1714 P.n2450 P.n2449 0.00113959
R1715 P.n3523 P.n3522 0.00113959
R1716 P.n3525 P.n3524 0.00113959
R1717 P.n3518 P.n3517 0.00113959
R1718 P.n2247 P.n2246 0.00113959
R1719 P.n2453 P.n2452 0.00113959
R1720 P.n2455 P.n2454 0.00113959
R1721 P.n2438 P.n2437 0.00113959
R1722 P.n2440 P.n2439 0.00113959
R1723 P.n2443 P.n2442 0.00113959
R1724 P.n2354 P.n2353 0.00113959
R1725 P.n3567 P.n3566 0.00113959
R1726 P.n2173 P.n2172 0.00113959
R1727 P.n2175 P.n2174 0.00113959
R1728 P.n3683 P.n3682 0.00113959
R1729 P.n2182 P.n2181 0.00113959
R1730 P.n2184 P.n2183 0.00113959
R1731 P.n2166 P.n2165 0.00113959
R1732 P.n2168 P.n2167 0.00113959
R1733 P.n2029 P.n2028 0.00113959
R1734 P.n2731 P.n2730 0.00113959
R1735 P.n3456 P.n3455 0.00113959
R1736 P.n3458 P.n3457 0.00113959
R1737 P.n3461 P.n3460 0.00113959
R1738 P.n2526 P.n2525 0.00113959
R1739 P.n2740 P.n2739 0.00113959
R1740 P.n2742 P.n2741 0.00113959
R1741 P.n2718 P.n2717 0.00113959
R1742 P.n2720 P.n2719 0.00113959
R1743 P.n2713 P.n2712 0.00113959
R1744 P.n2627 P.n2626 0.00113959
R1745 P.n2950 P.n2949 0.00113959
R1746 P.n2952 P.n2951 0.00113959
R1747 P.n2957 P.n2956 0.00113959
R1748 P.n2958 P.n2957 0.00113959
R1749 P.n3074 P.n3073 0.00113959
R1750 P.n3066 P.n3065 0.00113959
R1751 P.n3139 P.n3138 0.00113959
R1752 P.n3141 P.n3140 0.00113959
R1753 P.n3151 P.n3150 0.00113959
R1754 P.n3153 P.n3152 0.00113959
R1755 P.n3158 P.n3157 0.00113959
R1756 P.n3159 P.n3158 0.00113959
R1757 P.n3256 P.n3255 0.00113959
R1758 P.n3248 P.n3247 0.00113959
R1759 P.n83 P.n82 0.00112366
R1760 P.n85 P.n84 0.00112366
R1761 P.n101 P.n93 0.00112366
R1762 P.n103 P.n102 0.00112366
R1763 P.n311 P.n310 0.00112366
R1764 P.n638 P.n637 0.00112366
R1765 P.n1091 P.n1090 0.00112366
R1766 P.n1370 P.n1369 0.00112366
R1767 P.n1376 P.n1375 0.00112366
R1768 P.n3699 P.n3698 0.00112366
R1769 P.n3693 P.n3590 0.00112366
R1770 P.n3542 P.n3541 0.00112366
R1771 P.n3532 P.n3531 0.00112366
R1772 P.n3530 P.n3529 0.00112366
R1773 P.n3528 P.n3516 0.00112366
R1774 P.n3515 P.n3514 0.00112366
R1775 P.n3500 P.n3499 0.00112366
R1776 P.n3299 P.n3298 0.00112366
R1777 P.n1742 P.n1741 0.00111825
R1778 P.n1981 P.n1980 0.00111825
R1779 P.n1983 P.n1982 0.00111825
R1780 P.n1989 P.n1988 0.00111825
R1781 P.n1722 P.n1721 0.00111825
R1782 P.n1734 P.n1733 0.00111825
R1783 P.n1736 P.n1735 0.00111825
R1784 P.n1852 P.n1851 0.00111825
R1785 P.n1854 P.n1853 0.00111825
R1786 P.n1860 P.n1859 0.00111825
R1787 P.n1712 P.n1711 0.00111825
R1788 P.n1391 P.n1390 0.00111825
R1789 P.n1534 P.n1533 0.00111825
R1790 P.n1536 P.n1535 0.00111825
R1791 P.n1542 P.n1541 0.00111825
R1792 P.n1421 P.n1420 0.00111825
R1793 P.n1396 P.n1395 0.00111825
R1794 P.n1398 P.n1397 0.00111825
R1795 P.n1653 P.n1652 0.00111825
R1796 P.n1655 P.n1654 0.00111825
R1797 P.n1661 P.n1660 0.00111825
R1798 P.n1549 P.n1548 0.00111825
R1799 P.n1087 P.n1086 0.00111825
R1800 P.n1318 P.n1317 0.00111825
R1801 P.n1320 P.n1319 0.00111825
R1802 P.n1326 P.n1325 0.00111825
R1803 P.n1106 P.n1105 0.00111825
R1804 P.n1205 P.n1204 0.00111825
R1805 P.n1081 P.n1080 0.00111825
R1806 P.n1083 P.n1082 0.00111825
R1807 P.n1305 P.n1304 0.00111825
R1808 P.n1307 P.n1306 0.00111825
R1809 P.n1312 P.n1311 0.00111825
R1810 P.n1069 P.n1068 0.00111825
R1811 P.n779 P.n778 0.00111825
R1812 P.n1025 P.n1024 0.00111825
R1813 P.n1027 P.n1026 0.00111825
R1814 P.n1033 P.n1032 0.00111825
R1815 P.n759 P.n758 0.00111825
R1816 P.n770 P.n769 0.00111825
R1817 P.n772 P.n771 0.00111825
R1818 P.n887 P.n886 0.00111825
R1819 P.n889 P.n888 0.00111825
R1820 P.n895 P.n894 0.00111825
R1821 P.n747 P.n746 0.00111825
R1822 P.n307 P.n306 0.00111825
R1823 P.n95 P.n94 0.00111825
R1824 P.n97 P.n96 0.00111825
R1825 P.n371 P.n370 0.00111825
R1826 P.n286 P.n285 0.00111825
R1827 P.n298 P.n297 0.00111825
R1828 P.n300 P.n299 0.00111825
R1829 P.n87 P.n86 0.00111825
R1830 P.n89 P.n88 0.00111825
R1831 P.n341 P.n340 0.00111825
R1832 P.n109 P.n108 0.00111825
R1833 P.n633 P.n632 0.00111825
R1834 P.n420 P.n419 0.00111825
R1835 P.n422 P.n421 0.00111825
R1836 P.n699 P.n698 0.00111825
R1837 P.n527 P.n526 0.00111825
R1838 P.n518 P.n517 0.00111825
R1839 P.n520 P.n519 0.00111825
R1840 P.n56 P.n55 0.00111825
R1841 P.n58 P.n57 0.00111825
R1842 P.n665 P.n664 0.00111825
R1843 P.n505 P.n504 0.00111825
R1844 P.n74 P.n73 0.00110752
R1845 P.n1361 P.n1360 0.00110215
R1846 P.n1374 P.n1373 0.00110215
R1847 P.n3707 P.n3706 0.00110215
R1848 P.n3695 P.n3694 0.00110215
R1849 P.n3304 P.n3303 0.00109137
R1850 P.n3291 P.n3290 0.00109137
R1851 P.n2811 P.n2810 0.00109137
R1852 P.n2763 P.n2762 0.00109137
R1853 P.n2766 P.n2765 0.00109137
R1854 P.n2913 P.n2912 0.00109137
R1855 P.n3414 P.n3413 0.00109137
R1856 P.n2919 P.n2918 0.00109137
R1857 P.n2924 P.n2923 0.00109137
R1858 P.n2777 P.n2776 0.00109137
R1859 P.n2781 P.n2774 0.00109137
R1860 P.n3396 P.n3395 0.00109137
R1861 P.n2745 P.n2744 0.00109137
R1862 P.n2462 P.n2461 0.00109137
R1863 P.n3527 P.n3526 0.00109137
R1864 P.n2228 P.n2227 0.00109137
R1865 P.n2231 P.n2230 0.00109137
R1866 P.n2345 P.n2253 0.00109137
R1867 P.n2349 P.n2348 0.00109137
R1868 P.n2347 P.n2346 0.00109137
R1869 P.n2211 P.n2210 0.00109137
R1870 P.n2457 P.n2456 0.00109137
R1871 P.n2467 P.n2466 0.00109137
R1872 P.n2446 P.n2445 0.00109137
R1873 P.n2244 P.n2243 0.00109137
R1874 P.n2245 P.n2239 0.00109137
R1875 P.n2434 P.n2360 0.00109137
R1876 P.n2351 P.n2350 0.00109137
R1877 P.n3574 P.n3573 0.00109137
R1878 P.n3572 P.n3571 0.00109137
R1879 P.n2180 P.n2179 0.00109137
R1880 P.n2149 P.n2148 0.00109137
R1881 P.n2152 P.n2151 0.00109137
R1882 P.n2160 P.n2159 0.00109137
R1883 P.n3692 P.n3691 0.00109137
R1884 P.n2123 P.n2122 0.00109137
R1885 P.n2132 P.n2131 0.00109137
R1886 P.n2191 P.n2190 0.00109137
R1887 P.n2170 P.n2169 0.00109137
R1888 P.n2135 P.n2134 0.00109137
R1889 P.n2138 P.n2137 0.00109137
R1890 P.n2146 P.n2145 0.00109137
R1891 P.n2109 P.n2035 0.00109137
R1892 P.n2111 P.n2110 0.00109137
R1893 P.n2121 P.n2120 0.00109137
R1894 P.n3464 P.n3463 0.00109137
R1895 P.n2486 P.n2485 0.00109137
R1896 P.n2489 P.n2488 0.00109137
R1897 P.n2497 P.n2496 0.00109137
R1898 P.n2624 P.n2532 0.00109137
R1899 P.n2476 P.n2475 0.00109137
R1900 P.n2722 P.n2715 0.00109137
R1901 P.n2499 P.n2498 0.00109137
R1902 P.n2502 P.n2501 0.00109137
R1903 P.n2510 P.n2509 0.00109137
R1904 P.n2707 P.n2633 0.00109137
R1905 P.n2711 P.n2710 0.00109137
R1906 P.n2484 P.n2483 0.00109137
R1907 P.n2722 P.n2721 0.00109137
R1908 P.n2113 P.n2112 0.00109137
R1909 P.n2435 P.n2352 0.00109137
R1910 P.n2709 P.n2708 0.00109137
R1911 P.n2911 P.n2819 0.00109137
R1912 P.n2767 P.n2760 0.00109137
R1913 P.n3527 P.n3520 0.00109137
R1914 P.n2811 P.n2804 0.00109137
R1915 P.n2625 P.n2524 0.00109137
R1916 P.n2732 P.n2728 0.00109137
R1917 P.n2737 P.n2736 0.00109137
R1918 P.n2743 P.n2738 0.00109137
R1919 P.n2523 P.n2522 0.00109137
R1920 P.n2451 P.n2447 0.00109137
R1921 P.n3464 P.n3459 0.00109137
R1922 P.n2232 P.n2226 0.00109137
R1923 P.n3415 P.n3412 0.00109137
R1924 P.n2780 P.n2779 0.00109137
R1925 P.n3394 P.n3320 0.00109137
R1926 P.n3690 P.n3689 0.00109137
R1927 P.n2189 P.n2188 0.00109137
R1928 P.n2170 P.n2163 0.00109137
R1929 P.n2180 P.n2176 0.00109137
R1930 P.n2219 P.n2218 0.00109137
R1931 P.n2241 P.n2240 0.00109137
R1932 P.n2446 P.n2441 0.00109137
R1933 P.n2727 P.n2726 0.00109137
R1934 P.n1744 P.n1743 0.00108832
R1935 P.n2009 P.n2008 0.00108832
R1936 P.n1986 P.n1985 0.00108832
R1937 P.n1991 P.n1990 0.00108832
R1938 P.n2002 P.n2001 0.00108832
R1939 P.n2000 P.n1999 0.00108832
R1940 P.n1959 P.n1958 0.00108832
R1941 P.n1970 P.n1969 0.00108832
R1942 P.n1978 P.n1977 0.00108832
R1943 P.n1857 P.n1856 0.00108832
R1944 P.n1862 P.n1861 0.00108832
R1945 P.n1849 P.n1848 0.00108832
R1946 P.n1830 P.n1829 0.00108832
R1947 P.n1840 P.n1839 0.00108832
R1948 P.n1838 P.n1837 0.00108832
R1949 P.n1673 P.n1672 0.00108832
R1950 P.n1539 P.n1538 0.00108832
R1951 P.n1544 P.n1543 0.00108832
R1952 P.n1546 P.n1532 0.00108832
R1953 P.n1531 P.n1530 0.00108832
R1954 P.n1519 P.n1427 0.00108832
R1955 P.n1681 P.n1680 0.00108832
R1956 P.n1658 P.n1657 0.00108832
R1957 P.n1663 P.n1662 0.00108832
R1958 P.n1665 P.n1651 0.00108832
R1959 P.n1650 P.n1649 0.00108832
R1960 P.n1629 P.n1555 0.00108832
R1961 P.n1631 P.n1630 0.00108832
R1962 P.n1641 P.n1640 0.00108832
R1963 P.n1354 P.n1353 0.00108832
R1964 P.n1323 P.n1322 0.00108832
R1965 P.n1328 P.n1327 0.00108832
R1966 P.n1339 P.n1338 0.00108832
R1967 P.n1204 P.n1112 0.00108832
R1968 P.n1207 P.n1104 0.00108832
R1969 P.n1347 P.n1346 0.00108832
R1970 P.n1314 P.n1313 0.00108832
R1971 P.n1316 P.n1303 0.00108832
R1972 P.n1302 P.n1301 0.00108832
R1973 P.n1283 P.n1282 0.00108832
R1974 P.n1293 P.n1292 0.00108832
R1975 P.n1046 P.n1045 0.00108832
R1976 P.n1030 P.n1029 0.00108832
R1977 P.n1035 P.n1034 0.00108832
R1978 P.n1037 P.n1023 0.00108832
R1979 P.n1002 P.n1001 0.00108832
R1980 P.n1013 P.n1012 0.00108832
R1981 P.n891 P.n890 0.00108832
R1982 P.n897 P.n896 0.00108832
R1983 P.n899 P.n885 0.00108832
R1984 P.n884 P.n883 0.00108832
R1985 P.n874 P.n873 0.00108832
R1986 P.n797 P.n796 0.00108832
R1987 P.n394 P.n392 0.00108832
R1988 P.n100 P.n99 0.00108832
R1989 P.n373 P.n372 0.00108832
R1990 P.n384 P.n383 0.00108832
R1991 P.n382 P.n381 0.00108832
R1992 P.n356 P.n355 0.00108832
R1993 P.n367 P.n366 0.00108832
R1994 P.n365 P.n364 0.00108832
R1995 P.n92 P.n91 0.00108832
R1996 P.n343 P.n342 0.00108832
R1997 P.n345 P.n338 0.00108832
R1998 P.n189 P.n188 0.00108832
R1999 P.n318 P.n317 0.00108832
R2000 P.n328 P.n327 0.00108832
R2001 P.n635 P.n634 0.00108832
R2002 P.n701 P.n700 0.00108832
R2003 P.n712 P.n711 0.00108832
R2004 P.n625 P.n624 0.00108832
R2005 P.n695 P.n694 0.00108832
R2006 P.n692 P.n691 0.00108832
R2007 P.n522 P.n521 0.00108832
R2008 P.n667 P.n666 0.00108832
R2009 P.n662 P.n661 0.00108832
R2010 P.n643 P.n642 0.00108832
R2011 P.n653 P.n652 0.00108832
R2012 P.n719 P.n718 0.00108832
R2013 P.n875 P.n798 0.00108832
R2014 P.n1337 P.n1336 0.00108832
R2015 P.n1291 P.n1290 0.00108832
R2016 P.n1985 P.n1984 0.00108832
R2017 P.n1522 P.n1419 0.00108832
R2018 P.n1521 P.n1520 0.00108832
R2019 P.n1968 P.n1967 0.00108832
R2020 P.n1864 P.n1850 0.00108832
R2021 P.n1856 P.n1855 0.00108832
R2022 P.n1657 P.n1656 0.00108832
R2023 P.n1418 P.n1417 0.00108832
R2024 P.n1322 P.n1321 0.00108832
R2025 P.n1538 P.n1537 0.00108832
R2026 P.n1029 P.n1028 0.00108832
R2027 P.n1022 P.n1021 0.00108832
R2028 P.n1011 P.n1010 0.00108832
R2029 P.n907 P.n905 0.00108832
R2030 P.n892 P.n891 0.00108832
R2031 P.n292 P.n284 0.00108832
R2032 P.n353 P.n352 0.00108832
R2033 P.n100 P.n98 0.00108832
R2034 P.n696 P.n693 0.00108832
R2035 P.n676 P.n675 0.00108832
R2036 P.n511 P.n503 0.00108832
R2037 P.n1639 P.n1638 0.00108832
R2038 P.n669 P.n663 0.00108832
R2039 P.n301 P.n296 0.00108832
R2040 P.n92 P.n90 0.00108832
R2041 P.n337 P.n336 0.00108832
R2042 P.n403 P.n402 0.00108064
R2043 P.n406 P.n405 0.00108064
R2044 P.n409 P.n408 0.00108064
R2045 P.n2929 P.n2928 0.00105914
R2046 P.n3281 P.n3280 0.00105914
R2047 P.n3277 P.n3276 0.00105914
R2048 P.n80 P.n79 0.00105914
R2049 P.n417 P.n416 0.00105914
R2050 P.n3535 P.n3534 0.00105914
R2051 P.n2881 P.n2880 0.00104822
R2052 P.n2869 P.n2868 0.00104822
R2053 P.n3365 P.n3364 0.00104822
R2054 P.n3353 P.n3352 0.00104822
R2055 P.n2888 P.n2887 0.00104822
R2056 P.n3372 P.n3371 0.00104822
R2057 P.n2315 P.n2314 0.00104822
R2058 P.n2303 P.n2302 0.00104822
R2059 P.n2405 P.n2404 0.00104822
R2060 P.n2393 P.n2392 0.00104822
R2061 P.n2322 P.n2321 0.00104822
R2062 P.n2412 P.n2411 0.00104822
R2063 P.n3652 P.n3651 0.00104822
R2064 P.n3640 P.n3639 0.00104822
R2065 P.n2080 P.n2079 0.00104822
R2066 P.n2068 P.n2067 0.00104822
R2067 P.n3659 P.n3658 0.00104822
R2068 P.n2087 P.n2086 0.00104822
R2069 P.n2594 P.n2593 0.00104822
R2070 P.n2582 P.n2581 0.00104822
R2071 P.n2678 P.n2677 0.00104822
R2072 P.n2666 P.n2665 0.00104822
R2073 P.n2601 P.n2600 0.00104822
R2074 P.n2685 P.n2684 0.00104822
R2075 P.n3023 P.n3022 0.00104822
R2076 P.n3011 P.n3010 0.00104822
R2077 P.n3207 P.n3206 0.00104822
R2078 P.n3195 P.n3194 0.00104822
R2079 P.n3030 P.n3029 0.00104822
R2080 P.n3214 P.n3213 0.00104822
R2081 P.n76 P.n75 0.00103763
R2082 P.n3703 P.n3702 0.00103763
R2083 P.n3539 P.n3538 0.00103763
R2084 P.n1927 P.n1926 0.00102993
R2085 P.n1915 P.n1914 0.00102993
R2086 P.n1799 P.n1798 0.00102993
R2087 P.n1787 P.n1786 0.00102993
R2088 P.n1934 P.n1933 0.00102993
R2089 P.n1806 P.n1805 0.00102993
R2090 P.n1489 P.n1488 0.00102993
R2091 P.n1477 P.n1476 0.00102993
R2092 P.n1600 P.n1599 0.00102993
R2093 P.n1588 P.n1587 0.00102993
R2094 P.n1496 P.n1495 0.00102993
R2095 P.n1607 P.n1606 0.00102993
R2096 P.n1174 P.n1173 0.00102993
R2097 P.n1162 P.n1161 0.00102993
R2098 P.n1252 P.n1251 0.00102993
R2099 P.n1240 P.n1239 0.00102993
R2100 P.n1181 P.n1180 0.00102993
R2101 P.n1259 P.n1258 0.00102993
R2102 P.n970 P.n969 0.00102993
R2103 P.n958 P.n957 0.00102993
R2104 P.n843 P.n842 0.00102993
R2105 P.n831 P.n830 0.00102993
R2106 P.n977 P.n976 0.00102993
R2107 P.n850 P.n849 0.00102993
R2108 P.n254 P.n253 0.00102993
R2109 P.n242 P.n241 0.00102993
R2110 P.n159 P.n158 0.00102993
R2111 P.n147 P.n146 0.00102993
R2112 P.n261 P.n260 0.00102993
R2113 P.n166 P.n165 0.00102993
R2114 P.n594 P.n593 0.00102993
R2115 P.n582 P.n581 0.00102993
R2116 P.n474 P.n473 0.00102993
R2117 P.n462 P.n461 0.00102993
R2118 P.n601 P.n600 0.00102993
R2119 P.n481 P.n480 0.00102993
R2120 P.n3093 P.n3092 0.00101613
R2121 P.n3105 P.n3104 0.00101613
R2122 P.n3130 P.n3129 0.00101613
R2123 P.n3118 P.n3117 0.00101613
R2124 P.n630 P.n629 0.000994624
R2125 P.n725 P.n724 0.000994624
R2126 P.n735 P.n734 0.000994624
R2127 P.n737 P.n736 0.000994624
R2128 P.n739 P.n738 0.000994624
R2129 P.n784 P.n783 0.000994624
R2130 P.n1079 P.n1078 0.000994624
R2131 P.n1700 P.n1699 0.000994624
R2132 P.n1706 P.n1705 0.000994624
R2133 P.n3307 P.n3306 0.000994624
R2134 P.n3100 P.n3099 0.000973118
R2135 P.n3123 P.n3122 0.000973118
R2136 P.n512 P.n429 0.000973118
R2137 P.n1076 P.n1067 0.000973118
R2138 P.n1692 P.n1691 0.000973118
R2139 P.n1704 P.n1703 0.000973118
R2140 P.n3310 P.n3309 0.000973118
R2141 P.n2883 P.n2865 0.000956853
R2142 P.n2873 P.n2872 0.000956853
R2143 P.n3367 P.n3350 0.000956853
R2144 P.n3357 P.n3356 0.000956853
R2145 P.n2884 P.n2837 0.000956853
R2146 P.n2896 P.n2895 0.000956853
R2147 P.n2909 P.n2908 0.000956853
R2148 P.n2904 P.n2903 0.000956853
R2149 P.n3368 P.n3339 0.000956853
R2150 P.n3380 P.n3379 0.000956853
R2151 P.n3392 P.n3391 0.000956853
R2152 P.n3387 P.n3386 0.000956853
R2153 P.n2804 P.n2803 0.000956853
R2154 P.n3410 P.n3409 0.000956853
R2155 P.n2801 P.n2800 0.000956853
R2156 P.n2751 P.n2750 0.000956853
R2157 P.n2317 P.n2299 0.000956853
R2158 P.n2307 P.n2306 0.000956853
R2159 P.n2407 P.n2390 0.000956853
R2160 P.n2397 P.n2396 0.000956853
R2161 P.n2318 P.n2271 0.000956853
R2162 P.n2330 P.n2329 0.000956853
R2163 P.n2343 P.n2342 0.000956853
R2164 P.n2338 P.n2337 0.000956853
R2165 P.n2408 P.n2379 0.000956853
R2166 P.n2420 P.n2419 0.000956853
R2167 P.n2432 P.n2431 0.000956853
R2168 P.n2427 P.n2426 0.000956853
R2169 P.n3520 P.n3519 0.000956853
R2170 P.n2208 P.n2207 0.000956853
R2171 P.n2445 P.n2444 0.000956853
R2172 P.n2216 P.n2215 0.000956853
R2173 P.n3654 P.n3636 0.000956853
R2174 P.n3644 P.n3643 0.000956853
R2175 P.n2082 P.n2065 0.000956853
R2176 P.n2072 P.n2071 0.000956853
R2177 P.n3655 P.n3608 0.000956853
R2178 P.n3667 P.n3666 0.000956853
R2179 P.n3680 P.n3679 0.000956853
R2180 P.n3675 P.n3674 0.000956853
R2181 P.n2083 P.n2054 0.000956853
R2182 P.n2095 P.n2094 0.000956853
R2183 P.n2107 P.n2106 0.000956853
R2184 P.n2102 P.n2101 0.000956853
R2185 P.n2179 P.n2178 0.000956853
R2186 P.n2129 P.n2128 0.000956853
R2187 P.n2163 P.n2162 0.000956853
R2188 P.n2118 P.n2117 0.000956853
R2189 P.n2596 P.n2578 0.000956853
R2190 P.n2586 P.n2585 0.000956853
R2191 P.n2680 P.n2663 0.000956853
R2192 P.n2670 P.n2669 0.000956853
R2193 P.n2597 P.n2550 0.000956853
R2194 P.n2609 P.n2608 0.000956853
R2195 P.n2622 P.n2621 0.000956853
R2196 P.n2617 P.n2616 0.000956853
R2197 P.n2681 P.n2652 0.000956853
R2198 P.n2693 P.n2692 0.000956853
R2199 P.n2705 P.n2704 0.000956853
R2200 P.n2700 P.n2699 0.000956853
R2201 P.n3463 P.n3462 0.000956853
R2202 P.n2473 P.n2472 0.000956853
R2203 P.n2715 P.n2714 0.000956853
R2204 P.n2481 P.n2480 0.000956853
R2205 P.n3025 P.n3007 0.000956853
R2206 P.n3015 P.n3014 0.000956853
R2207 P.n3209 P.n3192 0.000956853
R2208 P.n3199 P.n3198 0.000956853
R2209 P.n3026 P.n2979 0.000956853
R2210 P.n3038 P.n3037 0.000956853
R2211 P.n3051 P.n3050 0.000956853
R2212 P.n3046 P.n3045 0.000956853
R2213 P.n3210 P.n3181 0.000956853
R2214 P.n3222 P.n3221 0.000956853
R2215 P.n3234 P.n3233 0.000956853
R2216 P.n3229 P.n3228 0.000956853
R2217 P.n2955 P.n2954 0.000956853
R2218 P.n3068 P.n3067 0.000956853
R2219 P.n3058 P.n3057 0.000956853
R2220 P.n3156 P.n3155 0.000956853
R2221 P.n3250 P.n3249 0.000956853
R2222 P.n3240 P.n3239 0.000956853
R2223 P.n1366 P.n1365 0.000951613
R2224 P.n1929 P.n1911 0.000941609
R2225 P.n1919 P.n1918 0.000941609
R2226 P.n1801 P.n1784 0.000941609
R2227 P.n1791 P.n1790 0.000941609
R2228 P.n1930 P.n1883 0.000941609
R2229 P.n1942 P.n1941 0.000941609
R2230 P.n1955 P.n1954 0.000941609
R2231 P.n1950 P.n1949 0.000941609
R2232 P.n1802 P.n1773 0.000941609
R2233 P.n1814 P.n1813 0.000941609
R2234 P.n1826 P.n1825 0.000941609
R2235 P.n1821 P.n1820 0.000941609
R2236 P.n1987 P.n1986 0.000941609
R2237 P.n1965 P.n1964 0.000941609
R2238 P.n1858 P.n1857 0.000941609
R2239 P.n1835 P.n1834 0.000941609
R2240 P.n1491 P.n1473 0.000941609
R2241 P.n1481 P.n1480 0.000941609
R2242 P.n1602 P.n1585 0.000941609
R2243 P.n1592 P.n1591 0.000941609
R2244 P.n1492 P.n1445 0.000941609
R2245 P.n1504 P.n1503 0.000941609
R2246 P.n1517 P.n1516 0.000941609
R2247 P.n1512 P.n1511 0.000941609
R2248 P.n1603 P.n1574 0.000941609
R2249 P.n1615 P.n1614 0.000941609
R2250 P.n1627 P.n1626 0.000941609
R2251 P.n1622 P.n1621 0.000941609
R2252 P.n1540 P.n1539 0.000941609
R2253 P.n1415 P.n1414 0.000941609
R2254 P.n1659 P.n1658 0.000941609
R2255 P.n1636 P.n1635 0.000941609
R2256 P.n1176 P.n1158 0.000941609
R2257 P.n1166 P.n1165 0.000941609
R2258 P.n1254 P.n1237 0.000941609
R2259 P.n1244 P.n1243 0.000941609
R2260 P.n1177 P.n1130 0.000941609
R2261 P.n1189 P.n1188 0.000941609
R2262 P.n1202 P.n1201 0.000941609
R2263 P.n1197 P.n1196 0.000941609
R2264 P.n1255 P.n1226 0.000941609
R2265 P.n1267 P.n1266 0.000941609
R2266 P.n1279 P.n1278 0.000941609
R2267 P.n1274 P.n1273 0.000941609
R2268 P.n1324 P.n1323 0.000941609
R2269 P.n1100 P.n1099 0.000941609
R2270 P.n1310 P.n1309 0.000941609
R2271 P.n1288 P.n1287 0.000941609
R2272 P.n972 P.n954 0.000941609
R2273 P.n962 P.n961 0.000941609
R2274 P.n845 P.n828 0.000941609
R2275 P.n835 P.n834 0.000941609
R2276 P.n973 P.n926 0.000941609
R2277 P.n985 P.n984 0.000941609
R2278 P.n998 P.n997 0.000941609
R2279 P.n993 P.n992 0.000941609
R2280 P.n846 P.n817 0.000941609
R2281 P.n858 P.n857 0.000941609
R2282 P.n870 P.n869 0.000941609
R2283 P.n865 P.n864 0.000941609
R2284 P.n1031 P.n1030 0.000941609
R2285 P.n1008 P.n1007 0.000941609
R2286 P.n893 P.n892 0.000941609
R2287 P.n794 P.n793 0.000941609
R2288 P.n256 P.n238 0.000941609
R2289 P.n246 P.n245 0.000941609
R2290 P.n161 P.n144 0.000941609
R2291 P.n151 P.n150 0.000941609
R2292 P.n257 P.n210 0.000941609
R2293 P.n269 P.n268 0.000941609
R2294 P.n282 P.n281 0.000941609
R2295 P.n277 P.n276 0.000941609
R2296 P.n162 P.n133 0.000941609
R2297 P.n174 P.n173 0.000941609
R2298 P.n186 P.n185 0.000941609
R2299 P.n181 P.n180 0.000941609
R2300 P.n362 P.n361 0.000941609
R2301 P.n323 P.n322 0.000941609
R2302 P.n596 P.n578 0.000941609
R2303 P.n586 P.n585 0.000941609
R2304 P.n476 P.n459 0.000941609
R2305 P.n466 P.n465 0.000941609
R2306 P.n597 P.n550 0.000941609
R2307 P.n609 P.n608 0.000941609
R2308 P.n622 P.n621 0.000941609
R2309 P.n617 P.n616 0.000941609
R2310 P.n477 P.n448 0.000941609
R2311 P.n489 P.n488 0.000941609
R2312 P.n501 P.n500 0.000941609
R2313 P.n496 P.n495 0.000941609
R2314 P.n425 P.n424 0.000941609
R2315 P.n689 P.n688 0.000941609
R2316 P.n61 P.n60 0.000941609
R2317 P.n648 P.n647 0.000941609
R2318 P.n3089 P.n3088 0.000930108
R2319 P.n3134 P.n3133 0.000930108
R2320 P.n721 P.n720 0.000930108
R2321 P.n732 P.n731 0.000930108
R2322 P.n1356 P.n1355 0.000930108
R2323 P.n3480 P.n3479 0.000930108
R2324 P.n3471 P.n3470 0.000930108
R2325 P.n3470 P.n3469 0.000930108
R2326 P.n3467 P.n3466 0.000930108
R2327 P.n3465 P.n3453 0.000930108
R2328 P.n3453 P.n3452 0.000930108
R2329 P.n3452 P.n3451 0.000930108
R2330 P.n3434 P.n3433 0.000930108
R2331 P.n3292 P.n3286 0.000930108
R2332 P.n639 P.n638 0.000908602
R2333 P.n654 P.n641 0.000908602
R2334 P.n728 P.n727 0.000908602
R2335 P.n1294 P.n1094 0.000908602
R2336 P.n1696 P.n1695 0.000908602
R2337 P.n3479 P.n3478 0.000908602
R2338 P.n3466 P.n3465 0.000908602
R2339 P.n3295 P.n3294 0.000908602
R2340 P.n2935 P.n2934 0.000887097
R2341 P.n3085 P.n3084 0.000887097
R2342 P.n3271 P.n3270 0.000887097
R2343 P.n3266 P.n3137 0.000887097
R2344 P.n1402 P.n1401 0.000887097
R2345 P.n3564 P.n3563 0.000887097
R2346 P.n3468 P.n3467 0.000887097
R2347 P.n106 P.n105 0.000865591
R2348 P.n429 P.n428 0.000865591
R2349 P.n734 P.n733 0.000865591
R2350 P.n740 P.n739 0.000865591
R2351 P.n744 P.n743 0.000865591
R2352 P.n1067 P.n1066 0.000865591
R2353 P.n1691 P.n1690 0.000865591
R2354 P.n1701 P.n1700 0.000865591
R2355 P.n1703 P.n1702 0.000865591
R2356 P.n1705 P.n1704 0.000865591
R2357 P.n1707 P.n1706 0.000865591
R2358 P.n1709 P.n1708 0.000865591
R2359 P.n1710 P.n1709 0.000865591
R2360 P.n1748 P.n1747 0.000865591
R2361 P.n3513 P.n3512 0.000865591
R2362 P.n3473 P.n3472 0.000865591
R2363 P.n3450 P.n3449 0.000865591
R2364 P.n3448 P.n3447 0.000865591
R2365 P.n3311 P.n3310 0.000865591
R2366 P.n2851 P.n2850 0.000865482
R2367 P.n2841 P.n2840 0.000865482
R2368 P.n2876 P.n2875 0.000865482
R2369 P.n2874 P.n2873 0.000865482
R2370 P.n2872 P.n2871 0.000865482
R2371 P.n2868 P.n2867 0.000865482
R2372 P.n3360 P.n3359 0.000865482
R2373 P.n3358 P.n3357 0.000865482
R2374 P.n3356 P.n3355 0.000865482
R2375 P.n3352 P.n3351 0.000865482
R2376 P.n2822 P.n2821 0.000865482
R2377 P.n2826 P.n2825 0.000865482
R2378 P.n2828 P.n2827 0.000865482
R2379 P.n2830 P.n2829 0.000865482
R2380 P.n2834 P.n2833 0.000865482
R2381 P.n2835 P.n2834 0.000865482
R2382 P.n2837 P.n2836 0.000865482
R2383 P.n2885 P.n2884 0.000865482
R2384 P.n2886 P.n2885 0.000865482
R2385 P.n2889 P.n2888 0.000865482
R2386 P.n2890 P.n2889 0.000865482
R2387 P.n2891 P.n2890 0.000865482
R2388 P.n2893 P.n2892 0.000865482
R2389 P.n2895 P.n2894 0.000865482
R2390 P.n2897 P.n2896 0.000865482
R2391 P.n2898 P.n2897 0.000865482
R2392 P.n2910 P.n2909 0.000865482
R2393 P.n2908 P.n2907 0.000865482
R2394 P.n2903 P.n2902 0.000865482
R2395 P.n2902 P.n2901 0.000865482
R2396 P.n2900 P.n2899 0.000865482
R2397 P.n3322 P.n3321 0.000865482
R2398 P.n3324 P.n3323 0.000865482
R2399 P.n3328 P.n3327 0.000865482
R2400 P.n3330 P.n3329 0.000865482
R2401 P.n3332 P.n3331 0.000865482
R2402 P.n3336 P.n3335 0.000865482
R2403 P.n3337 P.n3336 0.000865482
R2404 P.n3339 P.n3338 0.000865482
R2405 P.n3369 P.n3368 0.000865482
R2406 P.n3370 P.n3369 0.000865482
R2407 P.n3373 P.n3372 0.000865482
R2408 P.n3374 P.n3373 0.000865482
R2409 P.n3375 P.n3374 0.000865482
R2410 P.n3377 P.n3376 0.000865482
R2411 P.n3379 P.n3378 0.000865482
R2412 P.n3381 P.n3380 0.000865482
R2413 P.n3382 P.n3381 0.000865482
R2414 P.n3393 P.n3392 0.000865482
R2415 P.n3391 P.n3390 0.000865482
R2416 P.n3386 P.n3385 0.000865482
R2417 P.n3385 P.n3384 0.000865482
R2418 P.n3289 P.n3288 0.000865482
R2419 P.n2764 P.n2763 0.000865482
R2420 P.n2759 P.n2758 0.000865482
R2421 P.n2758 P.n2757 0.000865482
R2422 P.n2757 P.n2756 0.000865482
R2423 P.n2755 P.n2754 0.000865482
R2424 P.n2815 P.n2814 0.000865482
R2425 P.n2817 P.n2816 0.000865482
R2426 P.n3411 P.n3410 0.000865482
R2427 P.n3409 P.n3408 0.000865482
R2428 P.n3408 P.n3407 0.000865482
R2429 P.n3406 P.n3405 0.000865482
R2430 P.n2922 P.n2921 0.000865482
R2431 P.n2778 P.n2777 0.000865482
R2432 P.n2773 P.n2772 0.000865482
R2433 P.n2772 P.n2771 0.000865482
R2434 P.n2771 P.n2770 0.000865482
R2435 P.n2769 P.n2768 0.000865482
R2436 P.n3316 P.n3315 0.000865482
R2437 P.n3318 P.n3317 0.000865482
R2438 P.n2752 P.n2751 0.000865482
R2439 P.n2750 P.n2749 0.000865482
R2440 P.n2749 P.n2748 0.000865482
R2441 P.n2285 P.n2284 0.000865482
R2442 P.n2275 P.n2274 0.000865482
R2443 P.n2310 P.n2309 0.000865482
R2444 P.n2308 P.n2307 0.000865482
R2445 P.n2306 P.n2305 0.000865482
R2446 P.n2302 P.n2301 0.000865482
R2447 P.n2400 P.n2399 0.000865482
R2448 P.n2398 P.n2397 0.000865482
R2449 P.n2396 P.n2395 0.000865482
R2450 P.n2392 P.n2391 0.000865482
R2451 P.n2256 P.n2255 0.000865482
R2452 P.n2260 P.n2259 0.000865482
R2453 P.n2262 P.n2261 0.000865482
R2454 P.n2264 P.n2263 0.000865482
R2455 P.n2268 P.n2267 0.000865482
R2456 P.n2269 P.n2268 0.000865482
R2457 P.n2271 P.n2270 0.000865482
R2458 P.n2319 P.n2318 0.000865482
R2459 P.n2320 P.n2319 0.000865482
R2460 P.n2323 P.n2322 0.000865482
R2461 P.n2324 P.n2323 0.000865482
R2462 P.n2325 P.n2324 0.000865482
R2463 P.n2327 P.n2326 0.000865482
R2464 P.n2329 P.n2328 0.000865482
R2465 P.n2331 P.n2330 0.000865482
R2466 P.n2332 P.n2331 0.000865482
R2467 P.n2344 P.n2343 0.000865482
R2468 P.n2342 P.n2341 0.000865482
R2469 P.n2337 P.n2336 0.000865482
R2470 P.n2336 P.n2335 0.000865482
R2471 P.n2334 P.n2333 0.000865482
R2472 P.n2362 P.n2361 0.000865482
R2473 P.n2364 P.n2363 0.000865482
R2474 P.n2368 P.n2367 0.000865482
R2475 P.n2370 P.n2369 0.000865482
R2476 P.n2372 P.n2371 0.000865482
R2477 P.n2376 P.n2375 0.000865482
R2478 P.n2377 P.n2376 0.000865482
R2479 P.n2379 P.n2378 0.000865482
R2480 P.n2409 P.n2408 0.000865482
R2481 P.n2410 P.n2409 0.000865482
R2482 P.n2413 P.n2412 0.000865482
R2483 P.n2414 P.n2413 0.000865482
R2484 P.n2415 P.n2414 0.000865482
R2485 P.n2417 P.n2416 0.000865482
R2486 P.n2419 P.n2418 0.000865482
R2487 P.n2421 P.n2420 0.000865482
R2488 P.n2422 P.n2421 0.000865482
R2489 P.n2433 P.n2432 0.000865482
R2490 P.n2431 P.n2430 0.000865482
R2491 P.n2426 P.n2425 0.000865482
R2492 P.n2425 P.n2424 0.000865482
R2493 P.n2460 P.n2459 0.000865482
R2494 P.n2229 P.n2228 0.000865482
R2495 P.n2225 P.n2224 0.000865482
R2496 P.n2224 P.n2223 0.000865482
R2497 P.n2223 P.n2222 0.000865482
R2498 P.n2221 P.n2220 0.000865482
R2499 P.n2249 P.n2248 0.000865482
R2500 P.n2251 P.n2250 0.000865482
R2501 P.n2209 P.n2208 0.000865482
R2502 P.n2207 P.n2206 0.000865482
R2503 P.n2206 P.n2205 0.000865482
R2504 P.n2204 P.n2203 0.000865482
R2505 P.n2465 P.n2464 0.000865482
R2506 P.n2242 P.n2241 0.000865482
R2507 P.n2238 P.n2237 0.000865482
R2508 P.n2237 P.n2236 0.000865482
R2509 P.n2236 P.n2235 0.000865482
R2510 P.n2234 P.n2233 0.000865482
R2511 P.n2356 P.n2355 0.000865482
R2512 P.n2358 P.n2357 0.000865482
R2513 P.n2217 P.n2216 0.000865482
R2514 P.n2215 P.n2214 0.000865482
R2515 P.n2214 P.n2213 0.000865482
R2516 P.n3622 P.n3621 0.000865482
R2517 P.n3612 P.n3611 0.000865482
R2518 P.n3647 P.n3646 0.000865482
R2519 P.n3645 P.n3644 0.000865482
R2520 P.n3643 P.n3642 0.000865482
R2521 P.n3639 P.n3638 0.000865482
R2522 P.n2075 P.n2074 0.000865482
R2523 P.n2073 P.n2072 0.000865482
R2524 P.n2071 P.n2070 0.000865482
R2525 P.n2067 P.n2066 0.000865482
R2526 P.n3593 P.n3592 0.000865482
R2527 P.n3597 P.n3596 0.000865482
R2528 P.n3599 P.n3598 0.000865482
R2529 P.n3601 P.n3600 0.000865482
R2530 P.n3605 P.n3604 0.000865482
R2531 P.n3606 P.n3605 0.000865482
R2532 P.n3608 P.n3607 0.000865482
R2533 P.n3656 P.n3655 0.000865482
R2534 P.n3657 P.n3656 0.000865482
R2535 P.n3660 P.n3659 0.000865482
R2536 P.n3661 P.n3660 0.000865482
R2537 P.n3662 P.n3661 0.000865482
R2538 P.n3664 P.n3663 0.000865482
R2539 P.n3666 P.n3665 0.000865482
R2540 P.n3668 P.n3667 0.000865482
R2541 P.n3669 P.n3668 0.000865482
R2542 P.n3681 P.n3680 0.000865482
R2543 P.n3679 P.n3678 0.000865482
R2544 P.n3674 P.n3673 0.000865482
R2545 P.n3673 P.n3672 0.000865482
R2546 P.n3671 P.n3670 0.000865482
R2547 P.n2037 P.n2036 0.000865482
R2548 P.n2039 P.n2038 0.000865482
R2549 P.n2043 P.n2042 0.000865482
R2550 P.n2045 P.n2044 0.000865482
R2551 P.n2047 P.n2046 0.000865482
R2552 P.n2051 P.n2050 0.000865482
R2553 P.n2052 P.n2051 0.000865482
R2554 P.n2054 P.n2053 0.000865482
R2555 P.n2084 P.n2083 0.000865482
R2556 P.n2085 P.n2084 0.000865482
R2557 P.n2088 P.n2087 0.000865482
R2558 P.n2089 P.n2088 0.000865482
R2559 P.n2090 P.n2089 0.000865482
R2560 P.n2092 P.n2091 0.000865482
R2561 P.n2094 P.n2093 0.000865482
R2562 P.n2096 P.n2095 0.000865482
R2563 P.n2097 P.n2096 0.000865482
R2564 P.n2108 P.n2107 0.000865482
R2565 P.n2106 P.n2105 0.000865482
R2566 P.n2101 P.n2100 0.000865482
R2567 P.n2100 P.n2099 0.000865482
R2568 P.n3570 P.n3569 0.000865482
R2569 P.n2150 P.n2149 0.000865482
R2570 P.n2158 P.n2157 0.000865482
R2571 P.n2157 P.n2156 0.000865482
R2572 P.n2156 P.n2155 0.000865482
R2573 P.n2154 P.n2153 0.000865482
R2574 P.n3685 P.n3684 0.000865482
R2575 P.n3687 P.n3686 0.000865482
R2576 P.n2130 P.n2129 0.000865482
R2577 P.n2128 P.n2127 0.000865482
R2578 P.n2127 P.n2126 0.000865482
R2579 P.n2125 P.n2124 0.000865482
R2580 P.n2187 P.n2186 0.000865482
R2581 P.n2136 P.n2135 0.000865482
R2582 P.n2144 P.n2143 0.000865482
R2583 P.n2143 P.n2142 0.000865482
R2584 P.n2142 P.n2141 0.000865482
R2585 P.n2140 P.n2139 0.000865482
R2586 P.n2031 P.n2030 0.000865482
R2587 P.n2033 P.n2032 0.000865482
R2588 P.n2119 P.n2118 0.000865482
R2589 P.n2117 P.n2116 0.000865482
R2590 P.n2116 P.n2115 0.000865482
R2591 P.n2564 P.n2563 0.000865482
R2592 P.n2554 P.n2553 0.000865482
R2593 P.n2589 P.n2588 0.000865482
R2594 P.n2587 P.n2586 0.000865482
R2595 P.n2585 P.n2584 0.000865482
R2596 P.n2581 P.n2580 0.000865482
R2597 P.n2673 P.n2672 0.000865482
R2598 P.n2671 P.n2670 0.000865482
R2599 P.n2669 P.n2668 0.000865482
R2600 P.n2665 P.n2664 0.000865482
R2601 P.n2535 P.n2534 0.000865482
R2602 P.n2539 P.n2538 0.000865482
R2603 P.n2541 P.n2540 0.000865482
R2604 P.n2543 P.n2542 0.000865482
R2605 P.n2547 P.n2546 0.000865482
R2606 P.n2548 P.n2547 0.000865482
R2607 P.n2550 P.n2549 0.000865482
R2608 P.n2598 P.n2597 0.000865482
R2609 P.n2599 P.n2598 0.000865482
R2610 P.n2602 P.n2601 0.000865482
R2611 P.n2603 P.n2602 0.000865482
R2612 P.n2604 P.n2603 0.000865482
R2613 P.n2606 P.n2605 0.000865482
R2614 P.n2608 P.n2607 0.000865482
R2615 P.n2610 P.n2609 0.000865482
R2616 P.n2611 P.n2610 0.000865482
R2617 P.n2623 P.n2622 0.000865482
R2618 P.n2621 P.n2620 0.000865482
R2619 P.n2616 P.n2615 0.000865482
R2620 P.n2615 P.n2614 0.000865482
R2621 P.n2613 P.n2612 0.000865482
R2622 P.n2635 P.n2634 0.000865482
R2623 P.n2637 P.n2636 0.000865482
R2624 P.n2641 P.n2640 0.000865482
R2625 P.n2643 P.n2642 0.000865482
R2626 P.n2645 P.n2644 0.000865482
R2627 P.n2649 P.n2648 0.000865482
R2628 P.n2650 P.n2649 0.000865482
R2629 P.n2652 P.n2651 0.000865482
R2630 P.n2682 P.n2681 0.000865482
R2631 P.n2683 P.n2682 0.000865482
R2632 P.n2686 P.n2685 0.000865482
R2633 P.n2687 P.n2686 0.000865482
R2634 P.n2688 P.n2687 0.000865482
R2635 P.n2690 P.n2689 0.000865482
R2636 P.n2692 P.n2691 0.000865482
R2637 P.n2694 P.n2693 0.000865482
R2638 P.n2695 P.n2694 0.000865482
R2639 P.n2706 P.n2705 0.000865482
R2640 P.n2704 P.n2703 0.000865482
R2641 P.n2699 P.n2698 0.000865482
R2642 P.n2698 P.n2697 0.000865482
R2643 P.n2725 P.n2724 0.000865482
R2644 P.n2487 P.n2486 0.000865482
R2645 P.n2495 P.n2494 0.000865482
R2646 P.n2494 P.n2493 0.000865482
R2647 P.n2493 P.n2492 0.000865482
R2648 P.n2491 P.n2490 0.000865482
R2649 P.n2528 P.n2527 0.000865482
R2650 P.n2530 P.n2529 0.000865482
R2651 P.n2474 P.n2473 0.000865482
R2652 P.n2472 P.n2471 0.000865482
R2653 P.n2471 P.n2470 0.000865482
R2654 P.n2469 P.n2468 0.000865482
R2655 P.n2735 P.n2734 0.000865482
R2656 P.n2500 P.n2499 0.000865482
R2657 P.n2508 P.n2507 0.000865482
R2658 P.n2507 P.n2506 0.000865482
R2659 P.n2506 P.n2505 0.000865482
R2660 P.n2504 P.n2503 0.000865482
R2661 P.n2629 P.n2628 0.000865482
R2662 P.n2631 P.n2630 0.000865482
R2663 P.n2482 P.n2481 0.000865482
R2664 P.n2480 P.n2479 0.000865482
R2665 P.n2479 P.n2478 0.000865482
R2666 P.n2993 P.n2992 0.000865482
R2667 P.n2983 P.n2982 0.000865482
R2668 P.n3018 P.n3017 0.000865482
R2669 P.n3016 P.n3015 0.000865482
R2670 P.n3014 P.n3013 0.000865482
R2671 P.n3010 P.n3009 0.000865482
R2672 P.n3202 P.n3201 0.000865482
R2673 P.n3200 P.n3199 0.000865482
R2674 P.n3198 P.n3197 0.000865482
R2675 P.n3194 P.n3193 0.000865482
R2676 P.n2964 P.n2963 0.000865482
R2677 P.n2968 P.n2967 0.000865482
R2678 P.n2970 P.n2969 0.000865482
R2679 P.n2972 P.n2971 0.000865482
R2680 P.n2976 P.n2975 0.000865482
R2681 P.n2977 P.n2976 0.000865482
R2682 P.n2979 P.n2978 0.000865482
R2683 P.n3027 P.n3026 0.000865482
R2684 P.n3028 P.n3027 0.000865482
R2685 P.n3031 P.n3030 0.000865482
R2686 P.n3032 P.n3031 0.000865482
R2687 P.n3033 P.n3032 0.000865482
R2688 P.n3035 P.n3034 0.000865482
R2689 P.n3037 P.n3036 0.000865482
R2690 P.n3039 P.n3038 0.000865482
R2691 P.n3040 P.n3039 0.000865482
R2692 P.n3052 P.n3051 0.000865482
R2693 P.n3050 P.n3049 0.000865482
R2694 P.n3045 P.n3044 0.000865482
R2695 P.n3044 P.n3043 0.000865482
R2696 P.n3042 P.n3041 0.000865482
R2697 P.n3164 P.n3163 0.000865482
R2698 P.n3166 P.n3165 0.000865482
R2699 P.n3170 P.n3169 0.000865482
R2700 P.n3172 P.n3171 0.000865482
R2701 P.n3174 P.n3173 0.000865482
R2702 P.n3178 P.n3177 0.000865482
R2703 P.n3179 P.n3178 0.000865482
R2704 P.n3181 P.n3180 0.000865482
R2705 P.n3211 P.n3210 0.000865482
R2706 P.n3212 P.n3211 0.000865482
R2707 P.n3215 P.n3214 0.000865482
R2708 P.n3216 P.n3215 0.000865482
R2709 P.n3217 P.n3216 0.000865482
R2710 P.n3219 P.n3218 0.000865482
R2711 P.n3221 P.n3220 0.000865482
R2712 P.n3223 P.n3222 0.000865482
R2713 P.n3224 P.n3223 0.000865482
R2714 P.n3235 P.n3234 0.000865482
R2715 P.n3233 P.n3232 0.000865482
R2716 P.n3228 P.n3227 0.000865482
R2717 P.n3227 P.n3226 0.000865482
R2718 P.n2946 P.n2945 0.000865482
R2719 P.n2948 P.n2947 0.000865482
R2720 P.n2960 P.n2959 0.000865482
R2721 P.n3080 P.n3079 0.000865482
R2722 P.n3079 P.n3078 0.000865482
R2723 P.n3078 P.n3077 0.000865482
R2724 P.n3076 P.n3075 0.000865482
R2725 P.n3072 P.n3071 0.000865482
R2726 P.n3070 P.n3069 0.000865482
R2727 P.n3059 P.n3058 0.000865482
R2728 P.n3057 P.n3056 0.000865482
R2729 P.n3056 P.n3055 0.000865482
R2730 P.n3054 P.n3053 0.000865482
R2731 P.n3147 P.n3146 0.000865482
R2732 P.n3149 P.n3148 0.000865482
R2733 P.n3161 P.n3160 0.000865482
R2734 P.n3262 P.n3261 0.000865482
R2735 P.n3261 P.n3260 0.000865482
R2736 P.n3260 P.n3259 0.000865482
R2737 P.n3258 P.n3257 0.000865482
R2738 P.n3254 P.n3253 0.000865482
R2739 P.n3252 P.n3251 0.000865482
R2740 P.n3241 P.n3240 0.000865482
R2741 P.n3239 P.n3238 0.000865482
R2742 P.n3238 P.n3237 0.000865482
R2743 P.n1897 P.n1896 0.000853288
R2744 P.n1887 P.n1886 0.000853288
R2745 P.n1922 P.n1921 0.000853288
R2746 P.n1920 P.n1919 0.000853288
R2747 P.n1918 P.n1917 0.000853288
R2748 P.n1914 P.n1913 0.000853288
R2749 P.n1794 P.n1793 0.000853288
R2750 P.n1792 P.n1791 0.000853288
R2751 P.n1790 P.n1789 0.000853288
R2752 P.n1786 P.n1785 0.000853288
R2753 P.n1868 P.n1867 0.000853288
R2754 P.n1872 P.n1871 0.000853288
R2755 P.n1874 P.n1873 0.000853288
R2756 P.n1876 P.n1875 0.000853288
R2757 P.n1880 P.n1879 0.000853288
R2758 P.n1881 P.n1880 0.000853288
R2759 P.n1883 P.n1882 0.000853288
R2760 P.n1931 P.n1930 0.000853288
R2761 P.n1932 P.n1931 0.000853288
R2762 P.n1935 P.n1934 0.000853288
R2763 P.n1936 P.n1935 0.000853288
R2764 P.n1937 P.n1936 0.000853288
R2765 P.n1939 P.n1938 0.000853288
R2766 P.n1941 P.n1940 0.000853288
R2767 P.n1943 P.n1942 0.000853288
R2768 P.n1944 P.n1943 0.000853288
R2769 P.n1956 P.n1955 0.000853288
R2770 P.n1954 P.n1953 0.000853288
R2771 P.n1949 P.n1948 0.000853288
R2772 P.n1948 P.n1947 0.000853288
R2773 P.n1946 P.n1945 0.000853288
R2774 P.n1756 P.n1755 0.000853288
R2775 P.n1758 P.n1757 0.000853288
R2776 P.n1762 P.n1761 0.000853288
R2777 P.n1764 P.n1763 0.000853288
R2778 P.n1766 P.n1765 0.000853288
R2779 P.n1770 P.n1769 0.000853288
R2780 P.n1771 P.n1770 0.000853288
R2781 P.n1773 P.n1772 0.000853288
R2782 P.n1803 P.n1802 0.000853288
R2783 P.n1804 P.n1803 0.000853288
R2784 P.n1807 P.n1806 0.000853288
R2785 P.n1808 P.n1807 0.000853288
R2786 P.n1809 P.n1808 0.000853288
R2787 P.n1811 P.n1810 0.000853288
R2788 P.n1813 P.n1812 0.000853288
R2789 P.n1815 P.n1814 0.000853288
R2790 P.n1816 P.n1815 0.000853288
R2791 P.n1827 P.n1826 0.000853288
R2792 P.n1825 P.n1824 0.000853288
R2793 P.n1820 P.n1819 0.000853288
R2794 P.n1819 P.n1818 0.000853288
R2795 P.n2007 P.n2006 0.000853288
R2796 P.n2005 P.n2004 0.000853288
R2797 P.n1992 P.n1991 0.000853288
R2798 P.n1998 P.n1997 0.000853288
R2799 P.n1997 P.n1996 0.000853288
R2800 P.n1996 P.n1995 0.000853288
R2801 P.n1994 P.n1993 0.000853288
R2802 P.n1724 P.n1723 0.000853288
R2803 P.n1726 P.n1725 0.000853288
R2804 P.n1966 P.n1965 0.000853288
R2805 P.n1964 P.n1963 0.000853288
R2806 P.n1963 P.n1962 0.000853288
R2807 P.n1961 P.n1960 0.000853288
R2808 P.n1976 P.n1975 0.000853288
R2809 P.n1974 P.n1973 0.000853288
R2810 P.n1863 P.n1862 0.000853288
R2811 P.n1847 P.n1846 0.000853288
R2812 P.n1846 P.n1845 0.000853288
R2813 P.n1845 P.n1844 0.000853288
R2814 P.n1843 P.n1842 0.000853288
R2815 P.n1714 P.n1713 0.000853288
R2816 P.n1716 P.n1715 0.000853288
R2817 P.n1836 P.n1835 0.000853288
R2818 P.n1834 P.n1833 0.000853288
R2819 P.n1833 P.n1832 0.000853288
R2820 P.n1459 P.n1458 0.000853288
R2821 P.n1449 P.n1448 0.000853288
R2822 P.n1484 P.n1483 0.000853288
R2823 P.n1482 P.n1481 0.000853288
R2824 P.n1480 P.n1479 0.000853288
R2825 P.n1476 P.n1475 0.000853288
R2826 P.n1595 P.n1594 0.000853288
R2827 P.n1593 P.n1592 0.000853288
R2828 P.n1591 P.n1590 0.000853288
R2829 P.n1587 P.n1586 0.000853288
R2830 P.n1430 P.n1429 0.000853288
R2831 P.n1434 P.n1433 0.000853288
R2832 P.n1436 P.n1435 0.000853288
R2833 P.n1438 P.n1437 0.000853288
R2834 P.n1442 P.n1441 0.000853288
R2835 P.n1443 P.n1442 0.000853288
R2836 P.n1445 P.n1444 0.000853288
R2837 P.n1493 P.n1492 0.000853288
R2838 P.n1494 P.n1493 0.000853288
R2839 P.n1497 P.n1496 0.000853288
R2840 P.n1498 P.n1497 0.000853288
R2841 P.n1499 P.n1498 0.000853288
R2842 P.n1501 P.n1500 0.000853288
R2843 P.n1503 P.n1502 0.000853288
R2844 P.n1505 P.n1504 0.000853288
R2845 P.n1506 P.n1505 0.000853288
R2846 P.n1518 P.n1517 0.000853288
R2847 P.n1516 P.n1515 0.000853288
R2848 P.n1511 P.n1510 0.000853288
R2849 P.n1510 P.n1509 0.000853288
R2850 P.n1508 P.n1507 0.000853288
R2851 P.n1557 P.n1556 0.000853288
R2852 P.n1559 P.n1558 0.000853288
R2853 P.n1563 P.n1562 0.000853288
R2854 P.n1565 P.n1564 0.000853288
R2855 P.n1567 P.n1566 0.000853288
R2856 P.n1571 P.n1570 0.000853288
R2857 P.n1572 P.n1571 0.000853288
R2858 P.n1574 P.n1573 0.000853288
R2859 P.n1604 P.n1603 0.000853288
R2860 P.n1605 P.n1604 0.000853288
R2861 P.n1608 P.n1607 0.000853288
R2862 P.n1609 P.n1608 0.000853288
R2863 P.n1610 P.n1609 0.000853288
R2864 P.n1612 P.n1611 0.000853288
R2865 P.n1614 P.n1613 0.000853288
R2866 P.n1616 P.n1615 0.000853288
R2867 P.n1617 P.n1616 0.000853288
R2868 P.n1628 P.n1627 0.000853288
R2869 P.n1626 P.n1625 0.000853288
R2870 P.n1621 P.n1620 0.000853288
R2871 P.n1620 P.n1619 0.000853288
R2872 P.n1671 P.n1670 0.000853288
R2873 P.n1669 P.n1668 0.000853288
R2874 P.n1545 P.n1544 0.000853288
R2875 P.n1529 P.n1528 0.000853288
R2876 P.n1528 P.n1527 0.000853288
R2877 P.n1527 P.n1526 0.000853288
R2878 P.n1525 P.n1524 0.000853288
R2879 P.n1423 P.n1422 0.000853288
R2880 P.n1425 P.n1424 0.000853288
R2881 P.n1416 P.n1415 0.000853288
R2882 P.n1414 P.n1413 0.000853288
R2883 P.n1413 P.n1412 0.000853288
R2884 P.n1411 P.n1410 0.000853288
R2885 P.n1679 P.n1678 0.000853288
R2886 P.n1677 P.n1676 0.000853288
R2887 P.n1664 P.n1663 0.000853288
R2888 P.n1648 P.n1647 0.000853288
R2889 P.n1647 P.n1646 0.000853288
R2890 P.n1646 P.n1645 0.000853288
R2891 P.n1644 P.n1643 0.000853288
R2892 P.n1551 P.n1550 0.000853288
R2893 P.n1553 P.n1552 0.000853288
R2894 P.n1637 P.n1636 0.000853288
R2895 P.n1635 P.n1634 0.000853288
R2896 P.n1634 P.n1633 0.000853288
R2897 P.n1144 P.n1143 0.000853288
R2898 P.n1134 P.n1133 0.000853288
R2899 P.n1169 P.n1168 0.000853288
R2900 P.n1167 P.n1166 0.000853288
R2901 P.n1165 P.n1164 0.000853288
R2902 P.n1161 P.n1160 0.000853288
R2903 P.n1247 P.n1246 0.000853288
R2904 P.n1245 P.n1244 0.000853288
R2905 P.n1243 P.n1242 0.000853288
R2906 P.n1239 P.n1238 0.000853288
R2907 P.n1115 P.n1114 0.000853288
R2908 P.n1119 P.n1118 0.000853288
R2909 P.n1121 P.n1120 0.000853288
R2910 P.n1123 P.n1122 0.000853288
R2911 P.n1127 P.n1126 0.000853288
R2912 P.n1128 P.n1127 0.000853288
R2913 P.n1130 P.n1129 0.000853288
R2914 P.n1178 P.n1177 0.000853288
R2915 P.n1179 P.n1178 0.000853288
R2916 P.n1182 P.n1181 0.000853288
R2917 P.n1183 P.n1182 0.000853288
R2918 P.n1184 P.n1183 0.000853288
R2919 P.n1186 P.n1185 0.000853288
R2920 P.n1188 P.n1187 0.000853288
R2921 P.n1190 P.n1189 0.000853288
R2922 P.n1191 P.n1190 0.000853288
R2923 P.n1203 P.n1202 0.000853288
R2924 P.n1201 P.n1200 0.000853288
R2925 P.n1196 P.n1195 0.000853288
R2926 P.n1195 P.n1194 0.000853288
R2927 P.n1193 P.n1192 0.000853288
R2928 P.n1209 P.n1208 0.000853288
R2929 P.n1211 P.n1210 0.000853288
R2930 P.n1215 P.n1214 0.000853288
R2931 P.n1217 P.n1216 0.000853288
R2932 P.n1219 P.n1218 0.000853288
R2933 P.n1223 P.n1222 0.000853288
R2934 P.n1224 P.n1223 0.000853288
R2935 P.n1226 P.n1225 0.000853288
R2936 P.n1256 P.n1255 0.000853288
R2937 P.n1257 P.n1256 0.000853288
R2938 P.n1260 P.n1259 0.000853288
R2939 P.n1261 P.n1260 0.000853288
R2940 P.n1262 P.n1261 0.000853288
R2941 P.n1264 P.n1263 0.000853288
R2942 P.n1266 P.n1265 0.000853288
R2943 P.n1268 P.n1267 0.000853288
R2944 P.n1269 P.n1268 0.000853288
R2945 P.n1280 P.n1279 0.000853288
R2946 P.n1278 P.n1277 0.000853288
R2947 P.n1273 P.n1272 0.000853288
R2948 P.n1272 P.n1271 0.000853288
R2949 P.n1352 P.n1351 0.000853288
R2950 P.n1350 P.n1349 0.000853288
R2951 P.n1329 P.n1328 0.000853288
R2952 P.n1335 P.n1334 0.000853288
R2953 P.n1334 P.n1333 0.000853288
R2954 P.n1333 P.n1332 0.000853288
R2955 P.n1331 P.n1330 0.000853288
R2956 P.n1108 P.n1107 0.000853288
R2957 P.n1110 P.n1109 0.000853288
R2958 P.n1101 P.n1100 0.000853288
R2959 P.n1099 P.n1098 0.000853288
R2960 P.n1098 P.n1097 0.000853288
R2961 P.n1096 P.n1095 0.000853288
R2962 P.n1345 P.n1344 0.000853288
R2963 P.n1343 P.n1342 0.000853288
R2964 P.n1315 P.n1314 0.000853288
R2965 P.n1300 P.n1299 0.000853288
R2966 P.n1299 P.n1298 0.000853288
R2967 P.n1298 P.n1297 0.000853288
R2968 P.n1296 P.n1295 0.000853288
R2969 P.n1071 P.n1070 0.000853288
R2970 P.n1073 P.n1072 0.000853288
R2971 P.n1289 P.n1288 0.000853288
R2972 P.n1287 P.n1286 0.000853288
R2973 P.n1286 P.n1285 0.000853288
R2974 P.n940 P.n939 0.000853288
R2975 P.n930 P.n929 0.000853288
R2976 P.n965 P.n964 0.000853288
R2977 P.n963 P.n962 0.000853288
R2978 P.n961 P.n960 0.000853288
R2979 P.n957 P.n956 0.000853288
R2980 P.n838 P.n837 0.000853288
R2981 P.n836 P.n835 0.000853288
R2982 P.n834 P.n833 0.000853288
R2983 P.n830 P.n829 0.000853288
R2984 P.n911 P.n910 0.000853288
R2985 P.n915 P.n914 0.000853288
R2986 P.n917 P.n916 0.000853288
R2987 P.n919 P.n918 0.000853288
R2988 P.n923 P.n922 0.000853288
R2989 P.n924 P.n923 0.000853288
R2990 P.n926 P.n925 0.000853288
R2991 P.n974 P.n973 0.000853288
R2992 P.n975 P.n974 0.000853288
R2993 P.n978 P.n977 0.000853288
R2994 P.n979 P.n978 0.000853288
R2995 P.n980 P.n979 0.000853288
R2996 P.n982 P.n981 0.000853288
R2997 P.n984 P.n983 0.000853288
R2998 P.n986 P.n985 0.000853288
R2999 P.n987 P.n986 0.000853288
R3000 P.n999 P.n998 0.000853288
R3001 P.n997 P.n996 0.000853288
R3002 P.n992 P.n991 0.000853288
R3003 P.n991 P.n990 0.000853288
R3004 P.n989 P.n988 0.000853288
R3005 P.n800 P.n799 0.000853288
R3006 P.n802 P.n801 0.000853288
R3007 P.n806 P.n805 0.000853288
R3008 P.n808 P.n807 0.000853288
R3009 P.n810 P.n809 0.000853288
R3010 P.n814 P.n813 0.000853288
R3011 P.n815 P.n814 0.000853288
R3012 P.n817 P.n816 0.000853288
R3013 P.n847 P.n846 0.000853288
R3014 P.n848 P.n847 0.000853288
R3015 P.n851 P.n850 0.000853288
R3016 P.n852 P.n851 0.000853288
R3017 P.n853 P.n852 0.000853288
R3018 P.n855 P.n854 0.000853288
R3019 P.n857 P.n856 0.000853288
R3020 P.n859 P.n858 0.000853288
R3021 P.n860 P.n859 0.000853288
R3022 P.n871 P.n870 0.000853288
R3023 P.n869 P.n868 0.000853288
R3024 P.n864 P.n863 0.000853288
R3025 P.n863 P.n862 0.000853288
R3026 P.n1044 P.n1043 0.000853288
R3027 P.n1042 P.n1041 0.000853288
R3028 P.n1036 P.n1035 0.000853288
R3029 P.n1020 P.n1019 0.000853288
R3030 P.n1019 P.n1018 0.000853288
R3031 P.n1018 P.n1017 0.000853288
R3032 P.n1016 P.n1015 0.000853288
R3033 P.n761 P.n760 0.000853288
R3034 P.n763 P.n762 0.000853288
R3035 P.n1009 P.n1008 0.000853288
R3036 P.n1007 P.n1006 0.000853288
R3037 P.n1006 P.n1005 0.000853288
R3038 P.n1004 P.n1003 0.000853288
R3039 P.n904 P.n903 0.000853288
R3040 P.n902 P.n901 0.000853288
R3041 P.n898 P.n897 0.000853288
R3042 P.n882 P.n881 0.000853288
R3043 P.n881 P.n880 0.000853288
R3044 P.n880 P.n879 0.000853288
R3045 P.n878 P.n877 0.000853288
R3046 P.n749 P.n748 0.000853288
R3047 P.n751 P.n750 0.000853288
R3048 P.n795 P.n794 0.000853288
R3049 P.n793 P.n792 0.000853288
R3050 P.n792 P.n791 0.000853288
R3051 P.n224 P.n223 0.000853288
R3052 P.n214 P.n213 0.000853288
R3053 P.n249 P.n248 0.000853288
R3054 P.n247 P.n246 0.000853288
R3055 P.n245 P.n244 0.000853288
R3056 P.n241 P.n240 0.000853288
R3057 P.n154 P.n153 0.000853288
R3058 P.n152 P.n151 0.000853288
R3059 P.n150 P.n149 0.000853288
R3060 P.n146 P.n145 0.000853288
R3061 P.n195 P.n194 0.000853288
R3062 P.n199 P.n198 0.000853288
R3063 P.n201 P.n200 0.000853288
R3064 P.n203 P.n202 0.000853288
R3065 P.n207 P.n206 0.000853288
R3066 P.n208 P.n207 0.000853288
R3067 P.n210 P.n209 0.000853288
R3068 P.n258 P.n257 0.000853288
R3069 P.n259 P.n258 0.000853288
R3070 P.n262 P.n261 0.000853288
R3071 P.n263 P.n262 0.000853288
R3072 P.n264 P.n263 0.000853288
R3073 P.n266 P.n265 0.000853288
R3074 P.n268 P.n267 0.000853288
R3075 P.n270 P.n269 0.000853288
R3076 P.n271 P.n270 0.000853288
R3077 P.n283 P.n282 0.000853288
R3078 P.n281 P.n280 0.000853288
R3079 P.n276 P.n275 0.000853288
R3080 P.n275 P.n274 0.000853288
R3081 P.n273 P.n272 0.000853288
R3082 P.n116 P.n115 0.000853288
R3083 P.n118 P.n117 0.000853288
R3084 P.n122 P.n121 0.000853288
R3085 P.n124 P.n123 0.000853288
R3086 P.n126 P.n125 0.000853288
R3087 P.n130 P.n129 0.000853288
R3088 P.n131 P.n130 0.000853288
R3089 P.n133 P.n132 0.000853288
R3090 P.n163 P.n162 0.000853288
R3091 P.n164 P.n163 0.000853288
R3092 P.n167 P.n166 0.000853288
R3093 P.n168 P.n167 0.000853288
R3094 P.n169 P.n168 0.000853288
R3095 P.n171 P.n170 0.000853288
R3096 P.n173 P.n172 0.000853288
R3097 P.n175 P.n174 0.000853288
R3098 P.n176 P.n175 0.000853288
R3099 P.n187 P.n186 0.000853288
R3100 P.n185 P.n184 0.000853288
R3101 P.n180 P.n179 0.000853288
R3102 P.n179 P.n178 0.000853288
R3103 P.n391 P.n390 0.000853288
R3104 P.n389 P.n388 0.000853288
R3105 P.n374 P.n373 0.000853288
R3106 P.n380 P.n379 0.000853288
R3107 P.n379 P.n378 0.000853288
R3108 P.n378 P.n377 0.000853288
R3109 P.n376 P.n375 0.000853288
R3110 P.n288 P.n287 0.000853288
R3111 P.n290 P.n289 0.000853288
R3112 P.n363 P.n362 0.000853288
R3113 P.n361 P.n360 0.000853288
R3114 P.n360 P.n359 0.000853288
R3115 P.n358 P.n357 0.000853288
R3116 P.n351 P.n350 0.000853288
R3117 P.n349 P.n348 0.000853288
R3118 P.n344 P.n343 0.000853288
R3119 P.n335 P.n334 0.000853288
R3120 P.n334 P.n333 0.000853288
R3121 P.n333 P.n332 0.000853288
R3122 P.n331 P.n330 0.000853288
R3123 P.n111 P.n110 0.000853288
R3124 P.n113 P.n112 0.000853288
R3125 P.n324 P.n323 0.000853288
R3126 P.n322 P.n321 0.000853288
R3127 P.n321 P.n320 0.000853288
R3128 P.n564 P.n563 0.000853288
R3129 P.n554 P.n553 0.000853288
R3130 P.n589 P.n588 0.000853288
R3131 P.n587 P.n586 0.000853288
R3132 P.n585 P.n584 0.000853288
R3133 P.n581 P.n580 0.000853288
R3134 P.n469 P.n468 0.000853288
R3135 P.n467 P.n466 0.000853288
R3136 P.n465 P.n464 0.000853288
R3137 P.n461 P.n460 0.000853288
R3138 P.n535 P.n534 0.000853288
R3139 P.n539 P.n538 0.000853288
R3140 P.n541 P.n540 0.000853288
R3141 P.n543 P.n542 0.000853288
R3142 P.n547 P.n546 0.000853288
R3143 P.n548 P.n547 0.000853288
R3144 P.n550 P.n549 0.000853288
R3145 P.n598 P.n597 0.000853288
R3146 P.n599 P.n598 0.000853288
R3147 P.n602 P.n601 0.000853288
R3148 P.n603 P.n602 0.000853288
R3149 P.n604 P.n603 0.000853288
R3150 P.n606 P.n605 0.000853288
R3151 P.n608 P.n607 0.000853288
R3152 P.n610 P.n609 0.000853288
R3153 P.n611 P.n610 0.000853288
R3154 P.n623 P.n622 0.000853288
R3155 P.n621 P.n620 0.000853288
R3156 P.n616 P.n615 0.000853288
R3157 P.n615 P.n614 0.000853288
R3158 P.n613 P.n612 0.000853288
R3159 P.n431 P.n430 0.000853288
R3160 P.n433 P.n432 0.000853288
R3161 P.n437 P.n436 0.000853288
R3162 P.n439 P.n438 0.000853288
R3163 P.n441 P.n440 0.000853288
R3164 P.n445 P.n444 0.000853288
R3165 P.n446 P.n445 0.000853288
R3166 P.n448 P.n447 0.000853288
R3167 P.n478 P.n477 0.000853288
R3168 P.n479 P.n478 0.000853288
R3169 P.n482 P.n481 0.000853288
R3170 P.n483 P.n482 0.000853288
R3171 P.n484 P.n483 0.000853288
R3172 P.n486 P.n485 0.000853288
R3173 P.n488 P.n487 0.000853288
R3174 P.n490 P.n489 0.000853288
R3175 P.n491 P.n490 0.000853288
R3176 P.n502 P.n501 0.000853288
R3177 P.n500 P.n499 0.000853288
R3178 P.n495 P.n494 0.000853288
R3179 P.n494 P.n493 0.000853288
R3180 P.n717 P.n716 0.000853288
R3181 P.n715 P.n714 0.000853288
R3182 P.n702 P.n701 0.000853288
R3183 P.n708 P.n707 0.000853288
R3184 P.n707 P.n706 0.000853288
R3185 P.n706 P.n705 0.000853288
R3186 P.n704 P.n703 0.000853288
R3187 P.n529 P.n528 0.000853288
R3188 P.n531 P.n530 0.000853288
R3189 P.n690 P.n689 0.000853288
R3190 P.n688 P.n687 0.000853288
R3191 P.n687 P.n686 0.000853288
R3192 P.n685 P.n684 0.000853288
R3193 P.n674 P.n673 0.000853288
R3194 P.n672 P.n671 0.000853288
R3195 P.n668 P.n667 0.000853288
R3196 P.n660 P.n659 0.000853288
R3197 P.n659 P.n658 0.000853288
R3198 P.n658 P.n657 0.000853288
R3199 P.n656 P.n655 0.000853288
R3200 P.n507 P.n506 0.000853288
R3201 P.n509 P.n508 0.000853288
R3202 P.n649 P.n648 0.000853288
R3203 P.n647 P.n646 0.000853288
R3204 P.n646 P.n645 0.000853288
R3205 P.n2930 P.n2929 0.000844086
R3206 P.n3282 P.n3281 0.000844086
R3207 P.n3276 P.n3275 0.000844086
R3208 P.n314 P.n313 0.000844086
R3209 P.n399 P.n398 0.000844086
R3210 P.n641 P.n640 0.000844086
R3211 P.n677 P.n670 0.000844086
R3212 P.n720 P.n713 0.000844086
R3213 P.n723 P.n722 0.000844086
R3214 P.n726 P.n725 0.000844086
R3215 P.n738 P.n737 0.000844086
R3216 P.n754 P.n745 0.000844086
R3217 P.n787 P.n786 0.000844086
R3218 P.n908 P.n900 0.000844086
R3219 P.n1049 P.n1048 0.000844086
R3220 P.n1052 P.n1051 0.000844086
R3221 P.n1094 P.n1093 0.000844086
R3222 P.n1355 P.n1340 0.000844086
R3223 P.n1358 P.n1357 0.000844086
R3224 P.n1754 P.n1753 0.000844086
R3225 P.n2010 P.n2003 0.000844086
R3226 P.n2016 P.n2015 0.000844086
R3227 P.n3497 P.n3496 0.000844086
R3228 P.n3482 P.n3481 0.000844086
R3229 P.n3477 P.n3476 0.000844086
R3230 P.n3475 P.n3474 0.000844086
R3231 P.n3431 P.n3430 0.000844086
R3232 P.n3426 P.n3425 0.000844086
R3233 P.n3424 P.n3423 0.000844086
R3234 P.n3422 P.n3421 0.000844086
R3235 P.n3420 P.n3419 0.000844086
R3236 P.n3296 P.n3295 0.000844086
R3237 P.n3293 P.n3292 0.000844086
R3238 P.n3285 P.n3284 0.000844086
R3239 P.n3429 P.n3428 0.000822581
R3240 P.n2927 P.n2926 0.000801075
R3241 P.n2936 P.n2935 0.000801075
R3242 P.n3087 P.n3086 0.000801075
R3243 P.n3279 P.n3278 0.000801075
R3244 P.n3270 P.n3269 0.000801075
R3245 P.n3136 P.n3135 0.000801075
R3246 P.n515 P.n514 0.000801075
R3247 P.n742 P.n741 0.000801075
R3248 P.n1698 P.n1697 0.000801075
R3249 P.n626 P.n525 0.00077957
R3250 P.n730 P.n729 0.00077957
R3251 P.n1039 P.n1038 0.00077957
R3252 P.n1694 P.n1693 0.00077957
R3253 P.n1751 P.n1750 0.00077957
R3254 P.n1971 P.n1865 0.00077957
R3255 P.n2013 P.n2012 0.00077957
R3256 P.n2870 P.n2869 0.000774112
R3257 P.n3354 P.n3353 0.000774112
R3258 P.n2832 P.n2831 0.000774112
R3259 P.n2906 P.n2905 0.000774112
R3260 P.n3334 P.n3333 0.000774112
R3261 P.n3389 P.n3388 0.000774112
R3262 P.n2816 P.n2815 0.000774112
R3263 P.n3317 P.n3316 0.000774112
R3264 P.n2304 P.n2303 0.000774112
R3265 P.n2394 P.n2393 0.000774112
R3266 P.n2266 P.n2265 0.000774112
R3267 P.n2340 P.n2339 0.000774112
R3268 P.n2374 P.n2373 0.000774112
R3269 P.n2429 P.n2428 0.000774112
R3270 P.n2250 P.n2249 0.000774112
R3271 P.n2357 P.n2356 0.000774112
R3272 P.n3641 P.n3640 0.000774112
R3273 P.n2069 P.n2068 0.000774112
R3274 P.n3603 P.n3602 0.000774112
R3275 P.n3677 P.n3676 0.000774112
R3276 P.n2049 P.n2048 0.000774112
R3277 P.n2104 P.n2103 0.000774112
R3278 P.n3686 P.n3685 0.000774112
R3279 P.n2032 P.n2031 0.000774112
R3280 P.n2583 P.n2582 0.000774112
R3281 P.n2667 P.n2666 0.000774112
R3282 P.n2545 P.n2544 0.000774112
R3283 P.n2619 P.n2618 0.000774112
R3284 P.n2647 P.n2646 0.000774112
R3285 P.n2702 P.n2701 0.000774112
R3286 P.n2529 P.n2528 0.000774112
R3287 P.n2630 P.n2629 0.000774112
R3288 P.n3012 P.n3011 0.000774112
R3289 P.n3196 P.n3195 0.000774112
R3290 P.n2974 P.n2973 0.000774112
R3291 P.n3048 P.n3047 0.000774112
R3292 P.n3176 P.n3175 0.000774112
R3293 P.n3231 P.n3230 0.000774112
R3294 P.n3071 P.n3070 0.000774112
R3295 P.n3253 P.n3252 0.000774112
R3296 P.n1916 P.n1915 0.000764966
R3297 P.n1788 P.n1787 0.000764966
R3298 P.n1878 P.n1877 0.000764966
R3299 P.n1952 P.n1951 0.000764966
R3300 P.n1768 P.n1767 0.000764966
R3301 P.n1823 P.n1822 0.000764966
R3302 P.n1725 P.n1724 0.000764966
R3303 P.n1715 P.n1714 0.000764966
R3304 P.n1478 P.n1477 0.000764966
R3305 P.n1589 P.n1588 0.000764966
R3306 P.n1440 P.n1439 0.000764966
R3307 P.n1514 P.n1513 0.000764966
R3308 P.n1569 P.n1568 0.000764966
R3309 P.n1624 P.n1623 0.000764966
R3310 P.n1424 P.n1423 0.000764966
R3311 P.n1552 P.n1551 0.000764966
R3312 P.n1163 P.n1162 0.000764966
R3313 P.n1241 P.n1240 0.000764966
R3314 P.n1125 P.n1124 0.000764966
R3315 P.n1199 P.n1198 0.000764966
R3316 P.n1221 P.n1220 0.000764966
R3317 P.n1276 P.n1275 0.000764966
R3318 P.n1109 P.n1108 0.000764966
R3319 P.n1072 P.n1071 0.000764966
R3320 P.n959 P.n958 0.000764966
R3321 P.n832 P.n831 0.000764966
R3322 P.n921 P.n920 0.000764966
R3323 P.n995 P.n994 0.000764966
R3324 P.n812 P.n811 0.000764966
R3325 P.n867 P.n866 0.000764966
R3326 P.n762 P.n761 0.000764966
R3327 P.n750 P.n749 0.000764966
R3328 P.n243 P.n242 0.000764966
R3329 P.n148 P.n147 0.000764966
R3330 P.n205 P.n204 0.000764966
R3331 P.n279 P.n278 0.000764966
R3332 P.n128 P.n127 0.000764966
R3333 P.n183 P.n182 0.000764966
R3334 P.n289 P.n288 0.000764966
R3335 P.n112 P.n111 0.000764966
R3336 P.n583 P.n582 0.000764966
R3337 P.n463 P.n462 0.000764966
R3338 P.n545 P.n544 0.000764966
R3339 P.n619 P.n618 0.000764966
R3340 P.n443 P.n442 0.000764966
R3341 P.n498 P.n497 0.000764966
R3342 P.n530 P.n529 0.000764966
R3343 P.n508 P.n507 0.000764966
R3344 P.n107 P.n106 0.000758065
R3345 P.n293 P.n192 0.000758065
R3346 P.n304 P.n303 0.000758065
R3347 P.n876 P.n789 0.000758065
R3348 P.n1388 P.n1387 0.000758065
R3349 P.n1747 P.n1746 0.000758065
R3350 P.n3579 P.n3578 0.000758065
R3351 P.n3512 P.n3511 0.000758065
R3352 P.n3508 P.n3507 0.000758065
R3353 P.n3503 P.n3502 0.000758065
R3354 P.n82 P.n81 0.000736559
R3355 P.n102 P.n101 0.000736559
R3356 P.n303 P.n302 0.000736559
R3357 P.n310 P.n309 0.000736559
R3358 P.n396 P.n395 0.000736559
R3359 P.n637 P.n636 0.000736559
R3360 P.n678 P.n677 0.000736559
R3361 P.n775 P.n774 0.000736559
R3362 P.n782 P.n781 0.000736559
R3363 P.n1090 P.n1089 0.000736559
R3364 P.n1360 P.n1359 0.000736559
R3365 P.n1371 P.n1370 0.000736559
R3366 P.n1373 P.n1372 0.000736559
R3367 P.n1375 P.n1374 0.000736559
R3368 P.n1377 P.n1376 0.000736559
R3369 P.n1379 P.n1378 0.000736559
R3370 P.n1381 P.n1380 0.000736559
R3371 P.n1382 P.n1381 0.000736559
R3372 P.n1401 P.n1400 0.000736559
R3373 P.n1403 P.n1402 0.000736559
R3374 P.n1409 P.n1408 0.000736559
R3375 P.n1682 P.n1674 0.000736559
R3376 P.n1688 P.n1687 0.000736559
R3377 P.n1739 P.n1738 0.000736559
R3378 P.n1746 P.n1745 0.000736559
R3379 P.n3708 P.n3707 0.000736559
R3380 P.n3698 P.n3697 0.000736559
R3381 P.n3696 P.n3695 0.000736559
R3382 P.n3694 P.n3693 0.000736559
R3383 P.n3590 P.n3589 0.000736559
R3384 P.n3588 P.n3587 0.000736559
R3385 P.n3586 P.n3585 0.000736559
R3386 P.n3585 P.n3584 0.000736559
R3387 P.n3575 P.n3564 0.000736559
R3388 P.n3563 P.n3562 0.000736559
R3389 P.n3557 P.n3556 0.000736559
R3390 P.n3551 P.n3550 0.000736559
R3391 P.n3545 P.n3544 0.000736559
R3392 P.n3533 P.n3532 0.000736559
R3393 P.n3516 P.n3515 0.000736559
R3394 P.n3504 P.n3503 0.000736559
R3395 P.n3501 P.n3500 0.000736559
R3396 P.n3485 P.n3484 0.000736559
R3397 P.n3439 P.n3438 0.000736559
R3398 P.n3436 P.n3435 0.000736559
R3399 P.n3305 P.n3299 0.000736559
R3400 P.n93 P.n85 0.000715054
R3401 P.n190 P.n107 0.000715054
R3402 P.n192 P.n191 0.000715054
R3403 P.n354 P.n347 0.000715054
R3404 P.n514 P.n513 0.000715054
R3405 P.n697 P.n683 0.000715054
R3406 P.n757 P.n756 0.000715054
R3407 P.n768 P.n767 0.000715054
R3408 P.n1078 P.n1077 0.000715054
R3409 P.n1387 P.n1386 0.000715054
R3410 P.n1729 P.n1720 0.000715054
R3411 P.n1731 P.n1730 0.000715054
R3412 P.n3580 P.n3579 0.000715054
R3413 P.n3541 P.n3540 0.000715054
R3414 P.n3529 P.n3528 0.000715054
R3415 P.n3511 P.n3510 0.000715054
R3416 P.n3509 P.n3508 0.000715054
R3417 P.n3491 P.n3490 0.000715054
R3418 P.n3445 P.n3444 0.000715054
R3419 P.n3442 P.n3441 0.000715054
R3420 P.n3308 P.n3307 0.000715054
R3421 P.n3091 P.n3090 0.000693548
R3422 P.n3103 P.n3102 0.000693548
R3423 P.n3132 P.n3131 0.000693548
R3424 P.n3120 P.n3119 0.000693548
R3425 P.n315 P.n314 0.000693548
R3426 P.n368 P.n354 0.000693548
R3427 P.n397 P.n396 0.000693548
R3428 P.n404 P.n403 0.000693548
R3429 P.n408 P.n407 0.000693548
R3430 P.n416 P.n415 0.000693548
R3431 P.n516 P.n515 0.000693548
R3432 P.n525 P.n524 0.000693548
R3433 P.n628 P.n627 0.000693548
R3434 P.n683 P.n682 0.000693548
R3435 P.n741 P.n740 0.000693548
R3436 P.n1683 P.n1682 0.000693548
R3437 P.n3550 P.n3549 0.000693548
R3438 P.n3496 P.n3495 0.000693548
R3439 P.n3490 P.n3489 0.000693548
R3440 P.n3484 P.n3483 0.000693548
R3441 P.n3435 P.n3434 0.000693548
R3442 P.n2814 P.n2813 0.000682741
R3443 P.n2801 P.n2798 0.000682741
R3444 P.n3315 P.n3314 0.000682741
R3445 P.n2753 P.n2746 0.000682741
R3446 P.n2248 P.n2247 0.000682741
R3447 P.n2355 P.n2354 0.000682741
R3448 P.n3684 P.n3683 0.000682741
R3449 P.n2030 P.n2029 0.000682741
R3450 P.n2527 P.n2526 0.000682741
R3451 P.n2628 P.n2627 0.000682741
R3452 P.n2942 P.n2941 0.000682741
R3453 P.n2944 P.n2943 0.000682741
R3454 P.n2954 P.n2953 0.000682741
R3455 P.n2959 P.n2958 0.000682741
R3456 P.n2961 P.n2960 0.000682741
R3457 P.n3083 P.n2961 0.000682741
R3458 P.n3082 P.n3081 0.000682741
R3459 P.n3073 P.n3072 0.000682741
R3460 P.n3067 P.n3066 0.000682741
R3461 P.n3065 P.n3064 0.000682741
R3462 P.n3064 P.n3063 0.000682741
R3463 P.n3063 P.n3062 0.000682741
R3464 P.n3061 P.n3060 0.000682741
R3465 P.n3143 P.n3142 0.000682741
R3466 P.n3145 P.n3144 0.000682741
R3467 P.n3155 P.n3154 0.000682741
R3468 P.n3160 P.n3159 0.000682741
R3469 P.n3162 P.n3161 0.000682741
R3470 P.n3265 P.n3162 0.000682741
R3471 P.n3264 P.n3263 0.000682741
R3472 P.n3255 P.n3254 0.000682741
R3473 P.n3249 P.n3248 0.000682741
R3474 P.n3247 P.n3246 0.000682741
R3475 P.n3246 P.n3245 0.000682741
R3476 P.n3245 P.n3244 0.000682741
R3477 P.n3243 P.n3242 0.000682741
R3478 P.n1723 P.n1722 0.000676644
R3479 P.n1713 P.n1712 0.000676644
R3480 P.n1422 P.n1421 0.000676644
R3481 P.n1550 P.n1549 0.000676644
R3482 P.n1107 P.n1106 0.000676644
R3483 P.n1206 P.n1205 0.000676644
R3484 P.n1103 P.n1102 0.000676644
R3485 P.n1309 P.n1308 0.000676644
R3486 P.n1070 P.n1069 0.000676644
R3487 P.n760 P.n759 0.000676644
R3488 P.n748 P.n747 0.000676644
R3489 P.n287 P.n286 0.000676644
R3490 P.n110 P.n109 0.000676644
R3491 P.n326 P.n325 0.000676644
R3492 P.n425 P.n423 0.000676644
R3493 P.n710 P.n709 0.000676644
R3494 P.n528 P.n527 0.000676644
R3495 P.n61 P.n59 0.000676644
R3496 P.n506 P.n505 0.000676644
R3497 P.n651 P.n650 0.000676644
R3498 P.n2933 P.n2932 0.000672043
R3499 P.n3088 P.n3087 0.000672043
R3500 P.n3273 P.n3272 0.000672043
R3501 P.n3135 P.n3134 0.000672043
R3502 P.n1368 P.n1367 0.000672043
R3503 P.n1523 P.n1409 0.000672043
R3504 P.n3701 P.n3700 0.000672043
R3505 P.n3556 P.n3555 0.000672043
R3506 P.n3402 P.n3401 0.000672043
R3507 P.n3096 P.n3095 0.000650538
R3508 P.n3127 P.n3126 0.000650538
R3509 P.n78 P.n77 0.000650538
R3510 P.n191 P.n190 0.000650538
R3511 P.n294 P.n293 0.000650538
R3512 P.n386 P.n385 0.000650538
R3513 P.n513 P.n512 0.000650538
R3514 P.n627 P.n626 0.000650538
R3515 P.n682 P.n681 0.000650538
R3516 P.n767 P.n766 0.000650538
R3517 P.n1077 P.n1076 0.000650538
R3518 P.n1363 P.n1362 0.000650538
R3519 P.n1383 P.n1382 0.000650538
R3520 P.n1406 P.n1405 0.000650538
R3521 P.n1642 P.n1547 0.000650538
R3522 P.n1685 P.n1684 0.000650538
R3523 P.n1720 P.n1719 0.000650538
R3524 P.n1730 P.n1729 0.000650538
R3525 P.n3705 P.n3704 0.000650538
R3526 P.n3584 P.n3583 0.000650538
R3527 P.n3560 P.n3559 0.000650538
R3528 P.n3554 P.n3553 0.000650538
R3529 P.n3548 P.n3547 0.000650538
R3530 P.n3537 P.n3536 0.000650538
R3531 P.n3510 P.n3509 0.000650538
R3532 P.n3507 P.n3506 0.000650538
R3533 P.n3488 P.n3487 0.000650538
R3534 P.n3446 P.n3445 0.000650538
R3535 P.n3443 P.n3442 0.000650538
R3536 P.n3309 P.n3308 0.000650538
R3537 P.n2938 P.n2937 0.000629032
R3538 P.n3268 P.n3267 0.000629032
R3539 P.n302 P.n295 0.000629032
R3540 P.n309 P.n304 0.000629032
R3541 P.n329 P.n316 0.000629032
R3542 P.n347 P.n346 0.000629032
R3543 P.n523 P.n516 0.000629032
R3544 P.n636 P.n630 0.000629032
R3545 P.n745 P.n744 0.000629032
R3546 P.n756 P.n755 0.000629032
R3547 P.n766 P.n757 0.000629032
R3548 P.n774 P.n768 0.000629032
R3549 P.n776 P.n775 0.000629032
R3550 P.n781 P.n776 0.000629032
R3551 P.n783 P.n782 0.000629032
R3552 P.n1089 P.n1079 0.000629032
R3553 P.n1380 P.n1379 0.000629032
R3554 P.n1385 P.n1384 0.000629032
R3555 P.n1393 P.n1388 0.000629032
R3556 P.n1400 P.n1394 0.000629032
R3557 P.n1690 P.n1689 0.000629032
R3558 P.n1732 P.n1731 0.000629032
R3559 P.n1738 P.n1732 0.000629032
R3560 P.n1745 P.n1739 0.000629032
R3561 P.n3587 P.n3586 0.000629032
R3562 P.n3582 P.n3581 0.000629032
R3563 P.n3578 P.n3577 0.000629032
R3564 P.n3576 P.n3575 0.000629032
R3565 P.n3505 P.n3504 0.000629032
R3566 P.n3502 P.n3501 0.000629032
R3567 P.n3494 P.n3493 0.000629032
R3568 P.n3492 P.n3491 0.000629032
R3569 P.n3440 P.n3439 0.000629032
R3570 P.n3437 P.n3436 0.000629032
R3571 P.n3306 P.n3305 0.000629032
R3572 P.n3094 P.n3093 0.000607527
R3573 P.n3102 P.n3101 0.000607527
R3574 P.n3129 P.n3128 0.000607527
R3575 P.n3121 P.n3120 0.000607527
R3576 P.n395 P.n387 0.000607527
R3577 P.n680 P.n679 0.000607527
R3578 P.n1394 P.n1393 0.000607527
R3579 P.n1408 P.n1407 0.000607527
R3580 P.n1674 P.n1666 0.000607527
R3581 P.n1687 P.n1686 0.000607527
R3582 P.n1719 P.n1710 0.000607527
R3583 P.n3577 P.n3576 0.000607527
R3584 P.n3558 P.n3557 0.000607527
R3585 P.n3552 P.n3551 0.000607527
R3586 P.n3546 P.n3545 0.000607527
R3587 P.n3486 P.n3485 0.000607527
R3588 P.n2863 P.n2862 0.000591371
R3589 P.n3348 P.n3347 0.000591371
R3590 P.n2833 P.n2832 0.000591371
R3591 P.n2905 P.n2904 0.000591371
R3592 P.n3335 P.n3334 0.000591371
R3593 P.n3388 P.n3387 0.000591371
R3594 P.n2810 P.n2809 0.000591371
R3595 P.n3412 P.n3411 0.000591371
R3596 P.n2798 P.n2797 0.000591371
R3597 P.n2753 P.n2752 0.000591371
R3598 P.n2297 P.n2296 0.000591371
R3599 P.n2388 P.n2387 0.000591371
R3600 P.n2267 P.n2266 0.000591371
R3601 P.n2339 P.n2338 0.000591371
R3602 P.n2375 P.n2374 0.000591371
R3603 P.n2428 P.n2427 0.000591371
R3604 P.n3526 P.n3525 0.000591371
R3605 P.n2210 P.n2209 0.000591371
R3606 P.n2441 P.n2440 0.000591371
R3607 P.n2218 P.n2217 0.000591371
R3608 P.n3634 P.n3633 0.000591371
R3609 P.n2063 P.n2062 0.000591371
R3610 P.n3604 P.n3603 0.000591371
R3611 P.n3676 P.n3675 0.000591371
R3612 P.n2050 P.n2049 0.000591371
R3613 P.n2103 P.n2102 0.000591371
R3614 P.n2176 P.n2175 0.000591371
R3615 P.n2131 P.n2130 0.000591371
R3616 P.n2169 P.n2168 0.000591371
R3617 P.n2120 P.n2119 0.000591371
R3618 P.n2576 P.n2575 0.000591371
R3619 P.n2661 P.n2660 0.000591371
R3620 P.n2546 P.n2545 0.000591371
R3621 P.n2618 P.n2617 0.000591371
R3622 P.n2648 P.n2647 0.000591371
R3623 P.n2701 P.n2700 0.000591371
R3624 P.n3459 P.n3458 0.000591371
R3625 P.n2475 P.n2474 0.000591371
R3626 P.n2721 P.n2720 0.000591371
R3627 P.n2483 P.n2482 0.000591371
R3628 P.n3005 P.n3004 0.000591371
R3629 P.n3190 P.n3189 0.000591371
R3630 P.n2975 P.n2974 0.000591371
R3631 P.n3047 P.n3046 0.000591371
R3632 P.n3177 P.n3176 0.000591371
R3633 P.n3230 P.n3229 0.000591371
R3634 P.n2953 P.n2952 0.000591371
R3635 P.n3060 P.n3059 0.000591371
R3636 P.n3154 P.n3153 0.000591371
R3637 P.n3242 P.n3241 0.000591371
R3638 P.n1909 P.n1908 0.000588322
R3639 P.n1782 P.n1781 0.000588322
R3640 P.n1879 P.n1878 0.000588322
R3641 P.n1951 P.n1950 0.000588322
R3642 P.n1769 P.n1768 0.000588322
R3643 P.n1822 P.n1821 0.000588322
R3644 P.n1984 P.n1983 0.000588322
R3645 P.n1967 P.n1966 0.000588322
R3646 P.n1855 P.n1854 0.000588322
R3647 P.n1837 P.n1836 0.000588322
R3648 P.n1471 P.n1470 0.000588322
R3649 P.n1583 P.n1582 0.000588322
R3650 P.n1441 P.n1440 0.000588322
R3651 P.n1513 P.n1512 0.000588322
R3652 P.n1570 P.n1569 0.000588322
R3653 P.n1623 P.n1622 0.000588322
R3654 P.n1537 P.n1536 0.000588322
R3655 P.n1417 P.n1416 0.000588322
R3656 P.n1656 P.n1655 0.000588322
R3657 P.n1638 P.n1637 0.000588322
R3658 P.n1156 P.n1155 0.000588322
R3659 P.n1235 P.n1234 0.000588322
R3660 P.n1126 P.n1125 0.000588322
R3661 P.n1198 P.n1197 0.000588322
R3662 P.n1222 P.n1221 0.000588322
R3663 P.n1275 P.n1274 0.000588322
R3664 P.n1321 P.n1320 0.000588322
R3665 P.n1102 P.n1101 0.000588322
R3666 P.n1308 P.n1307 0.000588322
R3667 P.n1290 P.n1289 0.000588322
R3668 P.n952 P.n951 0.000588322
R3669 P.n826 P.n825 0.000588322
R3670 P.n922 P.n921 0.000588322
R3671 P.n994 P.n993 0.000588322
R3672 P.n813 P.n812 0.000588322
R3673 P.n866 P.n865 0.000588322
R3674 P.n1028 P.n1027 0.000588322
R3675 P.n1010 P.n1009 0.000588322
R3676 P.n890 P.n889 0.000588322
R3677 P.n796 P.n795 0.000588322
R3678 P.n236 P.n235 0.000588322
R3679 P.n142 P.n141 0.000588322
R3680 P.n206 P.n205 0.000588322
R3681 P.n278 P.n277 0.000588322
R3682 P.n129 P.n128 0.000588322
R3683 P.n182 P.n181 0.000588322
R3684 P.n98 P.n97 0.000588322
R3685 P.n364 P.n363 0.000588322
R3686 P.n90 P.n89 0.000588322
R3687 P.n325 P.n324 0.000588322
R3688 P.n576 P.n575 0.000588322
R3689 P.n457 P.n456 0.000588322
R3690 P.n546 P.n545 0.000588322
R3691 P.n618 P.n617 0.000588322
R3692 P.n444 P.n443 0.000588322
R3693 P.n497 P.n496 0.000588322
R3694 P.n423 P.n422 0.000588322
R3695 P.n691 P.n690 0.000588322
R3696 P.n59 P.n58 0.000588322
R3697 P.n650 P.n649 0.000588322
R3698 P.n3092 P.n3091 0.000586021
R3699 P.n3104 P.n3103 0.000586021
R3700 P.n3131 P.n3130 0.000586021
R3701 P.n3119 P.n3118 0.000586021
R3702 P.n75 P.n74 0.000586021
R3703 P.n77 P.n76 0.000586021
R3704 P.n295 P.n294 0.000586021
R3705 P.n313 P.n312 0.000586021
R3706 P.n316 P.n315 0.000586021
R3707 P.n346 P.n329 0.000586021
R3708 P.n385 P.n368 0.000586021
R3709 P.n387 P.n386 0.000586021
R3710 P.n398 P.n397 0.000586021
R3711 P.n402 P.n401 0.000586021
R3712 P.n407 P.n406 0.000586021
R3713 P.n418 P.n417 0.000586021
R3714 P.n640 P.n639 0.000586021
R3715 P.n670 P.n654 0.000586021
R3716 P.n679 P.n678 0.000586021
R3717 P.n681 P.n680 0.000586021
R3718 P.n713 P.n697 0.000586021
R3719 P.n722 P.n721 0.000586021
R3720 P.n727 P.n726 0.000586021
R3721 P.n729 P.n728 0.000586021
R3722 P.n786 P.n785 0.000586021
R3723 P.n789 P.n788 0.000586021
R3724 P.n900 P.n876 0.000586021
R3725 P.n1038 P.n1014 0.000586021
R3726 P.n1051 P.n1050 0.000586021
R3727 P.n1056 P.n1055 0.000586021
R3728 P.n1093 P.n1092 0.000586021
R3729 P.n1340 P.n1294 0.000586021
R3730 P.n1357 P.n1356 0.000586021
R3731 P.n1362 P.n1361 0.000586021
R3732 P.n1364 P.n1363 0.000586021
R3733 P.n1365 P.n1364 0.000586021
R3734 P.n1384 P.n1383 0.000586021
R3735 P.n1405 P.n1404 0.000586021
R3736 P.n1407 P.n1406 0.000586021
R3737 P.n1547 P.n1523 0.000586021
R3738 P.n1666 P.n1642 0.000586021
R3739 P.n1684 P.n1683 0.000586021
R3740 P.n1686 P.n1685 0.000586021
R3741 P.n1693 P.n1692 0.000586021
R3742 P.n1695 P.n1694 0.000586021
R3743 P.n1750 P.n1749 0.000586021
R3744 P.n1865 P.n1841 0.000586021
R3745 P.n2012 P.n2011 0.000586021
R3746 P.n3706 P.n3705 0.000586021
R3747 P.n3704 P.n3703 0.000586021
R3748 P.n3583 P.n3582 0.000586021
R3749 P.n3561 P.n3560 0.000586021
R3750 P.n3559 P.n3558 0.000586021
R3751 P.n3555 P.n3554 0.000586021
R3752 P.n3553 P.n3552 0.000586021
R3753 P.n3549 P.n3548 0.000586021
R3754 P.n3547 P.n3546 0.000586021
R3755 P.n3540 P.n3539 0.000586021
R3756 P.n3538 P.n3537 0.000586021
R3757 P.n3506 P.n3505 0.000586021
R3758 P.n3498 P.n3497 0.000586021
R3759 P.n3495 P.n3494 0.000586021
R3760 P.n3493 P.n3492 0.000586021
R3761 P.n3489 P.n3488 0.000586021
R3762 P.n3487 P.n3486 0.000586021
R3763 P.n3483 P.n3482 0.000586021
R3764 P.n3478 P.n3477 0.000586021
R3765 P.n3476 P.n3475 0.000586021
R3766 P.n3432 P.n3431 0.000586021
R3767 P.n3430 P.n3429 0.000586021
R3768 P.n3425 P.n3424 0.000586021
R3769 P.n3423 P.n3422 0.000586021
R3770 P.n3421 P.n3420 0.000586021
R3771 P.n3416 P.n3404 0.000586021
R3772 P.n3297 P.n3296 0.000586021
R3773 P.n3294 P.n3293 0.000586021
R3774 P.n3286 P.n3285 0.000586021
R3775 P.n79 P.n78 0.000564516
R3776 P.n81 P.n80 0.000564516
R3777 P.n405 P.n404 0.000564516
R3778 P.n410 P.n409 0.000564516
R3779 P.n731 P.n730 0.000564516
R3780 P.n733 P.n732 0.000564516
R3781 P.n788 P.n787 0.000564516
R3782 P.n1014 P.n908 0.000564516
R3783 P.n1047 P.n1039 0.000564516
R3784 P.n1050 P.n1049 0.000564516
R3785 P.n1058 P.n1057 0.000564516
R3786 P.n1367 P.n1366 0.000564516
R3787 P.n1369 P.n1368 0.000564516
R3788 P.n1697 P.n1696 0.000564516
R3789 P.n1699 P.n1698 0.000564516
R3790 P.n1752 P.n1751 0.000564516
R3791 P.n1979 P.n1971 0.000564516
R3792 P.n2011 P.n2010 0.000564516
R3793 P.n2014 P.n2013 0.000564516
R3794 P.n3702 P.n3701 0.000564516
R3795 P.n3700 P.n3699 0.000564516
R3796 P.n3536 P.n3535 0.000564516
R3797 P.n3534 P.n3533 0.000564516
R3798 P.n3474 P.n3473 0.000564516
R3799 P.n3472 P.n3471 0.000564516
R3800 P.n3449 P.n3448 0.000564516
R3801 P.n3444 P.n3443 0.000564516
R3802 P.n3441 P.n3440 0.000564516
R3803 P.n3438 P.n3437 0.000564516
R3804 P.n3427 P.n3426 0.000564516
R3805 P.n3403 P.n3402 0.000564516
R3806 P.n2926 P.n2925 0.000543011
R3807 P.n2928 P.n2927 0.000543011
R3808 P.n2934 P.n2933 0.000543011
R3809 P.n2937 P.n2936 0.000543011
R3810 P.n3084 P.n2938 0.000543011
R3811 P.n3086 P.n3085 0.000543011
R3812 P.n3095 P.n3094 0.000543011
R3813 P.n3097 P.n3096 0.000543011
R3814 P.n3098 P.n3097 0.000543011
R3815 P.n3099 P.n3098 0.000543011
R3816 P.n3101 P.n3100 0.000543011
R3817 P.n3280 P.n3279 0.000543011
R3818 P.n3278 P.n3277 0.000543011
R3819 P.n3272 P.n3271 0.000543011
R3820 P.n3269 P.n3268 0.000543011
R3821 P.n3267 P.n3266 0.000543011
R3822 P.n3137 P.n3136 0.000543011
R3823 P.n3128 P.n3127 0.000543011
R3824 P.n3126 P.n3125 0.000543011
R3825 P.n3125 P.n3124 0.000543011
R3826 P.n3124 P.n3123 0.000543011
R3827 P.n3122 P.n3121 0.000543011
R3828 P.n524 P.n523 0.000543011
R3829 P.n1841 P.n1754 0.000543011
R3830 P.n3447 P.n3446 0.000543011
R3831 P.n629 P.n628 0.000521505
R3832 P.n755 P.n754 0.000521505
R3833 P.n1048 P.n1047 0.000521505
R3834 P.n1386 P.n1385 0.000521505
R3835 P.n1753 P.n1752 0.000521505
R3836 P.n2003 P.n1979 0.000521505
R3837 P.n2015 P.n2014 0.000521505
R3838 P.n3581 P.n3580 0.000521505
R3839 P.n3543 P.n3542 0.000521505
R3840 P.n3428 P.n3427 0.000521505
R3841 M.n1173 M.t80 3.41655
R3842 M.n1162 M.t122 3.41655
R3843 M.n1151 M.t116 3.41655
R3844 M.n1126 M.t71 3.41655
R3845 M.n1115 M.t118 3.41655
R3846 M.n44 M.t20 3.41655
R3847 M.n55 M.t23 3.41655
R3848 M.n33 M.t65 3.41655
R3849 M.n22 M.t108 3.41655
R3850 M.n11 M.t61 3.41655
R3851 M.n0 M.t74 3.41655
R3852 M.n1495 M.n1470 2.26934
R3853 M.n1173 M.t101 2.25428
R3854 M.n1174 M.t58 2.25428
R3855 M.n1175 M.t9 2.25428
R3856 M.n1176 M.t17 2.25428
R3857 M.n1177 M.t128 2.25428
R3858 M.n1178 M.t81 2.25428
R3859 M.n1179 M.t47 2.25428
R3860 M.n1180 M.t127 2.25428
R3861 M.n1181 M.t5 2.25428
R3862 M.n1182 M.t111 2.25428
R3863 M.n1183 M.t57 2.25428
R3864 M.n1162 M.t44 2.25428
R3865 M.n1163 M.t115 2.25428
R3866 M.n1164 M.t59 2.25428
R3867 M.n1165 M.t75 2.25428
R3868 M.n1166 M.t41 2.25428
R3869 M.n1167 M.t130 2.25428
R3870 M.n1168 M.t102 2.25428
R3871 M.n1169 M.t39 2.25428
R3872 M.n1170 M.t51 2.25428
R3873 M.n1171 M.t28 2.25428
R3874 M.n1172 M.t113 2.25428
R3875 M.n1151 M.t94 2.25428
R3876 M.n1152 M.t97 2.25428
R3877 M.n1153 M.t40 2.25428
R3878 M.n1154 M.t53 2.25428
R3879 M.n1155 M.t29 2.25428
R3880 M.n1156 M.t114 2.25428
R3881 M.n1157 M.t91 2.25428
R3882 M.n1158 M.t27 2.25428
R3883 M.n1159 M.t34 2.25428
R3884 M.n1160 M.t18 2.25428
R3885 M.n1161 M.t95 2.25428
R3886 M.n1126 M.t64 2.25428
R3887 M.n1127 M.t14 2.25428
R3888 M.n1128 M.t92 2.25428
R3889 M.n1129 M.t99 2.25428
R3890 M.n1130 M.t83 2.25428
R3891 M.n1131 M.t24 2.25428
R3892 M.n1132 M.t7 2.25428
R3893 M.n1133 M.t82 2.25428
R3894 M.n1134 M.t88 2.25428
R3895 M.n1135 M.t60 2.25428
R3896 M.n1136 M.t12 2.25428
R3897 M.n1115 M.t10 2.25428
R3898 M.n1116 M.t69 2.25428
R3899 M.n1117 M.t15 2.25428
R3900 M.n1118 M.t22 2.25428
R3901 M.n1119 M.t3 2.25428
R3902 M.n1120 M.t85 2.25428
R3903 M.n1121 M.t54 2.25428
R3904 M.n1122 M.t1 2.25428
R3905 M.n1123 M.t8 2.25428
R3906 M.n1124 M.t119 2.25428
R3907 M.n1125 M.t67 2.25428
R3908 M.n44 M.t86 2.25428
R3909 M.n45 M.t4 2.25428
R3910 M.n46 M.t84 2.25428
R3911 M.n47 M.t90 2.25428
R3912 M.n48 M.t68 2.25428
R3913 M.n49 M.t16 2.25428
R3914 M.n50 M.t125 2.25428
R3915 M.n51 M.t63 2.25428
R3916 M.n52 M.t79 2.25428
R3917 M.n53 M.t46 2.25428
R3918 M.n54 M.t2 2.25428
R3919 M.n55 M.t73 2.25428
R3920 M.n56 M.t120 2.25428
R3921 M.n57 M.t62 2.25428
R3922 M.n58 M.t78 2.25428
R3923 M.n59 M.t45 2.25428
R3924 M.n60 M.t0 2.25428
R3925 M.n61 M.t105 2.25428
R3926 M.n62 M.t42 2.25428
R3927 M.n63 M.t55 2.25428
R3928 M.n64 M.t31 2.25428
R3929 M.n65 M.t117 2.25428
R3930 M.n33 M.t32 2.25428
R3931 M.n34 M.t21 2.25428
R3932 M.n35 M.t98 2.25428
R3933 M.n36 M.t109 2.25428
R3934 M.n37 M.t89 2.25428
R3935 M.n38 M.t30 2.25428
R3936 M.n39 M.t13 2.25428
R3937 M.n40 M.t87 2.25428
R3938 M.n41 M.t93 2.25428
R3939 M.n42 M.t76 2.25428
R3940 M.n43 M.t19 2.25428
R3941 M.n22 M.t77 2.25428
R3942 M.n23 M.t106 2.25428
R3943 M.n24 M.t52 2.25428
R3944 M.n25 M.t66 2.25428
R3945 M.n26 M.t35 2.25428
R3946 M.n27 M.t124 2.25428
R3947 M.n28 M.t96 2.25428
R3948 M.n29 M.t33 2.25428
R3949 M.n30 M.t43 2.25428
R3950 M.n31 M.t25 2.25428
R3951 M.n32 M.t104 2.25428
R3952 M.n11 M.t129 2.25428
R3953 M.n12 M.t50 2.25428
R3954 M.n13 M.t6 2.25428
R3955 M.n14 M.t11 2.25428
R3956 M.n15 M.t123 2.25428
R3957 M.n16 M.t72 2.25428
R3958 M.n17 M.t38 2.25428
R3959 M.n18 M.t121 2.25428
R3960 M.n19 M.t131 2.25428
R3961 M.n20 M.t103 2.25428
R3962 M.n21 M.t49 2.25428
R3963 M.n0 M.t110 2.25428
R3964 M.n1 M.t112 2.25428
R3965 M.n2 M.t56 2.25428
R3966 M.n3 M.t70 2.25428
R3967 M.n4 M.t37 2.25428
R3968 M.n5 M.t126 2.25428
R3969 M.n6 M.t100 2.25428
R3970 M.n7 M.t36 2.25428
R3971 M.n8 M.t48 2.25428
R3972 M.n9 M.t26 2.25428
R3973 M.n10 M.t107 2.25428
R3974 M.n1841 M.n1840 2.2505
R3975 M.n1980 M.n1979 2.2505
R3976 M.n1990 M.n1973 2.2505
R3977 M.n1982 M.n1981 2.2505
R3978 M.n1987 M.n1986 2.2505
R3979 M.n1976 M.n1974 2.2505
R3980 M.n1839 M.n1838 2.2505
R3981 M.n1993 M.n1972 2.2505
R3982 M.n1726 M.n1712 2.2505
R3983 M.n1809 M.n1808 2.2505
R3984 M.n1815 M.n1806 2.2505
R3985 M.n1759 M.n1758 2.2505
R3986 M.n1812 M.n1807 2.2505
R3987 M.n1720 M.n1715 2.2505
R3988 M.n1721 M.n1713 2.2505
R3989 M.n1519 M.n1518 2.2505
R3990 M.n1650 M.n1641 2.2505
R3991 M.n1655 M.n1639 2.2505
R3992 M.n1646 M.n1642 2.2505
R3993 M.n1517 M.n1516 2.2505
R3994 M.n1509 M.n1508 2.2505
R3995 M.n1651 M.n1640 2.2505
R3996 M.n1511 M.n1510 2.2505
R3997 M.n1481 M.n1480 2.2505
R3998 M.n1489 M.n1471 2.2505
R3999 M.n1486 M.n1472 2.2505
R4000 M.n1476 M.n1474 2.2505
R4001 M.n1340 M.n1339 2.2505
R4002 M.n1482 M.n1473 2.2505
R4003 M.n968 M.n939 2.2505
R4004 M.n971 M.n938 2.2505
R4005 M.n965 M.n940 2.2505
R4006 M.n957 M.n943 2.2505
R4007 M.n961 M.n941 2.2505
R4008 M.n952 M.n945 2.2505
R4009 M.n960 M.n942 2.2505
R4010 M.n950 M.n949 2.2505
R4011 M.n901 M.n900 2.2505
R4012 M.n926 M.n925 2.2505
R4013 M.n912 M.n911 2.2505
R4014 M.n910 M.n909 2.2505
R4015 M.n905 M.n904 2.2505
R4016 M.n916 M.n915 2.2505
R4017 M.n924 M.n923 2.2505
R4018 M.n897 M.n896 2.2505
R4019 M.n749 M.n748 2.2505
R4020 M.n737 M.n736 2.2505
R4021 M.n724 M.n723 2.2505
R4022 M.n745 M.n744 2.2505
R4023 M.n583 M.n582 2.2505
R4024 M.n733 M.n732 2.2505
R4025 M.n587 M.n581 2.2505
R4026 M.n729 M.n728 2.2505
R4027 M.n741 M.n740 2.2505
R4028 M.n413 M.n409 2.2505
R4029 M.n420 M.n407 2.2505
R4030 M.n431 M.n404 2.2505
R4031 M.n424 M.n405 2.2505
R4032 M.n416 M.n408 2.2505
R4033 M.n432 M.n402 2.2505
R4034 M.n422 M.n406 2.2505
R4035 M.n437 M.n401 2.2505
R4036 M.n1174 M.n1173 1.16276
R4037 M.n1175 M.n1174 1.16276
R4038 M.n1176 M.n1175 1.16276
R4039 M.n1177 M.n1176 1.16276
R4040 M.n1178 M.n1177 1.16276
R4041 M.n1179 M.n1178 1.16276
R4042 M.n1180 M.n1179 1.16276
R4043 M.n1181 M.n1180 1.16276
R4044 M.n1182 M.n1181 1.16276
R4045 M.n1183 M.n1182 1.16276
R4046 M.n1163 M.n1162 1.16276
R4047 M.n1164 M.n1163 1.16276
R4048 M.n1165 M.n1164 1.16276
R4049 M.n1166 M.n1165 1.16276
R4050 M.n1167 M.n1166 1.16276
R4051 M.n1168 M.n1167 1.16276
R4052 M.n1169 M.n1168 1.16276
R4053 M.n1170 M.n1169 1.16276
R4054 M.n1171 M.n1170 1.16276
R4055 M.n1172 M.n1171 1.16276
R4056 M.n1152 M.n1151 1.16276
R4057 M.n1153 M.n1152 1.16276
R4058 M.n1154 M.n1153 1.16276
R4059 M.n1155 M.n1154 1.16276
R4060 M.n1156 M.n1155 1.16276
R4061 M.n1157 M.n1156 1.16276
R4062 M.n1158 M.n1157 1.16276
R4063 M.n1159 M.n1158 1.16276
R4064 M.n1160 M.n1159 1.16276
R4065 M.n1161 M.n1160 1.16276
R4066 M.n1127 M.n1126 1.16276
R4067 M.n1128 M.n1127 1.16276
R4068 M.n1129 M.n1128 1.16276
R4069 M.n1130 M.n1129 1.16276
R4070 M.n1131 M.n1130 1.16276
R4071 M.n1132 M.n1131 1.16276
R4072 M.n1133 M.n1132 1.16276
R4073 M.n1134 M.n1133 1.16276
R4074 M.n1135 M.n1134 1.16276
R4075 M.n1136 M.n1135 1.16276
R4076 M.n1116 M.n1115 1.16276
R4077 M.n1117 M.n1116 1.16276
R4078 M.n1118 M.n1117 1.16276
R4079 M.n1119 M.n1118 1.16276
R4080 M.n1120 M.n1119 1.16276
R4081 M.n1121 M.n1120 1.16276
R4082 M.n1122 M.n1121 1.16276
R4083 M.n1123 M.n1122 1.16276
R4084 M.n1124 M.n1123 1.16276
R4085 M.n1125 M.n1124 1.16276
R4086 M.n45 M.n44 1.16276
R4087 M.n46 M.n45 1.16276
R4088 M.n47 M.n46 1.16276
R4089 M.n48 M.n47 1.16276
R4090 M.n49 M.n48 1.16276
R4091 M.n50 M.n49 1.16276
R4092 M.n51 M.n50 1.16276
R4093 M.n52 M.n51 1.16276
R4094 M.n53 M.n52 1.16276
R4095 M.n54 M.n53 1.16276
R4096 M.n56 M.n55 1.16276
R4097 M.n57 M.n56 1.16276
R4098 M.n58 M.n57 1.16276
R4099 M.n59 M.n58 1.16276
R4100 M.n60 M.n59 1.16276
R4101 M.n61 M.n60 1.16276
R4102 M.n62 M.n61 1.16276
R4103 M.n63 M.n62 1.16276
R4104 M.n64 M.n63 1.16276
R4105 M.n65 M.n64 1.16276
R4106 M.n34 M.n33 1.16276
R4107 M.n35 M.n34 1.16276
R4108 M.n36 M.n35 1.16276
R4109 M.n37 M.n36 1.16276
R4110 M.n38 M.n37 1.16276
R4111 M.n39 M.n38 1.16276
R4112 M.n40 M.n39 1.16276
R4113 M.n41 M.n40 1.16276
R4114 M.n42 M.n41 1.16276
R4115 M.n43 M.n42 1.16276
R4116 M.n23 M.n22 1.16276
R4117 M.n24 M.n23 1.16276
R4118 M.n25 M.n24 1.16276
R4119 M.n26 M.n25 1.16276
R4120 M.n27 M.n26 1.16276
R4121 M.n28 M.n27 1.16276
R4122 M.n29 M.n28 1.16276
R4123 M.n30 M.n29 1.16276
R4124 M.n31 M.n30 1.16276
R4125 M.n32 M.n31 1.16276
R4126 M.n12 M.n11 1.16276
R4127 M.n13 M.n12 1.16276
R4128 M.n14 M.n13 1.16276
R4129 M.n15 M.n14 1.16276
R4130 M.n16 M.n15 1.16276
R4131 M.n17 M.n16 1.16276
R4132 M.n18 M.n17 1.16276
R4133 M.n19 M.n18 1.16276
R4134 M.n20 M.n19 1.16276
R4135 M.n21 M.n20 1.16276
R4136 M.n1 M.n0 1.16276
R4137 M.n2 M.n1 1.16276
R4138 M.n3 M.n2 1.16276
R4139 M.n4 M.n3 1.16276
R4140 M.n5 M.n4 1.16276
R4141 M.n6 M.n5 1.16276
R4142 M.n7 M.n6 1.16276
R4143 M.n8 M.n7 1.16276
R4144 M.n9 M.n8 1.16276
R4145 M.n10 M.n9 1.16276
R4146 M.n205 M.n204 1.13934
R4147 M.n1295 M.n1294 1.12652
R4148 M.n1150 M.n1149 1.1255
R4149 M.n1316 M.n1315 1.1255
R4150 M.n1414 M.n1410 1.1255
R4151 M.n1448 M.n1443 1.1255
R4152 M.n1502 M.n1499 1.1255
R4153 M.n1371 M.n1370 1.1255
R4154 M.n1349 M.n1347 1.1255
R4155 M.n1386 M.n1385 1.1255
R4156 M.n1402 M.n1399 1.1255
R4157 M.n1435 M.n1434 1.1255
R4158 M.n1436 M.n1435 1.1255
R4159 M.n1403 M.n1402 1.1255
R4160 M.n1369 M.n1368 1.1255
R4161 M.n1368 M.n1367 1.1255
R4162 M.n1465 M.n1460 1.1255
R4163 M.n1425 M.n1424 1.1255
R4164 M.n1426 M.n1425 1.1255
R4165 M.n1466 M.n1465 1.1255
R4166 M.n1387 M.n1386 1.1255
R4167 M.n1350 M.n1349 1.1255
R4168 M.n1372 M.n1371 1.1255
R4169 M.n1503 M.n1502 1.1255
R4170 M.n1449 M.n1448 1.1255
R4171 M.n1415 M.n1414 1.1255
R4172 M.n1527 M.n1525 1.1255
R4173 M.n1579 M.n1578 1.1255
R4174 M.n1620 M.n1619 1.1255
R4175 M.n1665 M.n1662 1.1255
R4176 M.n1609 M.n1604 1.1255
R4177 M.n1569 M.n1568 1.1255
R4178 M.n1595 M.n1592 1.1255
R4179 M.n1554 M.n1553 1.1255
R4180 M.n1555 M.n1554 1.1255
R4181 M.n1596 M.n1595 1.1255
R4182 M.n1635 M.n1634 1.1255
R4183 M.n1634 M.n1633 1.1255
R4184 M.n1543 M.n1537 1.1255
R4185 M.n1544 M.n1543 1.1255
R4186 M.n1570 M.n1569 1.1255
R4187 M.n1610 M.n1609 1.1255
R4188 M.n1666 M.n1665 1.1255
R4189 M.n1621 M.n1620 1.1255
R4190 M.n1580 M.n1579 1.1255
R4191 M.n1528 M.n1527 1.1255
R4192 M.n1702 M.n1150 1.1255
R4193 M.n1825 M.n1822 1.1255
R4194 M.n1743 M.n1740 1.1255
R4195 M.n1678 M.n1676 1.1255
R4196 M.n1771 M.n1768 1.1255
R4197 M.n1697 M.n1690 1.1255
R4198 M.n1701 M.n1700 1.1255
R4199 M.n1700 M.n1699 1.1255
R4200 M.n1788 M.n1787 1.1255
R4201 M.n1787 M.n1786 1.1255
R4202 M.n1731 M.n1730 1.1255
R4203 M.n1732 M.n1731 1.1255
R4204 M.n1698 M.n1697 1.1255
R4205 M.n1772 M.n1771 1.1255
R4206 M.n1761 M.n1760 1.1255
R4207 M.n1762 M.n1761 1.1255
R4208 M.n1802 M.n1801 1.1255
R4209 M.n1801 M.n1800 1.1255
R4210 M.n1679 M.n1678 1.1255
R4211 M.n1744 M.n1743 1.1255
R4212 M.n1826 M.n1825 1.1255
R4213 M.n1869 M.n1862 1.1255
R4214 M.n1916 M.n1915 1.1255
R4215 M.n1951 M.n1946 1.1255
R4216 M.n2003 M.n2000 1.1255
R4217 M.n1850 M.n1848 1.1255
R4218 M.n1887 M.n1886 1.1255
R4219 M.n1872 M.n1871 1.1255
R4220 M.n1926 M.n1925 1.1255
R4221 M.n1968 M.n1967 1.1255
R4222 M.n1967 M.n1966 1.1255
R4223 M.n1940 M.n1939 1.1255
R4224 M.n1939 M.n1938 1.1255
R4225 M.n1904 M.n1903 1.1255
R4226 M.n1903 M.n1902 1.1255
R4227 M.n1873 M.n1872 1.1255
R4228 M.n1927 M.n1926 1.1255
R4229 M.n1888 M.n1887 1.1255
R4230 M.n1851 M.n1850 1.1255
R4231 M.n2004 M.n2003 1.1255
R4232 M.n1952 M.n1951 1.1255
R4233 M.n1917 M.n1916 1.1255
R4234 M.n1870 M.n1869 1.1255
R4235 M.n768 M.n767 1.1255
R4236 M.n303 M.n302 1.1255
R4237 M.n238 M.n236 1.1255
R4238 M.n175 M.n174 1.1255
R4239 M.n93 M.n92 1.1255
R4240 M.n120 M.n116 1.1255
R4241 M.n160 M.n155 1.1255
R4242 M.n161 M.n160 1.1255
R4243 M.n121 M.n120 1.1255
R4244 M.n81 M.n80 1.1255
R4245 M.n80 M.n79 1.1255
R4246 M.n72 M.n71 1.1255
R4247 M.n150 M.n149 1.1255
R4248 M.n149 M.n148 1.1255
R4249 M.n109 M.n108 1.1255
R4250 M.n110 M.n109 1.1255
R4251 M.n73 M.n72 1.1255
R4252 M.n187 M.n186 1.1255
R4253 M.n186 M.n185 1.1255
R4254 M.n131 M.n130 1.1255
R4255 M.n94 M.n93 1.1255
R4256 M.n132 M.n131 1.1255
R4257 M.n176 M.n175 1.1255
R4258 M.n239 M.n238 1.1255
R4259 M.n566 M.n565 1.1255
R4260 M.n538 M.n533 1.1255
R4261 M.n575 M.n571 1.1255
R4262 M.n522 M.n521 1.1255
R4263 M.n479 M.n478 1.1255
R4264 M.n518 M.n515 1.1255
R4265 M.n482 M.n481 1.1255
R4266 M.n483 M.n482 1.1255
R4267 M.n519 M.n518 1.1255
R4268 M.n549 M.n548 1.1255
R4269 M.n548 M.n547 1.1255
R4270 M.n497 M.n496 1.1255
R4271 M.n461 M.n460 1.1255
R4272 M.n460 M.n459 1.1255
R4273 M.n443 M.n442 1.1255
R4274 M.n444 M.n443 1.1255
R4275 M.n480 M.n479 1.1255
R4276 M.n523 M.n522 1.1255
R4277 M.n576 M.n575 1.1255
R4278 M.n498 M.n497 1.1255
R4279 M.n539 M.n538 1.1255
R4280 M.n567 M.n566 1.1255
R4281 M.n711 M.n710 1.1255
R4282 M.n674 M.n673 1.1255
R4283 M.n635 M.n630 1.1255
R4284 M.n593 M.n592 1.1255
R4285 M.n756 M.n754 1.1255
R4286 M.n685 M.n684 1.1255
R4287 M.n698 M.n697 1.1255
R4288 M.n609 M.n608 1.1255
R4289 M.n608 M.n607 1.1255
R4290 M.n645 M.n644 1.1255
R4291 M.n646 M.n645 1.1255
R4292 M.n625 M.n624 1.1255
R4293 M.n624 M.n623 1.1255
R4294 M.n665 M.n664 1.1255
R4295 M.n664 M.n663 1.1255
R4296 M.n699 M.n698 1.1255
R4297 M.n686 M.n685 1.1255
R4298 M.n757 M.n756 1.1255
R4299 M.n594 M.n593 1.1255
R4300 M.n636 M.n635 1.1255
R4301 M.n675 M.n674 1.1255
R4302 M.n712 M.n711 1.1255
R4303 M.n792 M.n791 1.1255
R4304 M.n885 M.n884 1.1255
R4305 M.n935 M.n933 1.1255
R4306 M.n867 M.n866 1.1255
R4307 M.n870 M.n869 1.1255
R4308 M.n833 M.n828 1.1255
R4309 M.n823 M.n822 1.1255
R4310 M.n780 M.n779 1.1255
R4311 M.n779 M.n778 1.1255
R4312 M.n806 M.n805 1.1255
R4313 M.n805 M.n804 1.1255
R4314 M.n848 M.n847 1.1255
R4315 M.n847 M.n846 1.1255
R4316 M.n871 M.n870 1.1255
R4317 M.n824 M.n823 1.1255
R4318 M.n868 M.n867 1.1255
R4319 M.n936 M.n935 1.1255
R4320 M.n834 M.n833 1.1255
R4321 M.n886 M.n885 1.1255
R4322 M.n793 M.n792 1.1255
R4323 M.n1070 M.n980 1.1255
R4324 M.n1060 M.n1059 1.1255
R4325 M.n1036 M.n986 1.1255
R4326 M.n1065 M.n985 1.1255
R4327 M.n1050 M.n1049 1.1255
R4328 M.n1028 M.n1027 1.1255
R4329 M.n1008 M.n1007 1.1255
R4330 M.n1112 M.n1110 1.1255
R4331 M.n1113 M.n1112 1.1255
R4332 M.n1010 M.n1009 1.1255
R4333 M.n1035 M.n992 1.1255
R4334 M.n1006 M.n1005 1.1255
R4335 M.n770 M.n769 1.12274
R4336 M.n1072 M.n1071 0.96098
R4337 M.n932 M.n931 0.900727
R4338 M.n753 M.n752 0.900727
R4339 M.n235 M.n234 0.900727
R4340 M.n1847 M.n1846 0.900647
R4341 M.n1730 M.n1726 0.9005
R4342 M.n1760 M.n1759 0.9005
R4343 M.n441 M.n440 0.900483
R4344 M.n1346 M.n1345 0.900467
R4345 M.n1496 M.n1495 0.900443
R4346 M.n591 M.n590 0.900443
R4347 M.n1675 M.n1674 0.900387
R4348 M.n1524 M.n1523 0.900387
R4349 M.n1109 M.n1108 0.900368
R4350 M.n1997 M.n1996 0.900365
R4351 M.n1819 M.n1818 0.900365
R4352 M.n1659 M.n1658 0.900365
R4353 M.n975 M.n974 0.900347
R4354 M.n766 M.n765 0.898241
R4355 M.n1893 M.n1125 0.615498
R4356 M.n1733 M.n1136 0.614262
R4357 M.n1571 M.n1161 0.609999
R4358 M.n383 M.n54 0.609008
R4359 M.n850 M.n21 0.608439
R4360 M.n111 M.n65 0.606848
R4361 M.n1392 M.n1172 0.606843
R4362 M.n649 M.n32 0.606489
R4363 M.n504 M.n43 0.605607
R4364 M.n1091 M.n10 0.601243
R4365 M.n1191 M.n1183 0.593624
R4366 M.n1317 M.n1316 0.563
R4367 M.n1318 M.n1317 0.563
R4368 M.n1319 M.n1318 0.563
R4369 M.n339 M.n303 0.563
R4370 M.n375 M.n339 0.563
R4371 M.n376 M.n375 0.563
R4372 M.n579 M.n578 0.473104
R4373 M.n1505 M.n1504 0.467151
R4374 M.n399 M.n398 0.465504
R4375 M.n1072 M.n937 0.458913
R4376 M.n1668 M.n1667 0.456584
R4377 M.n1828 M.n1827 0.451624
R4378 M.n1327 M.n1326 0.449946
R4379 M.n772 M.n758 0.443676
R4380 M.n241 M.n240 0.441768
R4381 M M.n2005 0.307487
R4382 M M.n1114 0.145448
R4383 M.n772 M.n771 0.0326212
R4384 M.n1315 M.n1314 0.0289279
R4385 M.n302 M.n296 0.028625
R4386 M.n1845 M.n1844 0.0262358
R4387 M.n1315 M.n1311 0.0249978
R4388 M.n761 M.n760 0.0243636
R4389 M.n199 M.n198 0.0233924
R4390 M.n765 M.n764 0.023
R4391 M.n767 M.n763 0.023
R4392 M.n930 M.n929 0.0228692
R4393 M.n301 M.n300 0.0228692
R4394 M.n1073 M.n1072 0.0203706
R4395 M.n1310 M.n1309 0.0201507
R4396 M.n273 M.n272 0.0198605
R4397 M.n1344 M.n1343 0.0195988
R4398 M.n1283 M.n1282 0.0193646
R4399 M.n266 M.n265 0.0190756
R4400 M.n1657 M.n1656 0.0190117
R4401 M.n233 M.n232 0.0189448
R4402 M.n1241 M.n1240 0.0185786
R4403 M.n255 M.n254 0.0182907
R4404 M.n298 M.n297 0.0176366
R4405 M.n773 M.n772 0.0164954
R4406 M.n1290 M.n1289 0.0162205
R4407 M.n436 M.n435 0.0160669
R4408 M.n956 M.n955 0.0155517
R4409 M.n1252 M.n1251 0.0154345
R4410 M.n1725 M.n1724 0.0153997
R4411 M.n1514 M.n1513 0.0152492
R4412 M.n202 M.n201 0.0150203
R4413 M.n427 M.n426 0.0148895
R4414 M.n1211 M.n1210 0.0146485
R4415 M.n227 M.n226 0.0146279
R4416 M.n1025 M.n1024 0.0146207
R4417 M.n973 M.n972 0.0144655
R4418 M.n292 M.n291 0.0141047
R4419 M.n1995 M.n1994 0.0140452
R4420 M.n1301 M.n1300 0.0137314
R4421 M.n1017 M.n1016 0.0136897
R4422 M.n978 M.n977 0.0135345
R4423 M.n332 M.n331 0.0133198
R4424 M.n771 M.n770 0.0132273
R4425 M.n918 M.n917 0.013189
R4426 M.n1268 M.n1267 0.0129454
R4427 M.n1068 M.n1067 0.0126034
R4428 M.n368 M.n367 0.0125349
R4429 M.n1226 M.n1225 0.0121594
R4430 M.n1817 M.n1816 0.0117876
R4431 M.n1853 M.n1852 0.0111355
R4432 M.n1494 M.n1493 0.0105727
R4433 M.n1754 M.n1753 0.0104331
R4434 M.n1648 M.n1647 0.0104331
R4435 M.n204 M.n203 0.0100494
R4436 M.n890 M.n889 0.00974419
R4437 M.n201 M.n200 0.00939535
R4438 M.n418 M.n417 0.00926454
R4439 M.n283 M.n282 0.00887209
R4440 M.n1485 M.n1484 0.00861047
R4441 M.n1102 M.n1101 0.00855063
R4442 M.n246 M.n245 0.00840698
R4443 M.n1201 M.n1200 0.00838571
R4444 M.n1352 M.n1351 0.0082907
R4445 M.n586 M.n585 0.00808721
R4446 M.n318 M.n317 0.00808721
R4447 M.n190 M.n189 0.00797826
R4448 M.n967 M.n966 0.00794828
R4449 M.n1989 M.n1988 0.00772408
R4450 M.n1654 M.n1653 0.00757358
R4451 M.n1637 M.n1636 0.00748113
R4452 M.n769 M.n768 0.00743292
R4453 M.n1681 M.n1680 0.0073277
R4454 M.n619 M.n618 0.00730233
R4455 M.n354 M.n353 0.00730233
R4456 M.n1057 M.n1056 0.00701724
R4457 M.n964 M.n963 0.00686207
R4458 M.n903 M.n902 0.00677907
R4459 M.n463 M.n462 0.00668497
R4460 M.n1321 M.n1320 0.00667143
R4461 M.n1985 M.n1984 0.00667057
R4462 M.n970 M.n969 0.00655172
R4463 M.n614 M.n613 0.00651744
R4464 M.n1992 M.n1991 0.00636957
R4465 M.n218 M.n217 0.00625581
R4466 M.n1070 M.n1069 0.00624138
R4467 M.n1065 M.n1064 0.00624138
R4468 M.n1060 M.n1054 0.00624138
R4469 M.n1050 M.n1042 0.00624138
R4470 M.n1028 M.n1018 0.00624138
R4471 M.n1112 M.n1111 0.00624138
R4472 M.n1892 M.n1891 0.00618562
R4473 M.n502 M.n501 0.00616474
R4474 M.n1706 M.n1705 0.00610386
R4475 M.n1066 M.n1065 0.00608621
R4476 M.n1061 M.n1060 0.00608621
R4477 M.n1053 M.n1052 0.00608621
R4478 M.n1051 M.n1050 0.00608621
R4479 M.n1112 M.n1104 0.00608621
R4480 M.n2003 M.n2002 0.00606856
R4481 M.n1967 M.n1960 0.00606856
R4482 M.n1951 M.n1950 0.00606856
R4483 M.n1939 M.n1933 0.00606856
R4484 M.n1903 M.n1897 0.00606856
R4485 M.n1850 M.n1849 0.00606856
R4486 M.n1825 M.n1824 0.00606856
R4487 M.n1771 M.n1770 0.00606856
R4488 M.n1678 M.n1677 0.00606856
R4489 M.n1665 M.n1664 0.00606856
R4490 M.n1634 M.n1628 0.00606856
R4491 M.n1527 M.n1526 0.00606856
R4492 M.n164 M.n163 0.00606522
R4493 M.n802 M.n801 0.00599419
R4494 M.n302 M.n301 0.00599419
R4495 M.n1047 M.n1046 0.00593103
R4496 M.n2003 M.n1971 0.00591806
R4497 M.n1967 M.n1956 0.00591806
R4498 M.n1949 M.n1948 0.00591806
R4499 M.n1850 M.n1830 0.00591806
R4500 M.n1825 M.n1805 0.00591806
R4501 M.n1801 M.n1792 0.00591806
R4502 M.n1678 M.n1670 0.00591806
R4503 M.n1665 M.n1638 0.00591806
R4504 M.n1634 M.n1626 0.00591806
R4505 M.n1595 M.n1585 0.00591806
R4506 M.n1558 M.n1557 0.0059088
R4507 M.n907 M.n906 0.00586337
R4508 M.n381 M.n380 0.00584884
R4509 M.n974 M.n973 0.00577586
R4510 M.n971 M.n970 0.00577586
R4511 M.n968 M.n967 0.00577586
R4512 M.n965 M.n964 0.00577586
R4513 M.n957 M.n956 0.00577586
R4514 M.n980 M.n979 0.00577586
R4515 M.n985 M.n984 0.00577586
R4516 M.n1059 M.n1058 0.00577586
R4517 M.n1049 M.n1048 0.00577586
R4518 M.n1027 M.n1026 0.00577586
R4519 M.n1970 M.n1969 0.00571739
R4520 M.n972 M.n971 0.00562069
R4521 M.n969 M.n968 0.00562069
R4522 M.n966 M.n965 0.00562069
R4523 M.n1108 M.n1107 0.00562069
R4524 M.n983 M.n982 0.00562069
R4525 M.n1110 M.n1106 0.00562069
R4526 M.n1996 M.n1995 0.00561706
R4527 M.n1993 M.n1992 0.00561706
R4528 M.n1990 M.n1989 0.00561706
R4529 M.n1987 M.n1985 0.00561706
R4530 M.n1976 M.n1975 0.00561706
R4531 M.n2000 M.n1999 0.00561706
R4532 M.n1966 M.n1965 0.00561706
R4533 M.n1946 M.n1945 0.00561706
R4534 M.n1938 M.n1937 0.00561706
R4535 M.n1902 M.n1901 0.00561706
R4536 M.n1818 M.n1817 0.00561706
R4537 M.n1726 M.n1725 0.00561706
R4538 M.n1822 M.n1821 0.00561706
R4539 M.n1768 M.n1767 0.00561706
R4540 M.n1658 M.n1657 0.00561706
R4541 M.n1655 M.n1654 0.00561706
R4542 M.n1662 M.n1661 0.00561706
R4543 M.n1633 M.n1632 0.00561706
R4544 M.n899 M.n898 0.00560174
R4545 M.n767 M.n766 0.00559846
R4546 M.n1994 M.n1993 0.00546656
R4547 M.n1991 M.n1990 0.00546656
R4548 M.n1988 M.n1987 0.00546656
R4549 M.n1846 M.n1845 0.00546656
R4550 M.n1966 M.n1962 0.00546656
R4551 M.n1964 M.n1963 0.00546656
R4552 M.n1946 M.n1943 0.00546656
R4553 M.n1938 M.n1935 0.00546656
R4554 M.n1848 M.n1832 0.00546656
R4555 M.n1758 M.n1757 0.00546656
R4556 M.n1816 M.n1815 0.00546656
R4557 M.n1759 M.n1754 0.00546656
R4558 M.n1759 M.n1756 0.00546656
R4559 M.n1674 M.n1673 0.00546656
R4560 M.n1800 M.n1796 0.00546656
R4561 M.n1676 M.n1672 0.00546656
R4562 M.n1656 M.n1655 0.00546656
R4563 M.n1647 M.n1646 0.00546656
R4564 M.n1633 M.n1630 0.00546656
R4565 M.n1592 M.n1587 0.00546656
R4566 M.n1191 M.n1190 0.00541429
R4567 M.n850 M.n849 0.00538372
R4568 M.n1209 M.n1208 0.00534716
R4569 M.n1318 M.n1242 0.00534716
R4570 M.n1502 M.n1501 0.00534012
R4571 M.n1435 M.n1431 0.00534012
R4572 M.n1402 M.n1401 0.00534012
R4573 M.n1349 M.n1348 0.00534012
R4574 M.n847 M.n841 0.00534012
R4575 M.n935 M.n934 0.00534012
R4576 M.n608 M.n601 0.00534012
R4577 M.n756 M.n755 0.00534012
R4578 M.n460 M.n452 0.00534012
R4579 M.n299 M.n298 0.00534012
R4580 M.n370 M.n369 0.00534012
R4581 M.n351 M.n350 0.00534012
R4582 M.n238 M.n237 0.00534012
R4583 M.n760 M.n759 0.00527273
R4584 M.n1203 M.n1202 0.00521616
R4585 M.n1318 M.n1212 0.00521616
R4586 M.n1502 M.n1469 0.0052093
R4587 M.n1465 M.n1453 0.0052093
R4588 M.n1349 M.n1329 0.0052093
R4589 M.n779 M.n775 0.0052093
R4590 M.n792 M.n786 0.0052093
R4591 M.n798 M.n797 0.0052093
R4592 M.n805 M.n799 0.0052093
R4593 M.n935 M.n892 0.0052093
R4594 M.n593 M.n580 0.0052093
R4595 M.n608 M.n600 0.0052093
R4596 M.n698 M.n692 0.0052093
R4597 M.n443 M.n400 0.0052093
R4598 M.n548 M.n544 0.0052093
R4599 M.n248 M.n247 0.0052093
R4600 M.n253 M.n252 0.0052093
R4601 M.n375 M.n256 0.0052093
R4602 M.n352 M.n351 0.0052093
R4603 M.n93 M.n88 0.0052093
R4604 M.n131 M.n127 0.0052093
R4605 M.n238 M.n192 0.0052093
R4606 M.n1729 M.n1728 0.00516555
R4607 M.n1710 M.n1709 0.00516555
R4608 M.n818 M.n817 0.00507849
R4609 M.n711 M.n705 0.00507849
R4610 M.n460 M.n450 0.00507849
R4611 M.n209 M.n208 0.00507849
R4612 M.n1752 M.n1751 0.00501505
R4613 M.n1748 M.n1747 0.00501505
R4614 M.n1041 M.n1040 0.005
R4615 M.n1289 M.n1288 0.00495415
R4616 M.n1316 M.n1310 0.00495415
R4617 M.n1250 M.n1249 0.00495415
R4618 M.n1317 M.n1284 0.00495415
R4619 M.n1495 M.n1494 0.00494767
R4620 M.n1492 M.n1491 0.00494767
R4621 M.n1486 M.n1485 0.00494767
R4622 M.n1476 M.n1475 0.00494767
R4623 M.n1499 M.n1498 0.00494767
R4624 M.n1434 M.n1433 0.00494767
R4625 M.n1399 M.n1398 0.00494767
R4626 M.n898 M.n897 0.00494767
R4627 M.n902 M.n901 0.00494767
R4628 M.n906 M.n905 0.00494767
R4629 M.n917 M.n916 0.00494767
R4630 M.n846 M.n845 0.00494767
R4631 M.n590 M.n589 0.00494767
R4632 M.n587 M.n586 0.00494767
R4633 M.n730 M.n729 0.00494767
R4634 M.n742 M.n741 0.00494767
R4635 M.n746 M.n745 0.00494767
R4636 M.n607 M.n606 0.00494767
R4637 M.n440 M.n439 0.00494767
R4638 M.n437 M.n436 0.00494767
R4639 M.n416 M.n415 0.00494767
R4640 M.n459 M.n458 0.00494767
R4641 M.n272 M.n271 0.00494767
R4642 M.n293 M.n292 0.00494767
R4643 M.n284 M.n283 0.00494767
R4644 M.n281 M.n280 0.00494767
R4645 M.n264 M.n263 0.00494767
R4646 M.n334 M.n333 0.00494767
R4647 M.n320 M.n319 0.00494767
R4648 M.n315 M.n314 0.00494767
R4649 M.n250 M.n249 0.00494767
R4650 M.n356 M.n355 0.00494767
R4651 M.n211 M.n210 0.00494767
R4652 M.n220 M.n219 0.00494767
R4653 M.n1932 M.n1931 0.00486455
R4654 M.n1316 M.n1290 0.00482314
R4655 M.n1317 M.n1253 0.00482314
R4656 M.n1493 M.n1492 0.00481686
R4657 M.n1490 M.n1489 0.00481686
R4658 M.n1345 M.n1344 0.00481686
R4659 M.n1460 M.n1455 0.00481686
R4660 M.n1460 M.n1459 0.00481686
R4661 M.n1347 M.n1331 0.00481686
R4662 M.n897 M.n895 0.00481686
R4663 M.n901 M.n899 0.00481686
R4664 M.n905 M.n903 0.00481686
R4665 M.n931 M.n930 0.00481686
R4666 M.n778 M.n777 0.00481686
R4667 M.n789 M.n788 0.00481686
R4668 M.n791 M.n790 0.00481686
R4669 M.n804 M.n803 0.00481686
R4670 M.n933 M.n894 0.00481686
R4671 M.n588 M.n587 0.00481686
R4672 M.n731 M.n730 0.00481686
R4673 M.n733 M.n731 0.00481686
R4674 M.n745 M.n743 0.00481686
R4675 M.n749 M.n747 0.00481686
R4676 M.n607 M.n605 0.00481686
R4677 M.n697 M.n696 0.00481686
R4678 M.n710 M.n709 0.00481686
R4679 M.n438 M.n437 0.00481686
R4680 M.n417 M.n416 0.00481686
R4681 M.n414 M.n413 0.00481686
R4682 M.n459 M.n456 0.00481686
R4683 M.n547 M.n546 0.00481686
R4684 M.n303 M.n273 0.00481686
R4685 M.n282 M.n281 0.00481686
R4686 M.n339 M.n267 0.00481686
R4687 M.n316 M.n315 0.00481686
R4688 M.n210 M.n209 0.00481686
R4689 M.n219 M.n218 0.00481686
R4690 M.n234 M.n233 0.00481686
R4691 M.n92 M.n91 0.00481686
R4692 M.n130 M.n129 0.00481686
R4693 M.n236 M.n194 0.00481686
R4694 M.n186 M.n180 0.00481686
R4695 M.n1093 M.n1092 0.0048038
R4696 M.n1391 M.n1390 0.00474419
R4697 M.n1812 M.n1811 0.00471405
R4698 M.n1063 M.n1062 0.00468966
R4699 M.n735 M.n734 0.00468605
R4700 M.n661 M.n660 0.00468605
R4701 M.n655 M.n654 0.00468605
R4702 M.n412 M.n411 0.00468605
R4703 M.n563 M.n562 0.00468605
R4704 M.n570 M.n569 0.00468605
R4705 M.n557 M.n556 0.00468605
R4706 M.n573 M.n572 0.00468605
R4707 M.n126 M.n125 0.00468605
R4708 M.n175 M.n169 0.00468605
R4709 M.n1959 M.n1958 0.00456355
R4710 M.n1810 M.n1809 0.00456355
R4711 M.n1804 M.n1803 0.00455797
R4712 M.n373 M.n372 0.00455523
R4713 M.n1074 M.n1073 0.00444937
R4714 M.n1206 M.n1205 0.00443013
R4715 M.n1465 M.n1464 0.00442442
R4716 M.n750 M.n749 0.00442442
R4717 M.n231 M.n230 0.00442442
R4718 M.n185 M.n184 0.00442442
R4719 M.n1313 M.n1312 0.00429913
R4720 M.n1302 M.n1301 0.00429913
R4721 M.n1484 M.n1483 0.0042936
R4722 M.n1482 M.n1481 0.0042936
R4723 M.n812 M.n811 0.0042936
R4724 M.n585 M.n584 0.0042936
R4725 M.n752 M.n751 0.0042936
R4726 M.n279 M.n278 0.0042936
R4727 M.n308 M.n307 0.0042936
R4728 M.n344 M.n343 0.0042936
R4729 M.n208 M.n207 0.0042936
R4730 M.n229 M.n228 0.0042936
R4731 M.n90 M.n89 0.0042936
R4732 M.n174 M.n173 0.0042936
R4733 M.n1468 M.n1467 0.00427907
R4734 M.n1786 M.n1785 0.00426254
R4735 M.n270 M.n269 0.00416279
R4736 M.n261 M.n260 0.00416279
R4737 M.n160 M.n159 0.00416279
R4738 M.n1609 M.n1608 0.00411204
R4739 M.n1489 M.n1488 0.00403198
R4740 M.n785 M.n784 0.00403198
R4741 M.n589 M.n588 0.00403198
R4742 M.n659 M.n658 0.00403198
R4743 M.n203 M.n202 0.00403198
R4744 M.n213 M.n212 0.00403198
R4745 M.n215 M.n214 0.00403198
R4746 M.n217 M.n216 0.00403198
R4747 M.n149 M.n141 0.00403198
R4748 M.n1765 M.n1764 0.00397826
R4749 M.n1620 M.n1614 0.00396154
R4750 M.n1270 M.n1269 0.00390611
R4751 M.n1228 M.n1227 0.00390611
R4752 M.n1487 M.n1486 0.00390116
R4753 M.n1422 M.n1421 0.00390116
R4754 M.n1418 M.n1417 0.00390116
R4755 M.n621 M.n620 0.00390116
R4756 M.n754 M.n722 0.00390116
R4757 M.n616 M.n615 0.00390116
R4758 M.n311 M.n310 0.00390116
R4759 M.n305 M.n304 0.00390116
R4760 M.n347 M.n346 0.00390116
R4761 M.n341 M.n340 0.00390116
R4762 M.n69 M.n68 0.00390116
R4763 M.n77 M.n76 0.00390116
R4764 M.n1598 M.n1597 0.00389623
R4765 M.n1787 M.n1780 0.00381104
R4766 M.n1697 M.n1696 0.00381104
R4767 M.n300 M.n299 0.00377035
R4768 M.n295 M.n294 0.00377035
R4769 M.n291 M.n290 0.00377035
R4770 M.n289 M.n288 0.00377035
R4771 M.n286 M.n285 0.00377035
R4772 M.n337 M.n336 0.00377035
R4773 M.n327 M.n326 0.00377035
R4774 M.n225 M.n224 0.00377035
R4775 M.n155 M.n154 0.00377035
R4776 M.n542 M.n541 0.00367919
R4777 M.n1815 M.n1814 0.00366054
R4778 M.n1150 M.n1142 0.00366054
R4779 M.n1650 M.n1649 0.00366054
R4780 M.n1646 M.n1645 0.00366054
R4781 M.n1604 M.n1603 0.00366054
R4782 M.n1287 M.n1286 0.0036441
R4783 M.n1247 M.n1246 0.0036441
R4784 M.n1443 M.n1442 0.00363953
R4785 M.n738 M.n737 0.00363953
R4786 M.n223 M.n222 0.00363953
R4787 M.n106 M.n105 0.00363953
R4788 M.n114 M.n113 0.00363953
R4789 M.n148 M.n147 0.00363953
R4790 M.n118 M.n117 0.00363953
R4791 M.n390 M.n389 0.00352326
R4792 M.n1813 M.n1812 0.00351003
R4793 M.n1652 M.n1651 0.00351003
R4794 M.n1619 M.n1618 0.00351003
R4795 M.n1569 M.n1563 0.00351003
R4796 M.n1554 M.n1548 0.00351003
R4797 M.n1478 M.n1477 0.00350872
R4798 M.n741 M.n739 0.00350872
R4799 M.n756 M.n718 0.00350872
R4800 M.n419 M.n418 0.00350872
R4801 M.n280 M.n279 0.00350872
R4802 M.n363 M.n362 0.00350872
R4803 M.n87 M.n86 0.00350872
R4804 M.n1037 M.n1036 0.00344828
R4805 M.n1429 M.n1428 0.00340698
R4806 M.n330 M.n329 0.00337791
R4807 M.n322 M.n321 0.00337791
R4808 M.n366 M.n365 0.00337791
R4809 M.n358 M.n357 0.00337791
R4810 M.n1926 M.n1920 0.00335953
R4811 M.n1719 M.n1718 0.00335953
R4812 M.n1690 M.n1689 0.00335953
R4813 M.n1448 M.n1447 0.00324709
R4814 M.n604 M.n603 0.00324709
R4815 M.n653 M.n652 0.00324709
R4816 M.n101 M.n100 0.00324709
R4817 M.n763 M.n762 0.00322727
R4818 M.n1722 M.n1721 0.00320903
R4819 M.n1800 M.n1799 0.00320903
R4820 M.n1149 M.n1148 0.00320903
R4821 M.n1592 M.n1591 0.00320903
R4822 M.n2004 M.n1970 0.00317559
R4823 M.n1968 M.n1954 0.00317559
R4824 M.n1952 M.n1942 0.00317559
R4825 M.n1940 M.n1930 0.00317559
R4826 M.n1851 M.n1828 0.00317559
R4827 M.n611 M.n610 0.00315896
R4828 M.n945 M.n944 0.00313793
R4829 M.n963 M.n962 0.00313793
R4830 M.n961 M.n960 0.00313793
R4831 M.n960 M.n959 0.00313793
R4832 M.n959 M.n958 0.00313793
R4833 M.n955 M.n954 0.00313793
R4834 M.n952 M.n951 0.00313793
R4835 M.n948 M.n947 0.00313793
R4836 M.n1036 M.n1035 0.00313793
R4837 M.n1010 M.n1008 0.00313793
R4838 M.n1233 M.n1232 0.00312009
R4839 M.n729 M.n727 0.00311628
R4840 M.n743 M.n742 0.00311628
R4841 M.n684 M.n683 0.00311628
R4842 M.n531 M.n530 0.00311628
R4843 M.n536 M.n535 0.00311628
R4844 M.n2005 M.n2004 0.0031087
R4845 M.n1969 M.n1968 0.0031087
R4846 M.n1953 M.n1952 0.0031087
R4847 M.n1941 M.n1940 0.0031087
R4848 M.n1852 M.n1851 0.0031087
R4849 M.n1826 M.n1804 0.00307649
R4850 M.n1772 M.n1765 0.00307649
R4851 M.n1679 M.n1668 0.00307649
R4852 M.n1838 M.n1837 0.00305853
R4853 M.n1984 M.n1983 0.00305853
R4854 M.n1982 M.n1980 0.00305853
R4855 M.n1980 M.n1978 0.00305853
R4856 M.n1978 M.n1977 0.00305853
R4857 M.n1834 M.n1833 0.00305853
R4858 M.n1839 M.n1836 0.00305853
R4859 M.n1843 M.n1842 0.00305853
R4860 M.n1786 M.n1781 0.00305853
R4861 M.n1511 M.n1509 0.00305853
R4862 M.n1512 M.n1511 0.00305853
R4863 M.n1513 M.n1512 0.00305853
R4864 M.n1517 M.n1515 0.00305853
R4865 M.n1568 M.n1567 0.00305853
R4866 M.n1553 M.n1552 0.00305853
R4867 M.n67 M.n66 0.00304301
R4868 M.n1666 M.n1637 0.00301572
R4869 M.n1635 M.n1624 0.00301572
R4870 M.n1528 M.n1505 0.00301572
R4871 M.n1827 M.n1826 0.00301208
R4872 M.n1803 M.n1802 0.00301208
R4873 M.n1680 M.n1679 0.00301208
R4874 M.n1237 M.n1236 0.00298908
R4875 M.n1339 M.n1338 0.00298547
R4876 M.n1334 M.n1333 0.00298547
R4877 M.n1340 M.n1336 0.00298547
R4878 M.n1343 M.n1342 0.00298547
R4879 M.n823 M.n815 0.00298547
R4880 M.n672 M.n671 0.00298547
R4881 M.n962 M.n961 0.00298276
R4882 M.n958 M.n957 0.00298276
R4883 M.n1006 M.n998 0.00298276
R4884 M.n1667 M.n1666 0.00295283
R4885 M.n1636 M.n1635 0.00295283
R4886 M.n1597 M.n1596 0.00295283
R4887 M.n1848 M.n1847 0.00292012
R4888 M.n1983 M.n1982 0.00290803
R4889 M.n1977 M.n1976 0.00290803
R4890 M.n1925 M.n1924 0.00290803
R4891 M.n1869 M.n1868 0.00290803
R4892 M.n1515 M.n1514 0.00290803
R4893 M.n1519 M.n1517 0.00290803
R4894 M.n1522 M.n1521 0.00290803
R4895 M.n1578 M.n1577 0.00290803
R4896 M.n1942 M.n1941 0.00290803
R4897 M.n276 M.n275 0.0028968
R4898 M.n205 M.n196 0.0028968
R4899 M.n277 M.n276 0.00289361
R4900 M.n206 M.n205 0.00289361
R4901 M.n426 M.n425 0.00285465
R4902 M.n518 M.n508 0.00285465
R4903 M.n1893 M.n1892 0.00284114
R4904 M.n1011 M.n1010 0.00282759
R4905 M.n1503 M.n1468 0.00282558
R4906 M.n1436 M.n1429 0.00282558
R4907 M.n1350 M.n1327 0.00282558
R4908 M.n380 M.n379 0.00282558
R4909 M.n392 M.n391 0.00282558
R4910 M.n781 M.n780 0.00282558
R4911 M.n794 M.n793 0.00282558
R4912 M.n807 M.n806 0.00282558
R4913 M.n849 M.n848 0.00282558
R4914 M.n937 M.n936 0.00282558
R4915 M.n240 M.n239 0.00281884
R4916 M.n462 M.n461 0.00281214
R4917 M.n550 M.n549 0.00281214
R4918 M.n595 M.n594 0.00281214
R4919 M.n610 M.n609 0.00281214
R4920 M.n647 M.n646 0.00281214
R4921 M.n687 M.n686 0.00281214
R4922 M.n758 M.n757 0.00281214
R4923 M.n933 M.n932 0.00278682
R4924 M.n754 M.n753 0.00278682
R4925 M.n236 M.n235 0.00278682
R4926 M.n1322 M.n1321 0.00278571
R4927 M.n1319 M.n1201 0.00278571
R4928 M.n1504 M.n1503 0.00276744
R4929 M.n1467 M.n1466 0.00276744
R4930 M.n1351 M.n1350 0.00276744
R4931 M.n242 M.n241 0.00276744
R4932 M.n243 M.n242 0.00276744
R4933 M.n245 M.n244 0.00276744
R4934 M.n376 M.n246 0.00276744
R4935 M.n391 M.n390 0.00276744
R4936 M.n780 M.n773 0.00276744
R4937 M.n793 M.n782 0.00276744
R4938 M.n806 M.n795 0.00276744
R4939 M.n936 M.n890 0.00276744
R4940 M.n94 M.n84 0.00276087
R4941 M.n132 M.n124 0.00276087
R4942 M.n239 M.n190 0.00276087
R4943 M.n1887 M.n1879 0.00275752
R4944 M.n1801 M.n1794 0.00275752
R4945 M.n1595 M.n1594 0.00275752
R4946 M.n444 M.n399 0.00275434
R4947 M.n549 M.n542 0.00275434
R4948 M.n594 M.n579 0.00275434
R4949 M.n609 M.n596 0.00275434
R4950 M.n699 M.n688 0.00275434
R4951 M.n1326 M.n1325 0.00272857
R4952 M.n1320 M.n1319 0.00272857
R4953 M.n1314 M.n1313 0.00272707
R4954 M.n1309 M.n1308 0.00272707
R4955 M.n1305 M.n1304 0.00272707
R4956 M.n1275 M.n1274 0.00272707
R4957 M.n1217 M.n1216 0.00272707
R4958 M.n923 M.n922 0.00272384
R4959 M.n908 M.n907 0.00272384
R4960 M.n912 M.n910 0.00272384
R4961 M.n913 M.n912 0.00272384
R4962 M.n914 M.n913 0.00272384
R4963 M.n919 M.n918 0.00272384
R4964 M.n924 M.n921 0.00272384
R4965 M.n928 M.n927 0.00272384
R4966 M.n644 M.n643 0.00272384
R4967 M.n685 M.n680 0.00272384
R4968 M.n313 M.n312 0.00272384
R4969 M.n1624 M.n1623 0.00270126
R4970 M.n1707 M.n1706 0.00269002
R4971 M.n1045 M.n1044 0.00267241
R4972 M.n992 M.n991 0.00267241
R4973 M.n989 M.n988 0.00267241
R4974 M.n1023 M.n1022 0.00267241
R4975 M.n1003 M.n1002 0.00267241
R4976 M.n1039 M.n1038 0.00267241
R4977 M.n1031 M.n1030 0.00267241
R4978 M.n1015 M.n1014 0.00267241
R4979 M.n997 M.n996 0.00267241
R4980 M.n378 M.n377 0.00265116
R4981 M.n389 M.n388 0.00265116
R4982 M.n1764 M.n1763 0.0026256
R4983 M.n1071 M.n1070 0.00261022
R4984 M.n1923 M.n1922 0.00260702
R4985 M.n1915 M.n1914 0.00260702
R4986 M.n1882 M.n1881 0.00260702
R4987 M.n1860 M.n1859 0.00260702
R4988 M.n1919 M.n1918 0.00260702
R4989 M.n1876 M.n1875 0.00260702
R4990 M.n1867 M.n1866 0.00260702
R4991 M.n1787 M.n1776 0.00260702
R4992 M.n1566 M.n1565 0.00260702
R4993 M.n1579 M.n1575 0.00260702
R4994 M.n1562 M.n1561 0.00260702
R4995 M.n1308 M.n1307 0.00259607
R4996 M.n1299 M.n1298 0.00259607
R4997 M.n1279 M.n1278 0.00259607
R4998 M.n1260 M.n1259 0.00259607
R4999 M.n1220 M.n1219 0.00259607
R5000 M.n1218 M.n1217 0.00259607
R5001 M.n1383 M.n1382 0.00259302
R5002 M.n1363 M.n1362 0.00259302
R5003 M.n1377 M.n1376 0.00259302
R5004 M.n1357 M.n1356 0.00259302
R5005 M.n910 M.n908 0.00259302
R5006 M.n916 M.n914 0.00259302
R5007 M.n822 M.n821 0.00259302
R5008 M.n885 M.n877 0.00259302
R5009 M.n726 M.n725 0.00259302
R5010 M.n422 M.n421 0.00259302
R5011 M.n795 M.n794 0.00259302
R5012 M.n188 M.n187 0.00258696
R5013 M.n445 M.n444 0.00258092
R5014 M.n700 M.n699 0.00258092
R5015 M.n1324 M.n1323 0.00255714
R5016 M.n176 M.n165 0.00252899
R5017 M.n1076 M.n1075 0.00252532
R5018 M.n1079 M.n1078 0.00252532
R5019 M.n1082 M.n1081 0.00252532
R5020 M.n1114 M.n1113 0.00252532
R5021 M.n461 M.n446 0.00252312
R5022 M.n552 M.n551 0.00252312
R5023 M.n576 M.n567 0.00252312
R5024 M.n578 M.n577 0.00252312
R5025 M.n675 M.n665 0.00252312
R5026 M.n712 M.n701 0.00252312
R5027 M.n950 M.n948 0.00251724
R5028 M.n1005 M.n1004 0.00251724
R5029 M.n1075 M.n1074 0.00247468
R5030 M.n1078 M.n1077 0.00247468
R5031 M.n1081 M.n1080 0.00247468
R5032 M.n1091 M.n1090 0.00247468
R5033 M.n1113 M.n1102 0.00247468
R5034 M.n95 M.n94 0.00247101
R5035 M.n867 M.n859 0.00246221
R5036 M.n599 M.n598 0.00246221
R5037 M.n425 M.n424 0.00246221
R5038 M.n511 M.n510 0.00246221
R5039 M.n515 M.n512 0.00246221
R5040 M.n507 M.n506 0.00246221
R5041 M.n1842 M.n1841 0.00245652
R5042 M.n1902 M.n1899 0.00245652
R5043 M.n1862 M.n1861 0.00245652
R5044 M.n1814 M.n1813 0.00245652
R5045 M.n1724 M.n1723 0.00245652
R5046 M.n1721 M.n1720 0.00245652
R5047 M.n1718 M.n1717 0.00245652
R5048 M.n1798 M.n1797 0.00245652
R5049 M.n1653 M.n1652 0.00245652
R5050 M.n1651 M.n1650 0.00245652
R5051 M.n1649 M.n1648 0.00245652
R5052 M.n1645 M.n1644 0.00245652
R5053 M.n1590 M.n1589 0.00245652
R5054 M.n1551 M.n1550 0.00245652
R5055 M.n1533 M.n1532 0.00245652
R5056 M.n1547 M.n1546 0.00245652
R5057 M.n1541 M.n1540 0.00245652
R5058 M.n1539 M.n1538 0.00245652
R5059 M.n1930 M.n1929 0.0024398
R5060 M.n953 M.n952 0.00236207
R5061 M.n124 M.n123 0.00235507
R5062 M.n1293 M.n1292 0.00233406
R5063 M.n1281 M.n1280 0.00233406
R5064 M.n1259 M.n1258 0.00233406
R5065 M.n1239 M.n1238 0.00233406
R5066 M.n1368 M.n1360 0.0023314
R5067 M.n820 M.n819 0.0023314
R5068 M.n828 M.n827 0.0023314
R5069 M.n862 M.n861 0.0023314
R5070 M.n882 M.n881 0.0023314
R5071 M.n814 M.n813 0.0023314
R5072 M.n856 M.n855 0.0023314
R5073 M.n876 M.n875 0.0023314
R5074 M.n695 M.n694 0.0023314
R5075 M.n645 M.n641 0.0023314
R5076 M.n415 M.n414 0.0023314
R5077 M.n538 M.n537 0.0023314
R5078 M.n1080 M.n1079 0.00232278
R5079 M.n1836 M.n1835 0.00230602
R5080 M.n1886 M.n1885 0.00230602
R5081 M.n1779 M.n1778 0.00230602
R5082 M.n1954 M.n1953 0.00230602
R5083 M.n1762 M.n1745 0.00230354
R5084 M.n162 M.n161 0.0022971
R5085 M.n1214 M.n1213 0.00224426
R5086 M.n1466 M.n1451 0.00224419
R5087 M.n980 M.n975 0.00222181
R5088 M.n1035 M.n1034 0.0022069
R5089 M.n1307 M.n1306 0.00220306
R5090 M.n1298 M.n1297 0.00220306
R5091 M.n1264 M.n1263 0.00220306
R5092 M.n1262 M.n1261 0.00220306
R5093 M.n1255 M.n1254 0.00220306
R5094 M.n1222 M.n1221 0.00220306
R5095 M.n1446 M.n1445 0.00220058
R5096 M.n1386 M.n1378 0.00220058
R5097 M.n927 M.n926 0.00220058
R5098 M.n846 M.n843 0.00220058
R5099 M.n884 M.n883 0.00220058
R5100 M.n727 M.n726 0.00220058
R5101 M.n668 M.n667 0.00220058
R5102 M.n404 M.n403 0.00220058
R5103 M.n434 M.n433 0.00220058
R5104 M.n431 M.n430 0.00220058
R5105 M.n428 M.n427 0.00220058
R5106 M.n1610 M.n1599 0.00219811
R5107 M.n2000 M.n1997 0.00219111
R5108 M.n1822 M.n1819 0.00219111
R5109 M.n1662 M.n1659 0.00219111
R5110 M.n1450 M.n1449 0.00218605
R5111 M.n1428 M.n1427 0.00218605
R5112 M.n1426 M.n1415 0.00218605
R5113 M.n1405 M.n1404 0.00218605
R5114 M.n394 M.n393 0.00218605
R5115 M.n396 M.n395 0.00218605
R5116 M.n398 M.n397 0.00218605
R5117 M.n808 M.n807 0.00218605
R5118 M.n81 M.n73 0.00218116
R5119 M.n83 M.n82 0.00218116
R5120 M.n133 M.n132 0.00218116
R5121 M.n612 M.n611 0.0021763
R5122 M.n636 M.n625 0.0021763
R5123 M.n1193 M.n1192 0.00215714
R5124 M.n1916 M.n1911 0.00215552
R5125 M.n1520 M.n1519 0.00215552
R5126 M.n1622 M.n1621 0.00213522
R5127 M.n150 M.n135 0.00212319
R5128 M.n649 M.n648 0.0021185
R5129 M.n1790 M.n1789 0.00211031
R5130 M.n1698 M.n1683 0.00211031
R5131 M.n1304 M.n1303 0.00207205
R5132 M.n921 M.n920 0.00206977
R5133 M.n866 M.n865 0.00206977
R5134 M.n435 M.n434 0.00206977
R5135 M.n432 M.n431 0.00206977
R5136 M.n429 M.n428 0.00206977
R5137 M.n497 M.n489 0.00206977
R5138 M.n782 M.n781 0.00206977
R5139 M.n123 M.n122 0.00206522
R5140 M.n1244 M.n1243 0.0020629
R5141 M.n1499 M.n1496 0.00206165
R5142 M.n592 M.n591 0.00206165
R5143 M.n258 M.n257 0.00206165
R5144 M.n1110 M.n1109 0.0020532
R5145 M.n1029 M.n1028 0.00205172
R5146 M.n1295 M.n1293 0.00204803
R5147 M.n1296 M.n1295 0.00204706
R5148 M.n1703 M.n1702 0.00204589
R5149 M.n1676 M.n1675 0.00202155
R5150 M.n1525 M.n1524 0.00202155
R5151 M.n1903 M.n1895 0.00200502
R5152 M.n1145 M.n1144 0.00200502
R5153 M.n1688 M.n1687 0.00200502
R5154 M.n1139 M.n1138 0.00200502
R5155 M.n1695 M.n1694 0.00200502
R5156 M.n1523 M.n1522 0.00200502
R5157 M.n1617 M.n1616 0.00200502
R5158 M.n1602 M.n1601 0.00200502
R5159 M.n1613 M.n1612 0.00200502
R5160 M.n1607 M.n1606 0.00200502
R5161 M.n1928 M.n1927 0.00197157
R5162 M.n1083 M.n1082 0.00196835
R5163 M.n382 M.n381 0.00195349
R5164 M.n1570 M.n1559 0.00194654
R5165 M.n1556 M.n1555 0.00194654
R5166 M.n639 M.n638 0.00194509
R5167 M.n1341 M.n1340 0.00193895
R5168 M.n1367 M.n1366 0.00193895
R5169 M.n833 M.n832 0.00193895
R5170 M.n420 M.n419 0.00193895
R5171 M.n533 M.n532 0.00193895
R5172 M.n479 M.n471 0.00193895
R5173 M.n364 M.n363 0.00193895
R5174 M.n360 M.n359 0.00193895
R5175 M.n349 M.n348 0.00193895
R5176 M.n1788 M.n1774 0.00191707
R5177 M.n1347 M.n1346 0.00188813
R5178 M.n713 M.n712 0.00188728
R5179 M.n1077 M.n1076 0.00186709
R5180 M.n768 M.n761 0.00186364
R5181 M.n442 M.n441 0.00186205
R5182 M.n1773 M.n1772 0.00185266
R5183 M.n384 M.n383 0.00183721
R5184 M.n84 M.n83 0.00183333
R5185 M.n541 M.n540 0.00182948
R5186 M.n757 M.n714 0.00182948
R5187 M.n1196 M.n1195 0.00181429
R5188 M.n1286 M.n1285 0.00181004
R5189 M.n1278 M.n1277 0.00181004
R5190 M.n1477 M.n1476 0.00180814
R5191 M.n1335 M.n1334 0.00180814
R5192 M.n1385 M.n1384 0.00180814
R5193 M.n847 M.n839 0.00180814
R5194 M.n739 M.n738 0.00180814
R5195 M.n628 M.n627 0.00180814
R5196 M.n682 M.n681 0.00180814
R5197 M.n717 M.n716 0.00180814
R5198 M.n423 M.n422 0.00180814
R5199 M.n476 M.n475 0.00180814
R5200 M.n492 M.n491 0.00180814
R5201 M.n470 M.n469 0.00180814
R5202 M.n486 M.n485 0.00180814
R5203 M.n120 M.n119 0.00180814
R5204 M.n1392 M.n1391 0.00177907
R5205 M.n387 M.n386 0.00177907
R5206 M.n824 M.n809 0.00177907
R5207 M.n524 M.n523 0.00177168
R5208 M.n678 M.n677 0.00177168
R5209 M.n1870 M.n1855 0.0017709
R5210 M.n1199 M.n1198 0.00175714
R5211 M.n1449 M.n1438 0.00172093
R5212 M.n97 M.n96 0.00171739
R5213 M.n648 M.n647 0.00171387
R5214 M.n1537 M.n1536 0.00170401
R5215 M.n1889 M.n1888 0.00170401
R5216 M.n1531 M.n1530 0.00169497
R5217 M.n1288 M.n1287 0.00167904
R5218 M.n1273 M.n1272 0.00167904
R5219 M.n430 M.n429 0.00167733
R5220 M.n474 M.n473 0.00167733
R5221 M.n496 M.n495 0.00167733
R5222 M.n494 M.n493 0.00167733
R5223 M.n468 M.n467 0.00167733
R5224 M.n488 M.n487 0.00167733
R5225 M.n303 M.n295 0.00167733
R5226 M.n200 M.n199 0.00167733
R5227 M.n222 M.n221 0.00167733
R5228 M.n224 M.n223 0.00167733
R5229 M.n226 M.n225 0.00167733
R5230 M.n109 M.n102 0.00167733
R5231 M.n1437 M.n1436 0.00166279
R5232 M.n1774 M.n1773 0.00165942
R5233 M.n1734 M.n1733 0.00165942
R5234 M.n519 M.n504 0.00165607
R5235 M.n1185 M.n1184 0.00164286
R5236 M.n1929 M.n1928 0.00163712
R5237 M.n1927 M.n1917 0.00163712
R5238 M.n1906 M.n1905 0.00163712
R5239 M.n1891 M.n1890 0.00163712
R5240 M.n1888 M.n1873 0.00163712
R5241 M.n1855 M.n1854 0.00163712
R5242 M.n1085 M.n1084 0.00161392
R5243 M.n1438 M.n1437 0.00160465
R5244 M.n1389 M.n1388 0.00160465
R5245 M.n1372 M.n1369 0.00160465
R5246 M.n1353 M.n1352 0.00160465
R5247 M.n887 M.n886 0.00160465
R5248 M.n111 M.n110 0.00160145
R5249 M.n1188 M.n1187 0.00158571
R5250 M.n1583 M.n1582 0.00156918
R5251 M.n1559 M.n1558 0.00156918
R5252 M.n1521 M.n1520 0.00155351
R5253 M.n1535 M.n1534 0.00155351
R5254 M.n1525 M.n1507 0.00155351
R5255 M.n1230 M.n1229 0.00154803
R5256 M.n1403 M.n1392 0.00154651
R5257 M.n747 M.n746 0.00154651
R5258 M.n635 M.n634 0.00154651
R5259 M.n691 M.n690 0.00154651
R5260 M.n439 M.n438 0.00154651
R5261 M.n433 M.n432 0.00154651
R5262 M.n424 M.n423 0.00154651
R5263 M.n478 M.n477 0.00154651
R5264 M.n561 M.n560 0.00154651
R5265 M.n294 M.n293 0.00154651
R5266 M.n290 M.n289 0.00154651
R5267 M.n328 M.n327 0.00154651
R5268 M.n343 M.n342 0.00154651
R5269 M.n80 M.n75 0.00154651
R5270 M.n868 M.n853 0.00154651
R5271 M.n503 M.n502 0.00154046
R5272 M.n1557 M.n1556 0.00150629
R5273 M.n1555 M.n1544 0.00150629
R5274 M.n1530 M.n1529 0.00150629
R5275 M.n1369 M.n1354 0.00148837
R5276 M.n809 M.n808 0.00148837
R5277 M.n834 M.n824 0.00148837
R5278 M.n837 M.n836 0.00148837
R5279 M.n852 M.n851 0.00148837
R5280 M.n871 M.n868 0.00148837
R5281 M.n888 M.n887 0.00148837
R5282 M.n540 M.n539 0.00148266
R5283 M.n686 M.n678 0.00148266
R5284 M.n1200 M.n1199 0.00147143
R5285 M.n1802 M.n1790 0.00146618
R5286 M.n1099 M.n1098 0.00146203
R5287 M.n1596 M.n1583 0.0014434
R5288 M.n1580 M.n1571 0.0014434
R5289 M.n1033 M.n1032 0.00143104
R5290 M.n1388 M.n1387 0.00143023
R5291 M.n523 M.n520 0.00142485
R5292 M.n714 M.n713 0.00142485
R5293 M.n1245 M.n1244 0.00141703
R5294 M.n1236 M.n1235 0.00141703
R5295 M.n1234 M.n1233 0.00141703
R5296 M.n1488 M.n1487 0.0014157
R5297 M.n1441 M.n1440 0.0014157
R5298 M.n1399 M.n1396 0.0014157
R5299 M.n1425 M.n1419 0.0014157
R5300 M.n624 M.n617 0.0014157
R5301 M.n421 M.n420 0.0014157
R5302 M.n345 M.n344 0.0014157
R5303 M.n216 M.n215 0.0014157
R5304 M.n116 M.n115 0.0014157
R5305 M.n72 M.n67 0.0014157
R5306 M.n1189 M.n1188 0.00141429
R5307 M.n1186 M.n1185 0.00141429
R5308 M.n1096 M.n1095 0.00141139
R5309 M.n1910 M.n1909 0.00140301
R5310 M.n1811 M.n1810 0.00140301
R5311 M.n1784 M.n1783 0.00140301
R5312 M.n1789 M.n1788 0.00140177
R5313 M.n1581 M.n1580 0.0013805
R5314 M.n386 M.n385 0.00137209
R5315 M.n499 M.n498 0.00136705
R5316 M.n596 M.n595 0.00136705
R5317 M.n1084 M.n1083 0.00136076
R5318 M.n1086 M.n1085 0.00136076
R5319 M.n1089 M.n1088 0.00136076
R5320 M.n1094 M.n1093 0.00136076
R5321 M.n1097 M.n1096 0.00136076
R5322 M.n1100 M.n1099 0.00136076
R5323 M.n1705 M.n1704 0.00133736
R5324 M.n1702 M.n1701 0.00133736
R5325 M.n1683 M.n1682 0.00133736
R5326 M.n1623 M.n1622 0.00131761
R5327 M.n1621 M.n1610 0.00131761
R5328 M.n1599 M.n1598 0.00131761
R5329 M.n383 M.n382 0.00131395
R5330 M.n480 M.n465 0.00130925
R5331 M.n646 M.n639 0.00130925
R5332 M.n1907 M.n1906 0.00130268
R5333 M.n1249 M.n1248 0.00128603
R5334 M.n1231 M.n1230 0.00128603
R5335 M.n1479 M.n1478 0.00128488
R5336 M.n831 M.n830 0.00128488
R5337 M.n269 M.n268 0.00128488
R5338 M.n339 M.n338 0.00128488
R5339 M.n212 M.n211 0.00128488
R5340 M.n214 M.n213 0.00128488
R5341 M.n108 M.n107 0.00128488
R5342 M.n153 M.n152 0.00128488
R5343 M.n158 M.n157 0.00128488
R5344 M.n122 M.n121 0.00125362
R5345 M.n1543 M.n1542 0.00125251
R5346 M.n465 M.n464 0.00125145
R5347 M.n498 M.n483 0.00125145
R5348 M.n501 M.n500 0.00125145
R5349 M.n677 M.n676 0.00125145
R5350 M.n1917 M.n1907 0.00123579
R5351 M.n836 M.n835 0.00119767
R5352 M.n110 M.n97 0.00119565
R5353 M.n464 M.n463 0.00119364
R5354 M.n483 M.n480 0.00119364
R5355 M.n500 M.n499 0.00119364
R5356 M.n1905 M.n1904 0.0011689
R5357 M.n1303 M.n1302 0.00115502
R5358 M.n1272 M.n1271 0.00115502
R5359 M.n1481 M.n1479 0.00115407
R5360 M.n1410 M.n1409 0.00115407
R5361 M.n1414 M.n1413 0.00115407
R5362 M.n725 M.n724 0.00115407
R5363 M.n630 M.n629 0.00115407
R5364 M.n515 M.n514 0.00115407
R5365 M.n271 M.n270 0.00115407
R5366 M.n287 M.n286 0.00115407
R5367 M.n275 M.n274 0.00115407
R5368 M.n335 M.n334 0.00115407
R5369 M.n324 M.n323 0.00115407
R5370 M.n307 M.n306 0.00115407
R5371 M.n207 M.n206 0.00115407
R5372 M.n79 M.n78 0.00115407
R5373 M.n138 M.n137 0.00115407
R5374 M.n393 M.n392 0.00113953
R5375 M.n397 M.n396 0.00113953
R5376 M.n835 M.n834 0.00113953
R5377 M.n82 M.n81 0.00113768
R5378 M.n637 M.n636 0.00113584
R5379 M.n1194 M.n1193 0.00112857
R5380 M.n954 M.n953 0.00112069
R5381 M.n951 M.n950 0.00112069
R5382 M.n947 M.n946 0.00112069
R5383 M.n1008 M.n1006 0.00112069
R5384 M.n1088 M.n1087 0.00110759
R5385 M.n1835 M.n1834 0.00110201
R5386 M.n1841 M.n1839 0.00110201
R5387 M.n1844 M.n1843 0.00110201
R5388 M.n1743 M.n1742 0.00110201
R5389 M.n1644 M.n1643 0.00110201
R5390 M.n1527 M.n1506 0.00110201
R5391 M.n1451 M.n1450 0.0010814
R5392 M.n1427 M.n1426 0.0010814
R5393 M.n395 M.n394 0.0010814
R5394 M.n848 M.n837 0.0010814
R5395 M.n1733 M.n1732 0.00107971
R5396 M.n625 M.n612 0.00107803
R5397 M.n1197 M.n1196 0.00107143
R5398 M.n1087 M.n1086 0.00105696
R5399 M.n1306 M.n1305 0.00102402
R5400 M.n1300 M.n1299 0.00102402
R5401 M.n1297 M.n1296 0.00102402
R5402 M.n1292 M.n1291 0.00102402
R5403 M.n1276 M.n1275 0.00102402
R5404 M.n1261 M.n1260 0.00102402
R5405 M.n1204 M.n1203 0.00102402
R5406 M.n1219 M.n1218 0.00102402
R5407 M.n1338 M.n1337 0.00102326
R5408 M.n1483 M.n1482 0.00102326
R5409 M.n1333 M.n1332 0.00102326
R5410 M.n1336 M.n1335 0.00102326
R5411 M.n1342 M.n1341 0.00102326
R5412 M.n1424 M.n1423 0.00102326
R5413 M.n1463 M.n1462 0.00102326
R5414 M.n1402 M.n1394 0.00102326
R5415 M.n920 M.n919 0.00102326
R5416 M.n926 M.n924 0.00102326
R5417 M.n929 M.n928 0.00102326
R5418 M.n584 M.n583 0.00102326
R5419 M.n751 M.n750 0.00102326
R5420 M.n623 M.n622 0.00102326
R5421 M.n721 M.n720 0.00102326
R5422 M.n633 M.n632 0.00102326
R5423 M.n533 M.n528 0.00102326
R5424 M.n288 M.n287 0.00102326
R5425 M.n278 M.n277 0.00102326
R5426 M.n309 M.n308 0.00102326
R5427 M.n198 M.n197 0.00102326
R5428 M.n196 M.n195 0.00102326
R5429 M.n228 M.n227 0.00102326
R5430 M.n230 M.n229 0.00102326
R5431 M.n232 M.n231 0.00102326
R5432 M.n71 M.n70 0.00102326
R5433 M.n146 M.n145 0.00102326
R5434 M.n134 M.n133 0.00102174
R5435 M.n161 M.n150 0.00102174
R5436 M.n163 M.n162 0.00102174
R5437 M.n1090 M.n1089 0.00100633
R5438 M.n1582 M.n1581 0.00100314
R5439 M.n979 M.n978 0.000965517
R5440 M.n977 M.n976 0.000965517
R5441 M.n984 M.n983 0.000965517
R5442 M.n982 M.n981 0.000965517
R5443 M.n1058 M.n1057 0.000965517
R5444 M.n1056 M.n1055 0.000965517
R5445 M.n1048 M.n1047 0.000965517
R5446 M.n1046 M.n1045 0.000965517
R5447 M.n1044 M.n1043 0.000965517
R5448 M.n991 M.n990 0.000965517
R5449 M.n990 M.n989 0.000965517
R5450 M.n988 M.n987 0.000965517
R5451 M.n1026 M.n1025 0.000965517
R5452 M.n1024 M.n1023 0.000965517
R5453 M.n1022 M.n1021 0.000965517
R5454 M.n1020 M.n1019 0.000965517
R5455 M.n1004 M.n1003 0.000965517
R5456 M.n1002 M.n1001 0.000965517
R5457 M.n1000 M.n999 0.000965517
R5458 M.n1106 M.n1105 0.000965517
R5459 M.n1069 M.n1068 0.000965517
R5460 M.n1067 M.n1066 0.000965517
R5461 M.n1064 M.n1063 0.000965517
R5462 M.n1062 M.n1061 0.000965517
R5463 M.n1054 M.n1053 0.000965517
R5464 M.n1052 M.n1051 0.000965517
R5465 M.n1042 M.n1041 0.000965517
R5466 M.n1040 M.n1039 0.000965517
R5467 M.n1038 M.n1037 0.000965517
R5468 M.n1034 M.n1033 0.000965517
R5469 M.n1032 M.n1031 0.000965517
R5470 M.n1030 M.n1029 0.000965517
R5471 M.n1018 M.n1017 0.000965517
R5472 M.n1016 M.n1015 0.000965517
R5473 M.n1014 M.n1013 0.000965517
R5474 M.n1012 M.n1011 0.000965517
R5475 M.n998 M.n997 0.000965517
R5476 M.n996 M.n995 0.000965517
R5477 M.n994 M.n993 0.000965517
R5478 M.n1104 M.n1103 0.000965517
R5479 M.n121 M.n111 0.000963768
R5480 M.n688 M.n687 0.000962428
R5481 M.n1999 M.n1998 0.000951505
R5482 M.n1962 M.n1961 0.000951505
R5483 M.n1965 M.n1964 0.000951505
R5484 M.n1945 M.n1944 0.000951505
R5485 M.n1935 M.n1934 0.000951505
R5486 M.n1937 M.n1936 0.000951505
R5487 M.n1922 M.n1921 0.000951505
R5488 M.n1924 M.n1923 0.000951505
R5489 M.n1914 M.n1913 0.000951505
R5490 M.n1913 M.n1912 0.000951505
R5491 M.n1899 M.n1898 0.000951505
R5492 M.n1901 M.n1900 0.000951505
R5493 M.n1881 M.n1880 0.000951505
R5494 M.n1883 M.n1882 0.000951505
R5495 M.n1885 M.n1884 0.000951505
R5496 M.n1861 M.n1860 0.000951505
R5497 M.n1859 M.n1858 0.000951505
R5498 M.n1857 M.n1856 0.000951505
R5499 M.n1832 M.n1831 0.000951505
R5500 M.n2002 M.n2001 0.000951505
R5501 M.n1956 M.n1955 0.000951505
R5502 M.n1960 M.n1959 0.000951505
R5503 M.n1958 M.n1957 0.000951505
R5504 M.n1950 M.n1949 0.000951505
R5505 M.n1948 M.n1947 0.000951505
R5506 M.n1933 M.n1932 0.000951505
R5507 M.n1920 M.n1919 0.000951505
R5508 M.n1911 M.n1910 0.000951505
R5509 M.n1909 M.n1908 0.000951505
R5510 M.n1895 M.n1894 0.000951505
R5511 M.n1897 M.n1896 0.000951505
R5512 M.n1875 M.n1874 0.000951505
R5513 M.n1877 M.n1876 0.000951505
R5514 M.n1879 M.n1878 0.000951505
R5515 M.n1868 M.n1867 0.000951505
R5516 M.n1866 M.n1865 0.000951505
R5517 M.n1864 M.n1863 0.000951505
R5518 M.n1830 M.n1829 0.000951505
R5519 M.n1821 M.n1820 0.000951505
R5520 M.n1796 M.n1795 0.000951505
R5521 M.n1799 M.n1798 0.000951505
R5522 M.n1785 M.n1784 0.000951505
R5523 M.n1783 M.n1782 0.000951505
R5524 M.n1767 M.n1766 0.000951505
R5525 M.n1751 M.n1750 0.000951505
R5526 M.n1760 M.n1752 0.000951505
R5527 M.n1739 M.n1738 0.000951505
R5528 M.n1730 M.n1729 0.000951505
R5529 M.n1728 M.n1727 0.000951505
R5530 M.n1144 M.n1143 0.000951505
R5531 M.n1689 M.n1688 0.000951505
R5532 M.n1672 M.n1671 0.000951505
R5533 M.n1824 M.n1823 0.000951505
R5534 M.n1792 M.n1791 0.000951505
R5535 M.n1794 M.n1793 0.000951505
R5536 M.n1776 M.n1775 0.000951505
R5537 M.n1780 M.n1779 0.000951505
R5538 M.n1778 M.n1777 0.000951505
R5539 M.n1770 M.n1769 0.000951505
R5540 M.n1747 M.n1746 0.000951505
R5541 M.n1749 M.n1748 0.000951505
R5542 M.n1761 M.n1749 0.000951505
R5543 M.n1736 M.n1735 0.000951505
R5544 M.n1742 M.n1741 0.000951505
R5545 M.n1731 M.n1711 0.000951505
R5546 M.n1711 M.n1710 0.000951505
R5547 M.n1709 M.n1708 0.000951505
R5548 M.n1138 M.n1137 0.000951505
R5549 M.n1696 M.n1695 0.000951505
R5550 M.n1670 M.n1669 0.000951505
R5551 M.n1661 M.n1660 0.000951505
R5552 M.n1630 M.n1629 0.000951505
R5553 M.n1632 M.n1631 0.000951505
R5554 M.n1616 M.n1615 0.000951505
R5555 M.n1618 M.n1617 0.000951505
R5556 M.n1603 M.n1602 0.000951505
R5557 M.n1601 M.n1600 0.000951505
R5558 M.n1587 M.n1586 0.000951505
R5559 M.n1591 M.n1590 0.000951505
R5560 M.n1567 M.n1566 0.000951505
R5561 M.n1565 M.n1564 0.000951505
R5562 M.n1550 M.n1549 0.000951505
R5563 M.n1552 M.n1551 0.000951505
R5564 M.n1536 M.n1535 0.000951505
R5565 M.n1534 M.n1533 0.000951505
R5566 M.n1664 M.n1663 0.000951505
R5567 M.n1626 M.n1625 0.000951505
R5568 M.n1628 M.n1627 0.000951505
R5569 M.n1612 M.n1611 0.000951505
R5570 M.n1614 M.n1613 0.000951505
R5571 M.n1608 M.n1607 0.000951505
R5572 M.n1606 M.n1605 0.000951505
R5573 M.n1585 M.n1584 0.000951505
R5574 M.n1594 M.n1593 0.000951505
R5575 M.n1573 M.n1572 0.000951505
R5576 M.n1575 M.n1574 0.000951505
R5577 M.n1563 M.n1562 0.000951505
R5578 M.n1561 M.n1560 0.000951505
R5579 M.n1546 M.n1545 0.000951505
R5580 M.n1548 M.n1547 0.000951505
R5581 M.n1542 M.n1541 0.000951505
R5582 M.n1540 M.n1539 0.000951505
R5583 M.n1744 M.n1734 0.000950886
R5584 M.n650 M.n649 0.000904624
R5585 M.n1198 M.n1197 0.0009
R5586 M.n1246 M.n1245 0.000893013
R5587 M.n1248 M.n1247 0.000893013
R5588 M.n1251 M.n1250 0.000893013
R5589 M.n1253 M.n1252 0.000893013
R5590 M.n1284 M.n1283 0.000893013
R5591 M.n1282 M.n1281 0.000893013
R5592 M.n1280 M.n1279 0.000893013
R5593 M.n1277 M.n1276 0.000893013
R5594 M.n1274 M.n1273 0.000893013
R5595 M.n1271 M.n1270 0.000893013
R5596 M.n1269 M.n1268 0.000893013
R5597 M.n1267 M.n1266 0.000893013
R5598 M.n1265 M.n1264 0.000893013
R5599 M.n1263 M.n1262 0.000893013
R5600 M.n1258 M.n1257 0.000893013
R5601 M.n1256 M.n1255 0.000893013
R5602 M.n1205 M.n1204 0.000893013
R5603 M.n1207 M.n1206 0.000893013
R5604 M.n1208 M.n1207 0.000893013
R5605 M.n1210 M.n1209 0.000893013
R5606 M.n1212 M.n1211 0.000893013
R5607 M.n1242 M.n1241 0.000893013
R5608 M.n1240 M.n1239 0.000893013
R5609 M.n1238 M.n1237 0.000893013
R5610 M.n1235 M.n1234 0.000893013
R5611 M.n1232 M.n1231 0.000893013
R5612 M.n1229 M.n1228 0.000893013
R5613 M.n1227 M.n1226 0.000893013
R5614 M.n1225 M.n1224 0.000893013
R5615 M.n1223 M.n1222 0.000893013
R5616 M.n1221 M.n1220 0.000893013
R5617 M.n1216 M.n1215 0.000893013
R5618 M.n1498 M.n1497 0.000892442
R5619 M.n1455 M.n1454 0.000892442
R5620 M.n1442 M.n1441 0.000892442
R5621 M.n1440 M.n1439 0.000892442
R5622 M.n1433 M.n1432 0.000892442
R5623 M.n1421 M.n1420 0.000892442
R5624 M.n1423 M.n1422 0.000892442
R5625 M.n1409 M.n1408 0.000892442
R5626 M.n1408 M.n1407 0.000892442
R5627 M.n1396 M.n1395 0.000892442
R5628 M.n1398 M.n1397 0.000892442
R5629 M.n1380 M.n1379 0.000892442
R5630 M.n1382 M.n1381 0.000892442
R5631 M.n1384 M.n1383 0.000892442
R5632 M.n1366 M.n1365 0.000892442
R5633 M.n1364 M.n1363 0.000892442
R5634 M.n1362 M.n1361 0.000892442
R5635 M.n1331 M.n1330 0.000892442
R5636 M.n1501 M.n1500 0.000892442
R5637 M.n1453 M.n1452 0.000892442
R5638 M.n1464 M.n1463 0.000892442
R5639 M.n1462 M.n1461 0.000892442
R5640 M.n1447 M.n1446 0.000892442
R5641 M.n1445 M.n1444 0.000892442
R5642 M.n1431 M.n1430 0.000892442
R5643 M.n1417 M.n1416 0.000892442
R5644 M.n1419 M.n1418 0.000892442
R5645 M.n1413 M.n1412 0.000892442
R5646 M.n1412 M.n1411 0.000892442
R5647 M.n1394 M.n1393 0.000892442
R5648 M.n1401 M.n1400 0.000892442
R5649 M.n1374 M.n1373 0.000892442
R5650 M.n1376 M.n1375 0.000892442
R5651 M.n1378 M.n1377 0.000892442
R5652 M.n1360 M.n1359 0.000892442
R5653 M.n1358 M.n1357 0.000892442
R5654 M.n1356 M.n1355 0.000892442
R5655 M.n1329 M.n1328 0.000892442
R5656 M.n777 M.n776 0.000892442
R5657 M.n788 M.n787 0.000892442
R5658 M.n790 M.n789 0.000892442
R5659 M.n801 M.n800 0.000892442
R5660 M.n803 M.n802 0.000892442
R5661 M.n817 M.n816 0.000892442
R5662 M.n819 M.n818 0.000892442
R5663 M.n821 M.n820 0.000892442
R5664 M.n827 M.n826 0.000892442
R5665 M.n826 M.n825 0.000892442
R5666 M.n843 M.n842 0.000892442
R5667 M.n845 M.n844 0.000892442
R5668 M.n861 M.n860 0.000892442
R5669 M.n863 M.n862 0.000892442
R5670 M.n865 M.n864 0.000892442
R5671 M.n883 M.n882 0.000892442
R5672 M.n881 M.n880 0.000892442
R5673 M.n879 M.n878 0.000892442
R5674 M.n894 M.n893 0.000892442
R5675 M.n775 M.n774 0.000892442
R5676 M.n784 M.n783 0.000892442
R5677 M.n786 M.n785 0.000892442
R5678 M.n797 M.n796 0.000892442
R5679 M.n799 M.n798 0.000892442
R5680 M.n811 M.n810 0.000892442
R5681 M.n813 M.n812 0.000892442
R5682 M.n815 M.n814 0.000892442
R5683 M.n832 M.n831 0.000892442
R5684 M.n830 M.n829 0.000892442
R5685 M.n839 M.n838 0.000892442
R5686 M.n841 M.n840 0.000892442
R5687 M.n855 M.n854 0.000892442
R5688 M.n857 M.n856 0.000892442
R5689 M.n859 M.n858 0.000892442
R5690 M.n877 M.n876 0.000892442
R5691 M.n875 M.n874 0.000892442
R5692 M.n873 M.n872 0.000892442
R5693 M.n892 M.n891 0.000892442
R5694 M.n603 M.n602 0.000892442
R5695 M.n605 M.n604 0.000892442
R5696 M.n620 M.n619 0.000892442
R5697 M.n622 M.n621 0.000892442
R5698 M.n629 M.n628 0.000892442
R5699 M.n627 M.n626 0.000892442
R5700 M.n643 M.n642 0.000892442
R5701 M.n658 M.n657 0.000892442
R5702 M.n660 M.n659 0.000892442
R5703 M.n683 M.n682 0.000892442
R5704 M.n694 M.n693 0.000892442
R5705 M.n696 M.n695 0.000892442
R5706 M.n707 M.n706 0.000892442
R5707 M.n709 M.n708 0.000892442
R5708 M.n720 M.n719 0.000892442
R5709 M.n722 M.n721 0.000892442
R5710 M.n598 M.n597 0.000892442
R5711 M.n600 M.n599 0.000892442
R5712 M.n615 M.n614 0.000892442
R5713 M.n617 M.n616 0.000892442
R5714 M.n634 M.n633 0.000892442
R5715 M.n632 M.n631 0.000892442
R5716 M.n641 M.n640 0.000892442
R5717 M.n652 M.n651 0.000892442
R5718 M.n654 M.n653 0.000892442
R5719 M.n656 M.n655 0.000892442
R5720 M.n669 M.n668 0.000892442
R5721 M.n667 M.n666 0.000892442
R5722 M.n680 M.n679 0.000892442
R5723 M.n690 M.n689 0.000892442
R5724 M.n692 M.n691 0.000892442
R5725 M.n716 M.n715 0.000892442
R5726 M.n718 M.n717 0.000892442
R5727 M.n454 M.n453 0.000892442
R5728 M.n456 M.n455 0.000892442
R5729 M.n458 M.n457 0.000892442
R5730 M.n473 M.n472 0.000892442
R5731 M.n475 M.n474 0.000892442
R5732 M.n477 M.n476 0.000892442
R5733 M.n495 M.n494 0.000892442
R5734 M.n493 M.n492 0.000892442
R5735 M.n491 M.n490 0.000892442
R5736 M.n510 M.n509 0.000892442
R5737 M.n512 M.n511 0.000892442
R5738 M.n514 M.n513 0.000892442
R5739 M.n528 M.n527 0.000892442
R5740 M.n532 M.n531 0.000892442
R5741 M.n530 M.n529 0.000892442
R5742 M.n546 M.n545 0.000892442
R5743 M.n560 M.n559 0.000892442
R5744 M.n562 M.n561 0.000892442
R5745 M.n452 M.n451 0.000892442
R5746 M.n467 M.n466 0.000892442
R5747 M.n469 M.n468 0.000892442
R5748 M.n471 M.n470 0.000892442
R5749 M.n489 M.n488 0.000892442
R5750 M.n487 M.n486 0.000892442
R5751 M.n485 M.n484 0.000892442
R5752 M.n506 M.n505 0.000892442
R5753 M.n508 M.n507 0.000892442
R5754 M.n517 M.n516 0.000892442
R5755 M.n526 M.n525 0.000892442
R5756 M.n537 M.n536 0.000892442
R5757 M.n535 M.n534 0.000892442
R5758 M.n544 M.n543 0.000892442
R5759 M.n554 M.n553 0.000892442
R5760 M.n556 M.n555 0.000892442
R5761 M.n558 M.n557 0.000892442
R5762 M.n574 M.n573 0.000892442
R5763 M.n285 M.n284 0.000892442
R5764 M.n259 M.n258 0.000892442
R5765 M.n260 M.n259 0.000892442
R5766 M.n262 M.n261 0.000892442
R5767 M.n265 M.n264 0.000892442
R5768 M.n267 M.n266 0.000892442
R5769 M.n338 M.n337 0.000892442
R5770 M.n336 M.n335 0.000892442
R5771 M.n333 M.n332 0.000892442
R5772 M.n331 M.n330 0.000892442
R5773 M.n329 M.n328 0.000892442
R5774 M.n325 M.n324 0.000892442
R5775 M.n323 M.n322 0.000892442
R5776 M.n321 M.n320 0.000892442
R5777 M.n319 M.n318 0.000892442
R5778 M.n317 M.n316 0.000892442
R5779 M.n314 M.n313 0.000892442
R5780 M.n312 M.n311 0.000892442
R5781 M.n310 M.n309 0.000892442
R5782 M.n306 M.n305 0.000892442
R5783 M.n249 M.n248 0.000892442
R5784 M.n254 M.n253 0.000892442
R5785 M.n256 M.n255 0.000892442
R5786 M.n375 M.n374 0.000892442
R5787 M.n374 M.n373 0.000892442
R5788 M.n372 M.n371 0.000892442
R5789 M.n369 M.n368 0.000892442
R5790 M.n367 M.n366 0.000892442
R5791 M.n365 M.n364 0.000892442
R5792 M.n359 M.n358 0.000892442
R5793 M.n357 M.n356 0.000892442
R5794 M.n355 M.n354 0.000892442
R5795 M.n353 M.n352 0.000892442
R5796 M.n350 M.n349 0.000892442
R5797 M.n348 M.n347 0.000892442
R5798 M.n346 M.n345 0.000892442
R5799 M.n342 M.n341 0.000892442
R5800 M.n70 M.n69 0.000892442
R5801 M.n78 M.n77 0.000892442
R5802 M.n91 M.n90 0.000892442
R5803 M.n104 M.n103 0.000892442
R5804 M.n105 M.n104 0.000892442
R5805 M.n107 M.n106 0.000892442
R5806 M.n115 M.n114 0.000892442
R5807 M.n113 M.n112 0.000892442
R5808 M.n129 M.n128 0.000892442
R5809 M.n147 M.n146 0.000892442
R5810 M.n154 M.n153 0.000892442
R5811 M.n152 M.n151 0.000892442
R5812 M.n171 M.n170 0.000892442
R5813 M.n173 M.n172 0.000892442
R5814 M.n184 M.n183 0.000892442
R5815 M.n182 M.n181 0.000892442
R5816 M.n194 M.n193 0.000892442
R5817 M.n75 M.n74 0.000892442
R5818 M.n86 M.n85 0.000892442
R5819 M.n88 M.n87 0.000892442
R5820 M.n99 M.n98 0.000892442
R5821 M.n100 M.n99 0.000892442
R5822 M.n102 M.n101 0.000892442
R5823 M.n119 M.n118 0.000892442
R5824 M.n127 M.n126 0.000892442
R5825 M.n137 M.n136 0.000892442
R5826 M.n159 M.n158 0.000892442
R5827 M.n157 M.n156 0.000892442
R5828 M.n167 M.n166 0.000892442
R5829 M.n169 M.n168 0.000892442
R5830 M.n180 M.n179 0.000892442
R5831 M.n178 M.n177 0.000892442
R5832 M.n192 M.n191 0.000892442
R5833 M.n1763 M.n1762 0.000886473
R5834 M.n1732 M.n1707 0.000886473
R5835 M.n1406 M.n1405 0.000848837
R5836 M.n96 M.n95 0.000847826
R5837 M.n1195 M.n1194 0.000842857
R5838 M.n1904 M.n1893 0.000834448
R5839 M.n1745 M.n1744 0.000822061
R5840 M.n1544 M.n1531 0.000814465
R5841 M.n1715 M.n1714 0.000801003
R5842 M.n1723 M.n1722 0.000801003
R5843 M.n1720 M.n1719 0.000801003
R5844 M.n1717 M.n1716 0.000801003
R5845 M.n1740 M.n1737 0.000801003
R5846 M.n1146 M.n1145 0.000801003
R5847 M.n1148 M.n1147 0.000801003
R5848 M.n1687 M.n1686 0.000801003
R5849 M.n1685 M.n1684 0.000801003
R5850 M.n1743 M.n1736 0.000801003
R5851 M.n1140 M.n1139 0.000801003
R5852 M.n1142 M.n1141 0.000801003
R5853 M.n1694 M.n1693 0.000801003
R5854 M.n1692 M.n1691 0.000801003
R5855 M.n1574 M.n1573 0.000801003
R5856 M.n1415 M.n1406 0.000790698
R5857 M.n577 M.n576 0.000789017
R5858 M.n676 M.n675 0.000789017
R5859 M.n1890 M.n1889 0.000767559
R5860 M.n1873 M.n1870 0.000767559
R5861 M.n1854 M.n1853 0.000767559
R5862 M.n1491 M.n1490 0.000761628
R5863 M.n1458 M.n1457 0.000761628
R5864 M.n734 M.n733 0.000761628
R5865 M.n663 M.n662 0.000761628
R5866 M.n673 M.n672 0.000761628
R5867 M.n708 M.n707 0.000761628
R5868 M.n674 M.n669 0.000761628
R5869 M.n704 M.n703 0.000761628
R5870 M.n413 M.n412 0.000761628
R5871 M.n455 M.n454 0.000761628
R5872 M.n565 M.n564 0.000761628
R5873 M.n571 M.n570 0.000761628
R5874 M.n449 M.n448 0.000761628
R5875 M.n518 M.n517 0.000761628
R5876 M.n555 M.n554 0.000761628
R5877 M.n575 M.n574 0.000761628
R5878 M.n263 M.n262 0.000761628
R5879 M.n251 M.n250 0.000761628
R5880 M.n371 M.n370 0.000761628
R5881 M.n362 M.n361 0.000761628
R5882 M.n143 M.n142 0.000761628
R5883 M.n145 M.n144 0.000761628
R5884 M.n140 M.n139 0.000761628
R5885 M.n1529 M.n1528 0.000751572
R5886 M.n1404 M.n1403 0.000732558
R5887 M.n1390 M.n1389 0.000732558
R5888 M.n1387 M.n1372 0.000732558
R5889 M.n1354 M.n1353 0.000732558
R5890 M.n853 M.n852 0.000732558
R5891 M.n886 M.n871 0.000732558
R5892 M.n889 M.n888 0.000732558
R5893 M.n165 M.n164 0.000731884
R5894 M.n187 M.n176 0.000731884
R5895 M.n189 M.n188 0.000731884
R5896 M.n446 M.n445 0.000731214
R5897 M.n567 M.n552 0.000731214
R5898 M.n638 M.n637 0.000731214
R5899 M.n665 M.n650 0.000731214
R5900 M.n701 M.n700 0.000731214
R5901 M.n1325 M.n1324 0.000728571
R5902 M.n1190 M.n1189 0.000728571
R5903 M.n1187 M.n1186 0.000728571
R5904 M.n1095 M.n1094 0.000702532
R5905 M.n1098 M.n1097 0.000702532
R5906 M.n1101 M.n1100 0.000702532
R5907 M.n377 M.n376 0.000674419
R5908 M.n388 M.n387 0.000674419
R5909 M.n1323 M.n1322 0.000671429
R5910 M.n1192 M.n1191 0.000671429
R5911 M.n1021 M.n1020 0.000655172
R5912 M.n1001 M.n1000 0.000655172
R5913 M.n1013 M.n1012 0.000655172
R5914 M.n995 M.n994 0.000655172
R5915 M.n1884 M.n1883 0.000650502
R5916 M.n1858 M.n1857 0.000650502
R5917 M.n1878 M.n1877 0.000650502
R5918 M.n1865 M.n1864 0.000650502
R5919 M.n1756 M.n1755 0.000650502
R5920 M.n1740 M.n1739 0.000650502
R5921 M.n1147 M.n1146 0.000650502
R5922 M.n1686 M.n1685 0.000650502
R5923 M.n1141 M.n1140 0.000650502
R5924 M.n1693 M.n1692 0.000650502
R5925 M.n1589 M.n1588 0.000650502
R5926 M.n1577 M.n1576 0.000650502
R5927 M.n1266 M.n1265 0.000631004
R5928 M.n1257 M.n1256 0.000631004
R5929 M.n1224 M.n1223 0.000631004
R5930 M.n1215 M.n1214 0.000631004
R5931 M.n1459 M.n1458 0.000630814
R5932 M.n1457 M.n1456 0.000630814
R5933 M.n1381 M.n1380 0.000630814
R5934 M.n1365 M.n1364 0.000630814
R5935 M.n1375 M.n1374 0.000630814
R5936 M.n1359 M.n1358 0.000630814
R5937 M.n864 M.n863 0.000630814
R5938 M.n880 M.n879 0.000630814
R5939 M.n858 M.n857 0.000630814
R5940 M.n874 M.n873 0.000630814
R5941 M.n737 M.n735 0.000630814
R5942 M.n663 M.n661 0.000630814
R5943 M.n673 M.n670 0.000630814
R5944 M.n664 M.n656 0.000630814
R5945 M.n703 M.n702 0.000630814
R5946 M.n705 M.n704 0.000630814
R5947 M.n411 M.n410 0.000630814
R5948 M.n565 M.n563 0.000630814
R5949 M.n571 M.n568 0.000630814
R5950 M.n448 M.n447 0.000630814
R5951 M.n450 M.n449 0.000630814
R5952 M.n538 M.n526 0.000630814
R5953 M.n566 M.n558 0.000630814
R5954 M.n326 M.n325 0.000630814
R5955 M.n252 M.n251 0.000630814
R5956 M.n361 M.n360 0.000630814
R5957 M.n221 M.n220 0.000630814
R5958 M.n144 M.n143 0.000630814
R5959 M.n172 M.n171 0.000630814
R5960 M.n183 M.n182 0.000630814
R5961 M.n139 M.n138 0.000630814
R5962 M.n141 M.n140 0.000630814
R5963 M.n168 M.n167 0.000630814
R5964 M.n179 M.n178 0.000630814
R5965 M.n1704 M.n1703 0.000628824
R5966 M.n1701 M.n1698 0.000628824
R5967 M.n1682 M.n1681 0.000628824
R5968 M.n1571 M.n1570 0.000625786
R5969 M.n379 M.n378 0.000616279
R5970 M.n385 M.n384 0.000616279
R5971 M.n135 M.n134 0.000615942
R5972 M.n520 M.n519 0.000615607
R5973 M.n551 M.n550 0.000615607
R5974 M.n244 M.n243 0.00055814
R5975 M.n851 M.n850 0.00055814
R5976 M.n504 M.n503 0.000557804
R5977 M.n539 M.n524 0.000557804
R5978 M.n1092 M.n1091 0.000550633
C0 m1_n36350_7190# P 0.782f
C1 P M 0.696p
C2 m1_n36350_7190# M 0.0433f
C3 M VSUBS 0.256p
C4 P VSUBS 1.08p
C5 m1_n36350_7190# VSUBS 3.7f $ **FLOATING
C6 M.t74 VSUBS 4.09f
C7 M.t110 VSUBS 3.72f
C8 M.n0 VSUBS 1.84f
C9 M.t112 VSUBS 3.72f
C10 M.n1 VSUBS 1.11f
C11 M.t56 VSUBS 3.72f
C12 M.n2 VSUBS 1.11f
C13 M.t70 VSUBS 3.72f
C14 M.n3 VSUBS 1.11f
C15 M.t37 VSUBS 3.72f
C16 M.n4 VSUBS 1.11f
C17 M.t126 VSUBS 3.72f
C18 M.n5 VSUBS 1.11f
C19 M.t100 VSUBS 3.72f
C20 M.n6 VSUBS 1.11f
C21 M.t36 VSUBS 3.72f
C22 M.n7 VSUBS 1.11f
C23 M.t48 VSUBS 3.72f
C24 M.n8 VSUBS 1.11f
C25 M.t26 VSUBS 3.72f
C26 M.n9 VSUBS 1.11f
C27 M.t107 VSUBS 3.72f
C28 M.n10 VSUBS 0.845f
C29 M.t61 VSUBS 4.09f
C30 M.t129 VSUBS 3.72f
C31 M.n11 VSUBS 1.84f
C32 M.t50 VSUBS 3.72f
C33 M.n12 VSUBS 1.11f
C34 M.t6 VSUBS 3.72f
C35 M.n13 VSUBS 1.11f
C36 M.t11 VSUBS 3.72f
C37 M.n14 VSUBS 1.11f
C38 M.t123 VSUBS 3.72f
C39 M.n15 VSUBS 1.11f
C40 M.t72 VSUBS 3.72f
C41 M.n16 VSUBS 1.11f
C42 M.t38 VSUBS 3.72f
C43 M.n17 VSUBS 1.11f
C44 M.t121 VSUBS 3.72f
C45 M.n18 VSUBS 1.11f
C46 M.t131 VSUBS 3.72f
C47 M.n19 VSUBS 1.11f
C48 M.t103 VSUBS 3.72f
C49 M.n20 VSUBS 1.11f
C50 M.t49 VSUBS 3.72f
C51 M.n21 VSUBS 0.851f
C52 M.t108 VSUBS 4.09f
C53 M.t77 VSUBS 3.72f
C54 M.n22 VSUBS 1.84f
C55 M.t106 VSUBS 3.72f
C56 M.n23 VSUBS 1.11f
C57 M.t52 VSUBS 3.72f
C58 M.n24 VSUBS 1.11f
C59 M.t66 VSUBS 3.72f
C60 M.n25 VSUBS 1.11f
C61 M.t35 VSUBS 3.72f
C62 M.n26 VSUBS 1.11f
C63 M.t124 VSUBS 3.72f
C64 M.n27 VSUBS 1.11f
C65 M.t96 VSUBS 3.72f
C66 M.n28 VSUBS 1.11f
C67 M.t33 VSUBS 3.72f
C68 M.n29 VSUBS 1.11f
C69 M.t43 VSUBS 3.72f
C70 M.n30 VSUBS 1.11f
C71 M.t25 VSUBS 3.72f
C72 M.n31 VSUBS 1.11f
C73 M.t104 VSUBS 3.72f
C74 M.n32 VSUBS 0.85f
C75 M.t65 VSUBS 4.09f
C76 M.t32 VSUBS 3.72f
C77 M.n33 VSUBS 1.84f
C78 M.t21 VSUBS 3.72f
C79 M.n34 VSUBS 1.11f
C80 M.t98 VSUBS 3.72f
C81 M.n35 VSUBS 1.11f
C82 M.t109 VSUBS 3.72f
C83 M.n36 VSUBS 1.11f
C84 M.t89 VSUBS 3.72f
C85 M.n37 VSUBS 1.11f
C86 M.t30 VSUBS 3.72f
C87 M.n38 VSUBS 1.11f
C88 M.t13 VSUBS 3.72f
C89 M.n39 VSUBS 1.11f
C90 M.t87 VSUBS 3.72f
C91 M.n40 VSUBS 1.11f
C92 M.t93 VSUBS 3.72f
C93 M.n41 VSUBS 1.11f
C94 M.t76 VSUBS 3.72f
C95 M.n42 VSUBS 1.11f
C96 M.t19 VSUBS 3.72f
C97 M.n43 VSUBS 0.85f
C98 M.t20 VSUBS 4.09f
C99 M.t86 VSUBS 3.72f
C100 M.n44 VSUBS 1.84f
C101 M.t4 VSUBS 3.72f
C102 M.n45 VSUBS 1.11f
C103 M.t84 VSUBS 3.72f
C104 M.n46 VSUBS 1.11f
C105 M.t90 VSUBS 3.72f
C106 M.n47 VSUBS 1.11f
C107 M.t68 VSUBS 3.72f
C108 M.n48 VSUBS 1.11f
C109 M.t16 VSUBS 3.72f
C110 M.n49 VSUBS 1.11f
C111 M.t125 VSUBS 3.72f
C112 M.n50 VSUBS 1.11f
C113 M.t63 VSUBS 3.72f
C114 M.n51 VSUBS 1.11f
C115 M.t79 VSUBS 3.72f
C116 M.n52 VSUBS 1.11f
C117 M.t46 VSUBS 3.72f
C118 M.n53 VSUBS 1.11f
C119 M.t2 VSUBS 3.72f
C120 M.n54 VSUBS 0.851f
C121 M.t23 VSUBS 4.09f
C122 M.t73 VSUBS 3.72f
C123 M.n55 VSUBS 1.84f
C124 M.t120 VSUBS 3.72f
C125 M.n56 VSUBS 1.11f
C126 M.t62 VSUBS 3.72f
C127 M.n57 VSUBS 1.11f
C128 M.t78 VSUBS 3.72f
C129 M.n58 VSUBS 1.11f
C130 M.t45 VSUBS 3.72f
C131 M.n59 VSUBS 1.11f
C132 M.t0 VSUBS 3.72f
C133 M.n60 VSUBS 1.11f
C134 M.t105 VSUBS 3.72f
C135 M.n61 VSUBS 1.11f
C136 M.t42 VSUBS 3.72f
C137 M.n62 VSUBS 1.11f
C138 M.t55 VSUBS 3.72f
C139 M.n63 VSUBS 1.11f
C140 M.t31 VSUBS 3.72f
C141 M.n64 VSUBS 1.11f
C142 M.t117 VSUBS 3.72f
C143 M.n65 VSUBS 0.85f
C144 M.n66 VSUBS 0.0314f
C145 M.n67 VSUBS 0.0101f
C146 M.n68 VSUBS 0.0315f
C147 M.n69 VSUBS 0.00845f
C148 M.n70 VSUBS 0.00204f
C149 M.n71 VSUBS 0.00962f
C150 M.n72 VSUBS 0.0105f
C151 M.n73 VSUBS 0.0512f
C152 M.n74 VSUBS 0.00845f
C153 M.n75 VSUBS 0.00321f
C154 M.n76 VSUBS 0.00845f
C155 M.n77 VSUBS 0.00845f
C156 M.n78 VSUBS 0.00233f
C157 M.n79 VSUBS 0.00991f
C158 M.n80 VSUBS 0.0108f
C159 M.n81 VSUBS 0.0117f
C160 M.n82 VSUBS 0.0117f
C161 M.n83 VSUBS 0.0152f
C162 M.n84 VSUBS 0.0181f
C163 M.n85 VSUBS 0.00845f
C164 M.n86 VSUBS 0.00758f
C165 M.n87 VSUBS 0.00758f
C166 M.n88 VSUBS 0.0114f
C167 M.n89 VSUBS 0.00933f
C168 M.n90 VSUBS 0.00933f
C169 M.n91 VSUBS 0.0105f
C170 M.n92 VSUBS 0.0195f
C171 M.n93 VSUBS 0.0204f
C172 M.n94 VSUBS 0.0213f
C173 M.n95 VSUBS 0.0117f
C174 M.n96 VSUBS 0.00789f
C175 M.n97 VSUBS 0.00965f
C176 M.n98 VSUBS 0.0108f
C177 M.n99 VSUBS 0.00175f
C178 M.n100 VSUBS 0.00699f
C179 M.n101 VSUBS 0.00699f
C180 M.n102 VSUBS 0.0035f
C181 M.n103 VSUBS 0.0108f
C182 M.n104 VSUBS 0.00175f
C183 M.n105 VSUBS 0.00787f
C184 M.n106 VSUBS 0.00787f
C185 M.n107 VSUBS 0.00262f
C186 M.n108 VSUBS 0.00962f
C187 M.n109 VSUBS 0.0105f
C188 M.n110 VSUBS 0.00906f
C189 M.n111 VSUBS 0.466f
C190 M.n112 VSUBS 0.0119f
C191 M.n113 VSUBS 0.00787f
C192 M.n114 VSUBS 0.00787f
C193 M.n115 VSUBS 0.00291f
C194 M.n116 VSUBS 0.00991f
C195 M.n117 VSUBS 0.00787f
C196 M.n118 VSUBS 0.00787f
C197 M.n119 VSUBS 0.00379f
C198 M.n120 VSUBS 0.0108f
C199 M.n121 VSUBS 0.00614f
C200 M.n122 VSUBS 0.0117f
C201 M.n123 VSUBS 0.0172f
C202 M.n124 VSUBS 0.0208f
C203 M.n125 VSUBS 0.0102f
C204 M.n126 VSUBS 0.0102f
C205 M.n127 VSUBS 0.0114f
C206 M.n128 VSUBS 0.0119f
C207 M.n129 VSUBS 0.0105f
C208 M.n130 VSUBS 0.0189f
C209 M.n131 VSUBS 0.0189f
C210 M.n132 VSUBS 0.0199f
C211 M.n133 VSUBS 0.0111f
C212 M.n134 VSUBS 0.00322f
C213 M.n135 VSUBS 0.00877f
C214 M.n136 VSUBS 0.00933f
C215 M.n137 VSUBS 0.00233f
C216 M.n138 VSUBS 0.00175f
C217 M.n139 VSUBS 8.74e-19
C218 M.n140 VSUBS 8.74e-19
C219 M.n141 VSUBS 0.00816f
C220 M.n142 VSUBS 0.00991f
C221 M.n143 VSUBS 8.74e-19
C222 M.n144 VSUBS 8.74e-19
C223 M.n145 VSUBS 0.00175f
C224 M.n146 VSUBS 0.00204f
C225 M.n147 VSUBS 0.00787f
C226 M.n148 VSUBS 0.00962f
C227 M.n149 VSUBS 0.0105f
C228 M.n150 VSUBS 0.0108f
C229 M.n151 VSUBS 0.0306f
C230 M.n152 VSUBS 0.00262f
C231 M.n153 VSUBS 0.00262f
C232 M.n154 VSUBS 0.00816f
C233 M.n155 VSUBS 0.00991f
C234 M.n156 VSUBS 0.0289f
C235 M.n157 VSUBS 0.00262f
C236 M.n158 VSUBS 0.00262f
C237 M.n159 VSUBS 0.00904f
C238 M.n160 VSUBS 0.0108f
C239 M.n161 VSUBS 0.0117f
C240 M.n162 VSUBS 0.0117f
C241 M.n163 VSUBS 0.0307f
C242 M.n164 VSUBS 0.0292f
C243 M.n165 VSUBS 0.0114f
C244 M.n166 VSUBS 0.0289f
C245 M.n167 VSUBS 0.00117f
C246 M.n168 VSUBS 0.00117f
C247 M.n169 VSUBS 0.0102f
C248 M.n170 VSUBS 0.0306f
C249 M.n171 VSUBS 0.00117f
C250 M.n172 VSUBS 0.00117f
C251 M.n173 VSUBS 0.00933f
C252 M.n174 VSUBS 0.00962f
C253 M.n175 VSUBS 0.0105f
C254 M.n176 VSUBS 0.0114f
C255 M.n177 VSUBS 0.0385f
C256 M.n178 VSUBS 0.00117f
C257 M.n179 VSUBS 0.00117f
C258 M.n180 VSUBS 0.0105f
C259 M.n181 VSUBS 0.0402f
C260 M.n182 VSUBS 0.00117f
C261 M.n183 VSUBS 0.00117f
C262 M.n184 VSUBS 0.00962f
C263 M.n185 VSUBS 0.00991f
C264 M.n186 VSUBS 0.0108f
C265 M.n187 VSUBS 0.0117f
C266 M.n188 VSUBS 0.0117f
C267 M.n189 VSUBS 0.0389f
C268 M.n190 VSUBS 0.0491f
C269 M.n191 VSUBS 0.0385f
C270 M.n192 VSUBS 0.0114f
C271 M.n193 VSUBS 0.0402f
C272 M.n194 VSUBS 0.0105f
C273 M.n195 VSUBS 0.0419f
C274 M.n196 VSUBS 0.0097f
C275 M.n197 VSUBS 0.193f
C276 M.n198 VSUBS 0.0522f
C277 M.n199 VSUBS 0.0536f
C278 M.n200 VSUBS 0.0224f
C279 M.n201 VSUBS 0.0522f
C280 M.n202 VSUBS 0.0402f
C281 M.n203 VSUBS 0.0291f
C282 M.n204 VSUBS 0.14f
C283 M.n205 VSUBS 0.00105f
C284 M.n206 VSUBS 0.00991f
C285 M.n207 VSUBS 0.00991f
C286 M.n208 VSUBS 0.0187f
C287 M.n209 VSUBS 0.0198f
C288 M.n210 VSUBS 0.0195f
C289 M.n211 VSUBS 0.0117f
C290 M.n212 VSUBS 0.00962f
C291 M.n213 VSUBS 0.00962f
C292 M.n214 VSUBS 0.00962f
C293 M.n215 VSUBS 0.00991f
C294 M.n216 VSUBS 0.00991f
C295 M.n217 VSUBS 0.0207f
C296 M.n218 VSUBS 0.0224f
C297 M.n219 VSUBS 0.0195f
C298 M.n220 VSUBS 0.0102f
C299 M.n221 VSUBS 0.00291f
C300 M.n222 VSUBS 0.00962f
C301 M.n223 VSUBS 0.00962f
C302 M.n224 VSUBS 0.00991f
C303 M.n225 VSUBS 0.00991f
C304 M.n226 VSUBS 0.0341f
C305 M.n227 VSUBS 0.0326f
C306 M.n228 VSUBS 0.00962f
C307 M.n229 VSUBS 0.00962f
C308 M.n230 VSUBS 0.00991f
C309 M.n231 VSUBS 0.00991f
C310 M.n232 VSUBS 0.0423f
C311 M.n233 VSUBS 0.0507f
C312 M.n234 VSUBS 0.0834f
C313 M.n235 VSUBS 0.0623f
C314 M.n236 VSUBS 0.0195f
C315 M.n237 VSUBS 0.0616f
C316 M.n238 VSUBS 0.0213f
C317 M.n239 VSUBS 0.0231f
C318 M.n240 VSUBS 1.25f
C319 M.n241 VSUBS 1.25f
C320 M.n242 VSUBS 0.0227f
C321 M.n243 VSUBS 0.0117f
C322 M.n244 VSUBS 0.0117f
C323 M.n245 VSUBS 0.051f
C324 M.n246 VSUBS 0.051f
C325 M.n247 VSUBS 0.0572f
C326 M.n248 VSUBS 0.0114f
C327 M.n249 VSUBS 0.0108f
C328 M.n250 VSUBS 0.0105f
C329 M.n251 VSUBS 8.74e-19
C330 M.n252 VSUBS 0.0108f
C331 M.n253 VSUBS 0.0114f
C332 M.n254 VSUBS 0.0405f
C333 M.n255 VSUBS 0.0405f
C334 M.n256 VSUBS 0.0114f
C335 M.n257 VSUBS 0.058f
C336 M.n258 VSUBS 0.0105f
C337 M.n259 VSUBS 0.00175f
C338 M.n260 VSUBS 0.00904f
C339 M.n261 VSUBS 0.00904f
C340 M.n262 VSUBS 0.00146f
C341 M.n263 VSUBS 0.0105f
C342 M.n264 VSUBS 0.0108f
C343 M.n265 VSUBS 0.0423f
C344 M.n266 VSUBS 0.0423f
C345 M.n267 VSUBS 0.0105f
C346 M.n268 VSUBS 0.0695f
C347 M.n269 VSUBS 0.00991f
C348 M.n270 VSUBS 0.00962f
C349 M.n271 VSUBS 0.0114f
C350 M.n272 VSUBS 0.053f
C351 M.n273 VSUBS 0.0528f
C352 M.n274 VSUBS 0.062f
C353 M.n275 VSUBS 0.01f
C354 M.n276 VSUBS 0.0011f
C355 M.n277 VSUBS 0.00962f
C356 M.n278 VSUBS 0.00962f
C357 M.n279 VSUBS 0.0152f
C358 M.n280 VSUBS 0.0166f
C359 M.n281 VSUBS 0.0195f
C360 M.n282 VSUBS 0.0283f
C361 M.n283 VSUBS 0.0286f
C362 M.n284 VSUBS 0.0108f
C363 M.n285 VSUBS 0.00816f
C364 M.n286 VSUBS 0.00874f
C365 M.n287 VSUBS 0.00262f
C366 M.n288 VSUBS 0.00845f
C367 M.n289 VSUBS 0.00962f
C368 M.n290 VSUBS 0.00962f
C369 M.n291 VSUBS 0.0376f
C370 M.n292 VSUBS 0.0402f
C371 M.n293 VSUBS 0.0122f
C372 M.n294 VSUBS 0.00962f
C373 M.n295 VSUBS 0.00991f
C374 M.n296 VSUBS 0.153f
C375 M.n297 VSUBS 0.17f
C376 M.n298 VSUBS 0.049f
C377 M.n299 VSUBS 0.0181f
C378 M.n300 VSUBS 0.0571f
C379 M.n301 VSUBS 0.0621f
C380 M.n302 VSUBS 0.0749f
C381 M.n303 VSUBS 0.0122f
C382 M.n304 VSUBS 0.0513f
C383 M.n305 VSUBS 0.00845f
C384 M.n306 VSUBS 0.00233f
C385 M.n307 VSUBS 0.00991f
C386 M.n308 VSUBS 0.00962f
C387 M.n309 VSUBS 0.00204f
C388 M.n310 VSUBS 0.00845f
C389 M.n311 VSUBS 0.00845f
C390 M.n312 VSUBS 0.00583f
C391 M.n313 VSUBS 0.00583f
C392 M.n314 VSUBS 0.0108f
C393 M.n315 VSUBS 0.0195f
C394 M.n316 VSUBS 0.0105f
C395 M.n317 VSUBS 0.0178f
C396 M.n318 VSUBS 0.0178f
C397 M.n319 VSUBS 0.0108f
C398 M.n320 VSUBS 0.0108f
C399 M.n321 VSUBS 0.00729f
C400 M.n322 VSUBS 0.00729f
C401 M.n323 VSUBS 0.00233f
C402 M.n324 VSUBS 0.00233f
C403 M.n325 VSUBS 0.00117f
C404 M.n326 VSUBS 0.00758f
C405 M.n327 VSUBS 0.00962f
C406 M.n328 VSUBS 0.00321f
C407 M.n329 VSUBS 0.00729f
C408 M.n330 VSUBS 0.00729f
C409 M.n331 VSUBS 0.0294f
C410 M.n332 VSUBS 0.0294f
C411 M.n333 VSUBS 0.0108f
C412 M.n334 VSUBS 0.0114f
C413 M.n335 VSUBS 0.00233f
C414 M.n336 VSUBS 0.00816f
C415 M.n337 VSUBS 0.00816f
C416 M.n338 VSUBS 0.00262f
C417 M.n339 VSUBS 0.0114f
C418 M.n340 VSUBS 0.0495f
C419 M.n341 VSUBS 0.00845f
C420 M.n342 VSUBS 0.00321f
C421 M.n343 VSUBS 0.0108f
C422 M.n344 VSUBS 0.0105f
C423 M.n345 VSUBS 0.00291f
C424 M.n346 VSUBS 0.00845f
C425 M.n347 VSUBS 0.00845f
C426 M.n348 VSUBS 0.00408f
C427 M.n349 VSUBS 0.00408f
C428 M.n350 VSUBS 0.0117f
C429 M.n351 VSUBS 0.0213f
C430 M.n352 VSUBS 0.0114f
C431 M.n353 VSUBS 0.016f
C432 M.n354 VSUBS 0.016f
C433 M.n355 VSUBS 0.0108f
C434 M.n356 VSUBS 0.0108f
C435 M.n357 VSUBS 0.00729f
C436 M.n358 VSUBS 0.00729f
C437 M.n359 VSUBS 0.00408f
C438 M.n360 VSUBS 0.0035f
C439 M.n361 VSUBS 8.74e-19
C440 M.n362 VSUBS 0.00729f
C441 M.n363 VSUBS 0.00991f
C442 M.n364 VSUBS 0.00408f
C443 M.n365 VSUBS 0.00729f
C444 M.n366 VSUBS 0.00729f
C445 M.n367 VSUBS 0.0277f
C446 M.n368 VSUBS 0.0277f
C447 M.n369 VSUBS 0.0117f
C448 M.n370 VSUBS 0.0114f
C449 M.n371 VSUBS 0.00146f
C450 M.n372 VSUBS 0.00991f
C451 M.n373 VSUBS 0.00991f
C452 M.n374 VSUBS 0.00175f
C453 M.n375 VSUBS 0.0114f
C454 M.n376 VSUBS 0.0122f
C455 M.n377 VSUBS 0.0117f
C456 M.n378 VSUBS 0.0114f
C457 M.n379 VSUBS 0.0122f
C458 M.n380 VSUBS 0.0385f
C459 M.n381 VSUBS 0.0341f
C460 M.n382 VSUBS 0.0114f
C461 M.n383 VSUBS 0.474f
C462 M.n384 VSUBS 0.00729f
C463 M.n385 VSUBS 0.00495f
C464 M.n386 VSUBS 0.0108f
C465 M.n387 VSUBS 0.00729f
C466 M.n388 VSUBS 0.0117f
C467 M.n389 VSUBS 0.0259f
C468 M.n390 VSUBS 0.0265f
C469 M.n391 VSUBS 0.023f
C470 M.n392 VSUBS 0.0149f
C471 M.n393 VSUBS 0.0117f
C472 M.n394 VSUBS 0.0114f
C473 M.n395 VSUBS 0.0114f
C474 M.n396 VSUBS 0.0117f
C475 M.n397 VSUBS 0.0117f
C476 M.n398 VSUBS 1.31f
C477 M.n399 VSUBS 1.32f
C478 M.n400 VSUBS 0.0729f
C479 M.n401 VSUBS 0.181f
C480 M.n402 VSUBS 0.0577f
C481 M.n403 VSUBS 0.0554f
C482 M.n404 VSUBS 0.00729f
C483 M.n405 VSUBS 0.0568f
C484 M.n406 VSUBS 0.0119f
C485 M.n407 VSUBS 0.0458f
C486 M.n408 VSUBS 0.0627f
C487 M.n409 VSUBS 0.106f
C488 M.n410 VSUBS 0.0628f
C489 M.n411 VSUBS 0.00962f
C490 M.n412 VSUBS 0.00991f
C491 M.n413 VSUBS 0.0102f
C492 M.n414 VSUBS 0.0137f
C493 M.n415 VSUBS 0.014f
C494 M.n416 VSUBS 0.0195f
C495 M.n417 VSUBS 0.0291f
C496 M.n418 VSUBS 0.0262f
C497 M.n419 VSUBS 0.00991f
C498 M.n420 VSUBS 0.00525f
C499 M.n421 VSUBS 0.0067f
C500 M.n422 VSUBS 0.00758f
C501 M.n423 VSUBS 0.00525f
C502 M.n424 VSUBS 0.0067f
C503 M.n425 VSUBS 0.00962f
C504 M.n426 VSUBS 0.0373f
C505 M.n427 VSUBS 0.0358f
C506 M.n428 VSUBS 0.00729f
C507 M.n429 VSUBS 0.00612f
C508 M.n430 VSUBS 0.00641f
C509 M.n431 VSUBS 0.00729f
C510 M.n432 VSUBS 0.00583f
C511 M.n433 VSUBS 0.00612f
C512 M.n434 VSUBS 0.00729f
C513 M.n435 VSUBS 0.0382f
C514 M.n436 VSUBS 0.0446f
C515 M.n437 VSUBS 0.0195f
C516 M.n438 VSUBS 0.0119f
C517 M.n439 VSUBS 0.0122f
C518 M.n440 VSUBS 0.0937f
C519 M.n441 VSUBS 0.0737f
C520 M.n442 VSUBS 0.0195f
C521 M.n443 VSUBS 0.021f
C522 M.n444 VSUBS 0.022f
C523 M.n445 VSUBS 0.0117f
C524 M.n446 VSUBS 0.0114f
C525 M.n447 VSUBS 0.0108f
C526 M.n448 VSUBS 8.74e-19
C527 M.n449 VSUBS 8.74e-19
C528 M.n450 VSUBS 0.0105f
C529 M.n451 VSUBS 0.0321f
C530 M.n452 VSUBS 0.0117f
C531 M.n453 VSUBS 0.0108f
C532 M.n454 VSUBS 0.00146f
C533 M.n455 VSUBS 0.00146f
C534 M.n456 VSUBS 0.0105f
C535 M.n457 VSUBS 0.0338f
C536 M.n458 VSUBS 0.0108f
C537 M.n459 VSUBS 0.0195f
C538 M.n460 VSUBS 0.021f
C539 M.n461 VSUBS 0.022f
C540 M.n462 VSUBS 0.0431f
C541 M.n463 VSUBS 0.0349f
C542 M.n464 VSUBS 0.00733f
C543 M.n465 VSUBS 0.00792f
C544 M.n466 VSUBS 0.0321f
C545 M.n467 VSUBS 0.0035f
C546 M.n468 VSUBS 0.0035f
C547 M.n469 VSUBS 0.00379f
C548 M.n470 VSUBS 0.00379f
C549 M.n471 VSUBS 0.00408f
C550 M.n472 VSUBS 0.0338f
C551 M.n473 VSUBS 0.0035f
C552 M.n474 VSUBS 0.0035f
C553 M.n475 VSUBS 0.00379f
C554 M.n476 VSUBS 0.00379f
C555 M.n477 VSUBS 0.00321f
C556 M.n478 VSUBS 0.00583f
C557 M.n479 VSUBS 0.0067f
C558 M.n480 VSUBS 0.00762f
C559 M.n481 VSUBS 0.00729f
C560 M.n482 VSUBS 0.00729f
C561 M.n483 VSUBS 0.00733f
C562 M.n484 VSUBS 0.0294f
C563 M.n485 VSUBS 0.00379f
C564 M.n486 VSUBS 0.00379f
C565 M.n487 VSUBS 0.0035f
C566 M.n488 VSUBS 0.0035f
C567 M.n489 VSUBS 0.00437f
C568 M.n490 VSUBS 0.0312f
C569 M.n491 VSUBS 0.00379f
C570 M.n492 VSUBS 0.00379f
C571 M.n493 VSUBS 0.0035f
C572 M.n494 VSUBS 0.0035f
C573 M.n495 VSUBS 0.0035f
C574 M.n496 VSUBS 0.00641f
C575 M.n497 VSUBS 0.00729f
C576 M.n498 VSUBS 0.00821f
C577 M.n499 VSUBS 0.00792f
C578 M.n500 VSUBS 0.00733f
C579 M.n501 VSUBS 0.0325f
C580 M.n502 VSUBS 0.034f
C581 M.n503 VSUBS 0.00557f
C582 M.n504 VSUBS 0.476f
C583 M.n505 VSUBS 0.0294f
C584 M.n506 VSUBS 0.00525f
C585 M.n507 VSUBS 0.00525f
C586 M.n508 VSUBS 0.00612f
C587 M.n509 VSUBS 0.0312f
C588 M.n510 VSUBS 0.00525f
C589 M.n511 VSUBS 0.00525f
C590 M.n512 VSUBS 0.00525f
C591 M.n513 VSUBS 0.00379f
C592 M.n514 VSUBS 0.00233f
C593 M.n515 VSUBS 0.00583f
C594 M.n516 VSUBS 0.00466f
C595 M.n517 VSUBS 0.00146f
C596 M.n518 VSUBS 0.00583f
C597 M.n519 VSUBS 0.00645f
C598 M.n520 VSUBS 0.00528f
C599 M.n521 VSUBS 0.00758f
C600 M.n522 VSUBS 0.00933f
C601 M.n523 VSUBS 0.0111f
C602 M.n524 VSUBS 0.00674f
C603 M.n525 VSUBS 0.00641f
C604 M.n526 VSUBS 0.00117f
C605 M.n527 VSUBS 0.00554f
C606 M.n528 VSUBS 0.00204f
C607 M.n529 VSUBS 0.0187f
C608 M.n530 VSUBS 0.0067f
C609 M.n531 VSUBS 0.0067f
C610 M.n532 VSUBS 0.00408f
C611 M.n533 VSUBS 0.00437f
C612 M.n534 VSUBS 0.0169f
C613 M.n535 VSUBS 0.0067f
C614 M.n536 VSUBS 0.0067f
C615 M.n537 VSUBS 0.00495f
C616 M.n538 VSUBS 0.00437f
C617 M.n539 VSUBS 0.00528f
C618 M.n540 VSUBS 0.0117f
C619 M.n541 VSUBS 0.0229f
C620 M.n542 VSUBS 0.0276f
C621 M.n543 VSUBS 0.0169f
C622 M.n544 VSUBS 0.0114f
C623 M.n545 VSUBS 0.0187f
C624 M.n546 VSUBS 0.0105f
C625 M.n547 VSUBS 0.0195f
C626 M.n548 VSUBS 0.0213f
C627 M.n549 VSUBS 0.0232f
C628 M.n550 VSUBS 0.0123f
C629 M.n551 VSUBS 0.0108f
C630 M.n552 VSUBS 0.0114f
C631 M.n553 VSUBS 0.0117f
C632 M.n554 VSUBS 0.00146f
C633 M.n555 VSUBS 0.00146f
C634 M.n556 VSUBS 0.0102f
C635 M.n557 VSUBS 0.0102f
C636 M.n558 VSUBS 0.00117f
C637 M.n559 VSUBS 0.0108f
C638 M.n560 VSUBS 0.00321f
C639 M.n561 VSUBS 0.00321f
C640 M.n562 VSUBS 0.0102f
C641 M.n563 VSUBS 0.00962f
C642 M.n564 VSUBS 0.00991f
C643 M.n565 VSUBS 8.74e-19
C644 M.n566 VSUBS 0.0105f
C645 M.n567 VSUBS 0.0114f
C646 M.n568 VSUBS 0.00962f
C647 M.n569 VSUBS 0.0519f
C648 M.n570 VSUBS 0.00991f
C649 M.n571 VSUBS 8.74e-19
C650 M.n572 VSUBS 0.0501f
C651 M.n573 VSUBS 0.0102f
C652 M.n574 VSUBS 0.00146f
C653 M.n575 VSUBS 0.0108f
C654 M.n576 VSUBS 0.0117f
C655 M.n577 VSUBS 0.0117f
C656 M.n578 VSUBS 1.33f
C657 M.n579 VSUBS 1.33f
C658 M.n580 VSUBS 0.0537f
C659 M.n581 VSUBS 0.155f
C660 M.n582 VSUBS 0.0449f
C661 M.n583 VSUBS 0.00962f
C662 M.n584 VSUBS 0.00962f
C663 M.n585 VSUBS 0.0254f
C664 M.n586 VSUBS 0.0268f
C665 M.n587 VSUBS 0.0195f
C666 M.n588 VSUBS 0.0175f
C667 M.n589 VSUBS 0.0178f
C668 M.n590 VSUBS 0.0745f
C669 M.n591 VSUBS 0.0545f
C670 M.n592 VSUBS 0.0195f
C671 M.n593 VSUBS 0.0213f
C672 M.n594 VSUBS 0.0232f
C673 M.n595 VSUBS 0.0161f
C674 M.n596 VSUBS 0.0158f
C675 M.n597 VSUBS 0.0117f
C676 M.n598 VSUBS 0.00525f
C677 M.n599 VSUBS 0.00525f
C678 M.n600 VSUBS 0.0114f
C679 M.n601 VSUBS 0.0117f
C680 M.n602 VSUBS 0.0108f
C681 M.n603 VSUBS 0.00699f
C682 M.n604 VSUBS 0.00699f
C683 M.n605 VSUBS 0.0105f
C684 M.n606 VSUBS 0.0108f
C685 M.n607 VSUBS 0.0195f
C686 M.n608 VSUBS 0.0213f
C687 M.n609 VSUBS 0.0232f
C688 M.n610 VSUBS 0.0252f
C689 M.n611 VSUBS 0.022f
C690 M.n612 VSUBS 0.0114f
C691 M.n613 VSUBS 0.0143f
C692 M.n614 VSUBS 0.0143f
C693 M.n615 VSUBS 0.00845f
C694 M.n616 VSUBS 0.00845f
C695 M.n617 VSUBS 0.00291f
C696 M.n618 VSUBS 0.016f
C697 M.n619 VSUBS 0.016f
C698 M.n620 VSUBS 0.00845f
C699 M.n621 VSUBS 0.00845f
C700 M.n622 VSUBS 0.00204f
C701 M.n623 VSUBS 0.00962f
C702 M.n624 VSUBS 0.0105f
C703 M.n625 VSUBS 0.0114f
C704 M.n626 VSUBS 0.00466f
C705 M.n627 VSUBS 0.00379f
C706 M.n628 VSUBS 0.00379f
C707 M.n629 VSUBS 0.00233f
C708 M.n630 VSUBS 0.00991f
C709 M.n631 VSUBS 0.00641f
C710 M.n632 VSUBS 0.00204f
C711 M.n633 VSUBS 0.00204f
C712 M.n634 VSUBS 0.00321f
C713 M.n635 VSUBS 0.0108f
C714 M.n636 VSUBS 0.0117f
C715 M.n637 VSUBS 0.0044f
C716 M.n638 VSUBS 0.0085f
C717 M.n639 VSUBS 0.0114f
C718 M.n640 VSUBS 0.00641f
C719 M.n641 VSUBS 0.00495f
C720 M.n642 VSUBS 0.00466f
C721 M.n643 VSUBS 0.00583f
C722 M.n644 VSUBS 0.0149f
C723 M.n645 VSUBS 0.0149f
C724 M.n646 VSUBS 0.0158f
C725 M.n647 VSUBS 0.0179f
C726 M.n648 VSUBS 0.0144f
C727 M.n649 VSUBS 0.478f
C728 M.n650 VSUBS 0.00322f
C729 M.n651 VSUBS 0.0117f
C730 M.n652 VSUBS 0.00699f
C731 M.n653 VSUBS 0.00699f
C732 M.n654 VSUBS 0.0102f
C733 M.n655 VSUBS 0.0102f
C734 M.n656 VSUBS 0.00117f
C735 M.n657 VSUBS 0.0108f
C736 M.n658 VSUBS 0.00874f
C737 M.n659 VSUBS 0.00874f
C738 M.n660 VSUBS 0.0102f
C739 M.n661 VSUBS 0.00962f
C740 M.n662 VSUBS 0.00991f
C741 M.n663 VSUBS 8.74e-19
C742 M.n664 VSUBS 0.0105f
C743 M.n665 VSUBS 0.0114f
C744 M.n666 VSUBS 0.00554f
C745 M.n667 VSUBS 0.00466f
C746 M.n668 VSUBS 0.00466f
C747 M.n669 VSUBS 0.00146f
C748 M.n670 VSUBS 0.00962f
C749 M.n671 VSUBS 0.00641f
C750 M.n672 VSUBS 0.00612f
C751 M.n673 VSUBS 8.74e-19
C752 M.n674 VSUBS 0.0108f
C753 M.n675 VSUBS 0.0117f
C754 M.n676 VSUBS 0.00528f
C755 M.n677 VSUBS 0.0103f
C756 M.n678 VSUBS 0.0114f
C757 M.n679 VSUBS 0.00554f
C758 M.n680 VSUBS 0.00583f
C759 M.n681 VSUBS 0.00379f
C760 M.n682 VSUBS 0.00379f
C761 M.n683 VSUBS 0.0067f
C762 M.n684 VSUBS 0.0157f
C763 M.n685 VSUBS 0.0157f
C764 M.n686 VSUBS 0.0167f
C765 M.n687 VSUBS 0.0141f
C766 M.n688 VSUBS 0.0138f
C767 M.n689 VSUBS 0.0117f
C768 M.n690 VSUBS 0.00321f
C769 M.n691 VSUBS 0.00321f
C770 M.n692 VSUBS 0.0114f
C771 M.n693 VSUBS 0.0108f
C772 M.n694 VSUBS 0.00495f
C773 M.n695 VSUBS 0.00495f
C774 M.n696 VSUBS 0.0105f
C775 M.n697 VSUBS 0.0195f
C776 M.n698 VSUBS 0.021f
C777 M.n699 VSUBS 0.022f
C778 M.n700 VSUBS 0.0117f
C779 M.n701 VSUBS 0.0114f
C780 M.n702 VSUBS 0.0108f
C781 M.n703 VSUBS 8.74e-19
C782 M.n704 VSUBS 8.74e-19
C783 M.n705 VSUBS 0.0105f
C784 M.n706 VSUBS 0.0108f
C785 M.n707 VSUBS 0.00146f
C786 M.n708 VSUBS 0.00146f
C787 M.n709 VSUBS 0.0105f
C788 M.n710 VSUBS 0.0175f
C789 M.n711 VSUBS 0.0172f
C790 M.n712 VSUBS 0.0173f
C791 M.n713 VSUBS 0.0117f
C792 M.n714 VSUBS 0.0114f
C793 M.n715 VSUBS 0.00787f
C794 M.n716 VSUBS 0.00379f
C795 M.n717 VSUBS 0.00379f
C796 M.n718 VSUBS 0.00758f
C797 M.n719 VSUBS 0.00874f
C798 M.n720 VSUBS 0.00204f
C799 M.n721 VSUBS 0.00204f
C800 M.n722 VSUBS 0.00845f
C801 M.n723 VSUBS 0.0242f
C802 M.n724 VSUBS 0.00991f
C803 M.n725 VSUBS 0.00612f
C804 M.n726 VSUBS 0.00845f
C805 M.n727 VSUBS 0.00962f
C806 M.n728 VSUBS 0.0449f
C807 M.n729 VSUBS 0.0157f
C808 M.n730 VSUBS 0.0195f
C809 M.n731 VSUBS 0.0192f
C810 M.n732 VSUBS 0.0393f
C811 M.n733 VSUBS 0.0102f
C812 M.n734 VSUBS 0.00991f
C813 M.n735 VSUBS 0.00962f
C814 M.n736 VSUBS 0.0268f
C815 M.n737 VSUBS 0.00729f
C816 M.n738 VSUBS 0.00991f
C817 M.n739 VSUBS 0.00962f
C818 M.n740 VSUBS 0.042f
C819 M.n741 VSUBS 0.0166f
C820 M.n742 VSUBS 0.0157f
C821 M.n743 VSUBS 0.0154f
C822 M.n744 VSUBS 0.0472f
C823 M.n745 VSUBS 0.0195f
C824 M.n746 VSUBS 0.0122f
C825 M.n747 VSUBS 0.0119f
C826 M.n748 VSUBS 0.16f
C827 M.n749 VSUBS 0.0184f
C828 M.n750 VSUBS 0.00991f
C829 M.n751 VSUBS 0.00962f
C830 M.n752 VSUBS 0.111f
C831 M.n753 VSUBS 0.0921f
C832 M.n754 VSUBS 0.0175f
C833 M.n755 VSUBS 0.0914f
C834 M.n756 VSUBS 0.0175f
C835 M.n757 VSUBS 0.0185f
C836 M.n758 VSUBS 1.27f
C837 M.n759 VSUBS 0.0125f
C838 M.n760 VSUBS 0.00235f
C839 M.n761 VSUBS 0.00207f
C840 M.n762 VSUBS 0.0128f
C841 M.n763 VSUBS 0.00207f
C842 M.n764 VSUBS 0.0149f
C843 M.n765 VSUBS 0.0133f
C844 M.n766 VSUBS 0.00798f
C845 M.n767 VSUBS 0.00375f
C846 M.n768 VSUBS 0.00224f
C847 M.n769 VSUBS 0.00775f
C848 M.n770 VSUBS 0.0143f
C849 M.n771 VSUBS 0.00828f
C850 M.n772 VSUBS 1.24f
C851 M.n773 VSUBS 0.0675f
C852 M.n774 VSUBS 0.0686f
C853 M.n775 VSUBS 0.0114f
C854 M.n776 VSUBS 0.0706f
C855 M.n777 VSUBS 0.0105f
C856 M.n778 VSUBS 0.0195f
C857 M.n779 VSUBS 0.0213f
C858 M.n780 VSUBS 0.023f
C859 M.n781 VSUBS 0.0195f
C860 M.n782 VSUBS 0.0192f
C861 M.n783 VSUBS 0.0117f
C862 M.n784 VSUBS 0.00874f
C863 M.n785 VSUBS 0.00874f
C864 M.n786 VSUBS 0.0114f
C865 M.n787 VSUBS 0.0108f
C866 M.n788 VSUBS 0.0105f
C867 M.n789 VSUBS 0.0105f
C868 M.n790 VSUBS 0.0105f
C869 M.n791 VSUBS 0.0195f
C870 M.n792 VSUBS 0.0213f
C871 M.n793 VSUBS 0.023f
C872 M.n794 VSUBS 0.0222f
C873 M.n795 VSUBS 0.0219f
C874 M.n796 VSUBS 0.0117f
C875 M.n797 VSUBS 0.0114f
C876 M.n798 VSUBS 0.0114f
C877 M.n799 VSUBS 0.0114f
C878 M.n800 VSUBS 0.0108f
C879 M.n801 VSUBS 0.0131f
C880 M.n802 VSUBS 0.0131f
C881 M.n803 VSUBS 0.0105f
C882 M.n804 VSUBS 0.0195f
C883 M.n805 VSUBS 0.0213f
C884 M.n806 VSUBS 0.023f
C885 M.n807 VSUBS 0.0201f
C886 M.n808 VSUBS 0.0134f
C887 M.n809 VSUBS 0.0114f
C888 M.n810 VSUBS 0.0117f
C889 M.n811 VSUBS 0.00933f
C890 M.n812 VSUBS 0.00933f
C891 M.n813 VSUBS 0.00495f
C892 M.n814 VSUBS 0.00495f
C893 M.n815 VSUBS 0.00641f
C894 M.n816 VSUBS 0.0108f
C895 M.n817 VSUBS 0.0111f
C896 M.n818 VSUBS 0.0111f
C897 M.n819 VSUBS 0.00495f
C898 M.n820 VSUBS 0.00495f
C899 M.n821 VSUBS 0.00554f
C900 M.n822 VSUBS 0.00962f
C901 M.n823 VSUBS 0.0105f
C902 M.n824 VSUBS 0.0114f
C903 M.n825 VSUBS 0.00495f
C904 M.n826 VSUBS 0.00175f
C905 M.n827 VSUBS 0.00495f
C906 M.n828 VSUBS 0.00904f
C907 M.n829 VSUBS 0.00495f
C908 M.n830 VSUBS 0.00262f
C909 M.n831 VSUBS 0.00262f
C910 M.n832 VSUBS 0.00408f
C911 M.n833 VSUBS 0.00816f
C912 M.n834 VSUBS 0.00816f
C913 M.n835 VSUBS 0.0067f
C914 M.n836 VSUBS 0.00845f
C915 M.n837 VSUBS 0.00787f
C916 M.n838 VSUBS 0.00495f
C917 M.n839 VSUBS 0.00379f
C918 M.n840 VSUBS 0.0256f
C919 M.n841 VSUBS 0.0117f
C920 M.n842 VSUBS 0.00495f
C921 M.n843 VSUBS 0.00466f
C922 M.n844 VSUBS 0.0274f
C923 M.n845 VSUBS 0.0108f
C924 M.n846 VSUBS 0.0137f
C925 M.n847 VSUBS 0.0137f
C926 M.n848 VSUBS 0.0146f
C927 M.n849 VSUBS 0.0361f
C928 M.n850 VSUBS 0.492f
C929 M.n851 VSUBS 0.00525f
C930 M.n852 VSUBS 0.00612f
C931 M.n853 VSUBS 0.00641f
C932 M.n854 VSUBS 0.0256f
C933 M.n855 VSUBS 0.00495f
C934 M.n856 VSUBS 0.00495f
C935 M.n857 VSUBS 0.00117f
C936 M.n858 VSUBS 0.00117f
C937 M.n859 VSUBS 0.00525f
C938 M.n860 VSUBS 0.0274f
C939 M.n861 VSUBS 0.00495f
C940 M.n862 VSUBS 0.00495f
C941 M.n863 VSUBS 0.00117f
C942 M.n864 VSUBS 0.00117f
C943 M.n865 VSUBS 0.00437f
C944 M.n866 VSUBS 0.00845f
C945 M.n867 VSUBS 0.00933f
C946 M.n868 VSUBS 0.0102f
C947 M.n869 VSUBS 0.00612f
C948 M.n870 VSUBS 0.00612f
C949 M.n871 VSUBS 0.00612f
C950 M.n872 VSUBS 0.0472f
C951 M.n873 VSUBS 0.00117f
C952 M.n874 VSUBS 0.00117f
C953 M.n875 VSUBS 0.00495f
C954 M.n876 VSUBS 0.00495f
C955 M.n877 VSUBS 0.00554f
C956 M.n878 VSUBS 0.049f
C957 M.n879 VSUBS 0.00117f
C958 M.n880 VSUBS 0.00117f
C959 M.n881 VSUBS 0.00495f
C960 M.n882 VSUBS 0.00495f
C961 M.n883 VSUBS 0.00466f
C962 M.n884 VSUBS 0.00495f
C963 M.n885 VSUBS 0.00583f
C964 M.n886 VSUBS 0.0067f
C965 M.n887 VSUBS 0.0105f
C966 M.n888 VSUBS 0.00612f
C967 M.n889 VSUBS 0.0475f
C968 M.n890 VSUBS 0.0577f
C969 M.n891 VSUBS 0.0472f
C970 M.n892 VSUBS 0.0114f
C971 M.n893 VSUBS 0.049f
C972 M.n894 VSUBS 0.0105f
C973 M.n895 VSUBS 0.0812f
C974 M.n896 VSUBS 0.147f
C975 M.n897 VSUBS 0.0195f
C976 M.n898 VSUBS 0.0213f
C977 M.n899 VSUBS 0.021f
C978 M.n900 VSUBS 0.0644f
C979 M.n901 VSUBS 0.0195f
C980 M.n902 VSUBS 0.0239f
C981 M.n903 VSUBS 0.0236f
C982 M.n904 VSUBS 0.065f
C983 M.n905 VSUBS 0.0195f
C984 M.n906 VSUBS 0.0219f
C985 M.n907 VSUBS 0.0169f
C986 M.n908 VSUBS 0.00962f
C987 M.n909 VSUBS 0.0364f
C988 M.n910 VSUBS 0.00962f
C989 M.n911 VSUBS 0.0195f
C990 M.n912 VSUBS 0.00991f
C991 M.n913 VSUBS 0.00991f
C992 M.n914 VSUBS 0.00962f
C993 M.n915 VSUBS 0.0624f
C994 M.n916 VSUBS 0.0146f
C995 M.n917 VSUBS 0.0382f
C996 M.n918 VSUBS 0.0332f
C997 M.n919 VSUBS 0.00612f
C998 M.n920 VSUBS 0.00466f
C999 M.n921 VSUBS 0.00845f
C1000 M.n922 VSUBS 0.0528f
C1001 M.n923 VSUBS 0.00612f
C1002 M.n924 VSUBS 0.00612f
C1003 M.n925 VSUBS 0.194f
C1004 M.n926 VSUBS 0.00495f
C1005 M.n927 VSUBS 0.00874f
C1006 M.n928 VSUBS 0.00612f
C1007 M.n929 VSUBS 0.051f
C1008 M.n930 VSUBS 0.0595f
C1009 M.n931 VSUBS 0.0667f
C1010 M.n932 VSUBS 0.0454f
C1011 M.n933 VSUBS 0.0195f
C1012 M.n934 VSUBS 0.0447f
C1013 M.n935 VSUBS 0.0213f
C1014 M.n936 VSUBS 0.023f
C1015 M.n937 VSUBS 1.29f
C1016 M.n938 VSUBS 0.134f
C1017 M.n939 VSUBS 0.0543f
C1018 M.n940 VSUBS 0.0548f
C1019 M.n941 VSUBS 0.0307f
C1020 M.n942 VSUBS 0.0165f
C1021 M.n943 VSUBS 0.0526f
C1022 M.n944 VSUBS 0.00516f
C1023 M.n945 VSUBS 0.0445f
C1024 M.n946 VSUBS 0.043f
C1025 M.n947 VSUBS 0.00516f
C1026 M.n948 VSUBS 0.00737f
C1027 M.n949 VSUBS 0.16f
C1028 M.n950 VSUBS 0.00418f
C1029 M.n951 VSUBS 0.00516f
C1030 M.n952 VSUBS 0.00713f
C1031 M.n953 VSUBS 0.00393f
C1032 M.n954 VSUBS 0.00516f
C1033 M.n955 VSUBS 0.028f
C1034 M.n956 VSUBS 0.0322f
C1035 M.n957 VSUBS 0.0123f
C1036 M.n958 VSUBS 0.00811f
C1037 M.n959 VSUBS 0.00835f
C1038 M.n960 VSUBS 0.00835f
C1039 M.n961 VSUBS 0.00811f
C1040 M.n962 VSUBS 0.00811f
C1041 M.n963 VSUBS 0.0143f
C1042 M.n964 VSUBS 0.0184f
C1043 M.n965 VSUBS 0.0165f
C1044 M.n966 VSUBS 0.0199f
C1045 M.n967 VSUBS 0.0201f
C1046 M.n968 VSUBS 0.0165f
C1047 M.n969 VSUBS 0.0177f
C1048 M.n970 VSUBS 0.0179f
C1049 M.n971 VSUBS 0.0165f
C1050 M.n972 VSUBS 0.0302f
C1051 M.n973 VSUBS 0.0305f
C1052 M.n974 VSUBS 0.041f
C1053 M.n975 VSUBS 0.0239f
C1054 M.n976 VSUBS 0.00885f
C1055 M.n977 VSUBS 0.0214f
C1056 M.n978 VSUBS 0.0214f
C1057 M.n979 VSUBS 0.00909f
C1058 M.n980 VSUBS 0.0165f
C1059 M.n981 VSUBS 0.00885f
C1060 M.n982 VSUBS 0.00885f
C1061 M.n983 VSUBS 0.00885f
C1062 M.n984 VSUBS 0.00909f
C1063 M.n985 VSUBS 0.0165f
C1064 M.n986 VSUBS 0.00811f
C1065 M.n987 VSUBS 0.00393f
C1066 M.n988 VSUBS 0.00418f
C1067 M.n989 VSUBS 0.00418f
C1068 M.n990 VSUBS 0.00147f
C1069 M.n991 VSUBS 0.00418f
C1070 M.n992 VSUBS 0.00762f
C1071 M.n993 VSUBS 0.0398f
C1072 M.n994 VSUBS 9.83e-19
C1073 M.n995 VSUBS 9.83e-19
C1074 M.n996 VSUBS 0.00418f
C1075 M.n997 VSUBS 0.00418f
C1076 M.n998 VSUBS 0.00467f
C1077 M.n999 VSUBS 0.0413f
C1078 M.n1000 VSUBS 9.83e-19
C1079 M.n1001 VSUBS 9.83e-19
C1080 M.n1002 VSUBS 0.00418f
C1081 M.n1003 VSUBS 0.00418f
C1082 M.n1004 VSUBS 0.00393f
C1083 M.n1005 VSUBS 0.00418f
C1084 M.n1006 VSUBS 0.00491f
C1085 M.n1007 VSUBS 0.00516f
C1086 M.n1008 VSUBS 0.00516f
C1087 M.n1009 VSUBS 0.00713f
C1088 M.n1010 VSUBS 0.00786f
C1089 M.n1011 VSUBS 0.00442f
C1090 M.n1012 VSUBS 9.83e-19
C1091 M.n1013 VSUBS 9.83e-19
C1092 M.n1014 VSUBS 0.00418f
C1093 M.n1015 VSUBS 0.00418f
C1094 M.n1016 VSUBS 0.0216f
C1095 M.n1017 VSUBS 0.0216f
C1096 M.n1018 VSUBS 0.00983f
C1097 M.n1019 VSUBS 0.00369f
C1098 M.n1020 VSUBS 9.83e-19
C1099 M.n1021 VSUBS 9.83e-19
C1100 M.n1022 VSUBS 0.00418f
C1101 M.n1023 VSUBS 0.00418f
C1102 M.n1024 VSUBS 0.0231f
C1103 M.n1025 VSUBS 0.0231f
C1104 M.n1026 VSUBS 0.00909f
C1105 M.n1027 VSUBS 0.0115f
C1106 M.n1028 VSUBS 0.0115f
C1107 M.n1029 VSUBS 0.00319f
C1108 M.n1030 VSUBS 0.00418f
C1109 M.n1031 VSUBS 0.00418f
C1110 M.n1032 VSUBS 0.00221f
C1111 M.n1033 VSUBS 0.00221f
C1112 M.n1034 VSUBS 0.00344f
C1113 M.n1035 VSUBS 0.00688f
C1114 M.n1036 VSUBS 0.00885f
C1115 M.n1037 VSUBS 0.00541f
C1116 M.n1038 VSUBS 0.00418f
C1117 M.n1039 VSUBS 0.00418f
C1118 M.n1040 VSUBS 0.00786f
C1119 M.n1041 VSUBS 0.00786f
C1120 M.n1042 VSUBS 0.00983f
C1121 M.n1043 VSUBS 0.00467f
C1122 M.n1044 VSUBS 0.00418f
C1123 M.n1045 VSUBS 0.00418f
C1124 M.n1046 VSUBS 0.00934f
C1125 M.n1047 VSUBS 0.00934f
C1126 M.n1048 VSUBS 0.00909f
C1127 M.n1049 VSUBS 0.0165f
C1128 M.n1050 VSUBS 0.0179f
C1129 M.n1051 VSUBS 0.00958f
C1130 M.n1052 VSUBS 0.00958f
C1131 M.n1053 VSUBS 0.00958f
C1132 M.n1054 VSUBS 0.00983f
C1133 M.n1055 VSUBS 0.00885f
C1134 M.n1056 VSUBS 0.0111f
C1135 M.n1057 VSUBS 0.0111f
C1136 M.n1058 VSUBS 0.00909f
C1137 M.n1059 VSUBS 0.0165f
C1138 M.n1060 VSUBS 0.0179f
C1139 M.n1061 VSUBS 0.00958f
C1140 M.n1062 VSUBS 0.00737f
C1141 M.n1063 VSUBS 0.00737f
C1142 M.n1064 VSUBS 0.00983f
C1143 M.n1065 VSUBS 0.0179f
C1144 M.n1066 VSUBS 0.00958f
C1145 M.n1067 VSUBS 0.0199f
C1146 M.n1068 VSUBS 0.0199f
C1147 M.n1069 VSUBS 0.00983f
C1148 M.n1070 VSUBS 0.018f
C1149 M.n1071 VSUBS 0.024f
C1150 M.n1072 VSUBS 1.28f
C1151 M.n1073 VSUBS 0.0595f
C1152 M.n1074 VSUBS 0.0392f
C1153 M.n1075 VSUBS 0.0264f
C1154 M.n1076 VSUBS 0.0224f
C1155 M.n1077 VSUBS 0.0221f
C1156 M.n1078 VSUBS 0.0264f
C1157 M.n1079 VSUBS 0.0254f
C1158 M.n1080 VSUBS 0.0251f
C1159 M.n1081 VSUBS 0.0264f
C1160 M.n1082 VSUBS 0.0231f
C1161 M.n1083 VSUBS 0.0154f
C1162 M.n1084 VSUBS 0.0131f
C1163 M.n1085 VSUBS 0.0131f
C1164 M.n1086 VSUBS 0.00937f
C1165 M.n1087 VSUBS 0.0077f
C1166 M.n1088 VSUBS 0.00971f
C1167 M.n1089 VSUBS 0.00904f
C1168 M.n1090 VSUBS 0.0164f
C1169 M.n1091 VSUBS 0.44f
C1170 M.n1092 VSUBS 0.0288f
C1171 M.n1093 VSUBS 0.0341f
C1172 M.n1094 VSUBS 0.00703f
C1173 M.n1095 VSUBS 0.00736f
C1174 M.n1096 VSUBS 0.0117f
C1175 M.n1097 VSUBS 0.00703f
C1176 M.n1098 VSUBS 0.0077f
C1177 M.n1099 VSUBS 0.012f
C1178 M.n1100 VSUBS 0.00703f
C1179 M.n1101 VSUBS 0.0546f
C1180 M.n1102 VSUBS 0.0663f
C1181 M.n1103 VSUBS 0.0398f
C1182 M.n1104 VSUBS 0.00958f
C1183 M.n1105 VSUBS 0.0413f
C1184 M.n1106 VSUBS 0.00885f
C1185 M.n1107 VSUBS 0.0501f
C1186 M.n1108 VSUBS 0.0535f
C1187 M.n1109 VSUBS 0.0354f
C1188 M.n1110 VSUBS 0.0165f
C1189 M.n1111 VSUBS 0.0347f
C1190 M.n1112 VSUBS 0.0179f
C1191 M.n1113 VSUBS 0.0264f
C1192 M.n1114 VSUBS 0.435f
C1193 M.t118 VSUBS 4.09f
C1194 M.t10 VSUBS 3.72f
C1195 M.n1115 VSUBS 1.84f
C1196 M.t69 VSUBS 3.72f
C1197 M.n1116 VSUBS 1.11f
C1198 M.t15 VSUBS 3.72f
C1199 M.n1117 VSUBS 1.11f
C1200 M.t22 VSUBS 3.72f
C1201 M.n1118 VSUBS 1.11f
C1202 M.t3 VSUBS 3.72f
C1203 M.n1119 VSUBS 1.11f
C1204 M.t85 VSUBS 3.72f
C1205 M.n1120 VSUBS 1.11f
C1206 M.t54 VSUBS 3.72f
C1207 M.n1121 VSUBS 1.11f
C1208 M.t1 VSUBS 3.72f
C1209 M.n1122 VSUBS 1.11f
C1210 M.t8 VSUBS 3.72f
C1211 M.n1123 VSUBS 1.11f
C1212 M.t119 VSUBS 3.72f
C1213 M.n1124 VSUBS 1.11f
C1214 M.t67 VSUBS 3.72f
C1215 M.n1125 VSUBS 0.856f
C1216 M.t71 VSUBS 4.09f
C1217 M.t64 VSUBS 3.72f
C1218 M.n1126 VSUBS 1.84f
C1219 M.t14 VSUBS 3.72f
C1220 M.n1127 VSUBS 1.11f
C1221 M.t92 VSUBS 3.72f
C1222 M.n1128 VSUBS 1.11f
C1223 M.t99 VSUBS 3.72f
C1224 M.n1129 VSUBS 1.11f
C1225 M.t83 VSUBS 3.72f
C1226 M.n1130 VSUBS 1.11f
C1227 M.t24 VSUBS 3.72f
C1228 M.n1131 VSUBS 1.11f
C1229 M.t7 VSUBS 3.72f
C1230 M.n1132 VSUBS 1.11f
C1231 M.t82 VSUBS 3.72f
C1232 M.n1133 VSUBS 1.11f
C1233 M.t88 VSUBS 3.72f
C1234 M.n1134 VSUBS 1.11f
C1235 M.t60 VSUBS 3.72f
C1236 M.n1135 VSUBS 1.11f
C1237 M.t12 VSUBS 3.72f
C1238 M.n1136 VSUBS 0.855f
C1239 M.n1137 VSUBS 0.0228f
C1240 M.n1138 VSUBS 0.00329f
C1241 M.n1139 VSUBS 0.00304f
C1242 M.n1140 VSUBS 7.6e-19
C1243 M.n1141 VSUBS 7.6e-19
C1244 M.n1142 VSUBS 0.00583f
C1245 M.n1143 VSUBS 0.0243f
C1246 M.n1144 VSUBS 0.00329f
C1247 M.n1145 VSUBS 0.00304f
C1248 M.n1146 VSUBS 7.6e-19
C1249 M.n1147 VSUBS 7.6e-19
C1250 M.n1148 VSUBS 0.00507f
C1251 M.n1149 VSUBS 0.00785f
C1252 M.n1150 VSUBS 0.00861f
C1253 M.t116 VSUBS 4.09f
C1254 M.t94 VSUBS 3.72f
C1255 M.n1151 VSUBS 1.84f
C1256 M.t97 VSUBS 3.72f
C1257 M.n1152 VSUBS 1.11f
C1258 M.t40 VSUBS 3.72f
C1259 M.n1153 VSUBS 1.11f
C1260 M.t53 VSUBS 3.72f
C1261 M.n1154 VSUBS 1.11f
C1262 M.t29 VSUBS 3.72f
C1263 M.n1155 VSUBS 1.11f
C1264 M.t114 VSUBS 3.72f
C1265 M.n1156 VSUBS 1.11f
C1266 M.t91 VSUBS 3.72f
C1267 M.n1157 VSUBS 1.11f
C1268 M.t27 VSUBS 3.72f
C1269 M.n1158 VSUBS 1.11f
C1270 M.t34 VSUBS 3.72f
C1271 M.n1159 VSUBS 1.11f
C1272 M.t18 VSUBS 3.72f
C1273 M.n1160 VSUBS 1.11f
C1274 M.t95 VSUBS 3.72f
C1275 M.n1161 VSUBS 0.853f
C1276 M.t122 VSUBS 4.09f
C1277 M.t44 VSUBS 3.72f
C1278 M.n1162 VSUBS 1.84f
C1279 M.t115 VSUBS 3.72f
C1280 M.n1163 VSUBS 1.11f
C1281 M.t59 VSUBS 3.72f
C1282 M.n1164 VSUBS 1.11f
C1283 M.t75 VSUBS 3.72f
C1284 M.n1165 VSUBS 1.11f
C1285 M.t41 VSUBS 3.72f
C1286 M.n1166 VSUBS 1.11f
C1287 M.t130 VSUBS 3.72f
C1288 M.n1167 VSUBS 1.11f
C1289 M.t102 VSUBS 3.72f
C1290 M.n1168 VSUBS 1.11f
C1291 M.t39 VSUBS 3.72f
C1292 M.n1169 VSUBS 1.11f
C1293 M.t51 VSUBS 3.72f
C1294 M.n1170 VSUBS 1.11f
C1295 M.t28 VSUBS 3.72f
C1296 M.n1171 VSUBS 1.11f
C1297 M.t113 VSUBS 3.72f
C1298 M.n1172 VSUBS 0.851f
C1299 M.t80 VSUBS 4.09f
C1300 M.t101 VSUBS 3.72f
C1301 M.n1173 VSUBS 1.84f
C1302 M.t58 VSUBS 3.72f
C1303 M.n1174 VSUBS 1.11f
C1304 M.t9 VSUBS 3.72f
C1305 M.n1175 VSUBS 1.11f
C1306 M.t17 VSUBS 3.72f
C1307 M.n1176 VSUBS 1.11f
C1308 M.t128 VSUBS 3.72f
C1309 M.n1177 VSUBS 1.11f
C1310 M.t81 VSUBS 3.72f
C1311 M.n1178 VSUBS 1.11f
C1312 M.t47 VSUBS 3.72f
C1313 M.n1179 VSUBS 1.11f
C1314 M.t127 VSUBS 3.72f
C1315 M.n1180 VSUBS 1.11f
C1316 M.t5 VSUBS 3.72f
C1317 M.n1181 VSUBS 1.11f
C1318 M.t111 VSUBS 3.72f
C1319 M.n1182 VSUBS 1.11f
C1320 M.t57 VSUBS 3.72f
C1321 M.n1183 VSUBS 0.847f
C1322 M.n1184 VSUBS 0.0593f
C1323 M.n1185 VSUBS 0.0107f
C1324 M.n1186 VSUBS 0.00593f
C1325 M.n1187 VSUBS 0.00682f
C1326 M.n1188 VSUBS 0.0104f
C1327 M.n1189 VSUBS 0.00593f
C1328 M.n1190 VSUBS 0.0267f
C1329 M.n1191 VSUBS 0.522f
C1330 M.n1192 VSUBS 0.00949f
C1331 M.n1193 VSUBS 0.0119f
C1332 M.n1194 VSUBS 0.00504f
C1333 M.n1195 VSUBS 0.0086f
C1334 M.n1196 VSUBS 0.00979f
C1335 M.n1197 VSUBS 0.00504f
C1336 M.n1198 VSUBS 0.0086f
C1337 M.n1199 VSUBS 0.0116f
C1338 M.n1200 VSUBS 0.046f
C1339 M.n1201 VSUBS 0.0528f
C1340 M.n1202 VSUBS 0.0373f
C1341 M.n1203 VSUBS 0.0116f
C1342 M.n1204 VSUBS 0.00204f
C1343 M.n1205 VSUBS 0.0096f
C1344 M.n1206 VSUBS 0.0096f
C1345 M.n1207 VSUBS 0.00175f
C1346 M.n1208 VSUBS 0.0116f
C1347 M.n1209 VSUBS 0.0116f
C1348 M.n1210 VSUBS 0.0323f
C1349 M.n1211 VSUBS 0.0323f
C1350 M.n1212 VSUBS 0.0113f
C1351 M.n1213 VSUBS 0.0421f
C1352 M.n1214 VSUBS 0.00477f
C1353 M.n1215 VSUBS 0.00116f
C1354 M.n1216 VSUBS 0.00582f
C1355 M.n1217 VSUBS 0.0096f
C1356 M.n1218 VSUBS 0.00582f
C1357 M.n1219 VSUBS 0.00582f
C1358 M.n1220 VSUBS 0.00553f
C1359 M.n1221 VSUBS 0.00466f
C1360 M.n1222 VSUBS 0.00466f
C1361 M.n1223 VSUBS 0.00116f
C1362 M.n1224 VSUBS 0.00116f
C1363 M.n1225 VSUBS 0.0268f
C1364 M.n1226 VSUBS 0.0268f
C1365 M.n1227 VSUBS 0.00844f
C1366 M.n1228 VSUBS 0.00844f
C1367 M.n1229 VSUBS 0.0032f
C1368 M.n1230 VSUBS 0.00407f
C1369 M.n1231 VSUBS 0.00262f
C1370 M.n1232 VSUBS 0.00669f
C1371 M.n1233 VSUBS 0.00786f
C1372 M.n1234 VSUBS 0.00291f
C1373 M.n1235 VSUBS 0.00291f
C1374 M.n1236 VSUBS 0.00757f
C1375 M.n1237 VSUBS 0.0064f
C1376 M.n1238 VSUBS 0.00495f
C1377 M.n1239 VSUBS 0.00495f
C1378 M.n1240 VSUBS 0.041f
C1379 M.n1241 VSUBS 0.041f
C1380 M.n1242 VSUBS 0.0116f
C1381 M.n1243 VSUBS 0.0381f
C1382 M.n1244 VSUBS 0.0116f
C1383 M.n1245 VSUBS 0.00291f
C1384 M.n1246 VSUBS 0.00786f
C1385 M.n1247 VSUBS 0.00786f
C1386 M.n1248 VSUBS 0.00262f
C1387 M.n1249 VSUBS 0.0116f
C1388 M.n1250 VSUBS 0.0108f
C1389 M.n1251 VSUBS 0.0341f
C1390 M.n1252 VSUBS 0.0341f
C1391 M.n1253 VSUBS 0.0105f
C1392 M.n1254 VSUBS 0.0428f
C1393 M.n1255 VSUBS 0.00466f
C1394 M.n1256 VSUBS 0.00116f
C1395 M.n1257 VSUBS 0.00116f
C1396 M.n1258 VSUBS 0.00495f
C1397 M.n1259 VSUBS 0.00873f
C1398 M.n1260 VSUBS 0.00582f
C1399 M.n1261 VSUBS 0.00495f
C1400 M.n1262 VSUBS 0.00466f
C1401 M.n1263 VSUBS 0.00466f
C1402 M.n1264 VSUBS 0.00466f
C1403 M.n1265 VSUBS 0.00116f
C1404 M.n1266 VSUBS 0.00116f
C1405 M.n1267 VSUBS 0.0285f
C1406 M.n1268 VSUBS 0.0285f
C1407 M.n1269 VSUBS 0.00844f
C1408 M.n1270 VSUBS 0.00844f
C1409 M.n1271 VSUBS 0.00233f
C1410 M.n1272 VSUBS 0.00407f
C1411 M.n1273 VSUBS 0.00349f
C1412 M.n1274 VSUBS 0.00582f
C1413 M.n1275 VSUBS 0.00611f
C1414 M.n1276 VSUBS 0.00204f
C1415 M.n1277 VSUBS 0.00378f
C1416 M.n1278 VSUBS 0.00757f
C1417 M.n1279 VSUBS 0.00553f
C1418 M.n1280 VSUBS 0.00495f
C1419 M.n1281 VSUBS 0.00495f
C1420 M.n1282 VSUBS 0.0428f
C1421 M.n1283 VSUBS 0.0428f
C1422 M.n1284 VSUBS 0.0108f
C1423 M.n1285 VSUBS 0.0508f
C1424 M.n1286 VSUBS 0.0099f
C1425 M.n1287 VSUBS 0.0096f
C1426 M.n1288 VSUBS 0.0125f
C1427 M.n1289 VSUBS 0.0448f
C1428 M.n1290 VSUBS 0.0445f
C1429 M.n1291 VSUBS 0.0495f
C1430 M.n1292 VSUBS 0.00524f
C1431 M.n1293 VSUBS 0.00879f
C1432 M.n1294 VSUBS 0.119f
C1433 M.n1295 VSUBS 3.22e-20
C1434 M.n1296 VSUBS 0.00582f
C1435 M.n1297 VSUBS 0.00495f
C1436 M.n1298 VSUBS 0.00844f
C1437 M.n1299 VSUBS 0.00582f
C1438 M.n1300 VSUBS 0.0306f
C1439 M.n1301 VSUBS 0.0378f
C1440 M.n1302 VSUBS 0.00989f
C1441 M.n1303 VSUBS 0.00495f
C1442 M.n1304 VSUBS 0.00844f
C1443 M.n1305 VSUBS 0.00611f
C1444 M.n1306 VSUBS 0.00495f
C1445 M.n1307 VSUBS 0.00844f
C1446 M.n1308 VSUBS 0.0096f
C1447 M.n1309 VSUBS 0.0486f
C1448 M.n1310 VSUBS 0.0536f
C1449 M.n1311 VSUBS 0.127f
C1450 M.n1312 VSUBS 0.0573f
C1451 M.n1313 VSUBS 0.0134f
C1452 M.n1314 VSUBS 0.0681f
C1453 M.n1315 VSUBS 0.118f
C1454 M.n1316 VSUBS 0.0195f
C1455 M.n1317 VSUBS 0.0195f
C1456 M.n1318 VSUBS 0.0212f
C1457 M.n1319 VSUBS 0.0234f
C1458 M.n1320 VSUBS 0.0436f
C1459 M.n1321 VSUBS 0.0439f
C1460 M.n1322 VSUBS 0.0128f
C1461 M.n1323 VSUBS 0.0116f
C1462 M.n1324 VSUBS 0.0119f
C1463 M.n1325 VSUBS 0.0128f
C1464 M.n1326 VSUBS 1.26f
C1465 M.n1327 VSUBS 1.27f
C1466 M.n1328 VSUBS 0.0399f
C1467 M.n1329 VSUBS 0.0114f
C1468 M.n1330 VSUBS 0.0417f
C1469 M.n1331 VSUBS 0.0105f
C1470 M.n1332 VSUBS 0.0259f
C1471 M.n1333 VSUBS 0.0067f
C1472 M.n1334 VSUBS 0.00845f
C1473 M.n1335 VSUBS 0.00408f
C1474 M.n1336 VSUBS 0.0067f
C1475 M.n1337 VSUBS 0.0455f
C1476 M.n1338 VSUBS 0.0067f
C1477 M.n1339 VSUBS 0.194f
C1478 M.n1340 VSUBS 0.00874f
C1479 M.n1341 VSUBS 0.00437f
C1480 M.n1342 VSUBS 0.0067f
C1481 M.n1343 VSUBS 0.0481f
C1482 M.n1344 VSUBS 0.0522f
C1483 M.n1345 VSUBS 0.077f
C1484 M.n1346 VSUBS 0.056f
C1485 M.n1347 VSUBS 0.0195f
C1486 M.n1348 VSUBS 0.0551f
C1487 M.n1349 VSUBS 0.0213f
C1488 M.n1350 VSUBS 0.023f
C1489 M.n1351 VSUBS 0.0504f
C1490 M.n1352 VSUBS 0.0446f
C1491 M.n1353 VSUBS 0.0067f
C1492 M.n1354 VSUBS 0.00612f
C1493 M.n1355 VSUBS 0.0399f
C1494 M.n1356 VSUBS 0.00554f
C1495 M.n1357 VSUBS 0.00554f
C1496 M.n1358 VSUBS 0.00117f
C1497 M.n1359 VSUBS 0.00117f
C1498 M.n1360 VSUBS 0.00495f
C1499 M.n1361 VSUBS 0.0417f
C1500 M.n1362 VSUBS 0.00554f
C1501 M.n1363 VSUBS 0.00554f
C1502 M.n1364 VSUBS 0.00117f
C1503 M.n1365 VSUBS 0.00117f
C1504 M.n1366 VSUBS 0.00408f
C1505 M.n1367 VSUBS 0.00874f
C1506 M.n1368 VSUBS 0.00962f
C1507 M.n1369 VSUBS 0.0105f
C1508 M.n1370 VSUBS 0.0067f
C1509 M.n1371 VSUBS 0.0067f
C1510 M.n1372 VSUBS 0.0067f
C1511 M.n1373 VSUBS 0.0222f
C1512 M.n1374 VSUBS 0.00117f
C1513 M.n1375 VSUBS 0.00117f
C1514 M.n1376 VSUBS 0.00554f
C1515 M.n1377 VSUBS 0.00554f
C1516 M.n1378 VSUBS 0.00466f
C1517 M.n1379 VSUBS 0.0239f
C1518 M.n1380 VSUBS 0.00117f
C1519 M.n1381 VSUBS 0.00117f
C1520 M.n1382 VSUBS 0.00554f
C1521 M.n1383 VSUBS 0.00554f
C1522 M.n1384 VSUBS 0.00379f
C1523 M.n1385 VSUBS 0.00408f
C1524 M.n1386 VSUBS 0.00495f
C1525 M.n1387 VSUBS 0.00583f
C1526 M.n1388 VSUBS 0.0102f
C1527 M.n1389 VSUBS 0.0067f
C1528 M.n1390 VSUBS 0.0224f
C1529 M.n1391 VSUBS 0.0277f
C1530 M.n1392 VSUBS 0.494f
C1531 M.n1393 VSUBS 0.00845f
C1532 M.n1394 VSUBS 0.00204f
C1533 M.n1395 VSUBS 0.00758f
C1534 M.n1396 VSUBS 0.00291f
C1535 M.n1397 VSUBS 0.0239f
C1536 M.n1398 VSUBS 0.0108f
C1537 M.n1399 VSUBS 0.0119f
C1538 M.n1400 VSUBS 0.0222f
C1539 M.n1401 VSUBS 0.0117f
C1540 M.n1402 VSUBS 0.0119f
C1541 M.n1403 VSUBS 0.00641f
C1542 M.n1404 VSUBS 0.00962f
C1543 M.n1405 VSUBS 0.0102f
C1544 M.n1406 VSUBS 0.00321f
C1545 M.n1407 VSUBS 0.00758f
C1546 M.n1408 VSUBS 0.00175f
C1547 M.n1409 VSUBS 0.00233f
C1548 M.n1410 VSUBS 0.00991f
C1549 M.n1411 VSUBS 0.00845f
C1550 M.n1412 VSUBS 0.00175f
C1551 M.n1413 VSUBS 0.00233f
C1552 M.n1414 VSUBS 0.00991f
C1553 M.n1415 VSUBS 0.00991f
C1554 M.n1416 VSUBS 0.0154f
C1555 M.n1417 VSUBS 0.00845f
C1556 M.n1418 VSUBS 0.00845f
C1557 M.n1419 VSUBS 0.00291f
C1558 M.n1420 VSUBS 0.0172f
C1559 M.n1421 VSUBS 0.00845f
C1560 M.n1422 VSUBS 0.00845f
C1561 M.n1423 VSUBS 0.00204f
C1562 M.n1424 VSUBS 0.00962f
C1563 M.n1425 VSUBS 0.0105f
C1564 M.n1426 VSUBS 0.0114f
C1565 M.n1427 VSUBS 0.0114f
C1566 M.n1428 VSUBS 0.023f
C1567 M.n1429 VSUBS 0.0262f
C1568 M.n1430 VSUBS 0.0154f
C1569 M.n1431 VSUBS 0.0117f
C1570 M.n1432 VSUBS 0.0172f
C1571 M.n1433 VSUBS 0.0108f
C1572 M.n1434 VSUBS 0.0166f
C1573 M.n1435 VSUBS 0.0166f
C1574 M.n1436 VSUBS 0.0175f
C1575 M.n1437 VSUBS 0.0114f
C1576 M.n1438 VSUBS 0.0117f
C1577 M.n1439 VSUBS 0.00758f
C1578 M.n1440 VSUBS 0.00291f
C1579 M.n1441 VSUBS 0.00291f
C1580 M.n1442 VSUBS 0.00787f
C1581 M.n1443 VSUBS 0.0163f
C1582 M.n1444 VSUBS 0.0067f
C1583 M.n1445 VSUBS 0.00466f
C1584 M.n1446 VSUBS 0.00466f
C1585 M.n1447 VSUBS 0.00699f
C1586 M.n1448 VSUBS 0.0146f
C1587 M.n1449 VSUBS 0.0146f
C1588 M.n1450 VSUBS 0.0114f
C1589 M.n1451 VSUBS 0.0117f
C1590 M.n1452 VSUBS 0.0198f
C1591 M.n1453 VSUBS 0.0114f
C1592 M.n1454 VSUBS 0.0216f
C1593 M.n1455 VSUBS 0.0105f
C1594 M.n1456 VSUBS 0.00962f
C1595 M.n1457 VSUBS 8.74e-19
C1596 M.n1458 VSUBS 8.74e-19
C1597 M.n1459 VSUBS 0.00991f
C1598 M.n1460 VSUBS 0.0192f
C1599 M.n1461 VSUBS 0.00933f
C1600 M.n1462 VSUBS 0.00204f
C1601 M.n1463 VSUBS 0.00204f
C1602 M.n1464 VSUBS 0.00962f
C1603 M.n1465 VSUBS 0.0192f
C1604 M.n1466 VSUBS 0.0201f
C1605 M.n1467 VSUBS 0.0303f
C1606 M.n1468 VSUBS 0.0306f
C1607 M.n1469 VSUBS 0.0362f
C1608 M.n1470 VSUBS 0.15f
C1609 M.n1471 VSUBS 0.0376f
C1610 M.n1472 VSUBS 0.0551f
C1611 M.n1473 VSUBS 0.0461f
C1612 M.n1474 VSUBS 0.0571f
C1613 M.n1475 VSUBS 0.0347f
C1614 M.n1476 VSUBS 0.0128f
C1615 M.n1477 VSUBS 0.00962f
C1616 M.n1478 VSUBS 0.00845f
C1617 M.n1479 VSUBS 0.00321f
C1618 M.n1480 VSUBS 0.0213f
C1619 M.n1481 VSUBS 0.00991f
C1620 M.n1482 VSUBS 0.00962f
C1621 M.n1483 VSUBS 0.00962f
C1622 M.n1484 VSUBS 0.0265f
C1623 M.n1485 VSUBS 0.028f
C1624 M.n1486 VSUBS 0.0175f
C1625 M.n1487 VSUBS 0.00962f
C1626 M.n1488 VSUBS 0.00991f
C1627 M.n1489 VSUBS 0.0175f
C1628 M.n1490 VSUBS 0.0102f
C1629 M.n1491 VSUBS 0.0105f
C1630 M.n1492 VSUBS 0.0195f
C1631 M.n1493 VSUBS 0.0321f
C1632 M.n1494 VSUBS 0.0324f
C1633 M.n1495 VSUBS 0.0572f
C1634 M.n1496 VSUBS 0.037f
C1635 M.n1497 VSUBS 0.0216f
C1636 M.n1498 VSUBS 0.0108f
C1637 M.n1499 VSUBS 0.0195f
C1638 M.n1500 VSUBS 0.0198f
C1639 M.n1501 VSUBS 0.0117f
C1640 M.n1502 VSUBS 0.0213f
C1641 M.n1503 VSUBS 0.023f
C1642 M.n1504 VSUBS 1.31f
C1643 M.n1505 VSUBS 1.34f
C1644 M.n1506 VSUBS 0.00177f
C1645 M.n1507 VSUBS 0.00253f
C1646 M.n1508 VSUBS 0.018f
C1647 M.n1509 VSUBS 0.00836f
C1648 M.n1510 VSUBS 0.0461f
C1649 M.n1511 VSUBS 0.00861f
C1650 M.n1512 VSUBS 0.00861f
C1651 M.n1513 VSUBS 0.0291f
C1652 M.n1514 VSUBS 0.0289f
C1653 M.n1515 VSUBS 0.00836f
C1654 M.n1516 VSUBS 0.0459f
C1655 M.n1517 VSUBS 0.00836f
C1656 M.n1518 VSUBS 0.155f
C1657 M.n1519 VSUBS 0.00684f
C1658 M.n1520 VSUBS 0.00456f
C1659 M.n1521 VSUBS 0.00583f
C1660 M.n1522 VSUBS 0.00659f
C1661 M.n1523 VSUBS 0.132f
C1662 M.n1524 VSUBS 0.121f
C1663 M.n1525 VSUBS 0.0104f
C1664 M.n1526 VSUBS 0.12f
C1665 M.n1527 VSUBS 0.0104f
C1666 M.n1528 VSUBS 0.0119f
C1667 M.n1529 VSUBS 0.00539f
C1668 M.n1530 VSUBS 0.00943f
C1669 M.n1531 VSUBS 0.00647f
C1670 M.n1532 VSUBS 0.00405f
C1671 M.n1533 VSUBS 0.00405f
C1672 M.n1534 VSUBS 0.00253f
C1673 M.n1535 VSUBS 0.00253f
C1674 M.n1536 VSUBS 0.00279f
C1675 M.n1537 VSUBS 0.00608f
C1676 M.n1538 VSUBS 0.00405f
C1677 M.n1539 VSUBS 0.00405f
C1678 M.n1540 VSUBS 0.00405f
C1679 M.n1541 VSUBS 0.00405f
C1680 M.n1542 VSUBS 0.00203f
C1681 M.n1543 VSUBS 0.00532f
C1682 M.n1544 VSUBS 0.00566f
C1683 M.n1545 VSUBS 0.0225f
C1684 M.n1546 VSUBS 0.00405f
C1685 M.n1547 VSUBS 0.00405f
C1686 M.n1548 VSUBS 0.00583f
C1687 M.n1549 VSUBS 0.0241f
C1688 M.n1550 VSUBS 0.00405f
C1689 M.n1551 VSUBS 0.00405f
C1690 M.n1552 VSUBS 0.00507f
C1691 M.n1553 VSUBS 0.00836f
C1692 M.n1554 VSUBS 0.00912f
C1693 M.n1555 VSUBS 0.0105f
C1694 M.n1556 VSUBS 0.0105f
C1695 M.n1557 VSUBS 0.0275f
C1696 M.n1558 VSUBS 0.0278f
C1697 M.n1559 VSUBS 0.0108f
C1698 M.n1560 VSUBS 0.0225f
C1699 M.n1561 VSUBS 0.00431f
C1700 M.n1562 VSUBS 0.00431f
C1701 M.n1563 VSUBS 0.00583f
C1702 M.n1564 VSUBS 0.0241f
C1703 M.n1565 VSUBS 0.00431f
C1704 M.n1566 VSUBS 0.00431f
C1705 M.n1567 VSUBS 0.00507f
C1706 M.n1568 VSUBS 0.00861f
C1707 M.n1569 VSUBS 0.00937f
C1708 M.n1570 VSUBS 0.00674f
C1709 M.n1571 VSUBS 0.495f
C1710 M.n1572 VSUBS 0.00431f
C1711 M.n1573 VSUBS 0.00127f
C1712 M.n1574 VSUBS 0.00127f
C1713 M.n1575 VSUBS 0.00431f
C1714 M.n1576 VSUBS 7.6e-19
C1715 M.n1577 VSUBS 0.00431f
C1716 M.n1578 VSUBS 0.00836f
C1717 M.n1579 VSUBS 0.00785f
C1718 M.n1580 VSUBS 0.00781f
C1719 M.n1581 VSUBS 0.00593f
C1720 M.n1582 VSUBS 0.00674f
C1721 M.n1583 VSUBS 0.00862f
C1722 M.n1584 VSUBS 0.0144f
C1723 M.n1585 VSUBS 0.00988f
C1724 M.n1586 VSUBS 0.016f
C1725 M.n1587 VSUBS 0.00912f
C1726 M.n1588 VSUBS 7.6e-19
C1727 M.n1589 VSUBS 0.00355f
C1728 M.n1590 VSUBS 0.00405f
C1729 M.n1591 VSUBS 0.00532f
C1730 M.n1592 VSUBS 0.0129f
C1731 M.n1593 VSUBS 0.00431f
C1732 M.n1594 VSUBS 0.00456f
C1733 M.n1595 VSUBS 0.0129f
C1734 M.n1596 VSUBS 0.0145f
C1735 M.n1597 VSUBS 0.0251f
C1736 M.n1598 VSUBS 0.0181f
C1737 M.n1599 VSUBS 0.0108f
C1738 M.n1600 VSUBS 0.016f
C1739 M.n1601 VSUBS 0.00329f
C1740 M.n1602 VSUBS 0.00329f
C1741 M.n1603 VSUBS 0.00608f
C1742 M.n1604 VSUBS 0.00861f
C1743 M.n1605 VSUBS 0.0144f
C1744 M.n1606 VSUBS 0.00329f
C1745 M.n1607 VSUBS 0.00329f
C1746 M.n1608 VSUBS 0.00684f
C1747 M.n1609 VSUBS 0.00937f
C1748 M.n1610 VSUBS 0.0108f
C1749 M.n1611 VSUBS 0.00963f
C1750 M.n1612 VSUBS 0.00329f
C1751 M.n1613 VSUBS 0.00329f
C1752 M.n1614 VSUBS 0.00659f
C1753 M.n1615 VSUBS 0.0111f
C1754 M.n1616 VSUBS 0.00329f
C1755 M.n1617 VSUBS 0.00329f
C1756 M.n1618 VSUBS 0.00583f
C1757 M.n1619 VSUBS 0.00836f
C1758 M.n1620 VSUBS 0.00912f
C1759 M.n1621 VSUBS 0.0105f
C1760 M.n1622 VSUBS 0.0105f
C1761 M.n1623 VSUBS 0.0129f
C1762 M.n1624 VSUBS 0.0202f
C1763 M.n1625 VSUBS 0.0289f
C1764 M.n1626 VSUBS 0.00988f
C1765 M.n1627 VSUBS 0.00963f
C1766 M.n1628 VSUBS 0.0101f
C1767 M.n1629 VSUBS 0.0304f
C1768 M.n1630 VSUBS 0.00912f
C1769 M.n1631 VSUBS 0.0111f
C1770 M.n1632 VSUBS 0.00937f
C1771 M.n1633 VSUBS 0.017f
C1772 M.n1634 VSUBS 0.0185f
C1773 M.n1635 VSUBS 0.0213f
C1774 M.n1636 VSUBS 0.0404f
C1775 M.n1637 VSUBS 0.0407f
C1776 M.n1638 VSUBS 0.0964f
C1777 M.n1639 VSUBS 0.229f
C1778 M.n1640 VSUBS 0.0322f
C1779 M.n1641 VSUBS 0.037f
C1780 M.n1642 VSUBS 0.0474f
C1781 M.n1643 VSUBS 0.00507f
C1782 M.n1644 VSUBS 0.00431f
C1783 M.n1645 VSUBS 0.00861f
C1784 M.n1646 VSUBS 0.0137f
C1785 M.n1647 VSUBS 0.0251f
C1786 M.n1648 VSUBS 0.02f
C1787 M.n1649 VSUBS 0.00861f
C1788 M.n1650 VSUBS 0.00861f
C1789 M.n1651 VSUBS 0.00836f
C1790 M.n1652 VSUBS 0.00836f
C1791 M.n1653 VSUBS 0.0152f
C1792 M.n1654 VSUBS 0.0205f
C1793 M.n1655 VSUBS 0.017f
C1794 M.n1656 VSUBS 0.0395f
C1795 M.n1657 VSUBS 0.0398f
C1796 M.n1658 VSUBS 0.116f
C1797 M.n1659 VSUBS 0.097f
C1798 M.n1660 VSUBS 0.0304f
C1799 M.n1661 VSUBS 0.00937f
C1800 M.n1662 VSUBS 0.017f
C1801 M.n1663 VSUBS 0.0289f
C1802 M.n1664 VSUBS 0.0101f
C1803 M.n1665 VSUBS 0.0185f
C1804 M.n1666 VSUBS 0.0213f
C1805 M.n1667 VSUBS 1.3f
C1806 M.n1668 VSUBS 1.29f
C1807 M.n1669 VSUBS 0.0276f
C1808 M.n1670 VSUBS 0.00988f
C1809 M.n1671 VSUBS 0.0291f
C1810 M.n1672 VSUBS 0.00912f
C1811 M.n1673 VSUBS 0.0383f
C1812 M.n1674 VSUBS 0.0909f
C1813 M.n1675 VSUBS 0.0725f
C1814 M.n1676 VSUBS 0.017f
C1815 M.n1677 VSUBS 0.0718f
C1816 M.n1678 VSUBS 0.0185f
C1817 M.n1679 VSUBS 0.0208f
C1818 M.n1680 VSUBS 0.0381f
C1819 M.n1681 VSUBS 0.0284f
C1820 M.n1682 VSUBS 0.00395f
C1821 M.n1683 VSUBS 0.01f
C1822 M.n1684 VSUBS 0.0289f
C1823 M.n1685 VSUBS 7.6e-19
C1824 M.n1686 VSUBS 7.6e-19
C1825 M.n1687 VSUBS 0.00304f
C1826 M.n1688 VSUBS 0.00329f
C1827 M.n1689 VSUBS 0.00557f
C1828 M.n1690 VSUBS 0.00532f
C1829 M.n1691 VSUBS 0.0274f
C1830 M.n1692 VSUBS 7.6e-19
C1831 M.n1693 VSUBS 7.6e-19
C1832 M.n1694 VSUBS 0.00304f
C1833 M.n1695 VSUBS 0.00329f
C1834 M.n1696 VSUBS 0.00633f
C1835 M.n1697 VSUBS 0.00608f
C1836 M.n1698 VSUBS 0.0071f
C1837 M.n1699 VSUBS 0.0038f
C1838 M.n1700 VSUBS 0.0038f
C1839 M.n1701 VSUBS 0.00395f
C1840 M.n1702 VSUBS 0.00973f
C1841 M.n1703 VSUBS 0.00684f
C1842 M.n1704 VSUBS 0.00395f
C1843 M.n1705 VSUBS 0.0263f
C1844 M.n1706 VSUBS 0.0318f
C1845 M.n1707 VSUBS 0.0105f
C1846 M.n1708 VSUBS 0.0228f
C1847 M.n1709 VSUBS 0.00861f
C1848 M.n1710 VSUBS 0.00861f
C1849 M.n1711 VSUBS 0.00152f
C1850 M.n1712 VSUBS 0.0507f
C1851 M.n1713 VSUBS 0.0453f
C1852 M.n1714 VSUBS 0.174f
C1853 M.n1715 VSUBS 0.0038f
C1854 M.n1716 VSUBS 0.0304f
C1855 M.n1717 VSUBS 0.0038f
C1856 M.n1718 VSUBS 0.00811f
C1857 M.n1719 VSUBS 0.00532f
C1858 M.n1720 VSUBS 0.0038f
C1859 M.n1721 VSUBS 0.00785f
C1860 M.n1722 VSUBS 0.00507f
C1861 M.n1723 VSUBS 0.0038f
C1862 M.n1724 VSUBS 0.0284f
C1863 M.n1725 VSUBS 0.0337f
C1864 M.n1726 VSUBS 0.017f
C1865 M.n1727 VSUBS 0.0243f
C1866 M.n1728 VSUBS 0.00861f
C1867 M.n1729 VSUBS 0.00861f
C1868 M.n1730 VSUBS 0.00836f
C1869 M.n1731 VSUBS 0.0076f
C1870 M.n1732 VSUBS 0.00395f
C1871 M.n1733 VSUBS 0.496f
C1872 M.n1734 VSUBS 0.00658f
C1873 M.n1735 VSUBS 0.00785f
C1874 M.n1736 VSUBS 0.00127f
C1875 M.n1737 VSUBS 0.00836f
C1876 M.n1738 VSUBS 0.00836f
C1877 M.n1739 VSUBS 0.00101f
C1878 M.n1740 VSUBS 7.6e-19
C1879 M.n1741 VSUBS 0.0076f
C1880 M.n1742 VSUBS 0.00177f
C1881 M.n1743 VSUBS 0.00152f
C1882 M.n1744 VSUBS 0.00316f
C1883 M.n1745 VSUBS 0.00868f
C1884 M.n1746 VSUBS 0.0144f
C1885 M.n1747 VSUBS 0.00836f
C1886 M.n1748 VSUBS 0.00836f
C1887 M.n1749 VSUBS 0.00152f
C1888 M.n1750 VSUBS 0.016f
C1889 M.n1751 VSUBS 0.00836f
C1890 M.n1752 VSUBS 0.00836f
C1891 M.n1753 VSUBS 0.0253f
C1892 M.n1754 VSUBS 0.0251f
C1893 M.n1755 VSUBS 0.00861f
C1894 M.n1756 VSUBS 0.00861f
C1895 M.n1757 VSUBS 0.017f
C1896 M.n1758 VSUBS 0.0421f
C1897 M.n1759 VSUBS 0.0167f
C1898 M.n1760 VSUBS 0.00861f
C1899 M.n1761 VSUBS 0.00785f
C1900 M.n1762 VSUBS 0.00894f
C1901 M.n1763 VSUBS 0.0103f
C1902 M.n1764 VSUBS 0.0229f
C1903 M.n1765 VSUBS 0.0247f
C1904 M.n1766 VSUBS 0.016f
C1905 M.n1767 VSUBS 0.00937f
C1906 M.n1768 VSUBS 0.0147f
C1907 M.n1769 VSUBS 0.0144f
C1908 M.n1770 VSUBS 0.0101f
C1909 M.n1771 VSUBS 0.0147f
C1910 M.n1772 VSUBS 0.016f
C1911 M.n1773 VSUBS 0.0103f
C1912 M.n1774 VSUBS 0.0105f
C1913 M.n1775 VSUBS 0.00557f
C1914 M.n1776 VSUBS 0.00431f
C1915 M.n1777 VSUBS 0.00608f
C1916 M.n1778 VSUBS 0.0038f
C1917 M.n1779 VSUBS 0.0038f
C1918 M.n1780 VSUBS 0.00633f
C1919 M.n1781 VSUBS 0.00507f
C1920 M.n1782 VSUBS 0.00684f
C1921 M.n1783 VSUBS 0.00228f
C1922 M.n1784 VSUBS 0.00228f
C1923 M.n1785 VSUBS 0.00709f
C1924 M.n1786 VSUBS 0.0106f
C1925 M.n1787 VSUBS 0.00912f
C1926 M.n1788 VSUBS 0.00947f
C1927 M.n1789 VSUBS 0.0103f
C1928 M.n1790 VSUBS 0.0105f
C1929 M.n1791 VSUBS 0.0167f
C1930 M.n1792 VSUBS 0.00988f
C1931 M.n1793 VSUBS 0.00557f
C1932 M.n1794 VSUBS 0.00456f
C1933 M.n1795 VSUBS 0.0182f
C1934 M.n1796 VSUBS 0.00912f
C1935 M.n1797 VSUBS 0.00405f
C1936 M.n1798 VSUBS 0.00405f
C1937 M.n1799 VSUBS 0.00532f
C1938 M.n1800 VSUBS 0.0129f
C1939 M.n1801 VSUBS 0.0129f
C1940 M.n1802 VSUBS 0.0142f
C1941 M.n1803 VSUBS 0.0268f
C1942 M.n1804 VSUBS 0.0271f
C1943 M.n1805 VSUBS 0.106f
C1944 M.n1806 VSUBS 0.199f
C1945 M.n1807 VSUBS 0.0291f
C1946 M.n1808 VSUBS 0.0491f
C1947 M.n1809 VSUBS 0.0155f
C1948 M.n1810 VSUBS 0.00836f
C1949 M.n1811 VSUBS 0.00861f
C1950 M.n1812 VSUBS 0.0122f
C1951 M.n1813 VSUBS 0.00836f
C1952 M.n1814 VSUBS 0.00861f
C1953 M.n1815 VSUBS 0.0137f
C1954 M.n1816 VSUBS 0.0274f
C1955 M.n1817 VSUBS 0.0276f
C1956 M.n1818 VSUBS 0.124f
C1957 M.n1819 VSUBS 0.106f
C1958 M.n1820 VSUBS 0.0182f
C1959 M.n1821 VSUBS 0.00937f
C1960 M.n1822 VSUBS 0.017f
C1961 M.n1823 VSUBS 0.0167f
C1962 M.n1824 VSUBS 0.0101f
C1963 M.n1825 VSUBS 0.0185f
C1964 M.n1826 VSUBS 0.0208f
C1965 M.n1827 VSUBS 1.28f
C1966 M.n1828 VSUBS 1.26f
C1967 M.n1829 VSUBS 0.041f
C1968 M.n1830 VSUBS 0.00988f
C1969 M.n1831 VSUBS 0.0426f
C1970 M.n1832 VSUBS 0.00912f
C1971 M.n1833 VSUBS 0.0289f
C1972 M.n1834 VSUBS 0.00532f
C1973 M.n1835 VSUBS 0.00405f
C1974 M.n1836 VSUBS 0.00735f
C1975 M.n1837 VSUBS 0.0459f
C1976 M.n1838 VSUBS 0.00532f
C1977 M.n1839 VSUBS 0.00532f
C1978 M.n1840 VSUBS 0.177f
C1979 M.n1841 VSUBS 0.00431f
C1980 M.n1842 VSUBS 0.0076f
C1981 M.n1843 VSUBS 0.00532f
C1982 M.n1844 VSUBS 0.0443f
C1983 M.n1845 VSUBS 0.0517f
C1984 M.n1846 VSUBS 0.0674f
C1985 M.n1847 VSUBS 0.0486f
C1986 M.n1848 VSUBS 0.017f
C1987 M.n1849 VSUBS 0.048f
C1988 M.n1850 VSUBS 0.0185f
C1989 M.n1851 VSUBS 0.02f
C1990 M.n1852 VSUBS 0.0502f
C1991 M.n1853 VSUBS 0.0413f
C1992 M.n1854 VSUBS 0.00532f
C1993 M.n1855 VSUBS 0.00912f
C1994 M.n1856 VSUBS 0.0426f
C1995 M.n1857 VSUBS 0.00101f
C1996 M.n1858 VSUBS 0.00101f
C1997 M.n1859 VSUBS 0.00431f
C1998 M.n1860 VSUBS 0.00431f
C1999 M.n1861 VSUBS 0.00405f
C2000 M.n1862 VSUBS 0.00431f
C2001 M.n1863 VSUBS 0.041f
C2002 M.n1864 VSUBS 0.00101f
C2003 M.n1865 VSUBS 0.00101f
C2004 M.n1866 VSUBS 0.00431f
C2005 M.n1867 VSUBS 0.00431f
C2006 M.n1868 VSUBS 0.00481f
C2007 M.n1869 VSUBS 0.00507f
C2008 M.n1870 VSUBS 0.00583f
C2009 M.n1871 VSUBS 0.00532f
C2010 M.n1872 VSUBS 0.00532f
C2011 M.n1873 VSUBS 0.00532f
C2012 M.n1874 VSUBS 0.0223f
C2013 M.n1875 VSUBS 0.00431f
C2014 M.n1876 VSUBS 0.00431f
C2015 M.n1877 VSUBS 0.00101f
C2016 M.n1878 VSUBS 0.00101f
C2017 M.n1879 VSUBS 0.00456f
C2018 M.n1880 VSUBS 0.0238f
C2019 M.n1881 VSUBS 0.00431f
C2020 M.n1882 VSUBS 0.00431f
C2021 M.n1883 VSUBS 0.00101f
C2022 M.n1884 VSUBS 0.00101f
C2023 M.n1885 VSUBS 0.0038f
C2024 M.n1886 VSUBS 0.00735f
C2025 M.n1887 VSUBS 0.00811f
C2026 M.n1888 VSUBS 0.00887f
C2027 M.n1889 VSUBS 0.00557f
C2028 M.n1890 VSUBS 0.00532f
C2029 M.n1891 VSUBS 0.0258f
C2030 M.n1892 VSUBS 0.0304f
C2031 M.n1893 VSUBS 0.511f
C2032 M.n1894 VSUBS 0.00431f
C2033 M.n1895 VSUBS 0.00329f
C2034 M.n1896 VSUBS 0.0223f
C2035 M.n1897 VSUBS 0.0101f
C2036 M.n1898 VSUBS 0.00431f
C2037 M.n1899 VSUBS 0.00405f
C2038 M.n1900 VSUBS 0.0238f
C2039 M.n1901 VSUBS 0.00937f
C2040 M.n1902 VSUBS 0.0119f
C2041 M.n1903 VSUBS 0.0119f
C2042 M.n1904 VSUBS 0.0038f
C2043 M.n1905 VSUBS 0.00684f
C2044 M.n1906 VSUBS 0.00735f
C2045 M.n1907 VSUBS 0.00583f
C2046 M.n1908 VSUBS 0.00431f
C2047 M.n1909 VSUBS 0.00228f
C2048 M.n1910 VSUBS 0.00228f
C2049 M.n1911 VSUBS 0.00355f
C2050 M.n1912 VSUBS 0.00431f
C2051 M.n1913 VSUBS 0.00152f
C2052 M.n1914 VSUBS 0.00431f
C2053 M.n1915 VSUBS 0.00785f
C2054 M.n1916 VSUBS 0.00709f
C2055 M.n1917 VSUBS 0.00709f
C2056 M.n1918 VSUBS 0.00431f
C2057 M.n1919 VSUBS 0.00431f
C2058 M.n1920 VSUBS 0.00557f
C2059 M.n1921 VSUBS 0.00963f
C2060 M.n1922 VSUBS 0.00431f
C2061 M.n1923 VSUBS 0.00431f
C2062 M.n1924 VSUBS 0.00481f
C2063 M.n1925 VSUBS 0.00836f
C2064 M.n1926 VSUBS 0.00912f
C2065 M.n1927 VSUBS 0.00988f
C2066 M.n1928 VSUBS 0.00988f
C2067 M.n1929 VSUBS 0.0117f
C2068 M.n1930 VSUBS 0.0175f
C2069 M.n1931 VSUBS 0.00811f
C2070 M.n1932 VSUBS 0.00811f
C2071 M.n1933 VSUBS 0.0101f
C2072 M.n1934 VSUBS 0.0114f
C2073 M.n1935 VSUBS 0.00912f
C2074 M.n1936 VSUBS 0.00963f
C2075 M.n1937 VSUBS 0.00937f
C2076 M.n1938 VSUBS 0.017f
C2077 M.n1939 VSUBS 0.0185f
C2078 M.n1940 VSUBS 0.02f
C2079 M.n1941 VSUBS 0.019f
C2080 M.n1942 VSUBS 0.0193f
C2081 M.n1943 VSUBS 0.00912f
C2082 M.n1944 VSUBS 0.0114f
C2083 M.n1945 VSUBS 0.00937f
C2084 M.n1946 VSUBS 0.017f
C2085 M.n1947 VSUBS 0.00988f
C2086 M.n1948 VSUBS 0.00988f
C2087 M.n1949 VSUBS 0.00988f
C2088 M.n1950 VSUBS 0.0101f
C2089 M.n1951 VSUBS 0.0185f
C2090 M.n1952 VSUBS 0.02f
C2091 M.n1953 VSUBS 0.0167f
C2092 M.n1954 VSUBS 0.017f
C2093 M.n1955 VSUBS 0.0205f
C2094 M.n1956 VSUBS 0.00988f
C2095 M.n1957 VSUBS 0.00988f
C2096 M.n1958 VSUBS 0.0076f
C2097 M.n1959 VSUBS 0.0076f
C2098 M.n1960 VSUBS 0.0101f
C2099 M.n1961 VSUBS 0.022f
C2100 M.n1962 VSUBS 0.00912f
C2101 M.n1963 VSUBS 0.00912f
C2102 M.n1964 VSUBS 0.00912f
C2103 M.n1965 VSUBS 0.00937f
C2104 M.n1966 VSUBS 0.017f
C2105 M.n1967 VSUBS 0.0185f
C2106 M.n1968 VSUBS 0.02f
C2107 M.n1969 VSUBS 0.0296f
C2108 M.n1970 VSUBS 0.0299f
C2109 M.n1971 VSUBS 0.0517f
C2110 M.n1972 VSUBS 0.166f
C2111 M.n1973 VSUBS 0.056f
C2112 M.n1974 VSUBS 0.0542f
C2113 M.n1975 VSUBS 0.0332f
C2114 M.n1976 VSUBS 0.0127f
C2115 M.n1977 VSUBS 0.00836f
C2116 M.n1978 VSUBS 0.00861f
C2117 M.n1979 VSUBS 0.017f
C2118 M.n1980 VSUBS 0.00861f
C2119 M.n1981 VSUBS 0.0317f
C2120 M.n1982 VSUBS 0.00836f
C2121 M.n1983 VSUBS 0.00836f
C2122 M.n1984 VSUBS 0.0147f
C2123 M.n1985 VSUBS 0.019f
C2124 M.n1986 VSUBS 0.0565f
C2125 M.n1987 VSUBS 0.017f
C2126 M.n1988 VSUBS 0.0205f
C2127 M.n1989 VSUBS 0.0208f
C2128 M.n1990 VSUBS 0.017f
C2129 M.n1991 VSUBS 0.0182f
C2130 M.n1992 VSUBS 0.0185f
C2131 M.n1993 VSUBS 0.017f
C2132 M.n1994 VSUBS 0.0312f
C2133 M.n1995 VSUBS 0.0314f
C2134 M.n1996 VSUBS 0.0704f
C2135 M.n1997 VSUBS 0.0524f
C2136 M.n1998 VSUBS 0.022f
C2137 M.n1999 VSUBS 0.00937f
C2138 M.n2000 VSUBS 0.017f
C2139 M.n2001 VSUBS 0.0205f
C2140 M.n2002 VSUBS 0.0101f
C2141 M.n2003 VSUBS 0.0185f
C2142 M.n2004 VSUBS 0.02f
C2143 M.n2005 VSUBS 0.867f
C2144 P.t57 VSUBS 2.64f
C2145 P.t21 VSUBS 2.64f
C2146 P.t19 VSUBS 2.64f
C2147 P.t75 VSUBS 2.64f
C2148 P.t61 VSUBS 2.64f
C2149 P.t94 VSUBS 2.64f
C2150 P.t5 VSUBS 2.64f
C2151 P.t31 VSUBS 2.64f
C2152 P.t95 VSUBS 2.64f
C2153 P.t83 VSUBS 2.64f
C2154 P.t105 VSUBS 2.64f
C2155 P.t24 VSUBS 2.78f
C2156 P.n0 VSUBS 4.87f
C2157 P.n1 VSUBS 2.51f
C2158 P.n2 VSUBS 2.51f
C2159 P.n3 VSUBS 2.51f
C2160 P.n4 VSUBS 2.51f
C2161 P.n5 VSUBS 2.51f
C2162 P.n6 VSUBS 2.51f
C2163 P.n7 VSUBS 2.51f
C2164 P.n8 VSUBS 2.51f
C2165 P.n9 VSUBS 2.51f
C2166 P.n10 VSUBS 2.18f
C2167 P.t70 VSUBS 2.64f
C2168 P.t2 VSUBS 2.64f
C2169 P.t81 VSUBS 2.64f
C2170 P.t125 VSUBS 2.64f
C2171 P.t120 VSUBS 2.64f
C2172 P.t8 VSUBS 2.64f
C2173 P.t59 VSUBS 2.64f
C2174 P.t93 VSUBS 2.64f
C2175 P.t10 VSUBS 2.64f
C2176 P.t0 VSUBS 2.64f
C2177 P.t28 VSUBS 2.64f
C2178 P.t82 VSUBS 2.78f
C2179 P.n11 VSUBS 4.87f
C2180 P.n12 VSUBS 2.51f
C2181 P.n13 VSUBS 2.51f
C2182 P.n14 VSUBS 2.51f
C2183 P.n15 VSUBS 2.51f
C2184 P.n16 VSUBS 2.51f
C2185 P.n17 VSUBS 2.51f
C2186 P.n18 VSUBS 2.51f
C2187 P.n19 VSUBS 2.51f
C2188 P.n20 VSUBS 2.51f
C2189 P.n21 VSUBS 2.18f
C2190 P.t23 VSUBS 2.64f
C2191 P.t54 VSUBS 2.64f
C2192 P.t25 VSUBS 2.64f
C2193 P.t79 VSUBS 2.64f
C2194 P.t65 VSUBS 2.64f
C2195 P.t96 VSUBS 2.64f
C2196 P.t7 VSUBS 2.64f
C2197 P.t35 VSUBS 2.64f
C2198 P.t98 VSUBS 2.64f
C2199 P.t88 VSUBS 2.64f
C2200 P.t106 VSUBS 2.64f
C2201 P.t27 VSUBS 2.78f
C2202 P.n22 VSUBS 4.87f
C2203 P.n23 VSUBS 2.51f
C2204 P.n24 VSUBS 2.51f
C2205 P.n25 VSUBS 2.51f
C2206 P.n26 VSUBS 2.51f
C2207 P.n27 VSUBS 2.51f
C2208 P.n28 VSUBS 2.51f
C2209 P.n29 VSUBS 2.51f
C2210 P.n30 VSUBS 2.51f
C2211 P.n31 VSUBS 2.51f
C2212 P.n32 VSUBS 2.18f
C2213 P.t66 VSUBS 2.64f
C2214 P.t99 VSUBS 2.64f
C2215 P.t110 VSUBS 2.64f
C2216 P.t33 VSUBS 2.64f
C2217 P.t22 VSUBS 2.64f
C2218 P.t42 VSUBS 2.64f
C2219 P.t101 VSUBS 2.64f
C2220 P.t118 VSUBS 2.64f
C2221 P.t44 VSUBS 2.64f
C2222 P.t38 VSUBS 2.64f
C2223 P.t55 VSUBS 2.64f
C2224 P.t112 VSUBS 2.78f
C2225 P.n33 VSUBS 4.87f
C2226 P.n34 VSUBS 2.51f
C2227 P.n35 VSUBS 2.51f
C2228 P.n36 VSUBS 2.51f
C2229 P.n37 VSUBS 2.51f
C2230 P.n38 VSUBS 2.51f
C2231 P.n39 VSUBS 2.51f
C2232 P.n40 VSUBS 2.51f
C2233 P.n41 VSUBS 2.51f
C2234 P.n42 VSUBS 2.51f
C2235 P.n43 VSUBS 2.18f
C2236 P.t111 VSUBS 2.64f
C2237 P.t45 VSUBS 2.64f
C2238 P.t127 VSUBS 2.64f
C2239 P.t47 VSUBS 2.64f
C2240 P.t41 VSUBS 2.64f
C2241 P.t63 VSUBS 2.64f
C2242 P.t115 VSUBS 2.64f
C2243 P.t6 VSUBS 2.64f
C2244 P.t68 VSUBS 2.64f
C2245 P.t52 VSUBS 2.64f
C2246 P.t85 VSUBS 2.64f
C2247 P.t129 VSUBS 2.78f
C2248 P.n44 VSUBS 4.87f
C2249 P.n45 VSUBS 2.51f
C2250 P.n46 VSUBS 2.51f
C2251 P.n47 VSUBS 2.51f
C2252 P.n48 VSUBS 2.51f
C2253 P.n49 VSUBS 2.51f
C2254 P.n50 VSUBS 2.51f
C2255 P.n51 VSUBS 2.51f
C2256 P.n52 VSUBS 2.51f
C2257 P.n53 VSUBS 2.51f
C2258 P.n54 VSUBS 2.18f
C2259 P.n55 VSUBS 0.0021f
C2260 P.n56 VSUBS 0.00127f
C2261 P.n57 VSUBS 0.00127f
C2262 P.n58 VSUBS 2.99e-19
C2263 P.n59 VSUBS 1.12e-19
C2264 P.n60 VSUBS 6.74e-19
C2265 P.n61 VSUBS 2.62e-19
C2266 P.t108 VSUBS 2.64f
C2267 P.t58 VSUBS 2.64f
C2268 P.t11 VSUBS 2.64f
C2269 P.t69 VSUBS 2.64f
C2270 P.t53 VSUBS 2.64f
C2271 P.t86 VSUBS 2.64f
C2272 P.t131 VSUBS 2.64f
C2273 P.t26 VSUBS 2.64f
C2274 P.t89 VSUBS 2.64f
C2275 P.t76 VSUBS 2.64f
C2276 P.t100 VSUBS 2.64f
C2277 P.t14 VSUBS 2.78f
C2278 P.n62 VSUBS 4.87f
C2279 P.n63 VSUBS 2.51f
C2280 P.n64 VSUBS 2.51f
C2281 P.n65 VSUBS 2.51f
C2282 P.n66 VSUBS 2.51f
C2283 P.n67 VSUBS 2.51f
C2284 P.n68 VSUBS 2.51f
C2285 P.n69 VSUBS 2.51f
C2286 P.n70 VSUBS 2.51f
C2287 P.n71 VSUBS 2.51f
C2288 P.n72 VSUBS 2.18f
C2289 P.n73 VSUBS 0.101f
C2290 P.n74 VSUBS 9.58e-19
C2291 P.n75 VSUBS 0.00198f
C2292 P.n76 VSUBS 0.00198f
C2293 P.n77 VSUBS 7.52e-19
C2294 P.n78 VSUBS 6.83e-19
C2295 P.n79 VSUBS 0.00198f
C2296 P.n80 VSUBS 0.00198f
C2297 P.n81 VSUBS 9.57e-19
C2298 P.n82 VSUBS 0.00273f
C2299 P.n83 VSUBS 0.00738f
C2300 P.n84 VSUBS 0.00738f
C2301 P.n85 VSUBS 0.00267f
C2302 P.n86 VSUBS 0.0021f
C2303 P.n87 VSUBS 0.00127f
C2304 P.n88 VSUBS 0.00127f
C2305 P.n89 VSUBS 2.99e-19
C2306 P.n90 VSUBS 1.12e-19
C2307 P.n91 VSUBS 2.62e-19
C2308 P.n93 VSUBS 0.00267f
C2309 P.n94 VSUBS 0.0021f
C2310 P.n95 VSUBS 0.00127f
C2311 P.n96 VSUBS 0.00127f
C2312 P.n97 VSUBS 2.99e-19
C2313 P.n98 VSUBS 1.12e-19
C2314 P.n99 VSUBS 2.62e-19
C2315 P.n101 VSUBS 0.00273f
C2316 P.n102 VSUBS 0.00273f
C2317 P.n103 VSUBS 0.00649f
C2318 P.n104 VSUBS 0.43f
C2319 P.n105 VSUBS 0.0041f
C2320 P.n106 VSUBS 0.00198f
C2321 P.n107 VSUBS 0.0015f
C2322 P.n108 VSUBS 0.00258f
C2323 P.n109 VSUBS 3.37e-19
C2324 P.n110 VSUBS 2.25e-19
C2325 P.n111 VSUBS 2.62e-19
C2326 P.n112 VSUBS 2.62e-19
C2327 P.n113 VSUBS 7.86e-19
C2328 P.n114 VSUBS 9.73e-19
C2329 P.n115 VSUBS 0.0208f
C2330 P.n116 VSUBS 5.99e-19
C2331 P.n117 VSUBS 5.99e-19
C2332 P.n118 VSUBS 7.86e-19
C2333 P.n119 VSUBS 0.00124f
C2334 P.n120 VSUBS 0.00127f
C2335 P.n121 VSUBS 8.24e-19
C2336 P.n122 VSUBS 5.99e-19
C2337 P.n123 VSUBS 5.99e-19
C2338 P.n124 VSUBS 0.0024f
C2339 P.n125 VSUBS 0.0024f
C2340 P.n126 VSUBS 0.00127f
C2341 P.n127 VSUBS 0.00124f
C2342 P.n128 VSUBS 1.5e-19
C2343 P.n129 VSUBS 1.87e-19
C2344 P.n130 VSUBS 3e-19
C2345 P.n131 VSUBS 7.49e-19
C2346 P.n132 VSUBS 7.49e-19
C2347 P.n133 VSUBS 3.37e-19
C2348 P.n134 VSUBS 0.0216f
C2349 P.n135 VSUBS 0.00124f
C2350 P.n136 VSUBS 0.00124f
C2351 P.n137 VSUBS 0.00127f
C2352 P.n138 VSUBS 0.00127f
C2353 P.n139 VSUBS 0.00314f
C2354 P.n140 VSUBS 0.00378f
C2355 P.n141 VSUBS 0.00127f
C2356 P.n142 VSUBS 3.37e-19
C2357 P.n143 VSUBS 0.00105f
C2358 P.n144 VSUBS 9.36e-19
C2359 P.n145 VSUBS 0.0201f
C2360 P.n146 VSUBS 3.74e-19
C2361 P.n147 VSUBS 3.57e-19
C2362 P.n148 VSUBS 8.98e-19
C2363 P.n149 VSUBS 9.36e-19
C2364 P.n150 VSUBS 3.37e-19
C2365 P.n151 VSUBS 3.37e-19
C2366 P.n152 VSUBS 8.99e-19
C2367 P.n153 VSUBS 8.99e-19
C2368 P.n154 VSUBS 4.87e-19
C2369 P.n155 VSUBS 0.00337f
C2370 P.n156 VSUBS 0.00378f
C2371 P.n157 VSUBS 0.00105f
C2372 P.n158 VSUBS 5.24e-19
C2373 P.n159 VSUBS 9.73e-19
C2374 P.n160 VSUBS 0.00105f
C2375 P.n161 VSUBS 4.87e-19
C2376 P.n162 VSUBS 3.37e-19
C2377 P.n163 VSUBS 3e-19
C2378 P.n164 VSUBS 8.99e-19
C2379 P.n165 VSUBS 9.73e-19
C2380 P.n166 VSUBS 3.74e-19
C2381 P.n167 VSUBS 3e-19
C2382 P.n168 VSUBS 3e-19
C2383 P.n169 VSUBS 7.49e-19
C2384 P.n170 VSUBS 7.49e-19
C2385 P.n171 VSUBS 0.00288f
C2386 P.n172 VSUBS 0.00288f
C2387 P.n173 VSUBS 3.37e-19
C2388 P.n174 VSUBS 3.37e-19
C2389 P.n175 VSUBS 3e-19
C2390 P.n176 VSUBS 8.99e-19
C2391 P.n177 VSUBS 0.0189f
C2392 P.n178 VSUBS 8.99e-19
C2393 P.n179 VSUBS 3e-19
C2394 P.n180 VSUBS 3.37e-19
C2395 P.n181 VSUBS 2.25e-19
C2396 P.n182 VSUBS 1.5e-19
C2397 P.n183 VSUBS 8.98e-19
C2398 P.n184 VSUBS 9.36e-19
C2399 P.n185 VSUBS 3.37e-19
C2400 P.n186 VSUBS 3.37e-19
C2401 P.n187 VSUBS 8.99e-19
C2402 P.n188 VSUBS 5.01e-19
C2403 P.n189 VSUBS 1.12e-19
C2404 P.n190 VSUBS 0.00116f
C2405 P.n191 VSUBS 0.00116f
C2406 P.n192 VSUBS 0.0015f
C2407 P.n193 VSUBS 0.00951f
C2408 P.n194 VSUBS 5.99e-19
C2409 P.n195 VSUBS 7.86e-19
C2410 P.n196 VSUBS 0.00124f
C2411 P.n197 VSUBS 0.00127f
C2412 P.n198 VSUBS 8.24e-19
C2413 P.n199 VSUBS 5.99e-19
C2414 P.n200 VSUBS 5.99e-19
C2415 P.n201 VSUBS 0.0024f
C2416 P.n202 VSUBS 0.0024f
C2417 P.n203 VSUBS 0.00127f
C2418 P.n204 VSUBS 0.00124f
C2419 P.n205 VSUBS 1.5e-19
C2420 P.n206 VSUBS 1.87e-19
C2421 P.n207 VSUBS 3e-19
C2422 P.n208 VSUBS 7.49e-19
C2423 P.n209 VSUBS 7.49e-19
C2424 P.n210 VSUBS 3.37e-19
C2425 P.n211 VSUBS 0.0109f
C2426 P.n212 VSUBS 0.00124f
C2427 P.n213 VSUBS 0.0226f
C2428 P.n214 VSUBS 4.87e-19
C2429 P.n215 VSUBS 0.00588f
C2430 P.n216 VSUBS 0.00629f
C2431 P.n217 VSUBS 0.00105f
C2432 P.n218 VSUBS 0.00157f
C2433 P.n219 VSUBS 0.00633f
C2434 P.n220 VSUBS 0.00565f
C2435 P.n221 VSUBS 0.0241f
C2436 P.n222 VSUBS 0.0244f
C2437 P.n223 VSUBS 0.00105f
C2438 P.n224 VSUBS 4.87e-19
C2439 P.n225 VSUBS 0.00588f
C2440 P.n226 VSUBS 0.00629f
C2441 P.n227 VSUBS 0.00105f
C2442 P.n228 VSUBS 0.00157f
C2443 P.n229 VSUBS 0.0239f
C2444 P.n230 VSUBS 1.86e-19
C2445 P.n231 VSUBS 0.00127f
C2446 P.n232 VSUBS 0.00127f
C2447 P.n233 VSUBS 0.00314f
C2448 P.n234 VSUBS 0.00378f
C2449 P.n235 VSUBS 0.00127f
C2450 P.n236 VSUBS 3.37e-19
C2451 P.n237 VSUBS 0.00105f
C2452 P.n238 VSUBS 9.36e-19
C2453 P.n239 VSUBS 0.0219f
C2454 P.n240 VSUBS 0.00105f
C2455 P.n241 VSUBS 3.74e-19
C2456 P.n242 VSUBS 3.37e-19
C2457 P.n243 VSUBS 8.98e-19
C2458 P.n244 VSUBS 9.36e-19
C2459 P.n245 VSUBS 3.37e-19
C2460 P.n246 VSUBS 3.37e-19
C2461 P.n247 VSUBS 8.99e-19
C2462 P.n248 VSUBS 8.99e-19
C2463 P.n249 VSUBS 4.87e-19
C2464 P.n250 VSUBS 0.00337f
C2465 P.n251 VSUBS 0.00378f
C2466 P.n252 VSUBS 0.00105f
C2467 P.n253 VSUBS 5.24e-19
C2468 P.n254 VSUBS 9.73e-19
C2469 P.n255 VSUBS 0.00105f
C2470 P.n256 VSUBS 4.87e-19
C2471 P.n257 VSUBS 3.37e-19
C2472 P.n258 VSUBS 3e-19
C2473 P.n259 VSUBS 8.99e-19
C2474 P.n260 VSUBS 9.73e-19
C2475 P.n261 VSUBS 3.74e-19
C2476 P.n262 VSUBS 3e-19
C2477 P.n263 VSUBS 3e-19
C2478 P.n264 VSUBS 7.49e-19
C2479 P.n265 VSUBS 7.49e-19
C2480 P.n266 VSUBS 0.00288f
C2481 P.n267 VSUBS 0.00288f
C2482 P.n268 VSUBS 3.37e-19
C2483 P.n269 VSUBS 3.37e-19
C2484 P.n270 VSUBS 3e-19
C2485 P.n271 VSUBS 8.99e-19
C2486 P.n272 VSUBS 0.0208f
C2487 P.n273 VSUBS 8.99e-19
C2488 P.n274 VSUBS 8.99e-19
C2489 P.n275 VSUBS 3e-19
C2490 P.n276 VSUBS 3.37e-19
C2491 P.n277 VSUBS 2.25e-19
C2492 P.n278 VSUBS 1.5e-19
C2493 P.n279 VSUBS 8.98e-19
C2494 P.n280 VSUBS 9.36e-19
C2495 P.n281 VSUBS 3.37e-19
C2496 P.n282 VSUBS 3.37e-19
C2497 P.n283 VSUBS 8.99e-19
C2498 P.n284 VSUBS 5.01e-19
C2499 P.n285 VSUBS 0.00258f
C2500 P.n286 VSUBS 3.37e-19
C2501 P.n287 VSUBS 2.25e-19
C2502 P.n288 VSUBS 2.62e-19
C2503 P.n289 VSUBS 2.62e-19
C2504 P.n290 VSUBS 7.86e-19
C2505 P.n291 VSUBS 9.73e-19
C2506 P.n292 VSUBS 1.12e-19
C2507 P.n293 VSUBS 0.0013f
C2508 P.n294 VSUBS 7.52e-19
C2509 P.n295 VSUBS 6.83e-19
C2510 P.n296 VSUBS 7.92e-19
C2511 P.n297 VSUBS 0.0205f
C2512 P.n298 VSUBS 5.99e-19
C2513 P.n299 VSUBS 5.99e-19
C2514 P.n300 VSUBS 0.00118f
C2515 P.n301 VSUBS 5.82e-19
C2516 P.n302 VSUBS 0.00116f
C2517 P.n303 VSUBS 0.00157f
C2518 P.n304 VSUBS 0.00123f
C2519 P.n305 VSUBS 0.0091f
C2520 P.n306 VSUBS 5.99e-19
C2521 P.n307 VSUBS 0.00118f
C2522 P.n308 VSUBS 5.82e-19
C2523 P.n309 VSUBS 0.00116f
C2524 P.n310 VSUBS 0.00273f
C2525 P.n311 VSUBS 0.00608f
C2526 P.n312 VSUBS 0.00437f
C2527 P.n313 VSUBS 0.00137f
C2528 P.n314 VSUBS 0.00171f
C2529 P.n315 VSUBS 8.88e-19
C2530 P.n316 VSUBS 6.83e-19
C2531 P.n317 VSUBS 1.73e-19
C2532 P.n318 VSUBS 2.65e-19
C2533 P.n319 VSUBS 0.0186f
C2534 P.n320 VSUBS 8.99e-19
C2535 P.n321 VSUBS 3e-19
C2536 P.n322 VSUBS 3.37e-19
C2537 P.n323 VSUBS 3.37e-19
C2538 P.n324 VSUBS 1.87e-19
C2539 P.n325 VSUBS 1.26e-19
C2540 P.n326 VSUBS 8.99e-19
C2541 P.n327 VSUBS 8.99e-19
C2542 P.n328 VSUBS 3.46e-20
C2543 P.n329 VSUBS 6.83e-19
C2544 P.n330 VSUBS 0.00247f
C2545 P.n331 VSUBS 7.49e-19
C2546 P.n332 VSUBS 7.49e-19
C2547 P.n333 VSUBS 3e-19
C2548 P.n334 VSUBS 3e-19
C2549 P.n335 VSUBS 5.24e-19
C2550 P.n336 VSUBS 4.49e-19
C2551 P.n337 VSUBS 5.47e-19
C2552 P.n338 VSUBS 9.51e-19
C2553 P.n339 VSUBS 6.74e-19
C2554 P.n340 VSUBS 7.49e-19
C2555 P.n341 VSUBS 6.88e-19
C2556 P.n342 VSUBS 1.73e-19
C2557 P.n343 VSUBS 2.25e-19
C2558 P.n344 VSUBS 3.4e-19
C2559 P.n345 VSUBS 3.46e-20
C2560 P.n346 VSUBS 6.83e-19
C2561 P.n347 VSUBS 0.00109f
C2562 P.n348 VSUBS 0.00198f
C2563 P.n349 VSUBS 5.99e-19
C2564 P.n350 VSUBS 5.99e-19
C2565 P.n351 VSUBS 9.73e-19
C2566 P.n352 VSUBS 8.99e-19
C2567 P.n353 VSUBS 4.06e-19
C2568 P.n354 VSUBS 0.0013f
C2569 P.n355 VSUBS 1.73e-19
C2570 P.n356 VSUBS 2.65e-19
C2571 P.n357 VSUBS 0.0204f
C2572 P.n358 VSUBS 8.99e-19
C2573 P.n359 VSUBS 8.99e-19
C2574 P.n360 VSUBS 3e-19
C2575 P.n361 VSUBS 3.37e-19
C2576 P.n362 VSUBS 3.37e-19
C2577 P.n363 VSUBS 1.87e-19
C2578 P.n364 VSUBS 1.26e-19
C2579 P.n365 VSUBS 6.9e-19
C2580 P.n366 VSUBS 0.00111f
C2581 P.n367 VSUBS 3.46e-20
C2582 P.n368 VSUBS 8.88e-19
C2583 P.n369 VSUBS 6.74e-19
C2584 P.n370 VSUBS 7.49e-19
C2585 P.n371 VSUBS 6.88e-19
C2586 P.n372 VSUBS 1.73e-19
C2587 P.n373 VSUBS 2.25e-19
C2588 P.n374 VSUBS 3.4e-19
C2589 P.n375 VSUBS 0.00247f
C2590 P.n376 VSUBS 7.49e-19
C2591 P.n377 VSUBS 7.49e-19
C2592 P.n378 VSUBS 3e-19
C2593 P.n379 VSUBS 3e-19
C2594 P.n380 VSUBS 5.24e-19
C2595 P.n381 VSUBS 4.49e-19
C2596 P.n382 VSUBS 5.47e-19
C2597 P.n383 VSUBS 9.51e-19
C2598 P.n384 VSUBS 3.46e-20
C2599 P.n385 VSUBS 7.52e-19
C2600 P.n386 VSUBS 7.52e-19
C2601 P.n387 VSUBS 6.15e-19
C2602 P.n388 VSUBS 0.00198f
C2603 P.n389 VSUBS 5.99e-19
C2604 P.n390 VSUBS 5.99e-19
C2605 P.n391 VSUBS 9.73e-19
C2606 P.n392 VSUBS 8.99e-19
C2607 P.n393 VSUBS 7.92e-19
C2608 P.n394 VSUBS 4.06e-19
C2609 P.n395 VSUBS 0.00109f
C2610 P.n396 VSUBS 0.00137f
C2611 P.n397 VSUBS 8.88e-19
C2612 P.n398 VSUBS 0.00137f
C2613 P.n399 VSUBS 0.338f
C2614 P.n400 VSUBS 0.333f
C2615 P.n401 VSUBS 0.00294f
C2616 P.n402 VSUBS 0.00212f
C2617 P.n403 VSUBS 0.00246f
C2618 P.n404 VSUBS 8.2e-19
C2619 P.n405 VSUBS 0.00205f
C2620 P.n406 VSUBS 0.00212f
C2621 P.n407 VSUBS 8.88e-19
C2622 P.n408 VSUBS 0.00246f
C2623 P.n409 VSUBS 0.00205f
C2624 P.n410 VSUBS 0.00294f
C2625 P.n411 VSUBS 0.00249f
C2626 P.n412 VSUBS 0.0081f
C2627 P.n414 VSUBS 0.00478f
C2628 P.n415 VSUBS 0.00273f
C2629 P.n416 VSUBS 0.00239f
C2630 P.n417 VSUBS 0.424f
C2631 P.n418 VSUBS 0.00301f
C2632 P.n419 VSUBS 0.0021f
C2633 P.n420 VSUBS 0.00127f
C2634 P.n421 VSUBS 0.00127f
C2635 P.n422 VSUBS 2.99e-19
C2636 P.n423 VSUBS 1.12e-19
C2637 P.n424 VSUBS 6.74e-19
C2638 P.n425 VSUBS 2.62e-19
C2639 P.n427 VSUBS 0.00738f
C2640 P.n428 VSUBS 0.00581f
C2641 P.n429 VSUBS 0.00267f
C2642 P.n430 VSUBS 0.0189f
C2643 P.n431 VSUBS 5.99e-19
C2644 P.n432 VSUBS 5.99e-19
C2645 P.n433 VSUBS 7.86e-19
C2646 P.n434 VSUBS 0.00124f
C2647 P.n435 VSUBS 0.00127f
C2648 P.n436 VSUBS 8.24e-19
C2649 P.n437 VSUBS 5.99e-19
C2650 P.n438 VSUBS 5.99e-19
C2651 P.n439 VSUBS 0.0024f
C2652 P.n440 VSUBS 0.0024f
C2653 P.n441 VSUBS 0.00127f
C2654 P.n442 VSUBS 0.00124f
C2655 P.n443 VSUBS 1.5e-19
C2656 P.n444 VSUBS 1.87e-19
C2657 P.n445 VSUBS 3e-19
C2658 P.n446 VSUBS 7.49e-19
C2659 P.n447 VSUBS 7.49e-19
C2660 P.n448 VSUBS 3.37e-19
C2661 P.n449 VSUBS 0.0196f
C2662 P.n450 VSUBS 0.00124f
C2663 P.n451 VSUBS 0.00124f
C2664 P.n452 VSUBS 0.00127f
C2665 P.n453 VSUBS 0.00127f
C2666 P.n454 VSUBS 0.00314f
C2667 P.n455 VSUBS 0.00378f
C2668 P.n456 VSUBS 0.00127f
C2669 P.n457 VSUBS 3.37e-19
C2670 P.n458 VSUBS 0.00105f
C2671 P.n459 VSUBS 9.36e-19
C2672 P.n460 VSUBS 0.024f
C2673 P.n461 VSUBS 3.74e-19
C2674 P.n462 VSUBS 3.61e-19
C2675 P.n463 VSUBS 8.98e-19
C2676 P.n464 VSUBS 9.36e-19
C2677 P.n465 VSUBS 3.37e-19
C2678 P.n466 VSUBS 3.37e-19
C2679 P.n467 VSUBS 8.99e-19
C2680 P.n468 VSUBS 8.99e-19
C2681 P.n469 VSUBS 4.87e-19
C2682 P.n470 VSUBS 0.00337f
C2683 P.n471 VSUBS 0.00378f
C2684 P.n472 VSUBS 0.00105f
C2685 P.n473 VSUBS 5.24e-19
C2686 P.n474 VSUBS 9.73e-19
C2687 P.n475 VSUBS 0.00105f
C2688 P.n476 VSUBS 4.87e-19
C2689 P.n477 VSUBS 3.37e-19
C2690 P.n478 VSUBS 3e-19
C2691 P.n479 VSUBS 8.99e-19
C2692 P.n480 VSUBS 9.73e-19
C2693 P.n481 VSUBS 3.74e-19
C2694 P.n482 VSUBS 3e-19
C2695 P.n483 VSUBS 3e-19
C2696 P.n484 VSUBS 7.49e-19
C2697 P.n485 VSUBS 7.49e-19
C2698 P.n486 VSUBS 0.00288f
C2699 P.n487 VSUBS 0.00288f
C2700 P.n488 VSUBS 3.37e-19
C2701 P.n489 VSUBS 3.37e-19
C2702 P.n490 VSUBS 3e-19
C2703 P.n491 VSUBS 8.99e-19
C2704 P.n492 VSUBS 0.0228f
C2705 P.n493 VSUBS 8.99e-19
C2706 P.n494 VSUBS 3e-19
C2707 P.n495 VSUBS 3.37e-19
C2708 P.n496 VSUBS 2.25e-19
C2709 P.n497 VSUBS 1.5e-19
C2710 P.n498 VSUBS 8.98e-19
C2711 P.n499 VSUBS 9.36e-19
C2712 P.n500 VSUBS 3.37e-19
C2713 P.n501 VSUBS 3.37e-19
C2714 P.n502 VSUBS 8.99e-19
C2715 P.n503 VSUBS 5.01e-19
C2716 P.n504 VSUBS 0.00258f
C2717 P.n505 VSUBS 3.37e-19
C2718 P.n506 VSUBS 2.25e-19
C2719 P.n507 VSUBS 2.62e-19
C2720 P.n508 VSUBS 2.62e-19
C2721 P.n509 VSUBS 7.86e-19
C2722 P.n510 VSUBS 9.73e-19
C2723 P.n511 VSUBS 1.12e-19
C2724 P.n512 VSUBS 0.00198f
C2725 P.n513 VSUBS 0.00116f
C2726 P.n514 VSUBS 0.00164f
C2727 P.n515 VSUBS 0.00157f
C2728 P.n516 VSUBS 0.00103f
C2729 P.n517 VSUBS 0.0186f
C2730 P.n518 VSUBS 5.99e-19
C2731 P.n519 VSUBS 5.99e-19
C2732 P.n520 VSUBS 0.00118f
C2733 P.n521 VSUBS 7.92e-19
C2734 P.n522 VSUBS 5.82e-19
C2735 P.n523 VSUBS 5.47e-19
C2736 P.n524 VSUBS 7.52e-19
C2737 P.n525 VSUBS 0.0015f
C2738 P.n526 VSUBS 0.00258f
C2739 P.n527 VSUBS 3.37e-19
C2740 P.n528 VSUBS 2.25e-19
C2741 P.n529 VSUBS 2.62e-19
C2742 P.n530 VSUBS 2.62e-19
C2743 P.n531 VSUBS 7.86e-19
C2744 P.n532 VSUBS 9.73e-19
C2745 P.n533 VSUBS 0.00951f
C2746 P.n534 VSUBS 5.99e-19
C2747 P.n535 VSUBS 7.86e-19
C2748 P.n536 VSUBS 0.00124f
C2749 P.n537 VSUBS 0.00127f
C2750 P.n538 VSUBS 8.24e-19
C2751 P.n539 VSUBS 5.99e-19
C2752 P.n540 VSUBS 5.99e-19
C2753 P.n541 VSUBS 0.0024f
C2754 P.n542 VSUBS 0.0024f
C2755 P.n543 VSUBS 0.00127f
C2756 P.n544 VSUBS 0.00124f
C2757 P.n545 VSUBS 1.5e-19
C2758 P.n546 VSUBS 1.87e-19
C2759 P.n547 VSUBS 3e-19
C2760 P.n548 VSUBS 7.49e-19
C2761 P.n549 VSUBS 7.49e-19
C2762 P.n550 VSUBS 3.37e-19
C2763 P.n551 VSUBS 0.0109f
C2764 P.n552 VSUBS 0.00124f
C2765 P.n553 VSUBS 0.0265f
C2766 P.n554 VSUBS 4.87e-19
C2767 P.n555 VSUBS 0.00588f
C2768 P.n556 VSUBS 0.00629f
C2769 P.n557 VSUBS 0.00105f
C2770 P.n558 VSUBS 0.00157f
C2771 P.n559 VSUBS 0.00633f
C2772 P.n560 VSUBS 0.00565f
C2773 P.n561 VSUBS 0.0221f
C2774 P.n562 VSUBS 0.0224f
C2775 P.n563 VSUBS 0.00105f
C2776 P.n564 VSUBS 4.87e-19
C2777 P.n565 VSUBS 0.00588f
C2778 P.n566 VSUBS 0.00629f
C2779 P.n567 VSUBS 0.00105f
C2780 P.n568 VSUBS 0.00157f
C2781 P.n569 VSUBS 0.0239f
C2782 P.n570 VSUBS 1.86e-19
C2783 P.n571 VSUBS 0.00127f
C2784 P.n572 VSUBS 0.00127f
C2785 P.n573 VSUBS 0.00314f
C2786 P.n574 VSUBS 0.00378f
C2787 P.n575 VSUBS 0.00127f
C2788 P.n576 VSUBS 3.37e-19
C2789 P.n577 VSUBS 0.00105f
C2790 P.n578 VSUBS 9.36e-19
C2791 P.n579 VSUBS 0.0199f
C2792 P.n580 VSUBS 0.00105f
C2793 P.n581 VSUBS 3.74e-19
C2794 P.n582 VSUBS 3.37e-19
C2795 P.n583 VSUBS 8.98e-19
C2796 P.n584 VSUBS 9.36e-19
C2797 P.n585 VSUBS 3.37e-19
C2798 P.n586 VSUBS 3.37e-19
C2799 P.n587 VSUBS 8.99e-19
C2800 P.n588 VSUBS 8.99e-19
C2801 P.n589 VSUBS 4.87e-19
C2802 P.n590 VSUBS 0.00337f
C2803 P.n591 VSUBS 0.00378f
C2804 P.n592 VSUBS 0.00105f
C2805 P.n593 VSUBS 5.24e-19
C2806 P.n594 VSUBS 9.73e-19
C2807 P.n595 VSUBS 0.00105f
C2808 P.n596 VSUBS 4.87e-19
C2809 P.n597 VSUBS 3.37e-19
C2810 P.n598 VSUBS 3e-19
C2811 P.n599 VSUBS 8.99e-19
C2812 P.n600 VSUBS 9.73e-19
C2813 P.n601 VSUBS 3.74e-19
C2814 P.n602 VSUBS 3e-19
C2815 P.n603 VSUBS 3e-19
C2816 P.n604 VSUBS 7.49e-19
C2817 P.n605 VSUBS 7.49e-19
C2818 P.n606 VSUBS 0.00288f
C2819 P.n607 VSUBS 0.00288f
C2820 P.n608 VSUBS 3.37e-19
C2821 P.n609 VSUBS 3.37e-19
C2822 P.n610 VSUBS 3e-19
C2823 P.n611 VSUBS 8.99e-19
C2824 P.n612 VSUBS 0.0189f
C2825 P.n613 VSUBS 8.99e-19
C2826 P.n614 VSUBS 8.99e-19
C2827 P.n615 VSUBS 3e-19
C2828 P.n616 VSUBS 3.37e-19
C2829 P.n617 VSUBS 2.25e-19
C2830 P.n618 VSUBS 1.5e-19
C2831 P.n619 VSUBS 8.98e-19
C2832 P.n620 VSUBS 9.36e-19
C2833 P.n621 VSUBS 3.37e-19
C2834 P.n622 VSUBS 3.37e-19
C2835 P.n623 VSUBS 8.99e-19
C2836 P.n624 VSUBS 5.01e-19
C2837 P.n625 VSUBS 1.12e-19
C2838 P.n626 VSUBS 0.00137f
C2839 P.n627 VSUBS 0.00109f
C2840 P.n628 VSUBS 6.83e-19
C2841 P.n629 VSUBS 0.00164f
C2842 P.n630 VSUBS 0.00198f
C2843 P.n631 VSUBS 0.0091f
C2844 P.n632 VSUBS 5.99e-19
C2845 P.n633 VSUBS 0.00118f
C2846 P.n634 VSUBS 7.92e-19
C2847 P.n635 VSUBS 5.82e-19
C2848 P.n636 VSUBS 0.00116f
C2849 P.n637 VSUBS 0.00273f
C2850 P.n638 VSUBS 0.00328f
C2851 P.n639 VSUBS 0.00157f
C2852 P.n640 VSUBS 0.00137f
C2853 P.n641 VSUBS 0.00239f
C2854 P.n642 VSUBS 1.73e-19
C2855 P.n643 VSUBS 2.65e-19
C2856 P.n644 VSUBS 0.0225f
C2857 P.n645 VSUBS 8.99e-19
C2858 P.n646 VSUBS 3e-19
C2859 P.n647 VSUBS 3.37e-19
C2860 P.n648 VSUBS 3.37e-19
C2861 P.n649 VSUBS 1.87e-19
C2862 P.n650 VSUBS 1.12e-19
C2863 P.n651 VSUBS 8.99e-19
C2864 P.n652 VSUBS 8.99e-19
C2865 P.n653 VSUBS 3.46e-20
C2866 P.n654 VSUBS 0.00157f
C2867 P.n655 VSUBS 0.00247f
C2868 P.n656 VSUBS 7.49e-19
C2869 P.n657 VSUBS 7.49e-19
C2870 P.n658 VSUBS 3e-19
C2871 P.n659 VSUBS 3e-19
C2872 P.n660 VSUBS 5.24e-19
C2873 P.n661 VSUBS 4.49e-19
C2874 P.n662 VSUBS 5.47e-19
C2875 P.n663 VSUBS 9.51e-19
C2876 P.n664 VSUBS 7.49e-19
C2877 P.n665 VSUBS 6.88e-19
C2878 P.n666 VSUBS 1.73e-19
C2879 P.n667 VSUBS 2.25e-19
C2880 P.n668 VSUBS 3.4e-19
C2881 P.n669 VSUBS 3.46e-20
C2882 P.n670 VSUBS 0.00137f
C2883 P.n671 VSUBS 0.00198f
C2884 P.n672 VSUBS 5.99e-19
C2885 P.n673 VSUBS 5.99e-19
C2886 P.n674 VSUBS 9.73e-19
C2887 P.n675 VSUBS 8.99e-19
C2888 P.n676 VSUBS 4.06e-19
C2889 P.n677 VSUBS 0.00185f
C2890 P.n678 VSUBS 0.00103f
C2891 P.n679 VSUBS 6.15e-19
C2892 P.n680 VSUBS 6.15e-19
C2893 P.n681 VSUBS 7.52e-19
C2894 P.n682 VSUBS 0.00109f
C2895 P.n683 VSUBS 0.0013f
C2896 P.n684 VSUBS 0.0185f
C2897 P.n685 VSUBS 8.99e-19
C2898 P.n686 VSUBS 8.99e-19
C2899 P.n687 VSUBS 3e-19
C2900 P.n688 VSUBS 3.37e-19
C2901 P.n689 VSUBS 3.37e-19
C2902 P.n690 VSUBS 1.87e-19
C2903 P.n691 VSUBS 1.12e-19
C2904 P.n692 VSUBS 6.9e-19
C2905 P.n693 VSUBS 0.00111f
C2906 P.n694 VSUBS 1.73e-19
C2907 P.n695 VSUBS 2.65e-19
C2908 P.n696 VSUBS 3.46e-20
C2909 P.n697 VSUBS 9.57e-19
C2910 P.n698 VSUBS 7.49e-19
C2911 P.n699 VSUBS 6.88e-19
C2912 P.n700 VSUBS 1.73e-19
C2913 P.n701 VSUBS 2.25e-19
C2914 P.n702 VSUBS 3.4e-19
C2915 P.n703 VSUBS 0.00247f
C2916 P.n704 VSUBS 7.49e-19
C2917 P.n705 VSUBS 7.49e-19
C2918 P.n706 VSUBS 3e-19
C2919 P.n707 VSUBS 3e-19
C2920 P.n708 VSUBS 5.24e-19
C2921 P.n709 VSUBS 4.49e-19
C2922 P.n710 VSUBS 7.49e-19
C2923 P.n711 VSUBS 7.49e-19
C2924 P.n712 VSUBS 3.46e-20
C2925 P.n713 VSUBS 0.00137f
C2926 P.n714 VSUBS 0.00198f
C2927 P.n715 VSUBS 5.99e-19
C2928 P.n716 VSUBS 5.99e-19
C2929 P.n717 VSUBS 9.73e-19
C2930 P.n718 VSUBS 8.99e-19
C2931 P.n719 VSUBS 4.06e-19
C2932 P.n720 VSUBS 0.00246f
C2933 P.n721 VSUBS 0.00164f
C2934 P.n722 VSUBS 0.00137f
C2935 P.n723 VSUBS 0.456f
C2936 P.n724 VSUBS 0.457f
C2937 P.n725 VSUBS 0.00267f
C2938 P.n726 VSUBS 0.00137f
C2939 P.n727 VSUBS 0.00157f
C2940 P.n728 VSUBS 0.00157f
C2941 P.n729 VSUBS 0.00116f
C2942 P.n730 VSUBS 0.00109f
C2943 P.n731 VSUBS 0.00157f
C2944 P.n732 VSUBS 0.00157f
C2945 P.n733 VSUBS 0.00137f
C2946 P.n734 VSUBS 0.00273f
C2947 P.n735 VSUBS 0.00738f
C2948 P.n736 VSUBS 0.00738f
C2949 P.n737 VSUBS 0.00267f
C2950 P.n738 VSUBS 0.00267f
C2951 P.n739 VSUBS 0.00273f
C2952 P.n740 VSUBS 0.00178f
C2953 P.n741 VSUBS 0.424f
C2954 P.n742 VSUBS 0.00882f
C2955 P.n743 VSUBS 0.00902f
C2956 P.n744 VSUBS 0.00157f
C2957 P.n745 VSUBS 0.0015f
C2958 P.n746 VSUBS 0.00258f
C2959 P.n747 VSUBS 3.37e-19
C2960 P.n748 VSUBS 2.25e-19
C2961 P.n749 VSUBS 2.62e-19
C2962 P.n750 VSUBS 2.62e-19
C2963 P.n751 VSUBS 7.86e-19
C2964 P.n752 VSUBS 9.73e-19
C2965 P.n753 VSUBS 1.12e-19
C2966 P.n754 VSUBS 0.00116f
C2967 P.n755 VSUBS 4.78e-19
C2968 P.n756 VSUBS 0.00109f
C2969 P.n757 VSUBS 0.00109f
C2970 P.n758 VSUBS 0.00258f
C2971 P.n759 VSUBS 3.37e-19
C2972 P.n760 VSUBS 2.25e-19
C2973 P.n761 VSUBS 2.62e-19
C2974 P.n762 VSUBS 2.62e-19
C2975 P.n763 VSUBS 7.86e-19
C2976 P.n764 VSUBS 9.73e-19
C2977 P.n765 VSUBS 1.12e-19
C2978 P.n766 VSUBS 8.88e-19
C2979 P.n767 VSUBS 0.00116f
C2980 P.n768 VSUBS 0.00109f
C2981 P.n769 VSUBS 0.019f
C2982 P.n770 VSUBS 5.99e-19
C2983 P.n771 VSUBS 5.99e-19
C2984 P.n772 VSUBS 0.00118f
C2985 P.n773 VSUBS 5.82e-19
C2986 P.n774 VSUBS 0.00116f
C2987 P.n775 VSUBS 0.00116f
C2988 P.n776 VSUBS 8.2e-19
C2989 P.n777 VSUBS 0.0091f
C2990 P.n778 VSUBS 5.99e-19
C2991 P.n779 VSUBS 0.00118f
C2992 P.n780 VSUBS 5.82e-19
C2993 P.n781 VSUBS 0.00116f
C2994 P.n782 VSUBS 0.00116f
C2995 P.n783 VSUBS 0.00198f
C2996 P.n784 VSUBS 0.00608f
C2997 P.n785 VSUBS 0.00478f
C2998 P.n786 VSUBS 0.00137f
C2999 P.n787 VSUBS 0.0013f
C3000 P.n788 VSUBS 4.78e-19
C3001 P.n789 VSUBS 0.00109f
C3002 P.n790 VSUBS 0.0216f
C3003 P.n791 VSUBS 8.99e-19
C3004 P.n792 VSUBS 3e-19
C3005 P.n793 VSUBS 3.37e-19
C3006 P.n794 VSUBS 3.37e-19
C3007 P.n795 VSUBS 1.87e-19
C3008 P.n796 VSUBS 1.12e-19
C3009 P.n797 VSUBS 6.9e-19
C3010 P.n798 VSUBS 0.00111f
C3011 P.n799 VSUBS 0.0193f
C3012 P.n800 VSUBS 5.99e-19
C3013 P.n801 VSUBS 5.99e-19
C3014 P.n802 VSUBS 7.86e-19
C3015 P.n803 VSUBS 0.00124f
C3016 P.n804 VSUBS 0.00127f
C3017 P.n805 VSUBS 8.24e-19
C3018 P.n806 VSUBS 5.99e-19
C3019 P.n807 VSUBS 5.99e-19
C3020 P.n808 VSUBS 0.0024f
C3021 P.n809 VSUBS 0.0024f
C3022 P.n810 VSUBS 0.00127f
C3023 P.n811 VSUBS 0.00124f
C3024 P.n812 VSUBS 1.5e-19
C3025 P.n813 VSUBS 1.87e-19
C3026 P.n814 VSUBS 3e-19
C3027 P.n815 VSUBS 7.49e-19
C3028 P.n816 VSUBS 7.49e-19
C3029 P.n817 VSUBS 3.37e-19
C3030 P.n818 VSUBS 0.0201f
C3031 P.n819 VSUBS 0.00124f
C3032 P.n820 VSUBS 0.00124f
C3033 P.n821 VSUBS 0.00127f
C3034 P.n822 VSUBS 0.00127f
C3035 P.n823 VSUBS 0.00314f
C3036 P.n824 VSUBS 0.00378f
C3037 P.n825 VSUBS 0.00127f
C3038 P.n826 VSUBS 3.37e-19
C3039 P.n827 VSUBS 0.00105f
C3040 P.n828 VSUBS 9.36e-19
C3041 P.n829 VSUBS 0.0231f
C3042 P.n830 VSUBS 3.74e-19
C3043 P.n831 VSUBS 3.6e-19
C3044 P.n832 VSUBS 8.98e-19
C3045 P.n833 VSUBS 9.36e-19
C3046 P.n834 VSUBS 3.37e-19
C3047 P.n835 VSUBS 3.37e-19
C3048 P.n836 VSUBS 8.99e-19
C3049 P.n837 VSUBS 8.99e-19
C3050 P.n838 VSUBS 4.87e-19
C3051 P.n839 VSUBS 0.00337f
C3052 P.n840 VSUBS 0.00378f
C3053 P.n841 VSUBS 0.00105f
C3054 P.n842 VSUBS 5.24e-19
C3055 P.n843 VSUBS 9.73e-19
C3056 P.n844 VSUBS 0.00105f
C3057 P.n845 VSUBS 4.87e-19
C3058 P.n846 VSUBS 3.37e-19
C3059 P.n847 VSUBS 3e-19
C3060 P.n848 VSUBS 8.99e-19
C3061 P.n849 VSUBS 9.73e-19
C3062 P.n850 VSUBS 3.74e-19
C3063 P.n851 VSUBS 3e-19
C3064 P.n852 VSUBS 3e-19
C3065 P.n853 VSUBS 7.49e-19
C3066 P.n854 VSUBS 7.49e-19
C3067 P.n855 VSUBS 0.00288f
C3068 P.n856 VSUBS 0.00288f
C3069 P.n857 VSUBS 3.37e-19
C3070 P.n858 VSUBS 3.37e-19
C3071 P.n859 VSUBS 3e-19
C3072 P.n860 VSUBS 8.99e-19
C3073 P.n861 VSUBS 0.0219f
C3074 P.n862 VSUBS 8.99e-19
C3075 P.n863 VSUBS 3e-19
C3076 P.n864 VSUBS 3.37e-19
C3077 P.n865 VSUBS 2.25e-19
C3078 P.n866 VSUBS 1.5e-19
C3079 P.n867 VSUBS 8.98e-19
C3080 P.n868 VSUBS 9.36e-19
C3081 P.n869 VSUBS 3.37e-19
C3082 P.n870 VSUBS 3.37e-19
C3083 P.n871 VSUBS 8.99e-19
C3084 P.n872 VSUBS 5.01e-19
C3085 P.n873 VSUBS 1.73e-19
C3086 P.n874 VSUBS 2.65e-19
C3087 P.n875 VSUBS 3.46e-20
C3088 P.n876 VSUBS 0.00109f
C3089 P.n877 VSUBS 0.00247f
C3090 P.n878 VSUBS 7.49e-19
C3091 P.n879 VSUBS 7.49e-19
C3092 P.n880 VSUBS 3e-19
C3093 P.n881 VSUBS 3e-19
C3094 P.n882 VSUBS 5.24e-19
C3095 P.n883 VSUBS 4.49e-19
C3096 P.n884 VSUBS 5.47e-19
C3097 P.n885 VSUBS 9.51e-19
C3098 P.n886 VSUBS 0.0021f
C3099 P.n887 VSUBS 0.00127f
C3100 P.n888 VSUBS 0.00127f
C3101 P.n889 VSUBS 2.99e-19
C3102 P.n890 VSUBS 1.12e-19
C3103 P.n892 VSUBS 2.62e-19
C3104 P.n893 VSUBS 6.74e-19
C3105 P.n894 VSUBS 7.49e-19
C3106 P.n895 VSUBS 6.88e-19
C3107 P.n896 VSUBS 1.73e-19
C3108 P.n897 VSUBS 2.25e-19
C3109 P.n898 VSUBS 3.4e-19
C3110 P.n899 VSUBS 3.46e-20
C3111 P.n900 VSUBS 0.00137f
C3112 P.n901 VSUBS 0.00198f
C3113 P.n902 VSUBS 5.99e-19
C3114 P.n903 VSUBS 5.99e-19
C3115 P.n904 VSUBS 9.73e-19
C3116 P.n905 VSUBS 8.99e-19
C3117 P.n906 VSUBS 7.92e-19
C3118 P.n907 VSUBS 4.06e-19
C3119 P.n908 VSUBS 0.0013f
C3120 P.n909 VSUBS 0.00951f
C3121 P.n910 VSUBS 5.99e-19
C3122 P.n911 VSUBS 7.86e-19
C3123 P.n912 VSUBS 0.00124f
C3124 P.n913 VSUBS 0.00127f
C3125 P.n914 VSUBS 8.24e-19
C3126 P.n915 VSUBS 5.99e-19
C3127 P.n916 VSUBS 5.99e-19
C3128 P.n917 VSUBS 0.0024f
C3129 P.n918 VSUBS 0.0024f
C3130 P.n919 VSUBS 0.00127f
C3131 P.n920 VSUBS 0.00124f
C3132 P.n921 VSUBS 1.5e-19
C3133 P.n922 VSUBS 1.87e-19
C3134 P.n923 VSUBS 3e-19
C3135 P.n924 VSUBS 7.49e-19
C3136 P.n925 VSUBS 7.49e-19
C3137 P.n926 VSUBS 3.37e-19
C3138 P.n927 VSUBS 0.0109f
C3139 P.n928 VSUBS 0.00124f
C3140 P.n929 VSUBS 0.0256f
C3141 P.n930 VSUBS 4.87e-19
C3142 P.n931 VSUBS 0.00588f
C3143 P.n932 VSUBS 0.00629f
C3144 P.n933 VSUBS 0.00105f
C3145 P.n934 VSUBS 0.00157f
C3146 P.n935 VSUBS 0.00633f
C3147 P.n936 VSUBS 0.00565f
C3148 P.n937 VSUBS 0.0226f
C3149 P.n938 VSUBS 0.0229f
C3150 P.n939 VSUBS 0.00105f
C3151 P.n940 VSUBS 4.87e-19
C3152 P.n941 VSUBS 0.00588f
C3153 P.n942 VSUBS 0.00629f
C3154 P.n943 VSUBS 0.00105f
C3155 P.n944 VSUBS 0.00157f
C3156 P.n945 VSUBS 0.0239f
C3157 P.n946 VSUBS 1.86e-19
C3158 P.n947 VSUBS 0.00127f
C3159 P.n948 VSUBS 0.00127f
C3160 P.n949 VSUBS 0.00314f
C3161 P.n950 VSUBS 0.00378f
C3162 P.n951 VSUBS 0.00127f
C3163 P.n952 VSUBS 3.37e-19
C3164 P.n953 VSUBS 0.00105f
C3165 P.n954 VSUBS 9.36e-19
C3166 P.n955 VSUBS 0.0204f
C3167 P.n956 VSUBS 0.00105f
C3168 P.n957 VSUBS 3.74e-19
C3169 P.n958 VSUBS 3.37e-19
C3170 P.n959 VSUBS 8.98e-19
C3171 P.n960 VSUBS 9.36e-19
C3172 P.n961 VSUBS 3.37e-19
C3173 P.n962 VSUBS 3.37e-19
C3174 P.n963 VSUBS 8.99e-19
C3175 P.n964 VSUBS 8.99e-19
C3176 P.n965 VSUBS 4.87e-19
C3177 P.n966 VSUBS 0.00337f
C3178 P.n967 VSUBS 0.00378f
C3179 P.n968 VSUBS 0.00105f
C3180 P.n969 VSUBS 5.24e-19
C3181 P.n970 VSUBS 9.73e-19
C3182 P.n971 VSUBS 0.00105f
C3183 P.n972 VSUBS 4.87e-19
C3184 P.n973 VSUBS 3.37e-19
C3185 P.n974 VSUBS 3e-19
C3186 P.n975 VSUBS 8.99e-19
C3187 P.n976 VSUBS 9.73e-19
C3188 P.n977 VSUBS 3.74e-19
C3189 P.n978 VSUBS 3e-19
C3190 P.n979 VSUBS 3e-19
C3191 P.n980 VSUBS 7.49e-19
C3192 P.n981 VSUBS 7.49e-19
C3193 P.n982 VSUBS 0.00288f
C3194 P.n983 VSUBS 0.00288f
C3195 P.n984 VSUBS 3.37e-19
C3196 P.n985 VSUBS 3.37e-19
C3197 P.n986 VSUBS 3e-19
C3198 P.n987 VSUBS 8.99e-19
C3199 P.n988 VSUBS 0.0193f
C3200 P.n989 VSUBS 8.99e-19
C3201 P.n990 VSUBS 8.99e-19
C3202 P.n991 VSUBS 3e-19
C3203 P.n992 VSUBS 3.37e-19
C3204 P.n993 VSUBS 2.25e-19
C3205 P.n994 VSUBS 1.5e-19
C3206 P.n995 VSUBS 8.98e-19
C3207 P.n996 VSUBS 9.36e-19
C3208 P.n997 VSUBS 3.37e-19
C3209 P.n998 VSUBS 3.37e-19
C3210 P.n999 VSUBS 8.99e-19
C3211 P.n1000 VSUBS 5.01e-19
C3212 P.n1001 VSUBS 1.73e-19
C3213 P.n1002 VSUBS 2.65e-19
C3214 P.n1003 VSUBS 0.0189f
C3215 P.n1004 VSUBS 8.99e-19
C3216 P.n1005 VSUBS 8.99e-19
C3217 P.n1006 VSUBS 3e-19
C3218 P.n1007 VSUBS 3.37e-19
C3219 P.n1008 VSUBS 3.37e-19
C3220 P.n1009 VSUBS 1.87e-19
C3221 P.n1010 VSUBS 1.12e-19
C3222 P.n1011 VSUBS 6.9e-19
C3223 P.n1012 VSUBS 0.00111f
C3224 P.n1013 VSUBS 3.46e-20
C3225 P.n1014 VSUBS 4.78e-19
C3226 P.n1015 VSUBS 0.00247f
C3227 P.n1016 VSUBS 7.49e-19
C3228 P.n1017 VSUBS 7.49e-19
C3229 P.n1018 VSUBS 3e-19
C3230 P.n1019 VSUBS 3e-19
C3231 P.n1020 VSUBS 5.24e-19
C3232 P.n1021 VSUBS 4.49e-19
C3233 P.n1022 VSUBS 5.47e-19
C3234 P.n1023 VSUBS 9.51e-19
C3235 P.n1024 VSUBS 0.0021f
C3236 P.n1025 VSUBS 0.00127f
C3237 P.n1026 VSUBS 0.00127f
C3238 P.n1027 VSUBS 2.99e-19
C3239 P.n1028 VSUBS 1.12e-19
C3240 P.n1030 VSUBS 2.62e-19
C3241 P.n1031 VSUBS 6.74e-19
C3242 P.n1032 VSUBS 7.49e-19
C3243 P.n1033 VSUBS 6.88e-19
C3244 P.n1034 VSUBS 1.73e-19
C3245 P.n1035 VSUBS 2.25e-19
C3246 P.n1036 VSUBS 3.4e-19
C3247 P.n1037 VSUBS 3.46e-20
C3248 P.n1038 VSUBS 0.00116f
C3249 P.n1039 VSUBS 0.00109f
C3250 P.n1040 VSUBS 7.92e-19
C3251 P.n1041 VSUBS 0.00198f
C3252 P.n1042 VSUBS 5.99e-19
C3253 P.n1043 VSUBS 5.99e-19
C3254 P.n1044 VSUBS 9.73e-19
C3255 P.n1045 VSUBS 8.99e-19
C3256 P.n1046 VSUBS 4.06e-19
C3257 P.n1047 VSUBS 2.73e-19
C3258 P.n1048 VSUBS 0.00116f
C3259 P.n1049 VSUBS 0.0013f
C3260 P.n1050 VSUBS 4.78e-19
C3261 P.n1051 VSUBS 0.00137f
C3262 P.n1052 VSUBS 0.427f
C3263 P.n1053 VSUBS 0.429f
C3264 P.n1055 VSUBS 0.00294f
C3265 P.n1056 VSUBS 0.00273f
C3266 P.n1057 VSUBS 0.00267f
C3267 P.n1058 VSUBS 0.00294f
C3268 P.n1059 VSUBS 0.00554f
C3269 P.n1060 VSUBS 0.43f
C3270 P.n1061 VSUBS 0.00724f
C3271 P.n1063 VSUBS 0.0054f
C3272 P.n1065 VSUBS 0.0122f
C3273 P.n1066 VSUBS 0.0106f
C3274 P.n1067 VSUBS 0.00267f
C3275 P.n1068 VSUBS 0.00258f
C3276 P.n1069 VSUBS 3.37e-19
C3277 P.n1070 VSUBS 2.25e-19
C3278 P.n1071 VSUBS 2.62e-19
C3279 P.n1072 VSUBS 2.62e-19
C3280 P.n1073 VSUBS 7.86e-19
C3281 P.n1074 VSUBS 9.73e-19
C3282 P.n1075 VSUBS 1.12e-19
C3283 P.n1076 VSUBS 0.00198f
C3284 P.n1077 VSUBS 0.00116f
C3285 P.n1078 VSUBS 0.00226f
C3286 P.n1079 VSUBS 0.00198f
C3287 P.n1080 VSUBS 0.0142f
C3288 P.n1081 VSUBS 5.99e-19
C3289 P.n1082 VSUBS 5.99e-19
C3290 P.n1083 VSUBS 0.00118f
C3291 P.n1084 VSUBS 5.82e-19
C3292 P.n1085 VSUBS 0.0182f
C3293 P.n1086 VSUBS 5.99e-19
C3294 P.n1087 VSUBS 0.00118f
C3295 P.n1088 VSUBS 5.82e-19
C3296 P.n1089 VSUBS 0.00116f
C3297 P.n1090 VSUBS 0.00273f
C3298 P.n1091 VSUBS 0.00806f
C3299 P.n1092 VSUBS 0.00636f
C3300 P.n1093 VSUBS 0.00137f
C3301 P.n1094 VSUBS 0.00239f
C3302 P.n1095 VSUBS 0.0141f
C3303 P.n1096 VSUBS 8.99e-19
C3304 P.n1097 VSUBS 8.99e-19
C3305 P.n1098 VSUBS 3e-19
C3306 P.n1099 VSUBS 3.37e-19
C3307 P.n1100 VSUBS 3.37e-19
C3308 P.n1101 VSUBS 1.87e-19
C3309 P.n1102 VSUBS 1.12e-19
C3310 P.n1103 VSUBS 8.99e-19
C3311 P.n1104 VSUBS 8.99e-19
C3312 P.n1105 VSUBS 0.00258f
C3313 P.n1106 VSUBS 3.37e-19
C3314 P.n1107 VSUBS 2.25e-19
C3315 P.n1108 VSUBS 2.62e-19
C3316 P.n1109 VSUBS 2.62e-19
C3317 P.n1110 VSUBS 7.86e-19
C3318 P.n1111 VSUBS 9.73e-19
C3319 P.n1112 VSUBS 1.12e-19
C3320 P.n1113 VSUBS 0.0186f
C3321 P.n1114 VSUBS 5.99e-19
C3322 P.n1115 VSUBS 7.86e-19
C3323 P.n1116 VSUBS 0.00124f
C3324 P.n1117 VSUBS 0.00127f
C3325 P.n1118 VSUBS 8.24e-19
C3326 P.n1119 VSUBS 5.99e-19
C3327 P.n1120 VSUBS 5.99e-19
C3328 P.n1121 VSUBS 0.0024f
C3329 P.n1122 VSUBS 0.0024f
C3330 P.n1123 VSUBS 0.00127f
C3331 P.n1124 VSUBS 0.00124f
C3332 P.n1125 VSUBS 1.5e-19
C3333 P.n1126 VSUBS 1.87e-19
C3334 P.n1127 VSUBS 3e-19
C3335 P.n1128 VSUBS 7.49e-19
C3336 P.n1129 VSUBS 7.49e-19
C3337 P.n1130 VSUBS 3.37e-19
C3338 P.n1131 VSUBS 0.02f
C3339 P.n1132 VSUBS 0.00125f
C3340 P.n1133 VSUBS 0.026f
C3341 P.n1134 VSUBS 4.87e-19
C3342 P.n1135 VSUBS 0.00588f
C3343 P.n1136 VSUBS 0.00629f
C3344 P.n1137 VSUBS 0.00105f
C3345 P.n1138 VSUBS 0.00157f
C3346 P.n1139 VSUBS 0.00633f
C3347 P.n1140 VSUBS 0.00565f
C3348 P.n1141 VSUBS 0.0178f
C3349 P.n1142 VSUBS 0.0181f
C3350 P.n1143 VSUBS 0.00105f
C3351 P.n1144 VSUBS 4.87e-19
C3352 P.n1145 VSUBS 0.00588f
C3353 P.n1146 VSUBS 0.00629f
C3354 P.n1147 VSUBS 0.00105f
C3355 P.n1148 VSUBS 0.00157f
C3356 P.n1149 VSUBS 0.033f
C3357 P.n1150 VSUBS 2.82e-19
C3358 P.n1151 VSUBS 0.00127f
C3359 P.n1152 VSUBS 0.00127f
C3360 P.n1153 VSUBS 0.00314f
C3361 P.n1154 VSUBS 0.00378f
C3362 P.n1155 VSUBS 0.00127f
C3363 P.n1156 VSUBS 3.37e-19
C3364 P.n1157 VSUBS 0.00105f
C3365 P.n1158 VSUBS 9.36e-19
C3366 P.n1159 VSUBS 0.0156f
C3367 P.n1160 VSUBS 0.00105f
C3368 P.n1161 VSUBS 3.74e-19
C3369 P.n1162 VSUBS 3.37e-19
C3370 P.n1163 VSUBS 8.98e-19
C3371 P.n1164 VSUBS 9.36e-19
C3372 P.n1165 VSUBS 3.37e-19
C3373 P.n1166 VSUBS 3.37e-19
C3374 P.n1167 VSUBS 8.99e-19
C3375 P.n1168 VSUBS 8.99e-19
C3376 P.n1169 VSUBS 4.87e-19
C3377 P.n1170 VSUBS 0.00337f
C3378 P.n1171 VSUBS 0.00378f
C3379 P.n1172 VSUBS 0.00105f
C3380 P.n1173 VSUBS 5.24e-19
C3381 P.n1174 VSUBS 9.73e-19
C3382 P.n1175 VSUBS 0.00105f
C3383 P.n1176 VSUBS 4.87e-19
C3384 P.n1177 VSUBS 3.37e-19
C3385 P.n1178 VSUBS 3e-19
C3386 P.n1179 VSUBS 8.99e-19
C3387 P.n1180 VSUBS 9.73e-19
C3388 P.n1181 VSUBS 3.74e-19
C3389 P.n1182 VSUBS 3e-19
C3390 P.n1183 VSUBS 3e-19
C3391 P.n1184 VSUBS 7.49e-19
C3392 P.n1185 VSUBS 7.49e-19
C3393 P.n1186 VSUBS 0.00288f
C3394 P.n1187 VSUBS 0.00288f
C3395 P.n1188 VSUBS 3.37e-19
C3396 P.n1189 VSUBS 3.37e-19
C3397 P.n1190 VSUBS 3e-19
C3398 P.n1191 VSUBS 8.99e-19
C3399 P.n1192 VSUBS 0.0145f
C3400 P.n1193 VSUBS 8.99e-19
C3401 P.n1194 VSUBS 8.99e-19
C3402 P.n1195 VSUBS 3e-19
C3403 P.n1196 VSUBS 3.37e-19
C3404 P.n1197 VSUBS 2.25e-19
C3405 P.n1198 VSUBS 1.5e-19
C3406 P.n1199 VSUBS 8.98e-19
C3407 P.n1200 VSUBS 9.36e-19
C3408 P.n1201 VSUBS 3.37e-19
C3409 P.n1202 VSUBS 3.37e-19
C3410 P.n1203 VSUBS 8.99e-19
C3411 P.n1204 VSUBS 3.37e-19
C3412 P.n1205 VSUBS 3.37e-19
C3413 P.n1206 VSUBS 2.65e-19
C3414 P.n1207 VSUBS 3.46e-20
C3415 P.n1208 VSUBS 0.0145f
C3416 P.n1209 VSUBS 5.99e-19
C3417 P.n1210 VSUBS 5.99e-19
C3418 P.n1211 VSUBS 7.86e-19
C3419 P.n1212 VSUBS 0.00124f
C3420 P.n1213 VSUBS 0.00127f
C3421 P.n1214 VSUBS 8.24e-19
C3422 P.n1215 VSUBS 5.99e-19
C3423 P.n1216 VSUBS 5.99e-19
C3424 P.n1217 VSUBS 0.0024f
C3425 P.n1218 VSUBS 0.0024f
C3426 P.n1219 VSUBS 0.00127f
C3427 P.n1220 VSUBS 0.00124f
C3428 P.n1221 VSUBS 1.5e-19
C3429 P.n1222 VSUBS 1.87e-19
C3430 P.n1223 VSUBS 3e-19
C3431 P.n1224 VSUBS 7.49e-19
C3432 P.n1225 VSUBS 7.49e-19
C3433 P.n1226 VSUBS 3.37e-19
C3434 P.n1227 VSUBS 0.0153f
C3435 P.n1228 VSUBS 0.00124f
C3436 P.n1229 VSUBS 0.00124f
C3437 P.n1230 VSUBS 0.00127f
C3438 P.n1231 VSUBS 0.00127f
C3439 P.n1232 VSUBS 0.00314f
C3440 P.n1233 VSUBS 0.00378f
C3441 P.n1234 VSUBS 0.00127f
C3442 P.n1235 VSUBS 3.37e-19
C3443 P.n1236 VSUBS 0.00105f
C3444 P.n1237 VSUBS 9.36e-19
C3445 P.n1238 VSUBS 0.0235f
C3446 P.n1239 VSUBS 3.74e-19
C3447 P.n1240 VSUBS 3.6e-19
C3448 P.n1241 VSUBS 8.98e-19
C3449 P.n1242 VSUBS 9.36e-19
C3450 P.n1243 VSUBS 3.37e-19
C3451 P.n1244 VSUBS 3.37e-19
C3452 P.n1245 VSUBS 8.99e-19
C3453 P.n1246 VSUBS 8.99e-19
C3454 P.n1247 VSUBS 4.87e-19
C3455 P.n1248 VSUBS 0.00337f
C3456 P.n1249 VSUBS 0.00378f
C3457 P.n1250 VSUBS 0.00105f
C3458 P.n1251 VSUBS 5.24e-19
C3459 P.n1252 VSUBS 9.73e-19
C3460 P.n1253 VSUBS 0.00105f
C3461 P.n1254 VSUBS 4.87e-19
C3462 P.n1255 VSUBS 3.37e-19
C3463 P.n1256 VSUBS 3e-19
C3464 P.n1257 VSUBS 8.99e-19
C3465 P.n1258 VSUBS 9.73e-19
C3466 P.n1259 VSUBS 3.74e-19
C3467 P.n1260 VSUBS 3e-19
C3468 P.n1261 VSUBS 3e-19
C3469 P.n1262 VSUBS 7.49e-19
C3470 P.n1263 VSUBS 7.49e-19
C3471 P.n1264 VSUBS 0.00288f
C3472 P.n1265 VSUBS 0.00288f
C3473 P.n1266 VSUBS 3.37e-19
C3474 P.n1267 VSUBS 3.37e-19
C3475 P.n1268 VSUBS 3e-19
C3476 P.n1269 VSUBS 8.99e-19
C3477 P.n1270 VSUBS 0.0223f
C3478 P.n1271 VSUBS 8.99e-19
C3479 P.n1272 VSUBS 3e-19
C3480 P.n1273 VSUBS 3.37e-19
C3481 P.n1274 VSUBS 2.25e-19
C3482 P.n1275 VSUBS 1.5e-19
C3483 P.n1276 VSUBS 8.98e-19
C3484 P.n1277 VSUBS 9.36e-19
C3485 P.n1278 VSUBS 3.37e-19
C3486 P.n1279 VSUBS 3.37e-19
C3487 P.n1280 VSUBS 8.99e-19
C3488 P.n1281 VSUBS 5.01e-19
C3489 P.n1282 VSUBS 1.73e-19
C3490 P.n1283 VSUBS 2.65e-19
C3491 P.n1284 VSUBS 0.022f
C3492 P.n1285 VSUBS 8.99e-19
C3493 P.n1286 VSUBS 3e-19
C3494 P.n1287 VSUBS 3.37e-19
C3495 P.n1288 VSUBS 3.37e-19
C3496 P.n1289 VSUBS 1.87e-19
C3497 P.n1290 VSUBS 1.12e-19
C3498 P.n1291 VSUBS 6.9e-19
C3499 P.n1292 VSUBS 0.00111f
C3500 P.n1293 VSUBS 3.46e-20
C3501 P.n1294 VSUBS 0.00157f
C3502 P.n1295 VSUBS 0.00247f
C3503 P.n1296 VSUBS 7.49e-19
C3504 P.n1297 VSUBS 7.49e-19
C3505 P.n1298 VSUBS 3e-19
C3506 P.n1299 VSUBS 3e-19
C3507 P.n1300 VSUBS 5.24e-19
C3508 P.n1301 VSUBS 4.49e-19
C3509 P.n1302 VSUBS 5.47e-19
C3510 P.n1303 VSUBS 9.51e-19
C3511 P.n1304 VSUBS 0.0021f
C3512 P.n1305 VSUBS 0.00127f
C3513 P.n1306 VSUBS 0.00127f
C3514 P.n1307 VSUBS 2.99e-19
C3515 P.n1308 VSUBS 1.12e-19
C3516 P.n1309 VSUBS 2.62e-19
C3517 P.n1310 VSUBS 6.74e-19
C3518 P.n1311 VSUBS 7.49e-19
C3519 P.n1312 VSUBS 6.88e-19
C3520 P.n1313 VSUBS 1.73e-19
C3521 P.n1314 VSUBS 2.25e-19
C3522 P.n1315 VSUBS 3.4e-19
C3523 P.n1316 VSUBS 3.46e-20
C3524 P.n1317 VSUBS 0.0021f
C3525 P.n1318 VSUBS 0.00127f
C3526 P.n1319 VSUBS 0.00127f
C3527 P.n1320 VSUBS 2.99e-19
C3528 P.n1321 VSUBS 1.12e-19
C3529 P.n1323 VSUBS 2.62e-19
C3530 P.n1324 VSUBS 6.74e-19
C3531 P.n1325 VSUBS 7.49e-19
C3532 P.n1326 VSUBS 6.88e-19
C3533 P.n1327 VSUBS 1.73e-19
C3534 P.n1328 VSUBS 2.25e-19
C3535 P.n1329 VSUBS 3.4e-19
C3536 P.n1330 VSUBS 0.00247f
C3537 P.n1331 VSUBS 7.49e-19
C3538 P.n1332 VSUBS 7.49e-19
C3539 P.n1333 VSUBS 3e-19
C3540 P.n1334 VSUBS 3e-19
C3541 P.n1335 VSUBS 5.24e-19
C3542 P.n1336 VSUBS 4.49e-19
C3543 P.n1337 VSUBS 5.47e-19
C3544 P.n1338 VSUBS 9.51e-19
C3545 P.n1339 VSUBS 3.46e-20
C3546 P.n1340 VSUBS 0.00137f
C3547 P.n1341 VSUBS 7.92e-19
C3548 P.n1342 VSUBS 0.00198f
C3549 P.n1343 VSUBS 5.99e-19
C3550 P.n1344 VSUBS 5.99e-19
C3551 P.n1345 VSUBS 9.73e-19
C3552 P.n1346 VSUBS 8.99e-19
C3553 P.n1347 VSUBS 4.06e-19
C3554 P.n1348 VSUBS 7.92e-19
C3555 P.n1349 VSUBS 0.00198f
C3556 P.n1350 VSUBS 5.99e-19
C3557 P.n1351 VSUBS 5.99e-19
C3558 P.n1352 VSUBS 9.73e-19
C3559 P.n1353 VSUBS 8.99e-19
C3560 P.n1354 VSUBS 4.06e-19
C3561 P.n1355 VSUBS 0.00246f
C3562 P.n1356 VSUBS 0.00164f
C3563 P.n1357 VSUBS 0.00137f
C3564 P.n1358 VSUBS 0.416f
C3565 P.n1359 VSUBS 0.416f
C3566 P.n1360 VSUBS 0.00267f
C3567 P.n1361 VSUBS 0.00219f
C3568 P.n1362 VSUBS 7.52e-19
C3569 P.n1363 VSUBS 7.54e-19
C3570 P.n1364 VSUBS 5.47e-19
C3571 P.n1365 VSUBS 0.424f
C3572 P.n1366 VSUBS 0.00164f
C3573 P.n1367 VSUBS 7.52e-19
C3574 P.n1368 VSUBS 7.52e-19
C3575 P.n1369 VSUBS 0.00219f
C3576 P.n1370 VSUBS 0.00273f
C3577 P.n1371 VSUBS 0.00738f
C3578 P.n1372 VSUBS 0.00738f
C3579 P.n1373 VSUBS 0.00267f
C3580 P.n1374 VSUBS 0.00267f
C3581 P.n1375 VSUBS 0.00273f
C3582 P.n1376 VSUBS 0.00273f
C3583 P.n1377 VSUBS 0.00943f
C3584 P.n1378 VSUBS 0.00943f
C3585 P.n1379 VSUBS 0.00116f
C3586 P.n1380 VSUBS 0.00116f
C3587 P.n1381 VSUBS 0.0015f
C3588 P.n1382 VSUBS 0.00123f
C3589 P.n1383 VSUBS 7.52e-19
C3590 P.n1384 VSUBS 6.83e-19
C3591 P.n1385 VSUBS 4.78e-19
C3592 P.n1386 VSUBS 7.52e-19
C3593 P.n1387 VSUBS 0.0015f
C3594 P.n1388 VSUBS 0.00123f
C3595 P.n1389 VSUBS 0.0157f
C3596 P.n1390 VSUBS 5.99e-19
C3597 P.n1391 VSUBS 0.00118f
C3598 P.n1392 VSUBS 5.82e-19
C3599 P.n1393 VSUBS 7.54e-19
C3600 P.n1394 VSUBS 7.52e-19
C3601 P.n1395 VSUBS 0.0133f
C3602 P.n1396 VSUBS 5.99e-19
C3603 P.n1397 VSUBS 5.99e-19
C3604 P.n1398 VSUBS 0.00118f
C3605 P.n1399 VSUBS 5.82e-19
C3606 P.n1400 VSUBS 0.00116f
C3607 P.n1401 VSUBS 0.00198f
C3608 P.n1402 VSUBS 0.00198f
C3609 P.n1403 VSUBS 0.00608f
C3610 P.n1404 VSUBS 0.0056f
C3611 P.n1405 VSUBS 7.52e-19
C3612 P.n1406 VSUBS 7.52e-19
C3613 P.n1407 VSUBS 6.15e-19
C3614 P.n1408 VSUBS 0.00109f
C3615 P.n1409 VSUBS 0.0013f
C3616 P.n1410 VSUBS 0.0132f
C3617 P.n1411 VSUBS 8.99e-19
C3618 P.n1412 VSUBS 8.99e-19
C3619 P.n1413 VSUBS 3e-19
C3620 P.n1414 VSUBS 3.37e-19
C3621 P.n1415 VSUBS 3.37e-19
C3622 P.n1416 VSUBS 1.87e-19
C3623 P.n1417 VSUBS 1.12e-19
C3624 P.n1418 VSUBS 6.9e-19
C3625 P.n1419 VSUBS 0.00111f
C3626 P.n1420 VSUBS 0.00258f
C3627 P.n1421 VSUBS 3.37e-19
C3628 P.n1422 VSUBS 2.25e-19
C3629 P.n1423 VSUBS 2.62e-19
C3630 P.n1424 VSUBS 2.62e-19
C3631 P.n1425 VSUBS 7.86e-19
C3632 P.n1426 VSUBS 9.73e-19
C3633 P.n1427 VSUBS 1.12e-19
C3634 P.n1428 VSUBS 0.0161f
C3635 P.n1429 VSUBS 5.99e-19
C3636 P.n1430 VSUBS 7.86e-19
C3637 P.n1431 VSUBS 0.00124f
C3638 P.n1432 VSUBS 0.00127f
C3639 P.n1433 VSUBS 8.24e-19
C3640 P.n1434 VSUBS 5.99e-19
C3641 P.n1435 VSUBS 5.99e-19
C3642 P.n1436 VSUBS 0.0024f
C3643 P.n1437 VSUBS 0.0024f
C3644 P.n1438 VSUBS 0.00127f
C3645 P.n1439 VSUBS 0.00124f
C3646 P.n1440 VSUBS 1.5e-19
C3647 P.n1441 VSUBS 1.87e-19
C3648 P.n1442 VSUBS 3e-19
C3649 P.n1443 VSUBS 7.49e-19
C3650 P.n1444 VSUBS 7.49e-19
C3651 P.n1445 VSUBS 3.37e-19
C3652 P.n1446 VSUBS 0.0175f
C3653 P.n1447 VSUBS 0.00125f
C3654 P.n1448 VSUBS 0.0304f
C3655 P.n1449 VSUBS 4.87e-19
C3656 P.n1450 VSUBS 0.00588f
C3657 P.n1451 VSUBS 0.00629f
C3658 P.n1452 VSUBS 0.00105f
C3659 P.n1453 VSUBS 0.00157f
C3660 P.n1454 VSUBS 0.00633f
C3661 P.n1455 VSUBS 0.00565f
C3662 P.n1456 VSUBS 0.0169f
C3663 P.n1457 VSUBS 0.0172f
C3664 P.n1458 VSUBS 0.00105f
C3665 P.n1459 VSUBS 4.87e-19
C3666 P.n1460 VSUBS 0.00588f
C3667 P.n1461 VSUBS 0.00629f
C3668 P.n1462 VSUBS 0.00105f
C3669 P.n1463 VSUBS 0.00157f
C3670 P.n1464 VSUBS 0.0304f
C3671 P.n1465 VSUBS 2.55e-19
C3672 P.n1466 VSUBS 0.00127f
C3673 P.n1467 VSUBS 0.00127f
C3674 P.n1468 VSUBS 0.00314f
C3675 P.n1469 VSUBS 0.00378f
C3676 P.n1470 VSUBS 0.00127f
C3677 P.n1471 VSUBS 3.37e-19
C3678 P.n1472 VSUBS 0.00105f
C3679 P.n1473 VSUBS 9.36e-19
C3680 P.n1474 VSUBS 0.0147f
C3681 P.n1475 VSUBS 0.00105f
C3682 P.n1476 VSUBS 3.74e-19
C3683 P.n1477 VSUBS 3.37e-19
C3684 P.n1478 VSUBS 8.98e-19
C3685 P.n1479 VSUBS 9.36e-19
C3686 P.n1480 VSUBS 3.37e-19
C3687 P.n1481 VSUBS 3.37e-19
C3688 P.n1482 VSUBS 8.99e-19
C3689 P.n1483 VSUBS 8.99e-19
C3690 P.n1484 VSUBS 4.87e-19
C3691 P.n1485 VSUBS 0.00337f
C3692 P.n1486 VSUBS 0.00378f
C3693 P.n1487 VSUBS 0.00105f
C3694 P.n1488 VSUBS 5.24e-19
C3695 P.n1489 VSUBS 9.73e-19
C3696 P.n1490 VSUBS 0.00105f
C3697 P.n1491 VSUBS 4.87e-19
C3698 P.n1492 VSUBS 3.37e-19
C3699 P.n1493 VSUBS 3e-19
C3700 P.n1494 VSUBS 8.99e-19
C3701 P.n1495 VSUBS 9.73e-19
C3702 P.n1496 VSUBS 3.74e-19
C3703 P.n1497 VSUBS 3e-19
C3704 P.n1498 VSUBS 3e-19
C3705 P.n1499 VSUBS 7.49e-19
C3706 P.n1500 VSUBS 7.49e-19
C3707 P.n1501 VSUBS 0.00288f
C3708 P.n1502 VSUBS 0.00288f
C3709 P.n1503 VSUBS 3.37e-19
C3710 P.n1504 VSUBS 3.37e-19
C3711 P.n1505 VSUBS 3e-19
C3712 P.n1506 VSUBS 8.99e-19
C3713 P.n1507 VSUBS 0.0136f
C3714 P.n1508 VSUBS 8.99e-19
C3715 P.n1509 VSUBS 8.99e-19
C3716 P.n1510 VSUBS 3e-19
C3717 P.n1511 VSUBS 3.37e-19
C3718 P.n1512 VSUBS 2.25e-19
C3719 P.n1513 VSUBS 1.5e-19
C3720 P.n1514 VSUBS 8.98e-19
C3721 P.n1515 VSUBS 9.36e-19
C3722 P.n1516 VSUBS 3.37e-19
C3723 P.n1517 VSUBS 3.37e-19
C3724 P.n1518 VSUBS 8.99e-19
C3725 P.n1519 VSUBS 5.01e-19
C3726 P.n1520 VSUBS 1.73e-19
C3727 P.n1521 VSUBS 2.65e-19
C3728 P.n1522 VSUBS 3.46e-20
C3729 P.n1523 VSUBS 8.2e-19
C3730 P.n1524 VSUBS 0.00247f
C3731 P.n1525 VSUBS 7.49e-19
C3732 P.n1526 VSUBS 7.49e-19
C3733 P.n1527 VSUBS 3e-19
C3734 P.n1528 VSUBS 3e-19
C3735 P.n1529 VSUBS 5.24e-19
C3736 P.n1530 VSUBS 4.49e-19
C3737 P.n1531 VSUBS 5.47e-19
C3738 P.n1532 VSUBS 9.51e-19
C3739 P.n1533 VSUBS 0.0021f
C3740 P.n1534 VSUBS 0.00127f
C3741 P.n1535 VSUBS 0.00127f
C3742 P.n1536 VSUBS 2.99e-19
C3743 P.n1537 VSUBS 1.12e-19
C3744 P.n1539 VSUBS 2.62e-19
C3745 P.n1540 VSUBS 6.74e-19
C3746 P.n1541 VSUBS 7.49e-19
C3747 P.n1542 VSUBS 6.88e-19
C3748 P.n1543 VSUBS 1.73e-19
C3749 P.n1544 VSUBS 2.25e-19
C3750 P.n1545 VSUBS 3.4e-19
C3751 P.n1546 VSUBS 3.46e-20
C3752 P.n1547 VSUBS 7.52e-19
C3753 P.n1548 VSUBS 0.00258f
C3754 P.n1549 VSUBS 3.37e-19
C3755 P.n1550 VSUBS 2.25e-19
C3756 P.n1551 VSUBS 2.62e-19
C3757 P.n1552 VSUBS 2.62e-19
C3758 P.n1553 VSUBS 7.86e-19
C3759 P.n1554 VSUBS 9.73e-19
C3760 P.n1555 VSUBS 1.12e-19
C3761 P.n1556 VSUBS 0.0136f
C3762 P.n1557 VSUBS 5.99e-19
C3763 P.n1558 VSUBS 5.99e-19
C3764 P.n1559 VSUBS 7.86e-19
C3765 P.n1560 VSUBS 0.00124f
C3766 P.n1561 VSUBS 0.00127f
C3767 P.n1562 VSUBS 8.24e-19
C3768 P.n1563 VSUBS 5.99e-19
C3769 P.n1564 VSUBS 5.99e-19
C3770 P.n1565 VSUBS 0.0024f
C3771 P.n1566 VSUBS 0.0024f
C3772 P.n1567 VSUBS 0.00127f
C3773 P.n1568 VSUBS 0.00124f
C3774 P.n1569 VSUBS 1.5e-19
C3775 P.n1570 VSUBS 1.87e-19
C3776 P.n1571 VSUBS 3e-19
C3777 P.n1572 VSUBS 7.49e-19
C3778 P.n1573 VSUBS 7.49e-19
C3779 P.n1574 VSUBS 3.37e-19
C3780 P.n1575 VSUBS 0.0144f
C3781 P.n1576 VSUBS 0.00124f
C3782 P.n1577 VSUBS 0.00124f
C3783 P.n1578 VSUBS 0.00127f
C3784 P.n1579 VSUBS 0.00127f
C3785 P.n1580 VSUBS 0.00314f
C3786 P.n1581 VSUBS 0.00378f
C3787 P.n1582 VSUBS 0.00127f
C3788 P.n1583 VSUBS 3.37e-19
C3789 P.n1584 VSUBS 0.00105f
C3790 P.n1585 VSUBS 9.36e-19
C3791 P.n1586 VSUBS 0.0278f
C3792 P.n1587 VSUBS 3.74e-19
C3793 P.n1588 VSUBS 3.65e-19
C3794 P.n1589 VSUBS 8.98e-19
C3795 P.n1590 VSUBS 9.36e-19
C3796 P.n1591 VSUBS 3.37e-19
C3797 P.n1592 VSUBS 3.37e-19
C3798 P.n1593 VSUBS 8.99e-19
C3799 P.n1594 VSUBS 8.99e-19
C3800 P.n1595 VSUBS 4.87e-19
C3801 P.n1596 VSUBS 0.00337f
C3802 P.n1597 VSUBS 0.00378f
C3803 P.n1598 VSUBS 0.00105f
C3804 P.n1599 VSUBS 5.24e-19
C3805 P.n1600 VSUBS 9.73e-19
C3806 P.n1601 VSUBS 0.00105f
C3807 P.n1602 VSUBS 4.87e-19
C3808 P.n1603 VSUBS 3.37e-19
C3809 P.n1604 VSUBS 3e-19
C3810 P.n1605 VSUBS 8.99e-19
C3811 P.n1606 VSUBS 9.73e-19
C3812 P.n1607 VSUBS 3.74e-19
C3813 P.n1608 VSUBS 3e-19
C3814 P.n1609 VSUBS 3e-19
C3815 P.n1610 VSUBS 7.49e-19
C3816 P.n1611 VSUBS 7.49e-19
C3817 P.n1612 VSUBS 0.00288f
C3818 P.n1613 VSUBS 0.00288f
C3819 P.n1614 VSUBS 3.37e-19
C3820 P.n1615 VSUBS 3.37e-19
C3821 P.n1616 VSUBS 3e-19
C3822 P.n1617 VSUBS 8.99e-19
C3823 P.n1618 VSUBS 0.0267f
C3824 P.n1619 VSUBS 8.99e-19
C3825 P.n1620 VSUBS 3e-19
C3826 P.n1621 VSUBS 3.37e-19
C3827 P.n1622 VSUBS 2.25e-19
C3828 P.n1623 VSUBS 1.5e-19
C3829 P.n1624 VSUBS 8.98e-19
C3830 P.n1625 VSUBS 9.36e-19
C3831 P.n1626 VSUBS 3.37e-19
C3832 P.n1627 VSUBS 3.37e-19
C3833 P.n1628 VSUBS 8.99e-19
C3834 P.n1629 VSUBS 5.01e-19
C3835 P.n1630 VSUBS 1.73e-19
C3836 P.n1631 VSUBS 2.65e-19
C3837 P.n1632 VSUBS 0.0264f
C3838 P.n1633 VSUBS 8.99e-19
C3839 P.n1634 VSUBS 3e-19
C3840 P.n1635 VSUBS 3.37e-19
C3841 P.n1636 VSUBS 3.37e-19
C3842 P.n1637 VSUBS 1.87e-19
C3843 P.n1638 VSUBS 1.12e-19
C3844 P.n1639 VSUBS 6.9e-19
C3845 P.n1640 VSUBS 0.00111f
C3846 P.n1641 VSUBS 3.46e-20
C3847 P.n1642 VSUBS 7.52e-19
C3848 P.n1643 VSUBS 0.00247f
C3849 P.n1644 VSUBS 7.49e-19
C3850 P.n1645 VSUBS 7.49e-19
C3851 P.n1646 VSUBS 3e-19
C3852 P.n1647 VSUBS 3e-19
C3853 P.n1648 VSUBS 5.24e-19
C3854 P.n1649 VSUBS 4.49e-19
C3855 P.n1650 VSUBS 5.47e-19
C3856 P.n1651 VSUBS 9.51e-19
C3857 P.n1652 VSUBS 0.0021f
C3858 P.n1653 VSUBS 0.00127f
C3859 P.n1654 VSUBS 0.00127f
C3860 P.n1655 VSUBS 2.99e-19
C3861 P.n1656 VSUBS 1.12e-19
C3862 P.n1658 VSUBS 2.62e-19
C3863 P.n1659 VSUBS 6.74e-19
C3864 P.n1660 VSUBS 7.49e-19
C3865 P.n1661 VSUBS 6.88e-19
C3866 P.n1662 VSUBS 1.73e-19
C3867 P.n1663 VSUBS 2.25e-19
C3868 P.n1664 VSUBS 3.4e-19
C3869 P.n1665 VSUBS 3.46e-20
C3870 P.n1666 VSUBS 6.15e-19
C3871 P.n1667 VSUBS 7.92e-19
C3872 P.n1668 VSUBS 0.00198f
C3873 P.n1669 VSUBS 5.99e-19
C3874 P.n1670 VSUBS 5.99e-19
C3875 P.n1671 VSUBS 9.73e-19
C3876 P.n1672 VSUBS 8.99e-19
C3877 P.n1673 VSUBS 4.06e-19
C3878 P.n1674 VSUBS 0.00109f
C3879 P.n1675 VSUBS 7.92e-19
C3880 P.n1676 VSUBS 0.00198f
C3881 P.n1677 VSUBS 5.99e-19
C3882 P.n1678 VSUBS 5.99e-19
C3883 P.n1679 VSUBS 9.73e-19
C3884 P.n1680 VSUBS 8.99e-19
C3885 P.n1681 VSUBS 4.06e-19
C3886 P.n1682 VSUBS 0.00137f
C3887 P.n1683 VSUBS 8.88e-19
C3888 P.n1684 VSUBS 7.52e-19
C3889 P.n1685 VSUBS 7.52e-19
C3890 P.n1686 VSUBS 6.15e-19
C3891 P.n1687 VSUBS 0.00109f
C3892 P.n1688 VSUBS 0.415f
C3893 P.n1689 VSUBS 0.836f
C3894 P.n1690 VSUBS 0.00157f
C3895 P.n1691 VSUBS 0.00267f
C3896 P.n1692 VSUBS 0.00178f
C3897 P.n1693 VSUBS 0.00116f
C3898 P.n1694 VSUBS 0.00116f
C3899 P.n1695 VSUBS 0.00157f
C3900 P.n1696 VSUBS 0.0015f
C3901 P.n1697 VSUBS 0.00116f
C3902 P.n1698 VSUBS 0.00116f
C3903 P.n1699 VSUBS 0.00178f
C3904 P.n1700 VSUBS 0.00273f
C3905 P.n1701 VSUBS 0.00738f
C3906 P.n1702 VSUBS 0.00738f
C3907 P.n1703 VSUBS 0.00267f
C3908 P.n1704 VSUBS 0.00267f
C3909 P.n1705 VSUBS 0.00273f
C3910 P.n1706 VSUBS 0.00273f
C3911 P.n1707 VSUBS 0.00943f
C3912 P.n1708 VSUBS 0.00943f
C3913 P.n1709 VSUBS 0.00232f
C3914 P.n1710 VSUBS 0.0015f
C3915 P.n1711 VSUBS 0.00258f
C3916 P.n1712 VSUBS 3.37e-19
C3917 P.n1713 VSUBS 2.25e-19
C3918 P.n1714 VSUBS 2.62e-19
C3919 P.n1715 VSUBS 2.62e-19
C3920 P.n1716 VSUBS 7.86e-19
C3921 P.n1717 VSUBS 9.73e-19
C3922 P.n1718 VSUBS 1.12e-19
C3923 P.n1719 VSUBS 8.2e-19
C3924 P.n1720 VSUBS 0.00116f
C3925 P.n1721 VSUBS 0.00258f
C3926 P.n1722 VSUBS 3.37e-19
C3927 P.n1723 VSUBS 2.25e-19
C3928 P.n1724 VSUBS 2.62e-19
C3929 P.n1725 VSUBS 2.62e-19
C3930 P.n1726 VSUBS 7.86e-19
C3931 P.n1727 VSUBS 9.73e-19
C3932 P.n1728 VSUBS 1.12e-19
C3933 P.n1729 VSUBS 0.00116f
C3934 P.n1730 VSUBS 0.00116f
C3935 P.n1731 VSUBS 0.00109f
C3936 P.n1732 VSUBS 8.2e-19
C3937 P.n1733 VSUBS 0.0155f
C3938 P.n1734 VSUBS 5.99e-19
C3939 P.n1735 VSUBS 5.99e-19
C3940 P.n1736 VSUBS 0.00118f
C3941 P.n1737 VSUBS 5.82e-19
C3942 P.n1738 VSUBS 0.00116f
C3943 P.n1739 VSUBS 0.00116f
C3944 P.n1740 VSUBS 0.0156f
C3945 P.n1741 VSUBS 5.99e-19
C3946 P.n1742 VSUBS 0.00118f
C3947 P.n1743 VSUBS 7.92e-19
C3948 P.n1744 VSUBS 5.82e-19
C3949 P.n1745 VSUBS 0.00116f
C3950 P.n1746 VSUBS 0.00157f
C3951 P.n1747 VSUBS 0.00198f
C3952 P.n1748 VSUBS 0.00608f
C3953 P.n1749 VSUBS 0.00519f
C3954 P.n1750 VSUBS 0.00116f
C3955 P.n1751 VSUBS 0.00109f
C3956 P.n1752 VSUBS 2.73e-19
C3957 P.n1753 VSUBS 0.00116f
C3958 P.n1754 VSUBS 0.00123f
C3959 P.n1755 VSUBS 0.0158f
C3960 P.n1756 VSUBS 5.99e-19
C3961 P.n1757 VSUBS 5.99e-19
C3962 P.n1758 VSUBS 7.86e-19
C3963 P.n1759 VSUBS 0.00124f
C3964 P.n1760 VSUBS 0.00127f
C3965 P.n1761 VSUBS 8.24e-19
C3966 P.n1762 VSUBS 5.99e-19
C3967 P.n1763 VSUBS 5.99e-19
C3968 P.n1764 VSUBS 0.0024f
C3969 P.n1765 VSUBS 0.0024f
C3970 P.n1766 VSUBS 0.00127f
C3971 P.n1767 VSUBS 0.00124f
C3972 P.n1768 VSUBS 1.5e-19
C3973 P.n1769 VSUBS 1.87e-19
C3974 P.n1770 VSUBS 3e-19
C3975 P.n1771 VSUBS 7.49e-19
C3976 P.n1772 VSUBS 7.49e-19
C3977 P.n1773 VSUBS 3.37e-19
C3978 P.n1774 VSUBS 0.0166f
C3979 P.n1775 VSUBS 0.00124f
C3980 P.n1776 VSUBS 0.00124f
C3981 P.n1777 VSUBS 0.00127f
C3982 P.n1778 VSUBS 0.00127f
C3983 P.n1779 VSUBS 0.00314f
C3984 P.n1780 VSUBS 0.00378f
C3985 P.n1781 VSUBS 0.00127f
C3986 P.n1782 VSUBS 3.37e-19
C3987 P.n1783 VSUBS 0.00105f
C3988 P.n1784 VSUBS 9.36e-19
C3989 P.n1785 VSUBS 0.0235f
C3990 P.n1786 VSUBS 3.74e-19
C3991 P.n1787 VSUBS 3.6e-19
C3992 P.n1788 VSUBS 8.98e-19
C3993 P.n1789 VSUBS 9.36e-19
C3994 P.n1790 VSUBS 3.37e-19
C3995 P.n1791 VSUBS 3.37e-19
C3996 P.n1792 VSUBS 8.99e-19
C3997 P.n1793 VSUBS 8.99e-19
C3998 P.n1794 VSUBS 4.87e-19
C3999 P.n1795 VSUBS 0.00337f
C4000 P.n1796 VSUBS 0.00378f
C4001 P.n1797 VSUBS 0.00105f
C4002 P.n1798 VSUBS 5.24e-19
C4003 P.n1799 VSUBS 9.73e-19
C4004 P.n1800 VSUBS 0.00105f
C4005 P.n1801 VSUBS 4.87e-19
C4006 P.n1802 VSUBS 3.37e-19
C4007 P.n1803 VSUBS 3e-19
C4008 P.n1804 VSUBS 8.99e-19
C4009 P.n1805 VSUBS 9.73e-19
C4010 P.n1806 VSUBS 3.74e-19
C4011 P.n1807 VSUBS 3e-19
C4012 P.n1808 VSUBS 3e-19
C4013 P.n1809 VSUBS 7.49e-19
C4014 P.n1810 VSUBS 7.49e-19
C4015 P.n1811 VSUBS 0.00288f
C4016 P.n1812 VSUBS 0.00288f
C4017 P.n1813 VSUBS 3.37e-19
C4018 P.n1814 VSUBS 3.37e-19
C4019 P.n1815 VSUBS 3e-19
C4020 P.n1816 VSUBS 8.99e-19
C4021 P.n1817 VSUBS 0.0223f
C4022 P.n1818 VSUBS 8.99e-19
C4023 P.n1819 VSUBS 3e-19
C4024 P.n1820 VSUBS 3.37e-19
C4025 P.n1821 VSUBS 2.25e-19
C4026 P.n1822 VSUBS 1.5e-19
C4027 P.n1823 VSUBS 8.98e-19
C4028 P.n1824 VSUBS 9.36e-19
C4029 P.n1825 VSUBS 3.37e-19
C4030 P.n1826 VSUBS 3.37e-19
C4031 P.n1827 VSUBS 8.99e-19
C4032 P.n1828 VSUBS 5.01e-19
C4033 P.n1829 VSUBS 1.73e-19
C4034 P.n1830 VSUBS 2.65e-19
C4035 P.n1831 VSUBS 0.022f
C4036 P.n1832 VSUBS 8.99e-19
C4037 P.n1833 VSUBS 3e-19
C4038 P.n1834 VSUBS 3.37e-19
C4039 P.n1835 VSUBS 3.37e-19
C4040 P.n1836 VSUBS 1.87e-19
C4041 P.n1837 VSUBS 1.12e-19
C4042 P.n1838 VSUBS 6.9e-19
C4043 P.n1839 VSUBS 0.00111f
C4044 P.n1840 VSUBS 3.46e-20
C4045 P.n1841 VSUBS 4.1e-19
C4046 P.n1842 VSUBS 0.00247f
C4047 P.n1843 VSUBS 7.49e-19
C4048 P.n1844 VSUBS 7.49e-19
C4049 P.n1845 VSUBS 3e-19
C4050 P.n1846 VSUBS 3e-19
C4051 P.n1847 VSUBS 5.24e-19
C4052 P.n1848 VSUBS 4.49e-19
C4053 P.n1849 VSUBS 5.47e-19
C4054 P.n1850 VSUBS 9.51e-19
C4055 P.n1851 VSUBS 0.0021f
C4056 P.n1852 VSUBS 0.00127f
C4057 P.n1853 VSUBS 0.00127f
C4058 P.n1854 VSUBS 2.99e-19
C4059 P.n1855 VSUBS 1.12e-19
C4060 P.n1857 VSUBS 2.62e-19
C4061 P.n1858 VSUBS 6.74e-19
C4062 P.n1859 VSUBS 7.49e-19
C4063 P.n1860 VSUBS 6.88e-19
C4064 P.n1861 VSUBS 1.73e-19
C4065 P.n1862 VSUBS 2.25e-19
C4066 P.n1863 VSUBS 3.4e-19
C4067 P.n1864 VSUBS 3.46e-20
C4068 P.n1865 VSUBS 0.00116f
C4069 P.n1866 VSUBS 0.016f
C4070 P.n1867 VSUBS 5.99e-19
C4071 P.n1868 VSUBS 7.86e-19
C4072 P.n1869 VSUBS 0.00124f
C4073 P.n1870 VSUBS 0.00127f
C4074 P.n1871 VSUBS 8.24e-19
C4075 P.n1872 VSUBS 5.99e-19
C4076 P.n1873 VSUBS 5.99e-19
C4077 P.n1874 VSUBS 0.0024f
C4078 P.n1875 VSUBS 0.0024f
C4079 P.n1876 VSUBS 0.00127f
C4080 P.n1877 VSUBS 0.00124f
C4081 P.n1878 VSUBS 1.5e-19
C4082 P.n1879 VSUBS 1.87e-19
C4083 P.n1880 VSUBS 3e-19
C4084 P.n1881 VSUBS 7.49e-19
C4085 P.n1882 VSUBS 7.49e-19
C4086 P.n1883 VSUBS 3.37e-19
C4087 P.n1884 VSUBS 0.0174f
C4088 P.n1885 VSUBS 0.00125f
C4089 P.n1886 VSUBS 0.026f
C4090 P.n1887 VSUBS 4.87e-19
C4091 P.n1888 VSUBS 0.00588f
C4092 P.n1889 VSUBS 0.00629f
C4093 P.n1890 VSUBS 0.00105f
C4094 P.n1891 VSUBS 0.00157f
C4095 P.n1892 VSUBS 0.00633f
C4096 P.n1893 VSUBS 0.00565f
C4097 P.n1894 VSUBS 0.0191f
C4098 P.n1895 VSUBS 0.0194f
C4099 P.n1896 VSUBS 0.00105f
C4100 P.n1897 VSUBS 4.87e-19
C4101 P.n1898 VSUBS 0.00588f
C4102 P.n1899 VSUBS 0.00629f
C4103 P.n1900 VSUBS 0.00105f
C4104 P.n1901 VSUBS 0.00157f
C4105 P.n1902 VSUBS 0.0304f
C4106 P.n1903 VSUBS 2.55e-19
C4107 P.n1904 VSUBS 0.00127f
C4108 P.n1905 VSUBS 0.00127f
C4109 P.n1906 VSUBS 0.00314f
C4110 P.n1907 VSUBS 0.00378f
C4111 P.n1908 VSUBS 0.00127f
C4112 P.n1909 VSUBS 3.37e-19
C4113 P.n1910 VSUBS 0.00105f
C4114 P.n1911 VSUBS 9.36e-19
C4115 P.n1912 VSUBS 0.0169f
C4116 P.n1913 VSUBS 0.00105f
C4117 P.n1914 VSUBS 3.74e-19
C4118 P.n1915 VSUBS 3.37e-19
C4119 P.n1916 VSUBS 8.98e-19
C4120 P.n1917 VSUBS 9.36e-19
C4121 P.n1918 VSUBS 3.37e-19
C4122 P.n1919 VSUBS 3.37e-19
C4123 P.n1920 VSUBS 8.99e-19
C4124 P.n1921 VSUBS 8.99e-19
C4125 P.n1922 VSUBS 4.87e-19
C4126 P.n1923 VSUBS 0.00337f
C4127 P.n1924 VSUBS 0.00378f
C4128 P.n1925 VSUBS 0.00105f
C4129 P.n1926 VSUBS 5.24e-19
C4130 P.n1927 VSUBS 9.73e-19
C4131 P.n1928 VSUBS 0.00105f
C4132 P.n1929 VSUBS 4.87e-19
C4133 P.n1930 VSUBS 3.37e-19
C4134 P.n1931 VSUBS 3e-19
C4135 P.n1932 VSUBS 8.99e-19
C4136 P.n1933 VSUBS 9.73e-19
C4137 P.n1934 VSUBS 3.74e-19
C4138 P.n1935 VSUBS 3e-19
C4139 P.n1936 VSUBS 3e-19
C4140 P.n1937 VSUBS 7.49e-19
C4141 P.n1938 VSUBS 7.49e-19
C4142 P.n1939 VSUBS 0.00288f
C4143 P.n1940 VSUBS 0.00288f
C4144 P.n1941 VSUBS 3.37e-19
C4145 P.n1942 VSUBS 3.37e-19
C4146 P.n1943 VSUBS 3e-19
C4147 P.n1944 VSUBS 8.99e-19
C4148 P.n1945 VSUBS 0.0158f
C4149 P.n1946 VSUBS 8.99e-19
C4150 P.n1947 VSUBS 8.99e-19
C4151 P.n1948 VSUBS 3e-19
C4152 P.n1949 VSUBS 3.37e-19
C4153 P.n1950 VSUBS 2.25e-19
C4154 P.n1951 VSUBS 1.5e-19
C4155 P.n1952 VSUBS 8.98e-19
C4156 P.n1953 VSUBS 9.36e-19
C4157 P.n1954 VSUBS 3.37e-19
C4158 P.n1955 VSUBS 3.37e-19
C4159 P.n1956 VSUBS 8.99e-19
C4160 P.n1957 VSUBS 5.01e-19
C4161 P.n1958 VSUBS 1.73e-19
C4162 P.n1959 VSUBS 2.65e-19
C4163 P.n1960 VSUBS 0.0154f
C4164 P.n1961 VSUBS 8.99e-19
C4165 P.n1962 VSUBS 8.99e-19
C4166 P.n1963 VSUBS 3e-19
C4167 P.n1964 VSUBS 3.37e-19
C4168 P.n1965 VSUBS 3.37e-19
C4169 P.n1966 VSUBS 1.87e-19
C4170 P.n1967 VSUBS 1.12e-19
C4171 P.n1968 VSUBS 6.9e-19
C4172 P.n1969 VSUBS 0.00111f
C4173 P.n1970 VSUBS 3.46e-20
C4174 P.n1971 VSUBS 0.00109f
C4175 P.n1972 VSUBS 7.92e-19
C4176 P.n1973 VSUBS 0.00198f
C4177 P.n1974 VSUBS 5.99e-19
C4178 P.n1975 VSUBS 5.99e-19
C4179 P.n1976 VSUBS 9.73e-19
C4180 P.n1977 VSUBS 8.99e-19
C4181 P.n1978 VSUBS 4.06e-19
C4182 P.n1979 VSUBS 2.73e-19
C4183 P.n1980 VSUBS 0.0021f
C4184 P.n1981 VSUBS 0.00127f
C4185 P.n1982 VSUBS 0.00127f
C4186 P.n1983 VSUBS 2.99e-19
C4187 P.n1984 VSUBS 1.12e-19
C4188 P.n1986 VSUBS 2.62e-19
C4189 P.n1987 VSUBS 6.74e-19
C4190 P.n1988 VSUBS 7.49e-19
C4191 P.n1989 VSUBS 6.88e-19
C4192 P.n1990 VSUBS 1.73e-19
C4193 P.n1991 VSUBS 2.25e-19
C4194 P.n1992 VSUBS 3.4e-19
C4195 P.n1993 VSUBS 0.00247f
C4196 P.n1994 VSUBS 7.49e-19
C4197 P.n1995 VSUBS 7.49e-19
C4198 P.n1996 VSUBS 3e-19
C4199 P.n1997 VSUBS 3e-19
C4200 P.n1998 VSUBS 5.24e-19
C4201 P.n1999 VSUBS 4.49e-19
C4202 P.n2000 VSUBS 5.47e-19
C4203 P.n2001 VSUBS 9.51e-19
C4204 P.n2002 VSUBS 3.46e-20
C4205 P.n2003 VSUBS 0.00116f
C4206 P.n2004 VSUBS 0.00198f
C4207 P.n2005 VSUBS 5.99e-19
C4208 P.n2006 VSUBS 5.99e-19
C4209 P.n2007 VSUBS 9.73e-19
C4210 P.n2008 VSUBS 8.99e-19
C4211 P.n2009 VSUBS 4.06e-19
C4212 P.n2010 VSUBS 0.0013f
C4213 P.n2011 VSUBS 4.78e-19
C4214 P.n2012 VSUBS 0.00116f
C4215 P.n2013 VSUBS 0.00109f
C4216 P.n2014 VSUBS 2.73e-19
C4217 P.n2015 VSUBS 0.00116f
C4218 P.n2016 VSUBS 0.246f
C4219 P.t13 VSUBS 2.64f
C4220 P.t121 VSUBS 2.64f
C4221 P.t62 VSUBS 2.64f
C4222 P.t116 VSUBS 2.64f
C4223 P.t109 VSUBS 2.64f
C4224 P.t128 VSUBS 2.64f
C4225 P.t46 VSUBS 2.64f
C4226 P.t77 VSUBS 2.64f
C4227 P.t130 VSUBS 2.64f
C4228 P.t123 VSUBS 2.64f
C4229 P.t12 VSUBS 2.64f
C4230 P.t64 VSUBS 2.78f
C4231 P.n2017 VSUBS 4.87f
C4232 P.n2018 VSUBS 2.51f
C4233 P.n2019 VSUBS 2.51f
C4234 P.n2020 VSUBS 2.51f
C4235 P.n2021 VSUBS 2.51f
C4236 P.n2022 VSUBS 2.51f
C4237 P.n2023 VSUBS 2.51f
C4238 P.n2024 VSUBS 2.51f
C4239 P.n2025 VSUBS 2.51f
C4240 P.n2026 VSUBS 2.51f
C4241 P.n2027 VSUBS 2.18f
C4242 P.n2028 VSUBS 0.0025f
C4243 P.n2029 VSUBS 3.26e-19
C4244 P.n2030 VSUBS 2.17e-19
C4245 P.n2031 VSUBS 2.53e-19
C4246 P.n2032 VSUBS 2.53e-19
C4247 P.n2033 VSUBS 7.6e-19
C4248 P.n2034 VSUBS 9.39e-19
C4249 P.n2035 VSUBS 1.1e-19
C4250 P.n2036 VSUBS 0.0134f
C4251 P.n2037 VSUBS 5.79e-19
C4252 P.n2038 VSUBS 5.79e-19
C4253 P.n2039 VSUBS 7.6e-19
C4254 P.n2040 VSUBS 0.00119f
C4255 P.n2041 VSUBS 0.00123f
C4256 P.n2042 VSUBS 7.96e-19
C4257 P.n2043 VSUBS 5.79e-19
C4258 P.n2044 VSUBS 5.79e-19
C4259 P.n2045 VSUBS 0.00232f
C4260 P.n2046 VSUBS 0.00232f
C4261 P.n2047 VSUBS 0.00123f
C4262 P.n2048 VSUBS 0.00119f
C4263 P.n2049 VSUBS 1.45e-19
C4264 P.n2050 VSUBS 1.81e-19
C4265 P.n2051 VSUBS 2.9e-19
C4266 P.n2052 VSUBS 7.24e-19
C4267 P.n2053 VSUBS 7.24e-19
C4268 P.n2054 VSUBS 3.26e-19
C4269 P.n2055 VSUBS 0.0141f
C4270 P.n2056 VSUBS 0.00119f
C4271 P.n2057 VSUBS 0.00119f
C4272 P.n2058 VSUBS 0.00123f
C4273 P.n2059 VSUBS 0.00123f
C4274 P.n2060 VSUBS 0.00304f
C4275 P.n2061 VSUBS 0.00366f
C4276 P.n2062 VSUBS 0.00123f
C4277 P.n2063 VSUBS 3.26e-19
C4278 P.n2064 VSUBS 0.00101f
C4279 P.n2065 VSUBS 9.05e-19
C4280 P.n2066 VSUBS 0.0198f
C4281 P.n2067 VSUBS 3.62e-19
C4282 P.n2068 VSUBS 3.46e-19
C4283 P.n2069 VSUBS 8.68e-19
C4284 P.n2070 VSUBS 9.05e-19
C4285 P.n2071 VSUBS 3.26e-19
C4286 P.n2072 VSUBS 3.26e-19
C4287 P.n2073 VSUBS 8.69e-19
C4288 P.n2074 VSUBS 8.69e-19
C4289 P.n2075 VSUBS 4.7e-19
C4290 P.n2076 VSUBS 0.00326f
C4291 P.n2077 VSUBS 0.00366f
C4292 P.n2078 VSUBS 0.00101f
C4293 P.n2079 VSUBS 5.07e-19
C4294 P.n2080 VSUBS 9.41e-19
C4295 P.n2081 VSUBS 0.00101f
C4296 P.n2082 VSUBS 4.7e-19
C4297 P.n2083 VSUBS 3.26e-19
C4298 P.n2084 VSUBS 2.9e-19
C4299 P.n2085 VSUBS 8.69e-19
C4300 P.n2086 VSUBS 9.41e-19
C4301 P.n2087 VSUBS 3.62e-19
C4302 P.n2088 VSUBS 2.9e-19
C4303 P.n2089 VSUBS 2.9e-19
C4304 P.n2090 VSUBS 7.24e-19
C4305 P.n2091 VSUBS 7.24e-19
C4306 P.n2092 VSUBS 0.00279f
C4307 P.n2093 VSUBS 0.00279f
C4308 P.n2094 VSUBS 3.26e-19
C4309 P.n2095 VSUBS 3.26e-19
C4310 P.n2096 VSUBS 2.9e-19
C4311 P.n2097 VSUBS 8.69e-19
C4312 P.n2098 VSUBS 0.0186f
C4313 P.n2099 VSUBS 8.69e-19
C4314 P.n2100 VSUBS 2.9e-19
C4315 P.n2101 VSUBS 3.26e-19
C4316 P.n2102 VSUBS 2.17e-19
C4317 P.n2103 VSUBS 1.45e-19
C4318 P.n2104 VSUBS 8.68e-19
C4319 P.n2105 VSUBS 9.05e-19
C4320 P.n2106 VSUBS 3.26e-19
C4321 P.n2107 VSUBS 3.26e-19
C4322 P.n2108 VSUBS 8.69e-19
C4323 P.n2109 VSUBS 4.82e-19
C4324 P.n2110 VSUBS 1.69e-19
C4325 P.n2111 VSUBS 2.55e-19
C4326 P.n2112 VSUBS 3.42e-20
C4327 P.n2113 VSUBS 0.00107f
C4328 P.n2114 VSUBS 0.0183f
C4329 P.n2115 VSUBS 8.69e-19
C4330 P.n2116 VSUBS 2.9e-19
C4331 P.n2117 VSUBS 3.26e-19
C4332 P.n2118 VSUBS 3.26e-19
C4333 P.n2119 VSUBS 1.81e-19
C4334 P.n2120 VSUBS 1.09e-19
C4335 P.n2121 VSUBS 6.71e-19
C4336 P.n2122 VSUBS 3.42e-20
C4337 P.n2123 VSUBS 0.00107f
C4338 P.n2124 VSUBS 0.013f
C4339 P.n2125 VSUBS 8.69e-19
C4340 P.n2126 VSUBS 8.69e-19
C4341 P.n2127 VSUBS 2.9e-19
C4342 P.n2128 VSUBS 3.26e-19
C4343 P.n2129 VSUBS 3.26e-19
C4344 P.n2130 VSUBS 1.81e-19
C4345 P.n2131 VSUBS 1.09e-19
C4346 P.n2132 VSUBS 6.71e-19
C4347 P.n2133 VSUBS 6.63e-19
C4348 P.n2134 VSUBS 1.69e-19
C4349 P.n2135 VSUBS 2.17e-19
C4350 P.n2136 VSUBS 3.28e-19
C4351 P.n2137 VSUBS 3.42e-20
C4352 P.n2138 VSUBS 9.15e-19
C4353 P.n2139 VSUBS 0.00239f
C4354 P.n2140 VSUBS 7.24e-19
C4355 P.n2141 VSUBS 7.24e-19
C4356 P.n2142 VSUBS 2.9e-19
C4357 P.n2143 VSUBS 2.9e-19
C4358 P.n2144 VSUBS 5.07e-19
C4359 P.n2145 VSUBS 4.34e-19
C4360 P.n2146 VSUBS 5.32e-19
C4361 P.n2147 VSUBS 6.63e-19
C4362 P.n2148 VSUBS 1.69e-19
C4363 P.n2149 VSUBS 2.17e-19
C4364 P.n2150 VSUBS 3.28e-19
C4365 P.n2151 VSUBS 3.42e-20
C4366 P.n2152 VSUBS 9.15e-19
C4367 P.n2153 VSUBS 0.00239f
C4368 P.n2154 VSUBS 7.24e-19
C4369 P.n2155 VSUBS 7.24e-19
C4370 P.n2156 VSUBS 2.9e-19
C4371 P.n2157 VSUBS 2.9e-19
C4372 P.n2158 VSUBS 5.07e-19
C4373 P.n2159 VSUBS 4.34e-19
C4374 P.n2160 VSUBS 5.32e-19
C4375 P.n2161 VSUBS 7.24e-19
C4376 P.n2162 VSUBS 6.51e-19
C4377 P.n2163 VSUBS 2.53e-19
C4378 P.n2164 VSUBS 0.00192f
C4379 P.n2165 VSUBS 0.00203f
C4380 P.n2166 VSUBS 0.00123f
C4381 P.n2167 VSUBS 0.00123f
C4382 P.n2168 VSUBS 2.89e-19
C4383 P.n2169 VSUBS 1.09e-19
C4384 P.n2171 VSUBS 0.00192f
C4385 P.n2172 VSUBS 0.00203f
C4386 P.n2173 VSUBS 0.00123f
C4387 P.n2174 VSUBS 0.00123f
C4388 P.n2175 VSUBS 2.89e-19
C4389 P.n2176 VSUBS 1.09e-19
C4390 P.n2177 VSUBS 7.24e-19
C4391 P.n2178 VSUBS 6.51e-19
C4392 P.n2179 VSUBS 2.53e-19
C4393 P.n2181 VSUBS 0.0131f
C4394 P.n2182 VSUBS 5.79e-19
C4395 P.n2183 VSUBS 5.79e-19
C4396 P.n2184 VSUBS 0.00113f
C4397 P.n2185 VSUBS 5.79e-19
C4398 P.n2186 VSUBS 5.79e-19
C4399 P.n2187 VSUBS 9.41e-19
C4400 P.n2188 VSUBS 8.69e-19
C4401 P.n2189 VSUBS 3.96e-19
C4402 P.n2190 VSUBS 7.62e-19
C4403 P.n2191 VSUBS 5.67e-19
C4404 P.t60 VSUBS 2.64f
C4405 P.t67 VSUBS 2.64f
C4406 P.t117 VSUBS 2.64f
C4407 P.t39 VSUBS 2.64f
C4408 P.t32 VSUBS 2.64f
C4409 P.t48 VSUBS 2.64f
C4410 P.t107 VSUBS 2.64f
C4411 P.t124 VSUBS 2.64f
C4412 P.t49 VSUBS 2.64f
C4413 P.t43 VSUBS 2.64f
C4414 P.t71 VSUBS 2.64f
C4415 P.t119 VSUBS 2.78f
C4416 P.n2192 VSUBS 4.87f
C4417 P.n2193 VSUBS 2.51f
C4418 P.n2194 VSUBS 2.51f
C4419 P.n2195 VSUBS 2.51f
C4420 P.n2196 VSUBS 2.51f
C4421 P.n2197 VSUBS 2.51f
C4422 P.n2198 VSUBS 2.51f
C4423 P.n2199 VSUBS 2.51f
C4424 P.n2200 VSUBS 2.51f
C4425 P.n2201 VSUBS 2.51f
C4426 P.n2202 VSUBS 2.18f
C4427 P.n2203 VSUBS 0.0164f
C4428 P.n2204 VSUBS 8.69e-19
C4429 P.n2205 VSUBS 8.69e-19
C4430 P.n2206 VSUBS 2.9e-19
C4431 P.n2207 VSUBS 3.26e-19
C4432 P.n2208 VSUBS 3.26e-19
C4433 P.n2209 VSUBS 1.81e-19
C4434 P.n2210 VSUBS 1.09e-19
C4435 P.n2211 VSUBS 6.71e-19
C4436 P.n2212 VSUBS 0.0154f
C4437 P.n2213 VSUBS 8.69e-19
C4438 P.n2214 VSUBS 2.9e-19
C4439 P.n2215 VSUBS 3.26e-19
C4440 P.n2216 VSUBS 3.26e-19
C4441 P.n2217 VSUBS 1.81e-19
C4442 P.n2218 VSUBS 1.09e-19
C4443 P.n2219 VSUBS 6.71e-19
C4444 P.n2220 VSUBS 0.00239f
C4445 P.n2221 VSUBS 7.24e-19
C4446 P.n2222 VSUBS 7.24e-19
C4447 P.n2223 VSUBS 2.9e-19
C4448 P.n2224 VSUBS 2.9e-19
C4449 P.n2225 VSUBS 5.07e-19
C4450 P.n2226 VSUBS 4.34e-19
C4451 P.n2227 VSUBS 1.69e-19
C4452 P.n2228 VSUBS 2.17e-19
C4453 P.n2229 VSUBS 3.28e-19
C4454 P.n2230 VSUBS 3.42e-20
C4455 P.n2231 VSUBS 9.15e-19
C4456 P.n2232 VSUBS 5.32e-19
C4457 P.n2233 VSUBS 0.00239f
C4458 P.n2234 VSUBS 7.24e-19
C4459 P.n2235 VSUBS 7.24e-19
C4460 P.n2236 VSUBS 2.9e-19
C4461 P.n2237 VSUBS 2.9e-19
C4462 P.n2238 VSUBS 5.07e-19
C4463 P.n2239 VSUBS 4.34e-19
C4464 P.n2240 VSUBS 1.69e-19
C4465 P.n2241 VSUBS 2.17e-19
C4466 P.n2242 VSUBS 3.28e-19
C4467 P.n2243 VSUBS 3.42e-20
C4468 P.n2244 VSUBS 9.15e-19
C4469 P.n2245 VSUBS 5.32e-19
C4470 P.n2246 VSUBS 0.0025f
C4471 P.n2247 VSUBS 3.26e-19
C4472 P.n2248 VSUBS 2.17e-19
C4473 P.n2249 VSUBS 2.53e-19
C4474 P.n2250 VSUBS 2.53e-19
C4475 P.n2251 VSUBS 7.6e-19
C4476 P.n2252 VSUBS 9.39e-19
C4477 P.n2253 VSUBS 1.1e-19
C4478 P.n2254 VSUBS 0.00702f
C4479 P.n2255 VSUBS 5.79e-19
C4480 P.n2256 VSUBS 7.6e-19
C4481 P.n2257 VSUBS 0.00119f
C4482 P.n2258 VSUBS 0.00123f
C4483 P.n2259 VSUBS 7.96e-19
C4484 P.n2260 VSUBS 5.79e-19
C4485 P.n2261 VSUBS 5.79e-19
C4486 P.n2262 VSUBS 0.00232f
C4487 P.n2263 VSUBS 0.00232f
C4488 P.n2264 VSUBS 0.00123f
C4489 P.n2265 VSUBS 0.00119f
C4490 P.n2266 VSUBS 1.45e-19
C4491 P.n2267 VSUBS 1.81e-19
C4492 P.n2268 VSUBS 2.9e-19
C4493 P.n2269 VSUBS 7.24e-19
C4494 P.n2270 VSUBS 7.24e-19
C4495 P.n2271 VSUBS 3.26e-19
C4496 P.n2272 VSUBS 0.00836f
C4497 P.n2273 VSUBS 0.0012f
C4498 P.n2274 VSUBS 0.0193f
C4499 P.n2275 VSUBS 4.7e-19
C4500 P.n2276 VSUBS 0.00568f
C4501 P.n2277 VSUBS 0.00608f
C4502 P.n2278 VSUBS 0.00101f
C4503 P.n2279 VSUBS 0.00152f
C4504 P.n2280 VSUBS 0.00612f
C4505 P.n2281 VSUBS 0.00546f
C4506 P.n2282 VSUBS 0.0199f
C4507 P.n2283 VSUBS 0.0202f
C4508 P.n2284 VSUBS 0.00101f
C4509 P.n2285 VSUBS 4.7e-19
C4510 P.n2286 VSUBS 0.00568f
C4511 P.n2287 VSUBS 0.00608f
C4512 P.n2288 VSUBS 0.00101f
C4513 P.n2289 VSUBS 0.00152f
C4514 P.n2290 VSUBS 0.021f
C4515 P.n2291 VSUBS 1.63e-19
C4516 P.n2292 VSUBS 0.00123f
C4517 P.n2293 VSUBS 0.00123f
C4518 P.n2294 VSUBS 0.00304f
C4519 P.n2295 VSUBS 0.00366f
C4520 P.n2296 VSUBS 0.00123f
C4521 P.n2297 VSUBS 3.26e-19
C4522 P.n2298 VSUBS 0.00101f
C4523 P.n2299 VSUBS 9.05e-19
C4524 P.n2300 VSUBS 0.0178f
C4525 P.n2301 VSUBS 0.00101f
C4526 P.n2302 VSUBS 3.62e-19
C4527 P.n2303 VSUBS 3.26e-19
C4528 P.n2304 VSUBS 8.68e-19
C4529 P.n2305 VSUBS 9.05e-19
C4530 P.n2306 VSUBS 3.26e-19
C4531 P.n2307 VSUBS 3.26e-19
C4532 P.n2308 VSUBS 8.69e-19
C4533 P.n2309 VSUBS 8.69e-19
C4534 P.n2310 VSUBS 4.7e-19
C4535 P.n2311 VSUBS 0.00326f
C4536 P.n2312 VSUBS 0.00366f
C4537 P.n2313 VSUBS 0.00101f
C4538 P.n2314 VSUBS 5.07e-19
C4539 P.n2315 VSUBS 9.41e-19
C4540 P.n2316 VSUBS 0.00101f
C4541 P.n2317 VSUBS 4.7e-19
C4542 P.n2318 VSUBS 3.26e-19
C4543 P.n2319 VSUBS 2.9e-19
C4544 P.n2320 VSUBS 8.69e-19
C4545 P.n2321 VSUBS 9.41e-19
C4546 P.n2322 VSUBS 3.62e-19
C4547 P.n2323 VSUBS 2.9e-19
C4548 P.n2324 VSUBS 2.9e-19
C4549 P.n2325 VSUBS 7.24e-19
C4550 P.n2326 VSUBS 7.24e-19
C4551 P.n2327 VSUBS 0.00279f
C4552 P.n2328 VSUBS 0.00279f
C4553 P.n2329 VSUBS 3.26e-19
C4554 P.n2330 VSUBS 3.26e-19
C4555 P.n2331 VSUBS 2.9e-19
C4556 P.n2332 VSUBS 8.69e-19
C4557 P.n2333 VSUBS 0.0168f
C4558 P.n2334 VSUBS 8.69e-19
C4559 P.n2335 VSUBS 8.69e-19
C4560 P.n2336 VSUBS 2.9e-19
C4561 P.n2337 VSUBS 3.26e-19
C4562 P.n2338 VSUBS 2.17e-19
C4563 P.n2339 VSUBS 1.45e-19
C4564 P.n2340 VSUBS 8.68e-19
C4565 P.n2341 VSUBS 9.05e-19
C4566 P.n2342 VSUBS 3.26e-19
C4567 P.n2343 VSUBS 3.26e-19
C4568 P.n2344 VSUBS 8.69e-19
C4569 P.n2345 VSUBS 4.82e-19
C4570 P.n2346 VSUBS 0.00107f
C4571 P.n2347 VSUBS 3.42e-20
C4572 P.n2348 VSUBS 2.55e-19
C4573 P.n2349 VSUBS 1.69e-19
C4574 P.n2350 VSUBS 0.00107f
C4575 P.n2351 VSUBS 3.42e-20
C4576 P.n2352 VSUBS 2.55e-19
C4577 P.n2353 VSUBS 0.0025f
C4578 P.n2354 VSUBS 3.26e-19
C4579 P.n2355 VSUBS 2.17e-19
C4580 P.n2356 VSUBS 2.53e-19
C4581 P.n2357 VSUBS 2.53e-19
C4582 P.n2358 VSUBS 7.6e-19
C4583 P.n2359 VSUBS 9.39e-19
C4584 P.n2360 VSUBS 1.1e-19
C4585 P.n2361 VSUBS 0.0168f
C4586 P.n2362 VSUBS 5.79e-19
C4587 P.n2363 VSUBS 5.79e-19
C4588 P.n2364 VSUBS 7.6e-19
C4589 P.n2365 VSUBS 0.00119f
C4590 P.n2366 VSUBS 0.00123f
C4591 P.n2367 VSUBS 7.96e-19
C4592 P.n2368 VSUBS 5.79e-19
C4593 P.n2369 VSUBS 5.79e-19
C4594 P.n2370 VSUBS 0.00232f
C4595 P.n2371 VSUBS 0.00232f
C4596 P.n2372 VSUBS 0.00123f
C4597 P.n2373 VSUBS 0.00119f
C4598 P.n2374 VSUBS 1.45e-19
C4599 P.n2375 VSUBS 1.81e-19
C4600 P.n2376 VSUBS 2.9e-19
C4601 P.n2377 VSUBS 7.24e-19
C4602 P.n2378 VSUBS 7.24e-19
C4603 P.n2379 VSUBS 3.26e-19
C4604 P.n2380 VSUBS 0.0175f
C4605 P.n2381 VSUBS 0.00119f
C4606 P.n2382 VSUBS 0.00119f
C4607 P.n2383 VSUBS 0.00123f
C4608 P.n2384 VSUBS 0.00123f
C4609 P.n2385 VSUBS 0.00304f
C4610 P.n2386 VSUBS 0.00366f
C4611 P.n2387 VSUBS 0.00123f
C4612 P.n2388 VSUBS 3.26e-19
C4613 P.n2389 VSUBS 0.00101f
C4614 P.n2390 VSUBS 9.05e-19
C4615 P.n2391 VSUBS 0.0169f
C4616 P.n2392 VSUBS 3.62e-19
C4617 P.n2393 VSUBS 3.44e-19
C4618 P.n2394 VSUBS 8.68e-19
C4619 P.n2395 VSUBS 9.05e-19
C4620 P.n2396 VSUBS 3.26e-19
C4621 P.n2397 VSUBS 3.26e-19
C4622 P.n2398 VSUBS 8.69e-19
C4623 P.n2399 VSUBS 8.69e-19
C4624 P.n2400 VSUBS 4.7e-19
C4625 P.n2401 VSUBS 0.00326f
C4626 P.n2402 VSUBS 0.00366f
C4627 P.n2403 VSUBS 0.00101f
C4628 P.n2404 VSUBS 5.07e-19
C4629 P.n2405 VSUBS 9.41e-19
C4630 P.n2406 VSUBS 0.00101f
C4631 P.n2407 VSUBS 4.7e-19
C4632 P.n2408 VSUBS 3.26e-19
C4633 P.n2409 VSUBS 2.9e-19
C4634 P.n2410 VSUBS 8.69e-19
C4635 P.n2411 VSUBS 9.41e-19
C4636 P.n2412 VSUBS 3.62e-19
C4637 P.n2413 VSUBS 2.9e-19
C4638 P.n2414 VSUBS 2.9e-19
C4639 P.n2415 VSUBS 7.24e-19
C4640 P.n2416 VSUBS 7.24e-19
C4641 P.n2417 VSUBS 0.00279f
C4642 P.n2418 VSUBS 0.00279f
C4643 P.n2419 VSUBS 3.26e-19
C4644 P.n2420 VSUBS 3.26e-19
C4645 P.n2421 VSUBS 2.9e-19
C4646 P.n2422 VSUBS 8.69e-19
C4647 P.n2423 VSUBS 0.0157f
C4648 P.n2424 VSUBS 8.69e-19
C4649 P.n2425 VSUBS 2.9e-19
C4650 P.n2426 VSUBS 3.26e-19
C4651 P.n2427 VSUBS 2.17e-19
C4652 P.n2428 VSUBS 1.45e-19
C4653 P.n2429 VSUBS 8.68e-19
C4654 P.n2430 VSUBS 9.05e-19
C4655 P.n2431 VSUBS 3.26e-19
C4656 P.n2432 VSUBS 3.26e-19
C4657 P.n2433 VSUBS 8.69e-19
C4658 P.n2434 VSUBS 4.82e-19
C4659 P.n2435 VSUBS 1.69e-19
C4660 P.n2436 VSUBS 0.00192f
C4661 P.n2437 VSUBS 0.00203f
C4662 P.n2438 VSUBS 0.00123f
C4663 P.n2439 VSUBS 0.00123f
C4664 P.n2440 VSUBS 2.89e-19
C4665 P.n2441 VSUBS 1.09e-19
C4666 P.n2442 VSUBS 6.63e-19
C4667 P.n2443 VSUBS 7.24e-19
C4668 P.n2444 VSUBS 6.51e-19
C4669 P.n2445 VSUBS 2.53e-19
C4670 P.n2447 VSUBS 7.62e-19
C4671 P.n2448 VSUBS 0.00662f
C4672 P.n2449 VSUBS 5.79e-19
C4673 P.n2450 VSUBS 0.00113f
C4674 P.n2451 VSUBS 5.67e-19
C4675 P.n2452 VSUBS 0.0165f
C4676 P.n2453 VSUBS 5.79e-19
C4677 P.n2454 VSUBS 5.79e-19
C4678 P.n2455 VSUBS 0.00113f
C4679 P.n2456 VSUBS 7.62e-19
C4680 P.n2457 VSUBS 5.67e-19
C4681 P.n2458 VSUBS 5.79e-19
C4682 P.n2459 VSUBS 5.79e-19
C4683 P.n2460 VSUBS 9.41e-19
C4684 P.n2461 VSUBS 8.69e-19
C4685 P.n2462 VSUBS 3.96e-19
C4686 P.n2463 VSUBS 5.79e-19
C4687 P.n2464 VSUBS 5.79e-19
C4688 P.n2465 VSUBS 9.41e-19
C4689 P.n2466 VSUBS 8.69e-19
C4690 P.n2467 VSUBS 3.96e-19
C4691 P.n2468 VSUBS 0.014f
C4692 P.n2469 VSUBS 8.69e-19
C4693 P.n2470 VSUBS 8.69e-19
C4694 P.n2471 VSUBS 2.9e-19
C4695 P.n2472 VSUBS 3.26e-19
C4696 P.n2473 VSUBS 3.26e-19
C4697 P.n2474 VSUBS 1.81e-19
C4698 P.n2475 VSUBS 1.09e-19
C4699 P.n2476 VSUBS 6.71e-19
C4700 P.n2477 VSUBS 0.0181f
C4701 P.n2478 VSUBS 8.69e-19
C4702 P.n2479 VSUBS 2.9e-19
C4703 P.n2480 VSUBS 3.26e-19
C4704 P.n2481 VSUBS 3.26e-19
C4705 P.n2482 VSUBS 1.81e-19
C4706 P.n2483 VSUBS 1.09e-19
C4707 P.n2484 VSUBS 6.71e-19
C4708 P.n2485 VSUBS 1.69e-19
C4709 P.n2486 VSUBS 2.17e-19
C4710 P.n2487 VSUBS 3.28e-19
C4711 P.n2488 VSUBS 3.42e-20
C4712 P.n2489 VSUBS 9.15e-19
C4713 P.n2490 VSUBS 0.00239f
C4714 P.n2491 VSUBS 7.24e-19
C4715 P.n2492 VSUBS 7.24e-19
C4716 P.n2493 VSUBS 2.9e-19
C4717 P.n2494 VSUBS 2.9e-19
C4718 P.n2495 VSUBS 5.07e-19
C4719 P.n2496 VSUBS 4.34e-19
C4720 P.n2497 VSUBS 5.32e-19
C4721 P.n2498 VSUBS 1.69e-19
C4722 P.n2499 VSUBS 2.17e-19
C4723 P.n2500 VSUBS 3.28e-19
C4724 P.n2501 VSUBS 3.42e-20
C4725 P.n2502 VSUBS 9.15e-19
C4726 P.n2503 VSUBS 0.00239f
C4727 P.n2504 VSUBS 7.24e-19
C4728 P.n2505 VSUBS 7.24e-19
C4729 P.n2506 VSUBS 2.9e-19
C4730 P.n2507 VSUBS 2.9e-19
C4731 P.n2508 VSUBS 5.07e-19
C4732 P.n2509 VSUBS 4.34e-19
C4733 P.n2510 VSUBS 5.32e-19
C4734 P.t15 VSUBS 2.64f
C4735 P.t37 VSUBS 2.64f
C4736 P.t34 VSUBS 2.64f
C4737 P.t91 VSUBS 2.64f
C4738 P.t78 VSUBS 2.64f
C4739 P.t102 VSUBS 2.64f
C4740 P.t17 VSUBS 2.64f
C4741 P.t40 VSUBS 2.64f
C4742 P.t104 VSUBS 2.64f
C4743 P.t97 VSUBS 2.64f
C4744 P.t113 VSUBS 2.64f
C4745 P.t36 VSUBS 2.78f
C4746 P.n2511 VSUBS 4.87f
C4747 P.n2512 VSUBS 2.51f
C4748 P.n2513 VSUBS 2.51f
C4749 P.n2514 VSUBS 2.51f
C4750 P.n2515 VSUBS 2.51f
C4751 P.n2516 VSUBS 2.51f
C4752 P.n2517 VSUBS 2.51f
C4753 P.n2518 VSUBS 2.51f
C4754 P.n2519 VSUBS 2.51f
C4755 P.n2520 VSUBS 2.51f
C4756 P.n2521 VSUBS 2.19f
C4757 P.n2522 VSUBS 0.00107f
C4758 P.n2523 VSUBS 3.42e-20
C4759 P.n2524 VSUBS 2.55e-19
C4760 P.n2525 VSUBS 0.0025f
C4761 P.n2526 VSUBS 3.26e-19
C4762 P.n2527 VSUBS 2.17e-19
C4763 P.n2528 VSUBS 2.53e-19
C4764 P.n2529 VSUBS 2.53e-19
C4765 P.n2530 VSUBS 7.6e-19
C4766 P.n2531 VSUBS 9.39e-19
C4767 P.n2532 VSUBS 1.1e-19
C4768 P.n2533 VSUBS 0.00912f
C4769 P.n2534 VSUBS 5.79e-19
C4770 P.n2535 VSUBS 7.6e-19
C4771 P.n2536 VSUBS 0.00119f
C4772 P.n2537 VSUBS 0.00123f
C4773 P.n2538 VSUBS 7.96e-19
C4774 P.n2539 VSUBS 5.79e-19
C4775 P.n2540 VSUBS 5.79e-19
C4776 P.n2541 VSUBS 0.00232f
C4777 P.n2542 VSUBS 0.00232f
C4778 P.n2543 VSUBS 0.00123f
C4779 P.n2544 VSUBS 0.00119f
C4780 P.n2545 VSUBS 1.45e-19
C4781 P.n2546 VSUBS 1.81e-19
C4782 P.n2547 VSUBS 2.9e-19
C4783 P.n2548 VSUBS 7.24e-19
C4784 P.n2549 VSUBS 7.24e-19
C4785 P.n2550 VSUBS 3.26e-19
C4786 P.n2551 VSUBS 0.0105f
C4787 P.n2552 VSUBS 0.0012f
C4788 P.n2553 VSUBS 0.022f
C4789 P.n2554 VSUBS 4.7e-19
C4790 P.n2555 VSUBS 0.00568f
C4791 P.n2556 VSUBS 0.00608f
C4792 P.n2557 VSUBS 0.00101f
C4793 P.n2558 VSUBS 0.00152f
C4794 P.n2559 VSUBS 0.00612f
C4795 P.n2560 VSUBS 0.00546f
C4796 P.n2561 VSUBS 0.0175f
C4797 P.n2562 VSUBS 0.0178f
C4798 P.n2563 VSUBS 0.00101f
C4799 P.n2564 VSUBS 4.7e-19
C4800 P.n2565 VSUBS 0.00568f
C4801 P.n2566 VSUBS 0.00608f
C4802 P.n2567 VSUBS 0.00101f
C4803 P.n2568 VSUBS 0.00152f
C4804 P.n2569 VSUBS 0.023f
C4805 P.n2570 VSUBS 1.85e-19
C4806 P.n2571 VSUBS 0.00123f
C4807 P.n2572 VSUBS 0.00123f
C4808 P.n2573 VSUBS 0.00304f
C4809 P.n2574 VSUBS 0.00366f
C4810 P.n2575 VSUBS 0.00123f
C4811 P.n2576 VSUBS 3.26e-19
C4812 P.n2577 VSUBS 0.00101f
C4813 P.n2578 VSUBS 9.05e-19
C4814 P.n2579 VSUBS 0.0154f
C4815 P.n2580 VSUBS 0.00101f
C4816 P.n2581 VSUBS 3.62e-19
C4817 P.n2582 VSUBS 3.26e-19
C4818 P.n2583 VSUBS 8.68e-19
C4819 P.n2584 VSUBS 9.05e-19
C4820 P.n2585 VSUBS 3.26e-19
C4821 P.n2586 VSUBS 3.26e-19
C4822 P.n2587 VSUBS 8.69e-19
C4823 P.n2588 VSUBS 8.69e-19
C4824 P.n2589 VSUBS 4.7e-19
C4825 P.n2590 VSUBS 0.00326f
C4826 P.n2591 VSUBS 0.00366f
C4827 P.n2592 VSUBS 0.00101f
C4828 P.n2593 VSUBS 5.07e-19
C4829 P.n2594 VSUBS 9.41e-19
C4830 P.n2595 VSUBS 0.00101f
C4831 P.n2596 VSUBS 4.7e-19
C4832 P.n2597 VSUBS 3.26e-19
C4833 P.n2598 VSUBS 2.9e-19
C4834 P.n2599 VSUBS 8.69e-19
C4835 P.n2600 VSUBS 9.41e-19
C4836 P.n2601 VSUBS 3.62e-19
C4837 P.n2602 VSUBS 2.9e-19
C4838 P.n2603 VSUBS 2.9e-19
C4839 P.n2604 VSUBS 7.24e-19
C4840 P.n2605 VSUBS 7.24e-19
C4841 P.n2606 VSUBS 0.00279f
C4842 P.n2607 VSUBS 0.00279f
C4843 P.n2608 VSUBS 3.26e-19
C4844 P.n2609 VSUBS 3.26e-19
C4845 P.n2610 VSUBS 2.9e-19
C4846 P.n2611 VSUBS 8.69e-19
C4847 P.n2612 VSUBS 0.0144f
C4848 P.n2613 VSUBS 8.69e-19
C4849 P.n2614 VSUBS 8.69e-19
C4850 P.n2615 VSUBS 2.9e-19
C4851 P.n2616 VSUBS 3.26e-19
C4852 P.n2617 VSUBS 2.17e-19
C4853 P.n2618 VSUBS 1.45e-19
C4854 P.n2619 VSUBS 8.68e-19
C4855 P.n2620 VSUBS 9.05e-19
C4856 P.n2621 VSUBS 3.26e-19
C4857 P.n2622 VSUBS 3.26e-19
C4858 P.n2623 VSUBS 8.69e-19
C4859 P.n2624 VSUBS 4.82e-19
C4860 P.n2625 VSUBS 1.69e-19
C4861 P.n2626 VSUBS 0.0025f
C4862 P.n2627 VSUBS 3.26e-19
C4863 P.n2628 VSUBS 2.17e-19
C4864 P.n2629 VSUBS 2.53e-19
C4865 P.n2630 VSUBS 2.53e-19
C4866 P.n2631 VSUBS 7.6e-19
C4867 P.n2632 VSUBS 9.39e-19
C4868 P.n2633 VSUBS 1.1e-19
C4869 P.n2634 VSUBS 0.0144f
C4870 P.n2635 VSUBS 5.79e-19
C4871 P.n2636 VSUBS 5.79e-19
C4872 P.n2637 VSUBS 7.6e-19
C4873 P.n2638 VSUBS 0.00119f
C4874 P.n2639 VSUBS 0.00123f
C4875 P.n2640 VSUBS 7.96e-19
C4876 P.n2641 VSUBS 5.79e-19
C4877 P.n2642 VSUBS 5.79e-19
C4878 P.n2643 VSUBS 0.00232f
C4879 P.n2644 VSUBS 0.00232f
C4880 P.n2645 VSUBS 0.00123f
C4881 P.n2646 VSUBS 0.00119f
C4882 P.n2647 VSUBS 1.45e-19
C4883 P.n2648 VSUBS 1.81e-19
C4884 P.n2649 VSUBS 2.9e-19
C4885 P.n2650 VSUBS 7.24e-19
C4886 P.n2651 VSUBS 7.24e-19
C4887 P.n2652 VSUBS 3.26e-19
C4888 P.n2653 VSUBS 0.0151f
C4889 P.n2654 VSUBS 0.00119f
C4890 P.n2655 VSUBS 0.00119f
C4891 P.n2656 VSUBS 0.00123f
C4892 P.n2657 VSUBS 0.00123f
C4893 P.n2658 VSUBS 0.00304f
C4894 P.n2659 VSUBS 0.00366f
C4895 P.n2660 VSUBS 0.00123f
C4896 P.n2661 VSUBS 3.26e-19
C4897 P.n2662 VSUBS 0.00101f
C4898 P.n2663 VSUBS 9.05e-19
C4899 P.n2664 VSUBS 0.0195f
C4900 P.n2665 VSUBS 3.62e-19
C4901 P.n2666 VSUBS 3.46e-19
C4902 P.n2667 VSUBS 8.68e-19
C4903 P.n2668 VSUBS 9.05e-19
C4904 P.n2669 VSUBS 3.26e-19
C4905 P.n2670 VSUBS 3.26e-19
C4906 P.n2671 VSUBS 8.69e-19
C4907 P.n2672 VSUBS 8.69e-19
C4908 P.n2673 VSUBS 4.7e-19
C4909 P.n2674 VSUBS 0.00326f
C4910 P.n2675 VSUBS 0.00366f
C4911 P.n2676 VSUBS 0.00101f
C4912 P.n2677 VSUBS 5.07e-19
C4913 P.n2678 VSUBS 9.41e-19
C4914 P.n2679 VSUBS 0.00101f
C4915 P.n2680 VSUBS 4.7e-19
C4916 P.n2681 VSUBS 3.26e-19
C4917 P.n2682 VSUBS 2.9e-19
C4918 P.n2683 VSUBS 8.69e-19
C4919 P.n2684 VSUBS 9.41e-19
C4920 P.n2685 VSUBS 3.62e-19
C4921 P.n2686 VSUBS 2.9e-19
C4922 P.n2687 VSUBS 2.9e-19
C4923 P.n2688 VSUBS 7.24e-19
C4924 P.n2689 VSUBS 7.24e-19
C4925 P.n2690 VSUBS 0.00279f
C4926 P.n2691 VSUBS 0.00279f
C4927 P.n2692 VSUBS 3.26e-19
C4928 P.n2693 VSUBS 3.26e-19
C4929 P.n2694 VSUBS 2.9e-19
C4930 P.n2695 VSUBS 8.69e-19
C4931 P.n2696 VSUBS 0.0184f
C4932 P.n2697 VSUBS 8.69e-19
C4933 P.n2698 VSUBS 2.9e-19
C4934 P.n2699 VSUBS 3.26e-19
C4935 P.n2700 VSUBS 2.17e-19
C4936 P.n2701 VSUBS 1.45e-19
C4937 P.n2702 VSUBS 8.68e-19
C4938 P.n2703 VSUBS 9.05e-19
C4939 P.n2704 VSUBS 3.26e-19
C4940 P.n2705 VSUBS 3.26e-19
C4941 P.n2706 VSUBS 8.69e-19
C4942 P.n2707 VSUBS 4.82e-19
C4943 P.n2708 VSUBS 0.00107f
C4944 P.n2709 VSUBS 3.42e-20
C4945 P.n2710 VSUBS 2.55e-19
C4946 P.n2711 VSUBS 1.69e-19
C4947 P.n2712 VSUBS 6.63e-19
C4948 P.n2713 VSUBS 7.24e-19
C4949 P.n2714 VSUBS 6.51e-19
C4950 P.n2715 VSUBS 2.53e-19
C4951 P.n2716 VSUBS 0.00192f
C4952 P.n2717 VSUBS 0.00203f
C4953 P.n2718 VSUBS 0.00123f
C4954 P.n2719 VSUBS 0.00123f
C4955 P.n2720 VSUBS 2.89e-19
C4956 P.n2721 VSUBS 1.09e-19
C4957 P.n2723 VSUBS 5.79e-19
C4958 P.n2724 VSUBS 5.79e-19
C4959 P.n2725 VSUBS 9.41e-19
C4960 P.n2726 VSUBS 8.69e-19
C4961 P.n2727 VSUBS 3.96e-19
C4962 P.n2728 VSUBS 7.62e-19
C4963 P.n2729 VSUBS 0.00872f
C4964 P.n2730 VSUBS 5.79e-19
C4965 P.n2731 VSUBS 0.00113f
C4966 P.n2732 VSUBS 5.67e-19
C4967 P.n2733 VSUBS 5.79e-19
C4968 P.n2734 VSUBS 5.79e-19
C4969 P.n2735 VSUBS 9.41e-19
C4970 P.n2736 VSUBS 8.69e-19
C4971 P.n2737 VSUBS 3.96e-19
C4972 P.n2738 VSUBS 7.62e-19
C4973 P.n2739 VSUBS 0.0141f
C4974 P.n2740 VSUBS 5.79e-19
C4975 P.n2741 VSUBS 5.79e-19
C4976 P.n2742 VSUBS 0.00113f
C4977 P.n2743 VSUBS 5.67e-19
C4978 P.n2744 VSUBS 3.42e-20
C4979 P.n2745 VSUBS 8.69e-19
C4980 P.n2746 VSUBS 8.69e-19
C4981 P.n2747 VSUBS 0.02f
C4982 P.n2748 VSUBS 8.69e-19
C4983 P.n2749 VSUBS 2.9e-19
C4984 P.n2750 VSUBS 3.26e-19
C4985 P.n2751 VSUBS 3.26e-19
C4986 P.n2752 VSUBS 1.81e-19
C4987 P.n2753 VSUBS 1.09e-19
C4988 P.n2754 VSUBS 0.00239f
C4989 P.n2755 VSUBS 7.24e-19
C4990 P.n2756 VSUBS 7.24e-19
C4991 P.n2757 VSUBS 2.9e-19
C4992 P.n2758 VSUBS 2.9e-19
C4993 P.n2759 VSUBS 5.07e-19
C4994 P.n2760 VSUBS 4.34e-19
C4995 P.n2761 VSUBS 6.63e-19
C4996 P.n2762 VSUBS 1.69e-19
C4997 P.n2763 VSUBS 2.17e-19
C4998 P.n2764 VSUBS 3.28e-19
C4999 P.n2765 VSUBS 3.42e-20
C5000 P.n2766 VSUBS 9.15e-19
C5001 P.n2767 VSUBS 5.32e-19
C5002 P.n2768 VSUBS 0.00239f
C5003 P.n2769 VSUBS 7.24e-19
C5004 P.n2770 VSUBS 7.24e-19
C5005 P.n2771 VSUBS 2.9e-19
C5006 P.n2772 VSUBS 2.9e-19
C5007 P.n2773 VSUBS 5.07e-19
C5008 P.n2774 VSUBS 4.34e-19
C5009 P.n2775 VSUBS 6.63e-19
C5010 P.n2776 VSUBS 1.69e-19
C5011 P.n2777 VSUBS 2.17e-19
C5012 P.n2778 VSUBS 3.28e-19
C5013 P.n2779 VSUBS 3.42e-20
C5014 P.n2780 VSUBS 9.15e-19
C5015 P.n2781 VSUBS 5.32e-19
C5016 P.t9 VSUBS 2.64f
C5017 P.t87 VSUBS 2.64f
C5018 P.t16 VSUBS 2.64f
C5019 P.t72 VSUBS 2.64f
C5020 P.t56 VSUBS 2.64f
C5021 P.t90 VSUBS 2.64f
C5022 P.t1 VSUBS 2.64f
C5023 P.t29 VSUBS 2.64f
C5024 P.t92 VSUBS 2.64f
C5025 P.t80 VSUBS 2.64f
C5026 P.t103 VSUBS 2.64f
C5027 P.t18 VSUBS 2.78f
C5028 P.n2782 VSUBS 4.87f
C5029 P.n2783 VSUBS 2.51f
C5030 P.n2784 VSUBS 2.51f
C5031 P.n2785 VSUBS 2.51f
C5032 P.n2786 VSUBS 2.51f
C5033 P.n2787 VSUBS 2.51f
C5034 P.n2788 VSUBS 2.51f
C5035 P.n2789 VSUBS 2.51f
C5036 P.n2790 VSUBS 2.51f
C5037 P.n2791 VSUBS 2.51f
C5038 P.n2792 VSUBS 2.18f
C5039 P.n2793 VSUBS 0.00192f
C5040 P.n2794 VSUBS 0.00203f
C5041 P.n2795 VSUBS 0.00123f
C5042 P.n2796 VSUBS 0.00123f
C5043 P.n2797 VSUBS 2.89e-19
C5044 P.n2798 VSUBS 1.09e-19
C5045 P.n2799 VSUBS 7.24e-19
C5046 P.n2800 VSUBS 6.51e-19
C5047 P.n2801 VSUBS 2.53e-19
C5048 P.n2802 VSUBS 7.24e-19
C5049 P.n2803 VSUBS 6.51e-19
C5050 P.n2804 VSUBS 2.53e-19
C5051 P.n2805 VSUBS 0.00192f
C5052 P.n2806 VSUBS 0.00203f
C5053 P.n2807 VSUBS 0.00123f
C5054 P.n2808 VSUBS 0.00123f
C5055 P.n2809 VSUBS 2.89e-19
C5056 P.n2810 VSUBS 1.09e-19
C5057 P.n2812 VSUBS 0.0025f
C5058 P.n2813 VSUBS 3.26e-19
C5059 P.n2814 VSUBS 2.17e-19
C5060 P.n2815 VSUBS 2.53e-19
C5061 P.n2816 VSUBS 2.53e-19
C5062 P.n2817 VSUBS 7.6e-19
C5063 P.n2818 VSUBS 9.39e-19
C5064 P.n2819 VSUBS 1.1e-19
C5065 P.n2820 VSUBS 0.00615f
C5066 P.n2821 VSUBS 5.79e-19
C5067 P.n2822 VSUBS 7.6e-19
C5068 P.n2823 VSUBS 0.00119f
C5069 P.n2824 VSUBS 0.00123f
C5070 P.n2825 VSUBS 7.96e-19
C5071 P.n2826 VSUBS 5.79e-19
C5072 P.n2827 VSUBS 5.79e-19
C5073 P.n2828 VSUBS 0.00232f
C5074 P.n2829 VSUBS 0.00232f
C5075 P.n2830 VSUBS 0.00123f
C5076 P.n2831 VSUBS 0.00119f
C5077 P.n2832 VSUBS 1.45e-19
C5078 P.n2833 VSUBS 1.81e-19
C5079 P.n2834 VSUBS 2.9e-19
C5080 P.n2835 VSUBS 7.24e-19
C5081 P.n2836 VSUBS 7.24e-19
C5082 P.n2837 VSUBS 3.26e-19
C5083 P.n2838 VSUBS 0.00749f
C5084 P.n2839 VSUBS 0.0012f
C5085 P.n2840 VSUBS 0.0239f
C5086 P.n2841 VSUBS 4.7e-19
C5087 P.n2842 VSUBS 0.00568f
C5088 P.n2843 VSUBS 0.00608f
C5089 P.n2844 VSUBS 0.00101f
C5090 P.n2845 VSUBS 0.00152f
C5091 P.n2846 VSUBS 0.00612f
C5092 P.n2847 VSUBS 0.00546f
C5093 P.n2848 VSUBS 0.018f
C5094 P.n2849 VSUBS 0.0183f
C5095 P.n2850 VSUBS 0.00101f
C5096 P.n2851 VSUBS 4.7e-19
C5097 P.n2852 VSUBS 0.00568f
C5098 P.n2853 VSUBS 0.00608f
C5099 P.n2854 VSUBS 0.00101f
C5100 P.n2855 VSUBS 0.00152f
C5101 P.n2856 VSUBS 0.0201f
C5102 P.n2857 VSUBS 1.53e-19
C5103 P.n2858 VSUBS 0.00123f
C5104 P.n2859 VSUBS 0.00123f
C5105 P.n2860 VSUBS 0.00304f
C5106 P.n2861 VSUBS 0.00366f
C5107 P.n2862 VSUBS 0.00123f
C5108 P.n2863 VSUBS 3.26e-19
C5109 P.n2864 VSUBS 0.00101f
C5110 P.n2865 VSUBS 9.05e-19
C5111 P.n2866 VSUBS 0.0159f
C5112 P.n2867 VSUBS 0.00101f
C5113 P.n2868 VSUBS 3.62e-19
C5114 P.n2869 VSUBS 3.26e-19
C5115 P.n2870 VSUBS 8.68e-19
C5116 P.n2871 VSUBS 9.05e-19
C5117 P.n2872 VSUBS 3.26e-19
C5118 P.n2873 VSUBS 3.26e-19
C5119 P.n2874 VSUBS 8.69e-19
C5120 P.n2875 VSUBS 8.69e-19
C5121 P.n2876 VSUBS 4.7e-19
C5122 P.n2877 VSUBS 0.00326f
C5123 P.n2878 VSUBS 0.00366f
C5124 P.n2879 VSUBS 0.00101f
C5125 P.n2880 VSUBS 5.07e-19
C5126 P.n2881 VSUBS 9.41e-19
C5127 P.n2882 VSUBS 0.00101f
C5128 P.n2883 VSUBS 4.7e-19
C5129 P.n2884 VSUBS 3.26e-19
C5130 P.n2885 VSUBS 2.9e-19
C5131 P.n2886 VSUBS 8.69e-19
C5132 P.n2887 VSUBS 9.41e-19
C5133 P.n2888 VSUBS 3.62e-19
C5134 P.n2889 VSUBS 2.9e-19
C5135 P.n2890 VSUBS 2.9e-19
C5136 P.n2891 VSUBS 7.24e-19
C5137 P.n2892 VSUBS 7.24e-19
C5138 P.n2893 VSUBS 0.00279f
C5139 P.n2894 VSUBS 0.00279f
C5140 P.n2895 VSUBS 3.26e-19
C5141 P.n2896 VSUBS 3.26e-19
C5142 P.n2897 VSUBS 2.9e-19
C5143 P.n2898 VSUBS 8.69e-19
C5144 P.n2899 VSUBS 0.0149f
C5145 P.n2900 VSUBS 8.69e-19
C5146 P.n2901 VSUBS 8.69e-19
C5147 P.n2902 VSUBS 2.9e-19
C5148 P.n2903 VSUBS 3.26e-19
C5149 P.n2904 VSUBS 2.17e-19
C5150 P.n2905 VSUBS 1.45e-19
C5151 P.n2906 VSUBS 8.68e-19
C5152 P.n2907 VSUBS 9.05e-19
C5153 P.n2908 VSUBS 3.26e-19
C5154 P.n2909 VSUBS 3.26e-19
C5155 P.n2910 VSUBS 8.69e-19
C5156 P.n2911 VSUBS 4.82e-19
C5157 P.n2912 VSUBS 2.55e-19
C5158 P.n2913 VSUBS 1.69e-19
C5159 P.n2914 VSUBS 0.0146f
C5160 P.n2915 VSUBS 5.79e-19
C5161 P.n2916 VSUBS 5.79e-19
C5162 P.n2917 VSUBS 0.00113f
C5163 P.n2918 VSUBS 7.62e-19
C5164 P.n2919 VSUBS 5.67e-19
C5165 P.n2920 VSUBS 5.79e-19
C5166 P.n2921 VSUBS 5.79e-19
C5167 P.n2922 VSUBS 9.41e-19
C5168 P.n2923 VSUBS 8.69e-19
C5169 P.n2924 VSUBS 3.96e-19
C5170 P.n2925 VSUBS 0.0593f
C5171 P.n2926 VSUBS 0.00109f
C5172 P.n2927 VSUBS 0.00109f
C5173 P.n2928 VSUBS 0.00191f
C5174 P.n2929 VSUBS 0.00287f
C5175 P.n2930 VSUBS 0.00444f
C5176 P.n2931 VSUBS 0.00567f
C5177 P.n2932 VSUBS 0.00287f
C5178 P.n2933 VSUBS 6.83e-19
C5179 P.n2934 VSUBS 0.00137f
C5180 P.n2935 VSUBS 0.00219f
C5181 P.n2936 VSUBS 0.00109f
C5182 P.n2937 VSUBS 5.47e-19
C5183 P.n2938 VSUBS 5.47e-19
C5184 P.n2939 VSUBS 0.0119f
C5185 P.n2940 VSUBS 0.00128f
C5186 P.n2941 VSUBS 7.6e-19
C5187 P.n2942 VSUBS 5.79e-19
C5188 P.n2943 VSUBS 5.79e-19
C5189 P.n2944 VSUBS 8.69e-19
C5190 P.n2945 VSUBS 9.41e-19
C5191 P.n2946 VSUBS 5.79e-19
C5192 P.n2947 VSUBS 5.79e-19
C5193 P.n2948 VSUBS 0.00192f
C5194 P.n2949 VSUBS 0.00203f
C5195 P.n2950 VSUBS 0.00123f
C5196 P.n2951 VSUBS 0.00123f
C5197 P.n2952 VSUBS 2.89e-19
C5198 P.n2953 VSUBS 1.09e-19
C5199 P.n2954 VSUBS 2.53e-19
C5200 P.n2955 VSUBS 6.51e-19
C5201 P.n2956 VSUBS 7.24e-19
C5202 P.n2957 VSUBS 5.07e-19
C5203 P.n2958 VSUBS 3.26e-19
C5204 P.n2959 VSUBS 2.17e-19
C5205 P.n2960 VSUBS 2.17e-19
C5206 P.n2961 VSUBS 1.45e-19
C5207 P.n2962 VSUBS 0.0121f
C5208 P.n2963 VSUBS 5.79e-19
C5209 P.n2964 VSUBS 7.6e-19
C5210 P.n2965 VSUBS 0.00119f
C5211 P.n2966 VSUBS 0.00123f
C5212 P.n2967 VSUBS 7.96e-19
C5213 P.n2968 VSUBS 5.79e-19
C5214 P.n2969 VSUBS 5.79e-19
C5215 P.n2970 VSUBS 0.00232f
C5216 P.n2971 VSUBS 0.00232f
C5217 P.n2972 VSUBS 0.00123f
C5218 P.n2973 VSUBS 0.00119f
C5219 P.n2974 VSUBS 1.45e-19
C5220 P.n2975 VSUBS 1.81e-19
C5221 P.n2976 VSUBS 2.9e-19
C5222 P.n2977 VSUBS 7.24e-19
C5223 P.n2978 VSUBS 7.24e-19
C5224 P.n2979 VSUBS 3.26e-19
C5225 P.n2980 VSUBS 0.0134f
C5226 P.n2981 VSUBS 0.0012f
C5227 P.n2982 VSUBS 0.0225f
C5228 P.n2983 VSUBS 4.7e-19
C5229 P.n2984 VSUBS 0.00568f
C5230 P.n2985 VSUBS 0.00608f
C5231 P.n2986 VSUBS 0.00101f
C5232 P.n2987 VSUBS 0.00152f
C5233 P.n2988 VSUBS 0.00612f
C5234 P.n2989 VSUBS 0.00546f
C5235 P.n2990 VSUBS 0.0158f
C5236 P.n2991 VSUBS 0.0161f
C5237 P.n2992 VSUBS 0.00101f
C5238 P.n2993 VSUBS 4.7e-19
C5239 P.n2994 VSUBS 0.00568f
C5240 P.n2995 VSUBS 0.00608f
C5241 P.n2996 VSUBS 0.00101f
C5242 P.n2997 VSUBS 0.00152f
C5243 P.n2998 VSUBS 0.026f
C5244 P.n2999 VSUBS 2.18e-19
C5245 P.n3000 VSUBS 0.00123f
C5246 P.n3001 VSUBS 0.00123f
C5247 P.n3002 VSUBS 0.00304f
C5248 P.n3003 VSUBS 0.00366f
C5249 P.n3004 VSUBS 0.00123f
C5250 P.n3005 VSUBS 3.26e-19
C5251 P.n3006 VSUBS 0.00101f
C5252 P.n3007 VSUBS 9.05e-19
C5253 P.n3008 VSUBS 0.0136f
C5254 P.n3009 VSUBS 0.00101f
C5255 P.n3010 VSUBS 3.62e-19
C5256 P.n3011 VSUBS 3.26e-19
C5257 P.n3012 VSUBS 8.68e-19
C5258 P.n3013 VSUBS 9.05e-19
C5259 P.n3014 VSUBS 3.26e-19
C5260 P.n3015 VSUBS 3.26e-19
C5261 P.n3016 VSUBS 8.69e-19
C5262 P.n3017 VSUBS 8.69e-19
C5263 P.n3018 VSUBS 4.7e-19
C5264 P.n3019 VSUBS 0.00326f
C5265 P.n3020 VSUBS 0.00366f
C5266 P.n3021 VSUBS 0.00101f
C5267 P.n3022 VSUBS 5.07e-19
C5268 P.n3023 VSUBS 9.41e-19
C5269 P.n3024 VSUBS 0.00101f
C5270 P.n3025 VSUBS 4.7e-19
C5271 P.n3026 VSUBS 3.26e-19
C5272 P.n3027 VSUBS 2.9e-19
C5273 P.n3028 VSUBS 8.69e-19
C5274 P.n3029 VSUBS 9.41e-19
C5275 P.n3030 VSUBS 3.62e-19
C5276 P.n3031 VSUBS 2.9e-19
C5277 P.n3032 VSUBS 2.9e-19
C5278 P.n3033 VSUBS 7.24e-19
C5279 P.n3034 VSUBS 7.24e-19
C5280 P.n3035 VSUBS 0.00279f
C5281 P.n3036 VSUBS 0.00279f
C5282 P.n3037 VSUBS 3.26e-19
C5283 P.n3038 VSUBS 3.26e-19
C5284 P.n3039 VSUBS 2.9e-19
C5285 P.n3040 VSUBS 8.69e-19
C5286 P.n3041 VSUBS 0.0126f
C5287 P.n3042 VSUBS 8.69e-19
C5288 P.n3043 VSUBS 8.69e-19
C5289 P.n3044 VSUBS 2.9e-19
C5290 P.n3045 VSUBS 3.26e-19
C5291 P.n3046 VSUBS 2.17e-19
C5292 P.n3047 VSUBS 1.45e-19
C5293 P.n3048 VSUBS 8.68e-19
C5294 P.n3049 VSUBS 9.05e-19
C5295 P.n3050 VSUBS 3.26e-19
C5296 P.n3051 VSUBS 3.26e-19
C5297 P.n3052 VSUBS 8.69e-19
C5298 P.n3053 VSUBS 0.0122f
C5299 P.n3054 VSUBS 8.69e-19
C5300 P.n3055 VSUBS 8.69e-19
C5301 P.n3056 VSUBS 2.9e-19
C5302 P.n3057 VSUBS 3.26e-19
C5303 P.n3058 VSUBS 3.26e-19
C5304 P.n3059 VSUBS 1.81e-19
C5305 P.n3060 VSUBS 1.09e-19
C5306 P.n3061 VSUBS 8.69e-19
C5307 P.n3062 VSUBS 8.69e-19
C5308 P.n3063 VSUBS 1.45e-19
C5309 P.n3064 VSUBS 1.45e-19
C5310 P.n3065 VSUBS 3.26e-19
C5311 P.n3066 VSUBS 3.26e-19
C5312 P.n3067 VSUBS 2.53e-19
C5313 P.n3068 VSUBS 7.96e-19
C5314 P.n3069 VSUBS 7.6e-19
C5315 P.n3070 VSUBS 2.53e-19
C5316 P.n3071 VSUBS 2.53e-19
C5317 P.n3072 VSUBS 2.17e-19
C5318 P.n3073 VSUBS 3.26e-19
C5319 P.n3074 VSUBS 0.0025f
C5320 P.n3075 VSUBS 0.00239f
C5321 P.n3076 VSUBS 7.24e-19
C5322 P.n3077 VSUBS 7.24e-19
C5323 P.n3078 VSUBS 2.9e-19
C5324 P.n3079 VSUBS 2.9e-19
C5325 P.n3080 VSUBS 5.07e-19
C5326 P.n3081 VSUBS 4.34e-19
C5327 P.n3082 VSUBS 7.24e-19
C5328 P.n3083 VSUBS 7.24e-19
C5329 P.n3084 VSUBS 0.00137f
C5330 P.n3085 VSUBS 0.00137f
C5331 P.n3086 VSUBS 0.00109f
C5332 P.n3087 VSUBS 0.0015f
C5333 P.n3088 VSUBS 0.00191f
C5334 P.n3089 VSUBS 0.0056f
C5335 P.n3090 VSUBS 0.00485f
C5336 P.n3091 VSUBS 8.88e-19
C5337 P.n3092 VSUBS 0.00191f
C5338 P.n3093 VSUBS 0.00198f
C5339 P.n3094 VSUBS 4.78e-19
C5340 P.n3095 VSUBS 6.15e-19
C5341 P.n3096 VSUBS 6.15e-19
C5342 P.n3097 VSUBS 2.73e-19
C5343 P.n3098 VSUBS 2.73e-19
C5344 P.n3099 VSUBS 0.00164f
C5345 P.n3100 VSUBS 0.00164f
C5346 P.n3101 VSUBS 4.78e-19
C5347 P.n3102 VSUBS 9.57e-19
C5348 P.n3103 VSUBS 8.88e-19
C5349 P.n3104 VSUBS 0.00191f
C5350 P.n3105 VSUBS 0.0054f
C5351 P.t51 VSUBS 2.64f
C5352 P.t30 VSUBS 2.64f
C5353 P.t73 VSUBS 2.64f
C5354 P.t122 VSUBS 2.64f
C5355 P.t114 VSUBS 2.64f
C5356 P.t3 VSUBS 2.64f
C5357 P.t50 VSUBS 2.64f
C5358 P.t84 VSUBS 2.64f
C5359 P.t4 VSUBS 2.64f
C5360 P.t126 VSUBS 2.64f
C5361 P.t20 VSUBS 2.64f
C5362 P.t74 VSUBS 2.78f
C5363 P.n3106 VSUBS 4.87f
C5364 P.n3107 VSUBS 2.51f
C5365 P.n3108 VSUBS 2.51f
C5366 P.n3109 VSUBS 2.51f
C5367 P.n3110 VSUBS 2.51f
C5368 P.n3111 VSUBS 2.51f
C5369 P.n3112 VSUBS 2.51f
C5370 P.n3113 VSUBS 2.51f
C5371 P.n3114 VSUBS 2.51f
C5372 P.n3115 VSUBS 2.51f
C5373 P.n3116 VSUBS 2.22f
C5374 P.n3117 VSUBS 0.405f
C5375 P.n3118 VSUBS 0.00191f
C5376 P.n3119 VSUBS 8.88e-19
C5377 P.n3120 VSUBS 9.57e-19
C5378 P.n3121 VSUBS 4.78e-19
C5379 P.n3122 VSUBS 0.00164f
C5380 P.n3123 VSUBS 0.00164f
C5381 P.n3124 VSUBS 2.73e-19
C5382 P.n3125 VSUBS 2.73e-19
C5383 P.n3126 VSUBS 6.15e-19
C5384 P.n3127 VSUBS 6.15e-19
C5385 P.n3128 VSUBS 4.78e-19
C5386 P.n3129 VSUBS 0.00198f
C5387 P.n3130 VSUBS 0.00191f
C5388 P.n3131 VSUBS 8.88e-19
C5389 P.n3132 VSUBS 0.00485f
C5390 P.n3133 VSUBS 0.0056f
C5391 P.n3134 VSUBS 0.00191f
C5392 P.n3135 VSUBS 0.0015f
C5393 P.n3136 VSUBS 0.00109f
C5394 P.n3137 VSUBS 0.00137f
C5395 P.n3138 VSUBS 0.0123f
C5396 P.n3139 VSUBS 5.79e-19
C5397 P.n3140 VSUBS 5.79e-19
C5398 P.n3141 VSUBS 9.41e-19
C5399 P.n3142 VSUBS 7.6e-19
C5400 P.n3143 VSUBS 5.79e-19
C5401 P.n3144 VSUBS 5.79e-19
C5402 P.n3145 VSUBS 8.69e-19
C5403 P.n3146 VSUBS 9.41e-19
C5404 P.n3147 VSUBS 5.79e-19
C5405 P.n3148 VSUBS 5.79e-19
C5406 P.n3149 VSUBS 0.00192f
C5407 P.n3150 VSUBS 0.00203f
C5408 P.n3151 VSUBS 0.00123f
C5409 P.n3152 VSUBS 0.00123f
C5410 P.n3153 VSUBS 2.89e-19
C5411 P.n3154 VSUBS 1.09e-19
C5412 P.n3155 VSUBS 2.53e-19
C5413 P.n3156 VSUBS 6.51e-19
C5414 P.n3157 VSUBS 7.24e-19
C5415 P.n3158 VSUBS 5.07e-19
C5416 P.n3159 VSUBS 3.26e-19
C5417 P.n3160 VSUBS 2.17e-19
C5418 P.n3161 VSUBS 2.17e-19
C5419 P.n3162 VSUBS 1.45e-19
C5420 P.n3163 VSUBS 0.0126f
C5421 P.n3164 VSUBS 5.79e-19
C5422 P.n3165 VSUBS 5.79e-19
C5423 P.n3166 VSUBS 7.6e-19
C5424 P.n3167 VSUBS 0.00119f
C5425 P.n3168 VSUBS 0.00123f
C5426 P.n3169 VSUBS 7.96e-19
C5427 P.n3170 VSUBS 5.79e-19
C5428 P.n3171 VSUBS 5.79e-19
C5429 P.n3172 VSUBS 0.00232f
C5430 P.n3173 VSUBS 0.00232f
C5431 P.n3174 VSUBS 0.00123f
C5432 P.n3175 VSUBS 0.00119f
C5433 P.n3176 VSUBS 1.45e-19
C5434 P.n3177 VSUBS 1.81e-19
C5435 P.n3178 VSUBS 2.9e-19
C5436 P.n3179 VSUBS 7.24e-19
C5437 P.n3180 VSUBS 7.24e-19
C5438 P.n3181 VSUBS 3.26e-19
C5439 P.n3182 VSUBS 0.0134f
C5440 P.n3183 VSUBS 0.00119f
C5441 P.n3184 VSUBS 0.00119f
C5442 P.n3185 VSUBS 0.00123f
C5443 P.n3186 VSUBS 0.00123f
C5444 P.n3187 VSUBS 0.00304f
C5445 P.n3188 VSUBS 0.00366f
C5446 P.n3189 VSUBS 0.00123f
C5447 P.n3190 VSUBS 3.26e-19
C5448 P.n3191 VSUBS 0.00101f
C5449 P.n3192 VSUBS 9.05e-19
C5450 P.n3193 VSUBS 0.02f
C5451 P.n3194 VSUBS 3.62e-19
C5452 P.n3195 VSUBS 3.47e-19
C5453 P.n3196 VSUBS 8.68e-19
C5454 P.n3197 VSUBS 9.05e-19
C5455 P.n3198 VSUBS 3.26e-19
C5456 P.n3199 VSUBS 3.26e-19
C5457 P.n3200 VSUBS 8.69e-19
C5458 P.n3201 VSUBS 8.69e-19
C5459 P.n3202 VSUBS 4.7e-19
C5460 P.n3203 VSUBS 0.00326f
C5461 P.n3204 VSUBS 0.00366f
C5462 P.n3205 VSUBS 0.00101f
C5463 P.n3206 VSUBS 5.07e-19
C5464 P.n3207 VSUBS 9.41e-19
C5465 P.n3208 VSUBS 0.00101f
C5466 P.n3209 VSUBS 4.7e-19
C5467 P.n3210 VSUBS 3.26e-19
C5468 P.n3211 VSUBS 2.9e-19
C5469 P.n3212 VSUBS 8.69e-19
C5470 P.n3213 VSUBS 9.41e-19
C5471 P.n3214 VSUBS 3.62e-19
C5472 P.n3215 VSUBS 2.9e-19
C5473 P.n3216 VSUBS 2.9e-19
C5474 P.n3217 VSUBS 7.24e-19
C5475 P.n3218 VSUBS 7.24e-19
C5476 P.n3219 VSUBS 0.00279f
C5477 P.n3220 VSUBS 0.00279f
C5478 P.n3221 VSUBS 3.26e-19
C5479 P.n3222 VSUBS 3.26e-19
C5480 P.n3223 VSUBS 2.9e-19
C5481 P.n3224 VSUBS 8.69e-19
C5482 P.n3225 VSUBS 0.0189f
C5483 P.n3226 VSUBS 8.69e-19
C5484 P.n3227 VSUBS 2.9e-19
C5485 P.n3228 VSUBS 3.26e-19
C5486 P.n3229 VSUBS 2.17e-19
C5487 P.n3230 VSUBS 1.45e-19
C5488 P.n3231 VSUBS 8.68e-19
C5489 P.n3232 VSUBS 9.05e-19
C5490 P.n3233 VSUBS 3.26e-19
C5491 P.n3234 VSUBS 3.26e-19
C5492 P.n3235 VSUBS 8.69e-19
C5493 P.n3236 VSUBS 0.0186f
C5494 P.n3237 VSUBS 8.69e-19
C5495 P.n3238 VSUBS 2.9e-19
C5496 P.n3239 VSUBS 3.26e-19
C5497 P.n3240 VSUBS 3.26e-19
C5498 P.n3241 VSUBS 1.81e-19
C5499 P.n3242 VSUBS 1.09e-19
C5500 P.n3243 VSUBS 8.69e-19
C5501 P.n3244 VSUBS 8.69e-19
C5502 P.n3245 VSUBS 1.45e-19
C5503 P.n3246 VSUBS 1.45e-19
C5504 P.n3247 VSUBS 3.26e-19
C5505 P.n3248 VSUBS 3.26e-19
C5506 P.n3249 VSUBS 2.53e-19
C5507 P.n3250 VSUBS 7.96e-19
C5508 P.n3251 VSUBS 7.6e-19
C5509 P.n3252 VSUBS 2.53e-19
C5510 P.n3253 VSUBS 2.53e-19
C5511 P.n3254 VSUBS 2.17e-19
C5512 P.n3255 VSUBS 3.26e-19
C5513 P.n3256 VSUBS 0.0025f
C5514 P.n3257 VSUBS 0.00239f
C5515 P.n3258 VSUBS 7.24e-19
C5516 P.n3259 VSUBS 7.24e-19
C5517 P.n3260 VSUBS 2.9e-19
C5518 P.n3261 VSUBS 2.9e-19
C5519 P.n3262 VSUBS 5.07e-19
C5520 P.n3263 VSUBS 4.34e-19
C5521 P.n3264 VSUBS 7.24e-19
C5522 P.n3265 VSUBS 7.24e-19
C5523 P.n3266 VSUBS 0.00137f
C5524 P.n3267 VSUBS 5.47e-19
C5525 P.n3268 VSUBS 5.47e-19
C5526 P.n3269 VSUBS 0.00109f
C5527 P.n3270 VSUBS 0.00219f
C5528 P.n3271 VSUBS 0.00137f
C5529 P.n3272 VSUBS 6.83e-19
C5530 P.n3273 VSUBS 0.00287f
C5531 P.n3274 VSUBS 0.00567f
C5532 P.n3275 VSUBS 0.00444f
C5533 P.n3276 VSUBS 0.00287f
C5534 P.n3277 VSUBS 0.00191f
C5535 P.n3278 VSUBS 0.00109f
C5536 P.n3279 VSUBS 0.00109f
C5537 P.n3280 VSUBS 0.00191f
C5538 P.n3281 VSUBS 0.00287f
C5539 P.n3282 VSUBS 0.0199f
C5540 P.n3283 VSUBS 0.326f
C5541 P.n3284 VSUBS 0.305f
C5542 P.n3285 VSUBS 0.00137f
C5543 P.n3286 VSUBS 0.00164f
C5544 P.n3287 VSUBS 5.79e-19
C5545 P.n3288 VSUBS 5.79e-19
C5546 P.n3289 VSUBS 9.41e-19
C5547 P.n3290 VSUBS 8.69e-19
C5548 P.n3291 VSUBS 3.96e-19
C5549 P.n3292 VSUBS 0.00246f
C5550 P.n3293 VSUBS 0.00137f
C5551 P.n3294 VSUBS 0.00157f
C5552 P.n3295 VSUBS 0.00239f
C5553 P.n3296 VSUBS 0.00137f
C5554 P.n3297 VSUBS 0.00636f
C5555 P.n3298 VSUBS 0.00806f
C5556 P.n3299 VSUBS 0.00273f
C5557 P.n3300 VSUBS 0.00575f
C5558 P.n3301 VSUBS 5.79e-19
C5559 P.n3302 VSUBS 0.00113f
C5560 P.n3303 VSUBS 7.62e-19
C5561 P.n3304 VSUBS 5.67e-19
C5562 P.n3305 VSUBS 0.00116f
C5563 P.n3306 VSUBS 0.00198f
C5564 P.n3307 VSUBS 0.00226f
C5565 P.n3308 VSUBS 0.00116f
C5566 P.n3309 VSUBS 0.00198f
C5567 P.n3310 VSUBS 0.00267f
C5568 P.n3311 VSUBS 0.0106f
C5569 P.n3312 VSUBS 0.0122f
C5570 P.n3313 VSUBS 0.0025f
C5571 P.n3314 VSUBS 3.26e-19
C5572 P.n3315 VSUBS 2.17e-19
C5573 P.n3316 VSUBS 2.53e-19
C5574 P.n3317 VSUBS 2.53e-19
C5575 P.n3318 VSUBS 7.6e-19
C5576 P.n3319 VSUBS 9.39e-19
C5577 P.n3320 VSUBS 1.1e-19
C5578 P.n3321 VSUBS 0.0149f
C5579 P.n3322 VSUBS 5.79e-19
C5580 P.n3323 VSUBS 5.79e-19
C5581 P.n3324 VSUBS 7.6e-19
C5582 P.n3325 VSUBS 0.00119f
C5583 P.n3326 VSUBS 0.00123f
C5584 P.n3327 VSUBS 7.96e-19
C5585 P.n3328 VSUBS 5.79e-19
C5586 P.n3329 VSUBS 5.79e-19
C5587 P.n3330 VSUBS 0.00232f
C5588 P.n3331 VSUBS 0.00232f
C5589 P.n3332 VSUBS 0.00123f
C5590 P.n3333 VSUBS 0.00119f
C5591 P.n3334 VSUBS 1.45e-19
C5592 P.n3335 VSUBS 1.81e-19
C5593 P.n3336 VSUBS 2.9e-19
C5594 P.n3337 VSUBS 7.24e-19
C5595 P.n3338 VSUBS 7.24e-19
C5596 P.n3339 VSUBS 3.26e-19
C5597 P.n3340 VSUBS 0.0156f
C5598 P.n3341 VSUBS 0.00119f
C5599 P.n3342 VSUBS 0.00119f
C5600 P.n3343 VSUBS 0.00123f
C5601 P.n3344 VSUBS 0.00123f
C5602 P.n3345 VSUBS 0.00304f
C5603 P.n3346 VSUBS 0.00366f
C5604 P.n3347 VSUBS 0.00123f
C5605 P.n3348 VSUBS 3.26e-19
C5606 P.n3349 VSUBS 0.00101f
C5607 P.n3350 VSUBS 9.05e-19
C5608 P.n3351 VSUBS 0.0215f
C5609 P.n3352 VSUBS 3.62e-19
C5610 P.n3353 VSUBS 3.48e-19
C5611 P.n3354 VSUBS 8.68e-19
C5612 P.n3355 VSUBS 9.05e-19
C5613 P.n3356 VSUBS 3.26e-19
C5614 P.n3357 VSUBS 3.26e-19
C5615 P.n3358 VSUBS 8.69e-19
C5616 P.n3359 VSUBS 8.69e-19
C5617 P.n3360 VSUBS 4.7e-19
C5618 P.n3361 VSUBS 0.00326f
C5619 P.n3362 VSUBS 0.00366f
C5620 P.n3363 VSUBS 0.00101f
C5621 P.n3364 VSUBS 5.07e-19
C5622 P.n3365 VSUBS 9.41e-19
C5623 P.n3366 VSUBS 0.00101f
C5624 P.n3367 VSUBS 4.7e-19
C5625 P.n3368 VSUBS 3.26e-19
C5626 P.n3369 VSUBS 2.9e-19
C5627 P.n3370 VSUBS 8.69e-19
C5628 P.n3371 VSUBS 9.41e-19
C5629 P.n3372 VSUBS 3.62e-19
C5630 P.n3373 VSUBS 2.9e-19
C5631 P.n3374 VSUBS 2.9e-19
C5632 P.n3375 VSUBS 7.24e-19
C5633 P.n3376 VSUBS 7.24e-19
C5634 P.n3377 VSUBS 0.00279f
C5635 P.n3378 VSUBS 0.00279f
C5636 P.n3379 VSUBS 3.26e-19
C5637 P.n3380 VSUBS 3.26e-19
C5638 P.n3381 VSUBS 2.9e-19
C5639 P.n3382 VSUBS 8.69e-19
C5640 P.n3383 VSUBS 0.0203f
C5641 P.n3384 VSUBS 8.69e-19
C5642 P.n3385 VSUBS 2.9e-19
C5643 P.n3386 VSUBS 3.26e-19
C5644 P.n3387 VSUBS 2.17e-19
C5645 P.n3388 VSUBS 1.45e-19
C5646 P.n3389 VSUBS 8.68e-19
C5647 P.n3390 VSUBS 9.05e-19
C5648 P.n3391 VSUBS 3.26e-19
C5649 P.n3392 VSUBS 3.26e-19
C5650 P.n3393 VSUBS 8.69e-19
C5651 P.n3394 VSUBS 4.82e-19
C5652 P.n3395 VSUBS 2.55e-19
C5653 P.n3396 VSUBS 1.69e-19
C5654 P.n3397 VSUBS 0.0054f
C5655 P.n3399 VSUBS 0.01f
C5656 P.n3400 VSUBS 0.00957f
C5657 P.n3401 VSUBS 0.425f
C5658 P.n3402 VSUBS 7.52e-19
C5659 P.n3403 VSUBS 0.00267f
C5660 P.n3404 VSUBS 0.00273f
C5661 P.n3405 VSUBS 0.0145f
C5662 P.n3406 VSUBS 8.69e-19
C5663 P.n3407 VSUBS 8.69e-19
C5664 P.n3408 VSUBS 2.9e-19
C5665 P.n3409 VSUBS 3.26e-19
C5666 P.n3410 VSUBS 3.26e-19
C5667 P.n3411 VSUBS 1.81e-19
C5668 P.n3412 VSUBS 1.09e-19
C5669 P.n3413 VSUBS 3.42e-20
C5670 P.n3414 VSUBS 0.00107f
C5671 P.n3415 VSUBS 6.71e-19
C5672 P.n3416 VSUBS 0.00294f
C5673 P.n3418 VSUBS 0.432f
C5674 P.n3419 VSUBS 0.43f
C5675 P.n3420 VSUBS 0.00137f
C5676 P.n3421 VSUBS 0.00137f
C5677 P.n3422 VSUBS 0.00137f
C5678 P.n3423 VSUBS 0.00137f
C5679 P.n3424 VSUBS 0.00137f
C5680 P.n3425 VSUBS 0.00137f
C5681 P.n3426 VSUBS 0.0013f
C5682 P.n3427 VSUBS 2.73e-19
C5683 P.n3428 VSUBS 0.00109f
C5684 P.n3429 VSUBS 0.0013f
C5685 P.n3430 VSUBS 0.00137f
C5686 P.n3431 VSUBS 0.00137f
C5687 P.n3432 VSUBS 0.00499f
C5688 P.n3433 VSUBS 0.00608f
C5689 P.n3434 VSUBS 0.00198f
C5690 P.n3435 VSUBS 0.00137f
C5691 P.n3436 VSUBS 0.00116f
C5692 P.n3437 VSUBS 6.15e-19
C5693 P.n3438 VSUBS 9.57e-19
C5694 P.n3439 VSUBS 0.00116f
C5695 P.n3440 VSUBS 6.15e-19
C5696 P.n3441 VSUBS 8.88e-19
C5697 P.n3442 VSUBS 0.00116f
C5698 P.n3443 VSUBS 6.83e-19
C5699 P.n3444 VSUBS 8.88e-19
C5700 P.n3445 VSUBS 0.00116f
C5701 P.n3446 VSUBS 6.15e-19
C5702 P.n3447 VSUBS 0.0013f
C5703 P.n3448 VSUBS 0.00137f
C5704 P.n3449 VSUBS 0.00137f
C5705 P.n3450 VSUBS 0.00748f
C5706 P.n3451 VSUBS 0.00835f
C5707 P.n3452 VSUBS 0.00273f
C5708 P.n3453 VSUBS 0.00273f
C5709 P.n3454 VSUBS 0.00192f
C5710 P.n3455 VSUBS 0.00203f
C5711 P.n3456 VSUBS 0.00123f
C5712 P.n3457 VSUBS 0.00123f
C5713 P.n3458 VSUBS 2.89e-19
C5714 P.n3459 VSUBS 1.09e-19
C5715 P.n3460 VSUBS 6.63e-19
C5716 P.n3461 VSUBS 7.24e-19
C5717 P.n3462 VSUBS 6.51e-19
C5718 P.n3463 VSUBS 2.53e-19
C5719 P.n3465 VSUBS 0.00267f
C5720 P.n3466 VSUBS 0.00267f
C5721 P.n3467 VSUBS 0.0026f
C5722 P.n3468 VSUBS 0.407f
C5723 P.n3469 VSUBS 0.00615f
C5724 P.n3470 VSUBS 0.00273f
C5725 P.n3471 VSUBS 0.00157f
C5726 P.n3472 VSUBS 0.00137f
C5727 P.n3473 VSUBS 0.00137f
C5728 P.n3474 VSUBS 0.0013f
C5729 P.n3475 VSUBS 0.00137f
C5730 P.n3476 VSUBS 0.00137f
C5731 P.n3477 VSUBS 0.00137f
C5732 P.n3478 VSUBS 0.00157f
C5733 P.n3479 VSUBS 0.00267f
C5734 P.n3480 VSUBS 0.394f
C5735 P.n3481 VSUBS 0.394f
C5736 P.n3482 VSUBS 0.00137f
C5737 P.n3483 VSUBS 8.88e-19
C5738 P.n3484 VSUBS 0.00137f
C5739 P.n3485 VSUBS 0.00109f
C5740 P.n3486 VSUBS 6.15e-19
C5741 P.n3487 VSUBS 7.52e-19
C5742 P.n3488 VSUBS 7.52e-19
C5743 P.n3489 VSUBS 8.88e-19
C5744 P.n3490 VSUBS 0.0013f
C5745 P.n3491 VSUBS 0.00109f
C5746 P.n3492 VSUBS 6.83e-19
C5747 P.n3493 VSUBS 6.83e-19
C5748 P.n3494 VSUBS 6.83e-19
C5749 P.n3495 VSUBS 8.88e-19
C5750 P.n3496 VSUBS 0.00171f
C5751 P.n3497 VSUBS 0.00137f
C5752 P.n3498 VSUBS 0.00437f
C5753 P.n3499 VSUBS 0.00608f
C5754 P.n3500 VSUBS 0.00273f
C5755 P.n3501 VSUBS 0.00116f
C5756 P.n3502 VSUBS 0.00123f
C5757 P.n3503 VSUBS 0.00157f
C5758 P.n3504 VSUBS 0.00116f
C5759 P.n3505 VSUBS 6.83e-19
C5760 P.n3506 VSUBS 7.52e-19
C5761 P.n3507 VSUBS 0.0013f
C5762 P.n3508 VSUBS 0.0015f
C5763 P.n3509 VSUBS 0.00116f
C5764 P.n3510 VSUBS 0.00116f
C5765 P.n3511 VSUBS 0.0015f
C5766 P.n3512 VSUBS 0.00198f
C5767 P.n3513 VSUBS 0.00861f
C5768 P.n3514 VSUBS 0.00943f
C5769 P.n3515 VSUBS 0.00273f
C5770 P.n3516 VSUBS 0.00273f
C5771 P.n3517 VSUBS 6.63e-19
C5772 P.n3518 VSUBS 7.24e-19
C5773 P.n3519 VSUBS 6.51e-19
C5774 P.n3520 VSUBS 2.53e-19
C5775 P.n3521 VSUBS 0.00192f
C5776 P.n3522 VSUBS 0.00203f
C5777 P.n3523 VSUBS 0.00123f
C5778 P.n3524 VSUBS 0.00123f
C5779 P.n3525 VSUBS 2.89e-19
C5780 P.n3526 VSUBS 1.09e-19
C5781 P.n3528 VSUBS 0.00267f
C5782 P.n3529 VSUBS 0.00267f
C5783 P.n3530 VSUBS 0.00738f
C5784 P.n3531 VSUBS 0.00738f
C5785 P.n3532 VSUBS 0.00273f
C5786 P.n3533 VSUBS 9.57e-19
C5787 P.n3534 VSUBS 0.00198f
C5788 P.n3535 VSUBS 0.00198f
C5789 P.n3536 VSUBS 6.83e-19
C5790 P.n3537 VSUBS 7.52e-19
C5791 P.n3538 VSUBS 0.00198f
C5792 P.n3539 VSUBS 0.00198f
C5793 P.n3540 VSUBS 9.57e-19
C5794 P.n3541 VSUBS 0.00267f
C5795 P.n3542 VSUBS 0.00205f
C5796 P.n3543 VSUBS 0.828f
C5797 P.n3544 VSUBS 0.407f
C5798 P.n3545 VSUBS 0.00109f
C5799 P.n3546 VSUBS 6.15e-19
C5800 P.n3547 VSUBS 7.52e-19
C5801 P.n3548 VSUBS 7.52e-19
C5802 P.n3549 VSUBS 8.88e-19
C5803 P.n3550 VSUBS 0.00137f
C5804 P.n3551 VSUBS 0.00109f
C5805 P.n3552 VSUBS 6.15e-19
C5806 P.n3553 VSUBS 7.52e-19
C5807 P.n3554 VSUBS 7.52e-19
C5808 P.n3555 VSUBS 8.2e-19
C5809 P.n3556 VSUBS 0.0013f
C5810 P.n3557 VSUBS 0.00109f
C5811 P.n3558 VSUBS 6.15e-19
C5812 P.n3559 VSUBS 7.52e-19
C5813 P.n3560 VSUBS 7.52e-19
C5814 P.n3561 VSUBS 0.0056f
C5815 P.n3562 VSUBS 0.00608f
C5816 P.n3563 VSUBS 0.00198f
C5817 P.n3564 VSUBS 0.00198f
C5818 P.n3565 VSUBS 0.0105f
C5819 P.n3566 VSUBS 5.79e-19
C5820 P.n3567 VSUBS 0.00113f
C5821 P.n3568 VSUBS 5.79e-19
C5822 P.n3569 VSUBS 5.79e-19
C5823 P.n3570 VSUBS 9.41e-19
C5824 P.n3571 VSUBS 8.69e-19
C5825 P.n3572 VSUBS 3.96e-19
C5826 P.n3573 VSUBS 7.62e-19
C5827 P.n3574 VSUBS 5.67e-19
C5828 P.n3575 VSUBS 0.00116f
C5829 P.n3576 VSUBS 7.52e-19
C5830 P.n3577 VSUBS 7.52e-19
C5831 P.n3578 VSUBS 0.00123f
C5832 P.n3579 VSUBS 0.0015f
C5833 P.n3580 VSUBS 7.52e-19
C5834 P.n3581 VSUBS 4.78e-19
C5835 P.n3582 VSUBS 6.83e-19
C5836 P.n3583 VSUBS 7.52e-19
C5837 P.n3584 VSUBS 0.00123f
C5838 P.n3585 VSUBS 0.0015f
C5839 P.n3586 VSUBS 0.00116f
C5840 P.n3587 VSUBS 0.00116f
C5841 P.n3588 VSUBS 0.00943f
C5842 P.n3589 VSUBS 0.00943f
C5843 P.n3590 VSUBS 0.00273f
C5844 P.n3591 VSUBS 0.0109f
C5845 P.n3592 VSUBS 5.79e-19
C5846 P.n3593 VSUBS 7.6e-19
C5847 P.n3594 VSUBS 0.00119f
C5848 P.n3595 VSUBS 0.00123f
C5849 P.n3596 VSUBS 7.96e-19
C5850 P.n3597 VSUBS 5.79e-19
C5851 P.n3598 VSUBS 5.79e-19
C5852 P.n3599 VSUBS 0.00232f
C5853 P.n3600 VSUBS 0.00232f
C5854 P.n3601 VSUBS 0.00123f
C5855 P.n3602 VSUBS 0.00119f
C5856 P.n3603 VSUBS 1.45e-19
C5857 P.n3604 VSUBS 1.81e-19
C5858 P.n3605 VSUBS 2.9e-19
C5859 P.n3606 VSUBS 7.24e-19
C5860 P.n3607 VSUBS 7.24e-19
C5861 P.n3608 VSUBS 3.26e-19
C5862 P.n3609 VSUBS 0.0122f
C5863 P.n3610 VSUBS 0.0012f
C5864 P.n3611 VSUBS 0.0222f
C5865 P.n3612 VSUBS 4.7e-19
C5866 P.n3613 VSUBS 0.00568f
C5867 P.n3614 VSUBS 0.00608f
C5868 P.n3615 VSUBS 0.00101f
C5869 P.n3616 VSUBS 0.00152f
C5870 P.n3617 VSUBS 0.00612f
C5871 P.n3618 VSUBS 0.00546f
C5872 P.n3619 VSUBS 0.0165f
C5873 P.n3620 VSUBS 0.0168f
C5874 P.n3621 VSUBS 0.00101f
C5875 P.n3622 VSUBS 4.7e-19
C5876 P.n3623 VSUBS 0.00568f
C5877 P.n3624 VSUBS 0.00608f
C5878 P.n3625 VSUBS 0.00101f
C5879 P.n3626 VSUBS 0.00152f
C5880 P.n3627 VSUBS 0.0248f
C5881 P.n3628 VSUBS 2.04e-19
C5882 P.n3629 VSUBS 0.00123f
C5883 P.n3630 VSUBS 0.00123f
C5884 P.n3631 VSUBS 0.00304f
C5885 P.n3632 VSUBS 0.00366f
C5886 P.n3633 VSUBS 0.00123f
C5887 P.n3634 VSUBS 3.26e-19
C5888 P.n3635 VSUBS 0.00101f
C5889 P.n3636 VSUBS 9.05e-19
C5890 P.n3637 VSUBS 0.0144f
C5891 P.n3638 VSUBS 0.00101f
C5892 P.n3639 VSUBS 3.62e-19
C5893 P.n3640 VSUBS 3.26e-19
C5894 P.n3641 VSUBS 8.68e-19
C5895 P.n3642 VSUBS 9.05e-19
C5896 P.n3643 VSUBS 3.26e-19
C5897 P.n3644 VSUBS 3.26e-19
C5898 P.n3645 VSUBS 8.69e-19
C5899 P.n3646 VSUBS 8.69e-19
C5900 P.n3647 VSUBS 4.7e-19
C5901 P.n3648 VSUBS 0.00326f
C5902 P.n3649 VSUBS 0.00366f
C5903 P.n3650 VSUBS 0.00101f
C5904 P.n3651 VSUBS 5.07e-19
C5905 P.n3652 VSUBS 9.41e-19
C5906 P.n3653 VSUBS 0.00101f
C5907 P.n3654 VSUBS 4.7e-19
C5908 P.n3655 VSUBS 3.26e-19
C5909 P.n3656 VSUBS 2.9e-19
C5910 P.n3657 VSUBS 8.69e-19
C5911 P.n3658 VSUBS 9.41e-19
C5912 P.n3659 VSUBS 3.62e-19
C5913 P.n3660 VSUBS 2.9e-19
C5914 P.n3661 VSUBS 2.9e-19
C5915 P.n3662 VSUBS 7.24e-19
C5916 P.n3663 VSUBS 7.24e-19
C5917 P.n3664 VSUBS 0.00279f
C5918 P.n3665 VSUBS 0.00279f
C5919 P.n3666 VSUBS 3.26e-19
C5920 P.n3667 VSUBS 3.26e-19
C5921 P.n3668 VSUBS 2.9e-19
C5922 P.n3669 VSUBS 8.69e-19
C5923 P.n3670 VSUBS 0.0134f
C5924 P.n3671 VSUBS 8.69e-19
C5925 P.n3672 VSUBS 8.69e-19
C5926 P.n3673 VSUBS 2.9e-19
C5927 P.n3674 VSUBS 3.26e-19
C5928 P.n3675 VSUBS 2.17e-19
C5929 P.n3676 VSUBS 1.45e-19
C5930 P.n3677 VSUBS 8.68e-19
C5931 P.n3678 VSUBS 9.05e-19
C5932 P.n3679 VSUBS 3.26e-19
C5933 P.n3680 VSUBS 3.26e-19
C5934 P.n3681 VSUBS 8.69e-19
C5935 P.n3682 VSUBS 0.0025f
C5936 P.n3683 VSUBS 3.26e-19
C5937 P.n3684 VSUBS 2.17e-19
C5938 P.n3685 VSUBS 2.53e-19
C5939 P.n3686 VSUBS 2.53e-19
C5940 P.n3687 VSUBS 7.6e-19
C5941 P.n3688 VSUBS 9.39e-19
C5942 P.n3689 VSUBS 1.1e-19
C5943 P.n3690 VSUBS 4.82e-19
C5944 P.n3691 VSUBS 2.55e-19
C5945 P.n3692 VSUBS 1.69e-19
C5946 P.n3693 VSUBS 0.00273f
C5947 P.n3694 VSUBS 0.00267f
C5948 P.n3695 VSUBS 0.00267f
C5949 P.n3696 VSUBS 0.00738f
C5950 P.n3697 VSUBS 0.00738f
C5951 P.n3698 VSUBS 0.00273f
C5952 P.n3699 VSUBS 0.00219f
C5953 P.n3700 VSUBS 7.52e-19
C5954 P.n3701 VSUBS 7.52e-19
C5955 P.n3702 VSUBS 0.00191f
C5956 P.n3703 VSUBS 0.00198f
C5957 P.n3704 VSUBS 7.52e-19
C5958 P.n3705 VSUBS 7.52e-19
C5959 P.n3706 VSUBS 0.00219f
C5960 P.n3707 VSUBS 0.425f
C5961 P.n3708 VSUBS 0.183f
.ends

