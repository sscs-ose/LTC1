magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2530 -2410 2530 2410
<< nwell >>
rect -530 -410 530 410
<< pmos >>
rect -356 -280 -256 280
rect -152 -280 -52 280
rect 52 -280 152 280
rect 256 -280 356 280
<< pdiff >>
rect -444 258 -356 280
rect -444 -258 -431 258
rect -385 -258 -356 258
rect -444 -280 -356 -258
rect -256 258 -152 280
rect -256 -258 -227 258
rect -181 -258 -152 258
rect -256 -280 -152 -258
rect -52 258 52 280
rect -52 -258 -23 258
rect 23 -258 52 258
rect -52 -280 52 -258
rect 152 258 256 280
rect 152 -258 181 258
rect 227 -258 256 258
rect 152 -280 256 -258
rect 356 258 444 280
rect 356 -258 385 258
rect 431 -258 444 258
rect 356 -280 444 -258
<< pdiffc >>
rect -431 -258 -385 258
rect -227 -258 -181 258
rect -23 -258 23 258
rect 181 -258 227 258
rect 385 -258 431 258
<< polysilicon >>
rect -356 280 -256 324
rect -152 280 -52 324
rect 52 280 152 324
rect 256 280 356 324
rect -356 -324 -256 -280
rect -152 -324 -52 -280
rect 52 -324 152 -280
rect 256 -324 356 -280
<< metal1 >>
rect -431 258 -385 278
rect -431 -278 -385 -258
rect -227 258 -181 278
rect -227 -278 -181 -258
rect -23 258 23 278
rect -23 -278 23 -258
rect 181 258 227 278
rect 181 -278 227 -258
rect 385 258 431 278
rect 385 -278 431 -258
<< end >>
