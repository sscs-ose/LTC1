magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2208 -2120 2348 3320
<< nwell >>
rect -208 -120 348 1320
<< mvpmos >>
rect 0 0 140 1200
<< mvpdiff >>
rect -88 1167 0 1200
rect -88 651 -75 1167
rect -29 651 0 1167
rect -88 574 0 651
rect -88 528 -75 574
rect -29 528 0 574
rect -88 471 0 528
rect -88 425 -75 471
rect -29 425 0 471
rect -88 368 0 425
rect -88 322 -75 368
rect -29 322 0 368
rect -88 265 0 322
rect -88 219 -75 265
rect -29 219 0 265
rect -88 162 0 219
rect -88 116 -75 162
rect -29 116 0 162
rect -88 59 0 116
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 1167 228 1200
rect 140 651 169 1167
rect 215 651 228 1167
rect 140 574 228 651
rect 140 528 169 574
rect 215 528 228 574
rect 140 471 228 528
rect 140 425 169 471
rect 215 425 228 471
rect 140 368 228 425
rect 140 322 169 368
rect 215 322 228 368
rect 140 265 228 322
rect 140 219 169 265
rect 215 219 228 265
rect 140 162 228 219
rect 140 116 169 162
rect 215 116 228 162
rect 140 59 228 116
rect 140 13 169 59
rect 215 13 228 59
rect 140 0 228 13
<< mvpdiffc >>
rect -75 651 -29 1167
rect -75 528 -29 574
rect -75 425 -29 471
rect -75 322 -29 368
rect -75 219 -29 265
rect -75 116 -29 162
rect -75 13 -29 59
rect 169 651 215 1167
rect 169 528 215 574
rect 169 425 215 471
rect 169 322 215 368
rect 169 219 215 265
rect 169 116 215 162
rect 169 13 215 59
<< polysilicon >>
rect 0 1200 140 1244
rect 0 -44 140 0
<< metal1 >>
rect -75 1167 -29 1200
rect -75 574 -29 651
rect -75 471 -29 528
rect -75 368 -29 425
rect -75 265 -29 322
rect -75 162 -29 219
rect -75 59 -29 116
rect -75 0 -29 13
rect 169 1167 215 1200
rect 169 574 215 651
rect 169 471 215 528
rect 169 368 215 425
rect 169 265 215 322
rect 169 162 215 219
rect 169 59 215 116
rect 169 0 215 13
<< labels >>
rlabel metal1 192 600 192 600 4 D
rlabel metal1 -52 600 -52 600 4 S
<< end >>
