magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1112 -1763 1112 1763
<< metal1 >>
rect -112 757 112 763
rect -112 731 -106 757
rect -80 731 -44 757
rect -18 731 18 757
rect 44 731 80 757
rect 106 731 112 757
rect -112 695 112 731
rect -112 669 -106 695
rect -80 669 -44 695
rect -18 669 18 695
rect 44 669 80 695
rect 106 669 112 695
rect -112 633 112 669
rect -112 607 -106 633
rect -80 607 -44 633
rect -18 607 18 633
rect 44 607 80 633
rect 106 607 112 633
rect -112 571 112 607
rect -112 545 -106 571
rect -80 545 -44 571
rect -18 545 18 571
rect 44 545 80 571
rect 106 545 112 571
rect -112 509 112 545
rect -112 483 -106 509
rect -80 483 -44 509
rect -18 483 18 509
rect 44 483 80 509
rect 106 483 112 509
rect -112 447 112 483
rect -112 421 -106 447
rect -80 421 -44 447
rect -18 421 18 447
rect 44 421 80 447
rect 106 421 112 447
rect -112 385 112 421
rect -112 359 -106 385
rect -80 359 -44 385
rect -18 359 18 385
rect 44 359 80 385
rect 106 359 112 385
rect -112 323 112 359
rect -112 297 -106 323
rect -80 297 -44 323
rect -18 297 18 323
rect 44 297 80 323
rect 106 297 112 323
rect -112 261 112 297
rect -112 235 -106 261
rect -80 235 -44 261
rect -18 235 18 261
rect 44 235 80 261
rect 106 235 112 261
rect -112 199 112 235
rect -112 173 -106 199
rect -80 173 -44 199
rect -18 173 18 199
rect 44 173 80 199
rect 106 173 112 199
rect -112 137 112 173
rect -112 111 -106 137
rect -80 111 -44 137
rect -18 111 18 137
rect 44 111 80 137
rect 106 111 112 137
rect -112 75 112 111
rect -112 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 112 75
rect -112 13 112 49
rect -112 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 112 13
rect -112 -49 112 -13
rect -112 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 112 -49
rect -112 -111 112 -75
rect -112 -137 -106 -111
rect -80 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 80 -111
rect 106 -137 112 -111
rect -112 -173 112 -137
rect -112 -199 -106 -173
rect -80 -199 -44 -173
rect -18 -199 18 -173
rect 44 -199 80 -173
rect 106 -199 112 -173
rect -112 -235 112 -199
rect -112 -261 -106 -235
rect -80 -261 -44 -235
rect -18 -261 18 -235
rect 44 -261 80 -235
rect 106 -261 112 -235
rect -112 -297 112 -261
rect -112 -323 -106 -297
rect -80 -323 -44 -297
rect -18 -323 18 -297
rect 44 -323 80 -297
rect 106 -323 112 -297
rect -112 -359 112 -323
rect -112 -385 -106 -359
rect -80 -385 -44 -359
rect -18 -385 18 -359
rect 44 -385 80 -359
rect 106 -385 112 -359
rect -112 -421 112 -385
rect -112 -447 -106 -421
rect -80 -447 -44 -421
rect -18 -447 18 -421
rect 44 -447 80 -421
rect 106 -447 112 -421
rect -112 -483 112 -447
rect -112 -509 -106 -483
rect -80 -509 -44 -483
rect -18 -509 18 -483
rect 44 -509 80 -483
rect 106 -509 112 -483
rect -112 -545 112 -509
rect -112 -571 -106 -545
rect -80 -571 -44 -545
rect -18 -571 18 -545
rect 44 -571 80 -545
rect 106 -571 112 -545
rect -112 -607 112 -571
rect -112 -633 -106 -607
rect -80 -633 -44 -607
rect -18 -633 18 -607
rect 44 -633 80 -607
rect 106 -633 112 -607
rect -112 -669 112 -633
rect -112 -695 -106 -669
rect -80 -695 -44 -669
rect -18 -695 18 -669
rect 44 -695 80 -669
rect 106 -695 112 -669
rect -112 -731 112 -695
rect -112 -757 -106 -731
rect -80 -757 -44 -731
rect -18 -757 18 -731
rect 44 -757 80 -731
rect 106 -757 112 -731
rect -112 -763 112 -757
<< via1 >>
rect -106 731 -80 757
rect -44 731 -18 757
rect 18 731 44 757
rect 80 731 106 757
rect -106 669 -80 695
rect -44 669 -18 695
rect 18 669 44 695
rect 80 669 106 695
rect -106 607 -80 633
rect -44 607 -18 633
rect 18 607 44 633
rect 80 607 106 633
rect -106 545 -80 571
rect -44 545 -18 571
rect 18 545 44 571
rect 80 545 106 571
rect -106 483 -80 509
rect -44 483 -18 509
rect 18 483 44 509
rect 80 483 106 509
rect -106 421 -80 447
rect -44 421 -18 447
rect 18 421 44 447
rect 80 421 106 447
rect -106 359 -80 385
rect -44 359 -18 385
rect 18 359 44 385
rect 80 359 106 385
rect -106 297 -80 323
rect -44 297 -18 323
rect 18 297 44 323
rect 80 297 106 323
rect -106 235 -80 261
rect -44 235 -18 261
rect 18 235 44 261
rect 80 235 106 261
rect -106 173 -80 199
rect -44 173 -18 199
rect 18 173 44 199
rect 80 173 106 199
rect -106 111 -80 137
rect -44 111 -18 137
rect 18 111 44 137
rect 80 111 106 137
rect -106 49 -80 75
rect -44 49 -18 75
rect 18 49 44 75
rect 80 49 106 75
rect -106 -13 -80 13
rect -44 -13 -18 13
rect 18 -13 44 13
rect 80 -13 106 13
rect -106 -75 -80 -49
rect -44 -75 -18 -49
rect 18 -75 44 -49
rect 80 -75 106 -49
rect -106 -137 -80 -111
rect -44 -137 -18 -111
rect 18 -137 44 -111
rect 80 -137 106 -111
rect -106 -199 -80 -173
rect -44 -199 -18 -173
rect 18 -199 44 -173
rect 80 -199 106 -173
rect -106 -261 -80 -235
rect -44 -261 -18 -235
rect 18 -261 44 -235
rect 80 -261 106 -235
rect -106 -323 -80 -297
rect -44 -323 -18 -297
rect 18 -323 44 -297
rect 80 -323 106 -297
rect -106 -385 -80 -359
rect -44 -385 -18 -359
rect 18 -385 44 -359
rect 80 -385 106 -359
rect -106 -447 -80 -421
rect -44 -447 -18 -421
rect 18 -447 44 -421
rect 80 -447 106 -421
rect -106 -509 -80 -483
rect -44 -509 -18 -483
rect 18 -509 44 -483
rect 80 -509 106 -483
rect -106 -571 -80 -545
rect -44 -571 -18 -545
rect 18 -571 44 -545
rect 80 -571 106 -545
rect -106 -633 -80 -607
rect -44 -633 -18 -607
rect 18 -633 44 -607
rect 80 -633 106 -607
rect -106 -695 -80 -669
rect -44 -695 -18 -669
rect 18 -695 44 -669
rect 80 -695 106 -669
rect -106 -757 -80 -731
rect -44 -757 -18 -731
rect 18 -757 44 -731
rect 80 -757 106 -731
<< metal2 >>
rect -112 757 112 763
rect -112 731 -106 757
rect -80 731 -44 757
rect -18 731 18 757
rect 44 731 80 757
rect 106 731 112 757
rect -112 695 112 731
rect -112 669 -106 695
rect -80 669 -44 695
rect -18 669 18 695
rect 44 669 80 695
rect 106 669 112 695
rect -112 633 112 669
rect -112 607 -106 633
rect -80 607 -44 633
rect -18 607 18 633
rect 44 607 80 633
rect 106 607 112 633
rect -112 571 112 607
rect -112 545 -106 571
rect -80 545 -44 571
rect -18 545 18 571
rect 44 545 80 571
rect 106 545 112 571
rect -112 509 112 545
rect -112 483 -106 509
rect -80 483 -44 509
rect -18 483 18 509
rect 44 483 80 509
rect 106 483 112 509
rect -112 447 112 483
rect -112 421 -106 447
rect -80 421 -44 447
rect -18 421 18 447
rect 44 421 80 447
rect 106 421 112 447
rect -112 385 112 421
rect -112 359 -106 385
rect -80 359 -44 385
rect -18 359 18 385
rect 44 359 80 385
rect 106 359 112 385
rect -112 323 112 359
rect -112 297 -106 323
rect -80 297 -44 323
rect -18 297 18 323
rect 44 297 80 323
rect 106 297 112 323
rect -112 261 112 297
rect -112 235 -106 261
rect -80 235 -44 261
rect -18 235 18 261
rect 44 235 80 261
rect 106 235 112 261
rect -112 199 112 235
rect -112 173 -106 199
rect -80 173 -44 199
rect -18 173 18 199
rect 44 173 80 199
rect 106 173 112 199
rect -112 137 112 173
rect -112 111 -106 137
rect -80 111 -44 137
rect -18 111 18 137
rect 44 111 80 137
rect 106 111 112 137
rect -112 75 112 111
rect -112 49 -106 75
rect -80 49 -44 75
rect -18 49 18 75
rect 44 49 80 75
rect 106 49 112 75
rect -112 13 112 49
rect -112 -13 -106 13
rect -80 -13 -44 13
rect -18 -13 18 13
rect 44 -13 80 13
rect 106 -13 112 13
rect -112 -49 112 -13
rect -112 -75 -106 -49
rect -80 -75 -44 -49
rect -18 -75 18 -49
rect 44 -75 80 -49
rect 106 -75 112 -49
rect -112 -111 112 -75
rect -112 -137 -106 -111
rect -80 -137 -44 -111
rect -18 -137 18 -111
rect 44 -137 80 -111
rect 106 -137 112 -111
rect -112 -173 112 -137
rect -112 -199 -106 -173
rect -80 -199 -44 -173
rect -18 -199 18 -173
rect 44 -199 80 -173
rect 106 -199 112 -173
rect -112 -235 112 -199
rect -112 -261 -106 -235
rect -80 -261 -44 -235
rect -18 -261 18 -235
rect 44 -261 80 -235
rect 106 -261 112 -235
rect -112 -297 112 -261
rect -112 -323 -106 -297
rect -80 -323 -44 -297
rect -18 -323 18 -297
rect 44 -323 80 -297
rect 106 -323 112 -297
rect -112 -359 112 -323
rect -112 -385 -106 -359
rect -80 -385 -44 -359
rect -18 -385 18 -359
rect 44 -385 80 -359
rect 106 -385 112 -359
rect -112 -421 112 -385
rect -112 -447 -106 -421
rect -80 -447 -44 -421
rect -18 -447 18 -421
rect 44 -447 80 -421
rect 106 -447 112 -421
rect -112 -483 112 -447
rect -112 -509 -106 -483
rect -80 -509 -44 -483
rect -18 -509 18 -483
rect 44 -509 80 -483
rect 106 -509 112 -483
rect -112 -545 112 -509
rect -112 -571 -106 -545
rect -80 -571 -44 -545
rect -18 -571 18 -545
rect 44 -571 80 -545
rect 106 -571 112 -545
rect -112 -607 112 -571
rect -112 -633 -106 -607
rect -80 -633 -44 -607
rect -18 -633 18 -607
rect 44 -633 80 -607
rect 106 -633 112 -607
rect -112 -669 112 -633
rect -112 -695 -106 -669
rect -80 -695 -44 -669
rect -18 -695 18 -669
rect 44 -695 80 -669
rect 106 -695 112 -669
rect -112 -731 112 -695
rect -112 -757 -106 -731
rect -80 -757 -44 -731
rect -18 -757 18 -731
rect 44 -757 80 -731
rect 106 -757 112 -731
rect -112 -763 112 -757
<< end >>
