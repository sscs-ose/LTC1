magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2360 -3465 15796 29678
<< isosubstrate >>
rect -257 10974 13760 27678
rect -39 -129 13470 10974
<< metal1 >>
rect -360 8855 61 10914
rect 843 10058 1780 10854
rect 11780 10058 12701 10854
rect 13375 8877 13796 10914
rect -360 8434 1108 8855
rect 1741 1243 2142 8863
rect 11290 1243 11732 8863
rect 12368 8456 13796 8877
rect 1741 510 2127 1243
rect 11316 770 11732 1243
rect 11290 510 11732 770
<< metal2 >>
rect 213 9051 313 26936
rect 393 9211 493 26936
rect 573 9371 673 26936
rect 753 9539 861 26936
rect 1697 26000 11781 26600
rect 1697 23319 2941 26000
rect 3465 23319 4709 26000
rect 5233 23319 6477 26000
rect 7001 23319 8245 26000
rect 8769 23319 10013 26000
rect 10537 23319 11781 26000
rect 1697 12658 2941 15319
rect 3465 12658 4709 15319
rect 5233 12658 6477 15319
rect 7001 12658 8245 15319
rect 8769 12658 10013 15319
rect 10537 12658 11781 15319
rect 753 9431 1206 9539
rect 573 9271 1206 9371
rect 393 9111 1206 9211
rect 213 8951 1206 9051
rect 1313 8943 12165 12658
rect 12617 9539 12725 26936
rect 12305 9431 12725 9539
rect 12805 9371 12905 26936
rect 12305 9271 12905 9371
rect 12985 9211 13085 26936
rect 12305 9111 13085 9211
rect 13165 9051 13265 26936
rect 12305 8951 13265 9051
rect 1313 -1210 1663 8943
rect 1741 510 2142 8863
rect 2372 -1210 4016 8943
rect 4720 -1210 6364 8943
rect 7069 -1210 8713 8943
rect 9416 -1210 11060 8943
rect 11290 510 11732 8863
rect 11831 -1465 12165 8943
use comp018green_out_paddrv_4T_NMOS_GROUP  comp018green_out_paddrv_4T_NMOS_GROUP_0
timestamp 1713338890
transform 1 0 1339 0 1 31
box -1367 -147 12129 10917
use comp018green_out_paddrv_4T_PMOS_GROUP  comp018green_out_paddrv_4T_PMOS_GROUP_0
timestamp 1713338890
transform 1 0 548 0 1 12347
box -767 -1312 13147 15294
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_0
timestamp 1713338890
transform 0 -1 1116 1 0 9158
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_1
timestamp 1713338890
transform 0 -1 1116 1 0 8992
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_2
timestamp 1713338890
transform 0 1 12395 1 0 8992
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_3
timestamp 1713338890
transform 0 1 12395 1 0 9158
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_4
timestamp 1713338890
transform 0 -1 1116 1 0 9318
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_5
timestamp 1713338890
transform 0 -1 1116 1 0 9484
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_6
timestamp 1713338890
transform 0 1 12395 1 0 9318
box -38 -90 38 90
use M2_M1_CDNS_69033583165570  M2_M1_CDNS_69033583165570_7
timestamp 1713338890
transform 0 1 12395 1 0 9484
box -38 -90 38 90
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_0
timestamp 1713338890
transform 1 0 1779 0 1 7701
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165579  M2_M1_CDNS_69033583165579_1
timestamp 1713338890
transform -1 0 11653 0 1 7701
box -38 -1130 38 1130
use M2_M1_CDNS_69033583165660  M2_M1_CDNS_69033583165660_0
timestamp 1713338890
transform 1 0 -150 0 1 10270
box -142 -506 142 506
use M2_M1_CDNS_69033583165660  M2_M1_CDNS_69033583165660_1
timestamp 1713338890
transform -1 0 13592 0 1 10270
box -142 -506 142 506
use M2_M1_CDNS_69033583165661  M2_M1_CDNS_69033583165661_0
timestamp 1713338890
transform 1 0 1089 0 1 10293
box -100 -534 100 534
use M2_M1_CDNS_69033583165661  M2_M1_CDNS_69033583165661_1
timestamp 1713338890
transform 1 0 12407 0 1 10293
box -100 -534 100 534
use M2_M1_CDNS_69033583165665  M2_M1_CDNS_69033583165665_0
timestamp 1713338890
transform 1 0 1779 0 1 1812
box -38 -1286 38 1286
use M2_M1_CDNS_69033583165665  M2_M1_CDNS_69033583165665_1
timestamp 1713338890
transform -1 0 11653 0 1 1812
box -38 -1286 38 1286
use M2_M1_CDNS_69033583165666  M2_M1_CDNS_69033583165666_0
timestamp 1713338890
transform 1 0 1779 0 1 4843
box -38 -1442 38 1442
use M2_M1_CDNS_69033583165666  M2_M1_CDNS_69033583165666_1
timestamp 1713338890
transform -1 0 11653 0 1 4843
box -38 -1442 38 1442
use M3_M2_CDNS_69033583165632  M3_M2_CDNS_69033583165632_0
timestamp 1713338890
transform 1 0 -146 0 1 10293
box -180 -535 180 535
use M3_M2_CDNS_69033583165632  M3_M2_CDNS_69033583165632_1
timestamp 1713338890
transform -1 0 13588 0 1 10293
box -180 -535 180 535
use M3_M2_CDNS_69033583165659  M3_M2_CDNS_69033583165659_0
timestamp 1713338890
transform 1 0 1089 0 1 10293
box -109 -535 109 535
use M3_M2_CDNS_69033583165659  M3_M2_CDNS_69033583165659_1
timestamp 1713338890
transform 1 0 12407 0 1 10293
box -109 -535 109 535
use M3_M2_CDNS_69033583165662  M3_M2_CDNS_69033583165662_0
timestamp 1713338890
transform 1 0 1779 0 1 1831
box -38 -870 38 870
use M3_M2_CDNS_69033583165662  M3_M2_CDNS_69033583165662_1
timestamp 1713338890
transform -1 0 11653 0 1 1831
box -38 -870 38 870
use M3_M2_CDNS_69033583165663  M3_M2_CDNS_69033583165663_0
timestamp 1713338890
transform 1 0 1779 0 1 4834
box -38 -1078 38 1078
use M3_M2_CDNS_69033583165663  M3_M2_CDNS_69033583165663_1
timestamp 1713338890
transform -1 0 11653 0 1 4834
box -38 -1078 38 1078
use M3_M2_CDNS_69033583165664  M3_M2_CDNS_69033583165664_0
timestamp 1713338890
transform 1 0 1779 0 1 7696
box -38 -818 38 818
use M3_M2_CDNS_69033583165664  M3_M2_CDNS_69033583165664_1
timestamp 1713338890
transform -1 0 11653 0 1 7696
box -38 -818 38 818
<< end >>
