magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2535 -2038 2535 2038
<< metal2 >>
rect -535 28 535 38
rect -535 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 535 28
rect -535 -38 535 -28
<< via2 >>
rect -525 -28 -469 28
rect -383 -28 -327 28
rect -241 -28 -185 28
rect -99 -28 -43 28
rect 43 -28 99 28
rect 185 -28 241 28
rect 327 -28 383 28
rect 469 -28 525 28
<< metal3 >>
rect -535 28 535 38
rect -535 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 535 28
rect -535 -38 535 -28
<< end >>
