magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3471 -2975 3471 2975
<< psubdiff >>
rect -1471 953 1471 975
rect -1471 907 -1449 953
rect -1403 907 -1325 953
rect -1279 907 -1201 953
rect -1155 907 -1077 953
rect -1031 907 -953 953
rect -907 907 -829 953
rect -783 907 -705 953
rect -659 907 -581 953
rect -535 907 -457 953
rect -411 907 -333 953
rect -287 907 -209 953
rect -163 907 -85 953
rect -39 907 39 953
rect 85 907 163 953
rect 209 907 287 953
rect 333 907 411 953
rect 457 907 535 953
rect 581 907 659 953
rect 705 907 783 953
rect 829 907 907 953
rect 953 907 1031 953
rect 1077 907 1155 953
rect 1201 907 1279 953
rect 1325 907 1403 953
rect 1449 907 1471 953
rect -1471 829 1471 907
rect -1471 783 -1449 829
rect -1403 783 -1325 829
rect -1279 783 -1201 829
rect -1155 783 -1077 829
rect -1031 783 -953 829
rect -907 783 -829 829
rect -783 783 -705 829
rect -659 783 -581 829
rect -535 783 -457 829
rect -411 783 -333 829
rect -287 783 -209 829
rect -163 783 -85 829
rect -39 783 39 829
rect 85 783 163 829
rect 209 783 287 829
rect 333 783 411 829
rect 457 783 535 829
rect 581 783 659 829
rect 705 783 783 829
rect 829 783 907 829
rect 953 783 1031 829
rect 1077 783 1155 829
rect 1201 783 1279 829
rect 1325 783 1403 829
rect 1449 783 1471 829
rect -1471 705 1471 783
rect -1471 659 -1449 705
rect -1403 659 -1325 705
rect -1279 659 -1201 705
rect -1155 659 -1077 705
rect -1031 659 -953 705
rect -907 659 -829 705
rect -783 659 -705 705
rect -659 659 -581 705
rect -535 659 -457 705
rect -411 659 -333 705
rect -287 659 -209 705
rect -163 659 -85 705
rect -39 659 39 705
rect 85 659 163 705
rect 209 659 287 705
rect 333 659 411 705
rect 457 659 535 705
rect 581 659 659 705
rect 705 659 783 705
rect 829 659 907 705
rect 953 659 1031 705
rect 1077 659 1155 705
rect 1201 659 1279 705
rect 1325 659 1403 705
rect 1449 659 1471 705
rect -1471 581 1471 659
rect -1471 535 -1449 581
rect -1403 535 -1325 581
rect -1279 535 -1201 581
rect -1155 535 -1077 581
rect -1031 535 -953 581
rect -907 535 -829 581
rect -783 535 -705 581
rect -659 535 -581 581
rect -535 535 -457 581
rect -411 535 -333 581
rect -287 535 -209 581
rect -163 535 -85 581
rect -39 535 39 581
rect 85 535 163 581
rect 209 535 287 581
rect 333 535 411 581
rect 457 535 535 581
rect 581 535 659 581
rect 705 535 783 581
rect 829 535 907 581
rect 953 535 1031 581
rect 1077 535 1155 581
rect 1201 535 1279 581
rect 1325 535 1403 581
rect 1449 535 1471 581
rect -1471 457 1471 535
rect -1471 411 -1449 457
rect -1403 411 -1325 457
rect -1279 411 -1201 457
rect -1155 411 -1077 457
rect -1031 411 -953 457
rect -907 411 -829 457
rect -783 411 -705 457
rect -659 411 -581 457
rect -535 411 -457 457
rect -411 411 -333 457
rect -287 411 -209 457
rect -163 411 -85 457
rect -39 411 39 457
rect 85 411 163 457
rect 209 411 287 457
rect 333 411 411 457
rect 457 411 535 457
rect 581 411 659 457
rect 705 411 783 457
rect 829 411 907 457
rect 953 411 1031 457
rect 1077 411 1155 457
rect 1201 411 1279 457
rect 1325 411 1403 457
rect 1449 411 1471 457
rect -1471 333 1471 411
rect -1471 287 -1449 333
rect -1403 287 -1325 333
rect -1279 287 -1201 333
rect -1155 287 -1077 333
rect -1031 287 -953 333
rect -907 287 -829 333
rect -783 287 -705 333
rect -659 287 -581 333
rect -535 287 -457 333
rect -411 287 -333 333
rect -287 287 -209 333
rect -163 287 -85 333
rect -39 287 39 333
rect 85 287 163 333
rect 209 287 287 333
rect 333 287 411 333
rect 457 287 535 333
rect 581 287 659 333
rect 705 287 783 333
rect 829 287 907 333
rect 953 287 1031 333
rect 1077 287 1155 333
rect 1201 287 1279 333
rect 1325 287 1403 333
rect 1449 287 1471 333
rect -1471 209 1471 287
rect -1471 163 -1449 209
rect -1403 163 -1325 209
rect -1279 163 -1201 209
rect -1155 163 -1077 209
rect -1031 163 -953 209
rect -907 163 -829 209
rect -783 163 -705 209
rect -659 163 -581 209
rect -535 163 -457 209
rect -411 163 -333 209
rect -287 163 -209 209
rect -163 163 -85 209
rect -39 163 39 209
rect 85 163 163 209
rect 209 163 287 209
rect 333 163 411 209
rect 457 163 535 209
rect 581 163 659 209
rect 705 163 783 209
rect 829 163 907 209
rect 953 163 1031 209
rect 1077 163 1155 209
rect 1201 163 1279 209
rect 1325 163 1403 209
rect 1449 163 1471 209
rect -1471 85 1471 163
rect -1471 39 -1449 85
rect -1403 39 -1325 85
rect -1279 39 -1201 85
rect -1155 39 -1077 85
rect -1031 39 -953 85
rect -907 39 -829 85
rect -783 39 -705 85
rect -659 39 -581 85
rect -535 39 -457 85
rect -411 39 -333 85
rect -287 39 -209 85
rect -163 39 -85 85
rect -39 39 39 85
rect 85 39 163 85
rect 209 39 287 85
rect 333 39 411 85
rect 457 39 535 85
rect 581 39 659 85
rect 705 39 783 85
rect 829 39 907 85
rect 953 39 1031 85
rect 1077 39 1155 85
rect 1201 39 1279 85
rect 1325 39 1403 85
rect 1449 39 1471 85
rect -1471 -39 1471 39
rect -1471 -85 -1449 -39
rect -1403 -85 -1325 -39
rect -1279 -85 -1201 -39
rect -1155 -85 -1077 -39
rect -1031 -85 -953 -39
rect -907 -85 -829 -39
rect -783 -85 -705 -39
rect -659 -85 -581 -39
rect -535 -85 -457 -39
rect -411 -85 -333 -39
rect -287 -85 -209 -39
rect -163 -85 -85 -39
rect -39 -85 39 -39
rect 85 -85 163 -39
rect 209 -85 287 -39
rect 333 -85 411 -39
rect 457 -85 535 -39
rect 581 -85 659 -39
rect 705 -85 783 -39
rect 829 -85 907 -39
rect 953 -85 1031 -39
rect 1077 -85 1155 -39
rect 1201 -85 1279 -39
rect 1325 -85 1403 -39
rect 1449 -85 1471 -39
rect -1471 -163 1471 -85
rect -1471 -209 -1449 -163
rect -1403 -209 -1325 -163
rect -1279 -209 -1201 -163
rect -1155 -209 -1077 -163
rect -1031 -209 -953 -163
rect -907 -209 -829 -163
rect -783 -209 -705 -163
rect -659 -209 -581 -163
rect -535 -209 -457 -163
rect -411 -209 -333 -163
rect -287 -209 -209 -163
rect -163 -209 -85 -163
rect -39 -209 39 -163
rect 85 -209 163 -163
rect 209 -209 287 -163
rect 333 -209 411 -163
rect 457 -209 535 -163
rect 581 -209 659 -163
rect 705 -209 783 -163
rect 829 -209 907 -163
rect 953 -209 1031 -163
rect 1077 -209 1155 -163
rect 1201 -209 1279 -163
rect 1325 -209 1403 -163
rect 1449 -209 1471 -163
rect -1471 -287 1471 -209
rect -1471 -333 -1449 -287
rect -1403 -333 -1325 -287
rect -1279 -333 -1201 -287
rect -1155 -333 -1077 -287
rect -1031 -333 -953 -287
rect -907 -333 -829 -287
rect -783 -333 -705 -287
rect -659 -333 -581 -287
rect -535 -333 -457 -287
rect -411 -333 -333 -287
rect -287 -333 -209 -287
rect -163 -333 -85 -287
rect -39 -333 39 -287
rect 85 -333 163 -287
rect 209 -333 287 -287
rect 333 -333 411 -287
rect 457 -333 535 -287
rect 581 -333 659 -287
rect 705 -333 783 -287
rect 829 -333 907 -287
rect 953 -333 1031 -287
rect 1077 -333 1155 -287
rect 1201 -333 1279 -287
rect 1325 -333 1403 -287
rect 1449 -333 1471 -287
rect -1471 -411 1471 -333
rect -1471 -457 -1449 -411
rect -1403 -457 -1325 -411
rect -1279 -457 -1201 -411
rect -1155 -457 -1077 -411
rect -1031 -457 -953 -411
rect -907 -457 -829 -411
rect -783 -457 -705 -411
rect -659 -457 -581 -411
rect -535 -457 -457 -411
rect -411 -457 -333 -411
rect -287 -457 -209 -411
rect -163 -457 -85 -411
rect -39 -457 39 -411
rect 85 -457 163 -411
rect 209 -457 287 -411
rect 333 -457 411 -411
rect 457 -457 535 -411
rect 581 -457 659 -411
rect 705 -457 783 -411
rect 829 -457 907 -411
rect 953 -457 1031 -411
rect 1077 -457 1155 -411
rect 1201 -457 1279 -411
rect 1325 -457 1403 -411
rect 1449 -457 1471 -411
rect -1471 -535 1471 -457
rect -1471 -581 -1449 -535
rect -1403 -581 -1325 -535
rect -1279 -581 -1201 -535
rect -1155 -581 -1077 -535
rect -1031 -581 -953 -535
rect -907 -581 -829 -535
rect -783 -581 -705 -535
rect -659 -581 -581 -535
rect -535 -581 -457 -535
rect -411 -581 -333 -535
rect -287 -581 -209 -535
rect -163 -581 -85 -535
rect -39 -581 39 -535
rect 85 -581 163 -535
rect 209 -581 287 -535
rect 333 -581 411 -535
rect 457 -581 535 -535
rect 581 -581 659 -535
rect 705 -581 783 -535
rect 829 -581 907 -535
rect 953 -581 1031 -535
rect 1077 -581 1155 -535
rect 1201 -581 1279 -535
rect 1325 -581 1403 -535
rect 1449 -581 1471 -535
rect -1471 -659 1471 -581
rect -1471 -705 -1449 -659
rect -1403 -705 -1325 -659
rect -1279 -705 -1201 -659
rect -1155 -705 -1077 -659
rect -1031 -705 -953 -659
rect -907 -705 -829 -659
rect -783 -705 -705 -659
rect -659 -705 -581 -659
rect -535 -705 -457 -659
rect -411 -705 -333 -659
rect -287 -705 -209 -659
rect -163 -705 -85 -659
rect -39 -705 39 -659
rect 85 -705 163 -659
rect 209 -705 287 -659
rect 333 -705 411 -659
rect 457 -705 535 -659
rect 581 -705 659 -659
rect 705 -705 783 -659
rect 829 -705 907 -659
rect 953 -705 1031 -659
rect 1077 -705 1155 -659
rect 1201 -705 1279 -659
rect 1325 -705 1403 -659
rect 1449 -705 1471 -659
rect -1471 -783 1471 -705
rect -1471 -829 -1449 -783
rect -1403 -829 -1325 -783
rect -1279 -829 -1201 -783
rect -1155 -829 -1077 -783
rect -1031 -829 -953 -783
rect -907 -829 -829 -783
rect -783 -829 -705 -783
rect -659 -829 -581 -783
rect -535 -829 -457 -783
rect -411 -829 -333 -783
rect -287 -829 -209 -783
rect -163 -829 -85 -783
rect -39 -829 39 -783
rect 85 -829 163 -783
rect 209 -829 287 -783
rect 333 -829 411 -783
rect 457 -829 535 -783
rect 581 -829 659 -783
rect 705 -829 783 -783
rect 829 -829 907 -783
rect 953 -829 1031 -783
rect 1077 -829 1155 -783
rect 1201 -829 1279 -783
rect 1325 -829 1403 -783
rect 1449 -829 1471 -783
rect -1471 -907 1471 -829
rect -1471 -953 -1449 -907
rect -1403 -953 -1325 -907
rect -1279 -953 -1201 -907
rect -1155 -953 -1077 -907
rect -1031 -953 -953 -907
rect -907 -953 -829 -907
rect -783 -953 -705 -907
rect -659 -953 -581 -907
rect -535 -953 -457 -907
rect -411 -953 -333 -907
rect -287 -953 -209 -907
rect -163 -953 -85 -907
rect -39 -953 39 -907
rect 85 -953 163 -907
rect 209 -953 287 -907
rect 333 -953 411 -907
rect 457 -953 535 -907
rect 581 -953 659 -907
rect 705 -953 783 -907
rect 829 -953 907 -907
rect 953 -953 1031 -907
rect 1077 -953 1155 -907
rect 1201 -953 1279 -907
rect 1325 -953 1403 -907
rect 1449 -953 1471 -907
rect -1471 -975 1471 -953
<< psubdiffcont >>
rect -1449 907 -1403 953
rect -1325 907 -1279 953
rect -1201 907 -1155 953
rect -1077 907 -1031 953
rect -953 907 -907 953
rect -829 907 -783 953
rect -705 907 -659 953
rect -581 907 -535 953
rect -457 907 -411 953
rect -333 907 -287 953
rect -209 907 -163 953
rect -85 907 -39 953
rect 39 907 85 953
rect 163 907 209 953
rect 287 907 333 953
rect 411 907 457 953
rect 535 907 581 953
rect 659 907 705 953
rect 783 907 829 953
rect 907 907 953 953
rect 1031 907 1077 953
rect 1155 907 1201 953
rect 1279 907 1325 953
rect 1403 907 1449 953
rect -1449 783 -1403 829
rect -1325 783 -1279 829
rect -1201 783 -1155 829
rect -1077 783 -1031 829
rect -953 783 -907 829
rect -829 783 -783 829
rect -705 783 -659 829
rect -581 783 -535 829
rect -457 783 -411 829
rect -333 783 -287 829
rect -209 783 -163 829
rect -85 783 -39 829
rect 39 783 85 829
rect 163 783 209 829
rect 287 783 333 829
rect 411 783 457 829
rect 535 783 581 829
rect 659 783 705 829
rect 783 783 829 829
rect 907 783 953 829
rect 1031 783 1077 829
rect 1155 783 1201 829
rect 1279 783 1325 829
rect 1403 783 1449 829
rect -1449 659 -1403 705
rect -1325 659 -1279 705
rect -1201 659 -1155 705
rect -1077 659 -1031 705
rect -953 659 -907 705
rect -829 659 -783 705
rect -705 659 -659 705
rect -581 659 -535 705
rect -457 659 -411 705
rect -333 659 -287 705
rect -209 659 -163 705
rect -85 659 -39 705
rect 39 659 85 705
rect 163 659 209 705
rect 287 659 333 705
rect 411 659 457 705
rect 535 659 581 705
rect 659 659 705 705
rect 783 659 829 705
rect 907 659 953 705
rect 1031 659 1077 705
rect 1155 659 1201 705
rect 1279 659 1325 705
rect 1403 659 1449 705
rect -1449 535 -1403 581
rect -1325 535 -1279 581
rect -1201 535 -1155 581
rect -1077 535 -1031 581
rect -953 535 -907 581
rect -829 535 -783 581
rect -705 535 -659 581
rect -581 535 -535 581
rect -457 535 -411 581
rect -333 535 -287 581
rect -209 535 -163 581
rect -85 535 -39 581
rect 39 535 85 581
rect 163 535 209 581
rect 287 535 333 581
rect 411 535 457 581
rect 535 535 581 581
rect 659 535 705 581
rect 783 535 829 581
rect 907 535 953 581
rect 1031 535 1077 581
rect 1155 535 1201 581
rect 1279 535 1325 581
rect 1403 535 1449 581
rect -1449 411 -1403 457
rect -1325 411 -1279 457
rect -1201 411 -1155 457
rect -1077 411 -1031 457
rect -953 411 -907 457
rect -829 411 -783 457
rect -705 411 -659 457
rect -581 411 -535 457
rect -457 411 -411 457
rect -333 411 -287 457
rect -209 411 -163 457
rect -85 411 -39 457
rect 39 411 85 457
rect 163 411 209 457
rect 287 411 333 457
rect 411 411 457 457
rect 535 411 581 457
rect 659 411 705 457
rect 783 411 829 457
rect 907 411 953 457
rect 1031 411 1077 457
rect 1155 411 1201 457
rect 1279 411 1325 457
rect 1403 411 1449 457
rect -1449 287 -1403 333
rect -1325 287 -1279 333
rect -1201 287 -1155 333
rect -1077 287 -1031 333
rect -953 287 -907 333
rect -829 287 -783 333
rect -705 287 -659 333
rect -581 287 -535 333
rect -457 287 -411 333
rect -333 287 -287 333
rect -209 287 -163 333
rect -85 287 -39 333
rect 39 287 85 333
rect 163 287 209 333
rect 287 287 333 333
rect 411 287 457 333
rect 535 287 581 333
rect 659 287 705 333
rect 783 287 829 333
rect 907 287 953 333
rect 1031 287 1077 333
rect 1155 287 1201 333
rect 1279 287 1325 333
rect 1403 287 1449 333
rect -1449 163 -1403 209
rect -1325 163 -1279 209
rect -1201 163 -1155 209
rect -1077 163 -1031 209
rect -953 163 -907 209
rect -829 163 -783 209
rect -705 163 -659 209
rect -581 163 -535 209
rect -457 163 -411 209
rect -333 163 -287 209
rect -209 163 -163 209
rect -85 163 -39 209
rect 39 163 85 209
rect 163 163 209 209
rect 287 163 333 209
rect 411 163 457 209
rect 535 163 581 209
rect 659 163 705 209
rect 783 163 829 209
rect 907 163 953 209
rect 1031 163 1077 209
rect 1155 163 1201 209
rect 1279 163 1325 209
rect 1403 163 1449 209
rect -1449 39 -1403 85
rect -1325 39 -1279 85
rect -1201 39 -1155 85
rect -1077 39 -1031 85
rect -953 39 -907 85
rect -829 39 -783 85
rect -705 39 -659 85
rect -581 39 -535 85
rect -457 39 -411 85
rect -333 39 -287 85
rect -209 39 -163 85
rect -85 39 -39 85
rect 39 39 85 85
rect 163 39 209 85
rect 287 39 333 85
rect 411 39 457 85
rect 535 39 581 85
rect 659 39 705 85
rect 783 39 829 85
rect 907 39 953 85
rect 1031 39 1077 85
rect 1155 39 1201 85
rect 1279 39 1325 85
rect 1403 39 1449 85
rect -1449 -85 -1403 -39
rect -1325 -85 -1279 -39
rect -1201 -85 -1155 -39
rect -1077 -85 -1031 -39
rect -953 -85 -907 -39
rect -829 -85 -783 -39
rect -705 -85 -659 -39
rect -581 -85 -535 -39
rect -457 -85 -411 -39
rect -333 -85 -287 -39
rect -209 -85 -163 -39
rect -85 -85 -39 -39
rect 39 -85 85 -39
rect 163 -85 209 -39
rect 287 -85 333 -39
rect 411 -85 457 -39
rect 535 -85 581 -39
rect 659 -85 705 -39
rect 783 -85 829 -39
rect 907 -85 953 -39
rect 1031 -85 1077 -39
rect 1155 -85 1201 -39
rect 1279 -85 1325 -39
rect 1403 -85 1449 -39
rect -1449 -209 -1403 -163
rect -1325 -209 -1279 -163
rect -1201 -209 -1155 -163
rect -1077 -209 -1031 -163
rect -953 -209 -907 -163
rect -829 -209 -783 -163
rect -705 -209 -659 -163
rect -581 -209 -535 -163
rect -457 -209 -411 -163
rect -333 -209 -287 -163
rect -209 -209 -163 -163
rect -85 -209 -39 -163
rect 39 -209 85 -163
rect 163 -209 209 -163
rect 287 -209 333 -163
rect 411 -209 457 -163
rect 535 -209 581 -163
rect 659 -209 705 -163
rect 783 -209 829 -163
rect 907 -209 953 -163
rect 1031 -209 1077 -163
rect 1155 -209 1201 -163
rect 1279 -209 1325 -163
rect 1403 -209 1449 -163
rect -1449 -333 -1403 -287
rect -1325 -333 -1279 -287
rect -1201 -333 -1155 -287
rect -1077 -333 -1031 -287
rect -953 -333 -907 -287
rect -829 -333 -783 -287
rect -705 -333 -659 -287
rect -581 -333 -535 -287
rect -457 -333 -411 -287
rect -333 -333 -287 -287
rect -209 -333 -163 -287
rect -85 -333 -39 -287
rect 39 -333 85 -287
rect 163 -333 209 -287
rect 287 -333 333 -287
rect 411 -333 457 -287
rect 535 -333 581 -287
rect 659 -333 705 -287
rect 783 -333 829 -287
rect 907 -333 953 -287
rect 1031 -333 1077 -287
rect 1155 -333 1201 -287
rect 1279 -333 1325 -287
rect 1403 -333 1449 -287
rect -1449 -457 -1403 -411
rect -1325 -457 -1279 -411
rect -1201 -457 -1155 -411
rect -1077 -457 -1031 -411
rect -953 -457 -907 -411
rect -829 -457 -783 -411
rect -705 -457 -659 -411
rect -581 -457 -535 -411
rect -457 -457 -411 -411
rect -333 -457 -287 -411
rect -209 -457 -163 -411
rect -85 -457 -39 -411
rect 39 -457 85 -411
rect 163 -457 209 -411
rect 287 -457 333 -411
rect 411 -457 457 -411
rect 535 -457 581 -411
rect 659 -457 705 -411
rect 783 -457 829 -411
rect 907 -457 953 -411
rect 1031 -457 1077 -411
rect 1155 -457 1201 -411
rect 1279 -457 1325 -411
rect 1403 -457 1449 -411
rect -1449 -581 -1403 -535
rect -1325 -581 -1279 -535
rect -1201 -581 -1155 -535
rect -1077 -581 -1031 -535
rect -953 -581 -907 -535
rect -829 -581 -783 -535
rect -705 -581 -659 -535
rect -581 -581 -535 -535
rect -457 -581 -411 -535
rect -333 -581 -287 -535
rect -209 -581 -163 -535
rect -85 -581 -39 -535
rect 39 -581 85 -535
rect 163 -581 209 -535
rect 287 -581 333 -535
rect 411 -581 457 -535
rect 535 -581 581 -535
rect 659 -581 705 -535
rect 783 -581 829 -535
rect 907 -581 953 -535
rect 1031 -581 1077 -535
rect 1155 -581 1201 -535
rect 1279 -581 1325 -535
rect 1403 -581 1449 -535
rect -1449 -705 -1403 -659
rect -1325 -705 -1279 -659
rect -1201 -705 -1155 -659
rect -1077 -705 -1031 -659
rect -953 -705 -907 -659
rect -829 -705 -783 -659
rect -705 -705 -659 -659
rect -581 -705 -535 -659
rect -457 -705 -411 -659
rect -333 -705 -287 -659
rect -209 -705 -163 -659
rect -85 -705 -39 -659
rect 39 -705 85 -659
rect 163 -705 209 -659
rect 287 -705 333 -659
rect 411 -705 457 -659
rect 535 -705 581 -659
rect 659 -705 705 -659
rect 783 -705 829 -659
rect 907 -705 953 -659
rect 1031 -705 1077 -659
rect 1155 -705 1201 -659
rect 1279 -705 1325 -659
rect 1403 -705 1449 -659
rect -1449 -829 -1403 -783
rect -1325 -829 -1279 -783
rect -1201 -829 -1155 -783
rect -1077 -829 -1031 -783
rect -953 -829 -907 -783
rect -829 -829 -783 -783
rect -705 -829 -659 -783
rect -581 -829 -535 -783
rect -457 -829 -411 -783
rect -333 -829 -287 -783
rect -209 -829 -163 -783
rect -85 -829 -39 -783
rect 39 -829 85 -783
rect 163 -829 209 -783
rect 287 -829 333 -783
rect 411 -829 457 -783
rect 535 -829 581 -783
rect 659 -829 705 -783
rect 783 -829 829 -783
rect 907 -829 953 -783
rect 1031 -829 1077 -783
rect 1155 -829 1201 -783
rect 1279 -829 1325 -783
rect 1403 -829 1449 -783
rect -1449 -953 -1403 -907
rect -1325 -953 -1279 -907
rect -1201 -953 -1155 -907
rect -1077 -953 -1031 -907
rect -953 -953 -907 -907
rect -829 -953 -783 -907
rect -705 -953 -659 -907
rect -581 -953 -535 -907
rect -457 -953 -411 -907
rect -333 -953 -287 -907
rect -209 -953 -163 -907
rect -85 -953 -39 -907
rect 39 -953 85 -907
rect 163 -953 209 -907
rect 287 -953 333 -907
rect 411 -953 457 -907
rect 535 -953 581 -907
rect 659 -953 705 -907
rect 783 -953 829 -907
rect 907 -953 953 -907
rect 1031 -953 1077 -907
rect 1155 -953 1201 -907
rect 1279 -953 1325 -907
rect 1403 -953 1449 -907
<< metal1 >>
rect -1460 953 1460 964
rect -1460 907 -1449 953
rect -1403 907 -1325 953
rect -1279 907 -1201 953
rect -1155 907 -1077 953
rect -1031 907 -953 953
rect -907 907 -829 953
rect -783 907 -705 953
rect -659 907 -581 953
rect -535 907 -457 953
rect -411 907 -333 953
rect -287 907 -209 953
rect -163 907 -85 953
rect -39 907 39 953
rect 85 907 163 953
rect 209 907 287 953
rect 333 907 411 953
rect 457 907 535 953
rect 581 907 659 953
rect 705 907 783 953
rect 829 907 907 953
rect 953 907 1031 953
rect 1077 907 1155 953
rect 1201 907 1279 953
rect 1325 907 1403 953
rect 1449 907 1460 953
rect -1460 829 1460 907
rect -1460 783 -1449 829
rect -1403 783 -1325 829
rect -1279 783 -1201 829
rect -1155 783 -1077 829
rect -1031 783 -953 829
rect -907 783 -829 829
rect -783 783 -705 829
rect -659 783 -581 829
rect -535 783 -457 829
rect -411 783 -333 829
rect -287 783 -209 829
rect -163 783 -85 829
rect -39 783 39 829
rect 85 783 163 829
rect 209 783 287 829
rect 333 783 411 829
rect 457 783 535 829
rect 581 783 659 829
rect 705 783 783 829
rect 829 783 907 829
rect 953 783 1031 829
rect 1077 783 1155 829
rect 1201 783 1279 829
rect 1325 783 1403 829
rect 1449 783 1460 829
rect -1460 705 1460 783
rect -1460 659 -1449 705
rect -1403 659 -1325 705
rect -1279 659 -1201 705
rect -1155 659 -1077 705
rect -1031 659 -953 705
rect -907 659 -829 705
rect -783 659 -705 705
rect -659 659 -581 705
rect -535 659 -457 705
rect -411 659 -333 705
rect -287 659 -209 705
rect -163 659 -85 705
rect -39 659 39 705
rect 85 659 163 705
rect 209 659 287 705
rect 333 659 411 705
rect 457 659 535 705
rect 581 659 659 705
rect 705 659 783 705
rect 829 659 907 705
rect 953 659 1031 705
rect 1077 659 1155 705
rect 1201 659 1279 705
rect 1325 659 1403 705
rect 1449 659 1460 705
rect -1460 581 1460 659
rect -1460 535 -1449 581
rect -1403 535 -1325 581
rect -1279 535 -1201 581
rect -1155 535 -1077 581
rect -1031 535 -953 581
rect -907 535 -829 581
rect -783 535 -705 581
rect -659 535 -581 581
rect -535 535 -457 581
rect -411 535 -333 581
rect -287 535 -209 581
rect -163 535 -85 581
rect -39 535 39 581
rect 85 535 163 581
rect 209 535 287 581
rect 333 535 411 581
rect 457 535 535 581
rect 581 535 659 581
rect 705 535 783 581
rect 829 535 907 581
rect 953 535 1031 581
rect 1077 535 1155 581
rect 1201 535 1279 581
rect 1325 535 1403 581
rect 1449 535 1460 581
rect -1460 457 1460 535
rect -1460 411 -1449 457
rect -1403 411 -1325 457
rect -1279 411 -1201 457
rect -1155 411 -1077 457
rect -1031 411 -953 457
rect -907 411 -829 457
rect -783 411 -705 457
rect -659 411 -581 457
rect -535 411 -457 457
rect -411 411 -333 457
rect -287 411 -209 457
rect -163 411 -85 457
rect -39 411 39 457
rect 85 411 163 457
rect 209 411 287 457
rect 333 411 411 457
rect 457 411 535 457
rect 581 411 659 457
rect 705 411 783 457
rect 829 411 907 457
rect 953 411 1031 457
rect 1077 411 1155 457
rect 1201 411 1279 457
rect 1325 411 1403 457
rect 1449 411 1460 457
rect -1460 333 1460 411
rect -1460 287 -1449 333
rect -1403 287 -1325 333
rect -1279 287 -1201 333
rect -1155 287 -1077 333
rect -1031 287 -953 333
rect -907 287 -829 333
rect -783 287 -705 333
rect -659 287 -581 333
rect -535 287 -457 333
rect -411 287 -333 333
rect -287 287 -209 333
rect -163 287 -85 333
rect -39 287 39 333
rect 85 287 163 333
rect 209 287 287 333
rect 333 287 411 333
rect 457 287 535 333
rect 581 287 659 333
rect 705 287 783 333
rect 829 287 907 333
rect 953 287 1031 333
rect 1077 287 1155 333
rect 1201 287 1279 333
rect 1325 287 1403 333
rect 1449 287 1460 333
rect -1460 209 1460 287
rect -1460 163 -1449 209
rect -1403 163 -1325 209
rect -1279 163 -1201 209
rect -1155 163 -1077 209
rect -1031 163 -953 209
rect -907 163 -829 209
rect -783 163 -705 209
rect -659 163 -581 209
rect -535 163 -457 209
rect -411 163 -333 209
rect -287 163 -209 209
rect -163 163 -85 209
rect -39 163 39 209
rect 85 163 163 209
rect 209 163 287 209
rect 333 163 411 209
rect 457 163 535 209
rect 581 163 659 209
rect 705 163 783 209
rect 829 163 907 209
rect 953 163 1031 209
rect 1077 163 1155 209
rect 1201 163 1279 209
rect 1325 163 1403 209
rect 1449 163 1460 209
rect -1460 85 1460 163
rect -1460 39 -1449 85
rect -1403 39 -1325 85
rect -1279 39 -1201 85
rect -1155 39 -1077 85
rect -1031 39 -953 85
rect -907 39 -829 85
rect -783 39 -705 85
rect -659 39 -581 85
rect -535 39 -457 85
rect -411 39 -333 85
rect -287 39 -209 85
rect -163 39 -85 85
rect -39 39 39 85
rect 85 39 163 85
rect 209 39 287 85
rect 333 39 411 85
rect 457 39 535 85
rect 581 39 659 85
rect 705 39 783 85
rect 829 39 907 85
rect 953 39 1031 85
rect 1077 39 1155 85
rect 1201 39 1279 85
rect 1325 39 1403 85
rect 1449 39 1460 85
rect -1460 -39 1460 39
rect -1460 -85 -1449 -39
rect -1403 -85 -1325 -39
rect -1279 -85 -1201 -39
rect -1155 -85 -1077 -39
rect -1031 -85 -953 -39
rect -907 -85 -829 -39
rect -783 -85 -705 -39
rect -659 -85 -581 -39
rect -535 -85 -457 -39
rect -411 -85 -333 -39
rect -287 -85 -209 -39
rect -163 -85 -85 -39
rect -39 -85 39 -39
rect 85 -85 163 -39
rect 209 -85 287 -39
rect 333 -85 411 -39
rect 457 -85 535 -39
rect 581 -85 659 -39
rect 705 -85 783 -39
rect 829 -85 907 -39
rect 953 -85 1031 -39
rect 1077 -85 1155 -39
rect 1201 -85 1279 -39
rect 1325 -85 1403 -39
rect 1449 -85 1460 -39
rect -1460 -163 1460 -85
rect -1460 -209 -1449 -163
rect -1403 -209 -1325 -163
rect -1279 -209 -1201 -163
rect -1155 -209 -1077 -163
rect -1031 -209 -953 -163
rect -907 -209 -829 -163
rect -783 -209 -705 -163
rect -659 -209 -581 -163
rect -535 -209 -457 -163
rect -411 -209 -333 -163
rect -287 -209 -209 -163
rect -163 -209 -85 -163
rect -39 -209 39 -163
rect 85 -209 163 -163
rect 209 -209 287 -163
rect 333 -209 411 -163
rect 457 -209 535 -163
rect 581 -209 659 -163
rect 705 -209 783 -163
rect 829 -209 907 -163
rect 953 -209 1031 -163
rect 1077 -209 1155 -163
rect 1201 -209 1279 -163
rect 1325 -209 1403 -163
rect 1449 -209 1460 -163
rect -1460 -287 1460 -209
rect -1460 -333 -1449 -287
rect -1403 -333 -1325 -287
rect -1279 -333 -1201 -287
rect -1155 -333 -1077 -287
rect -1031 -333 -953 -287
rect -907 -333 -829 -287
rect -783 -333 -705 -287
rect -659 -333 -581 -287
rect -535 -333 -457 -287
rect -411 -333 -333 -287
rect -287 -333 -209 -287
rect -163 -333 -85 -287
rect -39 -333 39 -287
rect 85 -333 163 -287
rect 209 -333 287 -287
rect 333 -333 411 -287
rect 457 -333 535 -287
rect 581 -333 659 -287
rect 705 -333 783 -287
rect 829 -333 907 -287
rect 953 -333 1031 -287
rect 1077 -333 1155 -287
rect 1201 -333 1279 -287
rect 1325 -333 1403 -287
rect 1449 -333 1460 -287
rect -1460 -411 1460 -333
rect -1460 -457 -1449 -411
rect -1403 -457 -1325 -411
rect -1279 -457 -1201 -411
rect -1155 -457 -1077 -411
rect -1031 -457 -953 -411
rect -907 -457 -829 -411
rect -783 -457 -705 -411
rect -659 -457 -581 -411
rect -535 -457 -457 -411
rect -411 -457 -333 -411
rect -287 -457 -209 -411
rect -163 -457 -85 -411
rect -39 -457 39 -411
rect 85 -457 163 -411
rect 209 -457 287 -411
rect 333 -457 411 -411
rect 457 -457 535 -411
rect 581 -457 659 -411
rect 705 -457 783 -411
rect 829 -457 907 -411
rect 953 -457 1031 -411
rect 1077 -457 1155 -411
rect 1201 -457 1279 -411
rect 1325 -457 1403 -411
rect 1449 -457 1460 -411
rect -1460 -535 1460 -457
rect -1460 -581 -1449 -535
rect -1403 -581 -1325 -535
rect -1279 -581 -1201 -535
rect -1155 -581 -1077 -535
rect -1031 -581 -953 -535
rect -907 -581 -829 -535
rect -783 -581 -705 -535
rect -659 -581 -581 -535
rect -535 -581 -457 -535
rect -411 -581 -333 -535
rect -287 -581 -209 -535
rect -163 -581 -85 -535
rect -39 -581 39 -535
rect 85 -581 163 -535
rect 209 -581 287 -535
rect 333 -581 411 -535
rect 457 -581 535 -535
rect 581 -581 659 -535
rect 705 -581 783 -535
rect 829 -581 907 -535
rect 953 -581 1031 -535
rect 1077 -581 1155 -535
rect 1201 -581 1279 -535
rect 1325 -581 1403 -535
rect 1449 -581 1460 -535
rect -1460 -659 1460 -581
rect -1460 -705 -1449 -659
rect -1403 -705 -1325 -659
rect -1279 -705 -1201 -659
rect -1155 -705 -1077 -659
rect -1031 -705 -953 -659
rect -907 -705 -829 -659
rect -783 -705 -705 -659
rect -659 -705 -581 -659
rect -535 -705 -457 -659
rect -411 -705 -333 -659
rect -287 -705 -209 -659
rect -163 -705 -85 -659
rect -39 -705 39 -659
rect 85 -705 163 -659
rect 209 -705 287 -659
rect 333 -705 411 -659
rect 457 -705 535 -659
rect 581 -705 659 -659
rect 705 -705 783 -659
rect 829 -705 907 -659
rect 953 -705 1031 -659
rect 1077 -705 1155 -659
rect 1201 -705 1279 -659
rect 1325 -705 1403 -659
rect 1449 -705 1460 -659
rect -1460 -783 1460 -705
rect -1460 -829 -1449 -783
rect -1403 -829 -1325 -783
rect -1279 -829 -1201 -783
rect -1155 -829 -1077 -783
rect -1031 -829 -953 -783
rect -907 -829 -829 -783
rect -783 -829 -705 -783
rect -659 -829 -581 -783
rect -535 -829 -457 -783
rect -411 -829 -333 -783
rect -287 -829 -209 -783
rect -163 -829 -85 -783
rect -39 -829 39 -783
rect 85 -829 163 -783
rect 209 -829 287 -783
rect 333 -829 411 -783
rect 457 -829 535 -783
rect 581 -829 659 -783
rect 705 -829 783 -783
rect 829 -829 907 -783
rect 953 -829 1031 -783
rect 1077 -829 1155 -783
rect 1201 -829 1279 -783
rect 1325 -829 1403 -783
rect 1449 -829 1460 -783
rect -1460 -907 1460 -829
rect -1460 -953 -1449 -907
rect -1403 -953 -1325 -907
rect -1279 -953 -1201 -907
rect -1155 -953 -1077 -907
rect -1031 -953 -953 -907
rect -907 -953 -829 -907
rect -783 -953 -705 -907
rect -659 -953 -581 -907
rect -535 -953 -457 -907
rect -411 -953 -333 -907
rect -287 -953 -209 -907
rect -163 -953 -85 -907
rect -39 -953 39 -907
rect 85 -953 163 -907
rect 209 -953 287 -907
rect 333 -953 411 -907
rect 457 -953 535 -907
rect 581 -953 659 -907
rect 705 -953 783 -907
rect 829 -953 907 -907
rect 953 -953 1031 -907
rect 1077 -953 1155 -907
rect 1201 -953 1279 -907
rect 1325 -953 1403 -907
rect 1449 -953 1460 -907
rect -1460 -964 1460 -953
<< end >>
