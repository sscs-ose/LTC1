magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -2938 2045 2938
<< psubdiff >>
rect -45 916 45 938
rect -45 -916 -23 916
rect 23 -916 45 916
rect -45 -938 45 -916
<< psubdiffcont >>
rect -23 -916 23 916
<< metal1 >>
rect -34 916 34 927
rect -34 -916 -23 916
rect 23 -916 34 916
rect -34 -927 34 -916
<< end >>
