magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1565 1019 1565
<< metal1 >>
rect -19 559 19 565
rect -19 -559 -13 559
rect 13 -559 19 559
rect -19 -565 19 -559
<< via1 >>
rect -13 -559 13 559
<< metal2 >>
rect -19 559 19 565
rect -19 -559 -13 559
rect 13 -559 19 559
rect -19 -565 19 -559
<< end >>
