magic
tech gf180mcuC
magscale 1 10
timestamp 1694434822
<< nwell >>
rect -984 -406 984 406
<< nsubdiff >>
rect -960 310 960 382
rect -960 -310 -888 310
rect 888 -310 960 310
rect -960 -382 960 -310
<< polysilicon >>
rect -800 209 -600 222
rect -800 163 -787 209
rect -613 163 -600 209
rect -800 120 -600 163
rect -800 -163 -600 -120
rect -800 -209 -787 -163
rect -613 -209 -600 -163
rect -800 -222 -600 -209
rect -520 209 -320 222
rect -520 163 -507 209
rect -333 163 -320 209
rect -520 120 -320 163
rect -520 -163 -320 -120
rect -520 -209 -507 -163
rect -333 -209 -320 -163
rect -520 -222 -320 -209
rect -240 209 -40 222
rect -240 163 -227 209
rect -53 163 -40 209
rect -240 120 -40 163
rect -240 -163 -40 -120
rect -240 -209 -227 -163
rect -53 -209 -40 -163
rect -240 -222 -40 -209
rect 40 209 240 222
rect 40 163 53 209
rect 227 163 240 209
rect 40 120 240 163
rect 40 -163 240 -120
rect 40 -209 53 -163
rect 227 -209 240 -163
rect 40 -222 240 -209
rect 320 209 520 222
rect 320 163 333 209
rect 507 163 520 209
rect 320 120 520 163
rect 320 -163 520 -120
rect 320 -209 333 -163
rect 507 -209 520 -163
rect 320 -222 520 -209
rect 600 209 800 222
rect 600 163 613 209
rect 787 163 800 209
rect 600 120 800 163
rect 600 -163 800 -120
rect 600 -209 613 -163
rect 787 -209 800 -163
rect 600 -222 800 -209
<< polycontact >>
rect -787 163 -613 209
rect -787 -209 -613 -163
rect -507 163 -333 209
rect -507 -209 -333 -163
rect -227 163 -53 209
rect -227 -209 -53 -163
rect 53 163 227 209
rect 53 -209 227 -163
rect 333 163 507 209
rect 333 -209 507 -163
rect 613 163 787 209
rect 613 -209 787 -163
<< ppolyres >>
rect -800 -120 -600 120
rect -520 -120 -320 120
rect -240 -120 -40 120
rect 40 -120 240 120
rect 320 -120 520 120
rect 600 -120 800 120
<< metal1 >>
rect -798 163 -787 209
rect -613 163 -602 209
rect -518 163 -507 209
rect -333 163 -322 209
rect -238 163 -227 209
rect -53 163 -42 209
rect 42 163 53 209
rect 227 163 238 209
rect 322 163 333 209
rect 507 163 518 209
rect 602 163 613 209
rect 787 163 798 209
rect -798 -209 -787 -163
rect -613 -209 -602 -163
rect -518 -209 -507 -163
rect -333 -209 -322 -163
rect -238 -209 -227 -163
rect -53 -209 -42 -163
rect 42 -209 53 -163
rect 227 -209 238 -163
rect 322 -209 333 -163
rect 507 -209 518 -163
rect 602 -209 613 -163
rect 787 -209 798 -163
<< properties >>
string FIXED_BBOX -924 -346 924 346
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.0 l 1.2 m 1 nx 6 wmin 0.80 lmin 1.00 rho 315 val 406.451 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
