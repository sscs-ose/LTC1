magic
tech gf180mcuC
magscale 1 10
timestamp 1691396512
<< error_p >>
rect -823 542 -777 638
rect -663 542 -617 638
rect -503 542 -457 638
rect -343 542 -297 638
rect -183 542 -137 638
rect -23 542 23 638
rect 137 542 183 638
rect 297 542 343 638
rect 457 542 503 638
rect 617 542 663 638
rect 777 542 823 638
rect -823 306 -777 402
rect -663 306 -617 402
rect -503 306 -457 402
rect -343 306 -297 402
rect -183 306 -137 402
rect -23 306 23 402
rect 137 306 183 402
rect 297 306 343 402
rect 457 306 503 402
rect 617 306 663 402
rect 777 306 823 402
rect -823 70 -777 166
rect -663 70 -617 166
rect -503 70 -457 166
rect -343 70 -297 166
rect -183 70 -137 166
rect -23 70 23 166
rect 137 70 183 166
rect 297 70 343 166
rect 457 70 503 166
rect 617 70 663 166
rect 777 70 823 166
rect -823 -166 -777 -70
rect -663 -166 -617 -70
rect -503 -166 -457 -70
rect -343 -166 -297 -70
rect -183 -166 -137 -70
rect -23 -166 23 -70
rect 137 -166 183 -70
rect 297 -166 343 -70
rect 457 -166 503 -70
rect 617 -166 663 -70
rect 777 -166 823 -70
rect -823 -402 -777 -306
rect -663 -402 -617 -306
rect -503 -402 -457 -306
rect -343 -402 -297 -306
rect -183 -402 -137 -306
rect -23 -402 23 -306
rect 137 -402 183 -306
rect 297 -402 343 -306
rect 457 -402 503 -306
rect 617 -402 663 -306
rect 777 -402 823 -306
rect -823 -638 -777 -542
rect -663 -638 -617 -542
rect -503 -638 -457 -542
rect -343 -638 -297 -542
rect -183 -638 -137 -542
rect -23 -638 23 -542
rect 137 -638 183 -542
rect 297 -638 343 -542
rect 457 -638 503 -542
rect 617 -638 663 -542
rect 777 -638 823 -542
<< pwell >>
rect -860 -708 860 708
<< nmos >>
rect -748 540 -692 640
rect -588 540 -532 640
rect -428 540 -372 640
rect -268 540 -212 640
rect -108 540 -52 640
rect 52 540 108 640
rect 212 540 268 640
rect 372 540 428 640
rect 532 540 588 640
rect 692 540 748 640
rect -748 304 -692 404
rect -588 304 -532 404
rect -428 304 -372 404
rect -268 304 -212 404
rect -108 304 -52 404
rect 52 304 108 404
rect 212 304 268 404
rect 372 304 428 404
rect 532 304 588 404
rect 692 304 748 404
rect -748 68 -692 168
rect -588 68 -532 168
rect -428 68 -372 168
rect -268 68 -212 168
rect -108 68 -52 168
rect 52 68 108 168
rect 212 68 268 168
rect 372 68 428 168
rect 532 68 588 168
rect 692 68 748 168
rect -748 -168 -692 -68
rect -588 -168 -532 -68
rect -428 -168 -372 -68
rect -268 -168 -212 -68
rect -108 -168 -52 -68
rect 52 -168 108 -68
rect 212 -168 268 -68
rect 372 -168 428 -68
rect 532 -168 588 -68
rect 692 -168 748 -68
rect -748 -404 -692 -304
rect -588 -404 -532 -304
rect -428 -404 -372 -304
rect -268 -404 -212 -304
rect -108 -404 -52 -304
rect 52 -404 108 -304
rect 212 -404 268 -304
rect 372 -404 428 -304
rect 532 -404 588 -304
rect 692 -404 748 -304
rect -748 -640 -692 -540
rect -588 -640 -532 -540
rect -428 -640 -372 -540
rect -268 -640 -212 -540
rect -108 -640 -52 -540
rect 52 -640 108 -540
rect 212 -640 268 -540
rect 372 -640 428 -540
rect 532 -640 588 -540
rect 692 -640 748 -540
<< ndiff >>
rect -836 627 -748 640
rect -836 553 -823 627
rect -777 553 -748 627
rect -836 540 -748 553
rect -692 627 -588 640
rect -692 553 -663 627
rect -617 553 -588 627
rect -692 540 -588 553
rect -532 627 -428 640
rect -532 553 -503 627
rect -457 553 -428 627
rect -532 540 -428 553
rect -372 627 -268 640
rect -372 553 -343 627
rect -297 553 -268 627
rect -372 540 -268 553
rect -212 627 -108 640
rect -212 553 -183 627
rect -137 553 -108 627
rect -212 540 -108 553
rect -52 627 52 640
rect -52 553 -23 627
rect 23 553 52 627
rect -52 540 52 553
rect 108 627 212 640
rect 108 553 137 627
rect 183 553 212 627
rect 108 540 212 553
rect 268 627 372 640
rect 268 553 297 627
rect 343 553 372 627
rect 268 540 372 553
rect 428 627 532 640
rect 428 553 457 627
rect 503 553 532 627
rect 428 540 532 553
rect 588 627 692 640
rect 588 553 617 627
rect 663 553 692 627
rect 588 540 692 553
rect 748 627 836 640
rect 748 553 777 627
rect 823 553 836 627
rect 748 540 836 553
rect -836 391 -748 404
rect -836 317 -823 391
rect -777 317 -748 391
rect -836 304 -748 317
rect -692 391 -588 404
rect -692 317 -663 391
rect -617 317 -588 391
rect -692 304 -588 317
rect -532 391 -428 404
rect -532 317 -503 391
rect -457 317 -428 391
rect -532 304 -428 317
rect -372 391 -268 404
rect -372 317 -343 391
rect -297 317 -268 391
rect -372 304 -268 317
rect -212 391 -108 404
rect -212 317 -183 391
rect -137 317 -108 391
rect -212 304 -108 317
rect -52 391 52 404
rect -52 317 -23 391
rect 23 317 52 391
rect -52 304 52 317
rect 108 391 212 404
rect 108 317 137 391
rect 183 317 212 391
rect 108 304 212 317
rect 268 391 372 404
rect 268 317 297 391
rect 343 317 372 391
rect 268 304 372 317
rect 428 391 532 404
rect 428 317 457 391
rect 503 317 532 391
rect 428 304 532 317
rect 588 391 692 404
rect 588 317 617 391
rect 663 317 692 391
rect 588 304 692 317
rect 748 391 836 404
rect 748 317 777 391
rect 823 317 836 391
rect 748 304 836 317
rect -836 155 -748 168
rect -836 81 -823 155
rect -777 81 -748 155
rect -836 68 -748 81
rect -692 155 -588 168
rect -692 81 -663 155
rect -617 81 -588 155
rect -692 68 -588 81
rect -532 155 -428 168
rect -532 81 -503 155
rect -457 81 -428 155
rect -532 68 -428 81
rect -372 155 -268 168
rect -372 81 -343 155
rect -297 81 -268 155
rect -372 68 -268 81
rect -212 155 -108 168
rect -212 81 -183 155
rect -137 81 -108 155
rect -212 68 -108 81
rect -52 155 52 168
rect -52 81 -23 155
rect 23 81 52 155
rect -52 68 52 81
rect 108 155 212 168
rect 108 81 137 155
rect 183 81 212 155
rect 108 68 212 81
rect 268 155 372 168
rect 268 81 297 155
rect 343 81 372 155
rect 268 68 372 81
rect 428 155 532 168
rect 428 81 457 155
rect 503 81 532 155
rect 428 68 532 81
rect 588 155 692 168
rect 588 81 617 155
rect 663 81 692 155
rect 588 68 692 81
rect 748 155 836 168
rect 748 81 777 155
rect 823 81 836 155
rect 748 68 836 81
rect -836 -81 -748 -68
rect -836 -155 -823 -81
rect -777 -155 -748 -81
rect -836 -168 -748 -155
rect -692 -81 -588 -68
rect -692 -155 -663 -81
rect -617 -155 -588 -81
rect -692 -168 -588 -155
rect -532 -81 -428 -68
rect -532 -155 -503 -81
rect -457 -155 -428 -81
rect -532 -168 -428 -155
rect -372 -81 -268 -68
rect -372 -155 -343 -81
rect -297 -155 -268 -81
rect -372 -168 -268 -155
rect -212 -81 -108 -68
rect -212 -155 -183 -81
rect -137 -155 -108 -81
rect -212 -168 -108 -155
rect -52 -81 52 -68
rect -52 -155 -23 -81
rect 23 -155 52 -81
rect -52 -168 52 -155
rect 108 -81 212 -68
rect 108 -155 137 -81
rect 183 -155 212 -81
rect 108 -168 212 -155
rect 268 -81 372 -68
rect 268 -155 297 -81
rect 343 -155 372 -81
rect 268 -168 372 -155
rect 428 -81 532 -68
rect 428 -155 457 -81
rect 503 -155 532 -81
rect 428 -168 532 -155
rect 588 -81 692 -68
rect 588 -155 617 -81
rect 663 -155 692 -81
rect 588 -168 692 -155
rect 748 -81 836 -68
rect 748 -155 777 -81
rect 823 -155 836 -81
rect 748 -168 836 -155
rect -836 -317 -748 -304
rect -836 -391 -823 -317
rect -777 -391 -748 -317
rect -836 -404 -748 -391
rect -692 -317 -588 -304
rect -692 -391 -663 -317
rect -617 -391 -588 -317
rect -692 -404 -588 -391
rect -532 -317 -428 -304
rect -532 -391 -503 -317
rect -457 -391 -428 -317
rect -532 -404 -428 -391
rect -372 -317 -268 -304
rect -372 -391 -343 -317
rect -297 -391 -268 -317
rect -372 -404 -268 -391
rect -212 -317 -108 -304
rect -212 -391 -183 -317
rect -137 -391 -108 -317
rect -212 -404 -108 -391
rect -52 -317 52 -304
rect -52 -391 -23 -317
rect 23 -391 52 -317
rect -52 -404 52 -391
rect 108 -317 212 -304
rect 108 -391 137 -317
rect 183 -391 212 -317
rect 108 -404 212 -391
rect 268 -317 372 -304
rect 268 -391 297 -317
rect 343 -391 372 -317
rect 268 -404 372 -391
rect 428 -317 532 -304
rect 428 -391 457 -317
rect 503 -391 532 -317
rect 428 -404 532 -391
rect 588 -317 692 -304
rect 588 -391 617 -317
rect 663 -391 692 -317
rect 588 -404 692 -391
rect 748 -317 836 -304
rect 748 -391 777 -317
rect 823 -391 836 -317
rect 748 -404 836 -391
rect -836 -553 -748 -540
rect -836 -627 -823 -553
rect -777 -627 -748 -553
rect -836 -640 -748 -627
rect -692 -553 -588 -540
rect -692 -627 -663 -553
rect -617 -627 -588 -553
rect -692 -640 -588 -627
rect -532 -553 -428 -540
rect -532 -627 -503 -553
rect -457 -627 -428 -553
rect -532 -640 -428 -627
rect -372 -553 -268 -540
rect -372 -627 -343 -553
rect -297 -627 -268 -553
rect -372 -640 -268 -627
rect -212 -553 -108 -540
rect -212 -627 -183 -553
rect -137 -627 -108 -553
rect -212 -640 -108 -627
rect -52 -553 52 -540
rect -52 -627 -23 -553
rect 23 -627 52 -553
rect -52 -640 52 -627
rect 108 -553 212 -540
rect 108 -627 137 -553
rect 183 -627 212 -553
rect 108 -640 212 -627
rect 268 -553 372 -540
rect 268 -627 297 -553
rect 343 -627 372 -553
rect 268 -640 372 -627
rect 428 -553 532 -540
rect 428 -627 457 -553
rect 503 -627 532 -553
rect 428 -640 532 -627
rect 588 -553 692 -540
rect 588 -627 617 -553
rect 663 -627 692 -553
rect 588 -640 692 -627
rect 748 -553 836 -540
rect 748 -627 777 -553
rect 823 -627 836 -553
rect 748 -640 836 -627
<< ndiffc >>
rect -823 553 -777 627
rect -663 553 -617 627
rect -503 553 -457 627
rect -343 553 -297 627
rect -183 553 -137 627
rect -23 553 23 627
rect 137 553 183 627
rect 297 553 343 627
rect 457 553 503 627
rect 617 553 663 627
rect 777 553 823 627
rect -823 317 -777 391
rect -663 317 -617 391
rect -503 317 -457 391
rect -343 317 -297 391
rect -183 317 -137 391
rect -23 317 23 391
rect 137 317 183 391
rect 297 317 343 391
rect 457 317 503 391
rect 617 317 663 391
rect 777 317 823 391
rect -823 81 -777 155
rect -663 81 -617 155
rect -503 81 -457 155
rect -343 81 -297 155
rect -183 81 -137 155
rect -23 81 23 155
rect 137 81 183 155
rect 297 81 343 155
rect 457 81 503 155
rect 617 81 663 155
rect 777 81 823 155
rect -823 -155 -777 -81
rect -663 -155 -617 -81
rect -503 -155 -457 -81
rect -343 -155 -297 -81
rect -183 -155 -137 -81
rect -23 -155 23 -81
rect 137 -155 183 -81
rect 297 -155 343 -81
rect 457 -155 503 -81
rect 617 -155 663 -81
rect 777 -155 823 -81
rect -823 -391 -777 -317
rect -663 -391 -617 -317
rect -503 -391 -457 -317
rect -343 -391 -297 -317
rect -183 -391 -137 -317
rect -23 -391 23 -317
rect 137 -391 183 -317
rect 297 -391 343 -317
rect 457 -391 503 -317
rect 617 -391 663 -317
rect 777 -391 823 -317
rect -823 -627 -777 -553
rect -663 -627 -617 -553
rect -503 -627 -457 -553
rect -343 -627 -297 -553
rect -183 -627 -137 -553
rect -23 -627 23 -553
rect 137 -627 183 -553
rect 297 -627 343 -553
rect 457 -627 503 -553
rect 617 -627 663 -553
rect 777 -627 823 -553
<< polysilicon >>
rect -748 640 -692 684
rect -588 640 -532 684
rect -428 640 -372 684
rect -268 640 -212 684
rect -108 640 -52 684
rect 52 640 108 684
rect 212 640 268 684
rect 372 640 428 684
rect 532 640 588 684
rect 692 640 748 684
rect -748 496 -692 540
rect -588 496 -532 540
rect -428 496 -372 540
rect -268 496 -212 540
rect -108 496 -52 540
rect 52 496 108 540
rect 212 496 268 540
rect 372 496 428 540
rect 532 496 588 540
rect 692 496 748 540
rect -748 404 -692 448
rect -588 404 -532 448
rect -428 404 -372 448
rect -268 404 -212 448
rect -108 404 -52 448
rect 52 404 108 448
rect 212 404 268 448
rect 372 404 428 448
rect 532 404 588 448
rect 692 404 748 448
rect -748 260 -692 304
rect -588 260 -532 304
rect -428 260 -372 304
rect -268 260 -212 304
rect -108 260 -52 304
rect 52 260 108 304
rect 212 260 268 304
rect 372 260 428 304
rect 532 260 588 304
rect 692 260 748 304
rect -748 168 -692 212
rect -588 168 -532 212
rect -428 168 -372 212
rect -268 168 -212 212
rect -108 168 -52 212
rect 52 168 108 212
rect 212 168 268 212
rect 372 168 428 212
rect 532 168 588 212
rect 692 168 748 212
rect -748 24 -692 68
rect -588 24 -532 68
rect -428 24 -372 68
rect -268 24 -212 68
rect -108 24 -52 68
rect 52 24 108 68
rect 212 24 268 68
rect 372 24 428 68
rect 532 24 588 68
rect 692 24 748 68
rect -748 -68 -692 -24
rect -588 -68 -532 -24
rect -428 -68 -372 -24
rect -268 -68 -212 -24
rect -108 -68 -52 -24
rect 52 -68 108 -24
rect 212 -68 268 -24
rect 372 -68 428 -24
rect 532 -68 588 -24
rect 692 -68 748 -24
rect -748 -212 -692 -168
rect -588 -212 -532 -168
rect -428 -212 -372 -168
rect -268 -212 -212 -168
rect -108 -212 -52 -168
rect 52 -212 108 -168
rect 212 -212 268 -168
rect 372 -212 428 -168
rect 532 -212 588 -168
rect 692 -212 748 -168
rect -748 -304 -692 -260
rect -588 -304 -532 -260
rect -428 -304 -372 -260
rect -268 -304 -212 -260
rect -108 -304 -52 -260
rect 52 -304 108 -260
rect 212 -304 268 -260
rect 372 -304 428 -260
rect 532 -304 588 -260
rect 692 -304 748 -260
rect -748 -448 -692 -404
rect -588 -448 -532 -404
rect -428 -448 -372 -404
rect -268 -448 -212 -404
rect -108 -448 -52 -404
rect 52 -448 108 -404
rect 212 -448 268 -404
rect 372 -448 428 -404
rect 532 -448 588 -404
rect 692 -448 748 -404
rect -748 -540 -692 -496
rect -588 -540 -532 -496
rect -428 -540 -372 -496
rect -268 -540 -212 -496
rect -108 -540 -52 -496
rect 52 -540 108 -496
rect 212 -540 268 -496
rect 372 -540 428 -496
rect 532 -540 588 -496
rect 692 -540 748 -496
rect -748 -684 -692 -640
rect -588 -684 -532 -640
rect -428 -684 -372 -640
rect -268 -684 -212 -640
rect -108 -684 -52 -640
rect 52 -684 108 -640
rect 212 -684 268 -640
rect 372 -684 428 -640
rect 532 -684 588 -640
rect 692 -684 748 -640
<< metal1 >>
rect -823 627 -777 638
rect -823 542 -777 553
rect -663 627 -617 638
rect -663 542 -617 553
rect -503 627 -457 638
rect -503 542 -457 553
rect -343 627 -297 638
rect -343 542 -297 553
rect -183 627 -137 638
rect -183 542 -137 553
rect -23 627 23 638
rect -23 542 23 553
rect 137 627 183 638
rect 137 542 183 553
rect 297 627 343 638
rect 297 542 343 553
rect 457 627 503 638
rect 457 542 503 553
rect 617 627 663 638
rect 617 542 663 553
rect 777 627 823 638
rect 777 542 823 553
rect -823 391 -777 402
rect -823 306 -777 317
rect -663 391 -617 402
rect -663 306 -617 317
rect -503 391 -457 402
rect -503 306 -457 317
rect -343 391 -297 402
rect -343 306 -297 317
rect -183 391 -137 402
rect -183 306 -137 317
rect -23 391 23 402
rect -23 306 23 317
rect 137 391 183 402
rect 137 306 183 317
rect 297 391 343 402
rect 297 306 343 317
rect 457 391 503 402
rect 457 306 503 317
rect 617 391 663 402
rect 617 306 663 317
rect 777 391 823 402
rect 777 306 823 317
rect -823 155 -777 166
rect -823 70 -777 81
rect -663 155 -617 166
rect -663 70 -617 81
rect -503 155 -457 166
rect -503 70 -457 81
rect -343 155 -297 166
rect -343 70 -297 81
rect -183 155 -137 166
rect -183 70 -137 81
rect -23 155 23 166
rect -23 70 23 81
rect 137 155 183 166
rect 137 70 183 81
rect 297 155 343 166
rect 297 70 343 81
rect 457 155 503 166
rect 457 70 503 81
rect 617 155 663 166
rect 617 70 663 81
rect 777 155 823 166
rect 777 70 823 81
rect -823 -81 -777 -70
rect -823 -166 -777 -155
rect -663 -81 -617 -70
rect -663 -166 -617 -155
rect -503 -81 -457 -70
rect -503 -166 -457 -155
rect -343 -81 -297 -70
rect -343 -166 -297 -155
rect -183 -81 -137 -70
rect -183 -166 -137 -155
rect -23 -81 23 -70
rect -23 -166 23 -155
rect 137 -81 183 -70
rect 137 -166 183 -155
rect 297 -81 343 -70
rect 297 -166 343 -155
rect 457 -81 503 -70
rect 457 -166 503 -155
rect 617 -81 663 -70
rect 617 -166 663 -155
rect 777 -81 823 -70
rect 777 -166 823 -155
rect -823 -317 -777 -306
rect -823 -402 -777 -391
rect -663 -317 -617 -306
rect -663 -402 -617 -391
rect -503 -317 -457 -306
rect -503 -402 -457 -391
rect -343 -317 -297 -306
rect -343 -402 -297 -391
rect -183 -317 -137 -306
rect -183 -402 -137 -391
rect -23 -317 23 -306
rect -23 -402 23 -391
rect 137 -317 183 -306
rect 137 -402 183 -391
rect 297 -317 343 -306
rect 297 -402 343 -391
rect 457 -317 503 -306
rect 457 -402 503 -391
rect 617 -317 663 -306
rect 617 -402 663 -391
rect 777 -317 823 -306
rect 777 -402 823 -391
rect -823 -553 -777 -542
rect -823 -638 -777 -627
rect -663 -553 -617 -542
rect -663 -638 -617 -627
rect -503 -553 -457 -542
rect -503 -638 -457 -627
rect -343 -553 -297 -542
rect -343 -638 -297 -627
rect -183 -553 -137 -542
rect -183 -638 -137 -627
rect -23 -553 23 -542
rect -23 -638 23 -627
rect 137 -553 183 -542
rect 137 -638 183 -627
rect 297 -553 343 -542
rect 297 -638 343 -627
rect 457 -553 503 -542
rect 457 -638 503 -627
rect 617 -553 663 -542
rect 617 -638 663 -627
rect 777 -553 823 -542
rect 777 -638 823 -627
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.5 l 0.280 m 6 nf 10 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
