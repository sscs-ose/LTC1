magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1123 1019 1123
<< metal2 >>
rect -19 118 19 123
rect -19 -118 -14 118
rect 14 -118 19 118
rect -19 -123 19 -118
<< via2 >>
rect -14 -118 14 118
<< metal3 >>
rect -19 118 19 123
rect -19 -118 -14 118
rect 14 -118 19 118
rect -19 -123 19 -118
<< end >>
