magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1217 -1316 1217 1316
<< metal1 >>
rect -217 310 217 316
rect -217 284 -211 310
rect -185 284 -145 310
rect -119 284 -79 310
rect -53 284 -13 310
rect 13 284 53 310
rect 79 284 119 310
rect 145 284 185 310
rect 211 284 217 310
rect -217 244 217 284
rect -217 218 -211 244
rect -185 218 -145 244
rect -119 218 -79 244
rect -53 218 -13 244
rect 13 218 53 244
rect 79 218 119 244
rect 145 218 185 244
rect 211 218 217 244
rect -217 178 217 218
rect -217 152 -211 178
rect -185 152 -145 178
rect -119 152 -79 178
rect -53 152 -13 178
rect 13 152 53 178
rect 79 152 119 178
rect 145 152 185 178
rect 211 152 217 178
rect -217 112 217 152
rect -217 86 -211 112
rect -185 86 -145 112
rect -119 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 119 112
rect 145 86 185 112
rect 211 86 217 112
rect -217 46 217 86
rect -217 20 -211 46
rect -185 20 -145 46
rect -119 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 119 46
rect 145 20 185 46
rect 211 20 217 46
rect -217 -20 217 20
rect -217 -46 -211 -20
rect -185 -46 -145 -20
rect -119 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 119 -20
rect 145 -46 185 -20
rect 211 -46 217 -20
rect -217 -86 217 -46
rect -217 -112 -211 -86
rect -185 -112 -145 -86
rect -119 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 119 -86
rect 145 -112 185 -86
rect 211 -112 217 -86
rect -217 -152 217 -112
rect -217 -178 -211 -152
rect -185 -178 -145 -152
rect -119 -178 -79 -152
rect -53 -178 -13 -152
rect 13 -178 53 -152
rect 79 -178 119 -152
rect 145 -178 185 -152
rect 211 -178 217 -152
rect -217 -218 217 -178
rect -217 -244 -211 -218
rect -185 -244 -145 -218
rect -119 -244 -79 -218
rect -53 -244 -13 -218
rect 13 -244 53 -218
rect 79 -244 119 -218
rect 145 -244 185 -218
rect 211 -244 217 -218
rect -217 -284 217 -244
rect -217 -310 -211 -284
rect -185 -310 -145 -284
rect -119 -310 -79 -284
rect -53 -310 -13 -284
rect 13 -310 53 -284
rect 79 -310 119 -284
rect 145 -310 185 -284
rect 211 -310 217 -284
rect -217 -316 217 -310
<< via1 >>
rect -211 284 -185 310
rect -145 284 -119 310
rect -79 284 -53 310
rect -13 284 13 310
rect 53 284 79 310
rect 119 284 145 310
rect 185 284 211 310
rect -211 218 -185 244
rect -145 218 -119 244
rect -79 218 -53 244
rect -13 218 13 244
rect 53 218 79 244
rect 119 218 145 244
rect 185 218 211 244
rect -211 152 -185 178
rect -145 152 -119 178
rect -79 152 -53 178
rect -13 152 13 178
rect 53 152 79 178
rect 119 152 145 178
rect 185 152 211 178
rect -211 86 -185 112
rect -145 86 -119 112
rect -79 86 -53 112
rect -13 86 13 112
rect 53 86 79 112
rect 119 86 145 112
rect 185 86 211 112
rect -211 20 -185 46
rect -145 20 -119 46
rect -79 20 -53 46
rect -13 20 13 46
rect 53 20 79 46
rect 119 20 145 46
rect 185 20 211 46
rect -211 -46 -185 -20
rect -145 -46 -119 -20
rect -79 -46 -53 -20
rect -13 -46 13 -20
rect 53 -46 79 -20
rect 119 -46 145 -20
rect 185 -46 211 -20
rect -211 -112 -185 -86
rect -145 -112 -119 -86
rect -79 -112 -53 -86
rect -13 -112 13 -86
rect 53 -112 79 -86
rect 119 -112 145 -86
rect 185 -112 211 -86
rect -211 -178 -185 -152
rect -145 -178 -119 -152
rect -79 -178 -53 -152
rect -13 -178 13 -152
rect 53 -178 79 -152
rect 119 -178 145 -152
rect 185 -178 211 -152
rect -211 -244 -185 -218
rect -145 -244 -119 -218
rect -79 -244 -53 -218
rect -13 -244 13 -218
rect 53 -244 79 -218
rect 119 -244 145 -218
rect 185 -244 211 -218
rect -211 -310 -185 -284
rect -145 -310 -119 -284
rect -79 -310 -53 -284
rect -13 -310 13 -284
rect 53 -310 79 -284
rect 119 -310 145 -284
rect 185 -310 211 -284
<< metal2 >>
rect -217 310 217 316
rect -217 284 -211 310
rect -185 284 -145 310
rect -119 284 -79 310
rect -53 284 -13 310
rect 13 284 53 310
rect 79 284 119 310
rect 145 284 185 310
rect 211 284 217 310
rect -217 244 217 284
rect -217 218 -211 244
rect -185 218 -145 244
rect -119 218 -79 244
rect -53 218 -13 244
rect 13 218 53 244
rect 79 218 119 244
rect 145 218 185 244
rect 211 218 217 244
rect -217 178 217 218
rect -217 152 -211 178
rect -185 152 -145 178
rect -119 152 -79 178
rect -53 152 -13 178
rect 13 152 53 178
rect 79 152 119 178
rect 145 152 185 178
rect 211 152 217 178
rect -217 112 217 152
rect -217 86 -211 112
rect -185 86 -145 112
rect -119 86 -79 112
rect -53 86 -13 112
rect 13 86 53 112
rect 79 86 119 112
rect 145 86 185 112
rect 211 86 217 112
rect -217 46 217 86
rect -217 20 -211 46
rect -185 20 -145 46
rect -119 20 -79 46
rect -53 20 -13 46
rect 13 20 53 46
rect 79 20 119 46
rect 145 20 185 46
rect 211 20 217 46
rect -217 -20 217 20
rect -217 -46 -211 -20
rect -185 -46 -145 -20
rect -119 -46 -79 -20
rect -53 -46 -13 -20
rect 13 -46 53 -20
rect 79 -46 119 -20
rect 145 -46 185 -20
rect 211 -46 217 -20
rect -217 -86 217 -46
rect -217 -112 -211 -86
rect -185 -112 -145 -86
rect -119 -112 -79 -86
rect -53 -112 -13 -86
rect 13 -112 53 -86
rect 79 -112 119 -86
rect 145 -112 185 -86
rect 211 -112 217 -86
rect -217 -152 217 -112
rect -217 -178 -211 -152
rect -185 -178 -145 -152
rect -119 -178 -79 -152
rect -53 -178 -13 -152
rect 13 -178 53 -152
rect 79 -178 119 -152
rect 145 -178 185 -152
rect 211 -178 217 -152
rect -217 -218 217 -178
rect -217 -244 -211 -218
rect -185 -244 -145 -218
rect -119 -244 -79 -218
rect -53 -244 -13 -218
rect 13 -244 53 -218
rect 79 -244 119 -218
rect 145 -244 185 -218
rect 211 -244 217 -218
rect -217 -284 217 -244
rect -217 -310 -211 -284
rect -185 -310 -145 -284
rect -119 -310 -79 -284
rect -53 -310 -13 -284
rect 13 -310 53 -284
rect 79 -310 119 -284
rect 145 -310 185 -284
rect 211 -310 217 -284
rect -217 -316 217 -310
<< end >>
