magic
tech gf180mcuC
magscale 1 10
timestamp 1714543819
<< nwell >>
rect -54 624 390 757
rect -54 609 -13 624
rect 63 609 390 624
rect -54 578 390 609
rect -54 349 -16 578
<< psubdiff >>
rect -126 10 499 23
rect -126 -40 -89 10
rect -39 -40 36 10
rect 86 -40 161 10
rect 211 -40 286 10
rect 336 -40 411 10
rect 461 -40 499 10
rect -126 -55 499 -40
<< nsubdiff >>
rect -30 687 49 733
rect -30 641 -10 687
rect 36 641 49 687
rect -30 624 49 641
<< psubdiffcont >>
rect -89 -40 -39 10
rect 36 -40 86 10
rect 161 -40 211 10
rect 286 -40 336 10
rect 411 -40 461 10
<< nsubdiffcont >>
rect -10 641 36 687
<< polysilicon >>
rect 142 423 212 436
rect 80 408 212 423
rect 80 342 95 408
rect 152 342 212 408
rect 80 329 212 342
rect 142 302 212 329
<< polycontact >>
rect 95 342 152 408
<< metal1 >>
rect -231 764 589 842
rect -231 23 -149 764
rect -30 687 330 694
rect -30 641 -10 687
rect 36 641 330 687
rect -30 624 330 641
rect 63 618 330 624
rect 63 492 120 618
rect 95 408 163 420
rect -40 342 95 389
rect 152 342 163 408
rect -40 330 163 342
rect 241 244 302 505
rect 66 23 113 158
rect 508 23 589 764
rect -231 10 589 23
rect -231 -40 -89 10
rect -39 -40 36 10
rect 86 -40 161 10
rect 211 -40 286 10
rect 336 -40 411 10
rect 461 -40 589 10
rect -231 -55 589 -40
use nmos_3p3_AQSZEK  nmos_3p3_AQSZEK_0
timestamp 1714126980
transform 1 0 177 0 1 188
box -147 -138 147 138
use pmos_3p3_HBGRPK  pmos_3p3_HBGRPK_0
timestamp 1714126980
transform 1 0 177 0 1 515
box -213 -166 213 166
<< labels >>
flabel metal1 112 662 112 662 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal1 -6 353 -6 353 0 FreeSans 320 0 0 0 IN
port 1 nsew
flabel metal1 273 357 273 357 0 FreeSans 320 0 0 0 OUT
port 2 nsew
flabel metal1 88 84 88 84 0 FreeSans 320 0 0 0 VSS
port 3 nsew
<< end >>
