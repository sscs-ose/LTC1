magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1729 1019 1729
<< metal2 >>
rect -19 724 19 729
rect -19 696 -14 724
rect 14 696 19 724
rect -19 653 19 696
rect -19 625 -14 653
rect 14 625 19 653
rect -19 582 19 625
rect -19 554 -14 582
rect 14 554 19 582
rect -19 511 19 554
rect -19 483 -14 511
rect 14 483 19 511
rect -19 440 19 483
rect -19 412 -14 440
rect 14 412 19 440
rect -19 369 19 412
rect -19 341 -14 369
rect 14 341 19 369
rect -19 298 19 341
rect -19 270 -14 298
rect 14 270 19 298
rect -19 227 19 270
rect -19 199 -14 227
rect 14 199 19 227
rect -19 156 19 199
rect -19 128 -14 156
rect 14 128 19 156
rect -19 85 19 128
rect -19 57 -14 85
rect 14 57 19 85
rect -19 14 19 57
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -57 19 -14
rect -19 -85 -14 -57
rect 14 -85 19 -57
rect -19 -128 19 -85
rect -19 -156 -14 -128
rect 14 -156 19 -128
rect -19 -199 19 -156
rect -19 -227 -14 -199
rect 14 -227 19 -199
rect -19 -270 19 -227
rect -19 -298 -14 -270
rect 14 -298 19 -270
rect -19 -341 19 -298
rect -19 -369 -14 -341
rect 14 -369 19 -341
rect -19 -412 19 -369
rect -19 -440 -14 -412
rect 14 -440 19 -412
rect -19 -483 19 -440
rect -19 -511 -14 -483
rect 14 -511 19 -483
rect -19 -554 19 -511
rect -19 -582 -14 -554
rect 14 -582 19 -554
rect -19 -625 19 -582
rect -19 -653 -14 -625
rect 14 -653 19 -625
rect -19 -696 19 -653
rect -19 -724 -14 -696
rect 14 -724 19 -696
rect -19 -729 19 -724
<< via2 >>
rect -14 696 14 724
rect -14 625 14 653
rect -14 554 14 582
rect -14 483 14 511
rect -14 412 14 440
rect -14 341 14 369
rect -14 270 14 298
rect -14 199 14 227
rect -14 128 14 156
rect -14 57 14 85
rect -14 -14 14 14
rect -14 -85 14 -57
rect -14 -156 14 -128
rect -14 -227 14 -199
rect -14 -298 14 -270
rect -14 -369 14 -341
rect -14 -440 14 -412
rect -14 -511 14 -483
rect -14 -582 14 -554
rect -14 -653 14 -625
rect -14 -724 14 -696
<< metal3 >>
rect -19 724 19 729
rect -19 696 -14 724
rect 14 696 19 724
rect -19 653 19 696
rect -19 625 -14 653
rect 14 625 19 653
rect -19 582 19 625
rect -19 554 -14 582
rect 14 554 19 582
rect -19 511 19 554
rect -19 483 -14 511
rect 14 483 19 511
rect -19 440 19 483
rect -19 412 -14 440
rect 14 412 19 440
rect -19 369 19 412
rect -19 341 -14 369
rect 14 341 19 369
rect -19 298 19 341
rect -19 270 -14 298
rect 14 270 19 298
rect -19 227 19 270
rect -19 199 -14 227
rect 14 199 19 227
rect -19 156 19 199
rect -19 128 -14 156
rect 14 128 19 156
rect -19 85 19 128
rect -19 57 -14 85
rect 14 57 19 85
rect -19 14 19 57
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -57 19 -14
rect -19 -85 -14 -57
rect 14 -85 19 -57
rect -19 -128 19 -85
rect -19 -156 -14 -128
rect 14 -156 19 -128
rect -19 -199 19 -156
rect -19 -227 -14 -199
rect 14 -227 19 -199
rect -19 -270 19 -227
rect -19 -298 -14 -270
rect 14 -298 19 -270
rect -19 -341 19 -298
rect -19 -369 -14 -341
rect 14 -369 19 -341
rect -19 -412 19 -369
rect -19 -440 -14 -412
rect 14 -440 19 -412
rect -19 -483 19 -440
rect -19 -511 -14 -483
rect 14 -511 19 -483
rect -19 -554 19 -511
rect -19 -582 -14 -554
rect 14 -582 19 -554
rect -19 -625 19 -582
rect -19 -653 -14 -625
rect 14 -653 19 -625
rect -19 -696 19 -653
rect -19 -724 -14 -696
rect 14 -724 19 -696
rect -19 -729 19 -724
<< end >>
