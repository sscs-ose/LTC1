magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1081 -1732 1081 1732
<< metal2 >>
rect -81 727 81 732
rect -81 699 -76 727
rect -48 699 -14 727
rect 14 699 48 727
rect 76 699 81 727
rect -81 665 81 699
rect -81 637 -76 665
rect -48 637 -14 665
rect 14 637 48 665
rect 76 637 81 665
rect -81 603 81 637
rect -81 575 -76 603
rect -48 575 -14 603
rect 14 575 48 603
rect 76 575 81 603
rect -81 541 81 575
rect -81 513 -76 541
rect -48 513 -14 541
rect 14 513 48 541
rect 76 513 81 541
rect -81 479 81 513
rect -81 451 -76 479
rect -48 451 -14 479
rect 14 451 48 479
rect 76 451 81 479
rect -81 417 81 451
rect -81 389 -76 417
rect -48 389 -14 417
rect 14 389 48 417
rect 76 389 81 417
rect -81 355 81 389
rect -81 327 -76 355
rect -48 327 -14 355
rect 14 327 48 355
rect 76 327 81 355
rect -81 293 81 327
rect -81 265 -76 293
rect -48 265 -14 293
rect 14 265 48 293
rect 76 265 81 293
rect -81 231 81 265
rect -81 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 81 231
rect -81 169 81 203
rect -81 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 81 169
rect -81 107 81 141
rect -81 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 81 107
rect -81 45 81 79
rect -81 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 81 45
rect -81 -17 81 17
rect -81 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 81 -17
rect -81 -79 81 -45
rect -81 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 81 -79
rect -81 -141 81 -107
rect -81 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 81 -141
rect -81 -203 81 -169
rect -81 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 81 -203
rect -81 -265 81 -231
rect -81 -293 -76 -265
rect -48 -293 -14 -265
rect 14 -293 48 -265
rect 76 -293 81 -265
rect -81 -327 81 -293
rect -81 -355 -76 -327
rect -48 -355 -14 -327
rect 14 -355 48 -327
rect 76 -355 81 -327
rect -81 -389 81 -355
rect -81 -417 -76 -389
rect -48 -417 -14 -389
rect 14 -417 48 -389
rect 76 -417 81 -389
rect -81 -451 81 -417
rect -81 -479 -76 -451
rect -48 -479 -14 -451
rect 14 -479 48 -451
rect 76 -479 81 -451
rect -81 -513 81 -479
rect -81 -541 -76 -513
rect -48 -541 -14 -513
rect 14 -541 48 -513
rect 76 -541 81 -513
rect -81 -575 81 -541
rect -81 -603 -76 -575
rect -48 -603 -14 -575
rect 14 -603 48 -575
rect 76 -603 81 -575
rect -81 -637 81 -603
rect -81 -665 -76 -637
rect -48 -665 -14 -637
rect 14 -665 48 -637
rect 76 -665 81 -637
rect -81 -699 81 -665
rect -81 -727 -76 -699
rect -48 -727 -14 -699
rect 14 -727 48 -699
rect 76 -727 81 -699
rect -81 -732 81 -727
<< via2 >>
rect -76 699 -48 727
rect -14 699 14 727
rect 48 699 76 727
rect -76 637 -48 665
rect -14 637 14 665
rect 48 637 76 665
rect -76 575 -48 603
rect -14 575 14 603
rect 48 575 76 603
rect -76 513 -48 541
rect -14 513 14 541
rect 48 513 76 541
rect -76 451 -48 479
rect -14 451 14 479
rect 48 451 76 479
rect -76 389 -48 417
rect -14 389 14 417
rect 48 389 76 417
rect -76 327 -48 355
rect -14 327 14 355
rect 48 327 76 355
rect -76 265 -48 293
rect -14 265 14 293
rect 48 265 76 293
rect -76 203 -48 231
rect -14 203 14 231
rect 48 203 76 231
rect -76 141 -48 169
rect -14 141 14 169
rect 48 141 76 169
rect -76 79 -48 107
rect -14 79 14 107
rect 48 79 76 107
rect -76 17 -48 45
rect -14 17 14 45
rect 48 17 76 45
rect -76 -45 -48 -17
rect -14 -45 14 -17
rect 48 -45 76 -17
rect -76 -107 -48 -79
rect -14 -107 14 -79
rect 48 -107 76 -79
rect -76 -169 -48 -141
rect -14 -169 14 -141
rect 48 -169 76 -141
rect -76 -231 -48 -203
rect -14 -231 14 -203
rect 48 -231 76 -203
rect -76 -293 -48 -265
rect -14 -293 14 -265
rect 48 -293 76 -265
rect -76 -355 -48 -327
rect -14 -355 14 -327
rect 48 -355 76 -327
rect -76 -417 -48 -389
rect -14 -417 14 -389
rect 48 -417 76 -389
rect -76 -479 -48 -451
rect -14 -479 14 -451
rect 48 -479 76 -451
rect -76 -541 -48 -513
rect -14 -541 14 -513
rect 48 -541 76 -513
rect -76 -603 -48 -575
rect -14 -603 14 -575
rect 48 -603 76 -575
rect -76 -665 -48 -637
rect -14 -665 14 -637
rect 48 -665 76 -637
rect -76 -727 -48 -699
rect -14 -727 14 -699
rect 48 -727 76 -699
<< metal3 >>
rect -81 727 81 732
rect -81 699 -76 727
rect -48 699 -14 727
rect 14 699 48 727
rect 76 699 81 727
rect -81 665 81 699
rect -81 637 -76 665
rect -48 637 -14 665
rect 14 637 48 665
rect 76 637 81 665
rect -81 603 81 637
rect -81 575 -76 603
rect -48 575 -14 603
rect 14 575 48 603
rect 76 575 81 603
rect -81 541 81 575
rect -81 513 -76 541
rect -48 513 -14 541
rect 14 513 48 541
rect 76 513 81 541
rect -81 479 81 513
rect -81 451 -76 479
rect -48 451 -14 479
rect 14 451 48 479
rect 76 451 81 479
rect -81 417 81 451
rect -81 389 -76 417
rect -48 389 -14 417
rect 14 389 48 417
rect 76 389 81 417
rect -81 355 81 389
rect -81 327 -76 355
rect -48 327 -14 355
rect 14 327 48 355
rect 76 327 81 355
rect -81 293 81 327
rect -81 265 -76 293
rect -48 265 -14 293
rect 14 265 48 293
rect 76 265 81 293
rect -81 231 81 265
rect -81 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 81 231
rect -81 169 81 203
rect -81 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 81 169
rect -81 107 81 141
rect -81 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 81 107
rect -81 45 81 79
rect -81 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 81 45
rect -81 -17 81 17
rect -81 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 81 -17
rect -81 -79 81 -45
rect -81 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 81 -79
rect -81 -141 81 -107
rect -81 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 81 -141
rect -81 -203 81 -169
rect -81 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 81 -203
rect -81 -265 81 -231
rect -81 -293 -76 -265
rect -48 -293 -14 -265
rect 14 -293 48 -265
rect 76 -293 81 -265
rect -81 -327 81 -293
rect -81 -355 -76 -327
rect -48 -355 -14 -327
rect 14 -355 48 -327
rect 76 -355 81 -327
rect -81 -389 81 -355
rect -81 -417 -76 -389
rect -48 -417 -14 -389
rect 14 -417 48 -389
rect 76 -417 81 -389
rect -81 -451 81 -417
rect -81 -479 -76 -451
rect -48 -479 -14 -451
rect 14 -479 48 -451
rect 76 -479 81 -451
rect -81 -513 81 -479
rect -81 -541 -76 -513
rect -48 -541 -14 -513
rect 14 -541 48 -513
rect 76 -541 81 -513
rect -81 -575 81 -541
rect -81 -603 -76 -575
rect -48 -603 -14 -575
rect 14 -603 48 -575
rect 76 -603 81 -575
rect -81 -637 81 -603
rect -81 -665 -76 -637
rect -48 -665 -14 -637
rect 14 -665 48 -637
rect 76 -665 81 -637
rect -81 -699 81 -665
rect -81 -727 -76 -699
rect -48 -727 -14 -699
rect 14 -727 48 -699
rect 76 -727 81 -699
rect -81 -732 81 -727
<< end >>
