** sch_path: /home/shahid/GF180Projects/GF_INV/DAC_low_curr/CM_LSB_V1_TB.sch
**.subckt CM_LSB_V1_TB
V2 VDD GND 3.3
.save i(v2)
I0 VDD ITAIL 2.5u
R1 OUT1 net1 2k m=1
R3 OUT2 net1 2k m=1
R4 OUT3 net1 2k m=1
R5 OUT4 net1 2k m=1
V1 net1 GND 3.3
.save i(v1)
R6 OUT5 net1 2k m=1
R2 OUT_6 net1 2k m=1
x1 ITAIL GND OUT1 OUT2 VDD OUT3 OUT4 OUT5 OUT_6 pex_CM_LSB_mod
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_CM_LSB_mod.spice
.option savecurrents
.control
save all
op

tran 10n 3u
plot v(ITAIL) v(OUT3)
write CM_LSB_V1_TB.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
