magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3099 -7873 3099 7873
<< psubdiff >>
rect -1099 5851 1099 5873
rect -1099 5805 -1077 5851
rect -1031 5805 -953 5851
rect -907 5805 -829 5851
rect -783 5805 -705 5851
rect -659 5805 -581 5851
rect -535 5805 -457 5851
rect -411 5805 -333 5851
rect -287 5805 -209 5851
rect -163 5805 -85 5851
rect -39 5805 39 5851
rect 85 5805 163 5851
rect 209 5805 287 5851
rect 333 5805 411 5851
rect 457 5805 535 5851
rect 581 5805 659 5851
rect 705 5805 783 5851
rect 829 5805 907 5851
rect 953 5805 1031 5851
rect 1077 5805 1099 5851
rect -1099 5727 1099 5805
rect -1099 5681 -1077 5727
rect -1031 5681 -953 5727
rect -907 5681 -829 5727
rect -783 5681 -705 5727
rect -659 5681 -581 5727
rect -535 5681 -457 5727
rect -411 5681 -333 5727
rect -287 5681 -209 5727
rect -163 5681 -85 5727
rect -39 5681 39 5727
rect 85 5681 163 5727
rect 209 5681 287 5727
rect 333 5681 411 5727
rect 457 5681 535 5727
rect 581 5681 659 5727
rect 705 5681 783 5727
rect 829 5681 907 5727
rect 953 5681 1031 5727
rect 1077 5681 1099 5727
rect -1099 5603 1099 5681
rect -1099 5557 -1077 5603
rect -1031 5557 -953 5603
rect -907 5557 -829 5603
rect -783 5557 -705 5603
rect -659 5557 -581 5603
rect -535 5557 -457 5603
rect -411 5557 -333 5603
rect -287 5557 -209 5603
rect -163 5557 -85 5603
rect -39 5557 39 5603
rect 85 5557 163 5603
rect 209 5557 287 5603
rect 333 5557 411 5603
rect 457 5557 535 5603
rect 581 5557 659 5603
rect 705 5557 783 5603
rect 829 5557 907 5603
rect 953 5557 1031 5603
rect 1077 5557 1099 5603
rect -1099 5479 1099 5557
rect -1099 5433 -1077 5479
rect -1031 5433 -953 5479
rect -907 5433 -829 5479
rect -783 5433 -705 5479
rect -659 5433 -581 5479
rect -535 5433 -457 5479
rect -411 5433 -333 5479
rect -287 5433 -209 5479
rect -163 5433 -85 5479
rect -39 5433 39 5479
rect 85 5433 163 5479
rect 209 5433 287 5479
rect 333 5433 411 5479
rect 457 5433 535 5479
rect 581 5433 659 5479
rect 705 5433 783 5479
rect 829 5433 907 5479
rect 953 5433 1031 5479
rect 1077 5433 1099 5479
rect -1099 5355 1099 5433
rect -1099 5309 -1077 5355
rect -1031 5309 -953 5355
rect -907 5309 -829 5355
rect -783 5309 -705 5355
rect -659 5309 -581 5355
rect -535 5309 -457 5355
rect -411 5309 -333 5355
rect -287 5309 -209 5355
rect -163 5309 -85 5355
rect -39 5309 39 5355
rect 85 5309 163 5355
rect 209 5309 287 5355
rect 333 5309 411 5355
rect 457 5309 535 5355
rect 581 5309 659 5355
rect 705 5309 783 5355
rect 829 5309 907 5355
rect 953 5309 1031 5355
rect 1077 5309 1099 5355
rect -1099 5231 1099 5309
rect -1099 5185 -1077 5231
rect -1031 5185 -953 5231
rect -907 5185 -829 5231
rect -783 5185 -705 5231
rect -659 5185 -581 5231
rect -535 5185 -457 5231
rect -411 5185 -333 5231
rect -287 5185 -209 5231
rect -163 5185 -85 5231
rect -39 5185 39 5231
rect 85 5185 163 5231
rect 209 5185 287 5231
rect 333 5185 411 5231
rect 457 5185 535 5231
rect 581 5185 659 5231
rect 705 5185 783 5231
rect 829 5185 907 5231
rect 953 5185 1031 5231
rect 1077 5185 1099 5231
rect -1099 5107 1099 5185
rect -1099 5061 -1077 5107
rect -1031 5061 -953 5107
rect -907 5061 -829 5107
rect -783 5061 -705 5107
rect -659 5061 -581 5107
rect -535 5061 -457 5107
rect -411 5061 -333 5107
rect -287 5061 -209 5107
rect -163 5061 -85 5107
rect -39 5061 39 5107
rect 85 5061 163 5107
rect 209 5061 287 5107
rect 333 5061 411 5107
rect 457 5061 535 5107
rect 581 5061 659 5107
rect 705 5061 783 5107
rect 829 5061 907 5107
rect 953 5061 1031 5107
rect 1077 5061 1099 5107
rect -1099 4983 1099 5061
rect -1099 4937 -1077 4983
rect -1031 4937 -953 4983
rect -907 4937 -829 4983
rect -783 4937 -705 4983
rect -659 4937 -581 4983
rect -535 4937 -457 4983
rect -411 4937 -333 4983
rect -287 4937 -209 4983
rect -163 4937 -85 4983
rect -39 4937 39 4983
rect 85 4937 163 4983
rect 209 4937 287 4983
rect 333 4937 411 4983
rect 457 4937 535 4983
rect 581 4937 659 4983
rect 705 4937 783 4983
rect 829 4937 907 4983
rect 953 4937 1031 4983
rect 1077 4937 1099 4983
rect -1099 4859 1099 4937
rect -1099 4813 -1077 4859
rect -1031 4813 -953 4859
rect -907 4813 -829 4859
rect -783 4813 -705 4859
rect -659 4813 -581 4859
rect -535 4813 -457 4859
rect -411 4813 -333 4859
rect -287 4813 -209 4859
rect -163 4813 -85 4859
rect -39 4813 39 4859
rect 85 4813 163 4859
rect 209 4813 287 4859
rect 333 4813 411 4859
rect 457 4813 535 4859
rect 581 4813 659 4859
rect 705 4813 783 4859
rect 829 4813 907 4859
rect 953 4813 1031 4859
rect 1077 4813 1099 4859
rect -1099 4735 1099 4813
rect -1099 4689 -1077 4735
rect -1031 4689 -953 4735
rect -907 4689 -829 4735
rect -783 4689 -705 4735
rect -659 4689 -581 4735
rect -535 4689 -457 4735
rect -411 4689 -333 4735
rect -287 4689 -209 4735
rect -163 4689 -85 4735
rect -39 4689 39 4735
rect 85 4689 163 4735
rect 209 4689 287 4735
rect 333 4689 411 4735
rect 457 4689 535 4735
rect 581 4689 659 4735
rect 705 4689 783 4735
rect 829 4689 907 4735
rect 953 4689 1031 4735
rect 1077 4689 1099 4735
rect -1099 4611 1099 4689
rect -1099 4565 -1077 4611
rect -1031 4565 -953 4611
rect -907 4565 -829 4611
rect -783 4565 -705 4611
rect -659 4565 -581 4611
rect -535 4565 -457 4611
rect -411 4565 -333 4611
rect -287 4565 -209 4611
rect -163 4565 -85 4611
rect -39 4565 39 4611
rect 85 4565 163 4611
rect 209 4565 287 4611
rect 333 4565 411 4611
rect 457 4565 535 4611
rect 581 4565 659 4611
rect 705 4565 783 4611
rect 829 4565 907 4611
rect 953 4565 1031 4611
rect 1077 4565 1099 4611
rect -1099 4487 1099 4565
rect -1099 4441 -1077 4487
rect -1031 4441 -953 4487
rect -907 4441 -829 4487
rect -783 4441 -705 4487
rect -659 4441 -581 4487
rect -535 4441 -457 4487
rect -411 4441 -333 4487
rect -287 4441 -209 4487
rect -163 4441 -85 4487
rect -39 4441 39 4487
rect 85 4441 163 4487
rect 209 4441 287 4487
rect 333 4441 411 4487
rect 457 4441 535 4487
rect 581 4441 659 4487
rect 705 4441 783 4487
rect 829 4441 907 4487
rect 953 4441 1031 4487
rect 1077 4441 1099 4487
rect -1099 4363 1099 4441
rect -1099 4317 -1077 4363
rect -1031 4317 -953 4363
rect -907 4317 -829 4363
rect -783 4317 -705 4363
rect -659 4317 -581 4363
rect -535 4317 -457 4363
rect -411 4317 -333 4363
rect -287 4317 -209 4363
rect -163 4317 -85 4363
rect -39 4317 39 4363
rect 85 4317 163 4363
rect 209 4317 287 4363
rect 333 4317 411 4363
rect 457 4317 535 4363
rect 581 4317 659 4363
rect 705 4317 783 4363
rect 829 4317 907 4363
rect 953 4317 1031 4363
rect 1077 4317 1099 4363
rect -1099 4239 1099 4317
rect -1099 4193 -1077 4239
rect -1031 4193 -953 4239
rect -907 4193 -829 4239
rect -783 4193 -705 4239
rect -659 4193 -581 4239
rect -535 4193 -457 4239
rect -411 4193 -333 4239
rect -287 4193 -209 4239
rect -163 4193 -85 4239
rect -39 4193 39 4239
rect 85 4193 163 4239
rect 209 4193 287 4239
rect 333 4193 411 4239
rect 457 4193 535 4239
rect 581 4193 659 4239
rect 705 4193 783 4239
rect 829 4193 907 4239
rect 953 4193 1031 4239
rect 1077 4193 1099 4239
rect -1099 4115 1099 4193
rect -1099 4069 -1077 4115
rect -1031 4069 -953 4115
rect -907 4069 -829 4115
rect -783 4069 -705 4115
rect -659 4069 -581 4115
rect -535 4069 -457 4115
rect -411 4069 -333 4115
rect -287 4069 -209 4115
rect -163 4069 -85 4115
rect -39 4069 39 4115
rect 85 4069 163 4115
rect 209 4069 287 4115
rect 333 4069 411 4115
rect 457 4069 535 4115
rect 581 4069 659 4115
rect 705 4069 783 4115
rect 829 4069 907 4115
rect 953 4069 1031 4115
rect 1077 4069 1099 4115
rect -1099 3991 1099 4069
rect -1099 3945 -1077 3991
rect -1031 3945 -953 3991
rect -907 3945 -829 3991
rect -783 3945 -705 3991
rect -659 3945 -581 3991
rect -535 3945 -457 3991
rect -411 3945 -333 3991
rect -287 3945 -209 3991
rect -163 3945 -85 3991
rect -39 3945 39 3991
rect 85 3945 163 3991
rect 209 3945 287 3991
rect 333 3945 411 3991
rect 457 3945 535 3991
rect 581 3945 659 3991
rect 705 3945 783 3991
rect 829 3945 907 3991
rect 953 3945 1031 3991
rect 1077 3945 1099 3991
rect -1099 3867 1099 3945
rect -1099 3821 -1077 3867
rect -1031 3821 -953 3867
rect -907 3821 -829 3867
rect -783 3821 -705 3867
rect -659 3821 -581 3867
rect -535 3821 -457 3867
rect -411 3821 -333 3867
rect -287 3821 -209 3867
rect -163 3821 -85 3867
rect -39 3821 39 3867
rect 85 3821 163 3867
rect 209 3821 287 3867
rect 333 3821 411 3867
rect 457 3821 535 3867
rect 581 3821 659 3867
rect 705 3821 783 3867
rect 829 3821 907 3867
rect 953 3821 1031 3867
rect 1077 3821 1099 3867
rect -1099 3743 1099 3821
rect -1099 3697 -1077 3743
rect -1031 3697 -953 3743
rect -907 3697 -829 3743
rect -783 3697 -705 3743
rect -659 3697 -581 3743
rect -535 3697 -457 3743
rect -411 3697 -333 3743
rect -287 3697 -209 3743
rect -163 3697 -85 3743
rect -39 3697 39 3743
rect 85 3697 163 3743
rect 209 3697 287 3743
rect 333 3697 411 3743
rect 457 3697 535 3743
rect 581 3697 659 3743
rect 705 3697 783 3743
rect 829 3697 907 3743
rect 953 3697 1031 3743
rect 1077 3697 1099 3743
rect -1099 3619 1099 3697
rect -1099 3573 -1077 3619
rect -1031 3573 -953 3619
rect -907 3573 -829 3619
rect -783 3573 -705 3619
rect -659 3573 -581 3619
rect -535 3573 -457 3619
rect -411 3573 -333 3619
rect -287 3573 -209 3619
rect -163 3573 -85 3619
rect -39 3573 39 3619
rect 85 3573 163 3619
rect 209 3573 287 3619
rect 333 3573 411 3619
rect 457 3573 535 3619
rect 581 3573 659 3619
rect 705 3573 783 3619
rect 829 3573 907 3619
rect 953 3573 1031 3619
rect 1077 3573 1099 3619
rect -1099 3495 1099 3573
rect -1099 3449 -1077 3495
rect -1031 3449 -953 3495
rect -907 3449 -829 3495
rect -783 3449 -705 3495
rect -659 3449 -581 3495
rect -535 3449 -457 3495
rect -411 3449 -333 3495
rect -287 3449 -209 3495
rect -163 3449 -85 3495
rect -39 3449 39 3495
rect 85 3449 163 3495
rect 209 3449 287 3495
rect 333 3449 411 3495
rect 457 3449 535 3495
rect 581 3449 659 3495
rect 705 3449 783 3495
rect 829 3449 907 3495
rect 953 3449 1031 3495
rect 1077 3449 1099 3495
rect -1099 3371 1099 3449
rect -1099 3325 -1077 3371
rect -1031 3325 -953 3371
rect -907 3325 -829 3371
rect -783 3325 -705 3371
rect -659 3325 -581 3371
rect -535 3325 -457 3371
rect -411 3325 -333 3371
rect -287 3325 -209 3371
rect -163 3325 -85 3371
rect -39 3325 39 3371
rect 85 3325 163 3371
rect 209 3325 287 3371
rect 333 3325 411 3371
rect 457 3325 535 3371
rect 581 3325 659 3371
rect 705 3325 783 3371
rect 829 3325 907 3371
rect 953 3325 1031 3371
rect 1077 3325 1099 3371
rect -1099 3247 1099 3325
rect -1099 3201 -1077 3247
rect -1031 3201 -953 3247
rect -907 3201 -829 3247
rect -783 3201 -705 3247
rect -659 3201 -581 3247
rect -535 3201 -457 3247
rect -411 3201 -333 3247
rect -287 3201 -209 3247
rect -163 3201 -85 3247
rect -39 3201 39 3247
rect 85 3201 163 3247
rect 209 3201 287 3247
rect 333 3201 411 3247
rect 457 3201 535 3247
rect 581 3201 659 3247
rect 705 3201 783 3247
rect 829 3201 907 3247
rect 953 3201 1031 3247
rect 1077 3201 1099 3247
rect -1099 3123 1099 3201
rect -1099 3077 -1077 3123
rect -1031 3077 -953 3123
rect -907 3077 -829 3123
rect -783 3077 -705 3123
rect -659 3077 -581 3123
rect -535 3077 -457 3123
rect -411 3077 -333 3123
rect -287 3077 -209 3123
rect -163 3077 -85 3123
rect -39 3077 39 3123
rect 85 3077 163 3123
rect 209 3077 287 3123
rect 333 3077 411 3123
rect 457 3077 535 3123
rect 581 3077 659 3123
rect 705 3077 783 3123
rect 829 3077 907 3123
rect 953 3077 1031 3123
rect 1077 3077 1099 3123
rect -1099 2999 1099 3077
rect -1099 2953 -1077 2999
rect -1031 2953 -953 2999
rect -907 2953 -829 2999
rect -783 2953 -705 2999
rect -659 2953 -581 2999
rect -535 2953 -457 2999
rect -411 2953 -333 2999
rect -287 2953 -209 2999
rect -163 2953 -85 2999
rect -39 2953 39 2999
rect 85 2953 163 2999
rect 209 2953 287 2999
rect 333 2953 411 2999
rect 457 2953 535 2999
rect 581 2953 659 2999
rect 705 2953 783 2999
rect 829 2953 907 2999
rect 953 2953 1031 2999
rect 1077 2953 1099 2999
rect -1099 2875 1099 2953
rect -1099 2829 -1077 2875
rect -1031 2829 -953 2875
rect -907 2829 -829 2875
rect -783 2829 -705 2875
rect -659 2829 -581 2875
rect -535 2829 -457 2875
rect -411 2829 -333 2875
rect -287 2829 -209 2875
rect -163 2829 -85 2875
rect -39 2829 39 2875
rect 85 2829 163 2875
rect 209 2829 287 2875
rect 333 2829 411 2875
rect 457 2829 535 2875
rect 581 2829 659 2875
rect 705 2829 783 2875
rect 829 2829 907 2875
rect 953 2829 1031 2875
rect 1077 2829 1099 2875
rect -1099 2751 1099 2829
rect -1099 2705 -1077 2751
rect -1031 2705 -953 2751
rect -907 2705 -829 2751
rect -783 2705 -705 2751
rect -659 2705 -581 2751
rect -535 2705 -457 2751
rect -411 2705 -333 2751
rect -287 2705 -209 2751
rect -163 2705 -85 2751
rect -39 2705 39 2751
rect 85 2705 163 2751
rect 209 2705 287 2751
rect 333 2705 411 2751
rect 457 2705 535 2751
rect 581 2705 659 2751
rect 705 2705 783 2751
rect 829 2705 907 2751
rect 953 2705 1031 2751
rect 1077 2705 1099 2751
rect -1099 2627 1099 2705
rect -1099 2581 -1077 2627
rect -1031 2581 -953 2627
rect -907 2581 -829 2627
rect -783 2581 -705 2627
rect -659 2581 -581 2627
rect -535 2581 -457 2627
rect -411 2581 -333 2627
rect -287 2581 -209 2627
rect -163 2581 -85 2627
rect -39 2581 39 2627
rect 85 2581 163 2627
rect 209 2581 287 2627
rect 333 2581 411 2627
rect 457 2581 535 2627
rect 581 2581 659 2627
rect 705 2581 783 2627
rect 829 2581 907 2627
rect 953 2581 1031 2627
rect 1077 2581 1099 2627
rect -1099 2503 1099 2581
rect -1099 2457 -1077 2503
rect -1031 2457 -953 2503
rect -907 2457 -829 2503
rect -783 2457 -705 2503
rect -659 2457 -581 2503
rect -535 2457 -457 2503
rect -411 2457 -333 2503
rect -287 2457 -209 2503
rect -163 2457 -85 2503
rect -39 2457 39 2503
rect 85 2457 163 2503
rect 209 2457 287 2503
rect 333 2457 411 2503
rect 457 2457 535 2503
rect 581 2457 659 2503
rect 705 2457 783 2503
rect 829 2457 907 2503
rect 953 2457 1031 2503
rect 1077 2457 1099 2503
rect -1099 2379 1099 2457
rect -1099 2333 -1077 2379
rect -1031 2333 -953 2379
rect -907 2333 -829 2379
rect -783 2333 -705 2379
rect -659 2333 -581 2379
rect -535 2333 -457 2379
rect -411 2333 -333 2379
rect -287 2333 -209 2379
rect -163 2333 -85 2379
rect -39 2333 39 2379
rect 85 2333 163 2379
rect 209 2333 287 2379
rect 333 2333 411 2379
rect 457 2333 535 2379
rect 581 2333 659 2379
rect 705 2333 783 2379
rect 829 2333 907 2379
rect 953 2333 1031 2379
rect 1077 2333 1099 2379
rect -1099 2255 1099 2333
rect -1099 2209 -1077 2255
rect -1031 2209 -953 2255
rect -907 2209 -829 2255
rect -783 2209 -705 2255
rect -659 2209 -581 2255
rect -535 2209 -457 2255
rect -411 2209 -333 2255
rect -287 2209 -209 2255
rect -163 2209 -85 2255
rect -39 2209 39 2255
rect 85 2209 163 2255
rect 209 2209 287 2255
rect 333 2209 411 2255
rect 457 2209 535 2255
rect 581 2209 659 2255
rect 705 2209 783 2255
rect 829 2209 907 2255
rect 953 2209 1031 2255
rect 1077 2209 1099 2255
rect -1099 2131 1099 2209
rect -1099 2085 -1077 2131
rect -1031 2085 -953 2131
rect -907 2085 -829 2131
rect -783 2085 -705 2131
rect -659 2085 -581 2131
rect -535 2085 -457 2131
rect -411 2085 -333 2131
rect -287 2085 -209 2131
rect -163 2085 -85 2131
rect -39 2085 39 2131
rect 85 2085 163 2131
rect 209 2085 287 2131
rect 333 2085 411 2131
rect 457 2085 535 2131
rect 581 2085 659 2131
rect 705 2085 783 2131
rect 829 2085 907 2131
rect 953 2085 1031 2131
rect 1077 2085 1099 2131
rect -1099 2007 1099 2085
rect -1099 1961 -1077 2007
rect -1031 1961 -953 2007
rect -907 1961 -829 2007
rect -783 1961 -705 2007
rect -659 1961 -581 2007
rect -535 1961 -457 2007
rect -411 1961 -333 2007
rect -287 1961 -209 2007
rect -163 1961 -85 2007
rect -39 1961 39 2007
rect 85 1961 163 2007
rect 209 1961 287 2007
rect 333 1961 411 2007
rect 457 1961 535 2007
rect 581 1961 659 2007
rect 705 1961 783 2007
rect 829 1961 907 2007
rect 953 1961 1031 2007
rect 1077 1961 1099 2007
rect -1099 1883 1099 1961
rect -1099 1837 -1077 1883
rect -1031 1837 -953 1883
rect -907 1837 -829 1883
rect -783 1837 -705 1883
rect -659 1837 -581 1883
rect -535 1837 -457 1883
rect -411 1837 -333 1883
rect -287 1837 -209 1883
rect -163 1837 -85 1883
rect -39 1837 39 1883
rect 85 1837 163 1883
rect 209 1837 287 1883
rect 333 1837 411 1883
rect 457 1837 535 1883
rect 581 1837 659 1883
rect 705 1837 783 1883
rect 829 1837 907 1883
rect 953 1837 1031 1883
rect 1077 1837 1099 1883
rect -1099 1759 1099 1837
rect -1099 1713 -1077 1759
rect -1031 1713 -953 1759
rect -907 1713 -829 1759
rect -783 1713 -705 1759
rect -659 1713 -581 1759
rect -535 1713 -457 1759
rect -411 1713 -333 1759
rect -287 1713 -209 1759
rect -163 1713 -85 1759
rect -39 1713 39 1759
rect 85 1713 163 1759
rect 209 1713 287 1759
rect 333 1713 411 1759
rect 457 1713 535 1759
rect 581 1713 659 1759
rect 705 1713 783 1759
rect 829 1713 907 1759
rect 953 1713 1031 1759
rect 1077 1713 1099 1759
rect -1099 1635 1099 1713
rect -1099 1589 -1077 1635
rect -1031 1589 -953 1635
rect -907 1589 -829 1635
rect -783 1589 -705 1635
rect -659 1589 -581 1635
rect -535 1589 -457 1635
rect -411 1589 -333 1635
rect -287 1589 -209 1635
rect -163 1589 -85 1635
rect -39 1589 39 1635
rect 85 1589 163 1635
rect 209 1589 287 1635
rect 333 1589 411 1635
rect 457 1589 535 1635
rect 581 1589 659 1635
rect 705 1589 783 1635
rect 829 1589 907 1635
rect 953 1589 1031 1635
rect 1077 1589 1099 1635
rect -1099 1511 1099 1589
rect -1099 1465 -1077 1511
rect -1031 1465 -953 1511
rect -907 1465 -829 1511
rect -783 1465 -705 1511
rect -659 1465 -581 1511
rect -535 1465 -457 1511
rect -411 1465 -333 1511
rect -287 1465 -209 1511
rect -163 1465 -85 1511
rect -39 1465 39 1511
rect 85 1465 163 1511
rect 209 1465 287 1511
rect 333 1465 411 1511
rect 457 1465 535 1511
rect 581 1465 659 1511
rect 705 1465 783 1511
rect 829 1465 907 1511
rect 953 1465 1031 1511
rect 1077 1465 1099 1511
rect -1099 1387 1099 1465
rect -1099 1341 -1077 1387
rect -1031 1341 -953 1387
rect -907 1341 -829 1387
rect -783 1341 -705 1387
rect -659 1341 -581 1387
rect -535 1341 -457 1387
rect -411 1341 -333 1387
rect -287 1341 -209 1387
rect -163 1341 -85 1387
rect -39 1341 39 1387
rect 85 1341 163 1387
rect 209 1341 287 1387
rect 333 1341 411 1387
rect 457 1341 535 1387
rect 581 1341 659 1387
rect 705 1341 783 1387
rect 829 1341 907 1387
rect 953 1341 1031 1387
rect 1077 1341 1099 1387
rect -1099 1263 1099 1341
rect -1099 1217 -1077 1263
rect -1031 1217 -953 1263
rect -907 1217 -829 1263
rect -783 1217 -705 1263
rect -659 1217 -581 1263
rect -535 1217 -457 1263
rect -411 1217 -333 1263
rect -287 1217 -209 1263
rect -163 1217 -85 1263
rect -39 1217 39 1263
rect 85 1217 163 1263
rect 209 1217 287 1263
rect 333 1217 411 1263
rect 457 1217 535 1263
rect 581 1217 659 1263
rect 705 1217 783 1263
rect 829 1217 907 1263
rect 953 1217 1031 1263
rect 1077 1217 1099 1263
rect -1099 1139 1099 1217
rect -1099 1093 -1077 1139
rect -1031 1093 -953 1139
rect -907 1093 -829 1139
rect -783 1093 -705 1139
rect -659 1093 -581 1139
rect -535 1093 -457 1139
rect -411 1093 -333 1139
rect -287 1093 -209 1139
rect -163 1093 -85 1139
rect -39 1093 39 1139
rect 85 1093 163 1139
rect 209 1093 287 1139
rect 333 1093 411 1139
rect 457 1093 535 1139
rect 581 1093 659 1139
rect 705 1093 783 1139
rect 829 1093 907 1139
rect 953 1093 1031 1139
rect 1077 1093 1099 1139
rect -1099 1015 1099 1093
rect -1099 969 -1077 1015
rect -1031 969 -953 1015
rect -907 969 -829 1015
rect -783 969 -705 1015
rect -659 969 -581 1015
rect -535 969 -457 1015
rect -411 969 -333 1015
rect -287 969 -209 1015
rect -163 969 -85 1015
rect -39 969 39 1015
rect 85 969 163 1015
rect 209 969 287 1015
rect 333 969 411 1015
rect 457 969 535 1015
rect 581 969 659 1015
rect 705 969 783 1015
rect 829 969 907 1015
rect 953 969 1031 1015
rect 1077 969 1099 1015
rect -1099 891 1099 969
rect -1099 845 -1077 891
rect -1031 845 -953 891
rect -907 845 -829 891
rect -783 845 -705 891
rect -659 845 -581 891
rect -535 845 -457 891
rect -411 845 -333 891
rect -287 845 -209 891
rect -163 845 -85 891
rect -39 845 39 891
rect 85 845 163 891
rect 209 845 287 891
rect 333 845 411 891
rect 457 845 535 891
rect 581 845 659 891
rect 705 845 783 891
rect 829 845 907 891
rect 953 845 1031 891
rect 1077 845 1099 891
rect -1099 767 1099 845
rect -1099 721 -1077 767
rect -1031 721 -953 767
rect -907 721 -829 767
rect -783 721 -705 767
rect -659 721 -581 767
rect -535 721 -457 767
rect -411 721 -333 767
rect -287 721 -209 767
rect -163 721 -85 767
rect -39 721 39 767
rect 85 721 163 767
rect 209 721 287 767
rect 333 721 411 767
rect 457 721 535 767
rect 581 721 659 767
rect 705 721 783 767
rect 829 721 907 767
rect 953 721 1031 767
rect 1077 721 1099 767
rect -1099 643 1099 721
rect -1099 597 -1077 643
rect -1031 597 -953 643
rect -907 597 -829 643
rect -783 597 -705 643
rect -659 597 -581 643
rect -535 597 -457 643
rect -411 597 -333 643
rect -287 597 -209 643
rect -163 597 -85 643
rect -39 597 39 643
rect 85 597 163 643
rect 209 597 287 643
rect 333 597 411 643
rect 457 597 535 643
rect 581 597 659 643
rect 705 597 783 643
rect 829 597 907 643
rect 953 597 1031 643
rect 1077 597 1099 643
rect -1099 519 1099 597
rect -1099 473 -1077 519
rect -1031 473 -953 519
rect -907 473 -829 519
rect -783 473 -705 519
rect -659 473 -581 519
rect -535 473 -457 519
rect -411 473 -333 519
rect -287 473 -209 519
rect -163 473 -85 519
rect -39 473 39 519
rect 85 473 163 519
rect 209 473 287 519
rect 333 473 411 519
rect 457 473 535 519
rect 581 473 659 519
rect 705 473 783 519
rect 829 473 907 519
rect 953 473 1031 519
rect 1077 473 1099 519
rect -1099 395 1099 473
rect -1099 349 -1077 395
rect -1031 349 -953 395
rect -907 349 -829 395
rect -783 349 -705 395
rect -659 349 -581 395
rect -535 349 -457 395
rect -411 349 -333 395
rect -287 349 -209 395
rect -163 349 -85 395
rect -39 349 39 395
rect 85 349 163 395
rect 209 349 287 395
rect 333 349 411 395
rect 457 349 535 395
rect 581 349 659 395
rect 705 349 783 395
rect 829 349 907 395
rect 953 349 1031 395
rect 1077 349 1099 395
rect -1099 271 1099 349
rect -1099 225 -1077 271
rect -1031 225 -953 271
rect -907 225 -829 271
rect -783 225 -705 271
rect -659 225 -581 271
rect -535 225 -457 271
rect -411 225 -333 271
rect -287 225 -209 271
rect -163 225 -85 271
rect -39 225 39 271
rect 85 225 163 271
rect 209 225 287 271
rect 333 225 411 271
rect 457 225 535 271
rect 581 225 659 271
rect 705 225 783 271
rect 829 225 907 271
rect 953 225 1031 271
rect 1077 225 1099 271
rect -1099 147 1099 225
rect -1099 101 -1077 147
rect -1031 101 -953 147
rect -907 101 -829 147
rect -783 101 -705 147
rect -659 101 -581 147
rect -535 101 -457 147
rect -411 101 -333 147
rect -287 101 -209 147
rect -163 101 -85 147
rect -39 101 39 147
rect 85 101 163 147
rect 209 101 287 147
rect 333 101 411 147
rect 457 101 535 147
rect 581 101 659 147
rect 705 101 783 147
rect 829 101 907 147
rect 953 101 1031 147
rect 1077 101 1099 147
rect -1099 23 1099 101
rect -1099 -23 -1077 23
rect -1031 -23 -953 23
rect -907 -23 -829 23
rect -783 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 783 23
rect 829 -23 907 23
rect 953 -23 1031 23
rect 1077 -23 1099 23
rect -1099 -101 1099 -23
rect -1099 -147 -1077 -101
rect -1031 -147 -953 -101
rect -907 -147 -829 -101
rect -783 -147 -705 -101
rect -659 -147 -581 -101
rect -535 -147 -457 -101
rect -411 -147 -333 -101
rect -287 -147 -209 -101
rect -163 -147 -85 -101
rect -39 -147 39 -101
rect 85 -147 163 -101
rect 209 -147 287 -101
rect 333 -147 411 -101
rect 457 -147 535 -101
rect 581 -147 659 -101
rect 705 -147 783 -101
rect 829 -147 907 -101
rect 953 -147 1031 -101
rect 1077 -147 1099 -101
rect -1099 -225 1099 -147
rect -1099 -271 -1077 -225
rect -1031 -271 -953 -225
rect -907 -271 -829 -225
rect -783 -271 -705 -225
rect -659 -271 -581 -225
rect -535 -271 -457 -225
rect -411 -271 -333 -225
rect -287 -271 -209 -225
rect -163 -271 -85 -225
rect -39 -271 39 -225
rect 85 -271 163 -225
rect 209 -271 287 -225
rect 333 -271 411 -225
rect 457 -271 535 -225
rect 581 -271 659 -225
rect 705 -271 783 -225
rect 829 -271 907 -225
rect 953 -271 1031 -225
rect 1077 -271 1099 -225
rect -1099 -349 1099 -271
rect -1099 -395 -1077 -349
rect -1031 -395 -953 -349
rect -907 -395 -829 -349
rect -783 -395 -705 -349
rect -659 -395 -581 -349
rect -535 -395 -457 -349
rect -411 -395 -333 -349
rect -287 -395 -209 -349
rect -163 -395 -85 -349
rect -39 -395 39 -349
rect 85 -395 163 -349
rect 209 -395 287 -349
rect 333 -395 411 -349
rect 457 -395 535 -349
rect 581 -395 659 -349
rect 705 -395 783 -349
rect 829 -395 907 -349
rect 953 -395 1031 -349
rect 1077 -395 1099 -349
rect -1099 -473 1099 -395
rect -1099 -519 -1077 -473
rect -1031 -519 -953 -473
rect -907 -519 -829 -473
rect -783 -519 -705 -473
rect -659 -519 -581 -473
rect -535 -519 -457 -473
rect -411 -519 -333 -473
rect -287 -519 -209 -473
rect -163 -519 -85 -473
rect -39 -519 39 -473
rect 85 -519 163 -473
rect 209 -519 287 -473
rect 333 -519 411 -473
rect 457 -519 535 -473
rect 581 -519 659 -473
rect 705 -519 783 -473
rect 829 -519 907 -473
rect 953 -519 1031 -473
rect 1077 -519 1099 -473
rect -1099 -597 1099 -519
rect -1099 -643 -1077 -597
rect -1031 -643 -953 -597
rect -907 -643 -829 -597
rect -783 -643 -705 -597
rect -659 -643 -581 -597
rect -535 -643 -457 -597
rect -411 -643 -333 -597
rect -287 -643 -209 -597
rect -163 -643 -85 -597
rect -39 -643 39 -597
rect 85 -643 163 -597
rect 209 -643 287 -597
rect 333 -643 411 -597
rect 457 -643 535 -597
rect 581 -643 659 -597
rect 705 -643 783 -597
rect 829 -643 907 -597
rect 953 -643 1031 -597
rect 1077 -643 1099 -597
rect -1099 -721 1099 -643
rect -1099 -767 -1077 -721
rect -1031 -767 -953 -721
rect -907 -767 -829 -721
rect -783 -767 -705 -721
rect -659 -767 -581 -721
rect -535 -767 -457 -721
rect -411 -767 -333 -721
rect -287 -767 -209 -721
rect -163 -767 -85 -721
rect -39 -767 39 -721
rect 85 -767 163 -721
rect 209 -767 287 -721
rect 333 -767 411 -721
rect 457 -767 535 -721
rect 581 -767 659 -721
rect 705 -767 783 -721
rect 829 -767 907 -721
rect 953 -767 1031 -721
rect 1077 -767 1099 -721
rect -1099 -845 1099 -767
rect -1099 -891 -1077 -845
rect -1031 -891 -953 -845
rect -907 -891 -829 -845
rect -783 -891 -705 -845
rect -659 -891 -581 -845
rect -535 -891 -457 -845
rect -411 -891 -333 -845
rect -287 -891 -209 -845
rect -163 -891 -85 -845
rect -39 -891 39 -845
rect 85 -891 163 -845
rect 209 -891 287 -845
rect 333 -891 411 -845
rect 457 -891 535 -845
rect 581 -891 659 -845
rect 705 -891 783 -845
rect 829 -891 907 -845
rect 953 -891 1031 -845
rect 1077 -891 1099 -845
rect -1099 -969 1099 -891
rect -1099 -1015 -1077 -969
rect -1031 -1015 -953 -969
rect -907 -1015 -829 -969
rect -783 -1015 -705 -969
rect -659 -1015 -581 -969
rect -535 -1015 -457 -969
rect -411 -1015 -333 -969
rect -287 -1015 -209 -969
rect -163 -1015 -85 -969
rect -39 -1015 39 -969
rect 85 -1015 163 -969
rect 209 -1015 287 -969
rect 333 -1015 411 -969
rect 457 -1015 535 -969
rect 581 -1015 659 -969
rect 705 -1015 783 -969
rect 829 -1015 907 -969
rect 953 -1015 1031 -969
rect 1077 -1015 1099 -969
rect -1099 -1093 1099 -1015
rect -1099 -1139 -1077 -1093
rect -1031 -1139 -953 -1093
rect -907 -1139 -829 -1093
rect -783 -1139 -705 -1093
rect -659 -1139 -581 -1093
rect -535 -1139 -457 -1093
rect -411 -1139 -333 -1093
rect -287 -1139 -209 -1093
rect -163 -1139 -85 -1093
rect -39 -1139 39 -1093
rect 85 -1139 163 -1093
rect 209 -1139 287 -1093
rect 333 -1139 411 -1093
rect 457 -1139 535 -1093
rect 581 -1139 659 -1093
rect 705 -1139 783 -1093
rect 829 -1139 907 -1093
rect 953 -1139 1031 -1093
rect 1077 -1139 1099 -1093
rect -1099 -1217 1099 -1139
rect -1099 -1263 -1077 -1217
rect -1031 -1263 -953 -1217
rect -907 -1263 -829 -1217
rect -783 -1263 -705 -1217
rect -659 -1263 -581 -1217
rect -535 -1263 -457 -1217
rect -411 -1263 -333 -1217
rect -287 -1263 -209 -1217
rect -163 -1263 -85 -1217
rect -39 -1263 39 -1217
rect 85 -1263 163 -1217
rect 209 -1263 287 -1217
rect 333 -1263 411 -1217
rect 457 -1263 535 -1217
rect 581 -1263 659 -1217
rect 705 -1263 783 -1217
rect 829 -1263 907 -1217
rect 953 -1263 1031 -1217
rect 1077 -1263 1099 -1217
rect -1099 -1341 1099 -1263
rect -1099 -1387 -1077 -1341
rect -1031 -1387 -953 -1341
rect -907 -1387 -829 -1341
rect -783 -1387 -705 -1341
rect -659 -1387 -581 -1341
rect -535 -1387 -457 -1341
rect -411 -1387 -333 -1341
rect -287 -1387 -209 -1341
rect -163 -1387 -85 -1341
rect -39 -1387 39 -1341
rect 85 -1387 163 -1341
rect 209 -1387 287 -1341
rect 333 -1387 411 -1341
rect 457 -1387 535 -1341
rect 581 -1387 659 -1341
rect 705 -1387 783 -1341
rect 829 -1387 907 -1341
rect 953 -1387 1031 -1341
rect 1077 -1387 1099 -1341
rect -1099 -1465 1099 -1387
rect -1099 -1511 -1077 -1465
rect -1031 -1511 -953 -1465
rect -907 -1511 -829 -1465
rect -783 -1511 -705 -1465
rect -659 -1511 -581 -1465
rect -535 -1511 -457 -1465
rect -411 -1511 -333 -1465
rect -287 -1511 -209 -1465
rect -163 -1511 -85 -1465
rect -39 -1511 39 -1465
rect 85 -1511 163 -1465
rect 209 -1511 287 -1465
rect 333 -1511 411 -1465
rect 457 -1511 535 -1465
rect 581 -1511 659 -1465
rect 705 -1511 783 -1465
rect 829 -1511 907 -1465
rect 953 -1511 1031 -1465
rect 1077 -1511 1099 -1465
rect -1099 -1589 1099 -1511
rect -1099 -1635 -1077 -1589
rect -1031 -1635 -953 -1589
rect -907 -1635 -829 -1589
rect -783 -1635 -705 -1589
rect -659 -1635 -581 -1589
rect -535 -1635 -457 -1589
rect -411 -1635 -333 -1589
rect -287 -1635 -209 -1589
rect -163 -1635 -85 -1589
rect -39 -1635 39 -1589
rect 85 -1635 163 -1589
rect 209 -1635 287 -1589
rect 333 -1635 411 -1589
rect 457 -1635 535 -1589
rect 581 -1635 659 -1589
rect 705 -1635 783 -1589
rect 829 -1635 907 -1589
rect 953 -1635 1031 -1589
rect 1077 -1635 1099 -1589
rect -1099 -1713 1099 -1635
rect -1099 -1759 -1077 -1713
rect -1031 -1759 -953 -1713
rect -907 -1759 -829 -1713
rect -783 -1759 -705 -1713
rect -659 -1759 -581 -1713
rect -535 -1759 -457 -1713
rect -411 -1759 -333 -1713
rect -287 -1759 -209 -1713
rect -163 -1759 -85 -1713
rect -39 -1759 39 -1713
rect 85 -1759 163 -1713
rect 209 -1759 287 -1713
rect 333 -1759 411 -1713
rect 457 -1759 535 -1713
rect 581 -1759 659 -1713
rect 705 -1759 783 -1713
rect 829 -1759 907 -1713
rect 953 -1759 1031 -1713
rect 1077 -1759 1099 -1713
rect -1099 -1837 1099 -1759
rect -1099 -1883 -1077 -1837
rect -1031 -1883 -953 -1837
rect -907 -1883 -829 -1837
rect -783 -1883 -705 -1837
rect -659 -1883 -581 -1837
rect -535 -1883 -457 -1837
rect -411 -1883 -333 -1837
rect -287 -1883 -209 -1837
rect -163 -1883 -85 -1837
rect -39 -1883 39 -1837
rect 85 -1883 163 -1837
rect 209 -1883 287 -1837
rect 333 -1883 411 -1837
rect 457 -1883 535 -1837
rect 581 -1883 659 -1837
rect 705 -1883 783 -1837
rect 829 -1883 907 -1837
rect 953 -1883 1031 -1837
rect 1077 -1883 1099 -1837
rect -1099 -1961 1099 -1883
rect -1099 -2007 -1077 -1961
rect -1031 -2007 -953 -1961
rect -907 -2007 -829 -1961
rect -783 -2007 -705 -1961
rect -659 -2007 -581 -1961
rect -535 -2007 -457 -1961
rect -411 -2007 -333 -1961
rect -287 -2007 -209 -1961
rect -163 -2007 -85 -1961
rect -39 -2007 39 -1961
rect 85 -2007 163 -1961
rect 209 -2007 287 -1961
rect 333 -2007 411 -1961
rect 457 -2007 535 -1961
rect 581 -2007 659 -1961
rect 705 -2007 783 -1961
rect 829 -2007 907 -1961
rect 953 -2007 1031 -1961
rect 1077 -2007 1099 -1961
rect -1099 -2085 1099 -2007
rect -1099 -2131 -1077 -2085
rect -1031 -2131 -953 -2085
rect -907 -2131 -829 -2085
rect -783 -2131 -705 -2085
rect -659 -2131 -581 -2085
rect -535 -2131 -457 -2085
rect -411 -2131 -333 -2085
rect -287 -2131 -209 -2085
rect -163 -2131 -85 -2085
rect -39 -2131 39 -2085
rect 85 -2131 163 -2085
rect 209 -2131 287 -2085
rect 333 -2131 411 -2085
rect 457 -2131 535 -2085
rect 581 -2131 659 -2085
rect 705 -2131 783 -2085
rect 829 -2131 907 -2085
rect 953 -2131 1031 -2085
rect 1077 -2131 1099 -2085
rect -1099 -2209 1099 -2131
rect -1099 -2255 -1077 -2209
rect -1031 -2255 -953 -2209
rect -907 -2255 -829 -2209
rect -783 -2255 -705 -2209
rect -659 -2255 -581 -2209
rect -535 -2255 -457 -2209
rect -411 -2255 -333 -2209
rect -287 -2255 -209 -2209
rect -163 -2255 -85 -2209
rect -39 -2255 39 -2209
rect 85 -2255 163 -2209
rect 209 -2255 287 -2209
rect 333 -2255 411 -2209
rect 457 -2255 535 -2209
rect 581 -2255 659 -2209
rect 705 -2255 783 -2209
rect 829 -2255 907 -2209
rect 953 -2255 1031 -2209
rect 1077 -2255 1099 -2209
rect -1099 -2333 1099 -2255
rect -1099 -2379 -1077 -2333
rect -1031 -2379 -953 -2333
rect -907 -2379 -829 -2333
rect -783 -2379 -705 -2333
rect -659 -2379 -581 -2333
rect -535 -2379 -457 -2333
rect -411 -2379 -333 -2333
rect -287 -2379 -209 -2333
rect -163 -2379 -85 -2333
rect -39 -2379 39 -2333
rect 85 -2379 163 -2333
rect 209 -2379 287 -2333
rect 333 -2379 411 -2333
rect 457 -2379 535 -2333
rect 581 -2379 659 -2333
rect 705 -2379 783 -2333
rect 829 -2379 907 -2333
rect 953 -2379 1031 -2333
rect 1077 -2379 1099 -2333
rect -1099 -2457 1099 -2379
rect -1099 -2503 -1077 -2457
rect -1031 -2503 -953 -2457
rect -907 -2503 -829 -2457
rect -783 -2503 -705 -2457
rect -659 -2503 -581 -2457
rect -535 -2503 -457 -2457
rect -411 -2503 -333 -2457
rect -287 -2503 -209 -2457
rect -163 -2503 -85 -2457
rect -39 -2503 39 -2457
rect 85 -2503 163 -2457
rect 209 -2503 287 -2457
rect 333 -2503 411 -2457
rect 457 -2503 535 -2457
rect 581 -2503 659 -2457
rect 705 -2503 783 -2457
rect 829 -2503 907 -2457
rect 953 -2503 1031 -2457
rect 1077 -2503 1099 -2457
rect -1099 -2581 1099 -2503
rect -1099 -2627 -1077 -2581
rect -1031 -2627 -953 -2581
rect -907 -2627 -829 -2581
rect -783 -2627 -705 -2581
rect -659 -2627 -581 -2581
rect -535 -2627 -457 -2581
rect -411 -2627 -333 -2581
rect -287 -2627 -209 -2581
rect -163 -2627 -85 -2581
rect -39 -2627 39 -2581
rect 85 -2627 163 -2581
rect 209 -2627 287 -2581
rect 333 -2627 411 -2581
rect 457 -2627 535 -2581
rect 581 -2627 659 -2581
rect 705 -2627 783 -2581
rect 829 -2627 907 -2581
rect 953 -2627 1031 -2581
rect 1077 -2627 1099 -2581
rect -1099 -2705 1099 -2627
rect -1099 -2751 -1077 -2705
rect -1031 -2751 -953 -2705
rect -907 -2751 -829 -2705
rect -783 -2751 -705 -2705
rect -659 -2751 -581 -2705
rect -535 -2751 -457 -2705
rect -411 -2751 -333 -2705
rect -287 -2751 -209 -2705
rect -163 -2751 -85 -2705
rect -39 -2751 39 -2705
rect 85 -2751 163 -2705
rect 209 -2751 287 -2705
rect 333 -2751 411 -2705
rect 457 -2751 535 -2705
rect 581 -2751 659 -2705
rect 705 -2751 783 -2705
rect 829 -2751 907 -2705
rect 953 -2751 1031 -2705
rect 1077 -2751 1099 -2705
rect -1099 -2829 1099 -2751
rect -1099 -2875 -1077 -2829
rect -1031 -2875 -953 -2829
rect -907 -2875 -829 -2829
rect -783 -2875 -705 -2829
rect -659 -2875 -581 -2829
rect -535 -2875 -457 -2829
rect -411 -2875 -333 -2829
rect -287 -2875 -209 -2829
rect -163 -2875 -85 -2829
rect -39 -2875 39 -2829
rect 85 -2875 163 -2829
rect 209 -2875 287 -2829
rect 333 -2875 411 -2829
rect 457 -2875 535 -2829
rect 581 -2875 659 -2829
rect 705 -2875 783 -2829
rect 829 -2875 907 -2829
rect 953 -2875 1031 -2829
rect 1077 -2875 1099 -2829
rect -1099 -2953 1099 -2875
rect -1099 -2999 -1077 -2953
rect -1031 -2999 -953 -2953
rect -907 -2999 -829 -2953
rect -783 -2999 -705 -2953
rect -659 -2999 -581 -2953
rect -535 -2999 -457 -2953
rect -411 -2999 -333 -2953
rect -287 -2999 -209 -2953
rect -163 -2999 -85 -2953
rect -39 -2999 39 -2953
rect 85 -2999 163 -2953
rect 209 -2999 287 -2953
rect 333 -2999 411 -2953
rect 457 -2999 535 -2953
rect 581 -2999 659 -2953
rect 705 -2999 783 -2953
rect 829 -2999 907 -2953
rect 953 -2999 1031 -2953
rect 1077 -2999 1099 -2953
rect -1099 -3077 1099 -2999
rect -1099 -3123 -1077 -3077
rect -1031 -3123 -953 -3077
rect -907 -3123 -829 -3077
rect -783 -3123 -705 -3077
rect -659 -3123 -581 -3077
rect -535 -3123 -457 -3077
rect -411 -3123 -333 -3077
rect -287 -3123 -209 -3077
rect -163 -3123 -85 -3077
rect -39 -3123 39 -3077
rect 85 -3123 163 -3077
rect 209 -3123 287 -3077
rect 333 -3123 411 -3077
rect 457 -3123 535 -3077
rect 581 -3123 659 -3077
rect 705 -3123 783 -3077
rect 829 -3123 907 -3077
rect 953 -3123 1031 -3077
rect 1077 -3123 1099 -3077
rect -1099 -3201 1099 -3123
rect -1099 -3247 -1077 -3201
rect -1031 -3247 -953 -3201
rect -907 -3247 -829 -3201
rect -783 -3247 -705 -3201
rect -659 -3247 -581 -3201
rect -535 -3247 -457 -3201
rect -411 -3247 -333 -3201
rect -287 -3247 -209 -3201
rect -163 -3247 -85 -3201
rect -39 -3247 39 -3201
rect 85 -3247 163 -3201
rect 209 -3247 287 -3201
rect 333 -3247 411 -3201
rect 457 -3247 535 -3201
rect 581 -3247 659 -3201
rect 705 -3247 783 -3201
rect 829 -3247 907 -3201
rect 953 -3247 1031 -3201
rect 1077 -3247 1099 -3201
rect -1099 -3325 1099 -3247
rect -1099 -3371 -1077 -3325
rect -1031 -3371 -953 -3325
rect -907 -3371 -829 -3325
rect -783 -3371 -705 -3325
rect -659 -3371 -581 -3325
rect -535 -3371 -457 -3325
rect -411 -3371 -333 -3325
rect -287 -3371 -209 -3325
rect -163 -3371 -85 -3325
rect -39 -3371 39 -3325
rect 85 -3371 163 -3325
rect 209 -3371 287 -3325
rect 333 -3371 411 -3325
rect 457 -3371 535 -3325
rect 581 -3371 659 -3325
rect 705 -3371 783 -3325
rect 829 -3371 907 -3325
rect 953 -3371 1031 -3325
rect 1077 -3371 1099 -3325
rect -1099 -3449 1099 -3371
rect -1099 -3495 -1077 -3449
rect -1031 -3495 -953 -3449
rect -907 -3495 -829 -3449
rect -783 -3495 -705 -3449
rect -659 -3495 -581 -3449
rect -535 -3495 -457 -3449
rect -411 -3495 -333 -3449
rect -287 -3495 -209 -3449
rect -163 -3495 -85 -3449
rect -39 -3495 39 -3449
rect 85 -3495 163 -3449
rect 209 -3495 287 -3449
rect 333 -3495 411 -3449
rect 457 -3495 535 -3449
rect 581 -3495 659 -3449
rect 705 -3495 783 -3449
rect 829 -3495 907 -3449
rect 953 -3495 1031 -3449
rect 1077 -3495 1099 -3449
rect -1099 -3573 1099 -3495
rect -1099 -3619 -1077 -3573
rect -1031 -3619 -953 -3573
rect -907 -3619 -829 -3573
rect -783 -3619 -705 -3573
rect -659 -3619 -581 -3573
rect -535 -3619 -457 -3573
rect -411 -3619 -333 -3573
rect -287 -3619 -209 -3573
rect -163 -3619 -85 -3573
rect -39 -3619 39 -3573
rect 85 -3619 163 -3573
rect 209 -3619 287 -3573
rect 333 -3619 411 -3573
rect 457 -3619 535 -3573
rect 581 -3619 659 -3573
rect 705 -3619 783 -3573
rect 829 -3619 907 -3573
rect 953 -3619 1031 -3573
rect 1077 -3619 1099 -3573
rect -1099 -3697 1099 -3619
rect -1099 -3743 -1077 -3697
rect -1031 -3743 -953 -3697
rect -907 -3743 -829 -3697
rect -783 -3743 -705 -3697
rect -659 -3743 -581 -3697
rect -535 -3743 -457 -3697
rect -411 -3743 -333 -3697
rect -287 -3743 -209 -3697
rect -163 -3743 -85 -3697
rect -39 -3743 39 -3697
rect 85 -3743 163 -3697
rect 209 -3743 287 -3697
rect 333 -3743 411 -3697
rect 457 -3743 535 -3697
rect 581 -3743 659 -3697
rect 705 -3743 783 -3697
rect 829 -3743 907 -3697
rect 953 -3743 1031 -3697
rect 1077 -3743 1099 -3697
rect -1099 -3821 1099 -3743
rect -1099 -3867 -1077 -3821
rect -1031 -3867 -953 -3821
rect -907 -3867 -829 -3821
rect -783 -3867 -705 -3821
rect -659 -3867 -581 -3821
rect -535 -3867 -457 -3821
rect -411 -3867 -333 -3821
rect -287 -3867 -209 -3821
rect -163 -3867 -85 -3821
rect -39 -3867 39 -3821
rect 85 -3867 163 -3821
rect 209 -3867 287 -3821
rect 333 -3867 411 -3821
rect 457 -3867 535 -3821
rect 581 -3867 659 -3821
rect 705 -3867 783 -3821
rect 829 -3867 907 -3821
rect 953 -3867 1031 -3821
rect 1077 -3867 1099 -3821
rect -1099 -3945 1099 -3867
rect -1099 -3991 -1077 -3945
rect -1031 -3991 -953 -3945
rect -907 -3991 -829 -3945
rect -783 -3991 -705 -3945
rect -659 -3991 -581 -3945
rect -535 -3991 -457 -3945
rect -411 -3991 -333 -3945
rect -287 -3991 -209 -3945
rect -163 -3991 -85 -3945
rect -39 -3991 39 -3945
rect 85 -3991 163 -3945
rect 209 -3991 287 -3945
rect 333 -3991 411 -3945
rect 457 -3991 535 -3945
rect 581 -3991 659 -3945
rect 705 -3991 783 -3945
rect 829 -3991 907 -3945
rect 953 -3991 1031 -3945
rect 1077 -3991 1099 -3945
rect -1099 -4069 1099 -3991
rect -1099 -4115 -1077 -4069
rect -1031 -4115 -953 -4069
rect -907 -4115 -829 -4069
rect -783 -4115 -705 -4069
rect -659 -4115 -581 -4069
rect -535 -4115 -457 -4069
rect -411 -4115 -333 -4069
rect -287 -4115 -209 -4069
rect -163 -4115 -85 -4069
rect -39 -4115 39 -4069
rect 85 -4115 163 -4069
rect 209 -4115 287 -4069
rect 333 -4115 411 -4069
rect 457 -4115 535 -4069
rect 581 -4115 659 -4069
rect 705 -4115 783 -4069
rect 829 -4115 907 -4069
rect 953 -4115 1031 -4069
rect 1077 -4115 1099 -4069
rect -1099 -4193 1099 -4115
rect -1099 -4239 -1077 -4193
rect -1031 -4239 -953 -4193
rect -907 -4239 -829 -4193
rect -783 -4239 -705 -4193
rect -659 -4239 -581 -4193
rect -535 -4239 -457 -4193
rect -411 -4239 -333 -4193
rect -287 -4239 -209 -4193
rect -163 -4239 -85 -4193
rect -39 -4239 39 -4193
rect 85 -4239 163 -4193
rect 209 -4239 287 -4193
rect 333 -4239 411 -4193
rect 457 -4239 535 -4193
rect 581 -4239 659 -4193
rect 705 -4239 783 -4193
rect 829 -4239 907 -4193
rect 953 -4239 1031 -4193
rect 1077 -4239 1099 -4193
rect -1099 -4317 1099 -4239
rect -1099 -4363 -1077 -4317
rect -1031 -4363 -953 -4317
rect -907 -4363 -829 -4317
rect -783 -4363 -705 -4317
rect -659 -4363 -581 -4317
rect -535 -4363 -457 -4317
rect -411 -4363 -333 -4317
rect -287 -4363 -209 -4317
rect -163 -4363 -85 -4317
rect -39 -4363 39 -4317
rect 85 -4363 163 -4317
rect 209 -4363 287 -4317
rect 333 -4363 411 -4317
rect 457 -4363 535 -4317
rect 581 -4363 659 -4317
rect 705 -4363 783 -4317
rect 829 -4363 907 -4317
rect 953 -4363 1031 -4317
rect 1077 -4363 1099 -4317
rect -1099 -4441 1099 -4363
rect -1099 -4487 -1077 -4441
rect -1031 -4487 -953 -4441
rect -907 -4487 -829 -4441
rect -783 -4487 -705 -4441
rect -659 -4487 -581 -4441
rect -535 -4487 -457 -4441
rect -411 -4487 -333 -4441
rect -287 -4487 -209 -4441
rect -163 -4487 -85 -4441
rect -39 -4487 39 -4441
rect 85 -4487 163 -4441
rect 209 -4487 287 -4441
rect 333 -4487 411 -4441
rect 457 -4487 535 -4441
rect 581 -4487 659 -4441
rect 705 -4487 783 -4441
rect 829 -4487 907 -4441
rect 953 -4487 1031 -4441
rect 1077 -4487 1099 -4441
rect -1099 -4565 1099 -4487
rect -1099 -4611 -1077 -4565
rect -1031 -4611 -953 -4565
rect -907 -4611 -829 -4565
rect -783 -4611 -705 -4565
rect -659 -4611 -581 -4565
rect -535 -4611 -457 -4565
rect -411 -4611 -333 -4565
rect -287 -4611 -209 -4565
rect -163 -4611 -85 -4565
rect -39 -4611 39 -4565
rect 85 -4611 163 -4565
rect 209 -4611 287 -4565
rect 333 -4611 411 -4565
rect 457 -4611 535 -4565
rect 581 -4611 659 -4565
rect 705 -4611 783 -4565
rect 829 -4611 907 -4565
rect 953 -4611 1031 -4565
rect 1077 -4611 1099 -4565
rect -1099 -4689 1099 -4611
rect -1099 -4735 -1077 -4689
rect -1031 -4735 -953 -4689
rect -907 -4735 -829 -4689
rect -783 -4735 -705 -4689
rect -659 -4735 -581 -4689
rect -535 -4735 -457 -4689
rect -411 -4735 -333 -4689
rect -287 -4735 -209 -4689
rect -163 -4735 -85 -4689
rect -39 -4735 39 -4689
rect 85 -4735 163 -4689
rect 209 -4735 287 -4689
rect 333 -4735 411 -4689
rect 457 -4735 535 -4689
rect 581 -4735 659 -4689
rect 705 -4735 783 -4689
rect 829 -4735 907 -4689
rect 953 -4735 1031 -4689
rect 1077 -4735 1099 -4689
rect -1099 -4813 1099 -4735
rect -1099 -4859 -1077 -4813
rect -1031 -4859 -953 -4813
rect -907 -4859 -829 -4813
rect -783 -4859 -705 -4813
rect -659 -4859 -581 -4813
rect -535 -4859 -457 -4813
rect -411 -4859 -333 -4813
rect -287 -4859 -209 -4813
rect -163 -4859 -85 -4813
rect -39 -4859 39 -4813
rect 85 -4859 163 -4813
rect 209 -4859 287 -4813
rect 333 -4859 411 -4813
rect 457 -4859 535 -4813
rect 581 -4859 659 -4813
rect 705 -4859 783 -4813
rect 829 -4859 907 -4813
rect 953 -4859 1031 -4813
rect 1077 -4859 1099 -4813
rect -1099 -4937 1099 -4859
rect -1099 -4983 -1077 -4937
rect -1031 -4983 -953 -4937
rect -907 -4983 -829 -4937
rect -783 -4983 -705 -4937
rect -659 -4983 -581 -4937
rect -535 -4983 -457 -4937
rect -411 -4983 -333 -4937
rect -287 -4983 -209 -4937
rect -163 -4983 -85 -4937
rect -39 -4983 39 -4937
rect 85 -4983 163 -4937
rect 209 -4983 287 -4937
rect 333 -4983 411 -4937
rect 457 -4983 535 -4937
rect 581 -4983 659 -4937
rect 705 -4983 783 -4937
rect 829 -4983 907 -4937
rect 953 -4983 1031 -4937
rect 1077 -4983 1099 -4937
rect -1099 -5061 1099 -4983
rect -1099 -5107 -1077 -5061
rect -1031 -5107 -953 -5061
rect -907 -5107 -829 -5061
rect -783 -5107 -705 -5061
rect -659 -5107 -581 -5061
rect -535 -5107 -457 -5061
rect -411 -5107 -333 -5061
rect -287 -5107 -209 -5061
rect -163 -5107 -85 -5061
rect -39 -5107 39 -5061
rect 85 -5107 163 -5061
rect 209 -5107 287 -5061
rect 333 -5107 411 -5061
rect 457 -5107 535 -5061
rect 581 -5107 659 -5061
rect 705 -5107 783 -5061
rect 829 -5107 907 -5061
rect 953 -5107 1031 -5061
rect 1077 -5107 1099 -5061
rect -1099 -5185 1099 -5107
rect -1099 -5231 -1077 -5185
rect -1031 -5231 -953 -5185
rect -907 -5231 -829 -5185
rect -783 -5231 -705 -5185
rect -659 -5231 -581 -5185
rect -535 -5231 -457 -5185
rect -411 -5231 -333 -5185
rect -287 -5231 -209 -5185
rect -163 -5231 -85 -5185
rect -39 -5231 39 -5185
rect 85 -5231 163 -5185
rect 209 -5231 287 -5185
rect 333 -5231 411 -5185
rect 457 -5231 535 -5185
rect 581 -5231 659 -5185
rect 705 -5231 783 -5185
rect 829 -5231 907 -5185
rect 953 -5231 1031 -5185
rect 1077 -5231 1099 -5185
rect -1099 -5309 1099 -5231
rect -1099 -5355 -1077 -5309
rect -1031 -5355 -953 -5309
rect -907 -5355 -829 -5309
rect -783 -5355 -705 -5309
rect -659 -5355 -581 -5309
rect -535 -5355 -457 -5309
rect -411 -5355 -333 -5309
rect -287 -5355 -209 -5309
rect -163 -5355 -85 -5309
rect -39 -5355 39 -5309
rect 85 -5355 163 -5309
rect 209 -5355 287 -5309
rect 333 -5355 411 -5309
rect 457 -5355 535 -5309
rect 581 -5355 659 -5309
rect 705 -5355 783 -5309
rect 829 -5355 907 -5309
rect 953 -5355 1031 -5309
rect 1077 -5355 1099 -5309
rect -1099 -5433 1099 -5355
rect -1099 -5479 -1077 -5433
rect -1031 -5479 -953 -5433
rect -907 -5479 -829 -5433
rect -783 -5479 -705 -5433
rect -659 -5479 -581 -5433
rect -535 -5479 -457 -5433
rect -411 -5479 -333 -5433
rect -287 -5479 -209 -5433
rect -163 -5479 -85 -5433
rect -39 -5479 39 -5433
rect 85 -5479 163 -5433
rect 209 -5479 287 -5433
rect 333 -5479 411 -5433
rect 457 -5479 535 -5433
rect 581 -5479 659 -5433
rect 705 -5479 783 -5433
rect 829 -5479 907 -5433
rect 953 -5479 1031 -5433
rect 1077 -5479 1099 -5433
rect -1099 -5557 1099 -5479
rect -1099 -5603 -1077 -5557
rect -1031 -5603 -953 -5557
rect -907 -5603 -829 -5557
rect -783 -5603 -705 -5557
rect -659 -5603 -581 -5557
rect -535 -5603 -457 -5557
rect -411 -5603 -333 -5557
rect -287 -5603 -209 -5557
rect -163 -5603 -85 -5557
rect -39 -5603 39 -5557
rect 85 -5603 163 -5557
rect 209 -5603 287 -5557
rect 333 -5603 411 -5557
rect 457 -5603 535 -5557
rect 581 -5603 659 -5557
rect 705 -5603 783 -5557
rect 829 -5603 907 -5557
rect 953 -5603 1031 -5557
rect 1077 -5603 1099 -5557
rect -1099 -5681 1099 -5603
rect -1099 -5727 -1077 -5681
rect -1031 -5727 -953 -5681
rect -907 -5727 -829 -5681
rect -783 -5727 -705 -5681
rect -659 -5727 -581 -5681
rect -535 -5727 -457 -5681
rect -411 -5727 -333 -5681
rect -287 -5727 -209 -5681
rect -163 -5727 -85 -5681
rect -39 -5727 39 -5681
rect 85 -5727 163 -5681
rect 209 -5727 287 -5681
rect 333 -5727 411 -5681
rect 457 -5727 535 -5681
rect 581 -5727 659 -5681
rect 705 -5727 783 -5681
rect 829 -5727 907 -5681
rect 953 -5727 1031 -5681
rect 1077 -5727 1099 -5681
rect -1099 -5805 1099 -5727
rect -1099 -5851 -1077 -5805
rect -1031 -5851 -953 -5805
rect -907 -5851 -829 -5805
rect -783 -5851 -705 -5805
rect -659 -5851 -581 -5805
rect -535 -5851 -457 -5805
rect -411 -5851 -333 -5805
rect -287 -5851 -209 -5805
rect -163 -5851 -85 -5805
rect -39 -5851 39 -5805
rect 85 -5851 163 -5805
rect 209 -5851 287 -5805
rect 333 -5851 411 -5805
rect 457 -5851 535 -5805
rect 581 -5851 659 -5805
rect 705 -5851 783 -5805
rect 829 -5851 907 -5805
rect 953 -5851 1031 -5805
rect 1077 -5851 1099 -5805
rect -1099 -5873 1099 -5851
<< psubdiffcont >>
rect -1077 5805 -1031 5851
rect -953 5805 -907 5851
rect -829 5805 -783 5851
rect -705 5805 -659 5851
rect -581 5805 -535 5851
rect -457 5805 -411 5851
rect -333 5805 -287 5851
rect -209 5805 -163 5851
rect -85 5805 -39 5851
rect 39 5805 85 5851
rect 163 5805 209 5851
rect 287 5805 333 5851
rect 411 5805 457 5851
rect 535 5805 581 5851
rect 659 5805 705 5851
rect 783 5805 829 5851
rect 907 5805 953 5851
rect 1031 5805 1077 5851
rect -1077 5681 -1031 5727
rect -953 5681 -907 5727
rect -829 5681 -783 5727
rect -705 5681 -659 5727
rect -581 5681 -535 5727
rect -457 5681 -411 5727
rect -333 5681 -287 5727
rect -209 5681 -163 5727
rect -85 5681 -39 5727
rect 39 5681 85 5727
rect 163 5681 209 5727
rect 287 5681 333 5727
rect 411 5681 457 5727
rect 535 5681 581 5727
rect 659 5681 705 5727
rect 783 5681 829 5727
rect 907 5681 953 5727
rect 1031 5681 1077 5727
rect -1077 5557 -1031 5603
rect -953 5557 -907 5603
rect -829 5557 -783 5603
rect -705 5557 -659 5603
rect -581 5557 -535 5603
rect -457 5557 -411 5603
rect -333 5557 -287 5603
rect -209 5557 -163 5603
rect -85 5557 -39 5603
rect 39 5557 85 5603
rect 163 5557 209 5603
rect 287 5557 333 5603
rect 411 5557 457 5603
rect 535 5557 581 5603
rect 659 5557 705 5603
rect 783 5557 829 5603
rect 907 5557 953 5603
rect 1031 5557 1077 5603
rect -1077 5433 -1031 5479
rect -953 5433 -907 5479
rect -829 5433 -783 5479
rect -705 5433 -659 5479
rect -581 5433 -535 5479
rect -457 5433 -411 5479
rect -333 5433 -287 5479
rect -209 5433 -163 5479
rect -85 5433 -39 5479
rect 39 5433 85 5479
rect 163 5433 209 5479
rect 287 5433 333 5479
rect 411 5433 457 5479
rect 535 5433 581 5479
rect 659 5433 705 5479
rect 783 5433 829 5479
rect 907 5433 953 5479
rect 1031 5433 1077 5479
rect -1077 5309 -1031 5355
rect -953 5309 -907 5355
rect -829 5309 -783 5355
rect -705 5309 -659 5355
rect -581 5309 -535 5355
rect -457 5309 -411 5355
rect -333 5309 -287 5355
rect -209 5309 -163 5355
rect -85 5309 -39 5355
rect 39 5309 85 5355
rect 163 5309 209 5355
rect 287 5309 333 5355
rect 411 5309 457 5355
rect 535 5309 581 5355
rect 659 5309 705 5355
rect 783 5309 829 5355
rect 907 5309 953 5355
rect 1031 5309 1077 5355
rect -1077 5185 -1031 5231
rect -953 5185 -907 5231
rect -829 5185 -783 5231
rect -705 5185 -659 5231
rect -581 5185 -535 5231
rect -457 5185 -411 5231
rect -333 5185 -287 5231
rect -209 5185 -163 5231
rect -85 5185 -39 5231
rect 39 5185 85 5231
rect 163 5185 209 5231
rect 287 5185 333 5231
rect 411 5185 457 5231
rect 535 5185 581 5231
rect 659 5185 705 5231
rect 783 5185 829 5231
rect 907 5185 953 5231
rect 1031 5185 1077 5231
rect -1077 5061 -1031 5107
rect -953 5061 -907 5107
rect -829 5061 -783 5107
rect -705 5061 -659 5107
rect -581 5061 -535 5107
rect -457 5061 -411 5107
rect -333 5061 -287 5107
rect -209 5061 -163 5107
rect -85 5061 -39 5107
rect 39 5061 85 5107
rect 163 5061 209 5107
rect 287 5061 333 5107
rect 411 5061 457 5107
rect 535 5061 581 5107
rect 659 5061 705 5107
rect 783 5061 829 5107
rect 907 5061 953 5107
rect 1031 5061 1077 5107
rect -1077 4937 -1031 4983
rect -953 4937 -907 4983
rect -829 4937 -783 4983
rect -705 4937 -659 4983
rect -581 4937 -535 4983
rect -457 4937 -411 4983
rect -333 4937 -287 4983
rect -209 4937 -163 4983
rect -85 4937 -39 4983
rect 39 4937 85 4983
rect 163 4937 209 4983
rect 287 4937 333 4983
rect 411 4937 457 4983
rect 535 4937 581 4983
rect 659 4937 705 4983
rect 783 4937 829 4983
rect 907 4937 953 4983
rect 1031 4937 1077 4983
rect -1077 4813 -1031 4859
rect -953 4813 -907 4859
rect -829 4813 -783 4859
rect -705 4813 -659 4859
rect -581 4813 -535 4859
rect -457 4813 -411 4859
rect -333 4813 -287 4859
rect -209 4813 -163 4859
rect -85 4813 -39 4859
rect 39 4813 85 4859
rect 163 4813 209 4859
rect 287 4813 333 4859
rect 411 4813 457 4859
rect 535 4813 581 4859
rect 659 4813 705 4859
rect 783 4813 829 4859
rect 907 4813 953 4859
rect 1031 4813 1077 4859
rect -1077 4689 -1031 4735
rect -953 4689 -907 4735
rect -829 4689 -783 4735
rect -705 4689 -659 4735
rect -581 4689 -535 4735
rect -457 4689 -411 4735
rect -333 4689 -287 4735
rect -209 4689 -163 4735
rect -85 4689 -39 4735
rect 39 4689 85 4735
rect 163 4689 209 4735
rect 287 4689 333 4735
rect 411 4689 457 4735
rect 535 4689 581 4735
rect 659 4689 705 4735
rect 783 4689 829 4735
rect 907 4689 953 4735
rect 1031 4689 1077 4735
rect -1077 4565 -1031 4611
rect -953 4565 -907 4611
rect -829 4565 -783 4611
rect -705 4565 -659 4611
rect -581 4565 -535 4611
rect -457 4565 -411 4611
rect -333 4565 -287 4611
rect -209 4565 -163 4611
rect -85 4565 -39 4611
rect 39 4565 85 4611
rect 163 4565 209 4611
rect 287 4565 333 4611
rect 411 4565 457 4611
rect 535 4565 581 4611
rect 659 4565 705 4611
rect 783 4565 829 4611
rect 907 4565 953 4611
rect 1031 4565 1077 4611
rect -1077 4441 -1031 4487
rect -953 4441 -907 4487
rect -829 4441 -783 4487
rect -705 4441 -659 4487
rect -581 4441 -535 4487
rect -457 4441 -411 4487
rect -333 4441 -287 4487
rect -209 4441 -163 4487
rect -85 4441 -39 4487
rect 39 4441 85 4487
rect 163 4441 209 4487
rect 287 4441 333 4487
rect 411 4441 457 4487
rect 535 4441 581 4487
rect 659 4441 705 4487
rect 783 4441 829 4487
rect 907 4441 953 4487
rect 1031 4441 1077 4487
rect -1077 4317 -1031 4363
rect -953 4317 -907 4363
rect -829 4317 -783 4363
rect -705 4317 -659 4363
rect -581 4317 -535 4363
rect -457 4317 -411 4363
rect -333 4317 -287 4363
rect -209 4317 -163 4363
rect -85 4317 -39 4363
rect 39 4317 85 4363
rect 163 4317 209 4363
rect 287 4317 333 4363
rect 411 4317 457 4363
rect 535 4317 581 4363
rect 659 4317 705 4363
rect 783 4317 829 4363
rect 907 4317 953 4363
rect 1031 4317 1077 4363
rect -1077 4193 -1031 4239
rect -953 4193 -907 4239
rect -829 4193 -783 4239
rect -705 4193 -659 4239
rect -581 4193 -535 4239
rect -457 4193 -411 4239
rect -333 4193 -287 4239
rect -209 4193 -163 4239
rect -85 4193 -39 4239
rect 39 4193 85 4239
rect 163 4193 209 4239
rect 287 4193 333 4239
rect 411 4193 457 4239
rect 535 4193 581 4239
rect 659 4193 705 4239
rect 783 4193 829 4239
rect 907 4193 953 4239
rect 1031 4193 1077 4239
rect -1077 4069 -1031 4115
rect -953 4069 -907 4115
rect -829 4069 -783 4115
rect -705 4069 -659 4115
rect -581 4069 -535 4115
rect -457 4069 -411 4115
rect -333 4069 -287 4115
rect -209 4069 -163 4115
rect -85 4069 -39 4115
rect 39 4069 85 4115
rect 163 4069 209 4115
rect 287 4069 333 4115
rect 411 4069 457 4115
rect 535 4069 581 4115
rect 659 4069 705 4115
rect 783 4069 829 4115
rect 907 4069 953 4115
rect 1031 4069 1077 4115
rect -1077 3945 -1031 3991
rect -953 3945 -907 3991
rect -829 3945 -783 3991
rect -705 3945 -659 3991
rect -581 3945 -535 3991
rect -457 3945 -411 3991
rect -333 3945 -287 3991
rect -209 3945 -163 3991
rect -85 3945 -39 3991
rect 39 3945 85 3991
rect 163 3945 209 3991
rect 287 3945 333 3991
rect 411 3945 457 3991
rect 535 3945 581 3991
rect 659 3945 705 3991
rect 783 3945 829 3991
rect 907 3945 953 3991
rect 1031 3945 1077 3991
rect -1077 3821 -1031 3867
rect -953 3821 -907 3867
rect -829 3821 -783 3867
rect -705 3821 -659 3867
rect -581 3821 -535 3867
rect -457 3821 -411 3867
rect -333 3821 -287 3867
rect -209 3821 -163 3867
rect -85 3821 -39 3867
rect 39 3821 85 3867
rect 163 3821 209 3867
rect 287 3821 333 3867
rect 411 3821 457 3867
rect 535 3821 581 3867
rect 659 3821 705 3867
rect 783 3821 829 3867
rect 907 3821 953 3867
rect 1031 3821 1077 3867
rect -1077 3697 -1031 3743
rect -953 3697 -907 3743
rect -829 3697 -783 3743
rect -705 3697 -659 3743
rect -581 3697 -535 3743
rect -457 3697 -411 3743
rect -333 3697 -287 3743
rect -209 3697 -163 3743
rect -85 3697 -39 3743
rect 39 3697 85 3743
rect 163 3697 209 3743
rect 287 3697 333 3743
rect 411 3697 457 3743
rect 535 3697 581 3743
rect 659 3697 705 3743
rect 783 3697 829 3743
rect 907 3697 953 3743
rect 1031 3697 1077 3743
rect -1077 3573 -1031 3619
rect -953 3573 -907 3619
rect -829 3573 -783 3619
rect -705 3573 -659 3619
rect -581 3573 -535 3619
rect -457 3573 -411 3619
rect -333 3573 -287 3619
rect -209 3573 -163 3619
rect -85 3573 -39 3619
rect 39 3573 85 3619
rect 163 3573 209 3619
rect 287 3573 333 3619
rect 411 3573 457 3619
rect 535 3573 581 3619
rect 659 3573 705 3619
rect 783 3573 829 3619
rect 907 3573 953 3619
rect 1031 3573 1077 3619
rect -1077 3449 -1031 3495
rect -953 3449 -907 3495
rect -829 3449 -783 3495
rect -705 3449 -659 3495
rect -581 3449 -535 3495
rect -457 3449 -411 3495
rect -333 3449 -287 3495
rect -209 3449 -163 3495
rect -85 3449 -39 3495
rect 39 3449 85 3495
rect 163 3449 209 3495
rect 287 3449 333 3495
rect 411 3449 457 3495
rect 535 3449 581 3495
rect 659 3449 705 3495
rect 783 3449 829 3495
rect 907 3449 953 3495
rect 1031 3449 1077 3495
rect -1077 3325 -1031 3371
rect -953 3325 -907 3371
rect -829 3325 -783 3371
rect -705 3325 -659 3371
rect -581 3325 -535 3371
rect -457 3325 -411 3371
rect -333 3325 -287 3371
rect -209 3325 -163 3371
rect -85 3325 -39 3371
rect 39 3325 85 3371
rect 163 3325 209 3371
rect 287 3325 333 3371
rect 411 3325 457 3371
rect 535 3325 581 3371
rect 659 3325 705 3371
rect 783 3325 829 3371
rect 907 3325 953 3371
rect 1031 3325 1077 3371
rect -1077 3201 -1031 3247
rect -953 3201 -907 3247
rect -829 3201 -783 3247
rect -705 3201 -659 3247
rect -581 3201 -535 3247
rect -457 3201 -411 3247
rect -333 3201 -287 3247
rect -209 3201 -163 3247
rect -85 3201 -39 3247
rect 39 3201 85 3247
rect 163 3201 209 3247
rect 287 3201 333 3247
rect 411 3201 457 3247
rect 535 3201 581 3247
rect 659 3201 705 3247
rect 783 3201 829 3247
rect 907 3201 953 3247
rect 1031 3201 1077 3247
rect -1077 3077 -1031 3123
rect -953 3077 -907 3123
rect -829 3077 -783 3123
rect -705 3077 -659 3123
rect -581 3077 -535 3123
rect -457 3077 -411 3123
rect -333 3077 -287 3123
rect -209 3077 -163 3123
rect -85 3077 -39 3123
rect 39 3077 85 3123
rect 163 3077 209 3123
rect 287 3077 333 3123
rect 411 3077 457 3123
rect 535 3077 581 3123
rect 659 3077 705 3123
rect 783 3077 829 3123
rect 907 3077 953 3123
rect 1031 3077 1077 3123
rect -1077 2953 -1031 2999
rect -953 2953 -907 2999
rect -829 2953 -783 2999
rect -705 2953 -659 2999
rect -581 2953 -535 2999
rect -457 2953 -411 2999
rect -333 2953 -287 2999
rect -209 2953 -163 2999
rect -85 2953 -39 2999
rect 39 2953 85 2999
rect 163 2953 209 2999
rect 287 2953 333 2999
rect 411 2953 457 2999
rect 535 2953 581 2999
rect 659 2953 705 2999
rect 783 2953 829 2999
rect 907 2953 953 2999
rect 1031 2953 1077 2999
rect -1077 2829 -1031 2875
rect -953 2829 -907 2875
rect -829 2829 -783 2875
rect -705 2829 -659 2875
rect -581 2829 -535 2875
rect -457 2829 -411 2875
rect -333 2829 -287 2875
rect -209 2829 -163 2875
rect -85 2829 -39 2875
rect 39 2829 85 2875
rect 163 2829 209 2875
rect 287 2829 333 2875
rect 411 2829 457 2875
rect 535 2829 581 2875
rect 659 2829 705 2875
rect 783 2829 829 2875
rect 907 2829 953 2875
rect 1031 2829 1077 2875
rect -1077 2705 -1031 2751
rect -953 2705 -907 2751
rect -829 2705 -783 2751
rect -705 2705 -659 2751
rect -581 2705 -535 2751
rect -457 2705 -411 2751
rect -333 2705 -287 2751
rect -209 2705 -163 2751
rect -85 2705 -39 2751
rect 39 2705 85 2751
rect 163 2705 209 2751
rect 287 2705 333 2751
rect 411 2705 457 2751
rect 535 2705 581 2751
rect 659 2705 705 2751
rect 783 2705 829 2751
rect 907 2705 953 2751
rect 1031 2705 1077 2751
rect -1077 2581 -1031 2627
rect -953 2581 -907 2627
rect -829 2581 -783 2627
rect -705 2581 -659 2627
rect -581 2581 -535 2627
rect -457 2581 -411 2627
rect -333 2581 -287 2627
rect -209 2581 -163 2627
rect -85 2581 -39 2627
rect 39 2581 85 2627
rect 163 2581 209 2627
rect 287 2581 333 2627
rect 411 2581 457 2627
rect 535 2581 581 2627
rect 659 2581 705 2627
rect 783 2581 829 2627
rect 907 2581 953 2627
rect 1031 2581 1077 2627
rect -1077 2457 -1031 2503
rect -953 2457 -907 2503
rect -829 2457 -783 2503
rect -705 2457 -659 2503
rect -581 2457 -535 2503
rect -457 2457 -411 2503
rect -333 2457 -287 2503
rect -209 2457 -163 2503
rect -85 2457 -39 2503
rect 39 2457 85 2503
rect 163 2457 209 2503
rect 287 2457 333 2503
rect 411 2457 457 2503
rect 535 2457 581 2503
rect 659 2457 705 2503
rect 783 2457 829 2503
rect 907 2457 953 2503
rect 1031 2457 1077 2503
rect -1077 2333 -1031 2379
rect -953 2333 -907 2379
rect -829 2333 -783 2379
rect -705 2333 -659 2379
rect -581 2333 -535 2379
rect -457 2333 -411 2379
rect -333 2333 -287 2379
rect -209 2333 -163 2379
rect -85 2333 -39 2379
rect 39 2333 85 2379
rect 163 2333 209 2379
rect 287 2333 333 2379
rect 411 2333 457 2379
rect 535 2333 581 2379
rect 659 2333 705 2379
rect 783 2333 829 2379
rect 907 2333 953 2379
rect 1031 2333 1077 2379
rect -1077 2209 -1031 2255
rect -953 2209 -907 2255
rect -829 2209 -783 2255
rect -705 2209 -659 2255
rect -581 2209 -535 2255
rect -457 2209 -411 2255
rect -333 2209 -287 2255
rect -209 2209 -163 2255
rect -85 2209 -39 2255
rect 39 2209 85 2255
rect 163 2209 209 2255
rect 287 2209 333 2255
rect 411 2209 457 2255
rect 535 2209 581 2255
rect 659 2209 705 2255
rect 783 2209 829 2255
rect 907 2209 953 2255
rect 1031 2209 1077 2255
rect -1077 2085 -1031 2131
rect -953 2085 -907 2131
rect -829 2085 -783 2131
rect -705 2085 -659 2131
rect -581 2085 -535 2131
rect -457 2085 -411 2131
rect -333 2085 -287 2131
rect -209 2085 -163 2131
rect -85 2085 -39 2131
rect 39 2085 85 2131
rect 163 2085 209 2131
rect 287 2085 333 2131
rect 411 2085 457 2131
rect 535 2085 581 2131
rect 659 2085 705 2131
rect 783 2085 829 2131
rect 907 2085 953 2131
rect 1031 2085 1077 2131
rect -1077 1961 -1031 2007
rect -953 1961 -907 2007
rect -829 1961 -783 2007
rect -705 1961 -659 2007
rect -581 1961 -535 2007
rect -457 1961 -411 2007
rect -333 1961 -287 2007
rect -209 1961 -163 2007
rect -85 1961 -39 2007
rect 39 1961 85 2007
rect 163 1961 209 2007
rect 287 1961 333 2007
rect 411 1961 457 2007
rect 535 1961 581 2007
rect 659 1961 705 2007
rect 783 1961 829 2007
rect 907 1961 953 2007
rect 1031 1961 1077 2007
rect -1077 1837 -1031 1883
rect -953 1837 -907 1883
rect -829 1837 -783 1883
rect -705 1837 -659 1883
rect -581 1837 -535 1883
rect -457 1837 -411 1883
rect -333 1837 -287 1883
rect -209 1837 -163 1883
rect -85 1837 -39 1883
rect 39 1837 85 1883
rect 163 1837 209 1883
rect 287 1837 333 1883
rect 411 1837 457 1883
rect 535 1837 581 1883
rect 659 1837 705 1883
rect 783 1837 829 1883
rect 907 1837 953 1883
rect 1031 1837 1077 1883
rect -1077 1713 -1031 1759
rect -953 1713 -907 1759
rect -829 1713 -783 1759
rect -705 1713 -659 1759
rect -581 1713 -535 1759
rect -457 1713 -411 1759
rect -333 1713 -287 1759
rect -209 1713 -163 1759
rect -85 1713 -39 1759
rect 39 1713 85 1759
rect 163 1713 209 1759
rect 287 1713 333 1759
rect 411 1713 457 1759
rect 535 1713 581 1759
rect 659 1713 705 1759
rect 783 1713 829 1759
rect 907 1713 953 1759
rect 1031 1713 1077 1759
rect -1077 1589 -1031 1635
rect -953 1589 -907 1635
rect -829 1589 -783 1635
rect -705 1589 -659 1635
rect -581 1589 -535 1635
rect -457 1589 -411 1635
rect -333 1589 -287 1635
rect -209 1589 -163 1635
rect -85 1589 -39 1635
rect 39 1589 85 1635
rect 163 1589 209 1635
rect 287 1589 333 1635
rect 411 1589 457 1635
rect 535 1589 581 1635
rect 659 1589 705 1635
rect 783 1589 829 1635
rect 907 1589 953 1635
rect 1031 1589 1077 1635
rect -1077 1465 -1031 1511
rect -953 1465 -907 1511
rect -829 1465 -783 1511
rect -705 1465 -659 1511
rect -581 1465 -535 1511
rect -457 1465 -411 1511
rect -333 1465 -287 1511
rect -209 1465 -163 1511
rect -85 1465 -39 1511
rect 39 1465 85 1511
rect 163 1465 209 1511
rect 287 1465 333 1511
rect 411 1465 457 1511
rect 535 1465 581 1511
rect 659 1465 705 1511
rect 783 1465 829 1511
rect 907 1465 953 1511
rect 1031 1465 1077 1511
rect -1077 1341 -1031 1387
rect -953 1341 -907 1387
rect -829 1341 -783 1387
rect -705 1341 -659 1387
rect -581 1341 -535 1387
rect -457 1341 -411 1387
rect -333 1341 -287 1387
rect -209 1341 -163 1387
rect -85 1341 -39 1387
rect 39 1341 85 1387
rect 163 1341 209 1387
rect 287 1341 333 1387
rect 411 1341 457 1387
rect 535 1341 581 1387
rect 659 1341 705 1387
rect 783 1341 829 1387
rect 907 1341 953 1387
rect 1031 1341 1077 1387
rect -1077 1217 -1031 1263
rect -953 1217 -907 1263
rect -829 1217 -783 1263
rect -705 1217 -659 1263
rect -581 1217 -535 1263
rect -457 1217 -411 1263
rect -333 1217 -287 1263
rect -209 1217 -163 1263
rect -85 1217 -39 1263
rect 39 1217 85 1263
rect 163 1217 209 1263
rect 287 1217 333 1263
rect 411 1217 457 1263
rect 535 1217 581 1263
rect 659 1217 705 1263
rect 783 1217 829 1263
rect 907 1217 953 1263
rect 1031 1217 1077 1263
rect -1077 1093 -1031 1139
rect -953 1093 -907 1139
rect -829 1093 -783 1139
rect -705 1093 -659 1139
rect -581 1093 -535 1139
rect -457 1093 -411 1139
rect -333 1093 -287 1139
rect -209 1093 -163 1139
rect -85 1093 -39 1139
rect 39 1093 85 1139
rect 163 1093 209 1139
rect 287 1093 333 1139
rect 411 1093 457 1139
rect 535 1093 581 1139
rect 659 1093 705 1139
rect 783 1093 829 1139
rect 907 1093 953 1139
rect 1031 1093 1077 1139
rect -1077 969 -1031 1015
rect -953 969 -907 1015
rect -829 969 -783 1015
rect -705 969 -659 1015
rect -581 969 -535 1015
rect -457 969 -411 1015
rect -333 969 -287 1015
rect -209 969 -163 1015
rect -85 969 -39 1015
rect 39 969 85 1015
rect 163 969 209 1015
rect 287 969 333 1015
rect 411 969 457 1015
rect 535 969 581 1015
rect 659 969 705 1015
rect 783 969 829 1015
rect 907 969 953 1015
rect 1031 969 1077 1015
rect -1077 845 -1031 891
rect -953 845 -907 891
rect -829 845 -783 891
rect -705 845 -659 891
rect -581 845 -535 891
rect -457 845 -411 891
rect -333 845 -287 891
rect -209 845 -163 891
rect -85 845 -39 891
rect 39 845 85 891
rect 163 845 209 891
rect 287 845 333 891
rect 411 845 457 891
rect 535 845 581 891
rect 659 845 705 891
rect 783 845 829 891
rect 907 845 953 891
rect 1031 845 1077 891
rect -1077 721 -1031 767
rect -953 721 -907 767
rect -829 721 -783 767
rect -705 721 -659 767
rect -581 721 -535 767
rect -457 721 -411 767
rect -333 721 -287 767
rect -209 721 -163 767
rect -85 721 -39 767
rect 39 721 85 767
rect 163 721 209 767
rect 287 721 333 767
rect 411 721 457 767
rect 535 721 581 767
rect 659 721 705 767
rect 783 721 829 767
rect 907 721 953 767
rect 1031 721 1077 767
rect -1077 597 -1031 643
rect -953 597 -907 643
rect -829 597 -783 643
rect -705 597 -659 643
rect -581 597 -535 643
rect -457 597 -411 643
rect -333 597 -287 643
rect -209 597 -163 643
rect -85 597 -39 643
rect 39 597 85 643
rect 163 597 209 643
rect 287 597 333 643
rect 411 597 457 643
rect 535 597 581 643
rect 659 597 705 643
rect 783 597 829 643
rect 907 597 953 643
rect 1031 597 1077 643
rect -1077 473 -1031 519
rect -953 473 -907 519
rect -829 473 -783 519
rect -705 473 -659 519
rect -581 473 -535 519
rect -457 473 -411 519
rect -333 473 -287 519
rect -209 473 -163 519
rect -85 473 -39 519
rect 39 473 85 519
rect 163 473 209 519
rect 287 473 333 519
rect 411 473 457 519
rect 535 473 581 519
rect 659 473 705 519
rect 783 473 829 519
rect 907 473 953 519
rect 1031 473 1077 519
rect -1077 349 -1031 395
rect -953 349 -907 395
rect -829 349 -783 395
rect -705 349 -659 395
rect -581 349 -535 395
rect -457 349 -411 395
rect -333 349 -287 395
rect -209 349 -163 395
rect -85 349 -39 395
rect 39 349 85 395
rect 163 349 209 395
rect 287 349 333 395
rect 411 349 457 395
rect 535 349 581 395
rect 659 349 705 395
rect 783 349 829 395
rect 907 349 953 395
rect 1031 349 1077 395
rect -1077 225 -1031 271
rect -953 225 -907 271
rect -829 225 -783 271
rect -705 225 -659 271
rect -581 225 -535 271
rect -457 225 -411 271
rect -333 225 -287 271
rect -209 225 -163 271
rect -85 225 -39 271
rect 39 225 85 271
rect 163 225 209 271
rect 287 225 333 271
rect 411 225 457 271
rect 535 225 581 271
rect 659 225 705 271
rect 783 225 829 271
rect 907 225 953 271
rect 1031 225 1077 271
rect -1077 101 -1031 147
rect -953 101 -907 147
rect -829 101 -783 147
rect -705 101 -659 147
rect -581 101 -535 147
rect -457 101 -411 147
rect -333 101 -287 147
rect -209 101 -163 147
rect -85 101 -39 147
rect 39 101 85 147
rect 163 101 209 147
rect 287 101 333 147
rect 411 101 457 147
rect 535 101 581 147
rect 659 101 705 147
rect 783 101 829 147
rect 907 101 953 147
rect 1031 101 1077 147
rect -1077 -23 -1031 23
rect -953 -23 -907 23
rect -829 -23 -783 23
rect -705 -23 -659 23
rect -581 -23 -535 23
rect -457 -23 -411 23
rect -333 -23 -287 23
rect -209 -23 -163 23
rect -85 -23 -39 23
rect 39 -23 85 23
rect 163 -23 209 23
rect 287 -23 333 23
rect 411 -23 457 23
rect 535 -23 581 23
rect 659 -23 705 23
rect 783 -23 829 23
rect 907 -23 953 23
rect 1031 -23 1077 23
rect -1077 -147 -1031 -101
rect -953 -147 -907 -101
rect -829 -147 -783 -101
rect -705 -147 -659 -101
rect -581 -147 -535 -101
rect -457 -147 -411 -101
rect -333 -147 -287 -101
rect -209 -147 -163 -101
rect -85 -147 -39 -101
rect 39 -147 85 -101
rect 163 -147 209 -101
rect 287 -147 333 -101
rect 411 -147 457 -101
rect 535 -147 581 -101
rect 659 -147 705 -101
rect 783 -147 829 -101
rect 907 -147 953 -101
rect 1031 -147 1077 -101
rect -1077 -271 -1031 -225
rect -953 -271 -907 -225
rect -829 -271 -783 -225
rect -705 -271 -659 -225
rect -581 -271 -535 -225
rect -457 -271 -411 -225
rect -333 -271 -287 -225
rect -209 -271 -163 -225
rect -85 -271 -39 -225
rect 39 -271 85 -225
rect 163 -271 209 -225
rect 287 -271 333 -225
rect 411 -271 457 -225
rect 535 -271 581 -225
rect 659 -271 705 -225
rect 783 -271 829 -225
rect 907 -271 953 -225
rect 1031 -271 1077 -225
rect -1077 -395 -1031 -349
rect -953 -395 -907 -349
rect -829 -395 -783 -349
rect -705 -395 -659 -349
rect -581 -395 -535 -349
rect -457 -395 -411 -349
rect -333 -395 -287 -349
rect -209 -395 -163 -349
rect -85 -395 -39 -349
rect 39 -395 85 -349
rect 163 -395 209 -349
rect 287 -395 333 -349
rect 411 -395 457 -349
rect 535 -395 581 -349
rect 659 -395 705 -349
rect 783 -395 829 -349
rect 907 -395 953 -349
rect 1031 -395 1077 -349
rect -1077 -519 -1031 -473
rect -953 -519 -907 -473
rect -829 -519 -783 -473
rect -705 -519 -659 -473
rect -581 -519 -535 -473
rect -457 -519 -411 -473
rect -333 -519 -287 -473
rect -209 -519 -163 -473
rect -85 -519 -39 -473
rect 39 -519 85 -473
rect 163 -519 209 -473
rect 287 -519 333 -473
rect 411 -519 457 -473
rect 535 -519 581 -473
rect 659 -519 705 -473
rect 783 -519 829 -473
rect 907 -519 953 -473
rect 1031 -519 1077 -473
rect -1077 -643 -1031 -597
rect -953 -643 -907 -597
rect -829 -643 -783 -597
rect -705 -643 -659 -597
rect -581 -643 -535 -597
rect -457 -643 -411 -597
rect -333 -643 -287 -597
rect -209 -643 -163 -597
rect -85 -643 -39 -597
rect 39 -643 85 -597
rect 163 -643 209 -597
rect 287 -643 333 -597
rect 411 -643 457 -597
rect 535 -643 581 -597
rect 659 -643 705 -597
rect 783 -643 829 -597
rect 907 -643 953 -597
rect 1031 -643 1077 -597
rect -1077 -767 -1031 -721
rect -953 -767 -907 -721
rect -829 -767 -783 -721
rect -705 -767 -659 -721
rect -581 -767 -535 -721
rect -457 -767 -411 -721
rect -333 -767 -287 -721
rect -209 -767 -163 -721
rect -85 -767 -39 -721
rect 39 -767 85 -721
rect 163 -767 209 -721
rect 287 -767 333 -721
rect 411 -767 457 -721
rect 535 -767 581 -721
rect 659 -767 705 -721
rect 783 -767 829 -721
rect 907 -767 953 -721
rect 1031 -767 1077 -721
rect -1077 -891 -1031 -845
rect -953 -891 -907 -845
rect -829 -891 -783 -845
rect -705 -891 -659 -845
rect -581 -891 -535 -845
rect -457 -891 -411 -845
rect -333 -891 -287 -845
rect -209 -891 -163 -845
rect -85 -891 -39 -845
rect 39 -891 85 -845
rect 163 -891 209 -845
rect 287 -891 333 -845
rect 411 -891 457 -845
rect 535 -891 581 -845
rect 659 -891 705 -845
rect 783 -891 829 -845
rect 907 -891 953 -845
rect 1031 -891 1077 -845
rect -1077 -1015 -1031 -969
rect -953 -1015 -907 -969
rect -829 -1015 -783 -969
rect -705 -1015 -659 -969
rect -581 -1015 -535 -969
rect -457 -1015 -411 -969
rect -333 -1015 -287 -969
rect -209 -1015 -163 -969
rect -85 -1015 -39 -969
rect 39 -1015 85 -969
rect 163 -1015 209 -969
rect 287 -1015 333 -969
rect 411 -1015 457 -969
rect 535 -1015 581 -969
rect 659 -1015 705 -969
rect 783 -1015 829 -969
rect 907 -1015 953 -969
rect 1031 -1015 1077 -969
rect -1077 -1139 -1031 -1093
rect -953 -1139 -907 -1093
rect -829 -1139 -783 -1093
rect -705 -1139 -659 -1093
rect -581 -1139 -535 -1093
rect -457 -1139 -411 -1093
rect -333 -1139 -287 -1093
rect -209 -1139 -163 -1093
rect -85 -1139 -39 -1093
rect 39 -1139 85 -1093
rect 163 -1139 209 -1093
rect 287 -1139 333 -1093
rect 411 -1139 457 -1093
rect 535 -1139 581 -1093
rect 659 -1139 705 -1093
rect 783 -1139 829 -1093
rect 907 -1139 953 -1093
rect 1031 -1139 1077 -1093
rect -1077 -1263 -1031 -1217
rect -953 -1263 -907 -1217
rect -829 -1263 -783 -1217
rect -705 -1263 -659 -1217
rect -581 -1263 -535 -1217
rect -457 -1263 -411 -1217
rect -333 -1263 -287 -1217
rect -209 -1263 -163 -1217
rect -85 -1263 -39 -1217
rect 39 -1263 85 -1217
rect 163 -1263 209 -1217
rect 287 -1263 333 -1217
rect 411 -1263 457 -1217
rect 535 -1263 581 -1217
rect 659 -1263 705 -1217
rect 783 -1263 829 -1217
rect 907 -1263 953 -1217
rect 1031 -1263 1077 -1217
rect -1077 -1387 -1031 -1341
rect -953 -1387 -907 -1341
rect -829 -1387 -783 -1341
rect -705 -1387 -659 -1341
rect -581 -1387 -535 -1341
rect -457 -1387 -411 -1341
rect -333 -1387 -287 -1341
rect -209 -1387 -163 -1341
rect -85 -1387 -39 -1341
rect 39 -1387 85 -1341
rect 163 -1387 209 -1341
rect 287 -1387 333 -1341
rect 411 -1387 457 -1341
rect 535 -1387 581 -1341
rect 659 -1387 705 -1341
rect 783 -1387 829 -1341
rect 907 -1387 953 -1341
rect 1031 -1387 1077 -1341
rect -1077 -1511 -1031 -1465
rect -953 -1511 -907 -1465
rect -829 -1511 -783 -1465
rect -705 -1511 -659 -1465
rect -581 -1511 -535 -1465
rect -457 -1511 -411 -1465
rect -333 -1511 -287 -1465
rect -209 -1511 -163 -1465
rect -85 -1511 -39 -1465
rect 39 -1511 85 -1465
rect 163 -1511 209 -1465
rect 287 -1511 333 -1465
rect 411 -1511 457 -1465
rect 535 -1511 581 -1465
rect 659 -1511 705 -1465
rect 783 -1511 829 -1465
rect 907 -1511 953 -1465
rect 1031 -1511 1077 -1465
rect -1077 -1635 -1031 -1589
rect -953 -1635 -907 -1589
rect -829 -1635 -783 -1589
rect -705 -1635 -659 -1589
rect -581 -1635 -535 -1589
rect -457 -1635 -411 -1589
rect -333 -1635 -287 -1589
rect -209 -1635 -163 -1589
rect -85 -1635 -39 -1589
rect 39 -1635 85 -1589
rect 163 -1635 209 -1589
rect 287 -1635 333 -1589
rect 411 -1635 457 -1589
rect 535 -1635 581 -1589
rect 659 -1635 705 -1589
rect 783 -1635 829 -1589
rect 907 -1635 953 -1589
rect 1031 -1635 1077 -1589
rect -1077 -1759 -1031 -1713
rect -953 -1759 -907 -1713
rect -829 -1759 -783 -1713
rect -705 -1759 -659 -1713
rect -581 -1759 -535 -1713
rect -457 -1759 -411 -1713
rect -333 -1759 -287 -1713
rect -209 -1759 -163 -1713
rect -85 -1759 -39 -1713
rect 39 -1759 85 -1713
rect 163 -1759 209 -1713
rect 287 -1759 333 -1713
rect 411 -1759 457 -1713
rect 535 -1759 581 -1713
rect 659 -1759 705 -1713
rect 783 -1759 829 -1713
rect 907 -1759 953 -1713
rect 1031 -1759 1077 -1713
rect -1077 -1883 -1031 -1837
rect -953 -1883 -907 -1837
rect -829 -1883 -783 -1837
rect -705 -1883 -659 -1837
rect -581 -1883 -535 -1837
rect -457 -1883 -411 -1837
rect -333 -1883 -287 -1837
rect -209 -1883 -163 -1837
rect -85 -1883 -39 -1837
rect 39 -1883 85 -1837
rect 163 -1883 209 -1837
rect 287 -1883 333 -1837
rect 411 -1883 457 -1837
rect 535 -1883 581 -1837
rect 659 -1883 705 -1837
rect 783 -1883 829 -1837
rect 907 -1883 953 -1837
rect 1031 -1883 1077 -1837
rect -1077 -2007 -1031 -1961
rect -953 -2007 -907 -1961
rect -829 -2007 -783 -1961
rect -705 -2007 -659 -1961
rect -581 -2007 -535 -1961
rect -457 -2007 -411 -1961
rect -333 -2007 -287 -1961
rect -209 -2007 -163 -1961
rect -85 -2007 -39 -1961
rect 39 -2007 85 -1961
rect 163 -2007 209 -1961
rect 287 -2007 333 -1961
rect 411 -2007 457 -1961
rect 535 -2007 581 -1961
rect 659 -2007 705 -1961
rect 783 -2007 829 -1961
rect 907 -2007 953 -1961
rect 1031 -2007 1077 -1961
rect -1077 -2131 -1031 -2085
rect -953 -2131 -907 -2085
rect -829 -2131 -783 -2085
rect -705 -2131 -659 -2085
rect -581 -2131 -535 -2085
rect -457 -2131 -411 -2085
rect -333 -2131 -287 -2085
rect -209 -2131 -163 -2085
rect -85 -2131 -39 -2085
rect 39 -2131 85 -2085
rect 163 -2131 209 -2085
rect 287 -2131 333 -2085
rect 411 -2131 457 -2085
rect 535 -2131 581 -2085
rect 659 -2131 705 -2085
rect 783 -2131 829 -2085
rect 907 -2131 953 -2085
rect 1031 -2131 1077 -2085
rect -1077 -2255 -1031 -2209
rect -953 -2255 -907 -2209
rect -829 -2255 -783 -2209
rect -705 -2255 -659 -2209
rect -581 -2255 -535 -2209
rect -457 -2255 -411 -2209
rect -333 -2255 -287 -2209
rect -209 -2255 -163 -2209
rect -85 -2255 -39 -2209
rect 39 -2255 85 -2209
rect 163 -2255 209 -2209
rect 287 -2255 333 -2209
rect 411 -2255 457 -2209
rect 535 -2255 581 -2209
rect 659 -2255 705 -2209
rect 783 -2255 829 -2209
rect 907 -2255 953 -2209
rect 1031 -2255 1077 -2209
rect -1077 -2379 -1031 -2333
rect -953 -2379 -907 -2333
rect -829 -2379 -783 -2333
rect -705 -2379 -659 -2333
rect -581 -2379 -535 -2333
rect -457 -2379 -411 -2333
rect -333 -2379 -287 -2333
rect -209 -2379 -163 -2333
rect -85 -2379 -39 -2333
rect 39 -2379 85 -2333
rect 163 -2379 209 -2333
rect 287 -2379 333 -2333
rect 411 -2379 457 -2333
rect 535 -2379 581 -2333
rect 659 -2379 705 -2333
rect 783 -2379 829 -2333
rect 907 -2379 953 -2333
rect 1031 -2379 1077 -2333
rect -1077 -2503 -1031 -2457
rect -953 -2503 -907 -2457
rect -829 -2503 -783 -2457
rect -705 -2503 -659 -2457
rect -581 -2503 -535 -2457
rect -457 -2503 -411 -2457
rect -333 -2503 -287 -2457
rect -209 -2503 -163 -2457
rect -85 -2503 -39 -2457
rect 39 -2503 85 -2457
rect 163 -2503 209 -2457
rect 287 -2503 333 -2457
rect 411 -2503 457 -2457
rect 535 -2503 581 -2457
rect 659 -2503 705 -2457
rect 783 -2503 829 -2457
rect 907 -2503 953 -2457
rect 1031 -2503 1077 -2457
rect -1077 -2627 -1031 -2581
rect -953 -2627 -907 -2581
rect -829 -2627 -783 -2581
rect -705 -2627 -659 -2581
rect -581 -2627 -535 -2581
rect -457 -2627 -411 -2581
rect -333 -2627 -287 -2581
rect -209 -2627 -163 -2581
rect -85 -2627 -39 -2581
rect 39 -2627 85 -2581
rect 163 -2627 209 -2581
rect 287 -2627 333 -2581
rect 411 -2627 457 -2581
rect 535 -2627 581 -2581
rect 659 -2627 705 -2581
rect 783 -2627 829 -2581
rect 907 -2627 953 -2581
rect 1031 -2627 1077 -2581
rect -1077 -2751 -1031 -2705
rect -953 -2751 -907 -2705
rect -829 -2751 -783 -2705
rect -705 -2751 -659 -2705
rect -581 -2751 -535 -2705
rect -457 -2751 -411 -2705
rect -333 -2751 -287 -2705
rect -209 -2751 -163 -2705
rect -85 -2751 -39 -2705
rect 39 -2751 85 -2705
rect 163 -2751 209 -2705
rect 287 -2751 333 -2705
rect 411 -2751 457 -2705
rect 535 -2751 581 -2705
rect 659 -2751 705 -2705
rect 783 -2751 829 -2705
rect 907 -2751 953 -2705
rect 1031 -2751 1077 -2705
rect -1077 -2875 -1031 -2829
rect -953 -2875 -907 -2829
rect -829 -2875 -783 -2829
rect -705 -2875 -659 -2829
rect -581 -2875 -535 -2829
rect -457 -2875 -411 -2829
rect -333 -2875 -287 -2829
rect -209 -2875 -163 -2829
rect -85 -2875 -39 -2829
rect 39 -2875 85 -2829
rect 163 -2875 209 -2829
rect 287 -2875 333 -2829
rect 411 -2875 457 -2829
rect 535 -2875 581 -2829
rect 659 -2875 705 -2829
rect 783 -2875 829 -2829
rect 907 -2875 953 -2829
rect 1031 -2875 1077 -2829
rect -1077 -2999 -1031 -2953
rect -953 -2999 -907 -2953
rect -829 -2999 -783 -2953
rect -705 -2999 -659 -2953
rect -581 -2999 -535 -2953
rect -457 -2999 -411 -2953
rect -333 -2999 -287 -2953
rect -209 -2999 -163 -2953
rect -85 -2999 -39 -2953
rect 39 -2999 85 -2953
rect 163 -2999 209 -2953
rect 287 -2999 333 -2953
rect 411 -2999 457 -2953
rect 535 -2999 581 -2953
rect 659 -2999 705 -2953
rect 783 -2999 829 -2953
rect 907 -2999 953 -2953
rect 1031 -2999 1077 -2953
rect -1077 -3123 -1031 -3077
rect -953 -3123 -907 -3077
rect -829 -3123 -783 -3077
rect -705 -3123 -659 -3077
rect -581 -3123 -535 -3077
rect -457 -3123 -411 -3077
rect -333 -3123 -287 -3077
rect -209 -3123 -163 -3077
rect -85 -3123 -39 -3077
rect 39 -3123 85 -3077
rect 163 -3123 209 -3077
rect 287 -3123 333 -3077
rect 411 -3123 457 -3077
rect 535 -3123 581 -3077
rect 659 -3123 705 -3077
rect 783 -3123 829 -3077
rect 907 -3123 953 -3077
rect 1031 -3123 1077 -3077
rect -1077 -3247 -1031 -3201
rect -953 -3247 -907 -3201
rect -829 -3247 -783 -3201
rect -705 -3247 -659 -3201
rect -581 -3247 -535 -3201
rect -457 -3247 -411 -3201
rect -333 -3247 -287 -3201
rect -209 -3247 -163 -3201
rect -85 -3247 -39 -3201
rect 39 -3247 85 -3201
rect 163 -3247 209 -3201
rect 287 -3247 333 -3201
rect 411 -3247 457 -3201
rect 535 -3247 581 -3201
rect 659 -3247 705 -3201
rect 783 -3247 829 -3201
rect 907 -3247 953 -3201
rect 1031 -3247 1077 -3201
rect -1077 -3371 -1031 -3325
rect -953 -3371 -907 -3325
rect -829 -3371 -783 -3325
rect -705 -3371 -659 -3325
rect -581 -3371 -535 -3325
rect -457 -3371 -411 -3325
rect -333 -3371 -287 -3325
rect -209 -3371 -163 -3325
rect -85 -3371 -39 -3325
rect 39 -3371 85 -3325
rect 163 -3371 209 -3325
rect 287 -3371 333 -3325
rect 411 -3371 457 -3325
rect 535 -3371 581 -3325
rect 659 -3371 705 -3325
rect 783 -3371 829 -3325
rect 907 -3371 953 -3325
rect 1031 -3371 1077 -3325
rect -1077 -3495 -1031 -3449
rect -953 -3495 -907 -3449
rect -829 -3495 -783 -3449
rect -705 -3495 -659 -3449
rect -581 -3495 -535 -3449
rect -457 -3495 -411 -3449
rect -333 -3495 -287 -3449
rect -209 -3495 -163 -3449
rect -85 -3495 -39 -3449
rect 39 -3495 85 -3449
rect 163 -3495 209 -3449
rect 287 -3495 333 -3449
rect 411 -3495 457 -3449
rect 535 -3495 581 -3449
rect 659 -3495 705 -3449
rect 783 -3495 829 -3449
rect 907 -3495 953 -3449
rect 1031 -3495 1077 -3449
rect -1077 -3619 -1031 -3573
rect -953 -3619 -907 -3573
rect -829 -3619 -783 -3573
rect -705 -3619 -659 -3573
rect -581 -3619 -535 -3573
rect -457 -3619 -411 -3573
rect -333 -3619 -287 -3573
rect -209 -3619 -163 -3573
rect -85 -3619 -39 -3573
rect 39 -3619 85 -3573
rect 163 -3619 209 -3573
rect 287 -3619 333 -3573
rect 411 -3619 457 -3573
rect 535 -3619 581 -3573
rect 659 -3619 705 -3573
rect 783 -3619 829 -3573
rect 907 -3619 953 -3573
rect 1031 -3619 1077 -3573
rect -1077 -3743 -1031 -3697
rect -953 -3743 -907 -3697
rect -829 -3743 -783 -3697
rect -705 -3743 -659 -3697
rect -581 -3743 -535 -3697
rect -457 -3743 -411 -3697
rect -333 -3743 -287 -3697
rect -209 -3743 -163 -3697
rect -85 -3743 -39 -3697
rect 39 -3743 85 -3697
rect 163 -3743 209 -3697
rect 287 -3743 333 -3697
rect 411 -3743 457 -3697
rect 535 -3743 581 -3697
rect 659 -3743 705 -3697
rect 783 -3743 829 -3697
rect 907 -3743 953 -3697
rect 1031 -3743 1077 -3697
rect -1077 -3867 -1031 -3821
rect -953 -3867 -907 -3821
rect -829 -3867 -783 -3821
rect -705 -3867 -659 -3821
rect -581 -3867 -535 -3821
rect -457 -3867 -411 -3821
rect -333 -3867 -287 -3821
rect -209 -3867 -163 -3821
rect -85 -3867 -39 -3821
rect 39 -3867 85 -3821
rect 163 -3867 209 -3821
rect 287 -3867 333 -3821
rect 411 -3867 457 -3821
rect 535 -3867 581 -3821
rect 659 -3867 705 -3821
rect 783 -3867 829 -3821
rect 907 -3867 953 -3821
rect 1031 -3867 1077 -3821
rect -1077 -3991 -1031 -3945
rect -953 -3991 -907 -3945
rect -829 -3991 -783 -3945
rect -705 -3991 -659 -3945
rect -581 -3991 -535 -3945
rect -457 -3991 -411 -3945
rect -333 -3991 -287 -3945
rect -209 -3991 -163 -3945
rect -85 -3991 -39 -3945
rect 39 -3991 85 -3945
rect 163 -3991 209 -3945
rect 287 -3991 333 -3945
rect 411 -3991 457 -3945
rect 535 -3991 581 -3945
rect 659 -3991 705 -3945
rect 783 -3991 829 -3945
rect 907 -3991 953 -3945
rect 1031 -3991 1077 -3945
rect -1077 -4115 -1031 -4069
rect -953 -4115 -907 -4069
rect -829 -4115 -783 -4069
rect -705 -4115 -659 -4069
rect -581 -4115 -535 -4069
rect -457 -4115 -411 -4069
rect -333 -4115 -287 -4069
rect -209 -4115 -163 -4069
rect -85 -4115 -39 -4069
rect 39 -4115 85 -4069
rect 163 -4115 209 -4069
rect 287 -4115 333 -4069
rect 411 -4115 457 -4069
rect 535 -4115 581 -4069
rect 659 -4115 705 -4069
rect 783 -4115 829 -4069
rect 907 -4115 953 -4069
rect 1031 -4115 1077 -4069
rect -1077 -4239 -1031 -4193
rect -953 -4239 -907 -4193
rect -829 -4239 -783 -4193
rect -705 -4239 -659 -4193
rect -581 -4239 -535 -4193
rect -457 -4239 -411 -4193
rect -333 -4239 -287 -4193
rect -209 -4239 -163 -4193
rect -85 -4239 -39 -4193
rect 39 -4239 85 -4193
rect 163 -4239 209 -4193
rect 287 -4239 333 -4193
rect 411 -4239 457 -4193
rect 535 -4239 581 -4193
rect 659 -4239 705 -4193
rect 783 -4239 829 -4193
rect 907 -4239 953 -4193
rect 1031 -4239 1077 -4193
rect -1077 -4363 -1031 -4317
rect -953 -4363 -907 -4317
rect -829 -4363 -783 -4317
rect -705 -4363 -659 -4317
rect -581 -4363 -535 -4317
rect -457 -4363 -411 -4317
rect -333 -4363 -287 -4317
rect -209 -4363 -163 -4317
rect -85 -4363 -39 -4317
rect 39 -4363 85 -4317
rect 163 -4363 209 -4317
rect 287 -4363 333 -4317
rect 411 -4363 457 -4317
rect 535 -4363 581 -4317
rect 659 -4363 705 -4317
rect 783 -4363 829 -4317
rect 907 -4363 953 -4317
rect 1031 -4363 1077 -4317
rect -1077 -4487 -1031 -4441
rect -953 -4487 -907 -4441
rect -829 -4487 -783 -4441
rect -705 -4487 -659 -4441
rect -581 -4487 -535 -4441
rect -457 -4487 -411 -4441
rect -333 -4487 -287 -4441
rect -209 -4487 -163 -4441
rect -85 -4487 -39 -4441
rect 39 -4487 85 -4441
rect 163 -4487 209 -4441
rect 287 -4487 333 -4441
rect 411 -4487 457 -4441
rect 535 -4487 581 -4441
rect 659 -4487 705 -4441
rect 783 -4487 829 -4441
rect 907 -4487 953 -4441
rect 1031 -4487 1077 -4441
rect -1077 -4611 -1031 -4565
rect -953 -4611 -907 -4565
rect -829 -4611 -783 -4565
rect -705 -4611 -659 -4565
rect -581 -4611 -535 -4565
rect -457 -4611 -411 -4565
rect -333 -4611 -287 -4565
rect -209 -4611 -163 -4565
rect -85 -4611 -39 -4565
rect 39 -4611 85 -4565
rect 163 -4611 209 -4565
rect 287 -4611 333 -4565
rect 411 -4611 457 -4565
rect 535 -4611 581 -4565
rect 659 -4611 705 -4565
rect 783 -4611 829 -4565
rect 907 -4611 953 -4565
rect 1031 -4611 1077 -4565
rect -1077 -4735 -1031 -4689
rect -953 -4735 -907 -4689
rect -829 -4735 -783 -4689
rect -705 -4735 -659 -4689
rect -581 -4735 -535 -4689
rect -457 -4735 -411 -4689
rect -333 -4735 -287 -4689
rect -209 -4735 -163 -4689
rect -85 -4735 -39 -4689
rect 39 -4735 85 -4689
rect 163 -4735 209 -4689
rect 287 -4735 333 -4689
rect 411 -4735 457 -4689
rect 535 -4735 581 -4689
rect 659 -4735 705 -4689
rect 783 -4735 829 -4689
rect 907 -4735 953 -4689
rect 1031 -4735 1077 -4689
rect -1077 -4859 -1031 -4813
rect -953 -4859 -907 -4813
rect -829 -4859 -783 -4813
rect -705 -4859 -659 -4813
rect -581 -4859 -535 -4813
rect -457 -4859 -411 -4813
rect -333 -4859 -287 -4813
rect -209 -4859 -163 -4813
rect -85 -4859 -39 -4813
rect 39 -4859 85 -4813
rect 163 -4859 209 -4813
rect 287 -4859 333 -4813
rect 411 -4859 457 -4813
rect 535 -4859 581 -4813
rect 659 -4859 705 -4813
rect 783 -4859 829 -4813
rect 907 -4859 953 -4813
rect 1031 -4859 1077 -4813
rect -1077 -4983 -1031 -4937
rect -953 -4983 -907 -4937
rect -829 -4983 -783 -4937
rect -705 -4983 -659 -4937
rect -581 -4983 -535 -4937
rect -457 -4983 -411 -4937
rect -333 -4983 -287 -4937
rect -209 -4983 -163 -4937
rect -85 -4983 -39 -4937
rect 39 -4983 85 -4937
rect 163 -4983 209 -4937
rect 287 -4983 333 -4937
rect 411 -4983 457 -4937
rect 535 -4983 581 -4937
rect 659 -4983 705 -4937
rect 783 -4983 829 -4937
rect 907 -4983 953 -4937
rect 1031 -4983 1077 -4937
rect -1077 -5107 -1031 -5061
rect -953 -5107 -907 -5061
rect -829 -5107 -783 -5061
rect -705 -5107 -659 -5061
rect -581 -5107 -535 -5061
rect -457 -5107 -411 -5061
rect -333 -5107 -287 -5061
rect -209 -5107 -163 -5061
rect -85 -5107 -39 -5061
rect 39 -5107 85 -5061
rect 163 -5107 209 -5061
rect 287 -5107 333 -5061
rect 411 -5107 457 -5061
rect 535 -5107 581 -5061
rect 659 -5107 705 -5061
rect 783 -5107 829 -5061
rect 907 -5107 953 -5061
rect 1031 -5107 1077 -5061
rect -1077 -5231 -1031 -5185
rect -953 -5231 -907 -5185
rect -829 -5231 -783 -5185
rect -705 -5231 -659 -5185
rect -581 -5231 -535 -5185
rect -457 -5231 -411 -5185
rect -333 -5231 -287 -5185
rect -209 -5231 -163 -5185
rect -85 -5231 -39 -5185
rect 39 -5231 85 -5185
rect 163 -5231 209 -5185
rect 287 -5231 333 -5185
rect 411 -5231 457 -5185
rect 535 -5231 581 -5185
rect 659 -5231 705 -5185
rect 783 -5231 829 -5185
rect 907 -5231 953 -5185
rect 1031 -5231 1077 -5185
rect -1077 -5355 -1031 -5309
rect -953 -5355 -907 -5309
rect -829 -5355 -783 -5309
rect -705 -5355 -659 -5309
rect -581 -5355 -535 -5309
rect -457 -5355 -411 -5309
rect -333 -5355 -287 -5309
rect -209 -5355 -163 -5309
rect -85 -5355 -39 -5309
rect 39 -5355 85 -5309
rect 163 -5355 209 -5309
rect 287 -5355 333 -5309
rect 411 -5355 457 -5309
rect 535 -5355 581 -5309
rect 659 -5355 705 -5309
rect 783 -5355 829 -5309
rect 907 -5355 953 -5309
rect 1031 -5355 1077 -5309
rect -1077 -5479 -1031 -5433
rect -953 -5479 -907 -5433
rect -829 -5479 -783 -5433
rect -705 -5479 -659 -5433
rect -581 -5479 -535 -5433
rect -457 -5479 -411 -5433
rect -333 -5479 -287 -5433
rect -209 -5479 -163 -5433
rect -85 -5479 -39 -5433
rect 39 -5479 85 -5433
rect 163 -5479 209 -5433
rect 287 -5479 333 -5433
rect 411 -5479 457 -5433
rect 535 -5479 581 -5433
rect 659 -5479 705 -5433
rect 783 -5479 829 -5433
rect 907 -5479 953 -5433
rect 1031 -5479 1077 -5433
rect -1077 -5603 -1031 -5557
rect -953 -5603 -907 -5557
rect -829 -5603 -783 -5557
rect -705 -5603 -659 -5557
rect -581 -5603 -535 -5557
rect -457 -5603 -411 -5557
rect -333 -5603 -287 -5557
rect -209 -5603 -163 -5557
rect -85 -5603 -39 -5557
rect 39 -5603 85 -5557
rect 163 -5603 209 -5557
rect 287 -5603 333 -5557
rect 411 -5603 457 -5557
rect 535 -5603 581 -5557
rect 659 -5603 705 -5557
rect 783 -5603 829 -5557
rect 907 -5603 953 -5557
rect 1031 -5603 1077 -5557
rect -1077 -5727 -1031 -5681
rect -953 -5727 -907 -5681
rect -829 -5727 -783 -5681
rect -705 -5727 -659 -5681
rect -581 -5727 -535 -5681
rect -457 -5727 -411 -5681
rect -333 -5727 -287 -5681
rect -209 -5727 -163 -5681
rect -85 -5727 -39 -5681
rect 39 -5727 85 -5681
rect 163 -5727 209 -5681
rect 287 -5727 333 -5681
rect 411 -5727 457 -5681
rect 535 -5727 581 -5681
rect 659 -5727 705 -5681
rect 783 -5727 829 -5681
rect 907 -5727 953 -5681
rect 1031 -5727 1077 -5681
rect -1077 -5851 -1031 -5805
rect -953 -5851 -907 -5805
rect -829 -5851 -783 -5805
rect -705 -5851 -659 -5805
rect -581 -5851 -535 -5805
rect -457 -5851 -411 -5805
rect -333 -5851 -287 -5805
rect -209 -5851 -163 -5805
rect -85 -5851 -39 -5805
rect 39 -5851 85 -5805
rect 163 -5851 209 -5805
rect 287 -5851 333 -5805
rect 411 -5851 457 -5805
rect 535 -5851 581 -5805
rect 659 -5851 705 -5805
rect 783 -5851 829 -5805
rect 907 -5851 953 -5805
rect 1031 -5851 1077 -5805
<< metal1 >>
rect -1088 5851 1088 5862
rect -1088 5805 -1077 5851
rect -1031 5805 -953 5851
rect -907 5805 -829 5851
rect -783 5805 -705 5851
rect -659 5805 -581 5851
rect -535 5805 -457 5851
rect -411 5805 -333 5851
rect -287 5805 -209 5851
rect -163 5805 -85 5851
rect -39 5805 39 5851
rect 85 5805 163 5851
rect 209 5805 287 5851
rect 333 5805 411 5851
rect 457 5805 535 5851
rect 581 5805 659 5851
rect 705 5805 783 5851
rect 829 5805 907 5851
rect 953 5805 1031 5851
rect 1077 5805 1088 5851
rect -1088 5727 1088 5805
rect -1088 5681 -1077 5727
rect -1031 5681 -953 5727
rect -907 5681 -829 5727
rect -783 5681 -705 5727
rect -659 5681 -581 5727
rect -535 5681 -457 5727
rect -411 5681 -333 5727
rect -287 5681 -209 5727
rect -163 5681 -85 5727
rect -39 5681 39 5727
rect 85 5681 163 5727
rect 209 5681 287 5727
rect 333 5681 411 5727
rect 457 5681 535 5727
rect 581 5681 659 5727
rect 705 5681 783 5727
rect 829 5681 907 5727
rect 953 5681 1031 5727
rect 1077 5681 1088 5727
rect -1088 5603 1088 5681
rect -1088 5557 -1077 5603
rect -1031 5557 -953 5603
rect -907 5557 -829 5603
rect -783 5557 -705 5603
rect -659 5557 -581 5603
rect -535 5557 -457 5603
rect -411 5557 -333 5603
rect -287 5557 -209 5603
rect -163 5557 -85 5603
rect -39 5557 39 5603
rect 85 5557 163 5603
rect 209 5557 287 5603
rect 333 5557 411 5603
rect 457 5557 535 5603
rect 581 5557 659 5603
rect 705 5557 783 5603
rect 829 5557 907 5603
rect 953 5557 1031 5603
rect 1077 5557 1088 5603
rect -1088 5479 1088 5557
rect -1088 5433 -1077 5479
rect -1031 5433 -953 5479
rect -907 5433 -829 5479
rect -783 5433 -705 5479
rect -659 5433 -581 5479
rect -535 5433 -457 5479
rect -411 5433 -333 5479
rect -287 5433 -209 5479
rect -163 5433 -85 5479
rect -39 5433 39 5479
rect 85 5433 163 5479
rect 209 5433 287 5479
rect 333 5433 411 5479
rect 457 5433 535 5479
rect 581 5433 659 5479
rect 705 5433 783 5479
rect 829 5433 907 5479
rect 953 5433 1031 5479
rect 1077 5433 1088 5479
rect -1088 5355 1088 5433
rect -1088 5309 -1077 5355
rect -1031 5309 -953 5355
rect -907 5309 -829 5355
rect -783 5309 -705 5355
rect -659 5309 -581 5355
rect -535 5309 -457 5355
rect -411 5309 -333 5355
rect -287 5309 -209 5355
rect -163 5309 -85 5355
rect -39 5309 39 5355
rect 85 5309 163 5355
rect 209 5309 287 5355
rect 333 5309 411 5355
rect 457 5309 535 5355
rect 581 5309 659 5355
rect 705 5309 783 5355
rect 829 5309 907 5355
rect 953 5309 1031 5355
rect 1077 5309 1088 5355
rect -1088 5231 1088 5309
rect -1088 5185 -1077 5231
rect -1031 5185 -953 5231
rect -907 5185 -829 5231
rect -783 5185 -705 5231
rect -659 5185 -581 5231
rect -535 5185 -457 5231
rect -411 5185 -333 5231
rect -287 5185 -209 5231
rect -163 5185 -85 5231
rect -39 5185 39 5231
rect 85 5185 163 5231
rect 209 5185 287 5231
rect 333 5185 411 5231
rect 457 5185 535 5231
rect 581 5185 659 5231
rect 705 5185 783 5231
rect 829 5185 907 5231
rect 953 5185 1031 5231
rect 1077 5185 1088 5231
rect -1088 5107 1088 5185
rect -1088 5061 -1077 5107
rect -1031 5061 -953 5107
rect -907 5061 -829 5107
rect -783 5061 -705 5107
rect -659 5061 -581 5107
rect -535 5061 -457 5107
rect -411 5061 -333 5107
rect -287 5061 -209 5107
rect -163 5061 -85 5107
rect -39 5061 39 5107
rect 85 5061 163 5107
rect 209 5061 287 5107
rect 333 5061 411 5107
rect 457 5061 535 5107
rect 581 5061 659 5107
rect 705 5061 783 5107
rect 829 5061 907 5107
rect 953 5061 1031 5107
rect 1077 5061 1088 5107
rect -1088 4983 1088 5061
rect -1088 4937 -1077 4983
rect -1031 4937 -953 4983
rect -907 4937 -829 4983
rect -783 4937 -705 4983
rect -659 4937 -581 4983
rect -535 4937 -457 4983
rect -411 4937 -333 4983
rect -287 4937 -209 4983
rect -163 4937 -85 4983
rect -39 4937 39 4983
rect 85 4937 163 4983
rect 209 4937 287 4983
rect 333 4937 411 4983
rect 457 4937 535 4983
rect 581 4937 659 4983
rect 705 4937 783 4983
rect 829 4937 907 4983
rect 953 4937 1031 4983
rect 1077 4937 1088 4983
rect -1088 4859 1088 4937
rect -1088 4813 -1077 4859
rect -1031 4813 -953 4859
rect -907 4813 -829 4859
rect -783 4813 -705 4859
rect -659 4813 -581 4859
rect -535 4813 -457 4859
rect -411 4813 -333 4859
rect -287 4813 -209 4859
rect -163 4813 -85 4859
rect -39 4813 39 4859
rect 85 4813 163 4859
rect 209 4813 287 4859
rect 333 4813 411 4859
rect 457 4813 535 4859
rect 581 4813 659 4859
rect 705 4813 783 4859
rect 829 4813 907 4859
rect 953 4813 1031 4859
rect 1077 4813 1088 4859
rect -1088 4735 1088 4813
rect -1088 4689 -1077 4735
rect -1031 4689 -953 4735
rect -907 4689 -829 4735
rect -783 4689 -705 4735
rect -659 4689 -581 4735
rect -535 4689 -457 4735
rect -411 4689 -333 4735
rect -287 4689 -209 4735
rect -163 4689 -85 4735
rect -39 4689 39 4735
rect 85 4689 163 4735
rect 209 4689 287 4735
rect 333 4689 411 4735
rect 457 4689 535 4735
rect 581 4689 659 4735
rect 705 4689 783 4735
rect 829 4689 907 4735
rect 953 4689 1031 4735
rect 1077 4689 1088 4735
rect -1088 4611 1088 4689
rect -1088 4565 -1077 4611
rect -1031 4565 -953 4611
rect -907 4565 -829 4611
rect -783 4565 -705 4611
rect -659 4565 -581 4611
rect -535 4565 -457 4611
rect -411 4565 -333 4611
rect -287 4565 -209 4611
rect -163 4565 -85 4611
rect -39 4565 39 4611
rect 85 4565 163 4611
rect 209 4565 287 4611
rect 333 4565 411 4611
rect 457 4565 535 4611
rect 581 4565 659 4611
rect 705 4565 783 4611
rect 829 4565 907 4611
rect 953 4565 1031 4611
rect 1077 4565 1088 4611
rect -1088 4487 1088 4565
rect -1088 4441 -1077 4487
rect -1031 4441 -953 4487
rect -907 4441 -829 4487
rect -783 4441 -705 4487
rect -659 4441 -581 4487
rect -535 4441 -457 4487
rect -411 4441 -333 4487
rect -287 4441 -209 4487
rect -163 4441 -85 4487
rect -39 4441 39 4487
rect 85 4441 163 4487
rect 209 4441 287 4487
rect 333 4441 411 4487
rect 457 4441 535 4487
rect 581 4441 659 4487
rect 705 4441 783 4487
rect 829 4441 907 4487
rect 953 4441 1031 4487
rect 1077 4441 1088 4487
rect -1088 4363 1088 4441
rect -1088 4317 -1077 4363
rect -1031 4317 -953 4363
rect -907 4317 -829 4363
rect -783 4317 -705 4363
rect -659 4317 -581 4363
rect -535 4317 -457 4363
rect -411 4317 -333 4363
rect -287 4317 -209 4363
rect -163 4317 -85 4363
rect -39 4317 39 4363
rect 85 4317 163 4363
rect 209 4317 287 4363
rect 333 4317 411 4363
rect 457 4317 535 4363
rect 581 4317 659 4363
rect 705 4317 783 4363
rect 829 4317 907 4363
rect 953 4317 1031 4363
rect 1077 4317 1088 4363
rect -1088 4239 1088 4317
rect -1088 4193 -1077 4239
rect -1031 4193 -953 4239
rect -907 4193 -829 4239
rect -783 4193 -705 4239
rect -659 4193 -581 4239
rect -535 4193 -457 4239
rect -411 4193 -333 4239
rect -287 4193 -209 4239
rect -163 4193 -85 4239
rect -39 4193 39 4239
rect 85 4193 163 4239
rect 209 4193 287 4239
rect 333 4193 411 4239
rect 457 4193 535 4239
rect 581 4193 659 4239
rect 705 4193 783 4239
rect 829 4193 907 4239
rect 953 4193 1031 4239
rect 1077 4193 1088 4239
rect -1088 4115 1088 4193
rect -1088 4069 -1077 4115
rect -1031 4069 -953 4115
rect -907 4069 -829 4115
rect -783 4069 -705 4115
rect -659 4069 -581 4115
rect -535 4069 -457 4115
rect -411 4069 -333 4115
rect -287 4069 -209 4115
rect -163 4069 -85 4115
rect -39 4069 39 4115
rect 85 4069 163 4115
rect 209 4069 287 4115
rect 333 4069 411 4115
rect 457 4069 535 4115
rect 581 4069 659 4115
rect 705 4069 783 4115
rect 829 4069 907 4115
rect 953 4069 1031 4115
rect 1077 4069 1088 4115
rect -1088 3991 1088 4069
rect -1088 3945 -1077 3991
rect -1031 3945 -953 3991
rect -907 3945 -829 3991
rect -783 3945 -705 3991
rect -659 3945 -581 3991
rect -535 3945 -457 3991
rect -411 3945 -333 3991
rect -287 3945 -209 3991
rect -163 3945 -85 3991
rect -39 3945 39 3991
rect 85 3945 163 3991
rect 209 3945 287 3991
rect 333 3945 411 3991
rect 457 3945 535 3991
rect 581 3945 659 3991
rect 705 3945 783 3991
rect 829 3945 907 3991
rect 953 3945 1031 3991
rect 1077 3945 1088 3991
rect -1088 3867 1088 3945
rect -1088 3821 -1077 3867
rect -1031 3821 -953 3867
rect -907 3821 -829 3867
rect -783 3821 -705 3867
rect -659 3821 -581 3867
rect -535 3821 -457 3867
rect -411 3821 -333 3867
rect -287 3821 -209 3867
rect -163 3821 -85 3867
rect -39 3821 39 3867
rect 85 3821 163 3867
rect 209 3821 287 3867
rect 333 3821 411 3867
rect 457 3821 535 3867
rect 581 3821 659 3867
rect 705 3821 783 3867
rect 829 3821 907 3867
rect 953 3821 1031 3867
rect 1077 3821 1088 3867
rect -1088 3743 1088 3821
rect -1088 3697 -1077 3743
rect -1031 3697 -953 3743
rect -907 3697 -829 3743
rect -783 3697 -705 3743
rect -659 3697 -581 3743
rect -535 3697 -457 3743
rect -411 3697 -333 3743
rect -287 3697 -209 3743
rect -163 3697 -85 3743
rect -39 3697 39 3743
rect 85 3697 163 3743
rect 209 3697 287 3743
rect 333 3697 411 3743
rect 457 3697 535 3743
rect 581 3697 659 3743
rect 705 3697 783 3743
rect 829 3697 907 3743
rect 953 3697 1031 3743
rect 1077 3697 1088 3743
rect -1088 3619 1088 3697
rect -1088 3573 -1077 3619
rect -1031 3573 -953 3619
rect -907 3573 -829 3619
rect -783 3573 -705 3619
rect -659 3573 -581 3619
rect -535 3573 -457 3619
rect -411 3573 -333 3619
rect -287 3573 -209 3619
rect -163 3573 -85 3619
rect -39 3573 39 3619
rect 85 3573 163 3619
rect 209 3573 287 3619
rect 333 3573 411 3619
rect 457 3573 535 3619
rect 581 3573 659 3619
rect 705 3573 783 3619
rect 829 3573 907 3619
rect 953 3573 1031 3619
rect 1077 3573 1088 3619
rect -1088 3495 1088 3573
rect -1088 3449 -1077 3495
rect -1031 3449 -953 3495
rect -907 3449 -829 3495
rect -783 3449 -705 3495
rect -659 3449 -581 3495
rect -535 3449 -457 3495
rect -411 3449 -333 3495
rect -287 3449 -209 3495
rect -163 3449 -85 3495
rect -39 3449 39 3495
rect 85 3449 163 3495
rect 209 3449 287 3495
rect 333 3449 411 3495
rect 457 3449 535 3495
rect 581 3449 659 3495
rect 705 3449 783 3495
rect 829 3449 907 3495
rect 953 3449 1031 3495
rect 1077 3449 1088 3495
rect -1088 3371 1088 3449
rect -1088 3325 -1077 3371
rect -1031 3325 -953 3371
rect -907 3325 -829 3371
rect -783 3325 -705 3371
rect -659 3325 -581 3371
rect -535 3325 -457 3371
rect -411 3325 -333 3371
rect -287 3325 -209 3371
rect -163 3325 -85 3371
rect -39 3325 39 3371
rect 85 3325 163 3371
rect 209 3325 287 3371
rect 333 3325 411 3371
rect 457 3325 535 3371
rect 581 3325 659 3371
rect 705 3325 783 3371
rect 829 3325 907 3371
rect 953 3325 1031 3371
rect 1077 3325 1088 3371
rect -1088 3247 1088 3325
rect -1088 3201 -1077 3247
rect -1031 3201 -953 3247
rect -907 3201 -829 3247
rect -783 3201 -705 3247
rect -659 3201 -581 3247
rect -535 3201 -457 3247
rect -411 3201 -333 3247
rect -287 3201 -209 3247
rect -163 3201 -85 3247
rect -39 3201 39 3247
rect 85 3201 163 3247
rect 209 3201 287 3247
rect 333 3201 411 3247
rect 457 3201 535 3247
rect 581 3201 659 3247
rect 705 3201 783 3247
rect 829 3201 907 3247
rect 953 3201 1031 3247
rect 1077 3201 1088 3247
rect -1088 3123 1088 3201
rect -1088 3077 -1077 3123
rect -1031 3077 -953 3123
rect -907 3077 -829 3123
rect -783 3077 -705 3123
rect -659 3077 -581 3123
rect -535 3077 -457 3123
rect -411 3077 -333 3123
rect -287 3077 -209 3123
rect -163 3077 -85 3123
rect -39 3077 39 3123
rect 85 3077 163 3123
rect 209 3077 287 3123
rect 333 3077 411 3123
rect 457 3077 535 3123
rect 581 3077 659 3123
rect 705 3077 783 3123
rect 829 3077 907 3123
rect 953 3077 1031 3123
rect 1077 3077 1088 3123
rect -1088 2999 1088 3077
rect -1088 2953 -1077 2999
rect -1031 2953 -953 2999
rect -907 2953 -829 2999
rect -783 2953 -705 2999
rect -659 2953 -581 2999
rect -535 2953 -457 2999
rect -411 2953 -333 2999
rect -287 2953 -209 2999
rect -163 2953 -85 2999
rect -39 2953 39 2999
rect 85 2953 163 2999
rect 209 2953 287 2999
rect 333 2953 411 2999
rect 457 2953 535 2999
rect 581 2953 659 2999
rect 705 2953 783 2999
rect 829 2953 907 2999
rect 953 2953 1031 2999
rect 1077 2953 1088 2999
rect -1088 2875 1088 2953
rect -1088 2829 -1077 2875
rect -1031 2829 -953 2875
rect -907 2829 -829 2875
rect -783 2829 -705 2875
rect -659 2829 -581 2875
rect -535 2829 -457 2875
rect -411 2829 -333 2875
rect -287 2829 -209 2875
rect -163 2829 -85 2875
rect -39 2829 39 2875
rect 85 2829 163 2875
rect 209 2829 287 2875
rect 333 2829 411 2875
rect 457 2829 535 2875
rect 581 2829 659 2875
rect 705 2829 783 2875
rect 829 2829 907 2875
rect 953 2829 1031 2875
rect 1077 2829 1088 2875
rect -1088 2751 1088 2829
rect -1088 2705 -1077 2751
rect -1031 2705 -953 2751
rect -907 2705 -829 2751
rect -783 2705 -705 2751
rect -659 2705 -581 2751
rect -535 2705 -457 2751
rect -411 2705 -333 2751
rect -287 2705 -209 2751
rect -163 2705 -85 2751
rect -39 2705 39 2751
rect 85 2705 163 2751
rect 209 2705 287 2751
rect 333 2705 411 2751
rect 457 2705 535 2751
rect 581 2705 659 2751
rect 705 2705 783 2751
rect 829 2705 907 2751
rect 953 2705 1031 2751
rect 1077 2705 1088 2751
rect -1088 2627 1088 2705
rect -1088 2581 -1077 2627
rect -1031 2581 -953 2627
rect -907 2581 -829 2627
rect -783 2581 -705 2627
rect -659 2581 -581 2627
rect -535 2581 -457 2627
rect -411 2581 -333 2627
rect -287 2581 -209 2627
rect -163 2581 -85 2627
rect -39 2581 39 2627
rect 85 2581 163 2627
rect 209 2581 287 2627
rect 333 2581 411 2627
rect 457 2581 535 2627
rect 581 2581 659 2627
rect 705 2581 783 2627
rect 829 2581 907 2627
rect 953 2581 1031 2627
rect 1077 2581 1088 2627
rect -1088 2503 1088 2581
rect -1088 2457 -1077 2503
rect -1031 2457 -953 2503
rect -907 2457 -829 2503
rect -783 2457 -705 2503
rect -659 2457 -581 2503
rect -535 2457 -457 2503
rect -411 2457 -333 2503
rect -287 2457 -209 2503
rect -163 2457 -85 2503
rect -39 2457 39 2503
rect 85 2457 163 2503
rect 209 2457 287 2503
rect 333 2457 411 2503
rect 457 2457 535 2503
rect 581 2457 659 2503
rect 705 2457 783 2503
rect 829 2457 907 2503
rect 953 2457 1031 2503
rect 1077 2457 1088 2503
rect -1088 2379 1088 2457
rect -1088 2333 -1077 2379
rect -1031 2333 -953 2379
rect -907 2333 -829 2379
rect -783 2333 -705 2379
rect -659 2333 -581 2379
rect -535 2333 -457 2379
rect -411 2333 -333 2379
rect -287 2333 -209 2379
rect -163 2333 -85 2379
rect -39 2333 39 2379
rect 85 2333 163 2379
rect 209 2333 287 2379
rect 333 2333 411 2379
rect 457 2333 535 2379
rect 581 2333 659 2379
rect 705 2333 783 2379
rect 829 2333 907 2379
rect 953 2333 1031 2379
rect 1077 2333 1088 2379
rect -1088 2255 1088 2333
rect -1088 2209 -1077 2255
rect -1031 2209 -953 2255
rect -907 2209 -829 2255
rect -783 2209 -705 2255
rect -659 2209 -581 2255
rect -535 2209 -457 2255
rect -411 2209 -333 2255
rect -287 2209 -209 2255
rect -163 2209 -85 2255
rect -39 2209 39 2255
rect 85 2209 163 2255
rect 209 2209 287 2255
rect 333 2209 411 2255
rect 457 2209 535 2255
rect 581 2209 659 2255
rect 705 2209 783 2255
rect 829 2209 907 2255
rect 953 2209 1031 2255
rect 1077 2209 1088 2255
rect -1088 2131 1088 2209
rect -1088 2085 -1077 2131
rect -1031 2085 -953 2131
rect -907 2085 -829 2131
rect -783 2085 -705 2131
rect -659 2085 -581 2131
rect -535 2085 -457 2131
rect -411 2085 -333 2131
rect -287 2085 -209 2131
rect -163 2085 -85 2131
rect -39 2085 39 2131
rect 85 2085 163 2131
rect 209 2085 287 2131
rect 333 2085 411 2131
rect 457 2085 535 2131
rect 581 2085 659 2131
rect 705 2085 783 2131
rect 829 2085 907 2131
rect 953 2085 1031 2131
rect 1077 2085 1088 2131
rect -1088 2007 1088 2085
rect -1088 1961 -1077 2007
rect -1031 1961 -953 2007
rect -907 1961 -829 2007
rect -783 1961 -705 2007
rect -659 1961 -581 2007
rect -535 1961 -457 2007
rect -411 1961 -333 2007
rect -287 1961 -209 2007
rect -163 1961 -85 2007
rect -39 1961 39 2007
rect 85 1961 163 2007
rect 209 1961 287 2007
rect 333 1961 411 2007
rect 457 1961 535 2007
rect 581 1961 659 2007
rect 705 1961 783 2007
rect 829 1961 907 2007
rect 953 1961 1031 2007
rect 1077 1961 1088 2007
rect -1088 1883 1088 1961
rect -1088 1837 -1077 1883
rect -1031 1837 -953 1883
rect -907 1837 -829 1883
rect -783 1837 -705 1883
rect -659 1837 -581 1883
rect -535 1837 -457 1883
rect -411 1837 -333 1883
rect -287 1837 -209 1883
rect -163 1837 -85 1883
rect -39 1837 39 1883
rect 85 1837 163 1883
rect 209 1837 287 1883
rect 333 1837 411 1883
rect 457 1837 535 1883
rect 581 1837 659 1883
rect 705 1837 783 1883
rect 829 1837 907 1883
rect 953 1837 1031 1883
rect 1077 1837 1088 1883
rect -1088 1759 1088 1837
rect -1088 1713 -1077 1759
rect -1031 1713 -953 1759
rect -907 1713 -829 1759
rect -783 1713 -705 1759
rect -659 1713 -581 1759
rect -535 1713 -457 1759
rect -411 1713 -333 1759
rect -287 1713 -209 1759
rect -163 1713 -85 1759
rect -39 1713 39 1759
rect 85 1713 163 1759
rect 209 1713 287 1759
rect 333 1713 411 1759
rect 457 1713 535 1759
rect 581 1713 659 1759
rect 705 1713 783 1759
rect 829 1713 907 1759
rect 953 1713 1031 1759
rect 1077 1713 1088 1759
rect -1088 1635 1088 1713
rect -1088 1589 -1077 1635
rect -1031 1589 -953 1635
rect -907 1589 -829 1635
rect -783 1589 -705 1635
rect -659 1589 -581 1635
rect -535 1589 -457 1635
rect -411 1589 -333 1635
rect -287 1589 -209 1635
rect -163 1589 -85 1635
rect -39 1589 39 1635
rect 85 1589 163 1635
rect 209 1589 287 1635
rect 333 1589 411 1635
rect 457 1589 535 1635
rect 581 1589 659 1635
rect 705 1589 783 1635
rect 829 1589 907 1635
rect 953 1589 1031 1635
rect 1077 1589 1088 1635
rect -1088 1511 1088 1589
rect -1088 1465 -1077 1511
rect -1031 1465 -953 1511
rect -907 1465 -829 1511
rect -783 1465 -705 1511
rect -659 1465 -581 1511
rect -535 1465 -457 1511
rect -411 1465 -333 1511
rect -287 1465 -209 1511
rect -163 1465 -85 1511
rect -39 1465 39 1511
rect 85 1465 163 1511
rect 209 1465 287 1511
rect 333 1465 411 1511
rect 457 1465 535 1511
rect 581 1465 659 1511
rect 705 1465 783 1511
rect 829 1465 907 1511
rect 953 1465 1031 1511
rect 1077 1465 1088 1511
rect -1088 1387 1088 1465
rect -1088 1341 -1077 1387
rect -1031 1341 -953 1387
rect -907 1341 -829 1387
rect -783 1341 -705 1387
rect -659 1341 -581 1387
rect -535 1341 -457 1387
rect -411 1341 -333 1387
rect -287 1341 -209 1387
rect -163 1341 -85 1387
rect -39 1341 39 1387
rect 85 1341 163 1387
rect 209 1341 287 1387
rect 333 1341 411 1387
rect 457 1341 535 1387
rect 581 1341 659 1387
rect 705 1341 783 1387
rect 829 1341 907 1387
rect 953 1341 1031 1387
rect 1077 1341 1088 1387
rect -1088 1263 1088 1341
rect -1088 1217 -1077 1263
rect -1031 1217 -953 1263
rect -907 1217 -829 1263
rect -783 1217 -705 1263
rect -659 1217 -581 1263
rect -535 1217 -457 1263
rect -411 1217 -333 1263
rect -287 1217 -209 1263
rect -163 1217 -85 1263
rect -39 1217 39 1263
rect 85 1217 163 1263
rect 209 1217 287 1263
rect 333 1217 411 1263
rect 457 1217 535 1263
rect 581 1217 659 1263
rect 705 1217 783 1263
rect 829 1217 907 1263
rect 953 1217 1031 1263
rect 1077 1217 1088 1263
rect -1088 1139 1088 1217
rect -1088 1093 -1077 1139
rect -1031 1093 -953 1139
rect -907 1093 -829 1139
rect -783 1093 -705 1139
rect -659 1093 -581 1139
rect -535 1093 -457 1139
rect -411 1093 -333 1139
rect -287 1093 -209 1139
rect -163 1093 -85 1139
rect -39 1093 39 1139
rect 85 1093 163 1139
rect 209 1093 287 1139
rect 333 1093 411 1139
rect 457 1093 535 1139
rect 581 1093 659 1139
rect 705 1093 783 1139
rect 829 1093 907 1139
rect 953 1093 1031 1139
rect 1077 1093 1088 1139
rect -1088 1015 1088 1093
rect -1088 969 -1077 1015
rect -1031 969 -953 1015
rect -907 969 -829 1015
rect -783 969 -705 1015
rect -659 969 -581 1015
rect -535 969 -457 1015
rect -411 969 -333 1015
rect -287 969 -209 1015
rect -163 969 -85 1015
rect -39 969 39 1015
rect 85 969 163 1015
rect 209 969 287 1015
rect 333 969 411 1015
rect 457 969 535 1015
rect 581 969 659 1015
rect 705 969 783 1015
rect 829 969 907 1015
rect 953 969 1031 1015
rect 1077 969 1088 1015
rect -1088 891 1088 969
rect -1088 845 -1077 891
rect -1031 845 -953 891
rect -907 845 -829 891
rect -783 845 -705 891
rect -659 845 -581 891
rect -535 845 -457 891
rect -411 845 -333 891
rect -287 845 -209 891
rect -163 845 -85 891
rect -39 845 39 891
rect 85 845 163 891
rect 209 845 287 891
rect 333 845 411 891
rect 457 845 535 891
rect 581 845 659 891
rect 705 845 783 891
rect 829 845 907 891
rect 953 845 1031 891
rect 1077 845 1088 891
rect -1088 767 1088 845
rect -1088 721 -1077 767
rect -1031 721 -953 767
rect -907 721 -829 767
rect -783 721 -705 767
rect -659 721 -581 767
rect -535 721 -457 767
rect -411 721 -333 767
rect -287 721 -209 767
rect -163 721 -85 767
rect -39 721 39 767
rect 85 721 163 767
rect 209 721 287 767
rect 333 721 411 767
rect 457 721 535 767
rect 581 721 659 767
rect 705 721 783 767
rect 829 721 907 767
rect 953 721 1031 767
rect 1077 721 1088 767
rect -1088 643 1088 721
rect -1088 597 -1077 643
rect -1031 597 -953 643
rect -907 597 -829 643
rect -783 597 -705 643
rect -659 597 -581 643
rect -535 597 -457 643
rect -411 597 -333 643
rect -287 597 -209 643
rect -163 597 -85 643
rect -39 597 39 643
rect 85 597 163 643
rect 209 597 287 643
rect 333 597 411 643
rect 457 597 535 643
rect 581 597 659 643
rect 705 597 783 643
rect 829 597 907 643
rect 953 597 1031 643
rect 1077 597 1088 643
rect -1088 519 1088 597
rect -1088 473 -1077 519
rect -1031 473 -953 519
rect -907 473 -829 519
rect -783 473 -705 519
rect -659 473 -581 519
rect -535 473 -457 519
rect -411 473 -333 519
rect -287 473 -209 519
rect -163 473 -85 519
rect -39 473 39 519
rect 85 473 163 519
rect 209 473 287 519
rect 333 473 411 519
rect 457 473 535 519
rect 581 473 659 519
rect 705 473 783 519
rect 829 473 907 519
rect 953 473 1031 519
rect 1077 473 1088 519
rect -1088 395 1088 473
rect -1088 349 -1077 395
rect -1031 349 -953 395
rect -907 349 -829 395
rect -783 349 -705 395
rect -659 349 -581 395
rect -535 349 -457 395
rect -411 349 -333 395
rect -287 349 -209 395
rect -163 349 -85 395
rect -39 349 39 395
rect 85 349 163 395
rect 209 349 287 395
rect 333 349 411 395
rect 457 349 535 395
rect 581 349 659 395
rect 705 349 783 395
rect 829 349 907 395
rect 953 349 1031 395
rect 1077 349 1088 395
rect -1088 271 1088 349
rect -1088 225 -1077 271
rect -1031 225 -953 271
rect -907 225 -829 271
rect -783 225 -705 271
rect -659 225 -581 271
rect -535 225 -457 271
rect -411 225 -333 271
rect -287 225 -209 271
rect -163 225 -85 271
rect -39 225 39 271
rect 85 225 163 271
rect 209 225 287 271
rect 333 225 411 271
rect 457 225 535 271
rect 581 225 659 271
rect 705 225 783 271
rect 829 225 907 271
rect 953 225 1031 271
rect 1077 225 1088 271
rect -1088 147 1088 225
rect -1088 101 -1077 147
rect -1031 101 -953 147
rect -907 101 -829 147
rect -783 101 -705 147
rect -659 101 -581 147
rect -535 101 -457 147
rect -411 101 -333 147
rect -287 101 -209 147
rect -163 101 -85 147
rect -39 101 39 147
rect 85 101 163 147
rect 209 101 287 147
rect 333 101 411 147
rect 457 101 535 147
rect 581 101 659 147
rect 705 101 783 147
rect 829 101 907 147
rect 953 101 1031 147
rect 1077 101 1088 147
rect -1088 23 1088 101
rect -1088 -23 -1077 23
rect -1031 -23 -953 23
rect -907 -23 -829 23
rect -783 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 783 23
rect 829 -23 907 23
rect 953 -23 1031 23
rect 1077 -23 1088 23
rect -1088 -101 1088 -23
rect -1088 -147 -1077 -101
rect -1031 -147 -953 -101
rect -907 -147 -829 -101
rect -783 -147 -705 -101
rect -659 -147 -581 -101
rect -535 -147 -457 -101
rect -411 -147 -333 -101
rect -287 -147 -209 -101
rect -163 -147 -85 -101
rect -39 -147 39 -101
rect 85 -147 163 -101
rect 209 -147 287 -101
rect 333 -147 411 -101
rect 457 -147 535 -101
rect 581 -147 659 -101
rect 705 -147 783 -101
rect 829 -147 907 -101
rect 953 -147 1031 -101
rect 1077 -147 1088 -101
rect -1088 -225 1088 -147
rect -1088 -271 -1077 -225
rect -1031 -271 -953 -225
rect -907 -271 -829 -225
rect -783 -271 -705 -225
rect -659 -271 -581 -225
rect -535 -271 -457 -225
rect -411 -271 -333 -225
rect -287 -271 -209 -225
rect -163 -271 -85 -225
rect -39 -271 39 -225
rect 85 -271 163 -225
rect 209 -271 287 -225
rect 333 -271 411 -225
rect 457 -271 535 -225
rect 581 -271 659 -225
rect 705 -271 783 -225
rect 829 -271 907 -225
rect 953 -271 1031 -225
rect 1077 -271 1088 -225
rect -1088 -349 1088 -271
rect -1088 -395 -1077 -349
rect -1031 -395 -953 -349
rect -907 -395 -829 -349
rect -783 -395 -705 -349
rect -659 -395 -581 -349
rect -535 -395 -457 -349
rect -411 -395 -333 -349
rect -287 -395 -209 -349
rect -163 -395 -85 -349
rect -39 -395 39 -349
rect 85 -395 163 -349
rect 209 -395 287 -349
rect 333 -395 411 -349
rect 457 -395 535 -349
rect 581 -395 659 -349
rect 705 -395 783 -349
rect 829 -395 907 -349
rect 953 -395 1031 -349
rect 1077 -395 1088 -349
rect -1088 -473 1088 -395
rect -1088 -519 -1077 -473
rect -1031 -519 -953 -473
rect -907 -519 -829 -473
rect -783 -519 -705 -473
rect -659 -519 -581 -473
rect -535 -519 -457 -473
rect -411 -519 -333 -473
rect -287 -519 -209 -473
rect -163 -519 -85 -473
rect -39 -519 39 -473
rect 85 -519 163 -473
rect 209 -519 287 -473
rect 333 -519 411 -473
rect 457 -519 535 -473
rect 581 -519 659 -473
rect 705 -519 783 -473
rect 829 -519 907 -473
rect 953 -519 1031 -473
rect 1077 -519 1088 -473
rect -1088 -597 1088 -519
rect -1088 -643 -1077 -597
rect -1031 -643 -953 -597
rect -907 -643 -829 -597
rect -783 -643 -705 -597
rect -659 -643 -581 -597
rect -535 -643 -457 -597
rect -411 -643 -333 -597
rect -287 -643 -209 -597
rect -163 -643 -85 -597
rect -39 -643 39 -597
rect 85 -643 163 -597
rect 209 -643 287 -597
rect 333 -643 411 -597
rect 457 -643 535 -597
rect 581 -643 659 -597
rect 705 -643 783 -597
rect 829 -643 907 -597
rect 953 -643 1031 -597
rect 1077 -643 1088 -597
rect -1088 -721 1088 -643
rect -1088 -767 -1077 -721
rect -1031 -767 -953 -721
rect -907 -767 -829 -721
rect -783 -767 -705 -721
rect -659 -767 -581 -721
rect -535 -767 -457 -721
rect -411 -767 -333 -721
rect -287 -767 -209 -721
rect -163 -767 -85 -721
rect -39 -767 39 -721
rect 85 -767 163 -721
rect 209 -767 287 -721
rect 333 -767 411 -721
rect 457 -767 535 -721
rect 581 -767 659 -721
rect 705 -767 783 -721
rect 829 -767 907 -721
rect 953 -767 1031 -721
rect 1077 -767 1088 -721
rect -1088 -845 1088 -767
rect -1088 -891 -1077 -845
rect -1031 -891 -953 -845
rect -907 -891 -829 -845
rect -783 -891 -705 -845
rect -659 -891 -581 -845
rect -535 -891 -457 -845
rect -411 -891 -333 -845
rect -287 -891 -209 -845
rect -163 -891 -85 -845
rect -39 -891 39 -845
rect 85 -891 163 -845
rect 209 -891 287 -845
rect 333 -891 411 -845
rect 457 -891 535 -845
rect 581 -891 659 -845
rect 705 -891 783 -845
rect 829 -891 907 -845
rect 953 -891 1031 -845
rect 1077 -891 1088 -845
rect -1088 -969 1088 -891
rect -1088 -1015 -1077 -969
rect -1031 -1015 -953 -969
rect -907 -1015 -829 -969
rect -783 -1015 -705 -969
rect -659 -1015 -581 -969
rect -535 -1015 -457 -969
rect -411 -1015 -333 -969
rect -287 -1015 -209 -969
rect -163 -1015 -85 -969
rect -39 -1015 39 -969
rect 85 -1015 163 -969
rect 209 -1015 287 -969
rect 333 -1015 411 -969
rect 457 -1015 535 -969
rect 581 -1015 659 -969
rect 705 -1015 783 -969
rect 829 -1015 907 -969
rect 953 -1015 1031 -969
rect 1077 -1015 1088 -969
rect -1088 -1093 1088 -1015
rect -1088 -1139 -1077 -1093
rect -1031 -1139 -953 -1093
rect -907 -1139 -829 -1093
rect -783 -1139 -705 -1093
rect -659 -1139 -581 -1093
rect -535 -1139 -457 -1093
rect -411 -1139 -333 -1093
rect -287 -1139 -209 -1093
rect -163 -1139 -85 -1093
rect -39 -1139 39 -1093
rect 85 -1139 163 -1093
rect 209 -1139 287 -1093
rect 333 -1139 411 -1093
rect 457 -1139 535 -1093
rect 581 -1139 659 -1093
rect 705 -1139 783 -1093
rect 829 -1139 907 -1093
rect 953 -1139 1031 -1093
rect 1077 -1139 1088 -1093
rect -1088 -1217 1088 -1139
rect -1088 -1263 -1077 -1217
rect -1031 -1263 -953 -1217
rect -907 -1263 -829 -1217
rect -783 -1263 -705 -1217
rect -659 -1263 -581 -1217
rect -535 -1263 -457 -1217
rect -411 -1263 -333 -1217
rect -287 -1263 -209 -1217
rect -163 -1263 -85 -1217
rect -39 -1263 39 -1217
rect 85 -1263 163 -1217
rect 209 -1263 287 -1217
rect 333 -1263 411 -1217
rect 457 -1263 535 -1217
rect 581 -1263 659 -1217
rect 705 -1263 783 -1217
rect 829 -1263 907 -1217
rect 953 -1263 1031 -1217
rect 1077 -1263 1088 -1217
rect -1088 -1341 1088 -1263
rect -1088 -1387 -1077 -1341
rect -1031 -1387 -953 -1341
rect -907 -1387 -829 -1341
rect -783 -1387 -705 -1341
rect -659 -1387 -581 -1341
rect -535 -1387 -457 -1341
rect -411 -1387 -333 -1341
rect -287 -1387 -209 -1341
rect -163 -1387 -85 -1341
rect -39 -1387 39 -1341
rect 85 -1387 163 -1341
rect 209 -1387 287 -1341
rect 333 -1387 411 -1341
rect 457 -1387 535 -1341
rect 581 -1387 659 -1341
rect 705 -1387 783 -1341
rect 829 -1387 907 -1341
rect 953 -1387 1031 -1341
rect 1077 -1387 1088 -1341
rect -1088 -1465 1088 -1387
rect -1088 -1511 -1077 -1465
rect -1031 -1511 -953 -1465
rect -907 -1511 -829 -1465
rect -783 -1511 -705 -1465
rect -659 -1511 -581 -1465
rect -535 -1511 -457 -1465
rect -411 -1511 -333 -1465
rect -287 -1511 -209 -1465
rect -163 -1511 -85 -1465
rect -39 -1511 39 -1465
rect 85 -1511 163 -1465
rect 209 -1511 287 -1465
rect 333 -1511 411 -1465
rect 457 -1511 535 -1465
rect 581 -1511 659 -1465
rect 705 -1511 783 -1465
rect 829 -1511 907 -1465
rect 953 -1511 1031 -1465
rect 1077 -1511 1088 -1465
rect -1088 -1589 1088 -1511
rect -1088 -1635 -1077 -1589
rect -1031 -1635 -953 -1589
rect -907 -1635 -829 -1589
rect -783 -1635 -705 -1589
rect -659 -1635 -581 -1589
rect -535 -1635 -457 -1589
rect -411 -1635 -333 -1589
rect -287 -1635 -209 -1589
rect -163 -1635 -85 -1589
rect -39 -1635 39 -1589
rect 85 -1635 163 -1589
rect 209 -1635 287 -1589
rect 333 -1635 411 -1589
rect 457 -1635 535 -1589
rect 581 -1635 659 -1589
rect 705 -1635 783 -1589
rect 829 -1635 907 -1589
rect 953 -1635 1031 -1589
rect 1077 -1635 1088 -1589
rect -1088 -1713 1088 -1635
rect -1088 -1759 -1077 -1713
rect -1031 -1759 -953 -1713
rect -907 -1759 -829 -1713
rect -783 -1759 -705 -1713
rect -659 -1759 -581 -1713
rect -535 -1759 -457 -1713
rect -411 -1759 -333 -1713
rect -287 -1759 -209 -1713
rect -163 -1759 -85 -1713
rect -39 -1759 39 -1713
rect 85 -1759 163 -1713
rect 209 -1759 287 -1713
rect 333 -1759 411 -1713
rect 457 -1759 535 -1713
rect 581 -1759 659 -1713
rect 705 -1759 783 -1713
rect 829 -1759 907 -1713
rect 953 -1759 1031 -1713
rect 1077 -1759 1088 -1713
rect -1088 -1837 1088 -1759
rect -1088 -1883 -1077 -1837
rect -1031 -1883 -953 -1837
rect -907 -1883 -829 -1837
rect -783 -1883 -705 -1837
rect -659 -1883 -581 -1837
rect -535 -1883 -457 -1837
rect -411 -1883 -333 -1837
rect -287 -1883 -209 -1837
rect -163 -1883 -85 -1837
rect -39 -1883 39 -1837
rect 85 -1883 163 -1837
rect 209 -1883 287 -1837
rect 333 -1883 411 -1837
rect 457 -1883 535 -1837
rect 581 -1883 659 -1837
rect 705 -1883 783 -1837
rect 829 -1883 907 -1837
rect 953 -1883 1031 -1837
rect 1077 -1883 1088 -1837
rect -1088 -1961 1088 -1883
rect -1088 -2007 -1077 -1961
rect -1031 -2007 -953 -1961
rect -907 -2007 -829 -1961
rect -783 -2007 -705 -1961
rect -659 -2007 -581 -1961
rect -535 -2007 -457 -1961
rect -411 -2007 -333 -1961
rect -287 -2007 -209 -1961
rect -163 -2007 -85 -1961
rect -39 -2007 39 -1961
rect 85 -2007 163 -1961
rect 209 -2007 287 -1961
rect 333 -2007 411 -1961
rect 457 -2007 535 -1961
rect 581 -2007 659 -1961
rect 705 -2007 783 -1961
rect 829 -2007 907 -1961
rect 953 -2007 1031 -1961
rect 1077 -2007 1088 -1961
rect -1088 -2085 1088 -2007
rect -1088 -2131 -1077 -2085
rect -1031 -2131 -953 -2085
rect -907 -2131 -829 -2085
rect -783 -2131 -705 -2085
rect -659 -2131 -581 -2085
rect -535 -2131 -457 -2085
rect -411 -2131 -333 -2085
rect -287 -2131 -209 -2085
rect -163 -2131 -85 -2085
rect -39 -2131 39 -2085
rect 85 -2131 163 -2085
rect 209 -2131 287 -2085
rect 333 -2131 411 -2085
rect 457 -2131 535 -2085
rect 581 -2131 659 -2085
rect 705 -2131 783 -2085
rect 829 -2131 907 -2085
rect 953 -2131 1031 -2085
rect 1077 -2131 1088 -2085
rect -1088 -2209 1088 -2131
rect -1088 -2255 -1077 -2209
rect -1031 -2255 -953 -2209
rect -907 -2255 -829 -2209
rect -783 -2255 -705 -2209
rect -659 -2255 -581 -2209
rect -535 -2255 -457 -2209
rect -411 -2255 -333 -2209
rect -287 -2255 -209 -2209
rect -163 -2255 -85 -2209
rect -39 -2255 39 -2209
rect 85 -2255 163 -2209
rect 209 -2255 287 -2209
rect 333 -2255 411 -2209
rect 457 -2255 535 -2209
rect 581 -2255 659 -2209
rect 705 -2255 783 -2209
rect 829 -2255 907 -2209
rect 953 -2255 1031 -2209
rect 1077 -2255 1088 -2209
rect -1088 -2333 1088 -2255
rect -1088 -2379 -1077 -2333
rect -1031 -2379 -953 -2333
rect -907 -2379 -829 -2333
rect -783 -2379 -705 -2333
rect -659 -2379 -581 -2333
rect -535 -2379 -457 -2333
rect -411 -2379 -333 -2333
rect -287 -2379 -209 -2333
rect -163 -2379 -85 -2333
rect -39 -2379 39 -2333
rect 85 -2379 163 -2333
rect 209 -2379 287 -2333
rect 333 -2379 411 -2333
rect 457 -2379 535 -2333
rect 581 -2379 659 -2333
rect 705 -2379 783 -2333
rect 829 -2379 907 -2333
rect 953 -2379 1031 -2333
rect 1077 -2379 1088 -2333
rect -1088 -2457 1088 -2379
rect -1088 -2503 -1077 -2457
rect -1031 -2503 -953 -2457
rect -907 -2503 -829 -2457
rect -783 -2503 -705 -2457
rect -659 -2503 -581 -2457
rect -535 -2503 -457 -2457
rect -411 -2503 -333 -2457
rect -287 -2503 -209 -2457
rect -163 -2503 -85 -2457
rect -39 -2503 39 -2457
rect 85 -2503 163 -2457
rect 209 -2503 287 -2457
rect 333 -2503 411 -2457
rect 457 -2503 535 -2457
rect 581 -2503 659 -2457
rect 705 -2503 783 -2457
rect 829 -2503 907 -2457
rect 953 -2503 1031 -2457
rect 1077 -2503 1088 -2457
rect -1088 -2581 1088 -2503
rect -1088 -2627 -1077 -2581
rect -1031 -2627 -953 -2581
rect -907 -2627 -829 -2581
rect -783 -2627 -705 -2581
rect -659 -2627 -581 -2581
rect -535 -2627 -457 -2581
rect -411 -2627 -333 -2581
rect -287 -2627 -209 -2581
rect -163 -2627 -85 -2581
rect -39 -2627 39 -2581
rect 85 -2627 163 -2581
rect 209 -2627 287 -2581
rect 333 -2627 411 -2581
rect 457 -2627 535 -2581
rect 581 -2627 659 -2581
rect 705 -2627 783 -2581
rect 829 -2627 907 -2581
rect 953 -2627 1031 -2581
rect 1077 -2627 1088 -2581
rect -1088 -2705 1088 -2627
rect -1088 -2751 -1077 -2705
rect -1031 -2751 -953 -2705
rect -907 -2751 -829 -2705
rect -783 -2751 -705 -2705
rect -659 -2751 -581 -2705
rect -535 -2751 -457 -2705
rect -411 -2751 -333 -2705
rect -287 -2751 -209 -2705
rect -163 -2751 -85 -2705
rect -39 -2751 39 -2705
rect 85 -2751 163 -2705
rect 209 -2751 287 -2705
rect 333 -2751 411 -2705
rect 457 -2751 535 -2705
rect 581 -2751 659 -2705
rect 705 -2751 783 -2705
rect 829 -2751 907 -2705
rect 953 -2751 1031 -2705
rect 1077 -2751 1088 -2705
rect -1088 -2829 1088 -2751
rect -1088 -2875 -1077 -2829
rect -1031 -2875 -953 -2829
rect -907 -2875 -829 -2829
rect -783 -2875 -705 -2829
rect -659 -2875 -581 -2829
rect -535 -2875 -457 -2829
rect -411 -2875 -333 -2829
rect -287 -2875 -209 -2829
rect -163 -2875 -85 -2829
rect -39 -2875 39 -2829
rect 85 -2875 163 -2829
rect 209 -2875 287 -2829
rect 333 -2875 411 -2829
rect 457 -2875 535 -2829
rect 581 -2875 659 -2829
rect 705 -2875 783 -2829
rect 829 -2875 907 -2829
rect 953 -2875 1031 -2829
rect 1077 -2875 1088 -2829
rect -1088 -2953 1088 -2875
rect -1088 -2999 -1077 -2953
rect -1031 -2999 -953 -2953
rect -907 -2999 -829 -2953
rect -783 -2999 -705 -2953
rect -659 -2999 -581 -2953
rect -535 -2999 -457 -2953
rect -411 -2999 -333 -2953
rect -287 -2999 -209 -2953
rect -163 -2999 -85 -2953
rect -39 -2999 39 -2953
rect 85 -2999 163 -2953
rect 209 -2999 287 -2953
rect 333 -2999 411 -2953
rect 457 -2999 535 -2953
rect 581 -2999 659 -2953
rect 705 -2999 783 -2953
rect 829 -2999 907 -2953
rect 953 -2999 1031 -2953
rect 1077 -2999 1088 -2953
rect -1088 -3077 1088 -2999
rect -1088 -3123 -1077 -3077
rect -1031 -3123 -953 -3077
rect -907 -3123 -829 -3077
rect -783 -3123 -705 -3077
rect -659 -3123 -581 -3077
rect -535 -3123 -457 -3077
rect -411 -3123 -333 -3077
rect -287 -3123 -209 -3077
rect -163 -3123 -85 -3077
rect -39 -3123 39 -3077
rect 85 -3123 163 -3077
rect 209 -3123 287 -3077
rect 333 -3123 411 -3077
rect 457 -3123 535 -3077
rect 581 -3123 659 -3077
rect 705 -3123 783 -3077
rect 829 -3123 907 -3077
rect 953 -3123 1031 -3077
rect 1077 -3123 1088 -3077
rect -1088 -3201 1088 -3123
rect -1088 -3247 -1077 -3201
rect -1031 -3247 -953 -3201
rect -907 -3247 -829 -3201
rect -783 -3247 -705 -3201
rect -659 -3247 -581 -3201
rect -535 -3247 -457 -3201
rect -411 -3247 -333 -3201
rect -287 -3247 -209 -3201
rect -163 -3247 -85 -3201
rect -39 -3247 39 -3201
rect 85 -3247 163 -3201
rect 209 -3247 287 -3201
rect 333 -3247 411 -3201
rect 457 -3247 535 -3201
rect 581 -3247 659 -3201
rect 705 -3247 783 -3201
rect 829 -3247 907 -3201
rect 953 -3247 1031 -3201
rect 1077 -3247 1088 -3201
rect -1088 -3325 1088 -3247
rect -1088 -3371 -1077 -3325
rect -1031 -3371 -953 -3325
rect -907 -3371 -829 -3325
rect -783 -3371 -705 -3325
rect -659 -3371 -581 -3325
rect -535 -3371 -457 -3325
rect -411 -3371 -333 -3325
rect -287 -3371 -209 -3325
rect -163 -3371 -85 -3325
rect -39 -3371 39 -3325
rect 85 -3371 163 -3325
rect 209 -3371 287 -3325
rect 333 -3371 411 -3325
rect 457 -3371 535 -3325
rect 581 -3371 659 -3325
rect 705 -3371 783 -3325
rect 829 -3371 907 -3325
rect 953 -3371 1031 -3325
rect 1077 -3371 1088 -3325
rect -1088 -3449 1088 -3371
rect -1088 -3495 -1077 -3449
rect -1031 -3495 -953 -3449
rect -907 -3495 -829 -3449
rect -783 -3495 -705 -3449
rect -659 -3495 -581 -3449
rect -535 -3495 -457 -3449
rect -411 -3495 -333 -3449
rect -287 -3495 -209 -3449
rect -163 -3495 -85 -3449
rect -39 -3495 39 -3449
rect 85 -3495 163 -3449
rect 209 -3495 287 -3449
rect 333 -3495 411 -3449
rect 457 -3495 535 -3449
rect 581 -3495 659 -3449
rect 705 -3495 783 -3449
rect 829 -3495 907 -3449
rect 953 -3495 1031 -3449
rect 1077 -3495 1088 -3449
rect -1088 -3573 1088 -3495
rect -1088 -3619 -1077 -3573
rect -1031 -3619 -953 -3573
rect -907 -3619 -829 -3573
rect -783 -3619 -705 -3573
rect -659 -3619 -581 -3573
rect -535 -3619 -457 -3573
rect -411 -3619 -333 -3573
rect -287 -3619 -209 -3573
rect -163 -3619 -85 -3573
rect -39 -3619 39 -3573
rect 85 -3619 163 -3573
rect 209 -3619 287 -3573
rect 333 -3619 411 -3573
rect 457 -3619 535 -3573
rect 581 -3619 659 -3573
rect 705 -3619 783 -3573
rect 829 -3619 907 -3573
rect 953 -3619 1031 -3573
rect 1077 -3619 1088 -3573
rect -1088 -3697 1088 -3619
rect -1088 -3743 -1077 -3697
rect -1031 -3743 -953 -3697
rect -907 -3743 -829 -3697
rect -783 -3743 -705 -3697
rect -659 -3743 -581 -3697
rect -535 -3743 -457 -3697
rect -411 -3743 -333 -3697
rect -287 -3743 -209 -3697
rect -163 -3743 -85 -3697
rect -39 -3743 39 -3697
rect 85 -3743 163 -3697
rect 209 -3743 287 -3697
rect 333 -3743 411 -3697
rect 457 -3743 535 -3697
rect 581 -3743 659 -3697
rect 705 -3743 783 -3697
rect 829 -3743 907 -3697
rect 953 -3743 1031 -3697
rect 1077 -3743 1088 -3697
rect -1088 -3821 1088 -3743
rect -1088 -3867 -1077 -3821
rect -1031 -3867 -953 -3821
rect -907 -3867 -829 -3821
rect -783 -3867 -705 -3821
rect -659 -3867 -581 -3821
rect -535 -3867 -457 -3821
rect -411 -3867 -333 -3821
rect -287 -3867 -209 -3821
rect -163 -3867 -85 -3821
rect -39 -3867 39 -3821
rect 85 -3867 163 -3821
rect 209 -3867 287 -3821
rect 333 -3867 411 -3821
rect 457 -3867 535 -3821
rect 581 -3867 659 -3821
rect 705 -3867 783 -3821
rect 829 -3867 907 -3821
rect 953 -3867 1031 -3821
rect 1077 -3867 1088 -3821
rect -1088 -3945 1088 -3867
rect -1088 -3991 -1077 -3945
rect -1031 -3991 -953 -3945
rect -907 -3991 -829 -3945
rect -783 -3991 -705 -3945
rect -659 -3991 -581 -3945
rect -535 -3991 -457 -3945
rect -411 -3991 -333 -3945
rect -287 -3991 -209 -3945
rect -163 -3991 -85 -3945
rect -39 -3991 39 -3945
rect 85 -3991 163 -3945
rect 209 -3991 287 -3945
rect 333 -3991 411 -3945
rect 457 -3991 535 -3945
rect 581 -3991 659 -3945
rect 705 -3991 783 -3945
rect 829 -3991 907 -3945
rect 953 -3991 1031 -3945
rect 1077 -3991 1088 -3945
rect -1088 -4069 1088 -3991
rect -1088 -4115 -1077 -4069
rect -1031 -4115 -953 -4069
rect -907 -4115 -829 -4069
rect -783 -4115 -705 -4069
rect -659 -4115 -581 -4069
rect -535 -4115 -457 -4069
rect -411 -4115 -333 -4069
rect -287 -4115 -209 -4069
rect -163 -4115 -85 -4069
rect -39 -4115 39 -4069
rect 85 -4115 163 -4069
rect 209 -4115 287 -4069
rect 333 -4115 411 -4069
rect 457 -4115 535 -4069
rect 581 -4115 659 -4069
rect 705 -4115 783 -4069
rect 829 -4115 907 -4069
rect 953 -4115 1031 -4069
rect 1077 -4115 1088 -4069
rect -1088 -4193 1088 -4115
rect -1088 -4239 -1077 -4193
rect -1031 -4239 -953 -4193
rect -907 -4239 -829 -4193
rect -783 -4239 -705 -4193
rect -659 -4239 -581 -4193
rect -535 -4239 -457 -4193
rect -411 -4239 -333 -4193
rect -287 -4239 -209 -4193
rect -163 -4239 -85 -4193
rect -39 -4239 39 -4193
rect 85 -4239 163 -4193
rect 209 -4239 287 -4193
rect 333 -4239 411 -4193
rect 457 -4239 535 -4193
rect 581 -4239 659 -4193
rect 705 -4239 783 -4193
rect 829 -4239 907 -4193
rect 953 -4239 1031 -4193
rect 1077 -4239 1088 -4193
rect -1088 -4317 1088 -4239
rect -1088 -4363 -1077 -4317
rect -1031 -4363 -953 -4317
rect -907 -4363 -829 -4317
rect -783 -4363 -705 -4317
rect -659 -4363 -581 -4317
rect -535 -4363 -457 -4317
rect -411 -4363 -333 -4317
rect -287 -4363 -209 -4317
rect -163 -4363 -85 -4317
rect -39 -4363 39 -4317
rect 85 -4363 163 -4317
rect 209 -4363 287 -4317
rect 333 -4363 411 -4317
rect 457 -4363 535 -4317
rect 581 -4363 659 -4317
rect 705 -4363 783 -4317
rect 829 -4363 907 -4317
rect 953 -4363 1031 -4317
rect 1077 -4363 1088 -4317
rect -1088 -4441 1088 -4363
rect -1088 -4487 -1077 -4441
rect -1031 -4487 -953 -4441
rect -907 -4487 -829 -4441
rect -783 -4487 -705 -4441
rect -659 -4487 -581 -4441
rect -535 -4487 -457 -4441
rect -411 -4487 -333 -4441
rect -287 -4487 -209 -4441
rect -163 -4487 -85 -4441
rect -39 -4487 39 -4441
rect 85 -4487 163 -4441
rect 209 -4487 287 -4441
rect 333 -4487 411 -4441
rect 457 -4487 535 -4441
rect 581 -4487 659 -4441
rect 705 -4487 783 -4441
rect 829 -4487 907 -4441
rect 953 -4487 1031 -4441
rect 1077 -4487 1088 -4441
rect -1088 -4565 1088 -4487
rect -1088 -4611 -1077 -4565
rect -1031 -4611 -953 -4565
rect -907 -4611 -829 -4565
rect -783 -4611 -705 -4565
rect -659 -4611 -581 -4565
rect -535 -4611 -457 -4565
rect -411 -4611 -333 -4565
rect -287 -4611 -209 -4565
rect -163 -4611 -85 -4565
rect -39 -4611 39 -4565
rect 85 -4611 163 -4565
rect 209 -4611 287 -4565
rect 333 -4611 411 -4565
rect 457 -4611 535 -4565
rect 581 -4611 659 -4565
rect 705 -4611 783 -4565
rect 829 -4611 907 -4565
rect 953 -4611 1031 -4565
rect 1077 -4611 1088 -4565
rect -1088 -4689 1088 -4611
rect -1088 -4735 -1077 -4689
rect -1031 -4735 -953 -4689
rect -907 -4735 -829 -4689
rect -783 -4735 -705 -4689
rect -659 -4735 -581 -4689
rect -535 -4735 -457 -4689
rect -411 -4735 -333 -4689
rect -287 -4735 -209 -4689
rect -163 -4735 -85 -4689
rect -39 -4735 39 -4689
rect 85 -4735 163 -4689
rect 209 -4735 287 -4689
rect 333 -4735 411 -4689
rect 457 -4735 535 -4689
rect 581 -4735 659 -4689
rect 705 -4735 783 -4689
rect 829 -4735 907 -4689
rect 953 -4735 1031 -4689
rect 1077 -4735 1088 -4689
rect -1088 -4813 1088 -4735
rect -1088 -4859 -1077 -4813
rect -1031 -4859 -953 -4813
rect -907 -4859 -829 -4813
rect -783 -4859 -705 -4813
rect -659 -4859 -581 -4813
rect -535 -4859 -457 -4813
rect -411 -4859 -333 -4813
rect -287 -4859 -209 -4813
rect -163 -4859 -85 -4813
rect -39 -4859 39 -4813
rect 85 -4859 163 -4813
rect 209 -4859 287 -4813
rect 333 -4859 411 -4813
rect 457 -4859 535 -4813
rect 581 -4859 659 -4813
rect 705 -4859 783 -4813
rect 829 -4859 907 -4813
rect 953 -4859 1031 -4813
rect 1077 -4859 1088 -4813
rect -1088 -4937 1088 -4859
rect -1088 -4983 -1077 -4937
rect -1031 -4983 -953 -4937
rect -907 -4983 -829 -4937
rect -783 -4983 -705 -4937
rect -659 -4983 -581 -4937
rect -535 -4983 -457 -4937
rect -411 -4983 -333 -4937
rect -287 -4983 -209 -4937
rect -163 -4983 -85 -4937
rect -39 -4983 39 -4937
rect 85 -4983 163 -4937
rect 209 -4983 287 -4937
rect 333 -4983 411 -4937
rect 457 -4983 535 -4937
rect 581 -4983 659 -4937
rect 705 -4983 783 -4937
rect 829 -4983 907 -4937
rect 953 -4983 1031 -4937
rect 1077 -4983 1088 -4937
rect -1088 -5061 1088 -4983
rect -1088 -5107 -1077 -5061
rect -1031 -5107 -953 -5061
rect -907 -5107 -829 -5061
rect -783 -5107 -705 -5061
rect -659 -5107 -581 -5061
rect -535 -5107 -457 -5061
rect -411 -5107 -333 -5061
rect -287 -5107 -209 -5061
rect -163 -5107 -85 -5061
rect -39 -5107 39 -5061
rect 85 -5107 163 -5061
rect 209 -5107 287 -5061
rect 333 -5107 411 -5061
rect 457 -5107 535 -5061
rect 581 -5107 659 -5061
rect 705 -5107 783 -5061
rect 829 -5107 907 -5061
rect 953 -5107 1031 -5061
rect 1077 -5107 1088 -5061
rect -1088 -5185 1088 -5107
rect -1088 -5231 -1077 -5185
rect -1031 -5231 -953 -5185
rect -907 -5231 -829 -5185
rect -783 -5231 -705 -5185
rect -659 -5231 -581 -5185
rect -535 -5231 -457 -5185
rect -411 -5231 -333 -5185
rect -287 -5231 -209 -5185
rect -163 -5231 -85 -5185
rect -39 -5231 39 -5185
rect 85 -5231 163 -5185
rect 209 -5231 287 -5185
rect 333 -5231 411 -5185
rect 457 -5231 535 -5185
rect 581 -5231 659 -5185
rect 705 -5231 783 -5185
rect 829 -5231 907 -5185
rect 953 -5231 1031 -5185
rect 1077 -5231 1088 -5185
rect -1088 -5309 1088 -5231
rect -1088 -5355 -1077 -5309
rect -1031 -5355 -953 -5309
rect -907 -5355 -829 -5309
rect -783 -5355 -705 -5309
rect -659 -5355 -581 -5309
rect -535 -5355 -457 -5309
rect -411 -5355 -333 -5309
rect -287 -5355 -209 -5309
rect -163 -5355 -85 -5309
rect -39 -5355 39 -5309
rect 85 -5355 163 -5309
rect 209 -5355 287 -5309
rect 333 -5355 411 -5309
rect 457 -5355 535 -5309
rect 581 -5355 659 -5309
rect 705 -5355 783 -5309
rect 829 -5355 907 -5309
rect 953 -5355 1031 -5309
rect 1077 -5355 1088 -5309
rect -1088 -5433 1088 -5355
rect -1088 -5479 -1077 -5433
rect -1031 -5479 -953 -5433
rect -907 -5479 -829 -5433
rect -783 -5479 -705 -5433
rect -659 -5479 -581 -5433
rect -535 -5479 -457 -5433
rect -411 -5479 -333 -5433
rect -287 -5479 -209 -5433
rect -163 -5479 -85 -5433
rect -39 -5479 39 -5433
rect 85 -5479 163 -5433
rect 209 -5479 287 -5433
rect 333 -5479 411 -5433
rect 457 -5479 535 -5433
rect 581 -5479 659 -5433
rect 705 -5479 783 -5433
rect 829 -5479 907 -5433
rect 953 -5479 1031 -5433
rect 1077 -5479 1088 -5433
rect -1088 -5557 1088 -5479
rect -1088 -5603 -1077 -5557
rect -1031 -5603 -953 -5557
rect -907 -5603 -829 -5557
rect -783 -5603 -705 -5557
rect -659 -5603 -581 -5557
rect -535 -5603 -457 -5557
rect -411 -5603 -333 -5557
rect -287 -5603 -209 -5557
rect -163 -5603 -85 -5557
rect -39 -5603 39 -5557
rect 85 -5603 163 -5557
rect 209 -5603 287 -5557
rect 333 -5603 411 -5557
rect 457 -5603 535 -5557
rect 581 -5603 659 -5557
rect 705 -5603 783 -5557
rect 829 -5603 907 -5557
rect 953 -5603 1031 -5557
rect 1077 -5603 1088 -5557
rect -1088 -5681 1088 -5603
rect -1088 -5727 -1077 -5681
rect -1031 -5727 -953 -5681
rect -907 -5727 -829 -5681
rect -783 -5727 -705 -5681
rect -659 -5727 -581 -5681
rect -535 -5727 -457 -5681
rect -411 -5727 -333 -5681
rect -287 -5727 -209 -5681
rect -163 -5727 -85 -5681
rect -39 -5727 39 -5681
rect 85 -5727 163 -5681
rect 209 -5727 287 -5681
rect 333 -5727 411 -5681
rect 457 -5727 535 -5681
rect 581 -5727 659 -5681
rect 705 -5727 783 -5681
rect 829 -5727 907 -5681
rect 953 -5727 1031 -5681
rect 1077 -5727 1088 -5681
rect -1088 -5805 1088 -5727
rect -1088 -5851 -1077 -5805
rect -1031 -5851 -953 -5805
rect -907 -5851 -829 -5805
rect -783 -5851 -705 -5805
rect -659 -5851 -581 -5805
rect -535 -5851 -457 -5805
rect -411 -5851 -333 -5805
rect -287 -5851 -209 -5805
rect -163 -5851 -85 -5805
rect -39 -5851 39 -5805
rect 85 -5851 163 -5805
rect 209 -5851 287 -5805
rect 333 -5851 411 -5805
rect 457 -5851 535 -5805
rect 581 -5851 659 -5805
rect 705 -5851 783 -5805
rect 829 -5851 907 -5805
rect 953 -5851 1031 -5805
rect 1077 -5851 1088 -5805
rect -1088 -5862 1088 -5851
<< end >>
