magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1247 -1133 1247 1133
<< metal2 >>
rect -247 128 247 133
rect -247 100 -242 128
rect -214 100 -166 128
rect -138 100 -90 128
rect -62 100 -14 128
rect 14 100 62 128
rect 90 100 138 128
rect 166 100 214 128
rect 242 100 247 128
rect -247 52 247 100
rect -247 24 -242 52
rect -214 24 -166 52
rect -138 24 -90 52
rect -62 24 -14 52
rect 14 24 62 52
rect 90 24 138 52
rect 166 24 214 52
rect 242 24 247 52
rect -247 -24 247 24
rect -247 -52 -242 -24
rect -214 -52 -166 -24
rect -138 -52 -90 -24
rect -62 -52 -14 -24
rect 14 -52 62 -24
rect 90 -52 138 -24
rect 166 -52 214 -24
rect 242 -52 247 -24
rect -247 -100 247 -52
rect -247 -128 -242 -100
rect -214 -128 -166 -100
rect -138 -128 -90 -100
rect -62 -128 -14 -100
rect 14 -128 62 -100
rect 90 -128 138 -100
rect 166 -128 214 -100
rect 242 -128 247 -100
rect -247 -133 247 -128
<< via2 >>
rect -242 100 -214 128
rect -166 100 -138 128
rect -90 100 -62 128
rect -14 100 14 128
rect 62 100 90 128
rect 138 100 166 128
rect 214 100 242 128
rect -242 24 -214 52
rect -166 24 -138 52
rect -90 24 -62 52
rect -14 24 14 52
rect 62 24 90 52
rect 138 24 166 52
rect 214 24 242 52
rect -242 -52 -214 -24
rect -166 -52 -138 -24
rect -90 -52 -62 -24
rect -14 -52 14 -24
rect 62 -52 90 -24
rect 138 -52 166 -24
rect 214 -52 242 -24
rect -242 -128 -214 -100
rect -166 -128 -138 -100
rect -90 -128 -62 -100
rect -14 -128 14 -100
rect 62 -128 90 -100
rect 138 -128 166 -100
rect 214 -128 242 -100
<< metal3 >>
rect -247 128 247 133
rect -247 100 -242 128
rect -214 100 -166 128
rect -138 100 -90 128
rect -62 100 -14 128
rect 14 100 62 128
rect 90 100 138 128
rect 166 100 214 128
rect 242 100 247 128
rect -247 52 247 100
rect -247 24 -242 52
rect -214 24 -166 52
rect -138 24 -90 52
rect -62 24 -14 52
rect 14 24 62 52
rect 90 24 138 52
rect 166 24 214 52
rect 242 24 247 52
rect -247 -24 247 24
rect -247 -52 -242 -24
rect -214 -52 -166 -24
rect -138 -52 -90 -24
rect -62 -52 -14 -24
rect 14 -52 62 -24
rect 90 -52 138 -24
rect 166 -52 214 -24
rect 242 -52 247 -24
rect -247 -100 247 -52
rect -247 -128 -242 -100
rect -214 -128 -166 -100
rect -138 -128 -90 -100
rect -62 -128 -14 -100
rect 14 -128 62 -100
rect 90 -128 138 -100
rect 166 -128 214 -100
rect 242 -128 247 -100
rect -247 -133 247 -128
<< end >>
