magic
tech gf180mcuC
magscale 1 10
timestamp 1694427317
<< psubdiff >>
rect -280 1977 3975 1994
rect -280 1911 -167 1977
rect -79 1911 -17 1977
rect 71 1911 133 1977
rect 221 1911 283 1977
rect 371 1911 433 1977
rect 521 1911 583 1977
rect 671 1911 733 1977
rect 821 1911 883 1977
rect 971 1911 1033 1977
rect 1121 1911 1183 1977
rect 1271 1911 1333 1977
rect 1421 1911 1483 1977
rect 1571 1911 1633 1977
rect 1721 1911 1783 1977
rect 1871 1911 1933 1977
rect 2021 1911 2083 1977
rect 2171 1911 2233 1977
rect 2321 1911 2383 1977
rect 2471 1911 2533 1977
rect 2621 1911 2683 1977
rect 2771 1911 2833 1977
rect 2921 1911 2983 1977
rect 3071 1911 3133 1977
rect 3221 1911 3283 1977
rect 3371 1911 3433 1977
rect 3521 1911 3583 1977
rect 3671 1911 3733 1977
rect 3821 1911 3975 1977
rect -280 1884 3975 1911
rect -280 1855 -170 1884
rect -280 1767 -258 1855
rect -191 1767 -170 1855
rect -280 1705 -170 1767
rect -280 1617 -258 1705
rect -191 1617 -170 1705
rect -280 1555 -170 1617
rect -280 1467 -258 1555
rect -191 1467 -170 1555
rect -280 1405 -170 1467
rect -280 1317 -258 1405
rect -191 1317 -170 1405
rect -280 1255 -170 1317
rect -280 1167 -258 1255
rect -191 1167 -170 1255
rect -280 1105 -170 1167
rect -280 1017 -258 1105
rect -191 1017 -170 1105
rect -280 955 -170 1017
rect -280 867 -258 955
rect -191 867 -170 955
rect -280 805 -170 867
rect -280 717 -258 805
rect -191 717 -170 805
rect -280 655 -170 717
rect -280 567 -258 655
rect -191 567 -170 655
rect -280 505 -170 567
rect -280 417 -258 505
rect -191 417 -170 505
rect -280 355 -170 417
rect -280 267 -258 355
rect -191 267 -170 355
rect -280 205 -170 267
rect -280 117 -258 205
rect -191 117 -170 205
rect -280 55 -170 117
rect -280 -33 -258 55
rect -191 -33 -170 55
rect -280 -79 -170 -33
rect 3865 1815 3975 1884
rect 3865 1727 3884 1815
rect 3951 1727 3975 1815
rect 3865 1665 3975 1727
rect 3865 1577 3884 1665
rect 3951 1577 3975 1665
rect 3865 1515 3975 1577
rect 3865 1427 3884 1515
rect 3951 1427 3975 1515
rect 3865 1365 3975 1427
rect 3865 1277 3884 1365
rect 3951 1277 3975 1365
rect 3865 1215 3975 1277
rect 3865 1127 3884 1215
rect 3951 1127 3975 1215
rect 3865 1065 3975 1127
rect 3865 977 3884 1065
rect 3951 977 3975 1065
rect 3865 915 3975 977
rect 3865 827 3884 915
rect 3951 827 3975 915
rect 3865 765 3975 827
rect 3865 677 3884 765
rect 3951 677 3975 765
rect 3865 615 3975 677
rect 3865 527 3884 615
rect 3951 527 3975 615
rect 3865 465 3975 527
rect 3865 377 3884 465
rect 3951 377 3975 465
rect 3865 315 3975 377
rect 3865 227 3884 315
rect 3951 227 3975 315
rect 3865 165 3975 227
rect 3865 77 3884 165
rect 3951 77 3975 165
rect 3865 15 3975 77
rect 3865 -73 3884 15
rect 3951 -73 3975 15
rect 3865 -79 3975 -73
rect -280 -102 3975 -79
rect -280 -168 -150 -102
rect -62 -168 0 -102
rect 88 -168 150 -102
rect 238 -168 300 -102
rect 388 -168 450 -102
rect 538 -168 600 -102
rect 688 -168 750 -102
rect 838 -168 900 -102
rect 988 -168 1050 -102
rect 1138 -168 1200 -102
rect 1288 -168 1350 -102
rect 1438 -168 1500 -102
rect 1588 -168 1650 -102
rect 1738 -168 1800 -102
rect 1888 -168 1950 -102
rect 2038 -168 2100 -102
rect 2188 -168 2250 -102
rect 2338 -168 2400 -102
rect 2488 -168 2550 -102
rect 2638 -168 2700 -102
rect 2788 -168 2850 -102
rect 2938 -168 3000 -102
rect 3088 -168 3150 -102
rect 3238 -168 3300 -102
rect 3388 -168 3450 -102
rect 3538 -168 3600 -102
rect 3688 -168 3750 -102
rect 3838 -168 3975 -102
rect -280 -189 3975 -168
<< psubdiffcont >>
rect -167 1911 -79 1977
rect -17 1911 71 1977
rect 133 1911 221 1977
rect 283 1911 371 1977
rect 433 1911 521 1977
rect 583 1911 671 1977
rect 733 1911 821 1977
rect 883 1911 971 1977
rect 1033 1911 1121 1977
rect 1183 1911 1271 1977
rect 1333 1911 1421 1977
rect 1483 1911 1571 1977
rect 1633 1911 1721 1977
rect 1783 1911 1871 1977
rect 1933 1911 2021 1977
rect 2083 1911 2171 1977
rect 2233 1911 2321 1977
rect 2383 1911 2471 1977
rect 2533 1911 2621 1977
rect 2683 1911 2771 1977
rect 2833 1911 2921 1977
rect 2983 1911 3071 1977
rect 3133 1911 3221 1977
rect 3283 1911 3371 1977
rect 3433 1911 3521 1977
rect 3583 1911 3671 1977
rect 3733 1911 3821 1977
rect -258 1767 -191 1855
rect -258 1617 -191 1705
rect -258 1467 -191 1555
rect -258 1317 -191 1405
rect -258 1167 -191 1255
rect -258 1017 -191 1105
rect -258 867 -191 955
rect -258 717 -191 805
rect -258 567 -191 655
rect -258 417 -191 505
rect -258 267 -191 355
rect -258 117 -191 205
rect -258 -33 -191 55
rect 3884 1727 3951 1815
rect 3884 1577 3951 1665
rect 3884 1427 3951 1515
rect 3884 1277 3951 1365
rect 3884 1127 3951 1215
rect 3884 977 3951 1065
rect 3884 827 3951 915
rect 3884 677 3951 765
rect 3884 527 3951 615
rect 3884 377 3951 465
rect 3884 227 3951 315
rect 3884 77 3951 165
rect 3884 -73 3951 15
rect -150 -168 -62 -102
rect 0 -168 88 -102
rect 150 -168 238 -102
rect 300 -168 388 -102
rect 450 -168 538 -102
rect 600 -168 688 -102
rect 750 -168 838 -102
rect 900 -168 988 -102
rect 1050 -168 1138 -102
rect 1200 -168 1288 -102
rect 1350 -168 1438 -102
rect 1500 -168 1588 -102
rect 1650 -168 1738 -102
rect 1800 -168 1888 -102
rect 1950 -168 2038 -102
rect 2100 -168 2188 -102
rect 2250 -168 2338 -102
rect 2400 -168 2488 -102
rect 2550 -168 2638 -102
rect 2700 -168 2788 -102
rect 2850 -168 2938 -102
rect 3000 -168 3088 -102
rect 3150 -168 3238 -102
rect 3300 -168 3388 -102
rect 3450 -168 3538 -102
rect 3600 -168 3688 -102
rect 3750 -168 3838 -102
<< metal1 >>
rect 1789 2209 1905 2227
rect 1686 2112 1799 2209
rect 1896 2112 1905 2209
rect 1789 2098 1905 2112
rect -285 1977 3979 1999
rect -285 1911 -167 1977
rect -79 1911 -17 1977
rect 71 1911 133 1977
rect 221 1911 283 1977
rect 371 1911 433 1977
rect 521 1911 583 1977
rect 671 1911 733 1977
rect 821 1911 883 1977
rect 971 1911 1033 1977
rect 1121 1911 1183 1977
rect 1271 1911 1333 1977
rect 1421 1911 1483 1977
rect 1571 1911 1633 1977
rect 1721 1911 1783 1977
rect 1871 1911 1933 1977
rect 2021 1911 2083 1977
rect 2171 1911 2233 1977
rect 2321 1911 2383 1977
rect 2471 1911 2533 1977
rect 2621 1911 2683 1977
rect 2771 1911 2833 1977
rect 2921 1911 2983 1977
rect 3071 1911 3133 1977
rect 3221 1911 3283 1977
rect 3371 1911 3433 1977
rect 3521 1911 3583 1977
rect 3671 1911 3733 1977
rect 3821 1911 3979 1977
rect -285 1879 3979 1911
rect -285 1855 -165 1879
rect -285 1767 -258 1855
rect -191 1767 -165 1855
rect 3859 1815 3979 1879
rect -285 1705 -165 1767
rect 1076 1708 2587 1786
rect 3859 1727 3884 1815
rect 3951 1727 3979 1815
rect -285 1617 -258 1705
rect -191 1617 -165 1705
rect -285 1555 -165 1617
rect -285 1467 -258 1555
rect -191 1467 -165 1555
rect -285 1405 -165 1467
rect -285 1317 -258 1405
rect -191 1317 -165 1405
rect -285 1255 -165 1317
rect -285 1167 -258 1255
rect -191 1167 -165 1255
rect -285 1105 -165 1167
rect -285 1017 -258 1105
rect -191 1017 -165 1105
rect -285 955 -165 1017
rect -82 1201 28 1217
rect -82 1139 -65 1201
rect -3 1139 28 1201
rect -82 1084 28 1139
rect 1374 1112 1452 1708
rect 1613 1106 1691 1708
rect 1852 1099 1930 1708
rect 2078 1108 2156 1708
rect 3859 1665 3979 1727
rect 3859 1577 3884 1665
rect 3951 1577 3979 1665
rect 3859 1515 3979 1577
rect 3859 1427 3884 1515
rect 3951 1427 3979 1515
rect 3691 1360 3810 1399
rect 3691 1265 3705 1360
rect 3800 1265 3810 1360
rect 3691 1190 3810 1265
rect 3692 1175 3810 1190
rect -82 1044 67 1084
rect 3692 1080 3703 1175
rect 3798 1080 3810 1175
rect 3648 1076 3810 1080
rect 3859 1365 3979 1427
rect 3859 1277 3884 1365
rect 3951 1277 3979 1365
rect 3859 1215 3979 1277
rect 3859 1127 3884 1215
rect 3951 1127 3979 1215
rect -82 982 -72 1044
rect -10 982 120 1044
rect 3648 983 3799 1076
rect 3859 1065 3979 1127
rect -82 971 67 982
rect 3859 977 3884 1065
rect 3951 977 3979 1065
rect -285 867 -258 955
rect -191 867 -165 955
rect -285 805 -165 867
rect -285 717 -258 805
rect -191 717 -165 805
rect -285 655 -165 717
rect -285 567 -258 655
rect -191 567 -165 655
rect 3859 915 3979 977
rect 3859 827 3884 915
rect 3951 827 3979 915
rect 3859 765 3979 827
rect 3859 677 3884 765
rect 3951 677 3979 765
rect 3859 615 3979 677
rect -285 505 -165 567
rect -285 417 -258 505
rect -191 417 -165 505
rect -285 355 -165 417
rect -285 267 -258 355
rect -191 267 -165 355
rect -3 529 98 543
rect 235 529 307 609
rect -3 528 307 529
rect -3 458 12 528
rect 82 458 307 528
rect 3735 524 3795 533
rect 3859 527 3884 615
rect 3951 527 3979 615
rect 3458 523 3736 524
rect -3 457 307 458
rect -3 373 98 457
rect -3 301 11 373
rect 83 301 98 373
rect 235 358 307 457
rect 1134 459 1232 512
rect 2385 488 2551 503
rect 1134 427 1453 459
rect 2336 442 2551 488
rect 3458 467 3619 523
rect 3675 467 3736 523
rect 3458 466 3736 467
rect 3794 466 3804 524
rect 3735 457 3804 466
rect 2385 430 2551 442
rect -3 296 98 301
rect 1134 353 1147 427
rect 1221 387 1453 427
rect 1221 353 1232 387
rect -285 205 -165 267
rect -285 117 -258 205
rect -191 117 -165 205
rect 1134 259 1232 353
rect 3746 367 3804 457
rect 3746 311 3747 367
rect 3803 311 3804 367
rect 3746 297 3804 311
rect 3859 465 3979 527
rect 3859 377 3884 465
rect 3951 377 3979 465
rect 3859 315 3979 377
rect 1134 183 1146 259
rect 1222 183 1232 259
rect 1134 174 1232 183
rect 3859 227 3884 315
rect 3951 227 3979 315
rect -285 55 -165 117
rect 3859 165 3979 227
rect -285 -33 -258 55
rect -191 -33 -165 55
rect -285 -73 -165 -33
rect -285 -74 46 -73
rect 197 -74 304 107
rect 681 -74 786 105
rect 1054 3 2632 91
rect 1657 -74 1747 3
rect 2451 -74 2539 3
rect 2926 -74 3031 107
rect 3859 77 3884 165
rect 3951 77 3979 165
rect 3859 15 3979 77
rect 3859 -73 3884 15
rect 3951 -73 3979 15
rect 3859 -74 3979 -73
rect -285 -102 3979 -74
rect -285 -168 -150 -102
rect -62 -168 0 -102
rect 88 -168 150 -102
rect 238 -168 300 -102
rect 388 -168 450 -102
rect 538 -168 600 -102
rect 688 -168 750 -102
rect 838 -168 900 -102
rect 988 -168 1050 -102
rect 1138 -168 1200 -102
rect 1288 -168 1350 -102
rect 1438 -168 1500 -102
rect 1588 -168 1650 -102
rect 1738 -168 1800 -102
rect 1888 -168 1950 -102
rect 2038 -168 2100 -102
rect 2188 -168 2250 -102
rect 2338 -168 2400 -102
rect 2488 -168 2550 -102
rect 2638 -168 2700 -102
rect 2788 -168 2850 -102
rect 2938 -168 3000 -102
rect 3088 -168 3150 -102
rect 3238 -168 3300 -102
rect 3388 -168 3450 -102
rect 3538 -168 3600 -102
rect 3688 -168 3750 -102
rect 3838 -168 3979 -102
rect -285 -193 3979 -168
rect -17 -314 392 -297
rect -17 -315 146 -314
rect -17 -387 11 -315
rect 83 -386 146 -315
rect 218 -316 392 -314
rect 218 -386 272 -316
rect 342 -386 392 -316
rect 83 -387 392 -386
rect -17 -403 392 -387
rect 794 -302 972 -301
rect 794 -314 1248 -302
rect 794 -315 995 -314
rect 794 -389 855 -315
rect 929 -389 995 -315
rect 794 -390 995 -389
rect 1071 -390 1146 -314
rect 1222 -390 1248 -314
rect 794 -410 1248 -390
rect 3327 -347 3845 -327
rect 3327 -349 3549 -347
rect 794 -413 972 -410
rect 3327 -438 3401 -349
rect 3490 -438 3549 -349
rect 3640 -349 3845 -347
rect 3640 -438 3731 -349
rect 3327 -440 3731 -438
rect 3822 -440 3845 -349
rect 3327 -452 3845 -440
<< via1 >>
rect 1799 2112 1896 2209
rect -65 1139 -3 1201
rect 3705 1265 3800 1360
rect 3703 1080 3798 1175
rect -72 982 -10 1044
rect 12 458 82 528
rect 11 301 83 373
rect 3619 467 3675 523
rect 3736 466 3794 524
rect 1147 353 1221 427
rect 3747 311 3803 367
rect 1146 183 1222 259
rect 11 -387 83 -315
rect 146 -386 218 -314
rect 272 -386 342 -316
rect 855 -389 929 -315
rect 995 -390 1071 -314
rect 1146 -390 1222 -314
rect 3401 -438 3490 -349
rect 3549 -438 3640 -347
rect 3731 -440 3822 -349
<< metal2 >>
rect 1789 2209 1905 2227
rect 1789 2112 1799 2209
rect 1896 2112 1905 2209
rect 1789 2098 1905 2112
rect 1799 1868 1896 2098
rect -73 1771 3799 1868
rect -69 1217 28 1771
rect 3702 1399 3799 1771
rect -82 1201 28 1217
rect -82 1139 -65 1201
rect -3 1139 28 1201
rect 3691 1360 3810 1399
rect 3691 1265 3705 1360
rect 3800 1265 3810 1360
rect 3691 1190 3810 1265
rect -82 1084 28 1139
rect 3692 1175 3810 1190
rect 3692 1099 3703 1175
rect -82 1044 67 1084
rect 3659 1080 3703 1099
rect 3798 1080 3810 1175
rect 3659 1076 3810 1080
rect -82 982 -72 1044
rect -10 982 78 1044
rect -82 971 67 982
rect 3659 969 3809 1076
rect -3 528 98 543
rect -3 458 12 528
rect 82 458 98 528
rect 3613 524 3816 539
rect 3613 523 3736 524
rect -3 373 98 458
rect -3 301 11 373
rect 83 301 98 373
rect -3 296 98 301
rect 1134 427 1232 512
rect 3613 467 3619 523
rect 3675 467 3736 523
rect 3613 466 3736 467
rect 3794 466 3816 524
rect 3613 455 3816 466
rect 1134 353 1147 427
rect 1221 353 1232 427
rect 3736 384 3816 455
rect 11 -297 83 296
rect 1134 259 1232 353
rect 1134 183 1146 259
rect 1222 183 1232 259
rect 1134 174 1232 183
rect 3731 367 3822 384
rect 3731 311 3747 367
rect 3803 311 3822 367
rect -17 -314 369 -297
rect 1146 -302 1222 174
rect -17 -315 146 -314
rect -17 -387 11 -315
rect 83 -386 146 -315
rect 218 -316 369 -314
rect 218 -386 272 -316
rect 342 -386 369 -316
rect 83 -387 369 -386
rect -17 -403 369 -387
rect 826 -314 1248 -302
rect 826 -315 995 -314
rect 826 -389 855 -315
rect 929 -389 995 -315
rect 826 -390 995 -389
rect 1071 -390 1146 -314
rect 1222 -390 1248 -314
rect 3731 -327 3822 311
rect 826 -410 1248 -390
rect 3378 -347 3845 -327
rect 3378 -349 3549 -347
rect 3378 -438 3401 -349
rect 3490 -438 3549 -349
rect 3640 -349 3845 -347
rect 3640 -438 3731 -349
rect 3378 -440 3731 -438
rect 3822 -440 3845 -349
rect 3378 -452 3845 -440
use INV_2  INV_2_0 ~/GF180Projects/Layout/Magic/VCO1/INV_2
timestamp 1693141036
transform 1 0 1311 0 1 486
box 21 -485 1081 648
use Tr_Gate  Tr_Gate_0 ~/GF180Projects/Layout/Magic/VCO1/Tr_Gate
timestamp 1692985371
transform -1 0 1154 0 1 1233
box -53 -1233 1187 569
use Tr_Gate  Tr_Gate_1
timestamp 1692985371
transform 1 0 2558 0 1 1235
box -53 -1233 1187 569
<< labels >>
flabel metal1 811 -359 811 -359 0 FreeSans 800 0 0 0 SEL
port 0 nsew
flabel metal1 3355 -397 3355 -397 0 FreeSans 800 0 0 0 IN1
port 1 nsew
flabel metal1 377 -354 377 -354 0 FreeSans 800 0 0 0 IN2
port 2 nsew
flabel metal1 1705 1747 1705 1747 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal1 1288 27 1288 27 0 FreeSans 800 0 0 0 VSS
port 4 nsew
flabel metal1 1728 2158 1728 2158 0 FreeSans 800 0 0 0 OUT
port 5 nsew
<< end >>
