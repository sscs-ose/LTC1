magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3690 -2045 3690 2045
<< psubdiff >>
rect -1690 23 1690 45
rect -1690 -23 -1668 23
rect 1668 -23 1690 23
rect -1690 -45 1690 -23
<< psubdiffcont >>
rect -1668 -23 1668 23
<< metal1 >>
rect -1679 23 1679 34
rect -1679 -23 -1668 23
rect 1668 -23 1679 23
rect -1679 -34 1679 -23
<< end >>
