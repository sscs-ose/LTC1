magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3245 -2180 3245 2180
<< metal2 >>
rect -1245 170 1245 180
rect -1245 114 -1235 170
rect -1179 114 -1093 170
rect -1037 114 -951 170
rect -895 114 -809 170
rect -753 114 -667 170
rect -611 114 -525 170
rect -469 114 -383 170
rect -327 114 -241 170
rect -185 114 -99 170
rect -43 114 43 170
rect 99 114 185 170
rect 241 114 327 170
rect 383 114 469 170
rect 525 114 611 170
rect 667 114 753 170
rect 809 114 895 170
rect 951 114 1037 170
rect 1093 114 1179 170
rect 1235 114 1245 170
rect -1245 28 1245 114
rect -1245 -28 -1235 28
rect -1179 -28 -1093 28
rect -1037 -28 -951 28
rect -895 -28 -809 28
rect -753 -28 -667 28
rect -611 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 611 28
rect 667 -28 753 28
rect 809 -28 895 28
rect 951 -28 1037 28
rect 1093 -28 1179 28
rect 1235 -28 1245 28
rect -1245 -114 1245 -28
rect -1245 -170 -1235 -114
rect -1179 -170 -1093 -114
rect -1037 -170 -951 -114
rect -895 -170 -809 -114
rect -753 -170 -667 -114
rect -611 -170 -525 -114
rect -469 -170 -383 -114
rect -327 -170 -241 -114
rect -185 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 185 -114
rect 241 -170 327 -114
rect 383 -170 469 -114
rect 525 -170 611 -114
rect 667 -170 753 -114
rect 809 -170 895 -114
rect 951 -170 1037 -114
rect 1093 -170 1179 -114
rect 1235 -170 1245 -114
rect -1245 -180 1245 -170
<< via2 >>
rect -1235 114 -1179 170
rect -1093 114 -1037 170
rect -951 114 -895 170
rect -809 114 -753 170
rect -667 114 -611 170
rect -525 114 -469 170
rect -383 114 -327 170
rect -241 114 -185 170
rect -99 114 -43 170
rect 43 114 99 170
rect 185 114 241 170
rect 327 114 383 170
rect 469 114 525 170
rect 611 114 667 170
rect 753 114 809 170
rect 895 114 951 170
rect 1037 114 1093 170
rect 1179 114 1235 170
rect -1235 -28 -1179 28
rect -1093 -28 -1037 28
rect -951 -28 -895 28
rect -809 -28 -753 28
rect -667 -28 -611 28
rect -525 -28 -469 28
rect -383 -28 -327 28
rect -241 -28 -185 28
rect -99 -28 -43 28
rect 43 -28 99 28
rect 185 -28 241 28
rect 327 -28 383 28
rect 469 -28 525 28
rect 611 -28 667 28
rect 753 -28 809 28
rect 895 -28 951 28
rect 1037 -28 1093 28
rect 1179 -28 1235 28
rect -1235 -170 -1179 -114
rect -1093 -170 -1037 -114
rect -951 -170 -895 -114
rect -809 -170 -753 -114
rect -667 -170 -611 -114
rect -525 -170 -469 -114
rect -383 -170 -327 -114
rect -241 -170 -185 -114
rect -99 -170 -43 -114
rect 43 -170 99 -114
rect 185 -170 241 -114
rect 327 -170 383 -114
rect 469 -170 525 -114
rect 611 -170 667 -114
rect 753 -170 809 -114
rect 895 -170 951 -114
rect 1037 -170 1093 -114
rect 1179 -170 1235 -114
<< metal3 >>
rect -1245 170 1245 180
rect -1245 114 -1235 170
rect -1179 114 -1093 170
rect -1037 114 -951 170
rect -895 114 -809 170
rect -753 114 -667 170
rect -611 114 -525 170
rect -469 114 -383 170
rect -327 114 -241 170
rect -185 114 -99 170
rect -43 114 43 170
rect 99 114 185 170
rect 241 114 327 170
rect 383 114 469 170
rect 525 114 611 170
rect 667 114 753 170
rect 809 114 895 170
rect 951 114 1037 170
rect 1093 114 1179 170
rect 1235 114 1245 170
rect -1245 28 1245 114
rect -1245 -28 -1235 28
rect -1179 -28 -1093 28
rect -1037 -28 -951 28
rect -895 -28 -809 28
rect -753 -28 -667 28
rect -611 -28 -525 28
rect -469 -28 -383 28
rect -327 -28 -241 28
rect -185 -28 -99 28
rect -43 -28 43 28
rect 99 -28 185 28
rect 241 -28 327 28
rect 383 -28 469 28
rect 525 -28 611 28
rect 667 -28 753 28
rect 809 -28 895 28
rect 951 -28 1037 28
rect 1093 -28 1179 28
rect 1235 -28 1245 28
rect -1245 -114 1245 -28
rect -1245 -170 -1235 -114
rect -1179 -170 -1093 -114
rect -1037 -170 -951 -114
rect -895 -170 -809 -114
rect -753 -170 -667 -114
rect -611 -170 -525 -114
rect -469 -170 -383 -114
rect -327 -170 -241 -114
rect -185 -170 -99 -114
rect -43 -170 43 -114
rect 99 -170 185 -114
rect 241 -170 327 -114
rect 383 -170 469 -114
rect 525 -170 611 -114
rect 667 -170 753 -114
rect 809 -170 895 -114
rect 951 -170 1037 -114
rect 1093 -170 1179 -114
rect 1235 -170 1245 -114
rect -1245 -180 1245 -170
<< end >>
