magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1484 -1298 1484 1298
<< metal2 >>
rect -484 293 484 298
rect -484 265 -479 293
rect -451 265 -417 293
rect -389 265 -355 293
rect -327 265 -293 293
rect -265 265 -231 293
rect -203 265 -169 293
rect -141 265 -107 293
rect -79 265 -45 293
rect -17 265 17 293
rect 45 265 79 293
rect 107 265 141 293
rect 169 265 203 293
rect 231 265 265 293
rect 293 265 327 293
rect 355 265 389 293
rect 417 265 451 293
rect 479 265 484 293
rect -484 231 484 265
rect -484 203 -479 231
rect -451 203 -417 231
rect -389 203 -355 231
rect -327 203 -293 231
rect -265 203 -231 231
rect -203 203 -169 231
rect -141 203 -107 231
rect -79 203 -45 231
rect -17 203 17 231
rect 45 203 79 231
rect 107 203 141 231
rect 169 203 203 231
rect 231 203 265 231
rect 293 203 327 231
rect 355 203 389 231
rect 417 203 451 231
rect 479 203 484 231
rect -484 169 484 203
rect -484 141 -479 169
rect -451 141 -417 169
rect -389 141 -355 169
rect -327 141 -293 169
rect -265 141 -231 169
rect -203 141 -169 169
rect -141 141 -107 169
rect -79 141 -45 169
rect -17 141 17 169
rect 45 141 79 169
rect 107 141 141 169
rect 169 141 203 169
rect 231 141 265 169
rect 293 141 327 169
rect 355 141 389 169
rect 417 141 451 169
rect 479 141 484 169
rect -484 107 484 141
rect -484 79 -479 107
rect -451 79 -417 107
rect -389 79 -355 107
rect -327 79 -293 107
rect -265 79 -231 107
rect -203 79 -169 107
rect -141 79 -107 107
rect -79 79 -45 107
rect -17 79 17 107
rect 45 79 79 107
rect 107 79 141 107
rect 169 79 203 107
rect 231 79 265 107
rect 293 79 327 107
rect 355 79 389 107
rect 417 79 451 107
rect 479 79 484 107
rect -484 45 484 79
rect -484 17 -479 45
rect -451 17 -417 45
rect -389 17 -355 45
rect -327 17 -293 45
rect -265 17 -231 45
rect -203 17 -169 45
rect -141 17 -107 45
rect -79 17 -45 45
rect -17 17 17 45
rect 45 17 79 45
rect 107 17 141 45
rect 169 17 203 45
rect 231 17 265 45
rect 293 17 327 45
rect 355 17 389 45
rect 417 17 451 45
rect 479 17 484 45
rect -484 -17 484 17
rect -484 -45 -479 -17
rect -451 -45 -417 -17
rect -389 -45 -355 -17
rect -327 -45 -293 -17
rect -265 -45 -231 -17
rect -203 -45 -169 -17
rect -141 -45 -107 -17
rect -79 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 79 -17
rect 107 -45 141 -17
rect 169 -45 203 -17
rect 231 -45 265 -17
rect 293 -45 327 -17
rect 355 -45 389 -17
rect 417 -45 451 -17
rect 479 -45 484 -17
rect -484 -79 484 -45
rect -484 -107 -479 -79
rect -451 -107 -417 -79
rect -389 -107 -355 -79
rect -327 -107 -293 -79
rect -265 -107 -231 -79
rect -203 -107 -169 -79
rect -141 -107 -107 -79
rect -79 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 79 -79
rect 107 -107 141 -79
rect 169 -107 203 -79
rect 231 -107 265 -79
rect 293 -107 327 -79
rect 355 -107 389 -79
rect 417 -107 451 -79
rect 479 -107 484 -79
rect -484 -141 484 -107
rect -484 -169 -479 -141
rect -451 -169 -417 -141
rect -389 -169 -355 -141
rect -327 -169 -293 -141
rect -265 -169 -231 -141
rect -203 -169 -169 -141
rect -141 -169 -107 -141
rect -79 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 79 -141
rect 107 -169 141 -141
rect 169 -169 203 -141
rect 231 -169 265 -141
rect 293 -169 327 -141
rect 355 -169 389 -141
rect 417 -169 451 -141
rect 479 -169 484 -141
rect -484 -203 484 -169
rect -484 -231 -479 -203
rect -451 -231 -417 -203
rect -389 -231 -355 -203
rect -327 -231 -293 -203
rect -265 -231 -231 -203
rect -203 -231 -169 -203
rect -141 -231 -107 -203
rect -79 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 79 -203
rect 107 -231 141 -203
rect 169 -231 203 -203
rect 231 -231 265 -203
rect 293 -231 327 -203
rect 355 -231 389 -203
rect 417 -231 451 -203
rect 479 -231 484 -203
rect -484 -265 484 -231
rect -484 -293 -479 -265
rect -451 -293 -417 -265
rect -389 -293 -355 -265
rect -327 -293 -293 -265
rect -265 -293 -231 -265
rect -203 -293 -169 -265
rect -141 -293 -107 -265
rect -79 -293 -45 -265
rect -17 -293 17 -265
rect 45 -293 79 -265
rect 107 -293 141 -265
rect 169 -293 203 -265
rect 231 -293 265 -265
rect 293 -293 327 -265
rect 355 -293 389 -265
rect 417 -293 451 -265
rect 479 -293 484 -265
rect -484 -298 484 -293
<< via2 >>
rect -479 265 -451 293
rect -417 265 -389 293
rect -355 265 -327 293
rect -293 265 -265 293
rect -231 265 -203 293
rect -169 265 -141 293
rect -107 265 -79 293
rect -45 265 -17 293
rect 17 265 45 293
rect 79 265 107 293
rect 141 265 169 293
rect 203 265 231 293
rect 265 265 293 293
rect 327 265 355 293
rect 389 265 417 293
rect 451 265 479 293
rect -479 203 -451 231
rect -417 203 -389 231
rect -355 203 -327 231
rect -293 203 -265 231
rect -231 203 -203 231
rect -169 203 -141 231
rect -107 203 -79 231
rect -45 203 -17 231
rect 17 203 45 231
rect 79 203 107 231
rect 141 203 169 231
rect 203 203 231 231
rect 265 203 293 231
rect 327 203 355 231
rect 389 203 417 231
rect 451 203 479 231
rect -479 141 -451 169
rect -417 141 -389 169
rect -355 141 -327 169
rect -293 141 -265 169
rect -231 141 -203 169
rect -169 141 -141 169
rect -107 141 -79 169
rect -45 141 -17 169
rect 17 141 45 169
rect 79 141 107 169
rect 141 141 169 169
rect 203 141 231 169
rect 265 141 293 169
rect 327 141 355 169
rect 389 141 417 169
rect 451 141 479 169
rect -479 79 -451 107
rect -417 79 -389 107
rect -355 79 -327 107
rect -293 79 -265 107
rect -231 79 -203 107
rect -169 79 -141 107
rect -107 79 -79 107
rect -45 79 -17 107
rect 17 79 45 107
rect 79 79 107 107
rect 141 79 169 107
rect 203 79 231 107
rect 265 79 293 107
rect 327 79 355 107
rect 389 79 417 107
rect 451 79 479 107
rect -479 17 -451 45
rect -417 17 -389 45
rect -355 17 -327 45
rect -293 17 -265 45
rect -231 17 -203 45
rect -169 17 -141 45
rect -107 17 -79 45
rect -45 17 -17 45
rect 17 17 45 45
rect 79 17 107 45
rect 141 17 169 45
rect 203 17 231 45
rect 265 17 293 45
rect 327 17 355 45
rect 389 17 417 45
rect 451 17 479 45
rect -479 -45 -451 -17
rect -417 -45 -389 -17
rect -355 -45 -327 -17
rect -293 -45 -265 -17
rect -231 -45 -203 -17
rect -169 -45 -141 -17
rect -107 -45 -79 -17
rect -45 -45 -17 -17
rect 17 -45 45 -17
rect 79 -45 107 -17
rect 141 -45 169 -17
rect 203 -45 231 -17
rect 265 -45 293 -17
rect 327 -45 355 -17
rect 389 -45 417 -17
rect 451 -45 479 -17
rect -479 -107 -451 -79
rect -417 -107 -389 -79
rect -355 -107 -327 -79
rect -293 -107 -265 -79
rect -231 -107 -203 -79
rect -169 -107 -141 -79
rect -107 -107 -79 -79
rect -45 -107 -17 -79
rect 17 -107 45 -79
rect 79 -107 107 -79
rect 141 -107 169 -79
rect 203 -107 231 -79
rect 265 -107 293 -79
rect 327 -107 355 -79
rect 389 -107 417 -79
rect 451 -107 479 -79
rect -479 -169 -451 -141
rect -417 -169 -389 -141
rect -355 -169 -327 -141
rect -293 -169 -265 -141
rect -231 -169 -203 -141
rect -169 -169 -141 -141
rect -107 -169 -79 -141
rect -45 -169 -17 -141
rect 17 -169 45 -141
rect 79 -169 107 -141
rect 141 -169 169 -141
rect 203 -169 231 -141
rect 265 -169 293 -141
rect 327 -169 355 -141
rect 389 -169 417 -141
rect 451 -169 479 -141
rect -479 -231 -451 -203
rect -417 -231 -389 -203
rect -355 -231 -327 -203
rect -293 -231 -265 -203
rect -231 -231 -203 -203
rect -169 -231 -141 -203
rect -107 -231 -79 -203
rect -45 -231 -17 -203
rect 17 -231 45 -203
rect 79 -231 107 -203
rect 141 -231 169 -203
rect 203 -231 231 -203
rect 265 -231 293 -203
rect 327 -231 355 -203
rect 389 -231 417 -203
rect 451 -231 479 -203
rect -479 -293 -451 -265
rect -417 -293 -389 -265
rect -355 -293 -327 -265
rect -293 -293 -265 -265
rect -231 -293 -203 -265
rect -169 -293 -141 -265
rect -107 -293 -79 -265
rect -45 -293 -17 -265
rect 17 -293 45 -265
rect 79 -293 107 -265
rect 141 -293 169 -265
rect 203 -293 231 -265
rect 265 -293 293 -265
rect 327 -293 355 -265
rect 389 -293 417 -265
rect 451 -293 479 -265
<< metal3 >>
rect -484 293 484 298
rect -484 265 -479 293
rect -451 265 -417 293
rect -389 265 -355 293
rect -327 265 -293 293
rect -265 265 -231 293
rect -203 265 -169 293
rect -141 265 -107 293
rect -79 265 -45 293
rect -17 265 17 293
rect 45 265 79 293
rect 107 265 141 293
rect 169 265 203 293
rect 231 265 265 293
rect 293 265 327 293
rect 355 265 389 293
rect 417 265 451 293
rect 479 265 484 293
rect -484 231 484 265
rect -484 203 -479 231
rect -451 203 -417 231
rect -389 203 -355 231
rect -327 203 -293 231
rect -265 203 -231 231
rect -203 203 -169 231
rect -141 203 -107 231
rect -79 203 -45 231
rect -17 203 17 231
rect 45 203 79 231
rect 107 203 141 231
rect 169 203 203 231
rect 231 203 265 231
rect 293 203 327 231
rect 355 203 389 231
rect 417 203 451 231
rect 479 203 484 231
rect -484 169 484 203
rect -484 141 -479 169
rect -451 141 -417 169
rect -389 141 -355 169
rect -327 141 -293 169
rect -265 141 -231 169
rect -203 141 -169 169
rect -141 141 -107 169
rect -79 141 -45 169
rect -17 141 17 169
rect 45 141 79 169
rect 107 141 141 169
rect 169 141 203 169
rect 231 141 265 169
rect 293 141 327 169
rect 355 141 389 169
rect 417 141 451 169
rect 479 141 484 169
rect -484 107 484 141
rect -484 79 -479 107
rect -451 79 -417 107
rect -389 79 -355 107
rect -327 79 -293 107
rect -265 79 -231 107
rect -203 79 -169 107
rect -141 79 -107 107
rect -79 79 -45 107
rect -17 79 17 107
rect 45 79 79 107
rect 107 79 141 107
rect 169 79 203 107
rect 231 79 265 107
rect 293 79 327 107
rect 355 79 389 107
rect 417 79 451 107
rect 479 79 484 107
rect -484 45 484 79
rect -484 17 -479 45
rect -451 17 -417 45
rect -389 17 -355 45
rect -327 17 -293 45
rect -265 17 -231 45
rect -203 17 -169 45
rect -141 17 -107 45
rect -79 17 -45 45
rect -17 17 17 45
rect 45 17 79 45
rect 107 17 141 45
rect 169 17 203 45
rect 231 17 265 45
rect 293 17 327 45
rect 355 17 389 45
rect 417 17 451 45
rect 479 17 484 45
rect -484 -17 484 17
rect -484 -45 -479 -17
rect -451 -45 -417 -17
rect -389 -45 -355 -17
rect -327 -45 -293 -17
rect -265 -45 -231 -17
rect -203 -45 -169 -17
rect -141 -45 -107 -17
rect -79 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 79 -17
rect 107 -45 141 -17
rect 169 -45 203 -17
rect 231 -45 265 -17
rect 293 -45 327 -17
rect 355 -45 389 -17
rect 417 -45 451 -17
rect 479 -45 484 -17
rect -484 -79 484 -45
rect -484 -107 -479 -79
rect -451 -107 -417 -79
rect -389 -107 -355 -79
rect -327 -107 -293 -79
rect -265 -107 -231 -79
rect -203 -107 -169 -79
rect -141 -107 -107 -79
rect -79 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 79 -79
rect 107 -107 141 -79
rect 169 -107 203 -79
rect 231 -107 265 -79
rect 293 -107 327 -79
rect 355 -107 389 -79
rect 417 -107 451 -79
rect 479 -107 484 -79
rect -484 -141 484 -107
rect -484 -169 -479 -141
rect -451 -169 -417 -141
rect -389 -169 -355 -141
rect -327 -169 -293 -141
rect -265 -169 -231 -141
rect -203 -169 -169 -141
rect -141 -169 -107 -141
rect -79 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 79 -141
rect 107 -169 141 -141
rect 169 -169 203 -141
rect 231 -169 265 -141
rect 293 -169 327 -141
rect 355 -169 389 -141
rect 417 -169 451 -141
rect 479 -169 484 -141
rect -484 -203 484 -169
rect -484 -231 -479 -203
rect -451 -231 -417 -203
rect -389 -231 -355 -203
rect -327 -231 -293 -203
rect -265 -231 -231 -203
rect -203 -231 -169 -203
rect -141 -231 -107 -203
rect -79 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 79 -203
rect 107 -231 141 -203
rect 169 -231 203 -203
rect 231 -231 265 -203
rect 293 -231 327 -203
rect 355 -231 389 -203
rect 417 -231 451 -203
rect 479 -231 484 -203
rect -484 -265 484 -231
rect -484 -293 -479 -265
rect -451 -293 -417 -265
rect -389 -293 -355 -265
rect -327 -293 -293 -265
rect -265 -293 -231 -265
rect -203 -293 -169 -265
rect -141 -293 -107 -265
rect -79 -293 -45 -265
rect -17 -293 17 -265
rect 45 -293 79 -265
rect 107 -293 141 -265
rect 169 -293 203 -265
rect 231 -293 265 -265
rect 293 -293 327 -265
rect 355 -293 389 -265
rect 417 -293 451 -265
rect 479 -293 484 -265
rect -484 -298 484 -293
<< end >>
