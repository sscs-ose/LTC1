magic
tech gf180mcuC
magscale 1 10
timestamp 1693222705
<< psubdiff >>
rect 596 7821 750 7838
rect 596 7766 610 7821
rect 734 7766 750 7821
rect 596 7753 750 7766
<< psubdiffcont >>
rect 610 7766 734 7821
<< polysilicon >>
rect 112 7950 212 7964
rect 112 7878 126 7950
rect 198 7878 212 7950
rect 112 7792 212 7878
rect 316 7960 416 7974
rect 316 7888 330 7960
rect 402 7888 416 7960
rect 316 7792 416 7888
<< polycontact >>
rect 126 7878 198 7950
rect 330 7888 402 7960
<< metal1 >>
rect 321 7960 411 7969
rect 117 7950 207 7959
rect 117 7878 126 7950
rect 198 7878 207 7950
rect 321 7888 330 7960
rect 402 7888 411 7960
rect 321 7879 411 7888
rect 117 7869 207 7878
rect 37 7735 83 7833
rect 445 7821 757 7844
rect 445 7766 610 7821
rect 734 7766 757 7821
rect 445 7750 757 7766
rect 445 7746 491 7750
use nmos_3p3_P8GAH7  nmos_3p3_P8GAH7_0
timestamp 1693222705
transform 1 0 366 0 1 3908
box -162 -3908 162 3908
use nmos_3p3_P8GAH7  nmos_3p3_P8GAH7_1
timestamp 1693222705
transform 1 0 162 0 1 3908
box -162 -3908 162 3908
<< labels >>
flabel polycontact 157 7907 157 7907 0 FreeSans 160 0 0 0 IM_T
port 0 nsew
flabel polycontact 375 7911 375 7911 0 FreeSans 160 0 0 0 IM
port 1 nsew
flabel metal1 60 7823 60 7823 0 FreeSans 160 0 0 0 OUT
port 2 nsew
flabel psubdiffcont 670 7795 670 7795 0 FreeSans 160 0 0 0 VSS
port 3 nsew
<< end >>
