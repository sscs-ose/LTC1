magic
tech gf180mcuC
magscale 1 10
timestamp 1693309239
<< pwell >>
rect 0 584 6648 960
rect 0 93 6648 469
<< nmos >>
rect 112 652 212 892
rect 316 652 416 892
rect 520 652 620 892
rect 724 652 824 892
rect 928 652 1028 892
rect 1132 652 1232 892
rect 1336 652 1436 892
rect 1540 652 1640 892
rect 1744 652 1844 892
rect 1948 652 2048 892
rect 2152 652 2252 892
rect 2356 652 2456 892
rect 2560 652 2660 892
rect 2764 652 2864 892
rect 2968 652 3068 892
rect 3172 652 3272 892
rect 3376 652 3476 892
rect 3580 652 3680 892
rect 3784 652 3884 892
rect 3988 652 4088 892
rect 4192 652 4292 892
rect 4396 652 4496 892
rect 4600 652 4700 892
rect 4804 652 4904 892
rect 5008 652 5108 892
rect 5212 652 5312 892
rect 5416 652 5516 892
rect 5620 652 5720 892
rect 5824 652 5924 892
rect 6028 652 6128 892
rect 6232 652 6332 892
rect 6436 652 6536 892
rect 112 161 212 401
rect 316 161 416 401
rect 520 161 620 401
rect 724 161 824 401
rect 928 161 1028 401
rect 1132 161 1232 401
rect 1336 161 1436 401
rect 1540 161 1640 401
rect 1744 161 1844 401
rect 1948 161 2048 401
rect 2152 161 2252 401
rect 2356 161 2456 401
rect 2560 161 2660 401
rect 2764 161 2864 401
rect 2968 161 3068 401
rect 3172 161 3272 401
rect 3376 161 3476 401
rect 3580 161 3680 401
rect 3784 161 3884 401
rect 3988 161 4088 401
rect 4192 161 4292 401
rect 4396 161 4496 401
rect 4600 161 4700 401
rect 4804 161 4904 401
rect 5008 161 5108 401
rect 5212 161 5312 401
rect 5416 161 5516 401
rect 5620 161 5720 401
rect 5824 161 5924 401
rect 6028 161 6128 401
rect 6232 161 6332 401
rect 6436 161 6536 401
<< ndiff >>
rect 24 879 112 892
rect 24 665 37 879
rect 83 665 112 879
rect 24 652 112 665
rect 212 879 316 892
rect 212 665 241 879
rect 287 665 316 879
rect 212 652 316 665
rect 416 879 520 892
rect 416 665 445 879
rect 491 665 520 879
rect 416 652 520 665
rect 620 879 724 892
rect 620 665 649 879
rect 695 665 724 879
rect 620 652 724 665
rect 824 879 928 892
rect 824 665 853 879
rect 899 665 928 879
rect 824 652 928 665
rect 1028 879 1132 892
rect 1028 665 1057 879
rect 1103 665 1132 879
rect 1028 652 1132 665
rect 1232 879 1336 892
rect 1232 665 1261 879
rect 1307 665 1336 879
rect 1232 652 1336 665
rect 1436 879 1540 892
rect 1436 665 1465 879
rect 1511 665 1540 879
rect 1436 652 1540 665
rect 1640 879 1744 892
rect 1640 665 1669 879
rect 1715 665 1744 879
rect 1640 652 1744 665
rect 1844 879 1948 892
rect 1844 665 1873 879
rect 1919 665 1948 879
rect 1844 652 1948 665
rect 2048 879 2152 892
rect 2048 665 2077 879
rect 2123 665 2152 879
rect 2048 652 2152 665
rect 2252 879 2356 892
rect 2252 665 2281 879
rect 2327 665 2356 879
rect 2252 652 2356 665
rect 2456 879 2560 892
rect 2456 665 2485 879
rect 2531 665 2560 879
rect 2456 652 2560 665
rect 2660 879 2764 892
rect 2660 665 2689 879
rect 2735 665 2764 879
rect 2660 652 2764 665
rect 2864 879 2968 892
rect 2864 665 2893 879
rect 2939 665 2968 879
rect 2864 652 2968 665
rect 3068 879 3172 892
rect 3068 665 3097 879
rect 3143 665 3172 879
rect 3068 652 3172 665
rect 3272 879 3376 892
rect 3272 665 3301 879
rect 3347 665 3376 879
rect 3272 652 3376 665
rect 3476 879 3580 892
rect 3476 665 3505 879
rect 3551 665 3580 879
rect 3476 652 3580 665
rect 3680 879 3784 892
rect 3680 665 3709 879
rect 3755 665 3784 879
rect 3680 652 3784 665
rect 3884 879 3988 892
rect 3884 665 3913 879
rect 3959 665 3988 879
rect 3884 652 3988 665
rect 4088 879 4192 892
rect 4088 665 4117 879
rect 4163 665 4192 879
rect 4088 652 4192 665
rect 4292 879 4396 892
rect 4292 665 4321 879
rect 4367 665 4396 879
rect 4292 652 4396 665
rect 4496 879 4600 892
rect 4496 665 4525 879
rect 4571 665 4600 879
rect 4496 652 4600 665
rect 4700 879 4804 892
rect 4700 665 4729 879
rect 4775 665 4804 879
rect 4700 652 4804 665
rect 4904 879 5008 892
rect 4904 665 4933 879
rect 4979 665 5008 879
rect 4904 652 5008 665
rect 5108 879 5212 892
rect 5108 665 5137 879
rect 5183 665 5212 879
rect 5108 652 5212 665
rect 5312 879 5416 892
rect 5312 665 5341 879
rect 5387 665 5416 879
rect 5312 652 5416 665
rect 5516 879 5620 892
rect 5516 665 5545 879
rect 5591 665 5620 879
rect 5516 652 5620 665
rect 5720 879 5824 892
rect 5720 665 5749 879
rect 5795 665 5824 879
rect 5720 652 5824 665
rect 5924 879 6028 892
rect 5924 665 5953 879
rect 5999 665 6028 879
rect 5924 652 6028 665
rect 6128 879 6232 892
rect 6128 665 6157 879
rect 6203 665 6232 879
rect 6128 652 6232 665
rect 6332 879 6436 892
rect 6332 665 6361 879
rect 6407 665 6436 879
rect 6332 652 6436 665
rect 6536 879 6624 892
rect 6536 665 6565 879
rect 6611 665 6624 879
rect 6536 652 6624 665
rect 24 388 112 401
rect 24 174 37 388
rect 83 174 112 388
rect 24 161 112 174
rect 212 388 316 401
rect 212 174 241 388
rect 287 174 316 388
rect 212 161 316 174
rect 416 388 520 401
rect 416 174 445 388
rect 491 174 520 388
rect 416 161 520 174
rect 620 388 724 401
rect 620 174 649 388
rect 695 174 724 388
rect 620 161 724 174
rect 824 388 928 401
rect 824 174 853 388
rect 899 174 928 388
rect 824 161 928 174
rect 1028 388 1132 401
rect 1028 174 1057 388
rect 1103 174 1132 388
rect 1028 161 1132 174
rect 1232 388 1336 401
rect 1232 174 1261 388
rect 1307 174 1336 388
rect 1232 161 1336 174
rect 1436 388 1540 401
rect 1436 174 1465 388
rect 1511 174 1540 388
rect 1436 161 1540 174
rect 1640 388 1744 401
rect 1640 174 1669 388
rect 1715 174 1744 388
rect 1640 161 1744 174
rect 1844 388 1948 401
rect 1844 174 1873 388
rect 1919 174 1948 388
rect 1844 161 1948 174
rect 2048 388 2152 401
rect 2048 174 2077 388
rect 2123 174 2152 388
rect 2048 161 2152 174
rect 2252 388 2356 401
rect 2252 174 2281 388
rect 2327 174 2356 388
rect 2252 161 2356 174
rect 2456 388 2560 401
rect 2456 174 2485 388
rect 2531 174 2560 388
rect 2456 161 2560 174
rect 2660 388 2764 401
rect 2660 174 2689 388
rect 2735 174 2764 388
rect 2660 161 2764 174
rect 2864 388 2968 401
rect 2864 174 2893 388
rect 2939 174 2968 388
rect 2864 161 2968 174
rect 3068 388 3172 401
rect 3068 174 3097 388
rect 3143 174 3172 388
rect 3068 161 3172 174
rect 3272 388 3376 401
rect 3272 174 3301 388
rect 3347 174 3376 388
rect 3272 161 3376 174
rect 3476 388 3580 401
rect 3476 174 3505 388
rect 3551 174 3580 388
rect 3476 161 3580 174
rect 3680 388 3784 401
rect 3680 174 3709 388
rect 3755 174 3784 388
rect 3680 161 3784 174
rect 3884 388 3988 401
rect 3884 174 3913 388
rect 3959 174 3988 388
rect 3884 161 3988 174
rect 4088 388 4192 401
rect 4088 174 4117 388
rect 4163 174 4192 388
rect 4088 161 4192 174
rect 4292 388 4396 401
rect 4292 174 4321 388
rect 4367 174 4396 388
rect 4292 161 4396 174
rect 4496 388 4600 401
rect 4496 174 4525 388
rect 4571 174 4600 388
rect 4496 161 4600 174
rect 4700 388 4804 401
rect 4700 174 4729 388
rect 4775 174 4804 388
rect 4700 161 4804 174
rect 4904 388 5008 401
rect 4904 174 4933 388
rect 4979 174 5008 388
rect 4904 161 5008 174
rect 5108 388 5212 401
rect 5108 174 5137 388
rect 5183 174 5212 388
rect 5108 161 5212 174
rect 5312 388 5416 401
rect 5312 174 5341 388
rect 5387 174 5416 388
rect 5312 161 5416 174
rect 5516 388 5620 401
rect 5516 174 5545 388
rect 5591 174 5620 388
rect 5516 161 5620 174
rect 5720 388 5824 401
rect 5720 174 5749 388
rect 5795 174 5824 388
rect 5720 161 5824 174
rect 5924 388 6028 401
rect 5924 174 5953 388
rect 5999 174 6028 388
rect 5924 161 6028 174
rect 6128 388 6232 401
rect 6128 174 6157 388
rect 6203 174 6232 388
rect 6128 161 6232 174
rect 6332 388 6436 401
rect 6332 174 6361 388
rect 6407 174 6436 388
rect 6332 161 6436 174
rect 6536 388 6624 401
rect 6536 174 6565 388
rect 6611 174 6624 388
rect 6536 161 6624 174
<< ndiffc >>
rect 37 665 83 879
rect 241 665 287 879
rect 445 665 491 879
rect 649 665 695 879
rect 853 665 899 879
rect 1057 665 1103 879
rect 1261 665 1307 879
rect 1465 665 1511 879
rect 1669 665 1715 879
rect 1873 665 1919 879
rect 2077 665 2123 879
rect 2281 665 2327 879
rect 2485 665 2531 879
rect 2689 665 2735 879
rect 2893 665 2939 879
rect 3097 665 3143 879
rect 3301 665 3347 879
rect 3505 665 3551 879
rect 3709 665 3755 879
rect 3913 665 3959 879
rect 4117 665 4163 879
rect 4321 665 4367 879
rect 4525 665 4571 879
rect 4729 665 4775 879
rect 4933 665 4979 879
rect 5137 665 5183 879
rect 5341 665 5387 879
rect 5545 665 5591 879
rect 5749 665 5795 879
rect 5953 665 5999 879
rect 6157 665 6203 879
rect 6361 665 6407 879
rect 6565 665 6611 879
rect 37 174 83 388
rect 241 174 287 388
rect 445 174 491 388
rect 649 174 695 388
rect 853 174 899 388
rect 1057 174 1103 388
rect 1261 174 1307 388
rect 1465 174 1511 388
rect 1669 174 1715 388
rect 1873 174 1919 388
rect 2077 174 2123 388
rect 2281 174 2327 388
rect 2485 174 2531 388
rect 2689 174 2735 388
rect 2893 174 2939 388
rect 3097 174 3143 388
rect 3301 174 3347 388
rect 3505 174 3551 388
rect 3709 174 3755 388
rect 3913 174 3959 388
rect 4117 174 4163 388
rect 4321 174 4367 388
rect 4525 174 4571 388
rect 4729 174 4775 388
rect 4933 174 4979 388
rect 5137 174 5183 388
rect 5341 174 5387 388
rect 5545 174 5591 388
rect 5749 174 5795 388
rect 5953 174 5999 388
rect 6157 174 6203 388
rect 6361 174 6407 388
rect 6565 174 6611 388
<< psubdiff >>
rect 0 1259 6715 1285
rect 0 1128 48 1259
rect 193 1128 348 1259
rect 493 1128 648 1259
rect 793 1128 948 1259
rect 1093 1128 1248 1259
rect 1393 1128 1548 1259
rect 1693 1128 1848 1259
rect 1993 1128 2148 1259
rect 2293 1128 2448 1259
rect 2593 1128 2748 1259
rect 2893 1128 3048 1259
rect 3193 1128 3348 1259
rect 3493 1128 3648 1259
rect 3793 1128 3948 1259
rect 4093 1128 4248 1259
rect 4393 1128 4548 1259
rect 4693 1128 4848 1259
rect 4993 1128 5148 1259
rect 5293 1128 5448 1259
rect 5593 1128 5748 1259
rect 5893 1128 6048 1259
rect 6193 1128 6348 1259
rect 6493 1128 6715 1259
rect 0 1098 6715 1128
rect 0 -50 6715 -21
rect 0 -181 44 -50
rect 189 -181 344 -50
rect 489 -181 644 -50
rect 789 -181 944 -50
rect 1089 -181 1244 -50
rect 1389 -181 1544 -50
rect 1689 -181 1844 -50
rect 1989 -181 2144 -50
rect 2289 -181 2444 -50
rect 2589 -181 2744 -50
rect 2889 -181 3044 -50
rect 3189 -181 3344 -50
rect 3489 -181 3644 -50
rect 3789 -181 3944 -50
rect 4089 -181 4244 -50
rect 4389 -181 4544 -50
rect 4689 -181 4844 -50
rect 4989 -181 5144 -50
rect 5289 -181 5444 -50
rect 5589 -181 5744 -50
rect 5889 -181 6044 -50
rect 6189 -181 6344 -50
rect 6489 -181 6715 -50
rect 0 -208 6715 -181
<< psubdiffcont >>
rect 48 1128 193 1259
rect 348 1128 493 1259
rect 648 1128 793 1259
rect 948 1128 1093 1259
rect 1248 1128 1393 1259
rect 1548 1128 1693 1259
rect 1848 1128 1993 1259
rect 2148 1128 2293 1259
rect 2448 1128 2593 1259
rect 2748 1128 2893 1259
rect 3048 1128 3193 1259
rect 3348 1128 3493 1259
rect 3648 1128 3793 1259
rect 3948 1128 4093 1259
rect 4248 1128 4393 1259
rect 4548 1128 4693 1259
rect 4848 1128 4993 1259
rect 5148 1128 5293 1259
rect 5448 1128 5593 1259
rect 5748 1128 5893 1259
rect 6048 1128 6193 1259
rect 6348 1128 6493 1259
rect 44 -181 189 -50
rect 344 -181 489 -50
rect 644 -181 789 -50
rect 944 -181 1089 -50
rect 1244 -181 1389 -50
rect 1544 -181 1689 -50
rect 1844 -181 1989 -50
rect 2144 -181 2289 -50
rect 2444 -181 2589 -50
rect 2744 -181 2889 -50
rect 3044 -181 3189 -50
rect 3344 -181 3489 -50
rect 3644 -181 3789 -50
rect 3944 -181 4089 -50
rect 4244 -181 4389 -50
rect 4544 -181 4689 -50
rect 4844 -181 4989 -50
rect 5144 -181 5289 -50
rect 5444 -181 5589 -50
rect 5744 -181 5889 -50
rect 6044 -181 6189 -50
rect 6344 -181 6489 -50
<< polysilicon >>
rect -168 1077 -82 1091
rect -168 1073 6536 1077
rect -168 1024 -150 1073
rect -102 1024 6536 1073
rect -168 1019 6536 1024
rect -168 1008 -82 1019
rect 112 892 212 1019
rect 316 892 416 936
rect 520 892 620 936
rect 724 892 824 1019
rect 928 892 1028 1019
rect 1132 892 1232 936
rect 1336 892 1436 936
rect 1540 892 1640 1019
rect 1744 892 1844 1019
rect 1948 892 2048 936
rect 2152 892 2252 936
rect 2356 892 2456 1019
rect 2560 892 2660 1019
rect 2764 892 2864 936
rect 2968 892 3068 936
rect 3172 892 3272 1019
rect 3376 892 3476 1019
rect 3580 892 3680 936
rect 3784 892 3884 936
rect 3988 892 4088 1019
rect 4192 892 4292 1019
rect 4396 892 4496 936
rect 4600 892 4700 936
rect 4804 892 4904 1019
rect 5008 892 5108 1019
rect 5212 892 5312 936
rect 5416 892 5516 936
rect 5620 892 5720 1019
rect 5824 892 5924 1019
rect 6028 892 6128 936
rect 6232 892 6332 936
rect 6436 892 6536 1019
rect 112 608 212 652
rect -171 553 -84 566
rect 316 553 416 652
rect 520 553 620 652
rect 724 608 824 652
rect 928 608 1028 652
rect 1132 553 1232 652
rect 1336 553 1436 652
rect 1540 608 1640 652
rect 1744 608 1844 652
rect 1948 553 2048 652
rect 2152 553 2252 652
rect 2356 608 2456 652
rect 2560 608 2660 652
rect 2764 553 2864 652
rect 2968 553 3068 652
rect 3172 608 3272 652
rect 3376 608 3476 652
rect 3580 553 3680 652
rect 3784 553 3884 652
rect 3988 608 4088 652
rect 4192 608 4292 652
rect 4396 553 4496 652
rect 4600 553 4700 652
rect 4804 608 4904 652
rect 5008 608 5108 652
rect 5212 553 5312 652
rect 5416 553 5516 652
rect 5620 608 5720 652
rect 5824 608 5924 652
rect 6028 553 6128 652
rect 6232 553 6332 652
rect 6436 608 6536 652
rect -171 552 6536 553
rect -171 499 -158 552
rect -102 499 6536 552
rect -171 494 6536 499
rect -171 485 -84 494
rect 112 401 212 494
rect 316 401 416 445
rect 520 401 620 445
rect 724 401 824 494
rect 928 401 1028 494
rect 1132 401 1232 445
rect 1336 401 1436 445
rect 1540 401 1640 494
rect 1744 401 1844 494
rect 1948 401 2048 445
rect 2152 401 2252 445
rect 2356 401 2456 494
rect 2560 401 2660 494
rect 2764 401 2864 445
rect 2968 401 3068 445
rect 3172 401 3272 494
rect 3376 401 3476 494
rect 3580 401 3680 445
rect 3784 401 3884 445
rect 3988 401 4088 494
rect 4192 401 4292 494
rect 4396 401 4496 445
rect 4600 401 4700 445
rect 4804 401 4904 494
rect 5008 401 5108 494
rect 5212 401 5312 445
rect 5416 401 5516 445
rect 5620 401 5720 494
rect 5824 401 5924 494
rect 6028 401 6128 445
rect 6232 401 6332 445
rect 6436 401 6536 494
rect 112 117 212 161
rect -166 58 -74 74
rect 316 58 416 161
rect 520 58 620 161
rect 724 117 824 161
rect 928 117 1028 161
rect 1132 58 1232 161
rect 1336 58 1436 161
rect 1540 117 1640 161
rect 1744 117 1844 161
rect 1948 58 2048 161
rect 2152 58 2252 161
rect 2356 117 2456 161
rect 2560 117 2660 161
rect 2764 58 2864 161
rect 2968 58 3068 161
rect 3172 117 3272 161
rect 3376 117 3476 161
rect 3580 58 3680 161
rect 3784 58 3884 161
rect 3988 117 4088 161
rect 4192 117 4292 161
rect 4396 58 4496 161
rect 4600 58 4700 161
rect 4804 117 4904 161
rect 5008 117 5108 161
rect 5212 58 5312 161
rect 5416 58 5516 161
rect 5620 117 5720 161
rect 5824 117 5924 161
rect 6028 58 6128 161
rect 6232 58 6332 161
rect 6436 117 6536 161
rect -166 53 6332 58
rect -166 2 -150 53
rect -102 2 6332 53
rect -166 -1 6332 2
rect -166 -14 -74 -1
<< polycontact >>
rect -150 1024 -102 1073
rect -158 499 -102 552
rect -150 2 -102 53
<< metal1 >>
rect 0 1259 6715 1285
rect 0 1128 48 1259
rect 193 1128 348 1259
rect 493 1128 648 1259
rect 793 1128 948 1259
rect 1093 1128 1248 1259
rect 1393 1128 1548 1259
rect 1693 1128 1848 1259
rect 1993 1128 2148 1259
rect 2293 1128 2448 1259
rect 2593 1128 2748 1259
rect 2893 1128 3048 1259
rect 3193 1128 3348 1259
rect 3493 1128 3648 1259
rect 3793 1128 3948 1259
rect 4093 1128 4248 1259
rect 4393 1128 4548 1259
rect 4693 1128 4848 1259
rect 4993 1128 5148 1259
rect 5293 1128 5448 1259
rect 5593 1128 5748 1259
rect 5893 1128 6048 1259
rect 6193 1128 6348 1259
rect 6493 1230 6715 1259
rect 6493 1158 6567 1230
rect 6656 1158 6715 1230
rect 6493 1128 6715 1158
rect 0 1098 6715 1128
rect -168 1076 -82 1091
rect -168 1020 -155 1076
rect -99 1020 -82 1076
rect -168 1008 -82 1020
rect 37 879 83 890
rect 241 879 287 890
rect 219 826 241 843
rect 445 879 491 1098
rect 287 826 304 843
rect 219 766 233 826
rect 290 766 304 826
rect 219 752 241 766
rect 37 591 83 665
rect 287 752 304 766
rect 241 654 287 665
rect 649 879 695 890
rect 632 830 649 844
rect 853 879 899 890
rect 695 830 717 844
rect 632 771 647 830
rect 702 771 717 830
rect 632 753 649 771
rect 445 654 491 665
rect 695 753 717 771
rect 649 654 695 665
rect 1057 879 1103 890
rect 1044 748 1057 838
rect 1261 879 1307 1098
rect 1103 824 1129 838
rect 1114 765 1129 824
rect 853 591 899 665
rect 1103 748 1129 765
rect 1057 654 1103 665
rect 1465 879 1511 890
rect 1444 830 1465 844
rect 1669 879 1715 890
rect 1511 830 1529 844
rect 1444 771 1459 830
rect 1514 771 1529 830
rect 1444 753 1465 771
rect 1261 654 1307 665
rect 1511 753 1529 771
rect 1465 654 1511 665
rect 1873 879 1919 890
rect 1857 812 1873 826
rect 2077 879 2123 1098
rect 1919 812 1942 826
rect 1857 753 1872 812
rect 1927 753 1942 812
rect 1857 735 1873 753
rect 1669 591 1715 665
rect 1919 735 1942 753
rect 1873 654 1919 665
rect 2281 879 2327 890
rect 2267 746 2281 837
rect 2485 879 2531 890
rect 2327 823 2352 837
rect 2337 764 2352 823
rect 2077 654 2123 665
rect 2327 746 2352 764
rect 2281 654 2327 665
rect 2689 879 2735 890
rect 2664 812 2689 826
rect 2893 879 2939 1098
rect 2664 753 2679 812
rect 2664 735 2689 753
rect 2485 591 2531 665
rect 2735 735 2749 826
rect 2689 654 2735 665
rect 3097 879 3143 890
rect 3079 817 3097 831
rect 3301 879 3347 890
rect 3143 817 3164 831
rect 3079 758 3094 817
rect 3149 758 3164 817
rect 3079 740 3097 758
rect 2893 654 2939 665
rect 3143 740 3164 758
rect 3097 654 3143 665
rect 3505 879 3551 890
rect 3490 743 3505 834
rect 3709 879 3755 1098
rect 3551 820 3575 834
rect 3560 761 3575 820
rect 3301 591 3347 665
rect 3551 743 3575 761
rect 3505 654 3551 665
rect 3913 879 3959 890
rect 3900 753 3913 844
rect 4117 879 4163 890
rect 3959 830 3985 844
rect 3970 771 3985 830
rect 3709 654 3755 665
rect 3959 753 3985 771
rect 3913 654 3959 665
rect 4321 879 4367 890
rect 4305 812 4321 826
rect 4525 879 4571 1098
rect 4367 812 4390 826
rect 4305 753 4320 812
rect 4375 753 4390 812
rect 4305 735 4321 753
rect 4117 591 4163 665
rect 4367 735 4390 753
rect 4321 654 4367 665
rect 4729 879 4775 890
rect 4707 812 4729 826
rect 4933 879 4979 890
rect 4775 812 4792 826
rect 4707 753 4722 812
rect 4777 753 4792 812
rect 4707 735 4729 753
rect 4525 654 4571 665
rect 4775 735 4792 753
rect 4729 654 4775 665
rect 5137 879 5183 890
rect 5123 748 5137 839
rect 5341 879 5387 1098
rect 5183 825 5208 839
rect 5193 766 5208 825
rect 4933 591 4979 665
rect 5183 748 5208 766
rect 5137 654 5183 665
rect 5545 879 5591 890
rect 5523 817 5545 831
rect 5749 879 5795 890
rect 5591 817 5608 831
rect 5523 758 5538 817
rect 5593 758 5608 817
rect 5523 740 5545 758
rect 5341 654 5387 665
rect 5591 740 5608 758
rect 5545 654 5591 665
rect 5953 879 5999 890
rect 5940 737 5953 828
rect 6157 879 6203 1098
rect 5999 814 6025 828
rect 6010 755 6025 814
rect 5749 591 5795 665
rect 5999 737 6025 755
rect 5953 654 5999 665
rect 6361 879 6407 890
rect 6328 820 6361 834
rect 6565 879 6611 890
rect 6328 761 6343 820
rect 6328 743 6361 761
rect 6157 654 6203 665
rect 6407 743 6413 834
rect 6361 654 6407 665
rect 6565 591 6611 665
rect -171 552 -84 566
rect -171 499 -158 552
rect -102 499 -84 552
rect 37 519 6915 591
rect -171 485 -84 499
rect 37 388 83 399
rect 241 388 287 399
rect 221 321 241 338
rect 445 388 491 519
rect 287 321 306 338
rect 221 262 235 321
rect 290 262 306 321
rect 221 247 241 262
rect -166 58 -74 74
rect -166 1 -151 58
rect -94 1 -74 58
rect -166 -14 -74 1
rect 37 -21 83 174
rect 287 247 306 262
rect 241 163 287 174
rect 649 388 695 399
rect 642 249 649 340
rect 853 388 899 399
rect 695 326 727 340
rect 712 267 727 326
rect 445 163 491 174
rect 695 249 727 267
rect 649 163 695 174
rect 1057 388 1103 399
rect 1038 342 1057 356
rect 1261 388 1307 519
rect 1103 342 1123 356
rect 1038 283 1053 342
rect 1108 283 1123 342
rect 1038 265 1057 283
rect 853 -21 899 174
rect 1103 265 1123 283
rect 1057 163 1103 174
rect 1465 388 1511 399
rect 1451 270 1465 361
rect 1669 388 1715 399
rect 1511 347 1536 361
rect 1521 288 1536 347
rect 1261 163 1307 174
rect 1511 270 1536 288
rect 1465 163 1511 174
rect 1873 388 1919 399
rect 1851 345 1873 359
rect 2077 388 2123 519
rect 1919 345 1936 359
rect 1851 286 1866 345
rect 1921 286 1936 345
rect 1851 268 1873 286
rect 1669 -21 1715 174
rect 1919 268 1936 286
rect 1873 163 1919 174
rect 2281 388 2327 399
rect 2254 335 2281 349
rect 2485 388 2531 399
rect 2254 276 2269 335
rect 2254 258 2281 276
rect 2077 163 2123 174
rect 2327 258 2339 349
rect 2281 163 2327 174
rect 2689 388 2735 399
rect 2677 260 2689 351
rect 2893 388 2939 519
rect 2735 337 2762 351
rect 2747 278 2762 337
rect 2485 -21 2531 174
rect 2735 260 2762 278
rect 2689 163 2735 174
rect 3097 388 3143 399
rect 3077 321 3097 335
rect 3301 388 3347 399
rect 3143 321 3162 335
rect 3077 262 3092 321
rect 3147 262 3162 321
rect 3077 244 3097 262
rect 2893 163 2939 174
rect 3143 244 3162 262
rect 3097 163 3143 174
rect 3505 388 3551 399
rect 3486 336 3505 338
rect 3479 322 3505 336
rect 3709 388 3755 519
rect 3551 336 3562 338
rect 3479 263 3494 322
rect 3479 245 3505 263
rect 3301 -21 3347 174
rect 3551 245 3564 336
rect 3505 163 3551 174
rect 3913 388 3959 399
rect 3892 337 3913 351
rect 4117 388 4163 399
rect 3959 337 3977 351
rect 3892 278 3907 337
rect 3962 278 3977 337
rect 3892 260 3913 278
rect 3709 163 3755 174
rect 3959 260 3977 278
rect 3913 163 3959 174
rect 4321 388 4367 399
rect 4295 306 4321 320
rect 4525 388 4571 519
rect 4295 247 4310 306
rect 4295 229 4321 247
rect 4117 -21 4163 174
rect 4367 229 4380 320
rect 4321 163 4367 174
rect 4729 388 4775 399
rect 4712 316 4729 330
rect 4933 388 4979 399
rect 4775 316 4797 330
rect 4712 257 4727 316
rect 4782 257 4797 316
rect 4712 239 4729 257
rect 4525 163 4571 174
rect 4775 239 4797 257
rect 4729 163 4775 174
rect 5137 388 5183 399
rect 5120 329 5137 343
rect 5341 388 5387 519
rect 5183 329 5205 343
rect 5120 270 5135 329
rect 5190 270 5205 329
rect 5120 252 5137 270
rect 4933 -21 4979 174
rect 5183 252 5205 270
rect 5137 163 5183 174
rect 5545 388 5591 399
rect 5520 331 5545 345
rect 5749 388 5795 399
rect 5520 272 5535 331
rect 5520 254 5545 272
rect 5341 163 5387 174
rect 5591 254 5605 345
rect 5545 163 5591 174
rect 5953 388 5999 399
rect 5935 332 5953 346
rect 6157 388 6203 519
rect 5999 332 6020 346
rect 5935 273 5950 332
rect 6005 273 6020 332
rect 5935 255 5953 273
rect 5749 -21 5795 174
rect 5999 255 6020 273
rect 5953 163 5999 174
rect 6361 388 6407 399
rect 6343 319 6361 333
rect 6565 388 6611 399
rect 6407 319 6428 333
rect 6343 260 6358 319
rect 6413 260 6428 319
rect 6343 242 6361 260
rect 6157 163 6203 174
rect 6407 242 6428 260
rect 6361 163 6407 174
rect 6565 -21 6611 174
rect 0 -50 6715 -21
rect 0 -181 44 -50
rect 189 -181 344 -50
rect 489 -181 644 -50
rect 789 -181 944 -50
rect 1089 -181 1244 -50
rect 1389 -181 1544 -50
rect 1689 -181 1844 -50
rect 1989 -181 2144 -50
rect 2289 -181 2444 -50
rect 2589 -181 2744 -50
rect 2889 -181 3044 -50
rect 3189 -181 3344 -50
rect 3489 -181 3644 -50
rect 3789 -181 3944 -50
rect 4089 -181 4244 -50
rect 4389 -181 4544 -50
rect 4689 -181 4844 -50
rect 4989 -181 5144 -50
rect 5289 -181 5444 -50
rect 5589 -181 5744 -50
rect 5889 -181 6044 -50
rect 6189 -181 6344 -50
rect 6489 -86 6715 -50
rect 6489 -153 6581 -86
rect 6648 -153 6715 -86
rect 6489 -181 6715 -153
rect 0 -208 6715 -181
<< via1 >>
rect 6567 1158 6656 1230
rect -155 1073 -99 1076
rect -155 1024 -150 1073
rect -150 1024 -102 1073
rect -102 1024 -99 1073
rect -155 1020 -99 1024
rect 233 766 241 826
rect 241 766 287 826
rect 287 766 290 826
rect 647 771 649 830
rect 649 771 695 830
rect 695 771 702 830
rect 1059 765 1103 824
rect 1103 765 1114 824
rect 1459 771 1465 830
rect 1465 771 1511 830
rect 1511 771 1514 830
rect 1872 753 1873 812
rect 1873 753 1919 812
rect 1919 753 1927 812
rect 2282 764 2327 823
rect 2327 764 2337 823
rect 2679 753 2689 812
rect 2689 753 2734 812
rect 3094 758 3097 817
rect 3097 758 3143 817
rect 3143 758 3149 817
rect 3505 761 3551 820
rect 3551 761 3560 820
rect 3915 771 3959 830
rect 3959 771 3970 830
rect 4320 753 4321 812
rect 4321 753 4367 812
rect 4367 753 4375 812
rect 4722 753 4729 812
rect 4729 753 4775 812
rect 4775 753 4777 812
rect 5138 766 5183 825
rect 5183 766 5193 825
rect 5538 758 5545 817
rect 5545 758 5591 817
rect 5591 758 5593 817
rect 5955 755 5999 814
rect 5999 755 6010 814
rect 6343 761 6361 820
rect 6361 761 6398 820
rect 235 262 241 321
rect 241 262 287 321
rect 287 262 290 321
rect -151 53 -94 58
rect -151 2 -150 53
rect -150 2 -102 53
rect -102 2 -94 53
rect -151 1 -94 2
rect 657 267 695 326
rect 695 267 712 326
rect 1053 283 1057 342
rect 1057 283 1103 342
rect 1103 283 1108 342
rect 1466 288 1511 347
rect 1511 288 1521 347
rect 1866 286 1873 345
rect 1873 286 1919 345
rect 1919 286 1921 345
rect 2269 276 2281 335
rect 2281 276 2324 335
rect 2692 278 2735 337
rect 2735 278 2747 337
rect 3092 262 3097 321
rect 3097 262 3143 321
rect 3143 262 3147 321
rect 3494 263 3505 322
rect 3505 263 3549 322
rect 3907 278 3913 337
rect 3913 278 3959 337
rect 3959 278 3962 337
rect 4310 247 4321 306
rect 4321 247 4365 306
rect 4727 257 4729 316
rect 4729 257 4775 316
rect 4775 257 4782 316
rect 5135 270 5137 329
rect 5137 270 5183 329
rect 5183 270 5190 329
rect 5535 272 5545 331
rect 5545 272 5590 331
rect 5950 273 5953 332
rect 5953 273 5999 332
rect 5999 273 6005 332
rect 6358 260 6361 319
rect 6361 260 6407 319
rect 6407 260 6413 319
rect 6581 -153 6648 -86
<< metal2 >>
rect 6547 1230 6686 1257
rect 6547 1158 6567 1230
rect 6656 1158 6686 1230
rect 6547 1133 6686 1158
rect -168 1076 -82 1091
rect -168 1020 -155 1076
rect -99 1020 -82 1076
rect -168 1008 -82 1020
rect -156 74 -98 1008
rect 219 826 304 843
rect 219 766 233 826
rect 290 766 304 826
rect 219 752 304 766
rect 632 830 717 844
rect 632 771 647 830
rect 702 771 717 830
rect 632 753 717 771
rect 1044 824 1129 838
rect 1044 765 1059 824
rect 1114 765 1129 824
rect 233 338 290 752
rect 650 340 707 753
rect 1044 748 1129 765
rect 1444 830 1529 844
rect 1444 771 1459 830
rect 1514 771 1529 830
rect 1444 753 1529 771
rect 1857 812 1942 826
rect 1857 753 1872 812
rect 1927 753 1942 812
rect 1058 356 1115 748
rect 1459 361 1516 753
rect 1857 735 1942 753
rect 2267 823 2352 837
rect 2267 764 2282 823
rect 2337 764 2352 823
rect 2267 746 2352 764
rect 2664 812 2749 826
rect 2664 753 2679 812
rect 2734 753 2749 812
rect 1038 342 1123 356
rect 221 336 306 338
rect 642 336 727 340
rect 1038 336 1053 342
rect 221 326 1053 336
rect 221 321 657 326
rect 221 262 235 321
rect 290 279 657 321
rect 290 262 306 279
rect 221 247 306 262
rect 642 267 657 279
rect 712 283 1053 326
rect 1108 336 1123 342
rect 1451 347 1536 361
rect 1867 359 1924 735
rect 1451 336 1466 347
rect 1108 288 1466 336
rect 1521 336 1536 347
rect 1851 345 1936 359
rect 2270 349 2327 746
rect 2664 735 2749 753
rect 3079 817 3164 831
rect 3079 758 3094 817
rect 3149 758 3164 817
rect 3079 740 3164 758
rect 3490 820 3575 834
rect 3490 761 3505 820
rect 3560 761 3575 820
rect 3490 743 3575 761
rect 3900 830 3985 844
rect 3900 771 3915 830
rect 3970 771 3985 830
rect 3900 753 3985 771
rect 4305 812 4390 826
rect 4305 753 4320 812
rect 4375 753 4390 812
rect 2684 351 2741 735
rect 1851 336 1866 345
rect 1521 288 1866 336
rect 1108 286 1866 288
rect 1921 336 1936 345
rect 2254 336 2339 349
rect 2677 337 2762 351
rect 2677 336 2692 337
rect 1921 335 2692 336
rect 1921 286 2269 335
rect 1108 283 2269 286
rect 712 279 2269 283
rect 712 267 727 279
rect 642 249 727 267
rect 1038 265 1123 279
rect 1451 270 1536 279
rect 1851 268 1936 279
rect 2254 276 2269 279
rect 2324 279 2692 335
rect 2324 276 2339 279
rect 2254 258 2339 276
rect 2677 278 2692 279
rect 2747 336 2762 337
rect 3093 336 3150 740
rect 3495 336 3552 743
rect 3909 351 3966 753
rect 4305 735 4390 753
rect 4707 812 4792 826
rect 4707 753 4722 812
rect 4777 753 4792 812
rect 4707 735 4792 753
rect 5123 825 5208 839
rect 5123 766 5138 825
rect 5193 766 5208 825
rect 5123 748 5208 766
rect 5523 817 5608 831
rect 5523 758 5538 817
rect 5593 758 5608 817
rect 3892 337 3977 351
rect 3892 336 3907 337
rect 2747 322 3907 336
rect 2747 321 3494 322
rect 2747 279 3092 321
rect 2747 278 2762 279
rect 2677 260 2762 278
rect 3077 262 3092 279
rect 3147 279 3494 321
rect 3147 262 3162 279
rect 3077 244 3162 262
rect 3479 263 3494 279
rect 3549 279 3907 322
rect 3549 263 3564 279
rect 3479 245 3564 263
rect 3892 278 3907 279
rect 3962 336 3977 337
rect 4311 336 4368 735
rect 4719 336 4776 735
rect 5128 343 5185 748
rect 5523 740 5608 758
rect 5940 814 6025 828
rect 5940 755 5955 814
rect 6010 755 6025 814
rect 5526 345 5583 740
rect 5940 737 6025 755
rect 6328 820 6413 834
rect 6328 761 6343 820
rect 6398 761 6413 820
rect 6328 743 6413 761
rect 5942 346 5999 737
rect 5120 336 5205 343
rect 5520 336 5605 345
rect 5935 336 6020 346
rect 6345 336 6402 743
rect 3962 333 6402 336
rect 3962 332 6428 333
rect 3962 331 5950 332
rect 3962 329 5535 331
rect 3962 316 5135 329
rect 3962 306 4727 316
rect 3962 279 4310 306
rect 3962 278 3977 279
rect 3892 260 3977 278
rect 4295 247 4310 279
rect 4365 279 4727 306
rect 4365 247 4380 279
rect 4295 229 4380 247
rect 4712 257 4727 279
rect 4782 279 5135 316
rect 4782 257 4797 279
rect 4712 239 4797 257
rect 5120 270 5135 279
rect 5190 279 5535 329
rect 5190 270 5205 279
rect 5120 252 5205 270
rect 5520 272 5535 279
rect 5590 279 5950 331
rect 5590 272 5605 279
rect 5520 254 5605 272
rect 5935 273 5950 279
rect 6005 319 6428 332
rect 6005 279 6358 319
rect 6005 273 6020 279
rect 5935 255 6020 273
rect 6343 260 6358 279
rect 6413 260 6428 319
rect 6343 242 6428 260
rect -166 58 -74 74
rect -166 1 -151 58
rect -94 1 -74 58
rect -166 -14 -74 1
rect 6581 -75 6648 1133
rect 6564 -86 6667 -75
rect 6564 -153 6581 -86
rect 6648 -153 6667 -86
rect 6564 -168 6667 -153
<< labels >>
flabel via1 -133 1049 -133 1049 0 FreeSans 1600 0 0 0 IM_T
port 0 nsew
flabel metal1 1480 1192 1480 1192 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 6857 556 6857 556 0 FreeSans 1600 0 0 0 OUT
port 3 nsew
flabel metal1 -164 520 -164 520 0 FreeSans 1600 0 0 0 IM
port 4 nsew
flabel via1 2290 310 2290 310 0 FreeSans 1600 0 0 0 SD
port 5 nsew
<< end >>
