* NGSPICE file created from CM_16_flat.ext - technology: gf180mcuC

.subckt CM_16_flat VSS OUT IM IM_T
X0 OUT IM_T.t0 a_312_430# VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X1 a_312_430# IM_T.t1 OUT.t14 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X2 a_312_430# IM_T.t2 OUT.t13 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X3 a_312_430# IM_T.t3 OUT.t12 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X4 a_312_430# IM.t0 VSS.t34 VSS.t33 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X5 a_312_430# IM.t1 VSS.t10 VSS.t9 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X6 a_312_430# IM.t2 VSS.t1 VSS.t0 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X7 OUT IM_T.t4 a_312_430# VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X8 VSS IM.t3 a_312_430# VSS.t4 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X9 OUT IM_T.t5 a_312_430# VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X10 VSS IM.t4 a_312_430# VSS.t28 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X11 a_312_430# IM_T.t6 OUT.t9 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X12 a_312_430# IM.t5 VSS.t39 VSS.t38 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X13 a_312_430# IM.t6 VSS.t8 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=1u
X14 a_312_430# IM_T.t7 OUT.t8 VSS.t7 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=1u
X15 OUT IM_T.t8 a_312_430# VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X16 OUT IM_T.t9 a_312_430# VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X17 VSS IM.t7 a_312_430# VSS.t19 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X18 VSS IM.t8 a_312_430# VSS.t22 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X19 a_312_430# IM.t9 VSS.t15 VSS.t14 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X20 a_312_430# IM_T.t10 OUT.t5 VSS.t14 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X21 a_312_430# IM.t10 VSS.t3 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X22 a_312_430# IM_T.t11 OUT.t4 VSS.t2 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X23 a_312_430# IM.t11 VSS.t32 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X24 VSS IM.t12 a_312_430# VSS.t25 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X25 a_312_430# IM_T.t12 OUT.t3 VSS.t31 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X26 OUT IM_T.t13 a_312_430# VSS.t25 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=1u
X27 VSS IM.t13 a_312_430# VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X28 VSS IM.t14 a_312_430# VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X29 OUT IM_T.t14 a_312_430# VSS.t35 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X30 OUT IM_T.t15 a_312_430# VSS.t16 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
X31 VSS IM.t15 a_312_430# VSS.t11 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=1u
R0 IM_T.n9 IM_T.n8 147.633
R1 IM_T.n11 IM_T.n10 147.633
R2 IM_T.n13 IM_T.n12 147.633
R3 IM_T.n0 IM_T.t13 60.7907
R4 IM_T.n2 IM_T.n1 54.4633
R5 IM_T.n4 IM_T.n3 54.4633
R6 IM_T.n6 IM_T.n5 51.6849
R7 IM_T IM_T.n14 44.1578
R8 IM_T.n8 IM_T.t1 33.0769
R9 IM_T.n10 IM_T.n9 27.6763
R10 IM_T.n12 IM_T.n11 27.6763
R11 IM_T.n14 IM_T.n13 27.6763
R12 IM_T.n1 IM_T.n0 12.9829
R13 IM_T.n3 IM_T.n2 12.9829
R14 IM_T.n5 IM_T.n4 12.9829
R15 IM_T.n6 IM_T.t7 8.96331
R16 IM_T IM_T.n7 4.5005
R17 IM_T IM_T.n7 4.5005
R18 IM_T.n8 IM_T.t4 2.1905
R19 IM_T.n9 IM_T.t3 2.1905
R20 IM_T.n10 IM_T.t8 2.1905
R21 IM_T.n11 IM_T.t6 2.1905
R22 IM_T.n12 IM_T.t9 2.1905
R23 IM_T.n13 IM_T.t2 2.1905
R24 IM_T.n14 IM_T.t5 2.1905
R25 IM_T.n0 IM_T.t10 2.1905
R26 IM_T.n1 IM_T.t14 2.1905
R27 IM_T.n2 IM_T.t11 2.1905
R28 IM_T.n3 IM_T.t15 2.1905
R29 IM_T.n4 IM_T.t12 2.1905
R30 IM_T.n5 IM_T.t0 2.1905
R31 IM_T.n7 IM_T.n6 1.06651
R32 OUT.n15 OUT.t8 6.79341
R33 OUT.n22 OUT.n0 6.10941
R34 OUT.n15 OUT.n14 3.51246
R35 OUT.n17 OUT.n10 3.51246
R36 OUT.n19 OUT.n6 3.51246
R37 OUT.n21 OUT.n2 3.51246
R38 OUT.n20 OUT.n4 3.37941
R39 OUT.n18 OUT.n8 3.37941
R40 OUT.n16 OUT.n12 3.37941
R41 OUT.n4 OUT.t5 2.7305
R42 OUT.n4 OUT.n3 2.7305
R43 OUT.n8 OUT.t4 2.7305
R44 OUT.n8 OUT.n7 2.7305
R45 OUT.n12 OUT.t3 2.7305
R46 OUT.n12 OUT.n11 2.7305
R47 OUT.n14 OUT.t13 2.7305
R48 OUT.n14 OUT.n13 2.7305
R49 OUT.n10 OUT.t9 2.7305
R50 OUT.n10 OUT.n9 2.7305
R51 OUT.n6 OUT.t12 2.7305
R52 OUT.n6 OUT.n5 2.7305
R53 OUT.n2 OUT.t14 2.7305
R54 OUT.n2 OUT.n1 2.7305
R55 OUT.n22 OUT.n21 0.6845
R56 OUT.n21 OUT.n20 0.6845
R57 OUT.n20 OUT.n19 0.6845
R58 OUT.n19 OUT.n18 0.6845
R59 OUT.n18 OUT.n17 0.6845
R60 OUT.n17 OUT.n16 0.6845
R61 OUT.n16 OUT.n15 0.6845
R62 OUT OUT.n22 0.27275
R63 VSS.n24 VSS.t25 299.599
R64 VSS.n74 VSS.t2 238.811
R65 VSS.n61 VSS.t22 210.589
R66 VSS.n31 VSS.t4 171.511
R67 VSS.n17 VSS.t14 160.655
R68 VSS.n51 VSS.t28 149.8
R69 VSS.n1 VSS.t19 138.946
R70 VSS.n86 VSS.t31 121.576
R71 VSS.n64 VSS.t38 110.722
R72 VSS.t2 VSS.n73 89.0119
R73 VSS.n80 VSS.t9 78.1568
R74 VSS.n28 VSS.t33 71.6438
R75 VSS.n14 VSS.t35 60.7887
R76 VSS.n48 VSS.t7 49.9337
R77 VSS.n11 VSS.t0 39.0787
R78 VSS.n83 VSS.t11 21.7106
R79 VSS.n75 VSS.n2 11.6672
R80 VSS.n94 VSS.n75 11.6672
R81 VSS.n67 VSS.t16 10.8555
R82 VSS.n50 VSS.t8 6.55042
R83 VSS.n27 VSS.n5 6.52684
R84 VSS VSS.n75 5.2005
R85 VSS VSS.n75 5.2005
R86 VSS.n82 VSS.n79 3.85174
R87 VSS.n92 VSS.n77 3.80202
R88 VSS.n10 VSS.n9 3.80202
R89 VSS.n23 VSS.n7 3.80202
R90 VSS.n37 VSS.n4 3.75507
R91 VSS.n70 VSS.n45 3.75507
R92 VSS.n57 VSS.n47 3.75507
R93 VSS.n4 VSS.t15 2.7305
R94 VSS.n4 VSS.n3 2.7305
R95 VSS.n45 VSS.t3 2.7305
R96 VSS.n45 VSS.n44 2.7305
R97 VSS.n47 VSS.t32 2.7305
R98 VSS.n47 VSS.n46 2.7305
R99 VSS.n79 VSS.t10 2.7305
R100 VSS.n79 VSS.n78 2.7305
R101 VSS.n77 VSS.t39 2.7305
R102 VSS.n77 VSS.n76 2.7305
R103 VSS.n9 VSS.t1 2.7305
R104 VSS.n9 VSS.n8 2.7305
R105 VSS.n7 VSS.t34 2.7305
R106 VSS.n7 VSS.n6 2.7305
R107 VSS.n33 VSS.n32 2.6005
R108 VSS.n32 VSS.n31 2.6005
R109 VSS.n36 VSS.n35 2.6005
R110 VSS.n35 VSS.n34 2.6005
R111 VSS.n40 VSS.n39 2.6005
R112 VSS.n39 VSS.n38 2.6005
R113 VSS.n43 VSS.n42 2.6005
R114 VSS.n42 VSS.n41 2.6005
R115 VSS.n72 VSS.n71 2.6005
R116 VSS.n73 VSS.n72 2.6005
R117 VSS.n69 VSS.n68 2.6005
R118 VSS.n68 VSS.n67 2.6005
R119 VSS.n66 VSS.n65 2.6005
R120 VSS.n65 VSS.n64 2.6005
R121 VSS.n63 VSS.n62 2.6005
R122 VSS.n62 VSS.n61 2.6005
R123 VSS.n60 VSS.n59 2.6005
R124 VSS.n59 VSS.n58 2.6005
R125 VSS.n56 VSS.n55 2.6005
R126 VSS.n55 VSS.n54 2.6005
R127 VSS.n53 VSS.n52 2.6005
R128 VSS.n52 VSS.n51 2.6005
R129 VSS.n50 VSS.n49 2.6005
R130 VSS.n49 VSS.n48 2.6005
R131 VSS.n30 VSS.n29 2.6005
R132 VSS.n29 VSS.n28 2.6005
R133 VSS.n26 VSS.n25 2.6005
R134 VSS.n25 VSS.n24 2.6005
R135 VSS.n22 VSS.n21 2.6005
R136 VSS.n21 VSS.n20 2.6005
R137 VSS.n19 VSS.n18 2.6005
R138 VSS.n18 VSS.n17 2.6005
R139 VSS.n16 VSS.n15 2.6005
R140 VSS.n15 VSS.n14 2.6005
R141 VSS.n13 VSS.n12 2.6005
R142 VSS.n12 VSS.n11 2.6005
R143 VSS.n2 VSS.n0 2.6005
R144 VSS.n2 VSS.n1 2.6005
R145 VSS.n75 VSS.n74 2.6005
R146 VSS.n95 VSS.n94 2.6005
R147 VSS.n94 VSS.n93 2.6005
R148 VSS.n91 VSS.n90 2.6005
R149 VSS.n90 VSS.n89 2.6005
R150 VSS.n88 VSS.n87 2.6005
R151 VSS.n87 VSS.n86 2.6005
R152 VSS.n85 VSS.n84 2.6005
R153 VSS.n84 VSS.n83 2.6005
R154 VSS.n82 VSS.n81 2.6005
R155 VSS.n81 VSS.n80 2.6005
R156 VSS.n27 VSS.n26 1.90126
R157 VSS.n22 VSS.n19 0.1505
R158 VSS.n19 VSS.n16 0.1505
R159 VSS.n16 VSS.n13 0.1505
R160 VSS VSS.n0 0.1505
R161 VSS VSS.n95 0.1505
R162 VSS.n91 VSS.n88 0.1505
R163 VSS.n88 VSS.n85 0.1505
R164 VSS.n85 VSS.n82 0.1505
R165 VSS.n30 VSS.n27 0.142302
R166 VSS.n26 VSS.n23 0.136786
R167 VSS.n33 VSS.n30 0.131205
R168 VSS.n36 VSS.n33 0.131205
R169 VSS.n43 VSS.n40 0.131205
R170 VSS.n71 VSS.n43 0.131205
R171 VSS.n69 VSS.n66 0.131205
R172 VSS.n66 VSS.n63 0.131205
R173 VSS.n63 VSS.n60 0.131205
R174 VSS.n56 VSS.n53 0.131205
R175 VSS.n53 VSS.n50 0.131205
R176 VSS.n95 VSS.n92 0.129071
R177 VSS.n57 VSS.n56 0.127844
R178 VSS.n40 VSS.n37 0.121122
R179 VSS.n10 VSS.n0 0.0930714
R180 VSS.n71 VSS.n70 0.0725747
R181 VSS.n70 VSS.n69 0.0591307
R182 VSS.n13 VSS.n10 0.0579286
R183 VSS.n92 VSS.n91 0.0219286
R184 VSS.n23 VSS.n22 0.0142143
R185 VSS.n37 VSS.n36 0.010583
R186 VSS.n60 VSS.n57 0.003861
R187 IM.n16 IM.n14 35.4095
R188 IM.n0 IM.t12 32.6004
R189 IM.n1 IM.n0 30.5194
R190 IM.n5 IM.n4 30.5194
R191 IM.n9 IM.n8 30.5194
R192 IM.n13 IM.n12 30.5194
R193 IM.n2 IM.n1 30.2907
R194 IM.n4 IM.n3 30.2907
R195 IM.n6 IM.n5 30.2907
R196 IM.n8 IM.n7 30.2907
R197 IM.n10 IM.n9 30.2907
R198 IM.n12 IM.n11 30.2907
R199 IM.n14 IM.n13 30.2907
R200 IM.n3 IM.n2 30.0619
R201 IM.n7 IM.n6 30.0619
R202 IM.n11 IM.n10 30.0619
R203 IM IM.n16 4.00981
R204 IM.n0 IM.t0 2.1905
R205 IM.n1 IM.t3 2.1905
R206 IM.n2 IM.t9 2.1905
R207 IM.n3 IM.t13 2.1905
R208 IM.n4 IM.t2 2.1905
R209 IM.n5 IM.t7 2.1905
R210 IM.n6 IM.t10 2.1905
R211 IM.n7 IM.t14 2.1905
R212 IM.n8 IM.t5 2.1905
R213 IM.n9 IM.t8 2.1905
R214 IM.n10 IM.t11 2.1905
R215 IM.n11 IM.t15 2.1905
R216 IM.n12 IM.t1 2.1905
R217 IM.n13 IM.t4 2.1905
R218 IM.n14 IM.t6 2.1905
R219 IM.n16 IM.n15 0.336132
C0 IM IM_T 1.27f
C1 IM_T OUT 0.742f
C2 IM_T a_312_430# 0.831f
C3 IM OUT 0.959f
C4 IM a_312_430# 0.588f
C5 a_312_430# OUT 1.94f
.ends

