magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1316 1019 1316
<< metal2 >>
rect -19 311 19 316
rect -19 283 -14 311
rect 14 283 19 311
rect -19 245 19 283
rect -19 217 -14 245
rect 14 217 19 245
rect -19 179 19 217
rect -19 151 -14 179
rect 14 151 19 179
rect -19 113 19 151
rect -19 85 -14 113
rect 14 85 19 113
rect -19 47 19 85
rect -19 19 -14 47
rect 14 19 19 47
rect -19 -19 19 19
rect -19 -47 -14 -19
rect 14 -47 19 -19
rect -19 -85 19 -47
rect -19 -113 -14 -85
rect 14 -113 19 -85
rect -19 -151 19 -113
rect -19 -179 -14 -151
rect 14 -179 19 -151
rect -19 -217 19 -179
rect -19 -245 -14 -217
rect 14 -245 19 -217
rect -19 -283 19 -245
rect -19 -311 -14 -283
rect 14 -311 19 -283
rect -19 -316 19 -311
<< via2 >>
rect -14 283 14 311
rect -14 217 14 245
rect -14 151 14 179
rect -14 85 14 113
rect -14 19 14 47
rect -14 -47 14 -19
rect -14 -113 14 -85
rect -14 -179 14 -151
rect -14 -245 14 -217
rect -14 -311 14 -283
<< metal3 >>
rect -19 311 19 316
rect -19 283 -14 311
rect 14 283 19 311
rect -19 245 19 283
rect -19 217 -14 245
rect 14 217 19 245
rect -19 179 19 217
rect -19 151 -14 179
rect 14 151 19 179
rect -19 113 19 151
rect -19 85 -14 113
rect 14 85 19 113
rect -19 47 19 85
rect -19 19 -14 47
rect 14 19 19 47
rect -19 -19 19 19
rect -19 -47 -14 -19
rect 14 -47 19 -19
rect -19 -85 19 -47
rect -19 -113 -14 -85
rect 14 -113 19 -85
rect -19 -151 19 -113
rect -19 -179 -14 -151
rect 14 -179 19 -151
rect -19 -217 19 -179
rect -19 -245 -14 -217
rect 14 -245 19 -217
rect -19 -283 19 -245
rect -19 -311 -14 -283
rect 14 -311 19 -283
rect -19 -316 19 -311
<< end >>
