magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 3448 2344
<< mvnmos >>
rect 0 0 140 300
rect 244 0 384 300
rect 488 0 628 300
rect 732 0 872 300
rect 976 0 1116 300
rect 1220 0 1360 300
<< mvndiff >>
rect -88 287 0 300
rect -88 241 -75 287
rect -29 241 0 287
rect -88 173 0 241
rect -88 127 -75 173
rect -29 127 0 173
rect -88 59 0 127
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 287 244 300
rect 140 241 169 287
rect 215 241 244 287
rect 140 173 244 241
rect 140 127 169 173
rect 215 127 244 173
rect 140 59 244 127
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 287 488 300
rect 384 241 413 287
rect 459 241 488 287
rect 384 173 488 241
rect 384 127 413 173
rect 459 127 488 173
rect 384 59 488 127
rect 384 13 413 59
rect 459 13 488 59
rect 384 0 488 13
rect 628 287 732 300
rect 628 241 657 287
rect 703 241 732 287
rect 628 173 732 241
rect 628 127 657 173
rect 703 127 732 173
rect 628 59 732 127
rect 628 13 657 59
rect 703 13 732 59
rect 628 0 732 13
rect 872 287 976 300
rect 872 241 901 287
rect 947 241 976 287
rect 872 173 976 241
rect 872 127 901 173
rect 947 127 976 173
rect 872 59 976 127
rect 872 13 901 59
rect 947 13 976 59
rect 872 0 976 13
rect 1116 287 1220 300
rect 1116 241 1145 287
rect 1191 241 1220 287
rect 1116 173 1220 241
rect 1116 127 1145 173
rect 1191 127 1220 173
rect 1116 59 1220 127
rect 1116 13 1145 59
rect 1191 13 1220 59
rect 1116 0 1220 13
rect 1360 287 1448 300
rect 1360 241 1389 287
rect 1435 241 1448 287
rect 1360 173 1448 241
rect 1360 127 1389 173
rect 1435 127 1448 173
rect 1360 59 1448 127
rect 1360 13 1389 59
rect 1435 13 1448 59
rect 1360 0 1448 13
<< mvndiffc >>
rect -75 241 -29 287
rect -75 127 -29 173
rect -75 13 -29 59
rect 169 241 215 287
rect 169 127 215 173
rect 169 13 215 59
rect 413 241 459 287
rect 413 127 459 173
rect 413 13 459 59
rect 657 241 703 287
rect 657 127 703 173
rect 657 13 703 59
rect 901 241 947 287
rect 901 127 947 173
rect 901 13 947 59
rect 1145 241 1191 287
rect 1145 127 1191 173
rect 1145 13 1191 59
rect 1389 241 1435 287
rect 1389 127 1435 173
rect 1389 13 1435 59
<< polysilicon >>
rect 0 300 140 344
rect 244 300 384 344
rect 488 300 628 344
rect 732 300 872 344
rect 976 300 1116 344
rect 1220 300 1360 344
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
rect 976 -44 1116 0
rect 1220 -44 1360 0
<< metal1 >>
rect -75 287 -29 300
rect -75 173 -29 241
rect -75 59 -29 127
rect -75 0 -29 13
rect 169 287 215 300
rect 169 173 215 241
rect 169 59 215 127
rect 169 0 215 13
rect 413 287 459 300
rect 413 173 459 241
rect 413 59 459 127
rect 413 0 459 13
rect 657 287 703 300
rect 657 173 703 241
rect 657 59 703 127
rect 657 0 703 13
rect 901 287 947 300
rect 901 173 947 241
rect 901 59 947 127
rect 901 0 947 13
rect 1145 287 1191 300
rect 1145 173 1191 241
rect 1145 59 1191 127
rect 1145 0 1191 13
rect 1389 287 1435 300
rect 1389 173 1435 241
rect 1389 59 1435 127
rect 1389 0 1435 13
<< labels >>
rlabel mvndiffc 1168 150 1168 150 4 D
rlabel mvndiffc 924 150 924 150 4 S
rlabel mvndiffc 680 150 680 150 4 D
rlabel mvndiffc 436 150 436 150 4 S
rlabel mvndiffc 192 150 192 150 4 D
rlabel mvndiffc 1412 150 1412 150 4 S
rlabel mvndiffc -52 150 -52 150 4 S
<< end >>
