magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6578 -2278 6578 2278
<< nwell >>
rect -4578 -278 4578 278
<< nsubdiff >>
rect -4495 173 4495 195
rect -4495 -173 -4473 173
rect 4473 -173 4495 173
rect -4495 -195 4495 -173
<< nsubdiffcont >>
rect -4473 -173 4473 173
<< metal1 >>
rect -4484 173 4484 184
rect -4484 -173 -4473 173
rect 4473 -173 4484 173
rect -4484 -184 4484 -173
<< end >>
