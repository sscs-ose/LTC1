magic
tech gf180mcuC
magscale 1 10
timestamp 1692183930
<< nwell >>
rect 114 386 838 945
<< pwell >>
rect 4 82 796 280
rect 873 82 1161 280
<< nmos >>
rect 120 156 176 206
rect 288 156 344 206
rect 456 156 512 206
rect 624 156 680 206
rect 989 156 1045 206
<< pmos >>
rect 288 516 344 616
rect 448 516 504 616
rect 608 516 664 616
<< ndiff >>
rect 28 206 100 217
rect 196 206 268 217
rect 364 206 436 217
rect 532 206 604 217
rect 700 206 772 217
rect 28 204 120 206
rect 28 158 41 204
rect 87 158 120 204
rect 28 156 120 158
rect 176 204 288 206
rect 176 158 209 204
rect 255 158 288 204
rect 176 156 288 158
rect 344 204 456 206
rect 344 158 377 204
rect 423 158 456 204
rect 344 156 456 158
rect 512 204 624 206
rect 512 158 545 204
rect 591 158 624 204
rect 512 156 624 158
rect 680 204 772 206
rect 680 158 713 204
rect 759 158 772 204
rect 680 156 772 158
rect 28 145 100 156
rect 196 145 268 156
rect 364 145 436 156
rect 532 145 604 156
rect 700 145 772 156
rect 897 206 969 217
rect 1065 206 1137 217
rect 897 204 989 206
rect 897 158 910 204
rect 956 158 989 204
rect 897 156 989 158
rect 1045 204 1137 206
rect 1045 158 1078 204
rect 1124 158 1137 204
rect 1045 156 1137 158
rect 897 145 969 156
rect 1065 145 1137 156
<< pdiff >>
rect 200 603 288 616
rect 200 529 213 603
rect 259 529 288 603
rect 200 516 288 529
rect 344 603 448 616
rect 344 529 373 603
rect 419 529 448 603
rect 344 516 448 529
rect 504 603 608 616
rect 504 529 533 603
rect 579 529 608 603
rect 504 516 608 529
rect 664 603 752 616
rect 664 529 693 603
rect 739 529 752 603
rect 664 516 752 529
<< ndiffc >>
rect 41 158 87 204
rect 209 158 255 204
rect 377 158 423 204
rect 545 158 591 204
rect 713 158 759 204
rect 910 158 956 204
rect 1078 158 1124 204
<< pdiffc >>
rect 213 529 259 603
rect 373 529 419 603
rect 533 529 579 603
rect 693 529 739 603
<< psubdiff >>
rect 38 -14 201 1
rect 38 -73 55 -14
rect 184 -73 201 -14
rect 38 -88 201 -73
rect 283 -8 446 7
rect 283 -67 300 -8
rect 429 -67 446 -8
rect 283 -82 446 -67
rect 515 -11 678 4
rect 515 -70 532 -11
rect 661 -70 678 -11
rect 515 -85 678 -70
rect 762 -12 925 3
rect 762 -71 779 -12
rect 908 -71 925 -12
rect 762 -86 925 -71
rect 986 -12 1149 3
rect 986 -71 1003 -12
rect 1132 -71 1149 -12
rect 986 -86 1149 -71
<< nsubdiff >>
rect 150 900 295 915
rect 150 849 166 900
rect 282 849 295 900
rect 150 833 295 849
rect 401 902 546 918
rect 401 851 417 902
rect 533 851 546 902
rect 401 837 546 851
rect 641 901 786 916
rect 641 850 657 901
rect 773 850 786 901
rect 641 835 786 850
<< psubdiffcont >>
rect 55 -73 184 -14
rect 300 -67 429 -8
rect 532 -70 661 -11
rect 779 -71 908 -12
rect 1003 -71 1132 -12
<< nsubdiffcont >>
rect 166 849 282 900
rect 417 851 533 902
rect 657 850 773 901
<< polysilicon >>
rect 87 756 161 771
rect 87 710 101 756
rect 147 710 504 756
rect 87 696 161 710
rect 288 616 344 660
rect 448 616 504 710
rect 608 616 664 660
rect 70 320 150 335
rect 288 320 344 516
rect 448 472 504 516
rect 70 316 344 320
rect 70 267 86 316
rect 134 267 344 316
rect 70 264 344 267
rect 70 253 176 264
rect 120 206 176 253
rect 288 206 344 264
rect 456 310 504 472
rect 608 472 664 516
rect 608 464 1045 472
rect 598 454 1045 464
rect 571 436 1045 454
rect 571 390 591 436
rect 637 416 1045 436
rect 637 390 664 416
rect 571 383 664 390
rect 571 376 648 383
rect 456 262 680 310
rect 456 206 512 262
rect 624 206 680 262
rect 120 112 176 156
rect 288 112 344 156
rect 456 112 512 156
rect 624 112 680 156
rect 989 206 1045 416
rect 989 112 1045 156
<< polycontact >>
rect 101 710 147 756
rect 86 267 134 316
rect 591 390 637 436
<< metal1 >>
rect 114 902 838 945
rect 114 900 417 902
rect 114 849 166 900
rect 282 851 417 900
rect 533 901 838 902
rect 533 851 657 901
rect 282 850 657 851
rect 773 850 838 901
rect 282 849 838 850
rect 114 822 838 849
rect 87 758 161 771
rect 26 756 161 758
rect 26 712 101 756
rect 87 710 101 712
rect 147 710 161 756
rect 87 696 161 710
rect 213 603 259 822
rect 213 518 259 529
rect 373 603 419 614
rect 373 435 419 529
rect 533 603 579 822
rect 533 518 579 529
rect 693 603 739 614
rect 693 519 739 529
rect 693 472 1174 519
rect 571 436 648 454
rect 571 435 591 436
rect 209 390 591 435
rect 637 390 648 436
rect 209 389 648 390
rect 70 316 150 335
rect 70 315 86 316
rect -4 268 86 315
rect 70 267 86 268
rect 134 267 150 316
rect 70 253 150 267
rect 209 204 255 389
rect 571 376 648 389
rect 377 253 759 299
rect 377 206 423 253
rect 713 206 759 253
rect 366 204 434 206
rect 702 204 770 206
rect 1077 204 1124 472
rect 30 158 41 204
rect 87 158 98 204
rect 198 158 209 204
rect 255 158 266 204
rect 366 158 377 204
rect 423 158 434 204
rect 534 158 545 204
rect 591 158 602 204
rect 702 158 713 204
rect 759 158 770 204
rect 899 158 910 204
rect 956 158 967 204
rect 1067 158 1078 204
rect 1124 158 1135 204
rect 41 108 87 158
rect 377 108 423 158
rect 41 62 423 108
rect 545 12 591 158
rect 910 12 956 158
rect 3 -8 1161 12
rect 3 -14 300 -8
rect 3 -73 55 -14
rect 184 -67 300 -14
rect 429 -11 1161 -8
rect 429 -67 532 -11
rect 184 -70 532 -67
rect 661 -12 1161 -11
rect 661 -70 779 -12
rect 184 -71 779 -70
rect 908 -71 1003 -12
rect 1132 -71 1161 -12
rect 184 -73 1161 -71
rect 3 -102 1161 -73
<< labels >>
flabel metal1 19 296 19 296 0 FreeSans 800 0 0 0 A
port 1 nsew
flabel metal1 50 724 50 724 0 FreeSans 800 0 0 0 B
port 3 nsew
flabel metal1 1126 494 1126 494 0 FreeSans 320 0 0 0 OUT
port 9 nsew
flabel nsubdiffcont 447 891 447 891 0 FreeSans 320 0 0 0 VDD
port 10 nsew
flabel metal1 483 -42 483 -42 0 FreeSans 320 0 0 0 VSS
port 11 nsew
<< end >>
