magic
tech gf180mcuC
magscale 1 10
timestamp 1694155088
<< nwell >>
rect -864 -954 864 954
<< nsubdiff >>
rect -840 917 840 930
rect -840 871 -724 917
rect 724 871 840 917
rect -840 858 840 871
rect -840 814 -768 858
rect -840 -814 -827 814
rect -781 -814 -768 814
rect 768 814 840 858
rect -840 -858 -768 -814
rect 768 -814 781 814
rect 827 -814 840 814
rect 768 -858 840 -814
rect -840 -871 840 -858
rect -840 -917 -724 -871
rect 724 -917 840 -871
rect -840 -930 840 -917
<< nsubdiffcont >>
rect -724 871 724 917
rect -827 -814 -781 814
rect 781 -814 827 814
rect -724 -917 724 -871
<< polysilicon >>
rect -680 757 -520 770
rect -680 711 -667 757
rect -533 711 -520 757
rect -680 667 -520 711
rect -680 -711 -520 -667
rect -680 -757 -667 -711
rect -533 -757 -520 -711
rect -680 -770 -520 -757
rect -440 757 -280 770
rect -440 711 -427 757
rect -293 711 -280 757
rect -440 667 -280 711
rect -440 -711 -280 -667
rect -440 -757 -427 -711
rect -293 -757 -280 -711
rect -440 -770 -280 -757
rect -200 757 -40 770
rect -200 711 -187 757
rect -53 711 -40 757
rect -200 667 -40 711
rect -200 -711 -40 -667
rect -200 -757 -187 -711
rect -53 -757 -40 -711
rect -200 -770 -40 -757
rect 40 757 200 770
rect 40 711 53 757
rect 187 711 200 757
rect 40 667 200 711
rect 40 -711 200 -667
rect 40 -757 53 -711
rect 187 -757 200 -711
rect 40 -770 200 -757
rect 280 757 440 770
rect 280 711 293 757
rect 427 711 440 757
rect 280 667 440 711
rect 280 -711 440 -667
rect 280 -757 293 -711
rect 427 -757 440 -711
rect 280 -770 440 -757
rect 520 757 680 770
rect 520 711 533 757
rect 667 711 680 757
rect 520 667 680 711
rect 520 -711 680 -667
rect 520 -757 533 -711
rect 667 -757 680 -711
rect 520 -770 680 -757
<< polycontact >>
rect -667 711 -533 757
rect -667 -757 -533 -711
rect -427 711 -293 757
rect -427 -757 -293 -711
rect -187 711 -53 757
rect -187 -757 -53 -711
rect 53 711 187 757
rect 53 -757 187 -711
rect 293 711 427 757
rect 293 -757 427 -711
rect 533 711 667 757
rect 533 -757 667 -711
<< ppolyres >>
rect -680 -667 -520 667
rect -440 -667 -280 667
rect -200 -667 -40 667
rect 40 -667 200 667
rect 280 -667 440 667
rect 520 -667 680 667
<< metal1 >>
rect -827 871 -724 917
rect 724 871 827 917
rect -827 814 -781 871
rect 781 814 827 871
rect -678 711 -667 757
rect -533 711 -522 757
rect -438 711 -427 757
rect -293 711 -282 757
rect -198 711 -187 757
rect -53 711 -42 757
rect 42 711 53 757
rect 187 711 198 757
rect 282 711 293 757
rect 427 711 438 757
rect 522 711 533 757
rect 667 711 678 757
rect -678 -757 -667 -711
rect -533 -757 -522 -711
rect -438 -757 -427 -711
rect -293 -757 -282 -711
rect -198 -757 -187 -711
rect -53 -757 -42 -711
rect 42 -757 53 -711
rect 187 -757 198 -711
rect 282 -757 293 -711
rect 427 -757 438 -711
rect 522 -757 533 -711
rect 667 -757 678 -711
rect -827 -871 -781 -814
rect 781 -871 827 -814
rect -827 -917 -724 -871
rect 724 -917 827 -871
<< properties >>
string FIXED_BBOX -804 -894 804 894
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 6.672 m 1 nx 6 wmin 0.80 lmin 1.00 rho 315 val 2.879k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1
<< end >>
