magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1184 -1580 1184 1580
<< metal1 >>
rect -184 574 184 580
rect -184 548 -178 574
rect -152 548 -112 574
rect -86 548 -46 574
rect -20 548 20 574
rect 46 548 86 574
rect 112 548 152 574
rect 178 548 184 574
rect -184 508 184 548
rect -184 482 -178 508
rect -152 482 -112 508
rect -86 482 -46 508
rect -20 482 20 508
rect 46 482 86 508
rect 112 482 152 508
rect 178 482 184 508
rect -184 442 184 482
rect -184 416 -178 442
rect -152 416 -112 442
rect -86 416 -46 442
rect -20 416 20 442
rect 46 416 86 442
rect 112 416 152 442
rect 178 416 184 442
rect -184 376 184 416
rect -184 350 -178 376
rect -152 350 -112 376
rect -86 350 -46 376
rect -20 350 20 376
rect 46 350 86 376
rect 112 350 152 376
rect 178 350 184 376
rect -184 310 184 350
rect -184 284 -178 310
rect -152 284 -112 310
rect -86 284 -46 310
rect -20 284 20 310
rect 46 284 86 310
rect 112 284 152 310
rect 178 284 184 310
rect -184 244 184 284
rect -184 218 -178 244
rect -152 218 -112 244
rect -86 218 -46 244
rect -20 218 20 244
rect 46 218 86 244
rect 112 218 152 244
rect 178 218 184 244
rect -184 178 184 218
rect -184 152 -178 178
rect -152 152 -112 178
rect -86 152 -46 178
rect -20 152 20 178
rect 46 152 86 178
rect 112 152 152 178
rect 178 152 184 178
rect -184 112 184 152
rect -184 86 -178 112
rect -152 86 -112 112
rect -86 86 -46 112
rect -20 86 20 112
rect 46 86 86 112
rect 112 86 152 112
rect 178 86 184 112
rect -184 46 184 86
rect -184 20 -178 46
rect -152 20 -112 46
rect -86 20 -46 46
rect -20 20 20 46
rect 46 20 86 46
rect 112 20 152 46
rect 178 20 184 46
rect -184 -20 184 20
rect -184 -46 -178 -20
rect -152 -46 -112 -20
rect -86 -46 -46 -20
rect -20 -46 20 -20
rect 46 -46 86 -20
rect 112 -46 152 -20
rect 178 -46 184 -20
rect -184 -86 184 -46
rect -184 -112 -178 -86
rect -152 -112 -112 -86
rect -86 -112 -46 -86
rect -20 -112 20 -86
rect 46 -112 86 -86
rect 112 -112 152 -86
rect 178 -112 184 -86
rect -184 -152 184 -112
rect -184 -178 -178 -152
rect -152 -178 -112 -152
rect -86 -178 -46 -152
rect -20 -178 20 -152
rect 46 -178 86 -152
rect 112 -178 152 -152
rect 178 -178 184 -152
rect -184 -218 184 -178
rect -184 -244 -178 -218
rect -152 -244 -112 -218
rect -86 -244 -46 -218
rect -20 -244 20 -218
rect 46 -244 86 -218
rect 112 -244 152 -218
rect 178 -244 184 -218
rect -184 -284 184 -244
rect -184 -310 -178 -284
rect -152 -310 -112 -284
rect -86 -310 -46 -284
rect -20 -310 20 -284
rect 46 -310 86 -284
rect 112 -310 152 -284
rect 178 -310 184 -284
rect -184 -350 184 -310
rect -184 -376 -178 -350
rect -152 -376 -112 -350
rect -86 -376 -46 -350
rect -20 -376 20 -350
rect 46 -376 86 -350
rect 112 -376 152 -350
rect 178 -376 184 -350
rect -184 -416 184 -376
rect -184 -442 -178 -416
rect -152 -442 -112 -416
rect -86 -442 -46 -416
rect -20 -442 20 -416
rect 46 -442 86 -416
rect 112 -442 152 -416
rect 178 -442 184 -416
rect -184 -482 184 -442
rect -184 -508 -178 -482
rect -152 -508 -112 -482
rect -86 -508 -46 -482
rect -20 -508 20 -482
rect 46 -508 86 -482
rect 112 -508 152 -482
rect 178 -508 184 -482
rect -184 -548 184 -508
rect -184 -574 -178 -548
rect -152 -574 -112 -548
rect -86 -574 -46 -548
rect -20 -574 20 -548
rect 46 -574 86 -548
rect 112 -574 152 -548
rect 178 -574 184 -548
rect -184 -580 184 -574
<< via1 >>
rect -178 548 -152 574
rect -112 548 -86 574
rect -46 548 -20 574
rect 20 548 46 574
rect 86 548 112 574
rect 152 548 178 574
rect -178 482 -152 508
rect -112 482 -86 508
rect -46 482 -20 508
rect 20 482 46 508
rect 86 482 112 508
rect 152 482 178 508
rect -178 416 -152 442
rect -112 416 -86 442
rect -46 416 -20 442
rect 20 416 46 442
rect 86 416 112 442
rect 152 416 178 442
rect -178 350 -152 376
rect -112 350 -86 376
rect -46 350 -20 376
rect 20 350 46 376
rect 86 350 112 376
rect 152 350 178 376
rect -178 284 -152 310
rect -112 284 -86 310
rect -46 284 -20 310
rect 20 284 46 310
rect 86 284 112 310
rect 152 284 178 310
rect -178 218 -152 244
rect -112 218 -86 244
rect -46 218 -20 244
rect 20 218 46 244
rect 86 218 112 244
rect 152 218 178 244
rect -178 152 -152 178
rect -112 152 -86 178
rect -46 152 -20 178
rect 20 152 46 178
rect 86 152 112 178
rect 152 152 178 178
rect -178 86 -152 112
rect -112 86 -86 112
rect -46 86 -20 112
rect 20 86 46 112
rect 86 86 112 112
rect 152 86 178 112
rect -178 20 -152 46
rect -112 20 -86 46
rect -46 20 -20 46
rect 20 20 46 46
rect 86 20 112 46
rect 152 20 178 46
rect -178 -46 -152 -20
rect -112 -46 -86 -20
rect -46 -46 -20 -20
rect 20 -46 46 -20
rect 86 -46 112 -20
rect 152 -46 178 -20
rect -178 -112 -152 -86
rect -112 -112 -86 -86
rect -46 -112 -20 -86
rect 20 -112 46 -86
rect 86 -112 112 -86
rect 152 -112 178 -86
rect -178 -178 -152 -152
rect -112 -178 -86 -152
rect -46 -178 -20 -152
rect 20 -178 46 -152
rect 86 -178 112 -152
rect 152 -178 178 -152
rect -178 -244 -152 -218
rect -112 -244 -86 -218
rect -46 -244 -20 -218
rect 20 -244 46 -218
rect 86 -244 112 -218
rect 152 -244 178 -218
rect -178 -310 -152 -284
rect -112 -310 -86 -284
rect -46 -310 -20 -284
rect 20 -310 46 -284
rect 86 -310 112 -284
rect 152 -310 178 -284
rect -178 -376 -152 -350
rect -112 -376 -86 -350
rect -46 -376 -20 -350
rect 20 -376 46 -350
rect 86 -376 112 -350
rect 152 -376 178 -350
rect -178 -442 -152 -416
rect -112 -442 -86 -416
rect -46 -442 -20 -416
rect 20 -442 46 -416
rect 86 -442 112 -416
rect 152 -442 178 -416
rect -178 -508 -152 -482
rect -112 -508 -86 -482
rect -46 -508 -20 -482
rect 20 -508 46 -482
rect 86 -508 112 -482
rect 152 -508 178 -482
rect -178 -574 -152 -548
rect -112 -574 -86 -548
rect -46 -574 -20 -548
rect 20 -574 46 -548
rect 86 -574 112 -548
rect 152 -574 178 -548
<< metal2 >>
rect -184 574 184 580
rect -184 548 -178 574
rect -152 548 -112 574
rect -86 548 -46 574
rect -20 548 20 574
rect 46 548 86 574
rect 112 548 152 574
rect 178 548 184 574
rect -184 508 184 548
rect -184 482 -178 508
rect -152 482 -112 508
rect -86 482 -46 508
rect -20 482 20 508
rect 46 482 86 508
rect 112 482 152 508
rect 178 482 184 508
rect -184 442 184 482
rect -184 416 -178 442
rect -152 416 -112 442
rect -86 416 -46 442
rect -20 416 20 442
rect 46 416 86 442
rect 112 416 152 442
rect 178 416 184 442
rect -184 376 184 416
rect -184 350 -178 376
rect -152 350 -112 376
rect -86 350 -46 376
rect -20 350 20 376
rect 46 350 86 376
rect 112 350 152 376
rect 178 350 184 376
rect -184 310 184 350
rect -184 284 -178 310
rect -152 284 -112 310
rect -86 284 -46 310
rect -20 284 20 310
rect 46 284 86 310
rect 112 284 152 310
rect 178 284 184 310
rect -184 244 184 284
rect -184 218 -178 244
rect -152 218 -112 244
rect -86 218 -46 244
rect -20 218 20 244
rect 46 218 86 244
rect 112 218 152 244
rect 178 218 184 244
rect -184 178 184 218
rect -184 152 -178 178
rect -152 152 -112 178
rect -86 152 -46 178
rect -20 152 20 178
rect 46 152 86 178
rect 112 152 152 178
rect 178 152 184 178
rect -184 112 184 152
rect -184 86 -178 112
rect -152 86 -112 112
rect -86 86 -46 112
rect -20 86 20 112
rect 46 86 86 112
rect 112 86 152 112
rect 178 86 184 112
rect -184 46 184 86
rect -184 20 -178 46
rect -152 20 -112 46
rect -86 20 -46 46
rect -20 20 20 46
rect 46 20 86 46
rect 112 20 152 46
rect 178 20 184 46
rect -184 -20 184 20
rect -184 -46 -178 -20
rect -152 -46 -112 -20
rect -86 -46 -46 -20
rect -20 -46 20 -20
rect 46 -46 86 -20
rect 112 -46 152 -20
rect 178 -46 184 -20
rect -184 -86 184 -46
rect -184 -112 -178 -86
rect -152 -112 -112 -86
rect -86 -112 -46 -86
rect -20 -112 20 -86
rect 46 -112 86 -86
rect 112 -112 152 -86
rect 178 -112 184 -86
rect -184 -152 184 -112
rect -184 -178 -178 -152
rect -152 -178 -112 -152
rect -86 -178 -46 -152
rect -20 -178 20 -152
rect 46 -178 86 -152
rect 112 -178 152 -152
rect 178 -178 184 -152
rect -184 -218 184 -178
rect -184 -244 -178 -218
rect -152 -244 -112 -218
rect -86 -244 -46 -218
rect -20 -244 20 -218
rect 46 -244 86 -218
rect 112 -244 152 -218
rect 178 -244 184 -218
rect -184 -284 184 -244
rect -184 -310 -178 -284
rect -152 -310 -112 -284
rect -86 -310 -46 -284
rect -20 -310 20 -284
rect 46 -310 86 -284
rect 112 -310 152 -284
rect 178 -310 184 -284
rect -184 -350 184 -310
rect -184 -376 -178 -350
rect -152 -376 -112 -350
rect -86 -376 -46 -350
rect -20 -376 20 -350
rect 46 -376 86 -350
rect 112 -376 152 -350
rect 178 -376 184 -350
rect -184 -416 184 -376
rect -184 -442 -178 -416
rect -152 -442 -112 -416
rect -86 -442 -46 -416
rect -20 -442 20 -416
rect 46 -442 86 -416
rect 112 -442 152 -416
rect 178 -442 184 -416
rect -184 -482 184 -442
rect -184 -508 -178 -482
rect -152 -508 -112 -482
rect -86 -508 -46 -482
rect -20 -508 20 -482
rect 46 -508 86 -482
rect 112 -508 152 -482
rect 178 -508 184 -482
rect -184 -548 184 -508
rect -184 -574 -178 -548
rect -152 -574 -112 -548
rect -86 -574 -46 -548
rect -20 -574 20 -548
rect 46 -574 86 -548
rect 112 -574 152 -548
rect 178 -574 184 -548
rect -184 -580 184 -574
<< end >>
