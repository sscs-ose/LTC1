magic
tech gf180mcuC
magscale 1 10
timestamp 1693309239
<< psubdiff >>
rect 0 1259 6715 1285
rect 0 1128 48 1259
rect 193 1128 348 1259
rect 493 1128 648 1259
rect 793 1128 948 1259
rect 1093 1128 1248 1259
rect 1393 1128 1548 1259
rect 1693 1128 1848 1259
rect 1993 1128 2148 1259
rect 2293 1128 2448 1259
rect 2593 1128 2748 1259
rect 2893 1128 3048 1259
rect 3193 1128 3348 1259
rect 3493 1128 3648 1259
rect 3793 1128 3948 1259
rect 4093 1128 4248 1259
rect 4393 1128 4548 1259
rect 4693 1128 4848 1259
rect 4993 1128 5148 1259
rect 5293 1128 5448 1259
rect 5593 1128 5748 1259
rect 5893 1128 6048 1259
rect 6193 1128 6348 1259
rect 6493 1128 6715 1259
rect 0 1098 6715 1128
rect 0 -50 6715 -21
rect 0 -181 44 -50
rect 189 -181 344 -50
rect 489 -181 644 -50
rect 789 -181 944 -50
rect 1089 -181 1244 -50
rect 1389 -181 1544 -50
rect 1689 -181 1844 -50
rect 1989 -181 2144 -50
rect 2289 -181 2444 -50
rect 2589 -181 2744 -50
rect 2889 -181 3044 -50
rect 3189 -181 3344 -50
rect 3489 -181 3644 -50
rect 3789 -181 3944 -50
rect 4089 -181 4244 -50
rect 4389 -181 4544 -50
rect 4689 -181 4844 -50
rect 4989 -181 5144 -50
rect 5289 -181 5444 -50
rect 5589 -181 5744 -50
rect 5889 -181 6044 -50
rect 6189 -181 6344 -50
rect 6489 -181 6715 -50
rect 0 -208 6715 -181
<< psubdiffcont >>
rect 48 1128 193 1259
rect 348 1128 493 1259
rect 648 1128 793 1259
rect 948 1128 1093 1259
rect 1248 1128 1393 1259
rect 1548 1128 1693 1259
rect 1848 1128 1993 1259
rect 2148 1128 2293 1259
rect 2448 1128 2593 1259
rect 2748 1128 2893 1259
rect 3048 1128 3193 1259
rect 3348 1128 3493 1259
rect 3648 1128 3793 1259
rect 3948 1128 4093 1259
rect 4248 1128 4393 1259
rect 4548 1128 4693 1259
rect 4848 1128 4993 1259
rect 5148 1128 5293 1259
rect 5448 1128 5593 1259
rect 5748 1128 5893 1259
rect 6048 1128 6193 1259
rect 6348 1128 6493 1259
rect 44 -181 189 -50
rect 344 -181 489 -50
rect 644 -181 789 -50
rect 944 -181 1089 -50
rect 1244 -181 1389 -50
rect 1544 -181 1689 -50
rect 1844 -181 1989 -50
rect 2144 -181 2289 -50
rect 2444 -181 2589 -50
rect 2744 -181 2889 -50
rect 3044 -181 3189 -50
rect 3344 -181 3489 -50
rect 3644 -181 3789 -50
rect 3944 -181 4089 -50
rect 4244 -181 4389 -50
rect 4544 -181 4689 -50
rect 4844 -181 4989 -50
rect 5144 -181 5289 -50
rect 5444 -181 5589 -50
rect 5744 -181 5889 -50
rect 6044 -181 6189 -50
rect 6344 -181 6489 -50
<< polysilicon >>
rect -168 1077 -82 1091
rect -168 1073 6536 1077
rect -168 1024 -150 1073
rect -102 1024 6536 1073
rect -168 1019 6536 1024
rect -168 1008 -82 1019
rect 112 925 212 1019
rect 724 936 824 1019
rect 928 936 1028 1019
rect 1540 936 1640 1019
rect 1744 936 1844 1019
rect 2356 936 2456 1019
rect 2560 936 2660 1019
rect 3172 936 3272 1019
rect 3376 936 3476 1019
rect 3988 936 4088 1019
rect 4192 936 4292 1019
rect 4804 936 4904 1019
rect 5008 936 5108 1019
rect 5620 936 5720 1019
rect 5824 936 5924 1019
rect 6436 936 6536 1019
rect -171 553 -84 566
rect 316 553 416 608
rect 520 553 620 608
rect 1132 553 1232 608
rect 1336 553 1436 608
rect 1948 553 2048 608
rect 2152 553 2252 608
rect 2764 553 2864 608
rect 2968 553 3068 608
rect 3580 553 3680 608
rect 3784 553 3884 608
rect 4396 553 4496 608
rect 4600 553 4700 608
rect 5212 553 5312 608
rect 5416 553 5516 608
rect 6028 553 6128 608
rect 6232 553 6332 608
rect -171 552 6536 553
rect -171 499 -158 552
rect -102 499 6536 552
rect -171 494 6536 499
rect -171 485 -84 494
rect 112 401 212 494
rect 724 445 824 494
rect 928 445 1028 494
rect 1540 445 1640 494
rect 1744 445 1844 494
rect 2356 445 2456 494
rect 2560 445 2660 494
rect 3172 445 3272 494
rect 3376 445 3476 494
rect 3988 445 4088 494
rect 4192 445 4292 494
rect 4804 445 4904 494
rect 5008 445 5108 494
rect 5620 445 5720 494
rect 5824 445 5924 494
rect 6436 445 6536 494
rect -166 58 -74 74
rect 316 58 416 129
rect 520 58 620 117
rect 1132 58 1232 117
rect 1336 58 1436 117
rect 1948 58 2048 117
rect 2152 58 2252 117
rect 2764 58 2864 117
rect 2968 58 3068 117
rect 3580 58 3680 117
rect 3784 58 3884 117
rect 4396 58 4496 117
rect 4600 58 4700 117
rect 5212 58 5312 117
rect 5416 58 5516 117
rect 6028 58 6128 117
rect 6232 58 6332 117
rect -166 53 6332 58
rect -166 2 -150 53
rect -102 2 6332 53
rect -166 -1 6332 2
rect -166 -14 -74 -1
<< polycontact >>
rect -150 1024 -102 1073
rect -158 499 -102 552
rect -150 2 -102 53
<< metal1 >>
rect 0 1259 6715 1285
rect 0 1128 48 1259
rect 193 1128 348 1259
rect 493 1128 648 1259
rect 793 1128 948 1259
rect 1093 1128 1248 1259
rect 1393 1128 1548 1259
rect 1693 1128 1848 1259
rect 1993 1128 2148 1259
rect 2293 1128 2448 1259
rect 2593 1128 2748 1259
rect 2893 1128 3048 1259
rect 3193 1128 3348 1259
rect 3493 1128 3648 1259
rect 3793 1128 3948 1259
rect 4093 1128 4248 1259
rect 4393 1128 4548 1259
rect 4693 1128 4848 1259
rect 4993 1128 5148 1259
rect 5293 1128 5448 1259
rect 5593 1128 5748 1259
rect 5893 1128 6048 1259
rect 6193 1128 6348 1259
rect 6493 1230 6715 1259
rect 6493 1158 6567 1230
rect 6656 1158 6715 1230
rect 6493 1128 6715 1158
rect 0 1098 6715 1128
rect -168 1076 -82 1091
rect -168 1020 -155 1076
rect -99 1020 -82 1076
rect -168 1008 -82 1020
rect 445 890 491 1098
rect 1261 890 1307 1098
rect 2077 890 2123 1098
rect 2893 890 2939 1098
rect 3709 890 3755 1098
rect 4525 890 4571 1098
rect 5341 890 5387 1098
rect 6157 890 6203 1098
rect 219 826 304 843
rect 219 766 233 826
rect 290 766 304 826
rect 219 752 304 766
rect 632 830 717 844
rect 632 771 647 830
rect 702 771 717 830
rect 632 753 717 771
rect 1044 824 1129 838
rect 1044 765 1059 824
rect 1114 765 1129 824
rect 1044 748 1129 765
rect 1444 830 1529 844
rect 1444 771 1459 830
rect 1514 771 1529 830
rect 1444 753 1529 771
rect 1857 812 1942 826
rect 1857 753 1872 812
rect 1927 753 1942 812
rect 1857 735 1942 753
rect 2267 823 2352 837
rect 2267 764 2282 823
rect 2337 764 2352 823
rect 2267 746 2352 764
rect 2664 812 2749 826
rect 2664 753 2679 812
rect 2734 753 2749 812
rect 2664 735 2749 753
rect 3079 817 3164 831
rect 3079 758 3094 817
rect 3149 758 3164 817
rect 3079 740 3164 758
rect 3490 820 3575 834
rect 3490 761 3505 820
rect 3560 761 3575 820
rect 3490 743 3575 761
rect 3900 830 3985 844
rect 3900 771 3915 830
rect 3970 771 3985 830
rect 3900 753 3985 771
rect 4305 812 4390 826
rect 4305 753 4320 812
rect 4375 753 4390 812
rect 4305 735 4390 753
rect 4707 812 4792 826
rect 4707 753 4722 812
rect 4777 753 4792 812
rect 4707 735 4792 753
rect 5123 825 5208 839
rect 5123 766 5138 825
rect 5193 766 5208 825
rect 5123 748 5208 766
rect 5523 817 5608 831
rect 5523 758 5538 817
rect 5593 758 5608 817
rect 5523 740 5608 758
rect 5940 814 6025 828
rect 5940 755 5955 814
rect 6010 755 6025 814
rect 5940 737 6025 755
rect 6328 820 6413 834
rect 6328 761 6343 820
rect 6398 761 6413 820
rect 6328 743 6413 761
rect 37 591 83 654
rect 853 591 899 654
rect 1669 591 1715 654
rect 2485 591 2531 654
rect 3301 591 3347 654
rect 4117 591 4163 654
rect 4933 591 4979 654
rect 5749 591 5795 654
rect 6565 591 6611 654
rect -171 552 -84 566
rect -171 499 -158 552
rect -102 499 -84 552
rect 37 519 6915 591
rect -171 485 -84 499
rect 445 399 491 519
rect 1261 399 1307 519
rect 2077 399 2123 519
rect 2893 399 2939 519
rect 3709 399 3755 519
rect 4525 399 4571 519
rect 5341 399 5387 519
rect 6157 399 6203 519
rect 1038 342 1123 356
rect 221 321 306 338
rect 221 262 235 321
rect 290 262 306 321
rect 221 247 306 262
rect 642 326 727 340
rect 642 267 657 326
rect 712 267 727 326
rect 642 249 727 267
rect 1038 283 1053 342
rect 1108 283 1123 342
rect 1038 265 1123 283
rect 1451 347 1536 361
rect 1451 288 1466 347
rect 1521 288 1536 347
rect 1451 270 1536 288
rect 1851 345 1936 359
rect 1851 286 1866 345
rect 1921 286 1936 345
rect 1851 268 1936 286
rect 2254 335 2339 349
rect 2254 276 2269 335
rect 2324 276 2339 335
rect 2254 258 2339 276
rect 2677 337 2762 351
rect 2677 278 2692 337
rect 2747 278 2762 337
rect 3486 336 3562 338
rect 3892 337 3977 351
rect 2677 260 2762 278
rect 3077 321 3162 335
rect 3077 262 3092 321
rect 3147 262 3162 321
rect 3077 244 3162 262
rect 3479 322 3564 336
rect 3479 263 3494 322
rect 3549 263 3564 322
rect 3479 245 3564 263
rect 3892 278 3907 337
rect 3962 278 3977 337
rect 3892 260 3977 278
rect 4295 306 4380 320
rect 4295 247 4310 306
rect 4365 247 4380 306
rect 4295 229 4380 247
rect 4712 316 4797 330
rect 4712 257 4727 316
rect 4782 257 4797 316
rect 4712 239 4797 257
rect 5120 329 5205 343
rect 5120 270 5135 329
rect 5190 270 5205 329
rect 5120 252 5205 270
rect 5520 331 5605 345
rect 5520 272 5535 331
rect 5590 272 5605 331
rect 5520 254 5605 272
rect 5935 332 6020 346
rect 5935 273 5950 332
rect 6005 273 6020 332
rect 5935 255 6020 273
rect 6343 319 6428 333
rect 6343 260 6358 319
rect 6413 260 6428 319
rect 6343 242 6428 260
rect -166 58 -74 74
rect -166 1 -151 58
rect -94 1 -74 58
rect -166 -14 -74 1
rect 37 -21 83 163
rect 853 -21 899 163
rect 1669 -21 1715 163
rect 2485 -21 2531 163
rect 3301 -21 3347 163
rect 4117 -21 4163 163
rect 4933 -21 4979 163
rect 5749 -21 5795 163
rect 6565 -21 6611 163
rect 0 -50 6715 -21
rect 0 -181 44 -50
rect 189 -181 344 -50
rect 489 -181 644 -50
rect 789 -181 944 -50
rect 1089 -181 1244 -50
rect 1389 -181 1544 -50
rect 1689 -181 1844 -50
rect 1989 -181 2144 -50
rect 2289 -181 2444 -50
rect 2589 -181 2744 -50
rect 2889 -181 3044 -50
rect 3189 -181 3344 -50
rect 3489 -181 3644 -50
rect 3789 -181 3944 -50
rect 4089 -181 4244 -50
rect 4389 -181 4544 -50
rect 4689 -181 4844 -50
rect 4989 -181 5144 -50
rect 5289 -181 5444 -50
rect 5589 -181 5744 -50
rect 5889 -181 6044 -50
rect 6189 -181 6344 -50
rect 6489 -86 6715 -50
rect 6489 -153 6581 -86
rect 6648 -153 6715 -86
rect 6489 -181 6715 -153
rect 0 -208 6715 -181
<< via1 >>
rect 6567 1158 6656 1230
rect -155 1073 -99 1076
rect -155 1024 -150 1073
rect -150 1024 -102 1073
rect -102 1024 -99 1073
rect -155 1020 -99 1024
rect 233 766 290 826
rect 647 771 702 830
rect 1059 765 1114 824
rect 1459 771 1514 830
rect 1872 753 1927 812
rect 2282 764 2337 823
rect 2679 753 2734 812
rect 3094 758 3149 817
rect 3505 761 3560 820
rect 3915 771 3970 830
rect 4320 753 4375 812
rect 4722 753 4777 812
rect 5138 766 5193 825
rect 5538 758 5593 817
rect 5955 755 6010 814
rect 6343 761 6398 820
rect 235 262 290 321
rect 657 267 712 326
rect 1053 283 1108 342
rect 1466 288 1521 347
rect 1866 286 1921 345
rect 2269 276 2324 335
rect 2692 278 2747 337
rect 3092 262 3147 321
rect 3494 263 3549 322
rect 3907 278 3962 337
rect 4310 247 4365 306
rect 4727 257 4782 316
rect 5135 270 5190 329
rect 5535 272 5590 331
rect 5950 273 6005 332
rect 6358 260 6413 319
rect -151 53 -94 58
rect -151 2 -150 53
rect -150 2 -102 53
rect -102 2 -94 53
rect -151 1 -94 2
rect 6581 -153 6648 -86
<< metal2 >>
rect 6547 1230 6686 1257
rect 6547 1158 6567 1230
rect 6656 1158 6686 1230
rect 6547 1133 6686 1158
rect -168 1076 -82 1091
rect -168 1020 -155 1076
rect -99 1020 -82 1076
rect -168 1008 -82 1020
rect -156 74 -98 1008
rect 219 826 304 843
rect 219 766 233 826
rect 290 766 304 826
rect 219 752 304 766
rect 632 830 717 844
rect 632 771 647 830
rect 702 771 717 830
rect 632 753 717 771
rect 1044 824 1129 838
rect 1044 765 1059 824
rect 1114 765 1129 824
rect 233 338 290 752
rect 650 340 707 753
rect 1044 748 1129 765
rect 1444 830 1529 844
rect 1444 771 1459 830
rect 1514 771 1529 830
rect 1444 753 1529 771
rect 1857 812 1942 826
rect 1857 753 1872 812
rect 1927 753 1942 812
rect 1058 356 1115 748
rect 1459 361 1516 753
rect 1857 735 1942 753
rect 2267 823 2352 837
rect 2267 764 2282 823
rect 2337 764 2352 823
rect 2267 746 2352 764
rect 2664 812 2749 826
rect 2664 753 2679 812
rect 2734 753 2749 812
rect 1038 342 1123 356
rect 221 336 306 338
rect 642 336 727 340
rect 1038 336 1053 342
rect 221 326 1053 336
rect 221 321 657 326
rect 221 262 235 321
rect 290 279 657 321
rect 290 262 306 279
rect 221 247 306 262
rect 642 267 657 279
rect 712 283 1053 326
rect 1108 336 1123 342
rect 1451 347 1536 361
rect 1867 359 1924 735
rect 1451 336 1466 347
rect 1108 288 1466 336
rect 1521 336 1536 347
rect 1851 345 1936 359
rect 2270 349 2327 746
rect 2664 735 2749 753
rect 3079 817 3164 831
rect 3079 758 3094 817
rect 3149 758 3164 817
rect 3079 740 3164 758
rect 3490 820 3575 834
rect 3490 761 3505 820
rect 3560 761 3575 820
rect 3490 743 3575 761
rect 3900 830 3985 844
rect 3900 771 3915 830
rect 3970 771 3985 830
rect 3900 753 3985 771
rect 4305 812 4390 826
rect 4305 753 4320 812
rect 4375 753 4390 812
rect 2684 351 2741 735
rect 1851 336 1866 345
rect 1521 288 1866 336
rect 1108 286 1866 288
rect 1921 336 1936 345
rect 2254 336 2339 349
rect 2677 337 2762 351
rect 2677 336 2692 337
rect 1921 335 2692 336
rect 1921 286 2269 335
rect 1108 283 2269 286
rect 712 279 2269 283
rect 712 267 727 279
rect 642 249 727 267
rect 1038 265 1123 279
rect 1451 270 1536 279
rect 1851 268 1936 279
rect 2254 276 2269 279
rect 2324 279 2692 335
rect 2324 276 2339 279
rect 2254 258 2339 276
rect 2677 278 2692 279
rect 2747 336 2762 337
rect 3093 336 3150 740
rect 3495 336 3552 743
rect 3909 351 3966 753
rect 4305 735 4390 753
rect 4707 812 4792 826
rect 4707 753 4722 812
rect 4777 753 4792 812
rect 4707 735 4792 753
rect 5123 825 5208 839
rect 5123 766 5138 825
rect 5193 766 5208 825
rect 5123 748 5208 766
rect 5523 817 5608 831
rect 5523 758 5538 817
rect 5593 758 5608 817
rect 3892 337 3977 351
rect 3892 336 3907 337
rect 2747 322 3907 336
rect 2747 321 3494 322
rect 2747 279 3092 321
rect 2747 278 2762 279
rect 2677 260 2762 278
rect 3077 262 3092 279
rect 3147 279 3494 321
rect 3147 262 3162 279
rect 3077 244 3162 262
rect 3479 263 3494 279
rect 3549 279 3907 322
rect 3549 263 3564 279
rect 3479 245 3564 263
rect 3892 278 3907 279
rect 3962 336 3977 337
rect 4311 336 4368 735
rect 4719 336 4776 735
rect 5128 343 5185 748
rect 5523 740 5608 758
rect 5940 814 6025 828
rect 5940 755 5955 814
rect 6010 755 6025 814
rect 5526 345 5583 740
rect 5940 737 6025 755
rect 6328 820 6413 834
rect 6328 761 6343 820
rect 6398 761 6413 820
rect 6328 743 6413 761
rect 5942 346 5999 737
rect 5120 336 5205 343
rect 5520 336 5605 345
rect 5935 336 6020 346
rect 6345 336 6402 743
rect 3962 333 6402 336
rect 3962 332 6428 333
rect 3962 331 5950 332
rect 3962 329 5535 331
rect 3962 316 5135 329
rect 3962 306 4727 316
rect 3962 279 4310 306
rect 3962 278 3977 279
rect 3892 260 3977 278
rect 4295 247 4310 279
rect 4365 279 4727 306
rect 4365 247 4380 279
rect 4295 229 4380 247
rect 4712 257 4727 279
rect 4782 279 5135 316
rect 4782 257 4797 279
rect 4712 239 4797 257
rect 5120 270 5135 279
rect 5190 279 5535 329
rect 5190 270 5205 279
rect 5120 252 5205 270
rect 5520 272 5535 279
rect 5590 279 5950 331
rect 5590 272 5605 279
rect 5520 254 5605 272
rect 5935 273 5950 279
rect 6005 319 6428 332
rect 6005 279 6358 319
rect 6005 273 6020 279
rect 5935 255 6020 273
rect 6343 260 6358 279
rect 6413 260 6428 319
rect 6343 242 6428 260
rect -166 58 -74 74
rect -166 1 -151 58
rect -94 1 -74 58
rect -166 -14 -74 1
rect 6581 -75 6648 1133
rect 6564 -86 6667 -75
rect 6564 -153 6581 -86
rect 6648 -153 6667 -86
rect 6564 -168 6667 -153
use nmos_3p3_LNPLVM  nmos_3p3_LNPLVM_0
timestamp 1693309239
transform 1 0 3324 0 1 772
box -3324 -188 3324 188
use nmos_3p3_LNPLVM  nmos_3p3_LNPLVM_1
timestamp 1693309239
transform 1 0 3324 0 1 281
box -3324 -188 3324 188
<< labels >>
flabel via1 -133 1049 -133 1049 0 FreeSans 1600 0 0 0 IM_T
port 0 nsew
flabel metal1 1480 1192 1480 1192 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 6857 556 6857 556 0 FreeSans 1600 0 0 0 OUT
port 3 nsew
flabel metal1 -164 520 -164 520 0 FreeSans 1600 0 0 0 IM
port 4 nsew
flabel via1 2290 310 2290 310 0 FreeSans 1600 0 0 0 SD
port 5 nsew
<< end >>
