magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2747 -2051 15709 27617
<< polysilicon >>
rect 1237 23733 1437 23873
rect 11525 23733 11725 23873
rect 1421 23489 1437 23629
rect 11525 23489 11541 23629
rect 1421 23245 1437 23385
rect 11525 23245 11541 23385
rect 1421 23001 1437 23141
rect 11525 23001 11541 23141
rect 1421 22757 1437 22897
rect 11525 22757 11541 22897
rect 1421 22513 1437 22653
rect 11525 22513 11541 22653
rect 1421 22269 1437 22409
rect 11525 22269 11541 22409
rect 1421 22025 1437 22165
rect 11525 22025 11541 22165
rect 1421 21781 1437 21921
rect 11525 21781 11541 21921
rect 1421 21537 1437 21677
rect 11525 21537 11541 21677
rect 1421 21293 1437 21433
rect 11525 21293 11541 21433
rect 1421 21049 1437 21189
rect 11525 21049 11541 21189
rect 1421 20805 1437 20945
rect 11525 20805 11541 20945
rect 1421 20561 1437 20701
rect 11525 20561 11541 20701
rect 1421 20317 1437 20457
rect 11525 20317 11541 20457
rect 1421 20073 1437 20213
rect 11525 20073 11541 20213
rect 1421 19829 1437 19969
rect 11525 19829 11541 19969
rect 1421 19585 1437 19725
rect 11525 19585 11541 19725
rect 1421 19341 1437 19481
rect 11525 19341 11541 19481
rect 1237 19097 1437 19237
rect 11525 19097 11725 19237
rect 1237 17861 1437 18001
rect 11525 17861 11725 18001
rect 1421 17617 1437 17757
rect 11525 17617 11541 17757
rect 1421 17373 1437 17513
rect 11525 17373 11541 17513
rect 1421 17129 1437 17269
rect 11525 17129 11541 17269
rect 1421 16885 1437 17025
rect 11525 16885 11541 17025
rect 1421 16641 1437 16781
rect 11525 16641 11541 16781
rect 1421 16397 1437 16537
rect 11525 16397 11541 16537
rect 1421 16153 1437 16293
rect 11525 16153 11541 16293
rect 1421 15909 1437 16049
rect 11525 15909 11541 16049
rect 1421 15665 1437 15805
rect 11525 15665 11541 15805
rect 1421 15421 1437 15561
rect 11525 15421 11541 15561
rect 1421 15177 1437 15317
rect 11525 15177 11541 15317
rect 1421 14933 1437 15073
rect 11525 14933 11541 15073
rect 1421 14689 1437 14829
rect 11525 14689 11541 14829
rect 1421 14445 1437 14585
rect 11525 14445 11541 14585
rect 1421 14201 1437 14341
rect 11525 14201 11541 14341
rect 1421 13957 1437 14097
rect 11525 13957 11541 14097
rect 1421 13713 1437 13853
rect 11525 13713 11541 13853
rect 1421 13469 1437 13609
rect 11525 13469 11541 13609
rect 1237 13225 1437 13365
rect 11525 13225 11725 13365
rect 1237 11989 1437 12129
rect 11525 11989 11725 12129
rect 1421 11745 1437 11885
rect 11525 11745 11541 11885
rect 1421 11501 1437 11641
rect 11525 11501 11541 11641
rect 1421 11257 1437 11397
rect 11525 11257 11541 11397
rect 1421 11013 1437 11153
rect 11525 11013 11541 11153
rect 1421 10769 1437 10909
rect 11525 10769 11541 10909
rect 1421 10525 1437 10665
rect 11525 10525 11541 10665
rect 1421 10281 1437 10421
rect 11525 10281 11541 10421
rect 1421 10037 1437 10177
rect 11525 10037 11541 10177
rect 1421 9793 1437 9933
rect 11525 9793 11541 9933
rect 1421 9549 1437 9689
rect 11525 9549 11541 9689
rect 1421 9305 1437 9445
rect 11525 9305 11541 9445
rect 1421 9061 1437 9201
rect 11525 9061 11541 9201
rect 1421 8817 1437 8957
rect 11525 8817 11541 8957
rect 1421 8573 1437 8713
rect 11525 8573 11541 8713
rect 1421 8329 1437 8469
rect 11525 8329 11541 8469
rect 1421 8085 1437 8225
rect 11525 8085 11541 8225
rect 1421 7841 1437 7981
rect 11525 7841 11541 7981
rect 1421 7597 1437 7737
rect 11525 7597 11541 7737
rect 1237 7353 1437 7493
rect 11525 7353 11725 7493
rect 1237 6117 1437 6257
rect 11525 6117 11725 6257
rect 1421 5873 1437 6013
rect 11525 5873 11541 6013
rect 1421 5629 1437 5769
rect 11525 5629 11541 5769
rect 1421 5385 1437 5525
rect 11525 5385 11541 5525
rect 1421 5141 1437 5281
rect 11525 5141 11541 5281
rect 1421 4897 1437 5037
rect 11525 4897 11541 5037
rect 1421 4653 1437 4793
rect 11525 4653 11541 4793
rect 1421 4409 1437 4549
rect 11525 4409 11541 4549
rect 1421 4165 1437 4305
rect 11525 4165 11541 4305
rect 1421 3921 1437 4061
rect 11525 3921 11541 4061
rect 1421 3677 1437 3817
rect 11525 3677 11541 3817
rect 1421 3433 1437 3573
rect 11525 3433 11541 3573
rect 1421 3189 1437 3329
rect 11525 3189 11541 3329
rect 1421 2945 1437 3085
rect 11525 2945 11541 3085
rect 1421 2701 1437 2841
rect 11525 2701 11541 2841
rect 1421 2457 1437 2597
rect 11525 2457 11541 2597
rect 1421 2213 1437 2353
rect 11525 2213 11541 2353
rect 1421 1969 1437 2109
rect 11525 1969 11541 2109
rect 1421 1725 1437 1865
rect 11525 1725 11541 1865
rect 1237 1481 1437 1621
rect 11525 1481 11725 1621
<< metal1 >>
rect 411 24943 497 25311
rect 12465 24943 12551 25311
rect 961 24343 1047 24711
rect 11915 24343 12001 24711
rect 1213 24053 11749 24253
rect 1213 18920 1413 24053
rect 1481 23887 11481 23963
rect 1481 23643 11481 23719
rect 1481 23399 11481 23475
rect 1481 23155 11481 23231
rect 1481 22911 11481 22987
rect 1481 22667 11481 22743
rect 1481 22423 11481 22499
rect 1481 22179 11481 22255
rect 1481 21935 11481 22011
rect 1481 21691 11481 21767
rect 1481 21447 11481 21523
rect 1481 21203 11481 21279
rect 1481 20959 11481 21035
rect 1481 20715 11481 20791
rect 1481 20471 11481 20547
rect 1481 20227 11481 20303
rect 1481 19983 11481 20059
rect 1481 19739 11481 19815
rect 1481 19495 11481 19571
rect 1481 19251 11481 19327
rect 1481 19007 11481 19083
rect 11549 18920 11749 24053
rect 1213 18720 11749 18920
rect 961 18457 12001 18641
rect 1213 18178 11749 18378
rect 1213 13048 1413 18178
rect 1481 18015 11481 18091
rect 1481 17771 11481 17847
rect 1481 17527 11481 17603
rect 1481 17283 11481 17359
rect 1481 17039 11481 17115
rect 1481 16795 11481 16871
rect 1481 16551 11481 16627
rect 1481 16307 11481 16383
rect 1481 16063 11481 16139
rect 1481 15819 11481 15895
rect 1481 15575 11481 15651
rect 1481 15331 11481 15407
rect 1481 15087 11481 15163
rect 1481 14843 11481 14919
rect 1481 14599 11481 14675
rect 1481 14355 11481 14431
rect 1481 14111 11481 14187
rect 1481 13867 11481 13943
rect 1481 13623 11481 13699
rect 1481 13379 11481 13455
rect 1481 13135 11481 13211
rect 11549 13048 11749 18178
rect 1213 12848 11749 13048
rect 961 12585 12001 12769
rect 1213 12306 11749 12506
rect 1213 7176 1413 12306
rect 1481 12143 11481 12219
rect 1481 11899 11481 11975
rect 1481 11655 11481 11731
rect 1481 11411 11481 11487
rect 1481 11167 11481 11243
rect 1481 10923 11481 10999
rect 1481 10679 11481 10755
rect 1481 10435 11481 10511
rect 1481 10191 11481 10267
rect 1481 9947 11481 10023
rect 1481 9703 11481 9779
rect 1481 9459 11481 9535
rect 1481 9215 11481 9291
rect 1481 8971 11481 9047
rect 1481 8727 11481 8803
rect 1481 8483 11481 8559
rect 1481 8239 11481 8315
rect 1481 7995 11481 8071
rect 1481 7751 11481 7827
rect 1481 7507 11481 7583
rect 1481 7263 11481 7339
rect 11549 7176 11749 12306
rect 1213 6976 11749 7176
rect 961 6713 12001 6897
rect 1213 6434 11749 6634
rect 1213 1298 1413 6434
rect 1481 6271 11481 6347
rect 1481 6027 11481 6103
rect 1481 5783 11481 5859
rect 1481 5539 11481 5615
rect 1481 5295 11481 5371
rect 1481 5051 11481 5127
rect 1481 4807 11481 4883
rect 1481 4563 11481 4639
rect 1481 4319 11481 4395
rect 1481 4075 11481 4151
rect 1481 3831 11481 3907
rect 1481 3587 11481 3663
rect 1481 3343 11481 3419
rect 1481 3099 11481 3175
rect 1481 2855 11481 2931
rect 1481 2611 11481 2687
rect 1481 2367 11481 2443
rect 1481 2123 11481 2199
rect 1481 1879 11481 1955
rect 1481 1635 11481 1711
rect 1481 1391 11481 1467
rect 11549 1298 11749 6434
rect 1213 1098 11749 1298
rect 961 643 1047 1011
rect 11915 643 12001 1011
rect 411 43 497 411
rect 12465 43 12551 411
<< metal2 >>
rect -747 43 1153 25617
rect 1213 1455 1413 25617
rect 1473 43 1673 25617
rect 1733 43 3783 25617
rect 3843 43 4043 25617
rect 4103 43 6153 25617
rect 6213 43 6749 25617
rect 6809 43 8859 25617
rect 8919 43 9119 25617
rect 9179 43 11229 25617
rect 11289 43 11489 25617
rect 11549 1455 11749 25617
rect 11809 43 13709 25617
use M1_NWELL_CDNS_40661953145131  M1_NWELL_CDNS_40661953145131_0
timestamp 1713338890
transform 1 0 12735 0 1 12677
box -278 -12728 278 12728
use M1_NWELL_CDNS_40661953145131  M1_NWELL_CDNS_40661953145131_1
timestamp 1713338890
transform 1 0 227 0 1 12677
box -278 -12728 278 12728
use M1_NWELL_CDNS_40661953145135  M1_NWELL_CDNS_40661953145135_0
timestamp 1713338890
transform 1 0 6481 0 1 227
box -6078 -278 6078 278
use M1_NWELL_CDNS_40661953145135  M1_NWELL_CDNS_40661953145135_1
timestamp 1713338890
transform 1 0 6481 0 1 25127
box -6078 -278 6078 278
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_0
timestamp 1713338890
transform 1 0 1329 0 1 3869
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_1
timestamp 1713338890
transform -1 0 11633 0 1 3869
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_2
timestamp 1713338890
transform 1 0 1329 0 1 9741
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_3
timestamp 1713338890
transform -1 0 11633 0 1 9741
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_4
timestamp 1713338890
transform 1 0 1329 0 1 15613
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_5
timestamp 1713338890
transform -1 0 11633 0 1 15613
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_6
timestamp 1713338890
transform 1 0 1329 0 1 21485
box -92 -2342 92 2342
use M1_POLY2_CDNS_69033583165361  M1_POLY2_CDNS_69033583165361_7
timestamp 1713338890
transform -1 0 11633 0 1 21485
box -92 -2342 92 2342
use M1_PSUB_CDNS_69033583165354  M1_PSUB_CDNS_69033583165354_0
timestamp 1713338890
transform 1 0 6481 0 1 827
box -5445 -195 5445 195
use M1_PSUB_CDNS_69033583165354  M1_PSUB_CDNS_69033583165354_1
timestamp 1713338890
transform 1 0 6481 0 1 24527
box -5445 -195 5445 195
use M1_PSUB_CDNS_69033583165355  M1_PSUB_CDNS_69033583165355_0
timestamp 1713338890
transform 1 0 777 0 1 12677
box -195 -12045 195 12045
use M1_PSUB_CDNS_69033583165355  M1_PSUB_CDNS_69033583165355_1
timestamp 1713338890
transform 1 0 12185 0 1 12677
box -195 -12045 195 12045
use M1_PSUB_CDNS_69033583165356  M1_PSUB_CDNS_69033583165356_0
timestamp 1713338890
transform 1 0 6481 0 1 6805
box -5445 -95 5445 95
use M1_PSUB_CDNS_69033583165356  M1_PSUB_CDNS_69033583165356_1
timestamp 1713338890
transform 1 0 6481 0 1 12677
box -5445 -95 5445 95
use M1_PSUB_CDNS_69033583165356  M1_PSUB_CDNS_69033583165356_2
timestamp 1713338890
transform 1 0 6481 0 1 18549
box -5445 -95 5445 95
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_0
timestamp 1713338890
transform 1 0 6481 0 1 227
box -254 -146 254 146
use M2_M1_CDNS_6903358316535  M2_M1_CDNS_6903358316535_1
timestamp 1713338890
transform 1 0 6481 0 1 25127
box -254 -146 254 146
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_0
timestamp 1713338890
transform 1 0 1313 0 1 3869
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_1
timestamp 1713338890
transform 1 0 11649 0 1 3869
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_2
timestamp 1713338890
transform 1 0 1313 0 1 9741
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_3
timestamp 1713338890
transform 1 0 11649 0 1 9741
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_4
timestamp 1713338890
transform 1 0 1313 0 1 15613
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_5
timestamp 1713338890
transform 1 0 11649 0 1 15613
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_6
timestamp 1713338890
transform 1 0 1313 0 1 21485
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165362  M2_M1_CDNS_69033583165362_7
timestamp 1713338890
transform 1 0 11649 0 1 21485
box -92 -2414 92 2414
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_0
timestamp 1713338890
transform 1 0 2758 0 1 6805
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_1
timestamp 1713338890
transform 1 0 5128 0 1 6805
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_2
timestamp 1713338890
transform -1 0 7834 0 1 6805
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_3
timestamp 1713338890
transform -1 0 10204 0 1 6805
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_4
timestamp 1713338890
transform 1 0 2758 0 1 12677
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_5
timestamp 1713338890
transform 1 0 5128 0 1 12677
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_6
timestamp 1713338890
transform -1 0 10204 0 1 12677
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_7
timestamp 1713338890
transform -1 0 7834 0 1 12677
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_8
timestamp 1713338890
transform 1 0 2758 0 1 18549
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_9
timestamp 1713338890
transform 1 0 5128 0 1 18549
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_10
timestamp 1713338890
transform -1 0 7834 0 1 18549
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165506  M2_M1_CDNS_69033583165506_11
timestamp 1713338890
transform -1 0 10204 0 1 18549
box -1010 -92 1010 92
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_0
timestamp 1713338890
transform 1 0 1573 0 1 227
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_1
timestamp 1713338890
transform -1 0 3943 0 1 227
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_2
timestamp 1713338890
transform -1 0 9019 0 1 227
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_3
timestamp 1713338890
transform -1 0 11389 0 1 227
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_4
timestamp 1713338890
transform -1 0 11389 0 1 25127
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_5
timestamp 1713338890
transform -1 0 9019 0 1 25127
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_6
timestamp 1713338890
transform 1 0 1573 0 1 25127
box -92 -146 92 146
use M2_M1_CDNS_69033583165507  M2_M1_CDNS_69033583165507_7
timestamp 1713338890
transform -1 0 3943 0 1 25127
box -92 -146 92 146
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_0
timestamp 1713338890
transform 1 0 2758 0 1 2405
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_1
timestamp 1713338890
transform 1 0 2758 0 1 1917
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_2
timestamp 1713338890
transform 1 0 2758 0 1 1429
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_3
timestamp 1713338890
transform 1 0 2758 0 1 2893
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_4
timestamp 1713338890
transform 1 0 2758 0 1 3381
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_5
timestamp 1713338890
transform 1 0 2758 0 1 3869
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_6
timestamp 1713338890
transform 1 0 2758 0 1 4357
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_7
timestamp 1713338890
transform 1 0 2758 0 1 4845
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_8
timestamp 1713338890
transform 1 0 5128 0 1 4357
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_9
timestamp 1713338890
transform 1 0 5128 0 1 3869
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_10
timestamp 1713338890
transform 1 0 5128 0 1 3381
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_11
timestamp 1713338890
transform 1 0 5128 0 1 2893
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_12
timestamp 1713338890
transform 1 0 5128 0 1 2405
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_13
timestamp 1713338890
transform 1 0 5128 0 1 1917
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_14
timestamp 1713338890
transform 1 0 5128 0 1 1429
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_15
timestamp 1713338890
transform 1 0 5128 0 1 4845
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_16
timestamp 1713338890
transform -1 0 7834 0 1 4845
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_17
timestamp 1713338890
transform -1 0 7834 0 1 4357
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_18
timestamp 1713338890
transform -1 0 7834 0 1 3869
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_19
timestamp 1713338890
transform -1 0 7834 0 1 3381
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_20
timestamp 1713338890
transform -1 0 7834 0 1 2893
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_21
timestamp 1713338890
transform -1 0 7834 0 1 2405
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_22
timestamp 1713338890
transform -1 0 7834 0 1 1429
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_23
timestamp 1713338890
transform -1 0 7834 0 1 1917
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_24
timestamp 1713338890
transform -1 0 10204 0 1 1429
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_25
timestamp 1713338890
transform -1 0 10204 0 1 1917
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_26
timestamp 1713338890
transform -1 0 10204 0 1 2405
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_27
timestamp 1713338890
transform -1 0 10204 0 1 2893
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_28
timestamp 1713338890
transform -1 0 10204 0 1 3381
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_29
timestamp 1713338890
transform -1 0 10204 0 1 3869
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_30
timestamp 1713338890
transform -1 0 10204 0 1 4357
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_31
timestamp 1713338890
transform -1 0 10204 0 1 4845
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_32
timestamp 1713338890
transform 1 0 2758 0 1 5821
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_33
timestamp 1713338890
transform 1 0 2758 0 1 5333
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_34
timestamp 1713338890
transform 1 0 2758 0 1 7301
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_35
timestamp 1713338890
transform 1 0 2758 0 1 6309
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_36
timestamp 1713338890
transform 1 0 2758 0 1 7789
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_37
timestamp 1713338890
transform 1 0 2758 0 1 8277
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_38
timestamp 1713338890
transform 1 0 2758 0 1 8765
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_39
timestamp 1713338890
transform 1 0 2758 0 1 9253
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_40
timestamp 1713338890
transform 1 0 2758 0 1 9741
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_41
timestamp 1713338890
transform 1 0 5128 0 1 5333
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_42
timestamp 1713338890
transform 1 0 5128 0 1 5821
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_43
timestamp 1713338890
transform 1 0 5128 0 1 6309
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_44
timestamp 1713338890
transform 1 0 5128 0 1 7301
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_45
timestamp 1713338890
transform 1 0 5128 0 1 7789
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_46
timestamp 1713338890
transform 1 0 5128 0 1 8277
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_47
timestamp 1713338890
transform 1 0 5128 0 1 8765
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_48
timestamp 1713338890
transform 1 0 5128 0 1 9253
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_49
timestamp 1713338890
transform 1 0 5128 0 1 9741
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_50
timestamp 1713338890
transform -1 0 7834 0 1 5333
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_51
timestamp 1713338890
transform -1 0 7834 0 1 5821
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_52
timestamp 1713338890
transform -1 0 7834 0 1 6309
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_53
timestamp 1713338890
transform -1 0 7834 0 1 7301
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_54
timestamp 1713338890
transform -1 0 7834 0 1 7789
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_55
timestamp 1713338890
transform -1 0 7834 0 1 8277
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_56
timestamp 1713338890
transform -1 0 7834 0 1 8765
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_57
timestamp 1713338890
transform -1 0 7834 0 1 9253
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_58
timestamp 1713338890
transform -1 0 7834 0 1 9741
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_59
timestamp 1713338890
transform -1 0 10204 0 1 5333
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_60
timestamp 1713338890
transform -1 0 10204 0 1 5821
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_61
timestamp 1713338890
transform -1 0 10204 0 1 6309
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_62
timestamp 1713338890
transform -1 0 10204 0 1 7301
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_63
timestamp 1713338890
transform -1 0 10204 0 1 7789
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_64
timestamp 1713338890
transform -1 0 10204 0 1 8277
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_65
timestamp 1713338890
transform -1 0 10204 0 1 8765
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_66
timestamp 1713338890
transform -1 0 10204 0 1 9253
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_67
timestamp 1713338890
transform -1 0 10204 0 1 9741
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_68
timestamp 1713338890
transform 1 0 5128 0 1 10229
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_69
timestamp 1713338890
transform 1 0 2758 0 1 10229
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_70
timestamp 1713338890
transform -1 0 7834 0 1 10229
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_71
timestamp 1713338890
transform -1 0 10204 0 1 10229
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_72
timestamp 1713338890
transform 1 0 5128 0 1 10717
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_73
timestamp 1713338890
transform 1 0 2758 0 1 10717
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_74
timestamp 1713338890
transform -1 0 7834 0 1 10717
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_75
timestamp 1713338890
transform -1 0 10204 0 1 10717
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_76
timestamp 1713338890
transform 1 0 5128 0 1 11205
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_77
timestamp 1713338890
transform 1 0 2758 0 1 11205
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_78
timestamp 1713338890
transform -1 0 7834 0 1 11205
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_79
timestamp 1713338890
transform -1 0 10204 0 1 11205
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_80
timestamp 1713338890
transform 1 0 5128 0 1 11693
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_81
timestamp 1713338890
transform 1 0 2758 0 1 11693
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_82
timestamp 1713338890
transform -1 0 7834 0 1 11693
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_83
timestamp 1713338890
transform -1 0 10204 0 1 11693
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_84
timestamp 1713338890
transform 1 0 5128 0 1 12181
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_85
timestamp 1713338890
transform 1 0 2758 0 1 12181
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_86
timestamp 1713338890
transform -1 0 7834 0 1 12181
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_87
timestamp 1713338890
transform -1 0 10204 0 1 12181
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_88
timestamp 1713338890
transform 1 0 2758 0 1 15125
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_89
timestamp 1713338890
transform 1 0 2758 0 1 14637
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_90
timestamp 1713338890
transform 1 0 2758 0 1 14149
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_91
timestamp 1713338890
transform 1 0 2758 0 1 13173
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_92
timestamp 1713338890
transform 1 0 2758 0 1 13661
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_93
timestamp 1713338890
transform 1 0 2758 0 1 15613
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_94
timestamp 1713338890
transform 1 0 2758 0 1 16101
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_95
timestamp 1713338890
transform 1 0 2758 0 1 16589
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_96
timestamp 1713338890
transform 1 0 2758 0 1 17077
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_97
timestamp 1713338890
transform 1 0 2758 0 1 17565
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_98
timestamp 1713338890
transform 1 0 5128 0 1 13173
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_99
timestamp 1713338890
transform 1 0 5128 0 1 13661
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_100
timestamp 1713338890
transform 1 0 5128 0 1 14149
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_101
timestamp 1713338890
transform 1 0 5128 0 1 14637
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_102
timestamp 1713338890
transform 1 0 5128 0 1 15125
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_103
timestamp 1713338890
transform 1 0 5128 0 1 15613
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_104
timestamp 1713338890
transform 1 0 5128 0 1 16101
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_105
timestamp 1713338890
transform 1 0 5128 0 1 16589
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_106
timestamp 1713338890
transform 1 0 5128 0 1 17077
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_107
timestamp 1713338890
transform 1 0 5128 0 1 17565
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_108
timestamp 1713338890
transform -1 0 7834 0 1 13173
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_109
timestamp 1713338890
transform -1 0 7834 0 1 13661
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_110
timestamp 1713338890
transform -1 0 7834 0 1 14149
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_111
timestamp 1713338890
transform -1 0 7834 0 1 14637
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_112
timestamp 1713338890
transform -1 0 7834 0 1 15125
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_113
timestamp 1713338890
transform -1 0 7834 0 1 15613
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_114
timestamp 1713338890
transform -1 0 7834 0 1 16101
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_115
timestamp 1713338890
transform -1 0 7834 0 1 16589
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_116
timestamp 1713338890
transform -1 0 7834 0 1 17077
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_117
timestamp 1713338890
transform -1 0 7834 0 1 17565
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_118
timestamp 1713338890
transform -1 0 10204 0 1 13173
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_119
timestamp 1713338890
transform -1 0 10204 0 1 13661
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_120
timestamp 1713338890
transform -1 0 10204 0 1 14149
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_121
timestamp 1713338890
transform -1 0 10204 0 1 14637
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_122
timestamp 1713338890
transform -1 0 10204 0 1 15125
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_123
timestamp 1713338890
transform -1 0 10204 0 1 15613
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_124
timestamp 1713338890
transform -1 0 10204 0 1 16101
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_125
timestamp 1713338890
transform -1 0 10204 0 1 16589
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_126
timestamp 1713338890
transform -1 0 10204 0 1 17077
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_127
timestamp 1713338890
transform -1 0 10204 0 1 17565
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_128
timestamp 1713338890
transform 1 0 2758 0 1 19533
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_129
timestamp 1713338890
transform 1 0 2758 0 1 18053
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_130
timestamp 1713338890
transform 1 0 2758 0 1 20021
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_131
timestamp 1713338890
transform 1 0 2758 0 1 19045
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_132
timestamp 1713338890
transform 1 0 2758 0 1 20509
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_133
timestamp 1713338890
transform 1 0 2758 0 1 20997
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_134
timestamp 1713338890
transform 1 0 2758 0 1 21485
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_135
timestamp 1713338890
transform 1 0 2758 0 1 21973
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_136
timestamp 1713338890
transform 1 0 2758 0 1 22461
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_137
timestamp 1713338890
transform 1 0 5128 0 1 18053
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_138
timestamp 1713338890
transform 1 0 5128 0 1 19045
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_139
timestamp 1713338890
transform 1 0 5128 0 1 19533
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_140
timestamp 1713338890
transform 1 0 5128 0 1 20021
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_141
timestamp 1713338890
transform 1 0 5128 0 1 20509
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_142
timestamp 1713338890
transform 1 0 5128 0 1 20997
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_143
timestamp 1713338890
transform 1 0 5128 0 1 21485
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_144
timestamp 1713338890
transform 1 0 5128 0 1 21973
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_145
timestamp 1713338890
transform 1 0 5128 0 1 22461
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_146
timestamp 1713338890
transform -1 0 7834 0 1 18053
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_147
timestamp 1713338890
transform -1 0 7834 0 1 19045
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_148
timestamp 1713338890
transform -1 0 7834 0 1 19533
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_149
timestamp 1713338890
transform -1 0 7834 0 1 20021
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_150
timestamp 1713338890
transform -1 0 7834 0 1 20509
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_151
timestamp 1713338890
transform -1 0 7834 0 1 20997
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_152
timestamp 1713338890
transform -1 0 7834 0 1 21485
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_153
timestamp 1713338890
transform -1 0 7834 0 1 21973
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_154
timestamp 1713338890
transform -1 0 7834 0 1 22461
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_155
timestamp 1713338890
transform -1 0 10204 0 1 18053
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_156
timestamp 1713338890
transform -1 0 10204 0 1 19045
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_157
timestamp 1713338890
transform -1 0 10204 0 1 19533
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_158
timestamp 1713338890
transform -1 0 10204 0 1 20021
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_159
timestamp 1713338890
transform -1 0 10204 0 1 20509
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_160
timestamp 1713338890
transform -1 0 10204 0 1 20997
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_161
timestamp 1713338890
transform -1 0 10204 0 1 21485
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_162
timestamp 1713338890
transform -1 0 10204 0 1 21973
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_163
timestamp 1713338890
transform -1 0 10204 0 1 22461
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_164
timestamp 1713338890
transform -1 0 7834 0 1 22949
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_165
timestamp 1713338890
transform -1 0 10204 0 1 22949
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_166
timestamp 1713338890
transform 1 0 2758 0 1 22949
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_167
timestamp 1713338890
transform 1 0 5128 0 1 22949
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_168
timestamp 1713338890
transform 1 0 2758 0 1 23437
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_169
timestamp 1713338890
transform 1 0 5128 0 1 23437
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_170
timestamp 1713338890
transform -1 0 7834 0 1 23437
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_171
timestamp 1713338890
transform -1 0 10204 0 1 23437
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_172
timestamp 1713338890
transform -1 0 7834 0 1 23925
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_173
timestamp 1713338890
transform -1 0 10204 0 1 23925
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_174
timestamp 1713338890
transform 1 0 5128 0 1 23925
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165509  M2_M1_CDNS_69033583165509_175
timestamp 1713338890
transform 1 0 2758 0 1 23925
box -1010 -38 1010 38
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_0
timestamp 1713338890
transform 1 0 2758 0 1 827
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_1
timestamp 1713338890
transform 1 0 5128 0 1 827
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_2
timestamp 1713338890
transform -1 0 7834 0 1 827
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_3
timestamp 1713338890
transform -1 0 10204 0 1 827
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_4
timestamp 1713338890
transform -1 0 10204 0 1 24527
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_5
timestamp 1713338890
transform -1 0 7834 0 1 24527
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_6
timestamp 1713338890
transform 1 0 2758 0 1 24527
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165510  M2_M1_CDNS_69033583165510_7
timestamp 1713338890
transform 1 0 5128 0 1 24527
box -1010 -146 1010 146
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_0
timestamp 1713338890
transform 1 0 1573 0 1 1673
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_1
timestamp 1713338890
transform 1 0 1573 0 1 2161
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_2
timestamp 1713338890
transform 1 0 1573 0 1 2649
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_3
timestamp 1713338890
transform 1 0 1573 0 1 3137
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_4
timestamp 1713338890
transform 1 0 1573 0 1 3625
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_5
timestamp 1713338890
transform 1 0 1573 0 1 4113
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_6
timestamp 1713338890
transform 1 0 1573 0 1 4601
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_7
timestamp 1713338890
transform -1 0 3943 0 1 4601
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_8
timestamp 1713338890
transform -1 0 3943 0 1 4113
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_9
timestamp 1713338890
transform -1 0 3943 0 1 3625
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_10
timestamp 1713338890
transform -1 0 3943 0 1 3137
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_11
timestamp 1713338890
transform -1 0 3943 0 1 2649
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_12
timestamp 1713338890
transform -1 0 3943 0 1 2161
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_13
timestamp 1713338890
transform -1 0 3943 0 1 1673
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_14
timestamp 1713338890
transform -1 0 9019 0 1 1673
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_15
timestamp 1713338890
transform -1 0 9019 0 1 2161
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_16
timestamp 1713338890
transform -1 0 9019 0 1 2649
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_17
timestamp 1713338890
transform -1 0 9019 0 1 3137
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_18
timestamp 1713338890
transform -1 0 9019 0 1 3625
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_19
timestamp 1713338890
transform -1 0 9019 0 1 4113
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_20
timestamp 1713338890
transform -1 0 9019 0 1 4601
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_21
timestamp 1713338890
transform -1 0 11389 0 1 4601
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_22
timestamp 1713338890
transform -1 0 11389 0 1 4113
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_23
timestamp 1713338890
transform -1 0 11389 0 1 3625
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_24
timestamp 1713338890
transform -1 0 11389 0 1 3137
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_25
timestamp 1713338890
transform -1 0 11389 0 1 1673
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_26
timestamp 1713338890
transform -1 0 11389 0 1 2161
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_27
timestamp 1713338890
transform -1 0 11389 0 1 2649
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_28
timestamp 1713338890
transform 1 0 1573 0 1 5089
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_29
timestamp 1713338890
transform 1 0 1573 0 1 5577
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_30
timestamp 1713338890
transform 1 0 1573 0 1 6065
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_31
timestamp 1713338890
transform 1 0 1573 0 1 7545
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_32
timestamp 1713338890
transform 1 0 1573 0 1 8033
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_33
timestamp 1713338890
transform 1 0 1573 0 1 8521
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_34
timestamp 1713338890
transform 1 0 1573 0 1 9009
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_35
timestamp 1713338890
transform 1 0 1573 0 1 9497
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_36
timestamp 1713338890
transform -1 0 3943 0 1 9497
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_37
timestamp 1713338890
transform -1 0 3943 0 1 9009
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_38
timestamp 1713338890
transform -1 0 3943 0 1 8521
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_39
timestamp 1713338890
transform -1 0 3943 0 1 8033
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_40
timestamp 1713338890
transform -1 0 3943 0 1 7545
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_41
timestamp 1713338890
transform -1 0 3943 0 1 6065
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_42
timestamp 1713338890
transform -1 0 3943 0 1 5577
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_43
timestamp 1713338890
transform -1 0 3943 0 1 5089
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_44
timestamp 1713338890
transform -1 0 9019 0 1 5089
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_45
timestamp 1713338890
transform -1 0 9019 0 1 5577
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_46
timestamp 1713338890
transform -1 0 9019 0 1 6065
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_47
timestamp 1713338890
transform -1 0 9019 0 1 7545
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_48
timestamp 1713338890
transform -1 0 9019 0 1 8033
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_49
timestamp 1713338890
transform -1 0 9019 0 1 8521
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_50
timestamp 1713338890
transform -1 0 9019 0 1 9009
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_51
timestamp 1713338890
transform -1 0 9019 0 1 9497
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_52
timestamp 1713338890
transform -1 0 11389 0 1 5089
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_53
timestamp 1713338890
transform -1 0 11389 0 1 9497
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_54
timestamp 1713338890
transform -1 0 11389 0 1 9009
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_55
timestamp 1713338890
transform -1 0 11389 0 1 8521
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_56
timestamp 1713338890
transform -1 0 11389 0 1 8033
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_57
timestamp 1713338890
transform -1 0 11389 0 1 7545
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_58
timestamp 1713338890
transform -1 0 11389 0 1 6065
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_59
timestamp 1713338890
transform -1 0 11389 0 1 5577
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_60
timestamp 1713338890
transform 1 0 1573 0 1 9985
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_61
timestamp 1713338890
transform -1 0 3943 0 1 9985
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_62
timestamp 1713338890
transform -1 0 9019 0 1 9985
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_63
timestamp 1713338890
transform -1 0 11389 0 1 9985
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_64
timestamp 1713338890
transform 1 0 1573 0 1 10473
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_65
timestamp 1713338890
transform -1 0 3943 0 1 10473
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_66
timestamp 1713338890
transform -1 0 9019 0 1 10473
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_67
timestamp 1713338890
transform -1 0 11389 0 1 10473
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_68
timestamp 1713338890
transform 1 0 1573 0 1 10961
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_69
timestamp 1713338890
transform -1 0 3943 0 1 10961
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_70
timestamp 1713338890
transform -1 0 9019 0 1 10961
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_71
timestamp 1713338890
transform -1 0 11389 0 1 10961
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_72
timestamp 1713338890
transform 1 0 1573 0 1 11449
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_73
timestamp 1713338890
transform -1 0 3943 0 1 11449
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_74
timestamp 1713338890
transform -1 0 9019 0 1 11449
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_75
timestamp 1713338890
transform -1 0 11389 0 1 11449
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_76
timestamp 1713338890
transform 1 0 1573 0 1 11937
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_77
timestamp 1713338890
transform -1 0 3943 0 1 11937
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_78
timestamp 1713338890
transform -1 0 9019 0 1 11937
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_79
timestamp 1713338890
transform -1 0 11389 0 1 11937
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_80
timestamp 1713338890
transform 1 0 1573 0 1 13905
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_81
timestamp 1713338890
transform 1 0 1573 0 1 14393
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_82
timestamp 1713338890
transform 1 0 1573 0 1 14881
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_83
timestamp 1713338890
transform 1 0 1573 0 1 13417
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_84
timestamp 1713338890
transform 1 0 1573 0 1 15369
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_85
timestamp 1713338890
transform 1 0 1573 0 1 15857
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_86
timestamp 1713338890
transform 1 0 1573 0 1 16345
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_87
timestamp 1713338890
transform 1 0 1573 0 1 16833
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_88
timestamp 1713338890
transform 1 0 1573 0 1 17321
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_89
timestamp 1713338890
transform -1 0 3943 0 1 17321
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_90
timestamp 1713338890
transform -1 0 3943 0 1 16833
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_91
timestamp 1713338890
transform -1 0 3943 0 1 16345
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_92
timestamp 1713338890
transform -1 0 3943 0 1 15857
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_93
timestamp 1713338890
transform -1 0 3943 0 1 15369
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_94
timestamp 1713338890
transform -1 0 3943 0 1 14881
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_95
timestamp 1713338890
transform -1 0 3943 0 1 14393
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_96
timestamp 1713338890
transform -1 0 3943 0 1 13905
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_97
timestamp 1713338890
transform -1 0 3943 0 1 13417
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_98
timestamp 1713338890
transform -1 0 9019 0 1 13417
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_99
timestamp 1713338890
transform -1 0 9019 0 1 13905
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_100
timestamp 1713338890
transform -1 0 9019 0 1 14393
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_101
timestamp 1713338890
transform -1 0 9019 0 1 14881
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_102
timestamp 1713338890
transform -1 0 9019 0 1 15369
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_103
timestamp 1713338890
transform -1 0 9019 0 1 15857
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_104
timestamp 1713338890
transform -1 0 9019 0 1 16345
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_105
timestamp 1713338890
transform -1 0 9019 0 1 16833
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_106
timestamp 1713338890
transform -1 0 9019 0 1 17321
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_107
timestamp 1713338890
transform -1 0 11389 0 1 14881
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_108
timestamp 1713338890
transform -1 0 11389 0 1 14393
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_109
timestamp 1713338890
transform -1 0 11389 0 1 13905
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_110
timestamp 1713338890
transform -1 0 11389 0 1 13417
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_111
timestamp 1713338890
transform -1 0 11389 0 1 17321
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_112
timestamp 1713338890
transform -1 0 11389 0 1 16833
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_113
timestamp 1713338890
transform -1 0 11389 0 1 16345
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_114
timestamp 1713338890
transform -1 0 11389 0 1 15857
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_115
timestamp 1713338890
transform -1 0 11389 0 1 15369
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_116
timestamp 1713338890
transform 1 0 1573 0 1 17809
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_117
timestamp 1713338890
transform 1 0 1573 0 1 19289
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_118
timestamp 1713338890
transform 1 0 1573 0 1 19777
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_119
timestamp 1713338890
transform 1 0 1573 0 1 20265
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_120
timestamp 1713338890
transform 1 0 1573 0 1 20753
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_121
timestamp 1713338890
transform 1 0 1573 0 1 21241
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_122
timestamp 1713338890
transform 1 0 1573 0 1 21729
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_123
timestamp 1713338890
transform 1 0 1573 0 1 22217
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_124
timestamp 1713338890
transform -1 0 3943 0 1 17809
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_125
timestamp 1713338890
transform -1 0 3943 0 1 19777
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_126
timestamp 1713338890
transform -1 0 3943 0 1 19289
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_127
timestamp 1713338890
transform -1 0 3943 0 1 20265
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_128
timestamp 1713338890
transform -1 0 3943 0 1 20753
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_129
timestamp 1713338890
transform -1 0 3943 0 1 21241
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_130
timestamp 1713338890
transform -1 0 3943 0 1 21729
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_131
timestamp 1713338890
transform -1 0 3943 0 1 22217
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_132
timestamp 1713338890
transform -1 0 9019 0 1 17809
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_133
timestamp 1713338890
transform -1 0 9019 0 1 19289
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_134
timestamp 1713338890
transform -1 0 9019 0 1 19777
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_135
timestamp 1713338890
transform -1 0 9019 0 1 20265
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_136
timestamp 1713338890
transform -1 0 9019 0 1 20753
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_137
timestamp 1713338890
transform -1 0 9019 0 1 21241
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_138
timestamp 1713338890
transform -1 0 9019 0 1 21729
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_139
timestamp 1713338890
transform -1 0 9019 0 1 22217
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_140
timestamp 1713338890
transform -1 0 11389 0 1 22217
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_141
timestamp 1713338890
transform -1 0 11389 0 1 21241
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_142
timestamp 1713338890
transform -1 0 11389 0 1 21729
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_143
timestamp 1713338890
transform -1 0 11389 0 1 20753
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_144
timestamp 1713338890
transform -1 0 11389 0 1 20265
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_145
timestamp 1713338890
transform -1 0 11389 0 1 19777
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_146
timestamp 1713338890
transform -1 0 11389 0 1 19289
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_147
timestamp 1713338890
transform -1 0 11389 0 1 17809
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_148
timestamp 1713338890
transform -1 0 9019 0 1 22705
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_149
timestamp 1713338890
transform -1 0 11389 0 1 22705
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_150
timestamp 1713338890
transform 1 0 1573 0 1 22705
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_151
timestamp 1713338890
transform -1 0 3943 0 1 22705
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_152
timestamp 1713338890
transform 1 0 1573 0 1 23193
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_153
timestamp 1713338890
transform -1 0 3943 0 1 23193
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_154
timestamp 1713338890
transform -1 0 9019 0 1 23193
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_155
timestamp 1713338890
transform -1 0 11389 0 1 23193
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_156
timestamp 1713338890
transform 1 0 1573 0 1 23681
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_157
timestamp 1713338890
transform -1 0 3943 0 1 23681
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_158
timestamp 1713338890
transform -1 0 9019 0 1 23681
box -92 -38 92 38
use M2_M1_CDNS_69033583165511  M2_M1_CDNS_69033583165511_159
timestamp 1713338890
transform -1 0 11389 0 1 23681
box -92 -38 92 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_0
timestamp 1713338890
transform 1 0 6481 0 1 1673
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_1
timestamp 1713338890
transform 1 0 6481 0 1 2161
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_2
timestamp 1713338890
transform 1 0 6481 0 1 2649
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_3
timestamp 1713338890
transform 1 0 6481 0 1 3137
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_4
timestamp 1713338890
transform 1 0 6481 0 1 3625
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_5
timestamp 1713338890
transform 1 0 6481 0 1 4113
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_6
timestamp 1713338890
transform 1 0 6481 0 1 4601
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_7
timestamp 1713338890
transform 1 0 6481 0 1 8521
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_8
timestamp 1713338890
transform 1 0 6481 0 1 5089
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_9
timestamp 1713338890
transform 1 0 6481 0 1 5577
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_10
timestamp 1713338890
transform 1 0 6481 0 1 7545
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_11
timestamp 1713338890
transform 1 0 6481 0 1 8033
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_12
timestamp 1713338890
transform 1 0 6481 0 1 9009
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_13
timestamp 1713338890
transform 1 0 6481 0 1 9497
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_14
timestamp 1713338890
transform 1 0 6481 0 1 6065
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_15
timestamp 1713338890
transform 1 0 6481 0 1 9985
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_16
timestamp 1713338890
transform 1 0 6481 0 1 10473
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_17
timestamp 1713338890
transform 1 0 6481 0 1 10961
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_18
timestamp 1713338890
transform 1 0 6481 0 1 11449
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_19
timestamp 1713338890
transform 1 0 6481 0 1 11937
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_20
timestamp 1713338890
transform 1 0 6481 0 1 13905
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_21
timestamp 1713338890
transform 1 0 6481 0 1 14393
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_22
timestamp 1713338890
transform 1 0 6481 0 1 14881
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_23
timestamp 1713338890
transform 1 0 6481 0 1 15369
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_24
timestamp 1713338890
transform 1 0 6481 0 1 15857
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_25
timestamp 1713338890
transform 1 0 6481 0 1 16345
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_26
timestamp 1713338890
transform 1 0 6481 0 1 16833
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_27
timestamp 1713338890
transform 1 0 6481 0 1 17321
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_28
timestamp 1713338890
transform 1 0 6481 0 1 13417
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_29
timestamp 1713338890
transform 1 0 6481 0 1 17809
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_30
timestamp 1713338890
transform 1 0 6481 0 1 19289
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_31
timestamp 1713338890
transform 1 0 6481 0 1 19777
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_32
timestamp 1713338890
transform 1 0 6481 0 1 20265
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_33
timestamp 1713338890
transform 1 0 6481 0 1 20753
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_34
timestamp 1713338890
transform 1 0 6481 0 1 21241
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_35
timestamp 1713338890
transform 1 0 6481 0 1 21729
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_36
timestamp 1713338890
transform 1 0 6481 0 1 22217
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_37
timestamp 1713338890
transform 1 0 6481 0 1 22705
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_38
timestamp 1713338890
transform 1 0 6481 0 1 23193
box -254 -38 254 38
use M2_M1_CDNS_69033583165526  M2_M1_CDNS_69033583165526_39
timestamp 1713338890
transform 1 0 6481 0 1 23681
box -254 -38 254 38
use M2_M1_CDNS_69033583165527  M2_M1_CDNS_69033583165527_0
timestamp 1713338890
transform 1 0 777 0 1 12677
box -146 -12026 146 12026
use M2_M1_CDNS_69033583165527  M2_M1_CDNS_69033583165527_1
timestamp 1713338890
transform 1 0 12185 0 1 12677
box -146 -12026 146 12026
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_0
timestamp 1713338890
transform 0 -1 11481 1 0 1481
box -88 -44 4864 10044
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_1
timestamp 1713338890
transform 0 -1 11481 1 0 7353
box -88 -44 4864 10044
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_2
timestamp 1713338890
transform 0 -1 11481 1 0 13225
box -88 -44 4864 10044
use nmos_6p0_CDNS_406619531457  nmos_6p0_CDNS_406619531457_3
timestamp 1713338890
transform 0 -1 11481 1 0 19097
box -88 -44 4864 10044
<< end >>
