magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1247 -1589 1247 1589
<< metal1 >>
rect -247 583 247 589
rect -247 557 -241 583
rect -215 557 -165 583
rect -139 557 -89 583
rect -63 557 -13 583
rect 13 557 63 583
rect 89 557 139 583
rect 165 557 215 583
rect 241 557 247 583
rect -247 507 247 557
rect -247 481 -241 507
rect -215 481 -165 507
rect -139 481 -89 507
rect -63 481 -13 507
rect 13 481 63 507
rect 89 481 139 507
rect 165 481 215 507
rect 241 481 247 507
rect -247 431 247 481
rect -247 405 -241 431
rect -215 405 -165 431
rect -139 405 -89 431
rect -63 405 -13 431
rect 13 405 63 431
rect 89 405 139 431
rect 165 405 215 431
rect 241 405 247 431
rect -247 355 247 405
rect -247 329 -241 355
rect -215 329 -165 355
rect -139 329 -89 355
rect -63 329 -13 355
rect 13 329 63 355
rect 89 329 139 355
rect 165 329 215 355
rect 241 329 247 355
rect -247 279 247 329
rect -247 253 -241 279
rect -215 253 -165 279
rect -139 253 -89 279
rect -63 253 -13 279
rect 13 253 63 279
rect 89 253 139 279
rect 165 253 215 279
rect 241 253 247 279
rect -247 203 247 253
rect -247 177 -241 203
rect -215 177 -165 203
rect -139 177 -89 203
rect -63 177 -13 203
rect 13 177 63 203
rect 89 177 139 203
rect 165 177 215 203
rect 241 177 247 203
rect -247 127 247 177
rect -247 101 -241 127
rect -215 101 -165 127
rect -139 101 -89 127
rect -63 101 -13 127
rect 13 101 63 127
rect 89 101 139 127
rect 165 101 215 127
rect 241 101 247 127
rect -247 51 247 101
rect -247 25 -241 51
rect -215 25 -165 51
rect -139 25 -89 51
rect -63 25 -13 51
rect 13 25 63 51
rect 89 25 139 51
rect 165 25 215 51
rect 241 25 247 51
rect -247 -25 247 25
rect -247 -51 -241 -25
rect -215 -51 -165 -25
rect -139 -51 -89 -25
rect -63 -51 -13 -25
rect 13 -51 63 -25
rect 89 -51 139 -25
rect 165 -51 215 -25
rect 241 -51 247 -25
rect -247 -101 247 -51
rect -247 -127 -241 -101
rect -215 -127 -165 -101
rect -139 -127 -89 -101
rect -63 -127 -13 -101
rect 13 -127 63 -101
rect 89 -127 139 -101
rect 165 -127 215 -101
rect 241 -127 247 -101
rect -247 -177 247 -127
rect -247 -203 -241 -177
rect -215 -203 -165 -177
rect -139 -203 -89 -177
rect -63 -203 -13 -177
rect 13 -203 63 -177
rect 89 -203 139 -177
rect 165 -203 215 -177
rect 241 -203 247 -177
rect -247 -253 247 -203
rect -247 -279 -241 -253
rect -215 -279 -165 -253
rect -139 -279 -89 -253
rect -63 -279 -13 -253
rect 13 -279 63 -253
rect 89 -279 139 -253
rect 165 -279 215 -253
rect 241 -279 247 -253
rect -247 -329 247 -279
rect -247 -355 -241 -329
rect -215 -355 -165 -329
rect -139 -355 -89 -329
rect -63 -355 -13 -329
rect 13 -355 63 -329
rect 89 -355 139 -329
rect 165 -355 215 -329
rect 241 -355 247 -329
rect -247 -405 247 -355
rect -247 -431 -241 -405
rect -215 -431 -165 -405
rect -139 -431 -89 -405
rect -63 -431 -13 -405
rect 13 -431 63 -405
rect 89 -431 139 -405
rect 165 -431 215 -405
rect 241 -431 247 -405
rect -247 -481 247 -431
rect -247 -507 -241 -481
rect -215 -507 -165 -481
rect -139 -507 -89 -481
rect -63 -507 -13 -481
rect 13 -507 63 -481
rect 89 -507 139 -481
rect 165 -507 215 -481
rect 241 -507 247 -481
rect -247 -557 247 -507
rect -247 -583 -241 -557
rect -215 -583 -165 -557
rect -139 -583 -89 -557
rect -63 -583 -13 -557
rect 13 -583 63 -557
rect 89 -583 139 -557
rect 165 -583 215 -557
rect 241 -583 247 -557
rect -247 -589 247 -583
<< via1 >>
rect -241 557 -215 583
rect -165 557 -139 583
rect -89 557 -63 583
rect -13 557 13 583
rect 63 557 89 583
rect 139 557 165 583
rect 215 557 241 583
rect -241 481 -215 507
rect -165 481 -139 507
rect -89 481 -63 507
rect -13 481 13 507
rect 63 481 89 507
rect 139 481 165 507
rect 215 481 241 507
rect -241 405 -215 431
rect -165 405 -139 431
rect -89 405 -63 431
rect -13 405 13 431
rect 63 405 89 431
rect 139 405 165 431
rect 215 405 241 431
rect -241 329 -215 355
rect -165 329 -139 355
rect -89 329 -63 355
rect -13 329 13 355
rect 63 329 89 355
rect 139 329 165 355
rect 215 329 241 355
rect -241 253 -215 279
rect -165 253 -139 279
rect -89 253 -63 279
rect -13 253 13 279
rect 63 253 89 279
rect 139 253 165 279
rect 215 253 241 279
rect -241 177 -215 203
rect -165 177 -139 203
rect -89 177 -63 203
rect -13 177 13 203
rect 63 177 89 203
rect 139 177 165 203
rect 215 177 241 203
rect -241 101 -215 127
rect -165 101 -139 127
rect -89 101 -63 127
rect -13 101 13 127
rect 63 101 89 127
rect 139 101 165 127
rect 215 101 241 127
rect -241 25 -215 51
rect -165 25 -139 51
rect -89 25 -63 51
rect -13 25 13 51
rect 63 25 89 51
rect 139 25 165 51
rect 215 25 241 51
rect -241 -51 -215 -25
rect -165 -51 -139 -25
rect -89 -51 -63 -25
rect -13 -51 13 -25
rect 63 -51 89 -25
rect 139 -51 165 -25
rect 215 -51 241 -25
rect -241 -127 -215 -101
rect -165 -127 -139 -101
rect -89 -127 -63 -101
rect -13 -127 13 -101
rect 63 -127 89 -101
rect 139 -127 165 -101
rect 215 -127 241 -101
rect -241 -203 -215 -177
rect -165 -203 -139 -177
rect -89 -203 -63 -177
rect -13 -203 13 -177
rect 63 -203 89 -177
rect 139 -203 165 -177
rect 215 -203 241 -177
rect -241 -279 -215 -253
rect -165 -279 -139 -253
rect -89 -279 -63 -253
rect -13 -279 13 -253
rect 63 -279 89 -253
rect 139 -279 165 -253
rect 215 -279 241 -253
rect -241 -355 -215 -329
rect -165 -355 -139 -329
rect -89 -355 -63 -329
rect -13 -355 13 -329
rect 63 -355 89 -329
rect 139 -355 165 -329
rect 215 -355 241 -329
rect -241 -431 -215 -405
rect -165 -431 -139 -405
rect -89 -431 -63 -405
rect -13 -431 13 -405
rect 63 -431 89 -405
rect 139 -431 165 -405
rect 215 -431 241 -405
rect -241 -507 -215 -481
rect -165 -507 -139 -481
rect -89 -507 -63 -481
rect -13 -507 13 -481
rect 63 -507 89 -481
rect 139 -507 165 -481
rect 215 -507 241 -481
rect -241 -583 -215 -557
rect -165 -583 -139 -557
rect -89 -583 -63 -557
rect -13 -583 13 -557
rect 63 -583 89 -557
rect 139 -583 165 -557
rect 215 -583 241 -557
<< metal2 >>
rect -247 583 247 589
rect -247 557 -241 583
rect -215 557 -165 583
rect -139 557 -89 583
rect -63 557 -13 583
rect 13 557 63 583
rect 89 557 139 583
rect 165 557 215 583
rect 241 557 247 583
rect -247 507 247 557
rect -247 481 -241 507
rect -215 481 -165 507
rect -139 481 -89 507
rect -63 481 -13 507
rect 13 481 63 507
rect 89 481 139 507
rect 165 481 215 507
rect 241 481 247 507
rect -247 431 247 481
rect -247 405 -241 431
rect -215 405 -165 431
rect -139 405 -89 431
rect -63 405 -13 431
rect 13 405 63 431
rect 89 405 139 431
rect 165 405 215 431
rect 241 405 247 431
rect -247 355 247 405
rect -247 329 -241 355
rect -215 329 -165 355
rect -139 329 -89 355
rect -63 329 -13 355
rect 13 329 63 355
rect 89 329 139 355
rect 165 329 215 355
rect 241 329 247 355
rect -247 279 247 329
rect -247 253 -241 279
rect -215 253 -165 279
rect -139 253 -89 279
rect -63 253 -13 279
rect 13 253 63 279
rect 89 253 139 279
rect 165 253 215 279
rect 241 253 247 279
rect -247 203 247 253
rect -247 177 -241 203
rect -215 177 -165 203
rect -139 177 -89 203
rect -63 177 -13 203
rect 13 177 63 203
rect 89 177 139 203
rect 165 177 215 203
rect 241 177 247 203
rect -247 127 247 177
rect -247 101 -241 127
rect -215 101 -165 127
rect -139 101 -89 127
rect -63 101 -13 127
rect 13 101 63 127
rect 89 101 139 127
rect 165 101 215 127
rect 241 101 247 127
rect -247 51 247 101
rect -247 25 -241 51
rect -215 25 -165 51
rect -139 25 -89 51
rect -63 25 -13 51
rect 13 25 63 51
rect 89 25 139 51
rect 165 25 215 51
rect 241 25 247 51
rect -247 -25 247 25
rect -247 -51 -241 -25
rect -215 -51 -165 -25
rect -139 -51 -89 -25
rect -63 -51 -13 -25
rect 13 -51 63 -25
rect 89 -51 139 -25
rect 165 -51 215 -25
rect 241 -51 247 -25
rect -247 -101 247 -51
rect -247 -127 -241 -101
rect -215 -127 -165 -101
rect -139 -127 -89 -101
rect -63 -127 -13 -101
rect 13 -127 63 -101
rect 89 -127 139 -101
rect 165 -127 215 -101
rect 241 -127 247 -101
rect -247 -177 247 -127
rect -247 -203 -241 -177
rect -215 -203 -165 -177
rect -139 -203 -89 -177
rect -63 -203 -13 -177
rect 13 -203 63 -177
rect 89 -203 139 -177
rect 165 -203 215 -177
rect 241 -203 247 -177
rect -247 -253 247 -203
rect -247 -279 -241 -253
rect -215 -279 -165 -253
rect -139 -279 -89 -253
rect -63 -279 -13 -253
rect 13 -279 63 -253
rect 89 -279 139 -253
rect 165 -279 215 -253
rect 241 -279 247 -253
rect -247 -329 247 -279
rect -247 -355 -241 -329
rect -215 -355 -165 -329
rect -139 -355 -89 -329
rect -63 -355 -13 -329
rect 13 -355 63 -329
rect 89 -355 139 -329
rect 165 -355 215 -329
rect 241 -355 247 -329
rect -247 -405 247 -355
rect -247 -431 -241 -405
rect -215 -431 -165 -405
rect -139 -431 -89 -405
rect -63 -431 -13 -405
rect 13 -431 63 -405
rect 89 -431 139 -405
rect 165 -431 215 -405
rect 241 -431 247 -405
rect -247 -481 247 -431
rect -247 -507 -241 -481
rect -215 -507 -165 -481
rect -139 -507 -89 -481
rect -63 -507 -13 -481
rect 13 -507 63 -481
rect 89 -507 139 -481
rect 165 -507 215 -481
rect 241 -507 247 -481
rect -247 -557 247 -507
rect -247 -583 -241 -557
rect -215 -583 -165 -557
rect -139 -583 -89 -557
rect -63 -583 -13 -557
rect 13 -583 63 -557
rect 89 -583 139 -557
rect 165 -583 215 -557
rect 241 -583 247 -557
rect -247 -589 247 -583
<< end >>
