magic
tech gf180mcuC
magscale 1 10
timestamp 1691495105
<< nwell >>
rect 61 1398 2865 2680
rect 260 573 664 1398
<< pwell >>
rect 322 263 602 499
rect 763 120 2163 1278
<< nmos >>
rect 875 960 931 1210
rect 1035 960 1091 1210
rect 1195 960 1251 1210
rect 1355 960 1411 1210
rect 1515 960 1571 1210
rect 1675 960 1731 1210
rect 1835 960 1891 1210
rect 1995 960 2051 1210
rect 875 574 931 824
rect 1035 574 1091 824
rect 1195 574 1251 824
rect 1355 574 1411 824
rect 1515 574 1571 824
rect 1675 574 1731 824
rect 1835 574 1891 824
rect 1995 574 2051 824
rect 434 331 490 431
rect 875 188 931 438
rect 1035 188 1091 438
rect 1195 188 1251 438
rect 1355 188 1411 438
rect 1515 188 1571 438
rect 1675 188 1731 438
rect 1835 188 1891 438
rect 1995 188 2051 438
<< pmos >>
rect 235 2300 291 2550
rect 395 2300 451 2550
rect 555 2300 611 2550
rect 715 2300 771 2550
rect 875 2300 931 2550
rect 1035 2300 1091 2550
rect 1195 2300 1251 2550
rect 1355 2300 1411 2550
rect 1515 2300 1571 2550
rect 1675 2300 1731 2550
rect 1835 2300 1891 2550
rect 1995 2300 2051 2550
rect 2155 2300 2211 2550
rect 2315 2300 2371 2550
rect 2475 2300 2531 2550
rect 2635 2300 2691 2550
rect 235 1914 291 2164
rect 395 1914 451 2164
rect 555 1914 611 2164
rect 715 1914 771 2164
rect 875 1914 931 2164
rect 1035 1914 1091 2164
rect 1195 1914 1251 2164
rect 1355 1914 1411 2164
rect 1515 1914 1571 2164
rect 1675 1914 1731 2164
rect 1835 1914 1891 2164
rect 1995 1914 2051 2164
rect 2155 1914 2211 2164
rect 2315 1914 2371 2164
rect 2475 1914 2531 2164
rect 2635 1914 2691 2164
rect 235 1528 291 1778
rect 395 1528 451 1778
rect 555 1528 611 1778
rect 715 1528 771 1778
rect 875 1528 931 1778
rect 1035 1528 1091 1778
rect 1195 1528 1251 1778
rect 1355 1528 1411 1778
rect 1515 1528 1571 1778
rect 1675 1528 1731 1778
rect 1835 1528 1891 1778
rect 1995 1528 2051 1778
rect 2155 1528 2211 1778
rect 2315 1528 2371 1778
rect 2475 1528 2531 1778
rect 2635 1528 2691 1778
rect 434 703 490 903
<< ndiff >>
rect 787 1197 875 1210
rect 787 973 800 1197
rect 846 973 875 1197
rect 787 960 875 973
rect 931 1197 1035 1210
rect 931 973 960 1197
rect 1006 973 1035 1197
rect 931 960 1035 973
rect 1091 1197 1195 1210
rect 1091 973 1120 1197
rect 1166 973 1195 1197
rect 1091 960 1195 973
rect 1251 1197 1355 1210
rect 1251 973 1280 1197
rect 1326 973 1355 1197
rect 1251 960 1355 973
rect 1411 1197 1515 1210
rect 1411 973 1440 1197
rect 1486 973 1515 1197
rect 1411 960 1515 973
rect 1571 1197 1675 1210
rect 1571 973 1600 1197
rect 1646 973 1675 1197
rect 1571 960 1675 973
rect 1731 1197 1835 1210
rect 1731 973 1760 1197
rect 1806 973 1835 1197
rect 1731 960 1835 973
rect 1891 1197 1995 1210
rect 1891 973 1920 1197
rect 1966 973 1995 1197
rect 1891 960 1995 973
rect 2051 1197 2139 1210
rect 2051 973 2080 1197
rect 2126 973 2139 1197
rect 2051 960 2139 973
rect 787 811 875 824
rect 787 587 800 811
rect 846 587 875 811
rect 787 574 875 587
rect 931 811 1035 824
rect 931 587 960 811
rect 1006 587 1035 811
rect 931 574 1035 587
rect 1091 811 1195 824
rect 1091 587 1120 811
rect 1166 587 1195 811
rect 1091 574 1195 587
rect 1251 811 1355 824
rect 1251 587 1280 811
rect 1326 587 1355 811
rect 1251 574 1355 587
rect 1411 811 1515 824
rect 1411 587 1440 811
rect 1486 587 1515 811
rect 1411 574 1515 587
rect 1571 811 1675 824
rect 1571 587 1600 811
rect 1646 587 1675 811
rect 1571 574 1675 587
rect 1731 811 1835 824
rect 1731 587 1760 811
rect 1806 587 1835 811
rect 1731 574 1835 587
rect 1891 811 1995 824
rect 1891 587 1920 811
rect 1966 587 1995 811
rect 1891 574 1995 587
rect 2051 811 2139 824
rect 2051 587 2080 811
rect 2126 587 2139 811
rect 2051 574 2139 587
rect 346 418 434 431
rect 346 344 359 418
rect 405 344 434 418
rect 346 331 434 344
rect 490 418 578 431
rect 490 344 519 418
rect 565 344 578 418
rect 787 425 875 438
rect 490 331 578 344
rect 787 201 800 425
rect 846 201 875 425
rect 787 188 875 201
rect 931 425 1035 438
rect 931 201 960 425
rect 1006 201 1035 425
rect 931 188 1035 201
rect 1091 425 1195 438
rect 1091 201 1120 425
rect 1166 201 1195 425
rect 1091 188 1195 201
rect 1251 425 1355 438
rect 1251 201 1280 425
rect 1326 201 1355 425
rect 1251 188 1355 201
rect 1411 425 1515 438
rect 1411 201 1440 425
rect 1486 201 1515 425
rect 1411 188 1515 201
rect 1571 425 1675 438
rect 1571 201 1600 425
rect 1646 201 1675 425
rect 1571 188 1675 201
rect 1731 425 1835 438
rect 1731 201 1760 425
rect 1806 201 1835 425
rect 1731 188 1835 201
rect 1891 425 1995 438
rect 1891 201 1920 425
rect 1966 201 1995 425
rect 1891 188 1995 201
rect 2051 425 2139 438
rect 2051 201 2080 425
rect 2126 201 2139 425
rect 2051 188 2139 201
<< pdiff >>
rect 147 2537 235 2550
rect 147 2313 160 2537
rect 206 2313 235 2537
rect 147 2300 235 2313
rect 291 2537 395 2550
rect 291 2313 320 2537
rect 366 2313 395 2537
rect 291 2300 395 2313
rect 451 2537 555 2550
rect 451 2313 480 2537
rect 526 2313 555 2537
rect 451 2300 555 2313
rect 611 2537 715 2550
rect 611 2313 640 2537
rect 686 2313 715 2537
rect 611 2300 715 2313
rect 771 2537 875 2550
rect 771 2313 800 2537
rect 846 2313 875 2537
rect 771 2300 875 2313
rect 931 2537 1035 2550
rect 931 2313 960 2537
rect 1006 2313 1035 2537
rect 931 2300 1035 2313
rect 1091 2537 1195 2550
rect 1091 2313 1120 2537
rect 1166 2313 1195 2537
rect 1091 2300 1195 2313
rect 1251 2537 1355 2550
rect 1251 2313 1280 2537
rect 1326 2313 1355 2537
rect 1251 2300 1355 2313
rect 1411 2537 1515 2550
rect 1411 2313 1440 2537
rect 1486 2313 1515 2537
rect 1411 2300 1515 2313
rect 1571 2537 1675 2550
rect 1571 2313 1600 2537
rect 1646 2313 1675 2537
rect 1571 2300 1675 2313
rect 1731 2537 1835 2550
rect 1731 2313 1760 2537
rect 1806 2313 1835 2537
rect 1731 2300 1835 2313
rect 1891 2537 1995 2550
rect 1891 2313 1920 2537
rect 1966 2313 1995 2537
rect 1891 2300 1995 2313
rect 2051 2537 2155 2550
rect 2051 2313 2080 2537
rect 2126 2313 2155 2537
rect 2051 2300 2155 2313
rect 2211 2537 2315 2550
rect 2211 2313 2240 2537
rect 2286 2313 2315 2537
rect 2211 2300 2315 2313
rect 2371 2537 2475 2550
rect 2371 2313 2400 2537
rect 2446 2313 2475 2537
rect 2371 2300 2475 2313
rect 2531 2537 2635 2550
rect 2531 2313 2560 2537
rect 2606 2313 2635 2537
rect 2531 2300 2635 2313
rect 2691 2537 2779 2550
rect 2691 2313 2720 2537
rect 2766 2313 2779 2537
rect 2691 2300 2779 2313
rect 147 2151 235 2164
rect 147 1927 160 2151
rect 206 1927 235 2151
rect 147 1914 235 1927
rect 291 2151 395 2164
rect 291 1927 320 2151
rect 366 1927 395 2151
rect 291 1914 395 1927
rect 451 2151 555 2164
rect 451 1927 480 2151
rect 526 1927 555 2151
rect 451 1914 555 1927
rect 611 2151 715 2164
rect 611 1927 640 2151
rect 686 1927 715 2151
rect 611 1914 715 1927
rect 771 2151 875 2164
rect 771 1927 800 2151
rect 846 1927 875 2151
rect 771 1914 875 1927
rect 931 2151 1035 2164
rect 931 1927 960 2151
rect 1006 1927 1035 2151
rect 931 1914 1035 1927
rect 1091 2151 1195 2164
rect 1091 1927 1120 2151
rect 1166 1927 1195 2151
rect 1091 1914 1195 1927
rect 1251 2151 1355 2164
rect 1251 1927 1280 2151
rect 1326 1927 1355 2151
rect 1251 1914 1355 1927
rect 1411 2151 1515 2164
rect 1411 1927 1440 2151
rect 1486 1927 1515 2151
rect 1411 1914 1515 1927
rect 1571 2151 1675 2164
rect 1571 1927 1600 2151
rect 1646 1927 1675 2151
rect 1571 1914 1675 1927
rect 1731 2151 1835 2164
rect 1731 1927 1760 2151
rect 1806 1927 1835 2151
rect 1731 1914 1835 1927
rect 1891 2151 1995 2164
rect 1891 1927 1920 2151
rect 1966 1927 1995 2151
rect 1891 1914 1995 1927
rect 2051 2151 2155 2164
rect 2051 1927 2080 2151
rect 2126 1927 2155 2151
rect 2051 1914 2155 1927
rect 2211 2151 2315 2164
rect 2211 1927 2240 2151
rect 2286 1927 2315 2151
rect 2211 1914 2315 1927
rect 2371 2151 2475 2164
rect 2371 1927 2400 2151
rect 2446 1927 2475 2151
rect 2371 1914 2475 1927
rect 2531 2151 2635 2164
rect 2531 1927 2560 2151
rect 2606 1927 2635 2151
rect 2531 1914 2635 1927
rect 2691 2151 2779 2164
rect 2691 1927 2720 2151
rect 2766 1927 2779 2151
rect 2691 1914 2779 1927
rect 147 1765 235 1778
rect 147 1541 160 1765
rect 206 1541 235 1765
rect 147 1528 235 1541
rect 291 1765 395 1778
rect 291 1541 320 1765
rect 366 1541 395 1765
rect 291 1528 395 1541
rect 451 1765 555 1778
rect 451 1541 480 1765
rect 526 1541 555 1765
rect 451 1528 555 1541
rect 611 1765 715 1778
rect 611 1541 640 1765
rect 686 1541 715 1765
rect 611 1528 715 1541
rect 771 1765 875 1778
rect 771 1541 800 1765
rect 846 1541 875 1765
rect 771 1528 875 1541
rect 931 1765 1035 1778
rect 931 1541 960 1765
rect 1006 1541 1035 1765
rect 931 1528 1035 1541
rect 1091 1765 1195 1778
rect 1091 1541 1120 1765
rect 1166 1541 1195 1765
rect 1091 1528 1195 1541
rect 1251 1765 1355 1778
rect 1251 1541 1280 1765
rect 1326 1541 1355 1765
rect 1251 1528 1355 1541
rect 1411 1765 1515 1778
rect 1411 1541 1440 1765
rect 1486 1541 1515 1765
rect 1411 1528 1515 1541
rect 1571 1765 1675 1778
rect 1571 1541 1600 1765
rect 1646 1541 1675 1765
rect 1571 1528 1675 1541
rect 1731 1765 1835 1778
rect 1731 1541 1760 1765
rect 1806 1541 1835 1765
rect 1731 1528 1835 1541
rect 1891 1765 1995 1778
rect 1891 1541 1920 1765
rect 1966 1541 1995 1765
rect 1891 1528 1995 1541
rect 2051 1765 2155 1778
rect 2051 1541 2080 1765
rect 2126 1541 2155 1765
rect 2051 1528 2155 1541
rect 2211 1765 2315 1778
rect 2211 1541 2240 1765
rect 2286 1541 2315 1765
rect 2211 1528 2315 1541
rect 2371 1765 2475 1778
rect 2371 1541 2400 1765
rect 2446 1541 2475 1765
rect 2371 1528 2475 1541
rect 2531 1765 2635 1778
rect 2531 1541 2560 1765
rect 2606 1541 2635 1765
rect 2531 1528 2635 1541
rect 2691 1765 2779 1778
rect 2691 1541 2720 1765
rect 2766 1541 2779 1765
rect 2691 1528 2779 1541
rect 346 890 434 903
rect 346 716 359 890
rect 405 716 434 890
rect 346 703 434 716
rect 490 890 578 903
rect 490 716 519 890
rect 565 716 578 890
rect 490 703 578 716
<< ndiffc >>
rect 800 973 846 1197
rect 960 973 1006 1197
rect 1120 973 1166 1197
rect 1280 973 1326 1197
rect 1440 973 1486 1197
rect 1600 973 1646 1197
rect 1760 973 1806 1197
rect 1920 973 1966 1197
rect 2080 973 2126 1197
rect 800 587 846 811
rect 960 587 1006 811
rect 1120 587 1166 811
rect 1280 587 1326 811
rect 1440 587 1486 811
rect 1600 587 1646 811
rect 1760 587 1806 811
rect 1920 587 1966 811
rect 2080 587 2126 811
rect 359 344 405 418
rect 519 344 565 418
rect 800 201 846 425
rect 960 201 1006 425
rect 1120 201 1166 425
rect 1280 201 1326 425
rect 1440 201 1486 425
rect 1600 201 1646 425
rect 1760 201 1806 425
rect 1920 201 1966 425
rect 2080 201 2126 425
<< pdiffc >>
rect 160 2313 206 2537
rect 320 2313 366 2537
rect 480 2313 526 2537
rect 640 2313 686 2537
rect 800 2313 846 2537
rect 960 2313 1006 2537
rect 1120 2313 1166 2537
rect 1280 2313 1326 2537
rect 1440 2313 1486 2537
rect 1600 2313 1646 2537
rect 1760 2313 1806 2537
rect 1920 2313 1966 2537
rect 2080 2313 2126 2537
rect 2240 2313 2286 2537
rect 2400 2313 2446 2537
rect 2560 2313 2606 2537
rect 2720 2313 2766 2537
rect 160 1927 206 2151
rect 320 1927 366 2151
rect 480 1927 526 2151
rect 640 1927 686 2151
rect 800 1927 846 2151
rect 960 1927 1006 2151
rect 1120 1927 1166 2151
rect 1280 1927 1326 2151
rect 1440 1927 1486 2151
rect 1600 1927 1646 2151
rect 1760 1927 1806 2151
rect 1920 1927 1966 2151
rect 2080 1927 2126 2151
rect 2240 1927 2286 2151
rect 2400 1927 2446 2151
rect 2560 1927 2606 2151
rect 2720 1927 2766 2151
rect 160 1541 206 1765
rect 320 1541 366 1765
rect 480 1541 526 1765
rect 640 1541 686 1765
rect 800 1541 846 1765
rect 960 1541 1006 1765
rect 1120 1541 1166 1765
rect 1280 1541 1326 1765
rect 1440 1541 1486 1765
rect 1600 1541 1646 1765
rect 1760 1541 1806 1765
rect 1920 1541 1966 1765
rect 2080 1541 2126 1765
rect 2240 1541 2286 1765
rect 2400 1541 2446 1765
rect 2560 1541 2606 1765
rect 2720 1541 2766 1765
rect 359 716 405 890
rect 519 716 565 890
<< psubdiff >>
rect 495 236 589 263
rect 495 190 519 236
rect 565 190 589 236
rect 495 166 589 190
<< nsubdiff >>
rect 495 1039 589 1063
rect 495 993 519 1039
rect 565 993 589 1039
rect 495 969 589 993
<< psubdiffcont >>
rect 519 190 565 236
<< nsubdiffcont >>
rect 519 993 565 1039
<< polysilicon >>
rect 235 2570 2691 2626
rect 235 2550 291 2570
rect 395 2550 451 2570
rect 555 2550 611 2570
rect 715 2550 771 2570
rect 875 2550 931 2570
rect 1035 2550 1091 2570
rect 1195 2550 1251 2570
rect 1355 2550 1411 2570
rect 1515 2550 1571 2570
rect 1675 2550 1731 2570
rect 1835 2550 1891 2570
rect 1995 2550 2051 2570
rect 2155 2550 2211 2570
rect 2315 2550 2371 2570
rect 2475 2550 2531 2570
rect 2635 2550 2691 2570
rect 235 2164 291 2300
rect 395 2164 451 2300
rect 555 2164 611 2300
rect 715 2164 771 2300
rect 875 2164 931 2300
rect 1035 2164 1091 2300
rect 1195 2164 1251 2300
rect 1355 2164 1411 2300
rect 1515 2164 1571 2300
rect 1675 2164 1731 2300
rect 1835 2164 1891 2300
rect 1995 2164 2051 2300
rect 2155 2164 2211 2300
rect 2315 2164 2371 2300
rect 2475 2164 2531 2300
rect 2635 2164 2691 2300
rect 235 1778 291 1914
rect 395 1778 451 1914
rect 555 1778 611 1914
rect 715 1778 771 1914
rect 875 1778 931 1914
rect 1035 1778 1091 1914
rect 1195 1778 1251 1914
rect 1355 1778 1411 1914
rect 1515 1778 1571 1914
rect 1675 1778 1731 1914
rect 1835 1778 1891 1914
rect 1995 1778 2051 1914
rect 2155 1778 2211 1914
rect 2315 1778 2371 1914
rect 2475 1778 2531 1914
rect 2635 1778 2691 1914
rect 235 1346 291 1528
rect 395 1484 451 1528
rect 555 1484 611 1528
rect 715 1484 771 1528
rect 875 1484 931 1528
rect 1035 1484 1091 1528
rect 1195 1484 1251 1528
rect 1355 1484 1411 1528
rect 1515 1484 1571 1528
rect 1675 1484 1731 1528
rect 1835 1484 1891 1528
rect 1995 1484 2051 1528
rect 2155 1484 2211 1528
rect 2315 1484 2371 1528
rect 2475 1484 2531 1528
rect 2635 1484 2691 1528
rect 227 1333 299 1346
rect 227 1287 240 1333
rect 286 1287 299 1333
rect 227 1274 299 1287
rect 875 1210 931 1254
rect 1035 1210 1091 1254
rect 1195 1210 1251 1254
rect 1355 1210 1411 1254
rect 1515 1210 1571 1254
rect 1675 1210 1731 1254
rect 1835 1210 1891 1254
rect 1995 1210 2051 1254
rect 434 903 490 947
rect 875 824 931 960
rect 1035 824 1091 960
rect 1195 824 1251 960
rect 1355 824 1411 960
rect 1515 824 1571 960
rect 1675 824 1731 960
rect 1835 824 1891 960
rect 1995 824 2051 960
rect 434 578 490 703
rect 538 578 610 586
rect 434 573 610 578
rect 434 527 551 573
rect 597 527 610 573
rect 434 522 610 527
rect 434 431 490 522
rect 538 514 610 522
rect 875 438 931 574
rect 1035 438 1091 574
rect 1195 438 1251 574
rect 1355 438 1411 574
rect 1515 438 1571 574
rect 1675 438 1731 574
rect 1835 438 1891 574
rect 1995 438 2051 574
rect 677 344 749 357
rect 434 287 490 331
rect 677 298 690 344
rect 736 298 749 344
rect 677 285 749 298
rect 685 168 741 285
rect 875 168 931 188
rect 1035 168 1091 188
rect 1195 168 1251 188
rect 1355 168 1411 188
rect 1515 168 1571 188
rect 1675 168 1731 188
rect 1835 168 1891 188
rect 1995 168 2051 188
rect 685 112 2051 168
<< polycontact >>
rect 240 1287 286 1333
rect 551 527 597 573
rect 690 298 736 344
<< metal1 >>
rect 160 2686 1166 2732
rect 160 2537 206 2686
rect 1120 2640 1166 2686
rect 1440 2686 2446 2732
rect 1440 2640 1486 2686
rect 2400 2640 2446 2686
rect 160 2151 206 2313
rect 160 1765 206 1927
rect 160 1484 206 1541
rect 320 2594 1006 2640
rect 320 2537 366 2594
rect 320 2151 366 2313
rect 320 1765 366 1927
rect 320 1530 366 1541
rect 480 2537 526 2548
rect 480 2151 526 2313
rect 480 1765 526 1927
rect 480 1484 526 1541
rect 160 1438 526 1484
rect 229 1333 297 1344
rect 229 1287 240 1333
rect 286 1287 297 1333
rect 229 1276 297 1287
rect 480 1300 526 1438
rect 640 2537 686 2594
rect 640 2151 686 2313
rect 640 1765 686 1927
rect 640 1392 686 1541
rect 800 2537 846 2548
rect 800 2151 846 2313
rect 800 1765 846 1927
rect 800 1484 846 1541
rect 960 2537 1006 2594
rect 960 2151 1006 2313
rect 960 1765 1006 1927
rect 960 1530 1006 1541
rect 1120 2594 1486 2640
rect 1120 2537 1166 2594
rect 1120 2151 1166 2313
rect 1120 1765 1166 1927
rect 1120 1484 1166 1541
rect 800 1438 1166 1484
rect 1280 2537 1326 2548
rect 1280 2151 1326 2313
rect 1280 1765 1326 1927
rect 1280 1392 1326 1541
rect 1440 2537 1486 2594
rect 1440 2151 1486 2313
rect 1440 1765 1486 1927
rect 1440 1484 1486 1541
rect 1600 2594 2286 2640
rect 1600 2537 1646 2594
rect 1600 2151 1646 2313
rect 1600 1765 1646 1927
rect 1600 1530 1646 1541
rect 1760 2537 1806 2548
rect 1760 2151 1806 2313
rect 1760 1765 1806 1927
rect 1760 1484 1806 1541
rect 1440 1438 1806 1484
rect 1920 2537 1966 2594
rect 1920 2151 1966 2313
rect 1920 1765 1966 1927
rect 1920 1392 1966 1541
rect 2080 2537 2126 2548
rect 2080 2151 2126 2313
rect 2080 1765 2126 1927
rect 2080 1484 2126 1541
rect 2240 2537 2286 2594
rect 2240 2151 2286 2313
rect 2240 1765 2286 1927
rect 2240 1530 2286 1541
rect 2400 2594 2766 2640
rect 2400 2537 2446 2594
rect 2400 2151 2446 2313
rect 2400 1765 2446 1927
rect 2400 1484 2446 1541
rect 2560 2537 2606 2548
rect 2560 2151 2606 2313
rect 2560 1765 2606 1927
rect 2080 1438 2447 1484
rect 2560 1392 2606 1541
rect 2720 2537 2766 2594
rect 2720 2151 2766 2313
rect 2720 1765 2766 1927
rect 2720 1530 2766 1541
rect 640 1346 2717 1392
rect 240 901 286 1276
rect 480 1254 1166 1300
rect 800 1197 846 1254
rect 440 1039 644 1050
rect 440 993 519 1039
rect 565 993 644 1039
rect 440 982 644 993
rect 240 890 405 901
rect 240 855 359 890
rect 359 573 405 716
rect 519 890 565 982
rect 519 705 565 716
rect 800 811 846 973
rect 262 527 405 573
rect 359 418 405 527
rect 540 573 608 584
rect 540 527 551 573
rect 597 527 736 573
rect 540 516 608 527
rect 359 333 405 344
rect 519 418 565 429
rect 690 355 736 527
rect 800 425 846 587
rect 519 247 565 344
rect 679 344 747 355
rect 679 298 690 344
rect 736 298 747 344
rect 679 287 747 298
rect 429 236 655 247
rect 429 190 519 236
rect 565 190 655 236
rect 429 179 503 190
rect 571 179 655 190
rect 800 52 846 201
rect 960 1197 1006 1208
rect 960 811 1006 973
rect 960 425 1006 587
rect 960 144 1006 201
rect 1120 1197 1166 1254
rect 1120 811 1166 973
rect 1120 425 1166 587
rect 1120 190 1166 201
rect 1280 1197 1326 1346
rect 1280 811 1326 973
rect 1280 425 1326 587
rect 1280 144 1326 201
rect 1440 1254 1806 1300
rect 1440 1197 1486 1254
rect 1440 811 1486 973
rect 1440 425 1486 587
rect 1440 190 1486 201
rect 1600 1197 1646 1208
rect 1600 811 1646 973
rect 1600 425 1646 587
rect 1600 144 1646 201
rect 960 98 1646 144
rect 1760 1197 1806 1254
rect 1760 811 1806 973
rect 1760 425 1806 587
rect 1760 144 1806 201
rect 1920 1197 1966 1346
rect 1920 811 1966 973
rect 1920 425 1966 587
rect 1920 190 1966 201
rect 2080 1239 2305 1285
rect 2080 1197 2126 1239
rect 2080 811 2126 973
rect 2080 425 2126 587
rect 2080 144 2126 201
rect 1760 98 2126 144
rect 1760 52 1806 98
rect 800 6 1806 52
<< labels >>
flabel metal1 542 1016 542 1016 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel metal1 542 213 542 213 0 FreeSans 320 0 0 0 VSS
port 1 nsew
flabel metal1 682 550 682 550 0 FreeSans 320 0 0 0 CLK
port 2 nsew
flabel metal1 2211 1262 2211 1262 0 FreeSans 320 0 0 0 VIN
port 5 nsew
flabel metal1 2628 1369 2628 1369 0 FreeSans 320 0 0 0 VOUT
port 7 nsew
flabel psubdiffcont 542 213 542 213 0 FreeSans 320 0 0 0 Inverter_Layout_0.VSS
flabel nsubdiffcont 542 1016 542 1016 0 FreeSans 320 0 0 0 Inverter_Layout_0.VDD
flabel metal1 642 550 642 550 0 FreeSans 320 0 0 0 Inverter_Layout_0.IN
flabel metal1 323 550 323 550 0 FreeSans 320 0 0 0 Inverter_Layout_0.OUT
<< end >>
