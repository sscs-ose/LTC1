magic
tech gf180mcuD
magscale 1 10
timestamp 1713971633
<< checkpaint >>
rect -2441 -12214 42218 14749
<< nwell >>
rect 498 10526 618 10604
rect 727 10526 845 10605
rect 18601 5998 18661 6058
rect 18724 6000 18784 6060
rect 18723 5891 18783 5951
rect 12010 5650 12900 5770
rect 15503 5747 15587 5750
rect 13937 5668 14487 5747
rect 15045 5668 15595 5747
rect 15503 5664 15587 5668
rect 230 5413 6491 5646
rect 12010 5644 12930 5650
rect 16049 5644 17452 5782
rect 22892 5663 22977 5669
rect 7129 5413 22403 5644
rect 23232 5413 24815 5644
rect 26829 5413 29492 5645
rect 389 5310 939 5390
rect 762 5309 939 5310
rect 26946 5251 28331 5413
rect 30279 5403 31387 5653
rect 28784 5310 29334 5389
rect 30927 5367 30960 5371
rect 30958 5310 31011 5366
rect 31146 5308 31199 5364
rect 13937 451 14487 530
rect 15045 451 15594 530
rect 22615 -995 23566 -415
rect 21773 -2726 21852 -2649
rect 21928 -2730 22007 -2653
rect 21894 -5021 21973 -4943
rect 22063 -5013 22142 -4935
rect 23369 -5018 23448 -4940
rect 23591 -5010 23670 -4932
rect 24094 -5002 24147 -4946
rect 24267 -5002 24320 -4946
<< psubdiff >>
rect -441 11406 40218 11422
rect -441 11405 -151 11406
rect -441 11386 -296 11405
rect -441 -9246 -426 11386
rect -380 11359 -296 11386
rect -250 11360 -151 11405
rect -105 11360 -34 11406
rect 12 11360 83 11406
rect 129 11360 200 11406
rect 246 11360 317 11406
rect 363 11360 434 11406
rect 480 11360 551 11406
rect 597 11360 668 11406
rect 714 11360 785 11406
rect 831 11360 902 11406
rect 948 11360 1019 11406
rect 1065 11360 1136 11406
rect 1182 11360 1253 11406
rect 1299 11360 1370 11406
rect 1416 11360 1487 11406
rect 1533 11360 1604 11406
rect 1650 11360 1721 11406
rect 1767 11360 1838 11406
rect 1884 11360 1955 11406
rect 2001 11360 2072 11406
rect 2118 11360 2189 11406
rect 2235 11360 2306 11406
rect 2352 11360 2423 11406
rect 2469 11360 2540 11406
rect 2586 11360 2657 11406
rect 2703 11360 2774 11406
rect 2820 11360 2891 11406
rect 2937 11360 3008 11406
rect 3054 11360 3125 11406
rect 3171 11360 3242 11406
rect 3288 11360 3359 11406
rect 3405 11360 3476 11406
rect 3522 11360 3593 11406
rect 3639 11360 3710 11406
rect 3756 11360 3827 11406
rect 3873 11360 3944 11406
rect 3990 11360 4061 11406
rect 4107 11360 4178 11406
rect 4224 11360 4295 11406
rect 4341 11360 4412 11406
rect 4458 11360 4529 11406
rect 4575 11360 4646 11406
rect 4692 11360 4763 11406
rect 4809 11360 4880 11406
rect 4926 11360 4997 11406
rect 5043 11360 5114 11406
rect 5160 11360 5231 11406
rect 5277 11360 5348 11406
rect 5394 11360 5465 11406
rect 5511 11360 5582 11406
rect 5628 11360 5699 11406
rect 5745 11360 5816 11406
rect 5862 11360 5933 11406
rect 5979 11360 6050 11406
rect 6096 11360 6167 11406
rect 6213 11360 6284 11406
rect 6330 11360 6401 11406
rect 6447 11360 6518 11406
rect 6564 11360 6635 11406
rect 6681 11360 6752 11406
rect 6798 11360 6869 11406
rect 6915 11360 6986 11406
rect 7032 11360 7103 11406
rect 7149 11360 7220 11406
rect 7266 11360 7337 11406
rect 7383 11360 7454 11406
rect 7500 11360 7571 11406
rect 7617 11360 7688 11406
rect 7734 11360 7805 11406
rect 7851 11360 7922 11406
rect 7968 11360 8039 11406
rect 8085 11360 8156 11406
rect 8202 11360 8273 11406
rect 8319 11360 8390 11406
rect 8436 11360 8507 11406
rect 8553 11360 8624 11406
rect 8670 11360 8741 11406
rect 8787 11360 8858 11406
rect 8904 11360 8975 11406
rect 9021 11360 9092 11406
rect 9138 11360 9209 11406
rect 9255 11360 9326 11406
rect 9372 11360 9443 11406
rect 9489 11360 9560 11406
rect 9606 11360 9677 11406
rect 9723 11360 9794 11406
rect 9840 11360 9911 11406
rect 9957 11360 10028 11406
rect 10074 11360 10145 11406
rect 10191 11360 10262 11406
rect 10308 11360 10379 11406
rect 10425 11360 10496 11406
rect 10542 11360 10613 11406
rect 10659 11360 10730 11406
rect 10776 11360 10847 11406
rect 10893 11360 10964 11406
rect 11010 11360 11081 11406
rect 11127 11360 11198 11406
rect 11244 11360 11315 11406
rect 11361 11360 11432 11406
rect 11478 11360 11549 11406
rect 11595 11360 11666 11406
rect 11712 11360 11783 11406
rect 11829 11360 11900 11406
rect 11946 11360 12017 11406
rect 12063 11360 12134 11406
rect 12180 11360 12251 11406
rect 12297 11360 12368 11406
rect 12414 11360 12485 11406
rect 12531 11360 12602 11406
rect 12648 11360 12719 11406
rect 12765 11360 12836 11406
rect 12882 11360 12953 11406
rect 12999 11360 13070 11406
rect 13116 11360 13187 11406
rect 13233 11360 13304 11406
rect 13350 11360 13421 11406
rect 13467 11360 13538 11406
rect 13584 11360 13655 11406
rect 13701 11360 13772 11406
rect 13818 11360 13889 11406
rect 13935 11360 14006 11406
rect 14052 11360 14123 11406
rect 14169 11360 14240 11406
rect 14286 11360 14357 11406
rect 14403 11360 14474 11406
rect 14520 11360 14591 11406
rect 14637 11360 14708 11406
rect 14754 11360 14825 11406
rect 14871 11360 14942 11406
rect 14988 11360 15059 11406
rect 15105 11360 15176 11406
rect 15222 11360 15293 11406
rect 15339 11360 15410 11406
rect 15456 11360 15527 11406
rect 15573 11360 15644 11406
rect 15690 11360 15761 11406
rect 15807 11360 15878 11406
rect 15924 11360 15995 11406
rect 16041 11360 16112 11406
rect 16158 11360 16229 11406
rect 16275 11360 16346 11406
rect 16392 11360 16463 11406
rect 16509 11360 16580 11406
rect 16626 11360 16697 11406
rect 16743 11360 16814 11406
rect 16860 11360 16931 11406
rect 16977 11360 17048 11406
rect 17094 11360 17165 11406
rect 17211 11360 17282 11406
rect 17328 11360 17399 11406
rect 17445 11360 17516 11406
rect 17562 11360 17633 11406
rect 17679 11360 17750 11406
rect 17796 11360 17867 11406
rect 17913 11360 17984 11406
rect 18030 11360 18101 11406
rect 18147 11360 18218 11406
rect 18264 11360 18335 11406
rect 18381 11360 18452 11406
rect 18498 11360 18569 11406
rect 18615 11360 18686 11406
rect 18732 11360 18803 11406
rect 18849 11360 18920 11406
rect 18966 11360 19037 11406
rect 19083 11360 19154 11406
rect 19200 11360 19271 11406
rect 19317 11360 19388 11406
rect 19434 11360 19505 11406
rect 19551 11360 19622 11406
rect 19668 11360 19739 11406
rect 19785 11360 19856 11406
rect 19902 11360 19973 11406
rect 20019 11360 20090 11406
rect 20136 11360 20207 11406
rect 20253 11360 20324 11406
rect 20370 11360 20441 11406
rect 20487 11360 20558 11406
rect 20604 11360 20675 11406
rect 20721 11360 20792 11406
rect 20838 11360 20909 11406
rect 20955 11360 21026 11406
rect 21072 11360 21143 11406
rect 21189 11360 21260 11406
rect 21306 11360 21377 11406
rect 21423 11360 21494 11406
rect 21540 11360 21611 11406
rect 21657 11360 21728 11406
rect 21774 11360 21845 11406
rect 21891 11360 21962 11406
rect 22008 11360 22079 11406
rect 22125 11360 22196 11406
rect 22242 11360 22313 11406
rect 22359 11360 22430 11406
rect 22476 11360 22547 11406
rect 22593 11360 22664 11406
rect 22710 11360 22781 11406
rect 22827 11360 22898 11406
rect 22944 11360 23015 11406
rect 23061 11360 23132 11406
rect 23178 11360 23249 11406
rect 23295 11360 23366 11406
rect 23412 11360 23483 11406
rect 23529 11360 23600 11406
rect 23646 11360 23717 11406
rect 23763 11360 23834 11406
rect 23880 11360 23951 11406
rect 23997 11360 24068 11406
rect 24114 11360 24185 11406
rect 24231 11360 24302 11406
rect 24348 11360 24419 11406
rect 24465 11360 24536 11406
rect 24582 11360 24653 11406
rect 24699 11360 24770 11406
rect 24816 11360 24887 11406
rect 24933 11360 25004 11406
rect 25050 11360 25121 11406
rect 25167 11360 25238 11406
rect 25284 11360 25355 11406
rect 25401 11360 25472 11406
rect 25518 11360 25589 11406
rect 25635 11360 25706 11406
rect 25752 11360 25823 11406
rect 25869 11360 25940 11406
rect 25986 11360 26057 11406
rect 26103 11360 26174 11406
rect 26220 11360 26291 11406
rect 26337 11360 26408 11406
rect 26454 11360 26525 11406
rect 26571 11360 26642 11406
rect 26688 11360 26759 11406
rect 26805 11360 26876 11406
rect 26922 11360 26993 11406
rect 27039 11360 27110 11406
rect 27156 11360 27227 11406
rect 27273 11360 27344 11406
rect 27390 11360 27461 11406
rect 27507 11360 27578 11406
rect 27624 11360 27695 11406
rect 27741 11360 27812 11406
rect 27858 11360 27929 11406
rect 27975 11360 28046 11406
rect 28092 11360 28163 11406
rect 28209 11360 28280 11406
rect 28326 11360 28397 11406
rect 28443 11360 28514 11406
rect 28560 11360 28631 11406
rect 28677 11360 28748 11406
rect 28794 11360 28865 11406
rect 28911 11360 28982 11406
rect 29028 11360 29099 11406
rect 29145 11360 29216 11406
rect 29262 11360 29333 11406
rect 29379 11360 29450 11406
rect 29496 11360 29567 11406
rect 29613 11360 29684 11406
rect 29730 11360 29801 11406
rect 29847 11360 29918 11406
rect 29964 11360 30035 11406
rect 30081 11360 30152 11406
rect 30198 11360 30269 11406
rect 30315 11360 30386 11406
rect 30432 11360 30503 11406
rect 30549 11360 30620 11406
rect 30666 11360 30737 11406
rect 30783 11360 30854 11406
rect 30900 11360 30971 11406
rect 31017 11360 31088 11406
rect 31134 11360 31205 11406
rect 31251 11360 31322 11406
rect 31368 11360 31439 11406
rect 31485 11360 31556 11406
rect 31602 11360 31673 11406
rect 31719 11360 31790 11406
rect 31836 11360 31907 11406
rect 31953 11360 32024 11406
rect 32070 11360 32141 11406
rect 32187 11360 32258 11406
rect 32304 11360 32375 11406
rect 32421 11360 32492 11406
rect 32538 11360 32609 11406
rect 32655 11360 32726 11406
rect 32772 11360 32843 11406
rect 32889 11360 32960 11406
rect 33006 11360 33077 11406
rect 33123 11360 33194 11406
rect 33240 11360 33311 11406
rect 33357 11360 33428 11406
rect 33474 11360 33545 11406
rect 33591 11360 33662 11406
rect 33708 11360 33779 11406
rect 33825 11360 33896 11406
rect 33942 11360 34013 11406
rect 34059 11360 34130 11406
rect 34176 11360 34247 11406
rect 34293 11360 34364 11406
rect 34410 11360 34481 11406
rect 34527 11360 34598 11406
rect 34644 11360 34715 11406
rect 34761 11360 34832 11406
rect 34878 11360 34949 11406
rect 34995 11360 35066 11406
rect 35112 11360 35183 11406
rect 35229 11360 35300 11406
rect 35346 11360 35417 11406
rect 35463 11360 35534 11406
rect 35580 11360 35651 11406
rect 35697 11360 35768 11406
rect 35814 11360 35885 11406
rect 35931 11360 36002 11406
rect 36048 11360 36119 11406
rect 36165 11360 36236 11406
rect 36282 11360 36353 11406
rect 36399 11360 36470 11406
rect 36516 11360 36587 11406
rect 36633 11360 36704 11406
rect 36750 11360 36821 11406
rect 36867 11360 36938 11406
rect 36984 11360 37055 11406
rect 37101 11360 37172 11406
rect 37218 11360 37289 11406
rect 37335 11360 37406 11406
rect 37452 11360 37523 11406
rect 37569 11360 37640 11406
rect 37686 11360 37757 11406
rect 37803 11360 37874 11406
rect 37920 11360 37991 11406
rect 38037 11360 38108 11406
rect 38154 11360 38225 11406
rect 38271 11360 38342 11406
rect 38388 11360 38459 11406
rect 38505 11360 38576 11406
rect 38622 11360 38693 11406
rect 38739 11360 38810 11406
rect 38856 11360 38927 11406
rect 38973 11360 39044 11406
rect 39090 11360 39161 11406
rect 39207 11360 39278 11406
rect 39324 11360 39395 11406
rect 39441 11360 39512 11406
rect 39558 11360 39629 11406
rect 39675 11360 39746 11406
rect 39792 11360 39863 11406
rect 39909 11360 39980 11406
rect 40026 11360 40096 11406
rect 40142 11360 40218 11406
rect -250 11359 40218 11360
rect -380 11344 40218 11359
rect -380 -9246 -341 11344
rect 40117 11232 40218 11344
rect -441 -9288 -341 -9246
rect 40117 -9212 40132 11232
rect 40178 -9212 40218 11232
rect 40117 -9288 40218 -9212
rect -441 -9304 40218 -9288
rect -441 -9350 -426 -9304
rect -185 -9350 -36 -9304
rect 40054 -9350 40132 -9304
rect 40178 -9350 40218 -9304
rect -441 -9366 40218 -9350
<< nsubdiff >>
rect 498 10526 618 10604
rect 727 10526 845 10605
rect 13937 5668 14487 5747
rect 15045 5668 15595 5747
rect 389 5310 939 5390
rect 28784 5310 29334 5389
rect 762 5309 939 5310
rect 13937 451 14487 530
rect 15045 451 15594 530
<< psubdiffcont >>
rect -426 -9246 -380 11386
rect -296 11359 -250 11405
rect -151 11360 -105 11406
rect -34 11360 12 11406
rect 83 11360 129 11406
rect 200 11360 246 11406
rect 317 11360 363 11406
rect 434 11360 480 11406
rect 551 11360 597 11406
rect 668 11360 714 11406
rect 785 11360 831 11406
rect 902 11360 948 11406
rect 1019 11360 1065 11406
rect 1136 11360 1182 11406
rect 1253 11360 1299 11406
rect 1370 11360 1416 11406
rect 1487 11360 1533 11406
rect 1604 11360 1650 11406
rect 1721 11360 1767 11406
rect 1838 11360 1884 11406
rect 1955 11360 2001 11406
rect 2072 11360 2118 11406
rect 2189 11360 2235 11406
rect 2306 11360 2352 11406
rect 2423 11360 2469 11406
rect 2540 11360 2586 11406
rect 2657 11360 2703 11406
rect 2774 11360 2820 11406
rect 2891 11360 2937 11406
rect 3008 11360 3054 11406
rect 3125 11360 3171 11406
rect 3242 11360 3288 11406
rect 3359 11360 3405 11406
rect 3476 11360 3522 11406
rect 3593 11360 3639 11406
rect 3710 11360 3756 11406
rect 3827 11360 3873 11406
rect 3944 11360 3990 11406
rect 4061 11360 4107 11406
rect 4178 11360 4224 11406
rect 4295 11360 4341 11406
rect 4412 11360 4458 11406
rect 4529 11360 4575 11406
rect 4646 11360 4692 11406
rect 4763 11360 4809 11406
rect 4880 11360 4926 11406
rect 4997 11360 5043 11406
rect 5114 11360 5160 11406
rect 5231 11360 5277 11406
rect 5348 11360 5394 11406
rect 5465 11360 5511 11406
rect 5582 11360 5628 11406
rect 5699 11360 5745 11406
rect 5816 11360 5862 11406
rect 5933 11360 5979 11406
rect 6050 11360 6096 11406
rect 6167 11360 6213 11406
rect 6284 11360 6330 11406
rect 6401 11360 6447 11406
rect 6518 11360 6564 11406
rect 6635 11360 6681 11406
rect 6752 11360 6798 11406
rect 6869 11360 6915 11406
rect 6986 11360 7032 11406
rect 7103 11360 7149 11406
rect 7220 11360 7266 11406
rect 7337 11360 7383 11406
rect 7454 11360 7500 11406
rect 7571 11360 7617 11406
rect 7688 11360 7734 11406
rect 7805 11360 7851 11406
rect 7922 11360 7968 11406
rect 8039 11360 8085 11406
rect 8156 11360 8202 11406
rect 8273 11360 8319 11406
rect 8390 11360 8436 11406
rect 8507 11360 8553 11406
rect 8624 11360 8670 11406
rect 8741 11360 8787 11406
rect 8858 11360 8904 11406
rect 8975 11360 9021 11406
rect 9092 11360 9138 11406
rect 9209 11360 9255 11406
rect 9326 11360 9372 11406
rect 9443 11360 9489 11406
rect 9560 11360 9606 11406
rect 9677 11360 9723 11406
rect 9794 11360 9840 11406
rect 9911 11360 9957 11406
rect 10028 11360 10074 11406
rect 10145 11360 10191 11406
rect 10262 11360 10308 11406
rect 10379 11360 10425 11406
rect 10496 11360 10542 11406
rect 10613 11360 10659 11406
rect 10730 11360 10776 11406
rect 10847 11360 10893 11406
rect 10964 11360 11010 11406
rect 11081 11360 11127 11406
rect 11198 11360 11244 11406
rect 11315 11360 11361 11406
rect 11432 11360 11478 11406
rect 11549 11360 11595 11406
rect 11666 11360 11712 11406
rect 11783 11360 11829 11406
rect 11900 11360 11946 11406
rect 12017 11360 12063 11406
rect 12134 11360 12180 11406
rect 12251 11360 12297 11406
rect 12368 11360 12414 11406
rect 12485 11360 12531 11406
rect 12602 11360 12648 11406
rect 12719 11360 12765 11406
rect 12836 11360 12882 11406
rect 12953 11360 12999 11406
rect 13070 11360 13116 11406
rect 13187 11360 13233 11406
rect 13304 11360 13350 11406
rect 13421 11360 13467 11406
rect 13538 11360 13584 11406
rect 13655 11360 13701 11406
rect 13772 11360 13818 11406
rect 13889 11360 13935 11406
rect 14006 11360 14052 11406
rect 14123 11360 14169 11406
rect 14240 11360 14286 11406
rect 14357 11360 14403 11406
rect 14474 11360 14520 11406
rect 14591 11360 14637 11406
rect 14708 11360 14754 11406
rect 14825 11360 14871 11406
rect 14942 11360 14988 11406
rect 15059 11360 15105 11406
rect 15176 11360 15222 11406
rect 15293 11360 15339 11406
rect 15410 11360 15456 11406
rect 15527 11360 15573 11406
rect 15644 11360 15690 11406
rect 15761 11360 15807 11406
rect 15878 11360 15924 11406
rect 15995 11360 16041 11406
rect 16112 11360 16158 11406
rect 16229 11360 16275 11406
rect 16346 11360 16392 11406
rect 16463 11360 16509 11406
rect 16580 11360 16626 11406
rect 16697 11360 16743 11406
rect 16814 11360 16860 11406
rect 16931 11360 16977 11406
rect 17048 11360 17094 11406
rect 17165 11360 17211 11406
rect 17282 11360 17328 11406
rect 17399 11360 17445 11406
rect 17516 11360 17562 11406
rect 17633 11360 17679 11406
rect 17750 11360 17796 11406
rect 17867 11360 17913 11406
rect 17984 11360 18030 11406
rect 18101 11360 18147 11406
rect 18218 11360 18264 11406
rect 18335 11360 18381 11406
rect 18452 11360 18498 11406
rect 18569 11360 18615 11406
rect 18686 11360 18732 11406
rect 18803 11360 18849 11406
rect 18920 11360 18966 11406
rect 19037 11360 19083 11406
rect 19154 11360 19200 11406
rect 19271 11360 19317 11406
rect 19388 11360 19434 11406
rect 19505 11360 19551 11406
rect 19622 11360 19668 11406
rect 19739 11360 19785 11406
rect 19856 11360 19902 11406
rect 19973 11360 20019 11406
rect 20090 11360 20136 11406
rect 20207 11360 20253 11406
rect 20324 11360 20370 11406
rect 20441 11360 20487 11406
rect 20558 11360 20604 11406
rect 20675 11360 20721 11406
rect 20792 11360 20838 11406
rect 20909 11360 20955 11406
rect 21026 11360 21072 11406
rect 21143 11360 21189 11406
rect 21260 11360 21306 11406
rect 21377 11360 21423 11406
rect 21494 11360 21540 11406
rect 21611 11360 21657 11406
rect 21728 11360 21774 11406
rect 21845 11360 21891 11406
rect 21962 11360 22008 11406
rect 22079 11360 22125 11406
rect 22196 11360 22242 11406
rect 22313 11360 22359 11406
rect 22430 11360 22476 11406
rect 22547 11360 22593 11406
rect 22664 11360 22710 11406
rect 22781 11360 22827 11406
rect 22898 11360 22944 11406
rect 23015 11360 23061 11406
rect 23132 11360 23178 11406
rect 23249 11360 23295 11406
rect 23366 11360 23412 11406
rect 23483 11360 23529 11406
rect 23600 11360 23646 11406
rect 23717 11360 23763 11406
rect 23834 11360 23880 11406
rect 23951 11360 23997 11406
rect 24068 11360 24114 11406
rect 24185 11360 24231 11406
rect 24302 11360 24348 11406
rect 24419 11360 24465 11406
rect 24536 11360 24582 11406
rect 24653 11360 24699 11406
rect 24770 11360 24816 11406
rect 24887 11360 24933 11406
rect 25004 11360 25050 11406
rect 25121 11360 25167 11406
rect 25238 11360 25284 11406
rect 25355 11360 25401 11406
rect 25472 11360 25518 11406
rect 25589 11360 25635 11406
rect 25706 11360 25752 11406
rect 25823 11360 25869 11406
rect 25940 11360 25986 11406
rect 26057 11360 26103 11406
rect 26174 11360 26220 11406
rect 26291 11360 26337 11406
rect 26408 11360 26454 11406
rect 26525 11360 26571 11406
rect 26642 11360 26688 11406
rect 26759 11360 26805 11406
rect 26876 11360 26922 11406
rect 26993 11360 27039 11406
rect 27110 11360 27156 11406
rect 27227 11360 27273 11406
rect 27344 11360 27390 11406
rect 27461 11360 27507 11406
rect 27578 11360 27624 11406
rect 27695 11360 27741 11406
rect 27812 11360 27858 11406
rect 27929 11360 27975 11406
rect 28046 11360 28092 11406
rect 28163 11360 28209 11406
rect 28280 11360 28326 11406
rect 28397 11360 28443 11406
rect 28514 11360 28560 11406
rect 28631 11360 28677 11406
rect 28748 11360 28794 11406
rect 28865 11360 28911 11406
rect 28982 11360 29028 11406
rect 29099 11360 29145 11406
rect 29216 11360 29262 11406
rect 29333 11360 29379 11406
rect 29450 11360 29496 11406
rect 29567 11360 29613 11406
rect 29684 11360 29730 11406
rect 29801 11360 29847 11406
rect 29918 11360 29964 11406
rect 30035 11360 30081 11406
rect 30152 11360 30198 11406
rect 30269 11360 30315 11406
rect 30386 11360 30432 11406
rect 30503 11360 30549 11406
rect 30620 11360 30666 11406
rect 30737 11360 30783 11406
rect 30854 11360 30900 11406
rect 30971 11360 31017 11406
rect 31088 11360 31134 11406
rect 31205 11360 31251 11406
rect 31322 11360 31368 11406
rect 31439 11360 31485 11406
rect 31556 11360 31602 11406
rect 31673 11360 31719 11406
rect 31790 11360 31836 11406
rect 31907 11360 31953 11406
rect 32024 11360 32070 11406
rect 32141 11360 32187 11406
rect 32258 11360 32304 11406
rect 32375 11360 32421 11406
rect 32492 11360 32538 11406
rect 32609 11360 32655 11406
rect 32726 11360 32772 11406
rect 32843 11360 32889 11406
rect 32960 11360 33006 11406
rect 33077 11360 33123 11406
rect 33194 11360 33240 11406
rect 33311 11360 33357 11406
rect 33428 11360 33474 11406
rect 33545 11360 33591 11406
rect 33662 11360 33708 11406
rect 33779 11360 33825 11406
rect 33896 11360 33942 11406
rect 34013 11360 34059 11406
rect 34130 11360 34176 11406
rect 34247 11360 34293 11406
rect 34364 11360 34410 11406
rect 34481 11360 34527 11406
rect 34598 11360 34644 11406
rect 34715 11360 34761 11406
rect 34832 11360 34878 11406
rect 34949 11360 34995 11406
rect 35066 11360 35112 11406
rect 35183 11360 35229 11406
rect 35300 11360 35346 11406
rect 35417 11360 35463 11406
rect 35534 11360 35580 11406
rect 35651 11360 35697 11406
rect 35768 11360 35814 11406
rect 35885 11360 35931 11406
rect 36002 11360 36048 11406
rect 36119 11360 36165 11406
rect 36236 11360 36282 11406
rect 36353 11360 36399 11406
rect 36470 11360 36516 11406
rect 36587 11360 36633 11406
rect 36704 11360 36750 11406
rect 36821 11360 36867 11406
rect 36938 11360 36984 11406
rect 37055 11360 37101 11406
rect 37172 11360 37218 11406
rect 37289 11360 37335 11406
rect 37406 11360 37452 11406
rect 37523 11360 37569 11406
rect 37640 11360 37686 11406
rect 37757 11360 37803 11406
rect 37874 11360 37920 11406
rect 37991 11360 38037 11406
rect 38108 11360 38154 11406
rect 38225 11360 38271 11406
rect 38342 11360 38388 11406
rect 38459 11360 38505 11406
rect 38576 11360 38622 11406
rect 38693 11360 38739 11406
rect 38810 11360 38856 11406
rect 38927 11360 38973 11406
rect 39044 11360 39090 11406
rect 39161 11360 39207 11406
rect 39278 11360 39324 11406
rect 39395 11360 39441 11406
rect 39512 11360 39558 11406
rect 39629 11360 39675 11406
rect 39746 11360 39792 11406
rect 39863 11360 39909 11406
rect 39980 11360 40026 11406
rect 40096 11360 40142 11406
rect 40132 -9212 40178 11232
rect -426 -9350 -185 -9304
rect -36 -9350 40054 -9304
rect 40132 -9350 40178 -9304
<< metal1 >>
rect 22622 12122 23188 12127
rect 22622 12081 23189 12122
rect 22622 12075 22921 12081
rect 22622 12072 22779 12075
rect 22622 12020 22655 12072
rect 22707 12023 22779 12072
rect 22831 12029 22921 12075
rect 22973 12079 23189 12081
rect 22973 12029 23065 12079
rect 22831 12027 23065 12029
rect 23117 12027 23189 12079
rect 22831 12023 23189 12027
rect 22707 12020 23189 12023
rect 4966 12006 5532 12011
rect 4966 11965 5533 12006
rect 4966 11959 5265 11965
rect 4966 11956 5123 11959
rect 4966 11904 4999 11956
rect 5051 11907 5123 11956
rect 5175 11913 5265 11959
rect 5317 11963 5533 11965
rect 5317 11913 5409 11963
rect 5175 11911 5409 11913
rect 5461 11911 5533 11963
rect 5175 11907 5533 11911
rect 5051 11904 5533 11907
rect 4966 11848 5533 11904
rect 4966 11846 5262 11848
rect 4966 11841 5122 11846
rect 4966 11789 4995 11841
rect 5047 11794 5122 11841
rect 5174 11796 5262 11846
rect 5314 11844 5533 11848
rect 5314 11796 5403 11844
rect 5174 11794 5403 11796
rect 5047 11792 5403 11794
rect 5455 11792 5533 11844
rect 5047 11789 5533 11792
rect 4966 11762 5533 11789
rect 15099 11996 15665 12001
rect 15099 11955 15666 11996
rect 15099 11949 15398 11955
rect 15099 11946 15256 11949
rect 15099 11894 15132 11946
rect 15184 11897 15256 11946
rect 15308 11903 15398 11949
rect 15450 11953 15666 11955
rect 15450 11903 15542 11953
rect 15308 11901 15542 11903
rect 15594 11901 15666 11953
rect 15308 11897 15666 11901
rect 15184 11894 15666 11897
rect 15099 11838 15666 11894
rect 22622 11964 23189 12020
rect 22622 11962 22918 11964
rect 22622 11957 22778 11962
rect 22622 11905 22651 11957
rect 22703 11910 22778 11957
rect 22830 11912 22918 11962
rect 22970 11960 23189 11964
rect 22970 11912 23059 11960
rect 22830 11910 23059 11912
rect 22703 11908 23059 11910
rect 23111 11908 23189 11960
rect 22703 11905 23189 11908
rect 22622 11878 23189 11905
rect 15099 11836 15395 11838
rect 15099 11831 15255 11836
rect 11263 11774 11829 11785
rect 11262 11744 11829 11774
rect 15099 11779 15128 11831
rect 15180 11784 15255 11831
rect 15307 11786 15395 11836
rect 15447 11834 15666 11838
rect 15447 11786 15536 11834
rect 15307 11784 15536 11786
rect 15180 11782 15536 11784
rect 15588 11782 15666 11834
rect 32982 11792 33548 11803
rect 15180 11779 15666 11782
rect 15099 11752 15666 11779
rect 32981 11762 33548 11792
rect 32981 11756 33280 11762
rect 32981 11753 33138 11756
rect 11262 11738 11561 11744
rect 11262 11735 11419 11738
rect 11262 11683 11295 11735
rect 11347 11686 11419 11735
rect 11471 11692 11561 11738
rect 11613 11742 11829 11744
rect 11613 11692 11705 11742
rect 11471 11690 11705 11692
rect 11757 11690 11829 11742
rect 19128 11738 19694 11749
rect 11471 11686 11829 11690
rect 11347 11683 11829 11686
rect 1604 11661 2170 11672
rect 1603 11631 2170 11661
rect 1603 11625 1902 11631
rect 1603 11622 1760 11625
rect 1603 11570 1636 11622
rect 1688 11573 1760 11622
rect 1812 11579 1902 11625
rect 1954 11629 2170 11631
rect 1954 11579 2046 11629
rect 1812 11577 2046 11579
rect 2098 11577 2170 11629
rect 1812 11573 2170 11577
rect 1688 11570 2170 11573
rect 1603 11514 2170 11570
rect 11262 11627 11829 11683
rect 11262 11625 11558 11627
rect 11262 11620 11418 11625
rect 11262 11568 11291 11620
rect 11343 11573 11418 11620
rect 11470 11575 11558 11625
rect 11610 11623 11829 11627
rect 11610 11575 11699 11623
rect 11470 11573 11699 11575
rect 11343 11571 11699 11573
rect 11751 11571 11829 11623
rect 11343 11568 11829 11571
rect 11262 11551 11829 11568
rect 1603 11512 1899 11514
rect 1603 11507 1759 11512
rect 1603 11455 1632 11507
rect 1684 11460 1759 11507
rect 1811 11462 1899 11512
rect 1951 11510 2170 11514
rect 1951 11462 2040 11510
rect 1811 11460 2040 11462
rect 1684 11458 2040 11460
rect 2092 11458 2170 11510
rect 1684 11455 2170 11458
rect 1603 11422 2170 11455
rect 11260 11422 11829 11551
rect 19127 11708 19694 11738
rect 26109 11720 26675 11731
rect 19127 11702 19426 11708
rect 19127 11699 19284 11702
rect 19127 11647 19160 11699
rect 19212 11650 19284 11699
rect 19336 11656 19426 11702
rect 19478 11706 19694 11708
rect 19478 11656 19570 11706
rect 19336 11654 19570 11656
rect 19622 11654 19694 11706
rect 19336 11650 19694 11654
rect 19212 11647 19694 11650
rect 19127 11591 19694 11647
rect 19127 11589 19423 11591
rect 19127 11584 19283 11589
rect 19127 11532 19156 11584
rect 19208 11537 19283 11584
rect 19335 11539 19423 11589
rect 19475 11587 19694 11591
rect 19475 11539 19564 11587
rect 19335 11537 19564 11539
rect 19208 11535 19564 11537
rect 19616 11535 19694 11587
rect 19208 11532 19694 11535
rect 19127 11422 19694 11532
rect 26108 11690 26675 11720
rect 26108 11684 26407 11690
rect 26108 11681 26265 11684
rect 26108 11629 26141 11681
rect 26193 11632 26265 11681
rect 26317 11638 26407 11684
rect 26459 11688 26675 11690
rect 26459 11638 26551 11688
rect 26317 11636 26551 11638
rect 26603 11636 26675 11688
rect 26317 11632 26675 11636
rect 26193 11629 26675 11632
rect 26108 11573 26675 11629
rect 26108 11571 26404 11573
rect 26108 11566 26264 11571
rect 26108 11514 26137 11566
rect 26189 11519 26264 11566
rect 26316 11521 26404 11571
rect 26456 11569 26675 11573
rect 26456 11521 26545 11569
rect 26316 11519 26545 11521
rect 26189 11517 26545 11519
rect 26597 11517 26675 11569
rect 26189 11514 26675 11517
rect 26108 11422 26675 11514
rect 32981 11701 33014 11753
rect 33066 11704 33138 11753
rect 33190 11710 33280 11756
rect 33332 11760 33548 11762
rect 33332 11710 33424 11760
rect 33190 11708 33424 11710
rect 33476 11708 33548 11760
rect 33190 11704 33548 11708
rect 33066 11701 33548 11704
rect 32981 11645 33548 11701
rect 32981 11643 33277 11645
rect 32981 11638 33137 11643
rect 32981 11586 33010 11638
rect 33062 11591 33137 11638
rect 33189 11593 33277 11643
rect 33329 11641 33548 11645
rect 33329 11593 33418 11641
rect 33189 11591 33418 11593
rect 33062 11589 33418 11591
rect 33470 11589 33548 11641
rect 33062 11586 33548 11589
rect 32981 11422 33548 11586
rect -441 11406 40218 11422
rect -441 11405 -151 11406
rect -441 11386 -296 11405
rect -441 -9246 -426 11386
rect -380 11359 -296 11386
rect -250 11360 -151 11405
rect -105 11360 -34 11406
rect 12 11360 83 11406
rect 129 11360 200 11406
rect 246 11360 317 11406
rect 363 11360 434 11406
rect 480 11360 551 11406
rect 597 11360 668 11406
rect 714 11360 785 11406
rect 831 11360 902 11406
rect 948 11360 1019 11406
rect 1065 11360 1136 11406
rect 1182 11360 1253 11406
rect 1299 11360 1370 11406
rect 1416 11360 1487 11406
rect 1533 11360 1604 11406
rect 1650 11360 1721 11406
rect 1767 11360 1838 11406
rect 1884 11360 1955 11406
rect 2001 11360 2072 11406
rect 2118 11360 2189 11406
rect 2235 11360 2306 11406
rect 2352 11360 2423 11406
rect 2469 11360 2540 11406
rect 2586 11360 2657 11406
rect 2703 11360 2774 11406
rect 2820 11360 2891 11406
rect 2937 11360 3008 11406
rect 3054 11360 3125 11406
rect 3171 11360 3242 11406
rect 3288 11360 3359 11406
rect 3405 11360 3476 11406
rect 3522 11360 3593 11406
rect 3639 11360 3710 11406
rect 3756 11360 3827 11406
rect 3873 11360 3944 11406
rect 3990 11360 4061 11406
rect 4107 11360 4178 11406
rect 4224 11360 4295 11406
rect 4341 11360 4412 11406
rect 4458 11360 4529 11406
rect 4575 11360 4646 11406
rect 4692 11360 4763 11406
rect 4809 11360 4880 11406
rect 4926 11360 4997 11406
rect 5043 11360 5114 11406
rect 5160 11360 5231 11406
rect 5277 11360 5348 11406
rect 5394 11360 5465 11406
rect 5511 11360 5582 11406
rect 5628 11360 5699 11406
rect 5745 11360 5816 11406
rect 5862 11360 5933 11406
rect 5979 11360 6050 11406
rect 6096 11360 6167 11406
rect 6213 11360 6284 11406
rect 6330 11360 6401 11406
rect 6447 11360 6518 11406
rect 6564 11360 6635 11406
rect 6681 11360 6752 11406
rect 6798 11360 6869 11406
rect 6915 11360 6986 11406
rect 7032 11360 7103 11406
rect 7149 11360 7220 11406
rect 7266 11360 7337 11406
rect 7383 11360 7454 11406
rect 7500 11360 7571 11406
rect 7617 11360 7688 11406
rect 7734 11360 7805 11406
rect 7851 11360 7922 11406
rect 7968 11360 8039 11406
rect 8085 11360 8156 11406
rect 8202 11360 8273 11406
rect 8319 11360 8390 11406
rect 8436 11360 8507 11406
rect 8553 11360 8624 11406
rect 8670 11360 8741 11406
rect 8787 11360 8858 11406
rect 8904 11360 8975 11406
rect 9021 11360 9092 11406
rect 9138 11360 9209 11406
rect 9255 11360 9326 11406
rect 9372 11360 9443 11406
rect 9489 11360 9560 11406
rect 9606 11360 9677 11406
rect 9723 11360 9794 11406
rect 9840 11360 9911 11406
rect 9957 11360 10028 11406
rect 10074 11360 10145 11406
rect 10191 11360 10262 11406
rect 10308 11360 10379 11406
rect 10425 11360 10496 11406
rect 10542 11360 10613 11406
rect 10659 11360 10730 11406
rect 10776 11360 10847 11406
rect 10893 11360 10964 11406
rect 11010 11360 11081 11406
rect 11127 11360 11198 11406
rect 11244 11360 11315 11406
rect 11361 11360 11432 11406
rect 11478 11360 11549 11406
rect 11595 11360 11666 11406
rect 11712 11360 11783 11406
rect 11829 11360 11900 11406
rect 11946 11360 12017 11406
rect 12063 11360 12134 11406
rect 12180 11360 12251 11406
rect 12297 11360 12368 11406
rect 12414 11360 12485 11406
rect 12531 11360 12602 11406
rect 12648 11360 12719 11406
rect 12765 11360 12836 11406
rect 12882 11360 12953 11406
rect 12999 11360 13070 11406
rect 13116 11360 13187 11406
rect 13233 11360 13304 11406
rect 13350 11360 13421 11406
rect 13467 11360 13538 11406
rect 13584 11360 13655 11406
rect 13701 11360 13772 11406
rect 13818 11360 13889 11406
rect 13935 11360 14006 11406
rect 14052 11360 14123 11406
rect 14169 11360 14240 11406
rect 14286 11360 14357 11406
rect 14403 11360 14474 11406
rect 14520 11360 14591 11406
rect 14637 11360 14708 11406
rect 14754 11360 14825 11406
rect 14871 11360 14942 11406
rect 14988 11360 15059 11406
rect 15105 11360 15176 11406
rect 15222 11360 15293 11406
rect 15339 11360 15410 11406
rect 15456 11360 15527 11406
rect 15573 11360 15644 11406
rect 15690 11360 15761 11406
rect 15807 11360 15878 11406
rect 15924 11360 15995 11406
rect 16041 11360 16112 11406
rect 16158 11360 16229 11406
rect 16275 11360 16346 11406
rect 16392 11360 16463 11406
rect 16509 11360 16580 11406
rect 16626 11360 16697 11406
rect 16743 11360 16814 11406
rect 16860 11360 16931 11406
rect 16977 11360 17048 11406
rect 17094 11360 17165 11406
rect 17211 11360 17282 11406
rect 17328 11360 17399 11406
rect 17445 11360 17516 11406
rect 17562 11360 17633 11406
rect 17679 11360 17750 11406
rect 17796 11360 17867 11406
rect 17913 11360 17984 11406
rect 18030 11360 18101 11406
rect 18147 11360 18218 11406
rect 18264 11360 18335 11406
rect 18381 11360 18452 11406
rect 18498 11360 18569 11406
rect 18615 11360 18686 11406
rect 18732 11360 18803 11406
rect 18849 11360 18920 11406
rect 18966 11360 19037 11406
rect 19083 11360 19154 11406
rect 19200 11360 19271 11406
rect 19317 11360 19388 11406
rect 19434 11360 19505 11406
rect 19551 11360 19622 11406
rect 19668 11360 19739 11406
rect 19785 11360 19856 11406
rect 19902 11360 19973 11406
rect 20019 11360 20090 11406
rect 20136 11360 20207 11406
rect 20253 11360 20324 11406
rect 20370 11360 20441 11406
rect 20487 11360 20558 11406
rect 20604 11360 20675 11406
rect 20721 11360 20792 11406
rect 20838 11360 20909 11406
rect 20955 11360 21026 11406
rect 21072 11360 21143 11406
rect 21189 11360 21260 11406
rect 21306 11360 21377 11406
rect 21423 11360 21494 11406
rect 21540 11360 21611 11406
rect 21657 11360 21728 11406
rect 21774 11360 21845 11406
rect 21891 11360 21962 11406
rect 22008 11360 22079 11406
rect 22125 11360 22196 11406
rect 22242 11360 22313 11406
rect 22359 11360 22430 11406
rect 22476 11360 22547 11406
rect 22593 11360 22664 11406
rect 22710 11360 22781 11406
rect 22827 11360 22898 11406
rect 22944 11360 23015 11406
rect 23061 11360 23132 11406
rect 23178 11360 23249 11406
rect 23295 11360 23366 11406
rect 23412 11360 23483 11406
rect 23529 11360 23600 11406
rect 23646 11360 23717 11406
rect 23763 11360 23834 11406
rect 23880 11360 23951 11406
rect 23997 11360 24068 11406
rect 24114 11360 24185 11406
rect 24231 11360 24302 11406
rect 24348 11360 24419 11406
rect 24465 11360 24536 11406
rect 24582 11360 24653 11406
rect 24699 11360 24770 11406
rect 24816 11360 24887 11406
rect 24933 11360 25004 11406
rect 25050 11360 25121 11406
rect 25167 11360 25238 11406
rect 25284 11360 25355 11406
rect 25401 11360 25472 11406
rect 25518 11360 25589 11406
rect 25635 11360 25706 11406
rect 25752 11360 25823 11406
rect 25869 11360 25940 11406
rect 25986 11360 26057 11406
rect 26103 11360 26174 11406
rect 26220 11360 26291 11406
rect 26337 11360 26408 11406
rect 26454 11360 26525 11406
rect 26571 11360 26642 11406
rect 26688 11360 26759 11406
rect 26805 11360 26876 11406
rect 26922 11360 26993 11406
rect 27039 11360 27110 11406
rect 27156 11360 27227 11406
rect 27273 11360 27344 11406
rect 27390 11360 27461 11406
rect 27507 11360 27578 11406
rect 27624 11360 27695 11406
rect 27741 11360 27812 11406
rect 27858 11360 27929 11406
rect 27975 11360 28046 11406
rect 28092 11360 28163 11406
rect 28209 11360 28280 11406
rect 28326 11360 28397 11406
rect 28443 11360 28514 11406
rect 28560 11360 28631 11406
rect 28677 11360 28748 11406
rect 28794 11360 28865 11406
rect 28911 11360 28982 11406
rect 29028 11360 29099 11406
rect 29145 11360 29216 11406
rect 29262 11360 29333 11406
rect 29379 11360 29450 11406
rect 29496 11360 29567 11406
rect 29613 11360 29684 11406
rect 29730 11360 29801 11406
rect 29847 11360 29918 11406
rect 29964 11360 30035 11406
rect 30081 11360 30152 11406
rect 30198 11360 30269 11406
rect 30315 11360 30386 11406
rect 30432 11360 30503 11406
rect 30549 11360 30620 11406
rect 30666 11360 30737 11406
rect 30783 11360 30854 11406
rect 30900 11360 30971 11406
rect 31017 11360 31088 11406
rect 31134 11360 31205 11406
rect 31251 11360 31322 11406
rect 31368 11360 31439 11406
rect 31485 11360 31556 11406
rect 31602 11360 31673 11406
rect 31719 11360 31790 11406
rect 31836 11360 31907 11406
rect 31953 11360 32024 11406
rect 32070 11360 32141 11406
rect 32187 11360 32258 11406
rect 32304 11360 32375 11406
rect 32421 11360 32492 11406
rect 32538 11360 32609 11406
rect 32655 11360 32726 11406
rect 32772 11360 32843 11406
rect 32889 11360 32960 11406
rect 33006 11360 33077 11406
rect 33123 11360 33194 11406
rect 33240 11360 33311 11406
rect 33357 11360 33428 11406
rect 33474 11360 33545 11406
rect 33591 11360 33662 11406
rect 33708 11360 33779 11406
rect 33825 11360 33896 11406
rect 33942 11360 34013 11406
rect 34059 11360 34130 11406
rect 34176 11360 34247 11406
rect 34293 11360 34364 11406
rect 34410 11360 34481 11406
rect 34527 11360 34598 11406
rect 34644 11360 34715 11406
rect 34761 11360 34832 11406
rect 34878 11360 34949 11406
rect 34995 11360 35066 11406
rect 35112 11360 35183 11406
rect 35229 11360 35300 11406
rect 35346 11360 35417 11406
rect 35463 11360 35534 11406
rect 35580 11360 35651 11406
rect 35697 11360 35768 11406
rect 35814 11360 35885 11406
rect 35931 11360 36002 11406
rect 36048 11360 36119 11406
rect 36165 11360 36236 11406
rect 36282 11360 36353 11406
rect 36399 11360 36470 11406
rect 36516 11360 36587 11406
rect 36633 11360 36704 11406
rect 36750 11360 36821 11406
rect 36867 11360 36938 11406
rect 36984 11360 37055 11406
rect 37101 11360 37172 11406
rect 37218 11360 37289 11406
rect 37335 11360 37406 11406
rect 37452 11360 37523 11406
rect 37569 11360 37640 11406
rect 37686 11360 37757 11406
rect 37803 11360 37874 11406
rect 37920 11360 37991 11406
rect 38037 11360 38108 11406
rect 38154 11360 38225 11406
rect 38271 11360 38342 11406
rect 38388 11360 38459 11406
rect 38505 11360 38576 11406
rect 38622 11360 38693 11406
rect 38739 11360 38810 11406
rect 38856 11360 38927 11406
rect 38973 11360 39044 11406
rect 39090 11360 39161 11406
rect 39207 11360 39278 11406
rect 39324 11360 39395 11406
rect 39441 11360 39512 11406
rect 39558 11360 39629 11406
rect 39675 11360 39746 11406
rect 39792 11360 39863 11406
rect 39909 11360 39980 11406
rect 40026 11360 40096 11406
rect 40142 11360 40218 11406
rect -250 11359 40218 11360
rect -380 11344 40218 11359
rect -380 -9246 -341 11344
rect 40117 11232 40218 11344
rect 606 10928 840 10942
rect 606 10876 619 10928
rect 671 10876 774 10928
rect 826 10926 840 10928
rect 826 10876 6921 10926
rect 606 10875 6921 10876
rect 606 10862 840 10875
rect 498 10526 618 10604
rect 727 10526 845 10605
rect 1132 10526 1254 10603
rect 5140 10570 5228 10587
rect 5140 10518 5158 10570
rect 5210 10518 5228 10570
rect 5140 10499 5228 10518
rect 38953 10472 39755 10915
rect 38953 10420 38985 10472
rect 39037 10420 39105 10472
rect 39157 10420 39225 10472
rect 39277 10420 39755 10472
rect 38953 10352 39755 10420
rect 38953 10300 38985 10352
rect 39037 10300 39105 10352
rect 39157 10300 39225 10352
rect 39277 10300 39755 10352
rect 38953 10232 39755 10300
rect 38953 10180 38985 10232
rect 39037 10180 39105 10232
rect 39157 10180 39225 10232
rect 39277 10180 39755 10232
rect 38953 10145 39755 10180
rect 1654 9573 1814 9622
rect 155 9204 202 9549
rect 1654 9521 1705 9573
rect 1757 9521 1814 9573
rect 6858 9567 6916 9857
rect 32754 9765 33766 9841
rect 22555 9525 22602 9558
rect 1654 9483 1814 9521
rect 22512 9281 22602 9525
rect 1052 8686 1151 8805
rect 19481 8804 19600 8830
rect 1053 8648 1151 8686
rect 1053 8596 1078 8648
rect 1130 8596 1151 8648
rect 1053 8535 1151 8596
rect 9843 8654 9935 8792
rect 19481 8752 19523 8804
rect 19575 8752 19600 8804
rect 19481 8722 19600 8752
rect 9843 8602 9850 8654
rect 9902 8602 9935 8654
rect 9843 8543 9935 8602
rect 1034 8486 1234 8535
rect 1053 8467 1151 8486
rect 9843 8476 9914 8543
rect 10183 8542 10411 8563
rect 10183 8490 10202 8542
rect 10254 8541 10411 8542
rect 10254 8490 10342 8541
rect 10183 8489 10342 8490
rect 10394 8489 10411 8541
rect 10183 8430 10411 8489
rect 10183 8378 10207 8430
rect 10259 8378 10411 8430
rect 10183 8332 10411 8378
rect 11451 8478 11632 8549
rect 11451 8426 11532 8478
rect 11584 8426 11632 8478
rect 11451 8372 11632 8426
rect 10184 8282 10411 8332
rect 1634 7999 1794 8048
rect 1634 7947 1685 7999
rect 1737 7947 1794 7999
rect 1634 7909 1794 7947
rect 10272 7904 10411 8282
rect 19390 7995 19455 8253
rect 20058 8159 21687 8236
rect 22555 8219 22602 9281
rect 26519 8415 26679 8472
rect 26519 8363 26570 8415
rect 26622 8363 26679 8415
rect 26519 8325 26679 8363
rect 22423 8172 22602 8219
rect 11515 7928 11575 7942
rect 19390 7930 19559 7995
rect 11475 7923 11592 7928
rect 10271 7846 10607 7904
rect 10271 7794 10301 7846
rect 10353 7794 10471 7846
rect 10523 7794 10607 7846
rect 10271 7740 10607 7794
rect 11475 7897 11594 7923
rect 11475 7845 11517 7897
rect 11569 7845 11594 7897
rect 11475 7815 11594 7845
rect 11475 7732 11592 7815
rect 13651 7738 13788 7787
rect 15677 7738 15909 7787
rect 19429 7609 19548 7635
rect 19429 7557 19471 7609
rect 19523 7557 19548 7609
rect 19429 7527 19548 7557
rect 19433 7436 19531 7527
rect 7931 7139 8009 7151
rect 7931 7087 7943 7139
rect 7995 7087 8009 7139
rect 7931 7075 8009 7087
rect 7938 6993 8016 7005
rect 7938 6941 7950 6993
rect 8002 6941 8016 6993
rect 7938 6929 8016 6941
rect 7744 6715 7974 6762
rect 15464 5747 15593 5762
rect 22850 5747 22976 5753
rect 13937 5668 14487 5747
rect 15045 5734 15595 5747
rect 15045 5682 15521 5734
rect 15573 5682 15595 5734
rect 15045 5668 15595 5682
rect 15788 5670 15912 5747
rect 22892 5669 22976 5747
rect 15496 5658 15593 5668
rect 389 5310 939 5390
rect 762 5309 939 5310
rect 5131 5348 5219 5364
rect 5131 5296 5153 5348
rect 5205 5296 5219 5348
rect 28490 5310 28616 5387
rect 30958 5364 31011 5366
rect 31010 5312 31011 5364
rect 30958 5310 31011 5312
rect 31146 5362 31199 5364
rect 31198 5310 31199 5362
rect 31146 5308 31199 5310
rect 5131 5276 5219 5296
rect 6867 4229 6915 4597
rect 22612 4387 22658 4716
rect 29985 4714 30375 4760
rect 6854 4214 6930 4229
rect 6854 4162 6867 4214
rect 6919 4162 6930 4214
rect 6854 4146 6930 4162
rect 6867 4064 6915 4146
rect 6854 4049 6930 4064
rect 6854 3997 6867 4049
rect 6919 3997 6930 4049
rect 6854 3981 6930 3997
rect 6867 3898 6915 3981
rect 19436 3612 19555 3638
rect 19436 3560 19478 3612
rect 19530 3560 19555 3612
rect 19436 3530 19555 3560
rect 9843 3431 9922 3467
rect 9843 3379 9851 3431
rect 9903 3379 9922 3431
rect 1085 3270 1221 3319
rect 9843 3250 9922 3379
rect 28484 3270 28685 3319
rect 11311 3233 11390 3237
rect 11727 3233 11806 3242
rect 11265 3229 11806 3233
rect 11265 3224 11740 3229
rect 11265 3221 11324 3224
rect 11183 3172 11324 3221
rect 11376 3219 11740 3224
rect 11376 3172 11545 3219
rect 11183 3167 11545 3172
rect 11597 3177 11740 3219
rect 11792 3177 11806 3229
rect 11597 3167 11806 3177
rect 11183 3164 11806 3167
rect 11183 3162 11799 3164
rect 3073 3009 3151 3021
rect 3073 2957 3085 3009
rect 3137 2957 3151 3009
rect 3073 2945 3151 2957
rect 3363 3010 3441 3022
rect 3363 2958 3375 3010
rect 3427 2958 3441 3010
rect 3363 2946 3441 2958
rect 1690 2803 1850 2852
rect 1690 2751 1741 2803
rect 1793 2751 1850 2803
rect 1690 2713 1850 2751
rect 11183 2652 11242 3162
rect 11311 3159 11390 3162
rect 11532 3154 11611 3162
rect 11496 2743 11556 2762
rect 11456 2742 11575 2743
rect 11036 2593 11242 2652
rect 11455 2717 11575 2742
rect 11455 2665 11498 2717
rect 11550 2665 11575 2717
rect 11036 2329 11095 2593
rect 11455 2512 11575 2665
rect 26416 2687 26576 2744
rect 26416 2635 26467 2687
rect 26519 2635 26576 2687
rect 26416 2597 26576 2635
rect 13674 2521 13824 2570
rect 15732 2521 15889 2570
rect 11023 2316 11102 2329
rect 11023 2264 11036 2316
rect 11088 2264 11102 2316
rect 11023 2251 11102 2264
rect 11036 2194 11095 2251
rect 11028 2181 11107 2194
rect 11028 2129 11041 2181
rect 11093 2129 11107 2181
rect 11028 2116 11107 2129
rect 11036 2108 11095 2116
rect 28945 1888 29008 1895
rect 28945 1836 28947 1888
rect 28999 1836 29008 1888
rect 28945 1835 29008 1836
rect 29228 1887 29284 1889
rect 29228 1835 29230 1887
rect 29282 1835 29284 1887
rect 29228 1834 29284 1835
rect 21760 1571 21812 1831
rect 7954 1199 8009 1401
rect 15199 530 15283 533
rect 13621 453 13761 530
rect 13937 451 14487 530
rect 15045 517 15594 530
rect 15045 465 15217 517
rect 15269 465 15594 517
rect 15045 451 15594 465
rect 15199 447 15283 451
rect 7651 390 7730 404
rect 7651 338 7663 390
rect 7715 338 7730 390
rect 7651 326 7730 338
rect 7806 400 7885 405
rect 7806 391 8203 400
rect 7806 339 7818 391
rect 7870 345 8203 391
rect 7870 339 7885 345
rect 7806 327 7885 339
rect 4500 113 4578 125
rect -210 13 829 76
rect 4500 61 4512 113
rect 4564 61 4578 113
rect 4500 49 4578 61
rect 6030 27 6093 33
rect -210 -8918 -147 13
rect 522 -192 600 -180
rect 522 -244 534 -192
rect 586 -244 600 -192
rect 522 -256 600 -244
rect 766 -285 829 13
rect 6025 13 6104 27
rect 6025 -39 6037 13
rect 6089 -39 6104 13
rect 21725 0 23055 52
rect 2356 -53 2434 -41
rect 6025 -51 6104 -39
rect 2356 -105 2368 -53
rect 2420 -105 2434 -53
rect 2967 -75 3045 -63
rect 2356 -117 2434 -105
rect 2543 -116 2621 -104
rect 2543 -168 2555 -116
rect 2607 -168 2621 -116
rect 2967 -127 2979 -75
rect 3031 -127 3045 -75
rect 2967 -139 3045 -127
rect 3171 -77 3249 -65
rect 3171 -129 3183 -77
rect 3235 -129 3249 -77
rect 3171 -141 3249 -129
rect 2543 -180 2621 -168
rect 6030 -174 6093 -51
rect 19485 -149 19531 -68
rect 3699 -237 6093 -174
rect 19480 -163 19559 -149
rect 19480 -215 19492 -163
rect 19544 -215 19559 -163
rect 19480 -227 19559 -215
rect 3699 -285 3762 -237
rect 518 -359 596 -347
rect 766 -348 3762 -285
rect 518 -411 530 -359
rect 582 -411 596 -359
rect 6030 -353 6093 -237
rect 518 -423 596 -411
rect 3916 -379 3994 -367
rect 3916 -431 3928 -379
rect 3980 -431 3994 -379
rect 3916 -443 3994 -431
rect 4139 -375 4217 -363
rect 4139 -427 4151 -375
rect 4203 -427 4217 -375
rect 4139 -439 4217 -427
rect 6030 -367 6112 -353
rect 6030 -419 6045 -367
rect 6097 -419 6112 -367
rect 6030 -431 6112 -419
rect 19485 -426 19531 -227
rect 6030 -476 6093 -431
rect 22708 -912 22802 -911
rect 22674 -957 22802 -912
rect 22674 -1049 22720 -957
rect 3812 -1209 3891 -1195
rect 316 -1348 395 -1334
rect 316 -1400 328 -1348
rect 380 -1400 395 -1348
rect 316 -1412 395 -1400
rect 2716 -1428 2762 -1216
rect 3812 -1261 3824 -1209
rect 3876 -1261 3891 -1209
rect 7400 -1205 7494 -1151
rect 6219 -1248 6265 -1216
rect 3812 -1273 3891 -1261
rect 6210 -1262 6289 -1248
rect 6210 -1314 6222 -1262
rect 6274 -1314 6289 -1262
rect 6210 -1326 6289 -1314
rect 7400 -1257 7427 -1205
rect 7479 -1257 7494 -1205
rect 22671 -1152 22742 -1140
rect 22671 -1204 22676 -1152
rect 22728 -1204 22742 -1152
rect 22671 -1216 22742 -1204
rect 6219 -1417 6265 -1326
rect 2716 -1442 2802 -1428
rect 2716 -1494 2735 -1442
rect 2787 -1494 2802 -1442
rect 2716 -1506 2802 -1494
rect 6215 -1431 6294 -1417
rect 6215 -1483 6227 -1431
rect 6279 -1483 6294 -1431
rect 6215 -1495 6294 -1483
rect 7400 -1455 7494 -1257
rect 9835 -1233 9914 -1219
rect 9835 -1285 9847 -1233
rect 9899 -1285 9914 -1233
rect 9835 -1297 9914 -1285
rect 22670 -1287 22742 -1275
rect 22670 -1339 22676 -1287
rect 22728 -1339 22742 -1287
rect 22670 -1351 22742 -1339
rect 323 -1532 402 -1518
rect 2716 -1520 2762 -1506
rect 3808 -1515 3887 -1501
rect 323 -1584 335 -1532
rect 387 -1584 402 -1532
rect 3808 -1567 3820 -1515
rect 3872 -1567 3887 -1515
rect 7400 -1507 7419 -1455
rect 7471 -1507 7494 -1455
rect 7400 -1557 7494 -1507
rect 3808 -1579 3887 -1567
rect 323 -1596 402 -1584
rect 1726 -2430 1886 -2381
rect 1726 -2482 1777 -2430
rect 1829 -2482 1886 -2430
rect 4344 -2387 4422 -2375
rect 4344 -2439 4356 -2387
rect 4408 -2439 4422 -2387
rect 4344 -2451 4422 -2439
rect 5238 -2425 6133 -2411
rect 1726 -2520 1886 -2482
rect 5238 -2477 5255 -2425
rect 5307 -2477 5484 -2425
rect 5536 -2477 6133 -2425
rect 5238 -2490 6133 -2477
rect 6054 -2511 6133 -2490
rect 6054 -2530 6534 -2511
rect 6054 -2533 6276 -2530
rect 3796 -2562 3875 -2557
rect 4056 -2562 4135 -2559
rect 3777 -2571 4139 -2562
rect 3777 -2623 3808 -2571
rect 3860 -2573 4139 -2571
rect 3860 -2623 4068 -2573
rect 3777 -2625 4068 -2623
rect 4120 -2625 4139 -2573
rect 6054 -2585 6100 -2533
rect 6152 -2582 6276 -2533
rect 6328 -2535 6534 -2530
rect 6328 -2582 6455 -2535
rect 6152 -2585 6455 -2582
rect 6054 -2587 6455 -2585
rect 6507 -2587 6534 -2535
rect 6054 -2592 6534 -2587
rect 9695 -2542 9773 -2530
rect 9695 -2594 9707 -2542
rect 9759 -2594 9773 -2542
rect 9695 -2606 9773 -2594
rect 9887 -2542 9965 -2530
rect 9887 -2594 9899 -2542
rect 9951 -2594 9965 -2542
rect 9887 -2606 9965 -2594
rect 3777 -2635 4139 -2625
rect 3792 -3029 3858 -2635
rect 4056 -2637 4135 -2635
rect 21773 -2662 21852 -2648
rect 21773 -2714 21785 -2662
rect 21837 -2714 21852 -2662
rect 21773 -2726 21852 -2714
rect 21928 -2666 22007 -2652
rect 21928 -2718 21940 -2666
rect 21992 -2718 22007 -2666
rect 21928 -2730 22007 -2718
rect 11603 -2772 11663 -2753
rect 11563 -2798 11682 -2772
rect 11563 -2850 11605 -2798
rect 11657 -2850 11682 -2798
rect 11563 -2880 11682 -2850
rect 17867 -2819 17946 -2813
rect 18125 -2819 18204 -2813
rect 23003 -2819 23055 0
rect 23480 -137 23559 -125
rect 23480 -189 23493 -137
rect 23545 -189 23559 -137
rect 23480 -202 23559 -189
rect 23485 -294 23531 -202
rect 23481 -306 23560 -294
rect 23481 -358 23494 -306
rect 23546 -358 23560 -306
rect 29985 -318 30031 4714
rect 31368 4284 31467 4331
rect 30204 3865 30482 3880
rect 30204 3813 30303 3865
rect 30355 3813 30482 3865
rect 30204 3790 30482 3813
rect 30204 3709 30294 3790
rect 30204 3657 30221 3709
rect 30273 3657 30294 3709
rect 30204 3578 30294 3657
rect 31420 3107 31467 4284
rect 33690 3374 33766 9765
rect 33690 3298 37314 3374
rect 37238 2972 37314 3298
rect 31692 2006 31786 2029
rect 31692 1954 31709 2006
rect 31761 1954 31786 2006
rect 31692 1941 31786 1954
rect 37119 1851 37200 1867
rect 37119 1799 37133 1851
rect 37185 1799 37200 1851
rect 37119 1782 37200 1799
rect 37354 1853 37435 1869
rect 37354 1801 37368 1853
rect 37420 1801 37435 1853
rect 37354 1784 37435 1801
rect 23481 -371 23560 -358
rect 23485 -430 23531 -371
rect 24011 -379 24479 -333
rect 29985 -364 31134 -318
rect 30469 -449 30548 -435
rect 30469 -501 30481 -449
rect 30533 -501 30548 -449
rect 30469 -513 30548 -501
rect 30666 -442 30745 -428
rect 30666 -494 30678 -442
rect 30730 -494 30745 -442
rect 30666 -506 30745 -494
rect 31088 -904 31134 -364
rect 31762 -436 31841 -422
rect 31762 -488 31774 -436
rect 31826 -488 31841 -436
rect 31762 -500 31841 -488
rect 31948 -434 32027 -420
rect 31948 -486 31960 -434
rect 32012 -486 32027 -434
rect 31948 -498 32027 -486
rect 32241 -504 32314 810
rect 38127 670 38173 1562
rect 32568 624 38173 670
rect 32568 143 32614 624
rect 32557 131 32633 143
rect 32557 79 32569 131
rect 32621 79 32633 131
rect 32557 67 32633 79
rect 32568 -68 32614 67
rect 32548 -80 32624 -68
rect 32548 -132 32560 -80
rect 32612 -132 32624 -80
rect 32548 -144 32624 -132
rect 17867 -2825 23055 -2819
rect 17867 -2877 17880 -2825
rect 17932 -2871 18138 -2825
rect 17932 -2877 17946 -2871
rect 11603 -2882 11663 -2880
rect 17867 -2890 17946 -2877
rect 18125 -2877 18138 -2871
rect 18190 -2871 23055 -2825
rect 23333 -966 23531 -920
rect 31001 -950 31135 -904
rect 23333 -2827 23379 -966
rect 32518 -1138 32567 -1083
rect 32505 -1150 32581 -1138
rect 23444 -1274 23525 -1164
rect 32505 -1202 32517 -1150
rect 32569 -1202 32581 -1150
rect 32505 -1214 32581 -1202
rect 23444 -1326 23454 -1274
rect 23506 -1326 23525 -1274
rect 23444 -1412 23525 -1326
rect 25533 -1355 25611 -1340
rect 25533 -1373 25546 -1355
rect 23444 -1464 23447 -1412
rect 23499 -1464 23525 -1412
rect 25505 -1407 25546 -1373
rect 25598 -1373 25611 -1355
rect 25692 -1354 25770 -1339
rect 25692 -1373 25705 -1354
rect 25598 -1406 25705 -1373
rect 25757 -1373 25770 -1354
rect 31554 -1347 31694 -1284
rect 32518 -1311 32567 -1214
rect 32510 -1323 32586 -1311
rect 25757 -1406 25869 -1373
rect 25598 -1407 25869 -1406
rect 25505 -1419 25869 -1407
rect 25533 -1422 25611 -1419
rect 25692 -1421 25770 -1419
rect 23444 -1483 23525 -1464
rect 23444 -1564 23798 -1483
rect 18190 -2877 18204 -2871
rect 18125 -2890 18204 -2877
rect 23111 -2873 23379 -2827
rect 7280 -2971 7359 -2957
rect 7280 -3023 7292 -2971
rect 7344 -3023 7359 -2971
rect 7280 -3035 7359 -3023
rect 492 -3274 558 -3272
rect 487 -3288 566 -3274
rect 487 -3340 499 -3288
rect 551 -3340 566 -3288
rect 11137 -3296 11203 -3257
rect 11118 -3310 11203 -3296
rect 487 -3352 566 -3340
rect 2712 -3334 2795 -3320
rect 492 -3483 558 -3352
rect 2712 -3386 2728 -3334
rect 2780 -3386 2795 -3334
rect 2712 -3400 2795 -3386
rect 6215 -3329 6290 -3315
rect 6215 -3381 6227 -3329
rect 6279 -3381 6290 -3329
rect 6215 -3394 6290 -3381
rect 7264 -3331 7343 -3317
rect 7264 -3383 7276 -3331
rect 7328 -3383 7343 -3331
rect 2722 -3475 2768 -3400
rect 483 -3497 562 -3483
rect 483 -3549 495 -3497
rect 547 -3549 562 -3497
rect 483 -3561 562 -3549
rect 2706 -3489 2789 -3475
rect 6233 -3488 6279 -3394
rect 7264 -3395 7343 -3383
rect 9700 -3358 9777 -3346
rect 9700 -3410 9712 -3358
rect 9764 -3410 9777 -3358
rect 11118 -3362 11130 -3310
rect 11182 -3362 11203 -3310
rect 11118 -3374 11203 -3362
rect 13352 -3304 13431 -3290
rect 13352 -3356 13364 -3304
rect 13416 -3356 13431 -3304
rect 13352 -3368 13431 -3356
rect 9700 -3422 9777 -3410
rect 2706 -3541 2722 -3489
rect 2774 -3541 2789 -3489
rect 2706 -3555 2789 -3541
rect 6218 -3502 6293 -3488
rect 6218 -3554 6230 -3502
rect 6282 -3554 6293 -3502
rect 9709 -3513 9755 -3422
rect 492 -3627 558 -3561
rect 395 -3693 558 -3627
rect 2722 -3683 2768 -3555
rect 6218 -3567 6293 -3554
rect 9699 -3525 9776 -3513
rect 6233 -3683 6279 -3567
rect 9699 -3577 9711 -3525
rect 9763 -3577 9776 -3525
rect 9699 -3589 9776 -3577
rect 9709 -3683 9755 -3589
rect 10930 -3627 10996 -3590
rect 11137 -3627 11203 -3374
rect 13357 -3451 13403 -3368
rect 13348 -3465 13427 -3451
rect 13348 -3517 13360 -3465
rect 13412 -3517 13427 -3465
rect 13348 -3529 13427 -3517
rect 10930 -3693 11203 -3627
rect 13357 -3683 13403 -3529
rect 5554 -4202 5648 -4184
rect 5554 -4254 5578 -4202
rect 5630 -4254 5648 -4202
rect 5554 -4267 5648 -4254
rect 15441 -4188 15541 -4171
rect 15441 -4240 15466 -4188
rect 15518 -4240 15541 -4188
rect 15441 -4262 15541 -4240
rect 23111 -4352 23157 -2873
rect 31024 -3181 31070 -1872
rect 31554 -2007 31617 -1347
rect 32510 -1375 32522 -1323
rect 32574 -1375 32586 -1323
rect 39210 -1326 39562 10145
rect 32510 -1387 32586 -1375
rect 32518 -1421 32567 -1387
rect 35219 -1678 39562 -1326
rect 32220 -1895 32411 -1798
rect 31549 -2019 31625 -2007
rect 31549 -2071 31561 -2019
rect 31613 -2071 31625 -2019
rect 31549 -2083 31625 -2071
rect 31554 -2220 31617 -2083
rect 31540 -2232 31617 -2220
rect 31540 -2284 31552 -2232
rect 31604 -2284 31617 -2232
rect 31540 -2296 31617 -2284
rect 31554 -2415 31617 -2296
rect 31536 -2427 31617 -2415
rect 31536 -2479 31548 -2427
rect 31600 -2479 31617 -2427
rect 31536 -2491 31617 -2479
rect 31554 -2502 31617 -2491
rect 32488 -2476 32564 -2464
rect 32488 -2502 32500 -2476
rect 32390 -2528 32500 -2502
rect 32552 -2502 32564 -2476
rect 32552 -2528 32656 -2502
rect 32390 -2551 32656 -2528
rect 32636 -2686 32717 -2670
rect 32636 -2738 32650 -2686
rect 32702 -2738 32717 -2686
rect 32636 -2755 32717 -2738
rect 32881 -2685 32962 -2669
rect 32881 -2737 32895 -2685
rect 32947 -2737 32962 -2685
rect 32881 -2754 32962 -2737
rect 34968 -2887 35059 -2412
rect 40117 -2887 40132 11232
rect 32198 -2947 32274 -2935
rect 32198 -2999 32210 -2947
rect 32262 -2999 32274 -2947
rect 32198 -3011 32274 -2999
rect 32212 -3107 32258 -3011
rect 34940 -3033 40132 -2887
rect 765 -4368 844 -4354
rect 765 -4370 777 -4368
rect 90 -4420 777 -4370
rect 829 -4370 844 -4368
rect 964 -4369 1043 -4355
rect 964 -4370 976 -4369
rect 829 -4420 976 -4370
rect 90 -4421 976 -4420
rect 1028 -4421 1043 -4369
rect 90 -4426 1043 -4421
rect 90 -4790 146 -4426
rect 765 -4432 844 -4426
rect 964 -4433 1043 -4426
rect 19378 -4398 23157 -4352
rect 23291 -3227 31070 -3181
rect 32198 -3119 32274 -3107
rect 32198 -3171 32210 -3119
rect 32262 -3171 32274 -3119
rect 32198 -3183 32274 -3171
rect 3278 -4529 3357 -4515
rect 3278 -4581 3290 -4529
rect 3342 -4581 3357 -4529
rect 3278 -4593 3357 -4581
rect 3612 -4523 3691 -4509
rect 3612 -4575 3624 -4523
rect 3676 -4575 3691 -4523
rect 3612 -4587 3691 -4575
rect 9562 -4542 9640 -4530
rect 9562 -4594 9574 -4542
rect 9626 -4594 9640 -4542
rect 9562 -4606 9640 -4594
rect 9799 -4533 9877 -4521
rect 9799 -4585 9811 -4533
rect 9863 -4585 9877 -4533
rect 9799 -4597 9877 -4585
rect 10397 -4542 10475 -4530
rect 10397 -4594 10409 -4542
rect 10461 -4594 10475 -4542
rect 10397 -4606 10475 -4594
rect 10644 -4542 10722 -4530
rect 10644 -4594 10656 -4542
rect 10708 -4594 10722 -4542
rect 10644 -4606 10722 -4594
rect 305 -4672 384 -4658
rect 305 -4724 317 -4672
rect 369 -4724 384 -4672
rect 305 -4736 384 -4724
rect 9565 -4708 9643 -4696
rect 9565 -4760 9577 -4708
rect 9629 -4760 9643 -4708
rect 9565 -4772 9643 -4760
rect 9813 -4706 9891 -4694
rect 9813 -4758 9825 -4706
rect 9877 -4758 9891 -4706
rect 9813 -4770 9891 -4758
rect 10407 -4695 10485 -4683
rect 10407 -4747 10419 -4695
rect 10471 -4747 10485 -4695
rect 10407 -4759 10485 -4747
rect 10656 -4691 10734 -4679
rect 10656 -4743 10668 -4691
rect 10720 -4743 10734 -4691
rect 10656 -4755 10734 -4743
rect -87 -4846 146 -4790
rect 303 -4829 382 -4815
rect -87 -5207 -31 -4846
rect 303 -4881 315 -4829
rect 367 -4881 382 -4829
rect 303 -4893 382 -4881
rect 2361 -4839 2440 -4825
rect 2361 -4891 2373 -4839
rect 2425 -4891 2440 -4839
rect 2361 -4903 2440 -4891
rect 2603 -4837 2682 -4823
rect 2603 -4889 2615 -4837
rect 2667 -4889 2682 -4837
rect 19378 -4852 19424 -4398
rect 19576 -4852 19622 -4398
rect 23291 -4763 23337 -3227
rect 23145 -4809 23337 -4763
rect 2603 -4901 2682 -4889
rect 21019 -4928 21098 -4914
rect 21019 -4980 21031 -4928
rect 21083 -4980 21098 -4928
rect 21019 -4992 21098 -4980
rect 21312 -4922 21391 -4908
rect 21312 -4974 21324 -4922
rect 21376 -4974 21391 -4922
rect 21312 -4986 21391 -4974
rect 21894 -4957 21973 -4943
rect 21894 -5009 21906 -4957
rect 21958 -5009 21973 -4957
rect 21894 -5021 21973 -5009
rect 22063 -4949 22142 -4935
rect 22063 -5001 22075 -4949
rect 22127 -5001 22142 -4949
rect 22063 -5013 22142 -5001
rect -88 -5221 -9 -5207
rect -88 -5273 -76 -5221
rect -24 -5273 -9 -5221
rect -88 -5285 -9 -5273
rect -87 -5386 -31 -5285
rect -96 -5400 -17 -5386
rect -96 -5452 -84 -5400
rect -32 -5452 -17 -5400
rect -96 -5464 -17 -5452
rect -87 -5465 -31 -5464
rect 3693 -5465 3759 -5336
rect 22733 -5455 22910 -5409
rect 3677 -5479 3759 -5465
rect 3677 -5531 3689 -5479
rect 3741 -5531 3759 -5479
rect 3677 -5543 3759 -5531
rect 317 -5753 379 -5751
rect 317 -5805 322 -5753
rect 374 -5805 379 -5753
rect 317 -5806 379 -5805
rect 2751 -5822 2797 -5714
rect 2750 -5836 2829 -5822
rect 2750 -5888 2762 -5836
rect 2814 -5888 2829 -5836
rect 2750 -5900 2829 -5888
rect 317 -5940 379 -5938
rect 317 -5992 322 -5940
rect 374 -5992 379 -5940
rect 317 -5993 379 -5992
rect 2751 -5995 2797 -5900
rect 3693 -5921 3759 -5543
rect 6265 -5810 6311 -5714
rect 6241 -5824 6320 -5810
rect 6241 -5876 6253 -5824
rect 6305 -5876 6320 -5824
rect 6241 -5888 6320 -5876
rect 7424 -5844 7503 -5830
rect 9829 -5841 9875 -5714
rect 3693 -5987 3876 -5921
rect 6265 -5986 6311 -5888
rect 7424 -5896 7436 -5844
rect 7488 -5896 7503 -5844
rect 7424 -5908 7503 -5896
rect 9815 -5855 9894 -5841
rect 9815 -5907 9827 -5855
rect 9879 -5907 9894 -5855
rect 9815 -5919 9894 -5907
rect 2748 -6009 2827 -5995
rect 2748 -6061 2760 -6009
rect 2812 -6061 2827 -6009
rect 2748 -6073 2827 -6061
rect 6239 -6000 6318 -5986
rect 6239 -6052 6251 -6000
rect 6303 -6052 6318 -6000
rect 9829 -6022 9875 -5919
rect 9814 -6036 9893 -6022
rect 6239 -6064 6318 -6052
rect 7415 -6061 7494 -6047
rect 2751 -6083 2797 -6073
rect 6265 -6077 6311 -6064
rect 7415 -6113 7427 -6061
rect 7479 -6113 7494 -6061
rect 9814 -6088 9826 -6036
rect 9878 -6088 9893 -6036
rect 9814 -6100 9893 -6088
rect 7415 -6125 7494 -6113
rect 22864 -6464 22910 -5455
rect 23145 -5545 23191 -4809
rect 23369 -4954 23448 -4940
rect 23369 -5006 23381 -4954
rect 23433 -5006 23448 -4954
rect 23369 -5018 23448 -5006
rect 23591 -4946 23670 -4932
rect 23591 -4998 23603 -4946
rect 23655 -4998 23670 -4946
rect 23591 -5010 23670 -4998
rect 24094 -4948 24147 -4946
rect 24146 -5000 24147 -4948
rect 24094 -5002 24147 -5000
rect 24267 -4948 24320 -4946
rect 24319 -5000 24320 -4948
rect 24267 -5002 24320 -5000
rect 24846 -5126 24892 -4975
rect 23145 -5591 23381 -5545
rect 24672 -5981 24719 -5499
rect 32212 -5530 32258 -3183
rect 24347 -6028 24719 -5981
rect 24781 -6066 25023 -5985
rect 26706 -5997 26785 -5983
rect 26706 -6049 26718 -5997
rect 26770 -6049 26785 -5997
rect 26706 -6061 26785 -6049
rect 27047 -5999 27126 -5985
rect 27047 -6051 27059 -5999
rect 27111 -6051 27126 -5999
rect 27047 -6063 27126 -6051
rect 31675 -5998 31756 -5982
rect 31675 -6050 31689 -5998
rect 31741 -6050 31756 -5998
rect 22864 -6510 23472 -6464
rect 24781 -6904 24862 -6066
rect 31675 -6067 31756 -6050
rect 31774 -5994 31936 -5978
rect 31774 -6046 31869 -5994
rect 31921 -6046 31936 -5994
rect 31774 -6059 31936 -6046
rect 31855 -6063 31936 -6059
rect 917 -6937 6408 -6922
rect 917 -6989 929 -6937
rect 981 -6940 6408 -6937
rect 981 -6984 1148 -6940
rect 981 -6989 996 -6984
rect 917 -7001 996 -6989
rect 1136 -6992 1148 -6984
rect 1200 -6984 6408 -6940
rect 1200 -6992 1215 -6984
rect 1136 -7004 1215 -6992
rect 6345 -7042 6408 -6984
rect 23326 -6928 23404 -6920
rect 24162 -6928 24862 -6904
rect 23326 -6985 24862 -6928
rect 6340 -7044 6417 -7042
rect 6686 -7044 6763 -7041
rect 6340 -7053 6763 -7044
rect 7125 -7045 7202 -7039
rect 7277 -7045 7354 -7039
rect 6340 -7054 6698 -7053
rect 6340 -7106 6352 -7054
rect 6404 -7057 6698 -7054
rect 6404 -7106 6513 -7057
rect 6340 -7109 6513 -7106
rect 6565 -7105 6698 -7057
rect 6750 -7105 6763 -7053
rect 6565 -7109 6763 -7105
rect 6340 -7111 6763 -7109
rect 7119 -7051 7354 -7045
rect 7119 -7103 7137 -7051
rect 7189 -7103 7289 -7051
rect 7341 -7103 7354 -7051
rect 7119 -7111 7354 -7103
rect 6340 -7118 6417 -7111
rect 6501 -7121 6578 -7111
rect 6686 -7117 6763 -7111
rect 7125 -7115 7202 -7111
rect 7277 -7115 7354 -7111
rect 23326 -7097 24219 -6985
rect 7279 -7544 7345 -7115
rect 11418 -7216 11478 -7197
rect 11378 -7242 11497 -7216
rect 11378 -7294 11420 -7242
rect 11472 -7294 11497 -7242
rect 11378 -7324 11497 -7294
rect 11418 -7348 11478 -7324
rect 23326 -7577 23506 -7097
rect 23102 -7590 23506 -7577
rect 20359 -7621 23506 -7590
rect 18682 -7699 23506 -7621
rect 20359 -7746 23506 -7699
rect 3773 -7763 3852 -7749
rect 20359 -7759 23271 -7746
rect 3773 -7815 3785 -7763
rect 3837 -7815 3852 -7763
rect 3773 -7827 3852 -7815
rect 6211 -7781 6291 -7767
rect 6211 -7833 6222 -7781
rect 6274 -7833 6291 -7781
rect 3768 -7945 3847 -7931
rect 3768 -7997 3780 -7945
rect 3832 -7997 3847 -7945
rect 6211 -7932 6291 -7833
rect 9689 -7783 9768 -7769
rect 9689 -7835 9701 -7783
rect 9753 -7835 9768 -7783
rect 9689 -7847 9768 -7835
rect 10932 -7785 11011 -7771
rect 10932 -7837 10944 -7785
rect 10996 -7837 11011 -7785
rect 6211 -7984 6225 -7932
rect 6277 -7984 6291 -7932
rect 9700 -7934 9746 -7847
rect 10932 -7849 11011 -7837
rect 13387 -7808 13466 -7794
rect 13387 -7860 13399 -7808
rect 13451 -7860 13466 -7808
rect 13387 -7872 13466 -7860
rect 6211 -7996 6291 -7984
rect 9693 -7948 9772 -7934
rect 3768 -8009 3847 -7997
rect 307 -8116 386 -8102
rect 307 -8168 319 -8116
rect 371 -8168 386 -8116
rect 307 -8180 386 -8168
rect 490 -8115 569 -8101
rect 490 -8167 502 -8115
rect 554 -8167 569 -8115
rect 490 -8179 569 -8167
rect 6222 -8135 6269 -7996
rect 9693 -8000 9705 -7948
rect 9757 -8000 9772 -7948
rect 9693 -8012 9772 -8000
rect 10930 -8003 11009 -7989
rect 6222 -8181 6337 -8135
rect 9700 -8181 9746 -8012
rect 10930 -8055 10942 -8003
rect 10994 -8055 11009 -8003
rect 13394 -8009 13440 -7872
rect 17898 -7947 17945 -7946
rect 17869 -7969 17945 -7947
rect 10930 -8067 11009 -8055
rect 13385 -8023 13464 -8009
rect 13385 -8075 13397 -8023
rect 13449 -8075 13464 -8023
rect 13385 -8087 13464 -8075
rect 17869 -8021 17877 -7969
rect 17929 -8021 17945 -7969
rect 17869 -8038 17945 -8021
rect 13394 -8135 13440 -8087
rect 13293 -8181 13440 -8135
rect 17869 -8115 17916 -8038
rect 17869 -8128 17967 -8115
rect 17869 -8180 17897 -8128
rect 17949 -8134 17967 -8128
rect 17949 -8135 18040 -8134
rect 17949 -8136 18113 -8135
rect 17949 -8180 18109 -8136
rect 17869 -8181 18109 -8180
rect 17882 -8193 17967 -8181
rect 634 -8918 713 -8914
rect 911 -8918 990 -8913
rect -210 -8927 990 -8918
rect -210 -8928 923 -8927
rect -210 -8980 646 -8928
rect 698 -8979 923 -8928
rect 975 -8979 990 -8927
rect 698 -8980 990 -8979
rect -210 -8981 990 -8980
rect 634 -8992 713 -8981
rect 911 -8991 990 -8981
rect 20360 -9233 20484 -7759
rect 21050 -9233 21174 -7759
rect -441 -9288 -341 -9246
rect 1480 -9248 2100 -9240
rect 1480 -9254 2012 -9248
rect 1480 -9257 1861 -9254
rect 1480 -9259 1734 -9257
rect 1480 -9264 1617 -9259
rect 1480 -9288 1502 -9264
rect -441 -9304 1502 -9288
rect 1554 -9304 1617 -9264
rect 1669 -9304 1734 -9259
rect 1786 -9304 1861 -9257
rect 1913 -9300 2012 -9254
rect 2064 -9288 2100 -9248
rect 20360 -9288 21174 -9233
rect 21965 -9288 22134 -7759
rect 23102 -9288 23271 -7759
rect 24050 -9288 24219 -7097
rect 40117 -9212 40132 -3033
rect 40178 -9212 40218 11232
rect 40117 -9288 40218 -9212
rect 2064 -9300 40218 -9288
rect 1913 -9304 40218 -9300
rect -441 -9350 -426 -9304
rect -185 -9350 -36 -9304
rect 40054 -9350 40132 -9304
rect 40178 -9350 40218 -9304
rect -441 -9366 40218 -9350
rect 1480 -9382 2100 -9366
rect 1480 -9384 1629 -9382
rect 1480 -9436 1514 -9384
rect 1566 -9434 1629 -9384
rect 1681 -9384 2100 -9382
rect 1681 -9434 1772 -9384
rect 1566 -9436 1772 -9434
rect 1824 -9436 1902 -9384
rect 1954 -9386 2100 -9384
rect 1954 -9436 2026 -9386
rect 1480 -9438 2026 -9436
rect 2078 -9438 2100 -9386
rect 11125 -9418 11693 -9366
rect 11125 -9430 11694 -9418
rect 19339 -9421 19907 -9366
rect 24050 -9394 24219 -9366
rect 1480 -9460 2100 -9438
rect 11127 -9459 11694 -9430
rect 11127 -9465 11426 -9459
rect 11127 -9468 11284 -9465
rect 11127 -9520 11160 -9468
rect 11212 -9517 11284 -9468
rect 11336 -9511 11426 -9465
rect 11478 -9461 11694 -9459
rect 11478 -9511 11570 -9461
rect 11336 -9513 11570 -9511
rect 11622 -9513 11694 -9461
rect 11336 -9517 11694 -9513
rect 11212 -9520 11694 -9517
rect 11127 -9576 11694 -9520
rect 11127 -9578 11423 -9576
rect 11127 -9583 11283 -9578
rect 11127 -9635 11156 -9583
rect 11208 -9630 11283 -9583
rect 11335 -9628 11423 -9578
rect 11475 -9580 11694 -9576
rect 11475 -9628 11564 -9580
rect 11335 -9630 11564 -9628
rect 11208 -9632 11564 -9630
rect 11616 -9632 11694 -9580
rect 11208 -9635 11694 -9632
rect 11127 -9662 11694 -9635
rect 19340 -9452 19907 -9421
rect 19340 -9458 19639 -9452
rect 19340 -9461 19497 -9458
rect 19340 -9513 19373 -9461
rect 19425 -9510 19497 -9461
rect 19549 -9504 19639 -9458
rect 19691 -9454 19907 -9452
rect 19691 -9504 19783 -9454
rect 19549 -9506 19783 -9504
rect 19835 -9506 19907 -9454
rect 19549 -9510 19907 -9506
rect 19425 -9513 19907 -9510
rect 19340 -9569 19907 -9513
rect 19340 -9571 19636 -9569
rect 19340 -9576 19496 -9571
rect 19340 -9628 19369 -9576
rect 19421 -9623 19496 -9576
rect 19548 -9621 19636 -9571
rect 19688 -9573 19907 -9569
rect 19688 -9621 19777 -9573
rect 19548 -9623 19777 -9621
rect 19421 -9625 19777 -9623
rect 19829 -9625 19907 -9573
rect 19421 -9628 19907 -9625
rect 19340 -9655 19907 -9628
rect 26402 -9433 26969 -9366
rect 26402 -9439 26701 -9433
rect 26402 -9442 26559 -9439
rect 26402 -9494 26435 -9442
rect 26487 -9491 26559 -9442
rect 26611 -9485 26701 -9439
rect 26753 -9435 26969 -9433
rect 26753 -9485 26845 -9435
rect 26611 -9487 26845 -9485
rect 26897 -9487 26969 -9435
rect 26611 -9491 26969 -9487
rect 26487 -9494 26969 -9491
rect 26402 -9550 26969 -9494
rect 26402 -9552 26698 -9550
rect 26402 -9557 26558 -9552
rect 26402 -9609 26431 -9557
rect 26483 -9604 26558 -9557
rect 26610 -9602 26698 -9552
rect 26750 -9554 26969 -9550
rect 26750 -9602 26839 -9554
rect 26610 -9604 26839 -9602
rect 26483 -9606 26839 -9604
rect 26891 -9606 26969 -9554
rect 26483 -9609 26969 -9606
rect 26402 -9636 26969 -9609
rect 33207 -9431 33774 -9366
rect 33207 -9437 33506 -9431
rect 33207 -9440 33364 -9437
rect 33207 -9492 33240 -9440
rect 33292 -9489 33364 -9440
rect 33416 -9483 33506 -9437
rect 33558 -9433 33774 -9431
rect 33558 -9483 33650 -9433
rect 33416 -9485 33650 -9483
rect 33702 -9485 33774 -9433
rect 33416 -9489 33774 -9485
rect 33292 -9492 33774 -9489
rect 33207 -9548 33774 -9492
rect 33207 -9550 33503 -9548
rect 33207 -9555 33363 -9550
rect 33207 -9607 33236 -9555
rect 33288 -9602 33363 -9555
rect 33415 -9600 33503 -9550
rect 33555 -9552 33774 -9548
rect 33555 -9600 33644 -9552
rect 33415 -9602 33644 -9600
rect 33288 -9604 33644 -9602
rect 33696 -9604 33774 -9552
rect 33288 -9607 33774 -9604
rect 33207 -9634 33774 -9607
rect 22630 -9811 23196 -9806
rect 15099 -9841 15665 -9836
rect 15099 -9882 15666 -9841
rect 15099 -9888 15398 -9882
rect 15099 -9891 15256 -9888
rect 5213 -9923 5779 -9918
rect 5213 -9964 5780 -9923
rect 5213 -9970 5512 -9964
rect 5213 -9973 5370 -9970
rect 5213 -10025 5246 -9973
rect 5298 -10022 5370 -9973
rect 5422 -10016 5512 -9970
rect 5564 -9966 5780 -9964
rect 5564 -10016 5656 -9966
rect 5422 -10018 5656 -10016
rect 5708 -10018 5780 -9966
rect 5422 -10022 5780 -10018
rect 5298 -10025 5780 -10022
rect 5213 -10081 5780 -10025
rect 5213 -10083 5509 -10081
rect 5213 -10088 5369 -10083
rect 5213 -10140 5242 -10088
rect 5294 -10135 5369 -10088
rect 5421 -10133 5509 -10083
rect 5561 -10085 5780 -10081
rect 15099 -9943 15132 -9891
rect 15184 -9940 15256 -9891
rect 15308 -9934 15398 -9888
rect 15450 -9884 15666 -9882
rect 15450 -9934 15542 -9884
rect 15308 -9936 15542 -9934
rect 15594 -9936 15666 -9884
rect 15308 -9940 15666 -9936
rect 15184 -9943 15666 -9940
rect 15099 -9999 15666 -9943
rect 15099 -10001 15395 -9999
rect 15099 -10006 15255 -10001
rect 15099 -10058 15128 -10006
rect 15180 -10053 15255 -10006
rect 15307 -10051 15395 -10001
rect 15447 -10003 15666 -9999
rect 15447 -10051 15536 -10003
rect 15307 -10053 15536 -10051
rect 15180 -10055 15536 -10053
rect 15588 -10055 15666 -10003
rect 22630 -9852 23197 -9811
rect 22630 -9858 22929 -9852
rect 22630 -9861 22787 -9858
rect 22630 -9913 22663 -9861
rect 22715 -9910 22787 -9861
rect 22839 -9904 22929 -9858
rect 22981 -9854 23197 -9852
rect 22981 -9904 23073 -9854
rect 22839 -9906 23073 -9904
rect 23125 -9906 23197 -9854
rect 22839 -9910 23197 -9906
rect 22715 -9913 23197 -9910
rect 22630 -9969 23197 -9913
rect 22630 -9971 22926 -9969
rect 22630 -9976 22786 -9971
rect 22630 -10028 22659 -9976
rect 22711 -10023 22786 -9976
rect 22838 -10021 22926 -9971
rect 22978 -9973 23197 -9969
rect 22978 -10021 23067 -9973
rect 22838 -10023 23067 -10021
rect 22711 -10025 23067 -10023
rect 23119 -10025 23197 -9973
rect 22711 -10028 23197 -10025
rect 22630 -10055 23197 -10028
rect 15180 -10058 15666 -10055
rect 15099 -10085 15666 -10058
rect 5561 -10133 5650 -10085
rect 5421 -10135 5650 -10133
rect 5294 -10137 5650 -10135
rect 5702 -10137 5780 -10085
rect 5294 -10140 5780 -10137
rect 5213 -10167 5780 -10140
<< via1 >>
rect 22655 12020 22707 12072
rect 22779 12023 22831 12075
rect 22921 12029 22973 12081
rect 23065 12027 23117 12079
rect 4999 11904 5051 11956
rect 5123 11907 5175 11959
rect 5265 11913 5317 11965
rect 5409 11911 5461 11963
rect 4995 11789 5047 11841
rect 5122 11794 5174 11846
rect 5262 11796 5314 11848
rect 5403 11792 5455 11844
rect 15132 11894 15184 11946
rect 15256 11897 15308 11949
rect 15398 11903 15450 11955
rect 15542 11901 15594 11953
rect 22651 11905 22703 11957
rect 22778 11910 22830 11962
rect 22918 11912 22970 11964
rect 23059 11908 23111 11960
rect 15128 11779 15180 11831
rect 15255 11784 15307 11836
rect 15395 11786 15447 11838
rect 15536 11782 15588 11834
rect 11295 11683 11347 11735
rect 11419 11686 11471 11738
rect 11561 11692 11613 11744
rect 11705 11690 11757 11742
rect 1636 11570 1688 11622
rect 1760 11573 1812 11625
rect 1902 11579 1954 11631
rect 2046 11577 2098 11629
rect 11291 11568 11343 11620
rect 11418 11573 11470 11625
rect 11558 11575 11610 11627
rect 11699 11571 11751 11623
rect 1632 11455 1684 11507
rect 1759 11460 1811 11512
rect 1899 11462 1951 11514
rect 2040 11458 2092 11510
rect 19160 11647 19212 11699
rect 19284 11650 19336 11702
rect 19426 11656 19478 11708
rect 19570 11654 19622 11706
rect 19156 11532 19208 11584
rect 19283 11537 19335 11589
rect 19423 11539 19475 11591
rect 19564 11535 19616 11587
rect 26141 11629 26193 11681
rect 26265 11632 26317 11684
rect 26407 11638 26459 11690
rect 26551 11636 26603 11688
rect 26137 11514 26189 11566
rect 26264 11519 26316 11571
rect 26404 11521 26456 11573
rect 26545 11517 26597 11569
rect 33014 11701 33066 11753
rect 33138 11704 33190 11756
rect 33280 11710 33332 11762
rect 33424 11708 33476 11760
rect 33010 11586 33062 11638
rect 33137 11591 33189 11643
rect 33277 11593 33329 11645
rect 33418 11589 33470 11641
rect 619 10876 671 10928
rect 774 10876 826 10928
rect 5158 10518 5210 10570
rect 38985 10420 39037 10472
rect 39105 10420 39157 10472
rect 39225 10420 39277 10472
rect 38985 10300 39037 10352
rect 39105 10300 39157 10352
rect 39225 10300 39277 10352
rect 38985 10180 39037 10232
rect 39105 10180 39157 10232
rect 39225 10180 39277 10232
rect 1705 9521 1757 9573
rect 1078 8596 1130 8648
rect 19523 8752 19575 8804
rect 9850 8602 9902 8654
rect 10202 8490 10254 8542
rect 10342 8489 10394 8541
rect 10207 8378 10259 8430
rect 11532 8426 11584 8478
rect 1685 7947 1737 7999
rect 26570 8363 26622 8415
rect 10301 7794 10353 7846
rect 10471 7794 10523 7846
rect 11517 7845 11569 7897
rect 19471 7557 19523 7609
rect 7943 7087 7995 7139
rect 7950 6941 8002 6993
rect 15521 5682 15573 5734
rect 5153 5296 5205 5348
rect 30958 5312 31010 5364
rect 31146 5310 31198 5362
rect 6867 4162 6919 4214
rect 6867 3997 6919 4049
rect 19478 3560 19530 3612
rect 9851 3379 9903 3431
rect 11324 3172 11376 3224
rect 11545 3167 11597 3219
rect 11740 3177 11792 3229
rect 3085 2957 3137 3009
rect 3375 2958 3427 3010
rect 1741 2751 1793 2803
rect 11498 2665 11550 2717
rect 26467 2635 26519 2687
rect 11036 2264 11088 2316
rect 11041 2129 11093 2181
rect 28947 1836 28999 1888
rect 29230 1835 29282 1887
rect 15217 465 15269 517
rect 7663 338 7715 390
rect 7818 339 7870 391
rect 4512 61 4564 113
rect 534 -244 586 -192
rect 6037 -39 6089 13
rect 2368 -105 2420 -53
rect 2555 -168 2607 -116
rect 2979 -127 3031 -75
rect 3183 -129 3235 -77
rect 19492 -215 19544 -163
rect 530 -411 582 -359
rect 3928 -431 3980 -379
rect 4151 -427 4203 -375
rect 6045 -419 6097 -367
rect 328 -1400 380 -1348
rect 3824 -1261 3876 -1209
rect 6222 -1314 6274 -1262
rect 7427 -1257 7479 -1205
rect 22676 -1204 22728 -1152
rect 2735 -1494 2787 -1442
rect 6227 -1483 6279 -1431
rect 9847 -1285 9899 -1233
rect 22676 -1339 22728 -1287
rect 335 -1584 387 -1532
rect 3820 -1567 3872 -1515
rect 7419 -1507 7471 -1455
rect 21890 -1701 21942 -1649
rect 22331 -1702 22383 -1650
rect 1777 -2482 1829 -2430
rect 4356 -2439 4408 -2387
rect 5255 -2477 5307 -2425
rect 5484 -2477 5536 -2425
rect 3808 -2623 3860 -2571
rect 4068 -2625 4120 -2573
rect 6100 -2585 6152 -2533
rect 6276 -2582 6328 -2530
rect 6455 -2587 6507 -2535
rect 9707 -2594 9759 -2542
rect 9899 -2594 9951 -2542
rect 21785 -2714 21837 -2662
rect 21940 -2718 21992 -2666
rect 11605 -2850 11657 -2798
rect 23493 -189 23545 -137
rect 23494 -358 23546 -306
rect 30303 3813 30355 3865
rect 30221 3657 30273 3709
rect 31709 1954 31761 2006
rect 37133 1799 37185 1851
rect 37368 1801 37420 1853
rect 30481 -501 30533 -449
rect 30678 -494 30730 -442
rect 31774 -488 31826 -436
rect 31960 -486 32012 -434
rect 32569 79 32621 131
rect 32560 -132 32612 -80
rect 17880 -2877 17932 -2825
rect 18138 -2877 18190 -2825
rect 32517 -1202 32569 -1150
rect 23454 -1326 23506 -1274
rect 23447 -1464 23499 -1412
rect 25546 -1407 25598 -1355
rect 25705 -1406 25757 -1354
rect 7292 -3023 7344 -2971
rect 499 -3340 551 -3288
rect 2728 -3386 2780 -3334
rect 6227 -3381 6279 -3329
rect 7276 -3383 7328 -3331
rect 495 -3549 547 -3497
rect 9712 -3410 9764 -3358
rect 11130 -3362 11182 -3310
rect 13364 -3356 13416 -3304
rect 2722 -3541 2774 -3489
rect 6230 -3554 6282 -3502
rect 9711 -3577 9763 -3525
rect 13360 -3517 13412 -3465
rect 5578 -4254 5630 -4202
rect 15466 -4240 15518 -4188
rect 32522 -1375 32574 -1323
rect 31561 -2071 31613 -2019
rect 31552 -2284 31604 -2232
rect 31548 -2479 31600 -2427
rect 32500 -2528 32552 -2476
rect 32650 -2738 32702 -2686
rect 32895 -2737 32947 -2685
rect 32210 -2999 32262 -2947
rect 777 -4420 829 -4368
rect 976 -4421 1028 -4369
rect 32210 -3171 32262 -3119
rect 3290 -4581 3342 -4529
rect 3624 -4575 3676 -4523
rect 9574 -4594 9626 -4542
rect 9811 -4585 9863 -4533
rect 10409 -4594 10461 -4542
rect 10656 -4594 10708 -4542
rect 317 -4724 369 -4672
rect 9577 -4760 9629 -4708
rect 9825 -4758 9877 -4706
rect 10419 -4747 10471 -4695
rect 10668 -4743 10720 -4691
rect 315 -4881 367 -4829
rect 2373 -4891 2425 -4839
rect 2615 -4889 2667 -4837
rect 21031 -4980 21083 -4928
rect 21324 -4974 21376 -4922
rect 21906 -5009 21958 -4957
rect 22075 -5001 22127 -4949
rect -76 -5273 -24 -5221
rect -84 -5452 -32 -5400
rect 3689 -5531 3741 -5479
rect 322 -5805 374 -5753
rect 2762 -5888 2814 -5836
rect 322 -5992 374 -5940
rect 6253 -5876 6305 -5824
rect 7436 -5896 7488 -5844
rect 9827 -5907 9879 -5855
rect 2760 -6061 2812 -6009
rect 6251 -6052 6303 -6000
rect 7427 -6113 7479 -6061
rect 9826 -6088 9878 -6036
rect 23381 -5006 23433 -4954
rect 23603 -4998 23655 -4946
rect 24094 -5000 24146 -4948
rect 24267 -5000 24319 -4948
rect 26718 -6049 26770 -5997
rect 27059 -6051 27111 -5999
rect 31689 -6050 31741 -5998
rect 31869 -6046 31921 -5994
rect 929 -6989 981 -6937
rect 1148 -6992 1200 -6940
rect 6352 -7106 6404 -7054
rect 6513 -7109 6565 -7057
rect 6698 -7105 6750 -7053
rect 7137 -7103 7189 -7051
rect 7289 -7103 7341 -7051
rect 11420 -7294 11472 -7242
rect 3785 -7815 3837 -7763
rect 6222 -7833 6274 -7781
rect 3780 -7997 3832 -7945
rect 9701 -7835 9753 -7783
rect 10944 -7837 10996 -7785
rect 6225 -7984 6277 -7932
rect 13399 -7860 13451 -7808
rect 319 -8168 371 -8116
rect 502 -8167 554 -8115
rect 9705 -8000 9757 -7948
rect 10942 -8055 10994 -8003
rect 13397 -8075 13449 -8023
rect 17877 -8021 17929 -7969
rect 17897 -8180 17949 -8128
rect 646 -8980 698 -8928
rect 923 -8979 975 -8927
rect 1502 -9304 1554 -9264
rect 1617 -9304 1669 -9259
rect 1734 -9304 1786 -9257
rect 1861 -9304 1913 -9254
rect 2012 -9300 2064 -9248
rect 1502 -9316 1554 -9304
rect 1617 -9311 1669 -9304
rect 1734 -9309 1786 -9304
rect 1861 -9306 1913 -9304
rect 1514 -9436 1566 -9384
rect 1629 -9434 1681 -9382
rect 1772 -9436 1824 -9384
rect 1902 -9436 1954 -9384
rect 2026 -9438 2078 -9386
rect 11160 -9520 11212 -9468
rect 11284 -9517 11336 -9465
rect 11426 -9511 11478 -9459
rect 11570 -9513 11622 -9461
rect 11156 -9635 11208 -9583
rect 11283 -9630 11335 -9578
rect 11423 -9628 11475 -9576
rect 11564 -9632 11616 -9580
rect 19373 -9513 19425 -9461
rect 19497 -9510 19549 -9458
rect 19639 -9504 19691 -9452
rect 19783 -9506 19835 -9454
rect 19369 -9628 19421 -9576
rect 19496 -9623 19548 -9571
rect 19636 -9621 19688 -9569
rect 19777 -9625 19829 -9573
rect 26435 -9494 26487 -9442
rect 26559 -9491 26611 -9439
rect 26701 -9485 26753 -9433
rect 26845 -9487 26897 -9435
rect 26431 -9609 26483 -9557
rect 26558 -9604 26610 -9552
rect 26698 -9602 26750 -9550
rect 26839 -9606 26891 -9554
rect 33240 -9492 33292 -9440
rect 33364 -9489 33416 -9437
rect 33506 -9483 33558 -9431
rect 33650 -9485 33702 -9433
rect 33236 -9607 33288 -9555
rect 33363 -9602 33415 -9550
rect 33503 -9600 33555 -9548
rect 33644 -9604 33696 -9552
rect 5246 -10025 5298 -9973
rect 5370 -10022 5422 -9970
rect 5512 -10016 5564 -9964
rect 5656 -10018 5708 -9966
rect 5242 -10140 5294 -10088
rect 5369 -10135 5421 -10083
rect 5509 -10133 5561 -10081
rect 15132 -9943 15184 -9891
rect 15256 -9940 15308 -9888
rect 15398 -9934 15450 -9882
rect 15542 -9936 15594 -9884
rect 15128 -10058 15180 -10006
rect 15255 -10053 15307 -10001
rect 15395 -10051 15447 -9999
rect 15536 -10055 15588 -10003
rect 22663 -9913 22715 -9861
rect 22787 -9910 22839 -9858
rect 22929 -9904 22981 -9852
rect 23073 -9906 23125 -9854
rect 22659 -10028 22711 -9976
rect 22786 -10023 22838 -9971
rect 22926 -10021 22978 -9969
rect 23067 -10025 23119 -9973
rect 5650 -10137 5702 -10085
<< metal2 >>
rect 22623 12083 23189 12122
rect 22623 12077 22919 12083
rect 22975 12081 23189 12083
rect 22623 12074 22777 12077
rect 22623 12018 22653 12074
rect 22709 12021 22777 12074
rect 22833 12027 22919 12077
rect 22975 12027 23063 12081
rect 22833 12025 23063 12027
rect 23119 12025 23189 12081
rect 22833 12021 23189 12025
rect 22709 12018 23189 12021
rect 4967 11967 5533 12006
rect 4967 11961 5263 11967
rect 5319 11965 5533 11967
rect 4967 11958 5121 11961
rect 4967 11902 4997 11958
rect 5053 11905 5121 11958
rect 5177 11911 5263 11961
rect 5319 11911 5407 11965
rect 5177 11909 5407 11911
rect 5463 11909 5533 11965
rect 5177 11905 5533 11909
rect 5053 11902 5533 11905
rect 4967 11850 5533 11902
rect 4967 11848 5260 11850
rect 4967 11843 5120 11848
rect 4967 11787 4993 11843
rect 5049 11792 5120 11843
rect 5176 11794 5260 11848
rect 5316 11846 5533 11850
rect 5316 11794 5401 11846
rect 5176 11792 5401 11794
rect 5049 11790 5401 11792
rect 5457 11790 5533 11846
rect 5049 11787 5533 11790
rect 4967 11768 5533 11787
rect 15100 11957 15666 11996
rect 15100 11951 15396 11957
rect 15452 11955 15666 11957
rect 15100 11948 15254 11951
rect 15100 11892 15130 11948
rect 15186 11895 15254 11948
rect 15310 11901 15396 11951
rect 15452 11901 15540 11955
rect 15310 11899 15540 11901
rect 15596 11899 15666 11955
rect 15310 11895 15666 11899
rect 15186 11892 15666 11895
rect 15100 11840 15666 11892
rect 22623 11966 23189 12018
rect 22623 11964 22916 11966
rect 22623 11959 22776 11964
rect 22623 11903 22649 11959
rect 22705 11908 22776 11959
rect 22832 11910 22916 11964
rect 22972 11962 23189 11966
rect 22972 11910 23057 11962
rect 22832 11908 23057 11910
rect 22705 11906 23057 11908
rect 23113 11906 23189 11962
rect 22705 11903 23189 11906
rect 22623 11884 23189 11903
rect 15100 11838 15393 11840
rect 15100 11833 15253 11838
rect 11263 11746 11829 11785
rect 15100 11777 15126 11833
rect 15182 11782 15253 11833
rect 15309 11784 15393 11838
rect 15449 11836 15666 11840
rect 15449 11784 15534 11836
rect 15309 11782 15534 11784
rect 15182 11780 15534 11782
rect 15590 11780 15666 11836
rect 15182 11777 15666 11780
rect 15100 11758 15666 11777
rect 32982 11764 33548 11803
rect 32982 11758 33278 11764
rect 33334 11762 33548 11764
rect 32982 11755 33136 11758
rect 11263 11740 11559 11746
rect 11615 11744 11829 11746
rect 11263 11737 11417 11740
rect 11263 11681 11293 11737
rect 11349 11684 11417 11737
rect 11473 11690 11559 11740
rect 11615 11690 11703 11744
rect 11473 11688 11703 11690
rect 11759 11688 11829 11744
rect 11473 11684 11829 11688
rect 11349 11681 11829 11684
rect 1604 11633 2170 11672
rect 1604 11627 1900 11633
rect 1956 11631 2170 11633
rect 1604 11624 1758 11627
rect 1604 11568 1634 11624
rect 1690 11571 1758 11624
rect 1814 11577 1900 11627
rect 1956 11577 2044 11631
rect 1814 11575 2044 11577
rect 2100 11575 2170 11631
rect 1814 11571 2170 11575
rect 1690 11568 2170 11571
rect 1604 11516 2170 11568
rect 11263 11629 11829 11681
rect 11263 11627 11556 11629
rect 11263 11622 11416 11627
rect 11263 11566 11289 11622
rect 11345 11571 11416 11622
rect 11472 11573 11556 11627
rect 11612 11625 11829 11629
rect 11612 11573 11697 11625
rect 11472 11571 11697 11573
rect 11345 11569 11697 11571
rect 11753 11569 11829 11625
rect 11345 11566 11829 11569
rect 11263 11547 11829 11566
rect 19128 11710 19694 11749
rect 19128 11704 19424 11710
rect 19480 11708 19694 11710
rect 19128 11701 19282 11704
rect 19128 11645 19158 11701
rect 19214 11648 19282 11701
rect 19338 11654 19424 11704
rect 19480 11654 19568 11708
rect 19338 11652 19568 11654
rect 19624 11652 19694 11708
rect 19338 11648 19694 11652
rect 19214 11645 19694 11648
rect 19128 11593 19694 11645
rect 19128 11591 19421 11593
rect 19128 11586 19281 11591
rect 1604 11514 1897 11516
rect 1604 11509 1757 11514
rect 1604 11453 1630 11509
rect 1686 11458 1757 11509
rect 1813 11460 1897 11514
rect 1953 11512 2170 11516
rect 1953 11460 2038 11512
rect 1813 11458 2038 11460
rect 1686 11456 2038 11458
rect 2094 11456 2170 11512
rect 19128 11530 19154 11586
rect 19210 11535 19281 11586
rect 19337 11537 19421 11591
rect 19477 11589 19694 11593
rect 19477 11537 19562 11589
rect 19337 11535 19562 11537
rect 19210 11533 19562 11535
rect 19618 11533 19694 11589
rect 19210 11530 19694 11533
rect 19128 11511 19694 11530
rect 26109 11692 26675 11731
rect 26109 11686 26405 11692
rect 26461 11690 26675 11692
rect 26109 11683 26263 11686
rect 26109 11627 26139 11683
rect 26195 11630 26263 11683
rect 26319 11636 26405 11686
rect 26461 11636 26549 11690
rect 26319 11634 26549 11636
rect 26605 11634 26675 11690
rect 26319 11630 26675 11634
rect 26195 11627 26675 11630
rect 26109 11575 26675 11627
rect 26109 11573 26402 11575
rect 26109 11568 26262 11573
rect 26109 11512 26135 11568
rect 26191 11517 26262 11568
rect 26318 11519 26402 11573
rect 26458 11571 26675 11575
rect 26458 11519 26543 11571
rect 26318 11517 26543 11519
rect 26191 11515 26543 11517
rect 26599 11515 26675 11571
rect 32982 11699 33012 11755
rect 33068 11702 33136 11755
rect 33192 11708 33278 11758
rect 33334 11708 33422 11762
rect 33192 11706 33422 11708
rect 33478 11706 33548 11762
rect 33192 11702 33548 11706
rect 33068 11699 33548 11702
rect 32982 11647 33548 11699
rect 32982 11645 33275 11647
rect 32982 11640 33135 11645
rect 32982 11584 33008 11640
rect 33064 11589 33135 11640
rect 33191 11591 33275 11645
rect 33331 11643 33548 11647
rect 33331 11591 33416 11643
rect 33191 11589 33416 11591
rect 33064 11587 33416 11589
rect 33472 11587 33548 11643
rect 33064 11584 33548 11587
rect 32982 11565 33548 11584
rect 26191 11512 26675 11515
rect 26109 11493 26675 11512
rect 1686 11453 2170 11456
rect 1604 11434 2170 11453
rect 18237 11328 18580 11336
rect -134 11326 18580 11328
rect -134 11324 18463 11326
rect -134 11268 18247 11324
rect 18303 11270 18463 11324
rect 18519 11270 18580 11326
rect 18303 11268 18580 11270
rect -134 11265 18580 11268
rect -118 -4526 -55 11265
rect 18237 11258 18580 11265
rect 606 10932 840 10942
rect 521 10928 840 10932
rect 39067 10931 39437 11939
rect 39026 10929 39479 10931
rect 521 10876 619 10928
rect 671 10876 774 10928
rect 826 10876 840 10928
rect 521 10862 840 10876
rect 534 -180 594 10862
rect 5140 10572 5228 10587
rect 5140 10516 5156 10572
rect 5212 10516 5228 10572
rect 5140 10499 5228 10516
rect 38953 10472 39755 10929
rect 38953 10420 38985 10472
rect 39037 10420 39105 10472
rect 39157 10420 39225 10472
rect 39277 10420 39755 10472
rect 38953 10352 39755 10420
rect 38953 10300 38985 10352
rect 39037 10300 39105 10352
rect 39157 10300 39225 10352
rect 39277 10300 39755 10352
rect 38953 10232 39755 10300
rect 38953 10180 38985 10232
rect 39037 10180 39105 10232
rect 39157 10180 39225 10232
rect 39277 10180 39755 10232
rect 38953 10145 39755 10180
rect 1654 9598 1814 9622
rect 1651 9575 1814 9598
rect 1651 9541 1703 9575
rect 1654 9519 1703 9541
rect 1759 9519 1814 9575
rect 1654 9483 1814 9519
rect 1670 9481 1748 9483
rect 19481 8806 19600 8830
rect 1052 8777 1151 8805
rect 1052 8721 1075 8777
rect 1131 8721 1151 8777
rect 1052 8686 1151 8721
rect 1053 8650 1151 8686
rect 1053 8594 1076 8650
rect 1132 8594 1151 8650
rect 1053 8390 1151 8594
rect 9843 8774 9935 8792
rect 9843 8718 9867 8774
rect 9923 8718 9935 8774
rect 19481 8750 19521 8806
rect 19577 8750 19600 8806
rect 19481 8722 19600 8750
rect 9843 8657 9935 8718
rect 9843 8654 9857 8657
rect 9843 8602 9850 8654
rect 9843 8601 9857 8602
rect 9913 8601 9935 8657
rect 9843 8543 9935 8601
rect 10183 8544 10411 8563
rect 9843 8539 9923 8543
rect 9843 8476 9914 8539
rect 10183 8488 10200 8544
rect 10256 8543 10411 8544
rect 10256 8488 10340 8543
rect 10183 8487 10340 8488
rect 10396 8487 10411 8543
rect 10183 8432 10411 8487
rect 10183 8376 10205 8432
rect 10261 8376 10411 8432
rect 11490 8480 11609 8504
rect 11490 8424 11530 8480
rect 11586 8424 11609 8480
rect 11490 8396 11609 8424
rect 26519 8439 26679 8472
rect 26519 8417 26711 8439
rect 10183 8332 10411 8376
rect 26519 8361 26568 8417
rect 26624 8414 26711 8417
rect 26624 8361 26679 8414
rect 26519 8325 26679 8361
rect 21686 8225 22426 8239
rect 702 8156 1133 8212
rect 21686 8169 21698 8225
rect 21754 8224 22426 8225
rect 21754 8169 21835 8224
rect 21686 8168 21835 8169
rect 21891 8168 22426 8224
rect 702 6528 758 8156
rect 18180 8109 18439 8119
rect 18180 8108 18373 8109
rect 11721 8088 11961 8098
rect 11721 8086 11895 8088
rect 1634 8024 1794 8048
rect 1631 8001 1794 8024
rect 11721 8030 11731 8086
rect 11787 8032 11895 8086
rect 11951 8032 11961 8088
rect 18180 8052 18190 8108
rect 18246 8053 18373 8108
rect 18429 8053 18439 8109
rect 18246 8052 18439 8053
rect 18180 8041 18439 8052
rect 11787 8030 11961 8032
rect 11721 8020 11961 8030
rect 1631 7967 1683 8001
rect 1634 7945 1683 7967
rect 1739 7945 1794 8001
rect 19981 7997 20058 8166
rect 21686 8158 22426 8168
rect 30989 8164 31058 9096
rect 30989 8095 33264 8164
rect 30989 8090 31058 8095
rect 1634 7909 1794 7945
rect 1650 7907 1728 7909
rect 10271 7848 10607 7903
rect 10271 7792 10299 7848
rect 10355 7792 10469 7848
rect 10525 7792 10607 7848
rect 11475 7899 11594 7923
rect 19551 7920 20058 7997
rect 11475 7843 11515 7899
rect 11571 7843 11594 7899
rect 11475 7815 11594 7843
rect 10271 7741 10607 7792
rect 19429 7611 19548 7635
rect 19429 7555 19469 7611
rect 19525 7555 19548 7611
rect 19429 7527 19548 7555
rect 7931 7141 8009 7151
rect 7931 7085 7942 7141
rect 7998 7085 8009 7141
rect 7931 7075 8009 7085
rect 7938 6995 8016 7005
rect 7938 6939 7949 6995
rect 8005 6939 8016 6995
rect 7938 6929 8016 6939
rect 702 6472 939 6528
rect 702 6462 758 6472
rect 883 -70 939 6472
rect 18585 6088 18796 6136
rect 18585 6058 19583 6088
rect 18585 6056 18726 6058
rect 18585 6000 18603 6056
rect 18659 6002 18726 6056
rect 18782 6002 19583 6058
rect 18659 6000 19583 6002
rect 18585 5955 19583 6000
rect 18585 5949 18796 5955
rect 18585 5942 18725 5949
rect 18585 5886 18604 5942
rect 18660 5893 18725 5942
rect 18781 5893 18796 5949
rect 18660 5886 18796 5893
rect 18585 5865 18796 5886
rect 18588 5864 18795 5865
rect 15496 5736 15593 5762
rect 15496 5680 15519 5736
rect 15575 5680 15593 5736
rect 15496 5658 15593 5680
rect 5131 5350 5219 5364
rect 5131 5294 5151 5350
rect 5207 5294 5219 5350
rect 5131 5276 5219 5294
rect 19450 5070 19583 5955
rect 22892 5733 22976 5753
rect 22892 5677 22904 5733
rect 22960 5677 22976 5733
rect 22892 5669 22976 5677
rect 33195 5547 33264 8095
rect 19172 4937 19583 5070
rect 29871 5478 33264 5547
rect 6854 4214 6930 4229
rect 6854 4162 6867 4214
rect 6919 4162 6930 4214
rect 6854 4146 6930 4162
rect 6857 4064 6926 4146
rect 6854 4049 6930 4064
rect 6854 3997 6867 4049
rect 6919 3997 6930 4049
rect 6854 3981 6930 3997
rect 1295 3012 1513 3024
rect 1295 2956 1424 3012
rect 1480 2956 1513 3012
rect 1295 2933 1513 2956
rect 3073 3011 3151 3021
rect 3073 2955 3084 3011
rect 3140 2955 3151 3011
rect 3073 2945 3151 2955
rect 3363 3012 3441 3022
rect 3363 2956 3374 3012
rect 3430 2956 3441 3012
rect 3363 2946 3441 2956
rect 1295 2877 1306 2933
rect 1362 2877 1513 2933
rect 1295 2874 1513 2877
rect 1295 2818 1425 2874
rect 1481 2818 1513 2874
rect 1690 2828 1850 2852
rect 1295 2802 1513 2818
rect 1687 2805 1850 2828
rect 6857 2820 6926 3981
rect 9843 3435 9922 3467
rect 9843 3431 9855 3435
rect 9843 3379 9851 3431
rect 9911 3379 9922 3435
rect 9843 3322 9922 3379
rect 9843 3266 9854 3322
rect 9910 3266 9922 3322
rect 9843 3259 9922 3266
rect 19172 3357 19305 4937
rect 19436 3614 19555 3638
rect 19436 3558 19476 3614
rect 19532 3558 19555 3614
rect 19436 3530 19555 3558
rect 9843 3250 9927 3259
rect 11311 3226 11390 3237
rect 11311 3170 11322 3226
rect 11378 3170 11390 3226
rect 11311 3159 11390 3170
rect 11532 3221 11611 3232
rect 11532 3165 11543 3221
rect 11599 3165 11611 3221
rect 11532 3154 11611 3165
rect 11727 3231 11806 3242
rect 11727 3175 11738 3231
rect 11794 3175 11806 3231
rect 19172 3224 19684 3357
rect 11727 3164 11806 3175
rect 25807 3004 26304 3021
rect 25807 3000 26136 3004
rect 1687 2771 1739 2805
rect 1690 2749 1739 2771
rect 1795 2749 1850 2805
rect 1690 2713 1850 2749
rect 6604 2740 6926 2820
rect 10084 2881 10163 2892
rect 10084 2825 10095 2881
rect 10151 2825 10163 2881
rect 10084 2815 10163 2825
rect 10322 2882 10401 2893
rect 10322 2826 10333 2882
rect 10389 2826 10401 2882
rect 13618 2844 14533 2900
rect 10322 2816 10401 2826
rect 1706 2711 1784 2713
rect 6604 395 6678 2740
rect 11456 2719 11575 2743
rect 11456 2663 11496 2719
rect 11552 2663 11575 2719
rect 11456 2635 11575 2663
rect 11023 2318 11102 2329
rect 11023 2262 11034 2318
rect 11090 2262 11102 2318
rect 11023 2251 11102 2262
rect 11028 2183 11107 2194
rect 11028 2127 11039 2183
rect 11095 2127 11107 2183
rect 11028 2116 11107 2127
rect 6604 340 6682 395
rect 4498 314 6682 340
rect 7651 393 7730 404
rect 7651 337 7662 393
rect 7718 337 7730 393
rect 7651 326 7730 337
rect 7806 394 7885 405
rect 7806 338 7817 394
rect 7873 338 7885 394
rect 7806 327 7885 338
rect 4498 266 6678 314
rect 4499 136 4577 266
rect 11249 162 11328 163
rect 11483 162 11562 167
rect 4500 125 4577 136
rect 4673 156 11562 162
rect 4673 152 11494 156
rect 4500 115 4578 125
rect 4500 59 4511 115
rect 4567 59 4578 115
rect 4500 49 4578 59
rect 4673 96 11260 152
rect 11316 100 11494 152
rect 11550 100 11562 156
rect 13917 113 13996 124
rect 13917 104 13928 113
rect 11316 96 11562 100
rect 4673 90 11562 96
rect 4503 47 4577 49
rect 2356 -51 2434 -41
rect 2356 -70 2367 -51
rect 883 -107 2367 -70
rect 2423 -70 2434 -51
rect 2423 -104 2605 -70
rect 2967 -73 3045 -63
rect 2967 -78 2978 -73
rect 2423 -107 2621 -104
rect 883 -114 2621 -107
rect 883 -126 2554 -114
rect 2543 -170 2554 -126
rect 2610 -170 2621 -114
rect 2943 -129 2978 -78
rect 3034 -78 3045 -73
rect 3171 -75 3249 -65
rect 3171 -78 3182 -75
rect 3034 -129 3182 -78
rect 3238 -78 3249 -75
rect 4673 -78 4745 90
rect 11249 86 11328 90
rect 13914 57 13928 104
rect 13984 104 13996 113
rect 14127 114 14206 125
rect 14127 104 14138 114
rect 13984 58 14138 104
rect 14194 104 14206 114
rect 14477 104 14533 2844
rect 15733 2573 15789 2663
rect 15442 2517 15789 2573
rect 15199 519 15283 533
rect 15199 463 15215 519
rect 15271 463 15283 519
rect 15199 447 15283 463
rect 14194 58 14533 104
rect 13984 57 14533 58
rect 13914 48 14533 57
rect 13917 47 13996 48
rect 6025 16 6104 27
rect 6025 -40 6036 16
rect 6092 -40 6104 16
rect 6290 -31 6369 -20
rect 6484 -30 6563 -19
rect 6484 -31 6495 -30
rect 6025 -51 6104 -40
rect 2943 -131 3182 -129
rect 3238 -131 4745 -78
rect 6247 -87 6301 -31
rect 6357 -86 6495 -31
rect 6551 -31 6563 -30
rect 14670 -31 14749 -22
rect 14873 -31 14952 -26
rect 15442 -31 15498 2517
rect 22504 376 22583 387
rect 22504 374 22515 376
rect 22442 320 22515 374
rect 22571 374 22583 376
rect 22679 374 22758 385
rect 24907 374 24963 2996
rect 25807 2944 25831 3000
rect 25887 2944 25979 3000
rect 26035 2948 26136 3000
rect 26192 2948 26304 3004
rect 26035 2944 26304 2948
rect 25807 2929 26304 2944
rect 26416 2712 26576 2744
rect 25748 2689 26576 2712
rect 25748 2655 26465 2689
rect 25748 2448 25805 2655
rect 26416 2633 26465 2655
rect 26521 2633 26576 2689
rect 26416 2597 26576 2633
rect 28898 1906 29204 1923
rect 28898 1893 29306 1906
rect 28898 1888 28948 1893
rect 29004 1892 29306 1893
rect 28898 1836 28947 1888
rect 29004 1887 29231 1892
rect 29004 1837 29230 1887
rect 28999 1836 29230 1837
rect 29287 1836 29306 1892
rect 28898 1835 29230 1836
rect 29282 1835 29306 1836
rect 28898 1821 29306 1835
rect 29173 1819 29306 1821
rect 22571 320 22690 374
rect 22442 318 22690 320
rect 22746 318 24963 374
rect 22504 310 22583 318
rect 22679 308 22758 318
rect 6551 -33 15498 -31
rect 6551 -86 14681 -33
rect 6357 -87 14681 -86
rect 6290 -97 6369 -87
rect 6484 -96 6563 -87
rect 14670 -89 14681 -87
rect 14737 -37 15498 -33
rect 14737 -87 14884 -37
rect 14737 -89 14749 -87
rect 14670 -99 14749 -89
rect 14873 -93 14884 -87
rect 14940 -87 15498 -37
rect 22720 189 25159 245
rect 14940 -93 14952 -87
rect 14873 -103 14952 -93
rect 2943 -150 4745 -131
rect 2543 -180 2621 -170
rect 19480 -160 19559 -149
rect 522 -190 600 -180
rect 522 -246 533 -190
rect 589 -246 600 -190
rect 19480 -216 19491 -160
rect 19547 -216 19559 -160
rect 522 -256 600 -246
rect 1185 -229 1417 -218
rect 19480 -227 19559 -216
rect 534 -347 594 -256
rect 1185 -285 1196 -229
rect 1252 -230 1417 -229
rect 1252 -285 1348 -230
rect 1185 -286 1348 -285
rect 1404 -238 1417 -230
rect 1404 -286 10079 -238
rect 1185 -294 10079 -286
rect 22720 -294 22776 189
rect 23480 -136 23559 -125
rect 23480 -192 23490 -136
rect 23546 -192 23559 -136
rect 23480 -202 23559 -192
rect 25681 -285 25750 -284
rect 29871 -285 29940 5478
rect 30960 5371 31023 5378
rect 30927 5367 31023 5371
rect 30927 5364 31229 5367
rect 30927 5312 30958 5364
rect 31010 5362 31229 5364
rect 31010 5312 31146 5362
rect 30927 5310 31146 5312
rect 31198 5310 31229 5362
rect 30927 5304 31229 5310
rect 30204 3865 30469 3880
rect 30204 3813 30303 3865
rect 30355 3813 30469 3865
rect 30204 3804 30469 3813
rect 30204 3801 30369 3804
rect 30204 3721 30276 3801
rect 30204 3709 30287 3721
rect 30204 3657 30221 3709
rect 30273 3657 30287 3709
rect 30204 3645 30287 3657
rect 30204 -103 30276 3645
rect 30960 3468 31023 5304
rect 30755 3405 31023 3468
rect 30755 2886 30818 3405
rect 31692 2011 31786 2029
rect 31692 2006 31710 2011
rect 31692 1954 31709 2006
rect 31766 1955 31786 2011
rect 31761 1954 31786 1955
rect 31692 1941 31786 1954
rect 37119 1861 37200 1867
rect 37354 1861 37435 1869
rect 37119 1853 37696 1861
rect 37119 1851 37368 1853
rect 37119 1799 37133 1851
rect 37185 1801 37368 1851
rect 37420 1801 37696 1853
rect 37185 1799 37696 1801
rect 37119 1782 37696 1799
rect 37119 475 37198 1782
rect 35781 396 37198 475
rect 32557 131 32633 143
rect 32557 79 32569 131
rect 32621 79 32633 131
rect 32557 67 32633 79
rect 32559 -68 32625 67
rect 32548 -80 32625 -68
rect 30204 -175 31359 -103
rect 32548 -132 32560 -80
rect 32612 -132 32625 -80
rect 32548 -144 32625 -132
rect 1185 -298 1417 -294
rect 518 -357 596 -347
rect 10023 -350 22776 -294
rect 23481 -305 23560 -294
rect 518 -413 529 -357
rect 585 -368 596 -357
rect 3916 -368 3994 -367
rect 4139 -368 4217 -363
rect 585 -373 4217 -368
rect 585 -377 4150 -373
rect 585 -413 3927 -377
rect 518 -423 3927 -413
rect 534 -428 3927 -423
rect 3916 -433 3927 -428
rect 3983 -428 4150 -377
rect 3983 -433 3994 -428
rect 3916 -443 3994 -433
rect 4139 -429 4150 -428
rect 4206 -429 4217 -373
rect 4139 -439 4217 -429
rect 6033 -364 6112 -353
rect 6033 -420 6044 -364
rect 6100 -420 6112 -364
rect 23481 -361 23491 -305
rect 23547 -361 23560 -305
rect 25680 -354 29940 -285
rect 23481 -371 23560 -361
rect 6033 -431 6112 -420
rect 25681 -710 25750 -354
rect 30469 -446 30548 -435
rect 30469 -502 30480 -446
rect 30536 -502 30548 -446
rect 30469 -513 30548 -502
rect 30666 -439 30745 -428
rect 30666 -495 30677 -439
rect 30733 -495 30745 -439
rect 30666 -506 30745 -495
rect 25499 -779 25750 -710
rect 22671 -1141 22742 -1140
rect 22670 -1152 22742 -1141
rect 3812 -1206 3891 -1195
rect 3812 -1262 3823 -1206
rect 3879 -1262 3891 -1206
rect 7415 -1202 7494 -1191
rect 3812 -1273 3891 -1262
rect 6210 -1259 6289 -1248
rect 6210 -1315 6221 -1259
rect 6277 -1315 6289 -1259
rect 7415 -1258 7426 -1202
rect 7482 -1258 7494 -1202
rect 22670 -1204 22676 -1152
rect 22728 -1204 22742 -1152
rect 7415 -1269 7494 -1258
rect 9835 -1230 9914 -1219
rect 9835 -1286 9846 -1230
rect 9902 -1286 9914 -1230
rect 9835 -1297 9914 -1286
rect 22670 -1287 22742 -1204
rect 6210 -1326 6289 -1315
rect 316 -1345 395 -1334
rect 316 -1401 327 -1345
rect 383 -1401 395 -1345
rect 22670 -1339 22676 -1287
rect 22728 -1339 22742 -1287
rect 316 -1412 395 -1401
rect 2718 -1428 2798 -1350
rect 6215 -1428 6294 -1417
rect 2718 -1439 2802 -1428
rect 2718 -1495 2734 -1439
rect 2790 -1495 2802 -1439
rect 6215 -1484 6226 -1428
rect 6282 -1484 6294 -1428
rect 6215 -1495 6294 -1484
rect 7407 -1452 7486 -1441
rect 2718 -1506 2802 -1495
rect 323 -1529 402 -1518
rect 323 -1585 334 -1529
rect 390 -1585 402 -1529
rect 323 -1596 402 -1585
rect 2718 -1654 2798 -1506
rect 3808 -1512 3887 -1501
rect 3808 -1568 3819 -1512
rect 3875 -1568 3887 -1512
rect 7407 -1508 7418 -1452
rect 7474 -1508 7486 -1452
rect 7407 -1519 7486 -1508
rect 3808 -1579 3887 -1568
rect 14890 -1596 14969 -1585
rect 14890 -1652 14901 -1596
rect 14957 -1652 14969 -1596
rect 2718 -1734 2863 -1654
rect 14890 -1662 14969 -1652
rect 21862 -1648 22410 -1635
rect 1726 -2405 1886 -2381
rect 1721 -2428 1886 -2405
rect 1721 -2462 1775 -2428
rect 1726 -2484 1775 -2462
rect 1831 -2484 1886 -2428
rect 1726 -2520 1886 -2484
rect 1742 -2780 1820 -2520
rect 2783 -2879 2863 -1734
rect 14901 -1746 14958 -1662
rect 21862 -1704 21886 -1648
rect 21942 -1649 22410 -1648
rect 21942 -1704 22328 -1649
rect 21862 -1705 22328 -1704
rect 22384 -1705 22410 -1649
rect 21862 -1717 22410 -1705
rect 14889 -1757 14968 -1746
rect 14889 -1813 14900 -1757
rect 14956 -1813 14968 -1757
rect 14889 -1823 14968 -1813
rect 14901 -1835 14968 -1823
rect 14901 -1891 15050 -1835
rect 4356 -2375 4421 -2263
rect 4344 -2385 4422 -2375
rect 4344 -2441 4355 -2385
rect 4411 -2420 4422 -2385
rect 4411 -2425 5670 -2420
rect 4411 -2441 5255 -2425
rect 4344 -2451 5255 -2441
rect 4356 -2477 5255 -2451
rect 5307 -2477 5484 -2425
rect 5536 -2477 5670 -2425
rect 4356 -2485 5670 -2477
rect 6054 -2530 6534 -2527
rect 6054 -2533 6276 -2530
rect 3796 -2568 3875 -2557
rect 3796 -2624 3807 -2568
rect 3863 -2624 3875 -2568
rect 3796 -2635 3875 -2624
rect 4056 -2570 4135 -2559
rect 4056 -2626 4067 -2570
rect 4123 -2626 4135 -2570
rect 6054 -2585 6100 -2533
rect 6152 -2582 6276 -2533
rect 6328 -2535 6534 -2530
rect 6328 -2582 6455 -2535
rect 6152 -2585 6455 -2582
rect 6054 -2587 6455 -2585
rect 6507 -2587 6534 -2535
rect 6054 -2592 6534 -2587
rect 9695 -2535 9773 -2530
rect 9887 -2535 9965 -2530
rect 9695 -2540 9971 -2535
rect 4056 -2637 4135 -2626
rect 2783 -2959 3059 -2879
rect 2783 -2962 2863 -2959
rect 487 -3285 566 -3274
rect 487 -3341 498 -3285
rect 554 -3341 566 -3285
rect 2712 -3322 2795 -3320
rect 487 -3352 566 -3341
rect 2707 -3334 2795 -3322
rect 2707 -3386 2728 -3334
rect 2780 -3386 2795 -3334
rect 2707 -3400 2795 -3386
rect 2707 -3475 2779 -3400
rect 483 -3494 562 -3483
rect 483 -3550 494 -3494
rect 550 -3550 562 -3494
rect 483 -3561 562 -3550
rect 2706 -3489 2789 -3475
rect 2706 -3541 2722 -3489
rect 2774 -3541 2789 -3489
rect 2706 -3555 2789 -3541
rect 765 -4365 844 -4354
rect 765 -4421 776 -4365
rect 832 -4421 844 -4365
rect 765 -4432 844 -4421
rect 964 -4366 1043 -4355
rect 964 -4422 975 -4366
rect 1031 -4422 1043 -4366
rect 964 -4433 1043 -4422
rect 2707 -4526 2779 -3555
rect -118 -4598 2779 -4526
rect 2979 -4504 3059 -2959
rect 6222 -3315 6287 -2592
rect 9695 -2596 9706 -2540
rect 9762 -2596 9898 -2540
rect 9954 -2596 9971 -2540
rect 9695 -2598 9971 -2596
rect 9695 -2606 9773 -2598
rect 9887 -2606 9965 -2598
rect 7280 -2968 7359 -2957
rect 7280 -3024 7291 -2968
rect 7347 -3024 7359 -2968
rect 7280 -3035 7359 -3024
rect 6215 -3329 6290 -3315
rect 6215 -3381 6227 -3329
rect 6279 -3381 6290 -3329
rect 6215 -3394 6290 -3381
rect 7264 -3328 7343 -3317
rect 7264 -3384 7275 -3328
rect 7331 -3384 7343 -3328
rect 9708 -3346 9771 -2606
rect 14749 -2715 14828 -2706
rect 14994 -2708 15050 -1891
rect 14935 -2715 15050 -2708
rect 14749 -2717 15050 -2715
rect 11563 -2796 11682 -2772
rect 14749 -2773 14760 -2717
rect 14816 -2719 15050 -2717
rect 14816 -2771 14946 -2719
rect 14816 -2773 14828 -2771
rect 14749 -2783 14828 -2773
rect 14935 -2775 14946 -2771
rect 15002 -2771 15050 -2719
rect 21773 -2659 21852 -2648
rect 21773 -2715 21784 -2659
rect 21840 -2715 21852 -2659
rect 21773 -2726 21852 -2715
rect 21928 -2663 22007 -2652
rect 21928 -2719 21939 -2663
rect 21995 -2719 22007 -2663
rect 21928 -2730 22007 -2719
rect 15002 -2775 15014 -2771
rect 14935 -2785 15014 -2775
rect 11563 -2852 11603 -2796
rect 11659 -2852 11682 -2796
rect 11563 -2880 11682 -2852
rect 17867 -2824 17946 -2813
rect 17867 -2880 17877 -2824
rect 17933 -2880 17946 -2824
rect 17867 -2890 17946 -2880
rect 18125 -2824 18204 -2813
rect 18125 -2880 18135 -2824
rect 18191 -2880 18204 -2824
rect 18125 -2890 18204 -2880
rect 22670 -2959 22742 -1339
rect 22848 -1142 23515 -1068
rect 22848 -1450 22922 -1142
rect 22848 -1506 22858 -1450
rect 22914 -1506 22922 -1450
rect 22848 -1621 22922 -1506
rect 23441 -1274 23515 -1142
rect 23441 -1326 23454 -1274
rect 23506 -1326 23515 -1274
rect 23441 -1412 23515 -1326
rect 23441 -1464 23447 -1412
rect 23499 -1464 23515 -1412
rect 25499 -1340 25568 -779
rect 25499 -1355 25611 -1340
rect 25499 -1407 25546 -1355
rect 25598 -1359 25611 -1355
rect 25692 -1354 25770 -1339
rect 25692 -1359 25705 -1354
rect 25598 -1406 25705 -1359
rect 25757 -1359 25770 -1354
rect 25757 -1406 25825 -1359
rect 25598 -1407 25825 -1406
rect 25499 -1428 25825 -1407
rect 23441 -1562 23515 -1464
rect 22848 -1677 22855 -1621
rect 22911 -1677 22922 -1621
rect 22848 -1697 22922 -1677
rect 31287 -2959 31359 -175
rect 32559 -263 32625 -144
rect 32493 -329 32625 -263
rect 31762 -433 31841 -422
rect 31762 -489 31773 -433
rect 31829 -489 31841 -433
rect 31762 -500 31841 -489
rect 31948 -431 32027 -420
rect 31948 -487 31959 -431
rect 32015 -487 32027 -431
rect 31948 -498 32027 -487
rect 32493 -1138 32559 -329
rect 32493 -1150 32581 -1138
rect 32493 -1202 32517 -1150
rect 32569 -1202 32581 -1150
rect 32493 -1214 32581 -1202
rect 32493 -1311 32559 -1214
rect 32493 -1323 32586 -1311
rect 32493 -1375 32522 -1323
rect 32574 -1375 32586 -1323
rect 32493 -1387 32586 -1375
rect 32493 -1393 32559 -1387
rect 31542 -2007 31614 -1993
rect 31542 -2019 31625 -2007
rect 31542 -2071 31561 -2019
rect 31613 -2071 31625 -2019
rect 31542 -2083 31625 -2071
rect 31542 -2220 31614 -2083
rect 31540 -2232 31616 -2220
rect 31540 -2284 31552 -2232
rect 31604 -2284 31616 -2232
rect 31540 -2296 31616 -2284
rect 31542 -2415 31614 -2296
rect 31536 -2427 31614 -2415
rect 31536 -2479 31548 -2427
rect 31600 -2479 31614 -2427
rect 31536 -2491 31614 -2479
rect 22670 -3031 31359 -2959
rect 11118 -3307 11197 -3296
rect 6222 -3488 6287 -3394
rect 7264 -3395 7343 -3384
rect 9700 -3358 9777 -3346
rect 9700 -3410 9712 -3358
rect 9764 -3410 9777 -3358
rect 11118 -3363 11129 -3307
rect 11185 -3363 11197 -3307
rect 11118 -3374 11197 -3363
rect 13352 -3301 13431 -3290
rect 13352 -3357 13363 -3301
rect 13419 -3357 13431 -3301
rect 13352 -3368 13431 -3357
rect 9700 -3422 9777 -3410
rect 6218 -3502 6293 -3488
rect 6218 -3554 6230 -3502
rect 6282 -3554 6293 -3502
rect 9708 -3513 9771 -3422
rect 13348 -3462 13427 -3451
rect 6218 -3567 6293 -3554
rect 9699 -3525 9776 -3513
rect 6222 -3572 6287 -3567
rect 9699 -3577 9711 -3525
rect 9763 -3577 9776 -3525
rect 13348 -3518 13359 -3462
rect 13415 -3518 13427 -3462
rect 13348 -3529 13427 -3518
rect 9699 -3589 9776 -3577
rect 9708 -3603 9771 -3589
rect 5554 -4200 5648 -4184
rect 5554 -4256 5576 -4200
rect 5632 -4256 5648 -4200
rect 5554 -4267 5648 -4256
rect 15441 -4186 15541 -4171
rect 15441 -4242 15464 -4186
rect 15520 -4242 15541 -4186
rect 15441 -4262 15541 -4242
rect 2979 -4520 3724 -4504
rect 2979 -4526 3623 -4520
rect 2979 -4582 3289 -4526
rect 3345 -4576 3623 -4526
rect 3679 -4576 3724 -4520
rect 9799 -4530 9877 -4521
rect 3345 -4582 3724 -4576
rect 2979 -4584 3724 -4582
rect 9550 -4531 10722 -4530
rect 9550 -4540 9810 -4531
rect 3278 -4593 3357 -4584
rect 3612 -4587 3691 -4584
rect 305 -4667 384 -4658
rect 305 -4669 387 -4667
rect 305 -4725 316 -4669
rect 372 -4725 387 -4669
rect 305 -4736 387 -4725
rect 311 -4815 387 -4736
rect 2707 -4672 2779 -4598
rect 9550 -4596 9573 -4540
rect 9629 -4587 9810 -4540
rect 9866 -4540 10722 -4531
rect 9866 -4587 10408 -4540
rect 9629 -4596 10408 -4587
rect 10464 -4596 10655 -4540
rect 10711 -4596 10722 -4540
rect 31542 -4583 31614 -2491
rect 32488 -2476 32564 -2464
rect 32488 -2506 32500 -2476
rect 32207 -2528 32500 -2506
rect 32552 -2506 32564 -2476
rect 32552 -2528 32612 -2506
rect 32207 -2563 32612 -2528
rect 32207 -2892 32264 -2563
rect 32636 -2684 32717 -2670
rect 32881 -2684 32962 -2669
rect 35781 -2684 35860 396
rect 32392 -2685 35860 -2684
rect 32392 -2686 32895 -2685
rect 32392 -2738 32650 -2686
rect 32702 -2737 32895 -2686
rect 32947 -2737 35860 -2685
rect 32702 -2738 35860 -2737
rect 32392 -2763 35860 -2738
rect 32207 -2935 32265 -2892
rect 32198 -2947 32274 -2935
rect 32198 -2999 32210 -2947
rect 32262 -2999 32274 -2947
rect 32198 -3011 32274 -2999
rect 32207 -3107 32265 -3011
rect 32198 -3119 32274 -3107
rect 32198 -3171 32210 -3119
rect 32262 -3171 32274 -3119
rect 32198 -3183 32274 -3171
rect 9550 -4603 10722 -4596
rect 9562 -4606 9640 -4603
rect 10397 -4606 10475 -4603
rect 10644 -4606 10722 -4603
rect 15336 -4655 31614 -4583
rect 2707 -4744 8089 -4672
rect 10407 -4687 10485 -4683
rect 10656 -4687 10734 -4679
rect 303 -4826 387 -4815
rect 303 -4882 314 -4826
rect 370 -4882 387 -4826
rect 2361 -4836 2440 -4825
rect 2361 -4839 2372 -4836
rect 2428 -4839 2440 -4836
rect 2603 -4834 2682 -4823
rect 2603 -4839 2614 -4834
rect 303 -4893 387 -4882
rect -88 -5218 -9 -5207
rect -88 -5274 -77 -5218
rect -21 -5274 -9 -5218
rect -88 -5285 -9 -5274
rect -96 -5397 -17 -5386
rect -96 -5453 -85 -5397
rect -29 -5453 -17 -5397
rect -96 -5464 -17 -5453
rect 311 -5753 387 -4893
rect 311 -5805 322 -5753
rect 374 -5805 387 -5753
rect 311 -5940 387 -5805
rect 311 -5992 322 -5940
rect 374 -5992 387 -5940
rect 311 -6012 387 -5992
rect 460 -4892 2372 -4839
rect 2428 -4890 2614 -4839
rect 2670 -4890 2682 -4834
rect 2428 -4892 2682 -4890
rect 460 -4901 2682 -4892
rect 8017 -4855 8089 -4744
rect 9540 -4689 10762 -4687
rect 9540 -4693 10667 -4689
rect 9540 -4704 10418 -4693
rect 9540 -4706 9824 -4704
rect 9540 -4762 9576 -4706
rect 9632 -4760 9824 -4706
rect 9880 -4749 10418 -4704
rect 10474 -4745 10667 -4693
rect 10723 -4745 10762 -4689
rect 10474 -4749 10762 -4745
rect 9880 -4760 10762 -4749
rect 9632 -4762 10762 -4760
rect 9540 -4771 10762 -4762
rect 15336 -4768 15408 -4655
rect 9565 -4772 9643 -4771
rect 11251 -4840 15408 -4768
rect 11251 -4855 11323 -4840
rect 460 -4904 2679 -4901
rect 460 -6069 525 -4904
rect 8017 -4927 11323 -4855
rect 21019 -4925 21098 -4914
rect 21019 -4981 21030 -4925
rect 21086 -4981 21098 -4925
rect 21019 -4992 21098 -4981
rect 21312 -4919 21391 -4908
rect 21312 -4975 21323 -4919
rect 21379 -4975 21391 -4919
rect 21312 -4986 21391 -4975
rect 21894 -4954 21973 -4943
rect 21894 -5010 21905 -4954
rect 21961 -5010 21973 -4954
rect 21894 -5021 21973 -5010
rect 22063 -4946 22142 -4935
rect 22063 -5002 22074 -4946
rect 22130 -5002 22142 -4946
rect 22063 -5013 22142 -5002
rect 3677 -5476 3756 -5465
rect 3677 -5532 3688 -5476
rect 3744 -5532 3756 -5476
rect 3677 -5543 3756 -5532
rect 6241 -5821 6320 -5810
rect 2750 -5833 2829 -5822
rect 2750 -5889 2761 -5833
rect 2817 -5889 2829 -5833
rect 6241 -5877 6252 -5821
rect 6308 -5877 6320 -5821
rect 6241 -5888 6320 -5877
rect 7424 -5841 7503 -5830
rect 2750 -5900 2829 -5889
rect 7424 -5897 7435 -5841
rect 7491 -5897 7503 -5841
rect 7424 -5908 7503 -5897
rect 9815 -5852 9894 -5841
rect 9815 -5908 9826 -5852
rect 9882 -5908 9894 -5852
rect 9815 -5919 9894 -5908
rect 112 -6132 525 -6069
rect 2748 -6006 2827 -5995
rect 2748 -6062 2759 -6006
rect 2815 -6062 2827 -6006
rect 2748 -6073 2827 -6062
rect 6239 -5997 6318 -5986
rect 6239 -6053 6250 -5997
rect 6306 -6053 6318 -5997
rect 9814 -6033 9893 -6022
rect 6239 -6064 6318 -6053
rect 7415 -6058 7494 -6047
rect 7415 -6114 7426 -6058
rect 7482 -6114 7494 -6058
rect 9814 -6089 9825 -6033
rect 9881 -6089 9893 -6033
rect 9814 -6100 9893 -6089
rect 7415 -6125 7494 -6114
rect 112 -6134 377 -6132
rect 112 -9090 177 -6134
rect 917 -6934 996 -6923
rect 917 -6990 928 -6934
rect 984 -6990 996 -6934
rect 917 -7001 996 -6990
rect 1136 -6937 1215 -6926
rect 1136 -6993 1147 -6937
rect 1203 -6993 1215 -6937
rect 1136 -7004 1215 -6993
rect 6340 -7045 6417 -7042
rect 6686 -7045 6763 -7041
rect 7125 -7045 7202 -7039
rect 7277 -7045 7354 -7039
rect 6340 -7051 7354 -7045
rect 6340 -7053 7137 -7051
rect 6340 -7054 6698 -7053
rect 6340 -7106 6352 -7054
rect 6404 -7057 6698 -7054
rect 6404 -7106 6513 -7057
rect 6340 -7109 6513 -7106
rect 6565 -7105 6698 -7057
rect 6750 -7103 7137 -7053
rect 7189 -7103 7289 -7051
rect 7341 -7103 7354 -7051
rect 6750 -7105 7354 -7103
rect 6565 -7109 7354 -7105
rect 6340 -7111 7354 -7109
rect 6340 -7118 6417 -7111
rect 6501 -7121 6578 -7111
rect 6686 -7117 6763 -7111
rect 7125 -7115 7202 -7111
rect 7277 -7115 7354 -7111
rect 11378 -7240 11497 -7216
rect 11378 -7296 11418 -7240
rect 11474 -7296 11497 -7240
rect 11378 -7324 11497 -7296
rect 22982 -7512 23054 -4655
rect 32392 -4747 32471 -2763
rect 31846 -4826 32471 -4747
rect 23369 -4951 23448 -4940
rect 23369 -5007 23380 -4951
rect 23436 -5007 23448 -4951
rect 23369 -5018 23448 -5007
rect 23591 -4943 23670 -4932
rect 23591 -4999 23602 -4943
rect 23658 -4999 23670 -4943
rect 23591 -5010 23670 -4999
rect 23980 -4948 24374 -4941
rect 23980 -5000 24094 -4948
rect 24146 -5000 24267 -4948
rect 24319 -4952 24374 -4948
rect 24319 -5000 24903 -4952
rect 23980 -5015 24903 -5000
rect 24840 -5109 24903 -5015
rect 31846 -5978 31925 -4826
rect 31846 -5981 31936 -5978
rect 26706 -5994 26785 -5983
rect 26706 -6050 26717 -5994
rect 26773 -6050 26785 -5994
rect 26706 -6061 26785 -6050
rect 27047 -5996 27126 -5985
rect 27047 -6052 27058 -5996
rect 27114 -6052 27126 -5996
rect 27047 -6063 27126 -6052
rect 31661 -5994 31936 -5981
rect 31661 -5998 31869 -5994
rect 31661 -6050 31689 -5998
rect 31741 -6046 31869 -5998
rect 31921 -6046 31936 -5994
rect 31741 -6050 31936 -6046
rect 31661 -6060 31936 -6050
rect 31675 -6067 31756 -6060
rect 31855 -6063 31936 -6060
rect 18969 -7584 23054 -7512
rect 3773 -7760 3852 -7749
rect 3773 -7816 3784 -7760
rect 3840 -7816 3852 -7760
rect 3773 -7827 3852 -7816
rect 6209 -7778 6291 -7767
rect 6209 -7834 6222 -7778
rect 6278 -7834 6291 -7778
rect 6209 -7844 6291 -7834
rect 9689 -7780 9768 -7769
rect 9689 -7836 9700 -7780
rect 9756 -7836 9768 -7780
rect 9689 -7847 9768 -7836
rect 10932 -7782 11011 -7771
rect 10932 -7838 10943 -7782
rect 10999 -7838 11011 -7782
rect 10932 -7849 11011 -7838
rect 13387 -7805 13466 -7794
rect 18969 -7799 19041 -7584
rect 13387 -7861 13398 -7805
rect 13454 -7861 13466 -7805
rect 13387 -7872 13466 -7861
rect 17862 -7871 19041 -7799
rect 6210 -7930 6292 -7919
rect 3768 -7942 3847 -7931
rect 3768 -7998 3779 -7942
rect 3835 -7998 3847 -7942
rect 6210 -7986 6223 -7930
rect 6279 -7986 6292 -7930
rect 6210 -7996 6292 -7986
rect 9693 -7945 9772 -7934
rect 3768 -8009 3847 -7998
rect 9693 -8001 9704 -7945
rect 9760 -8001 9772 -7945
rect 17862 -7969 17934 -7871
rect 9693 -8012 9772 -8001
rect 10930 -8000 11009 -7989
rect 10930 -8056 10941 -8000
rect 10997 -8056 11009 -8000
rect 10930 -8067 11009 -8056
rect 13385 -8020 13464 -8009
rect 13385 -8076 13396 -8020
rect 13452 -8076 13464 -8020
rect 13385 -8087 13464 -8076
rect 17862 -8021 17877 -7969
rect 17929 -8021 17934 -7969
rect 307 -8113 386 -8102
rect 307 -8169 318 -8113
rect 374 -8169 386 -8113
rect 307 -8180 386 -8169
rect 490 -8112 569 -8101
rect 490 -8168 501 -8112
rect 557 -8168 569 -8112
rect 490 -8179 569 -8168
rect 17862 -8113 17934 -8021
rect 17862 -8128 18113 -8113
rect 17862 -8180 17897 -8128
rect 17949 -8180 18113 -8128
rect 17862 -8185 18113 -8180
rect 2891 -8823 2973 -8812
rect 2891 -8826 2904 -8823
rect 2787 -8879 2904 -8826
rect 2960 -8826 2973 -8823
rect 3138 -8823 3220 -8812
rect 3138 -8826 3151 -8823
rect 2960 -8879 3151 -8826
rect 3207 -8826 3220 -8823
rect 3207 -8879 3264 -8826
rect 2787 -8891 3264 -8879
rect 634 -8925 713 -8914
rect 634 -8981 645 -8925
rect 701 -8981 713 -8925
rect 634 -8992 713 -8981
rect 911 -8924 990 -8913
rect 911 -8980 922 -8924
rect 978 -8980 990 -8924
rect 911 -8991 990 -8980
rect 2787 -9090 2852 -8891
rect 112 -9155 2852 -9090
rect 1480 -9246 2100 -9240
rect 1480 -9252 2010 -9246
rect 1480 -9255 1859 -9252
rect 1480 -9257 1732 -9255
rect 1480 -9262 1615 -9257
rect 1480 -9318 1500 -9262
rect 1556 -9313 1615 -9262
rect 1671 -9311 1732 -9257
rect 1788 -9308 1859 -9255
rect 1915 -9302 2010 -9252
rect 2066 -9302 2100 -9246
rect 1915 -9308 2100 -9302
rect 1788 -9311 2100 -9308
rect 1671 -9313 2100 -9311
rect 1556 -9318 2100 -9313
rect 1480 -9380 2100 -9318
rect 1480 -9382 1627 -9380
rect 1683 -9382 2100 -9380
rect 1480 -9438 1512 -9382
rect 1568 -9436 1627 -9382
rect 1683 -9436 1770 -9382
rect 1568 -9438 1770 -9436
rect 1826 -9438 1900 -9382
rect 1956 -9384 2100 -9382
rect 1956 -9438 2024 -9384
rect 1480 -9440 2024 -9438
rect 2080 -9440 2100 -9384
rect 1480 -9460 2100 -9440
rect 11128 -9457 11694 -9418
rect 11128 -9463 11424 -9457
rect 11480 -9459 11694 -9457
rect 11128 -9466 11282 -9463
rect 11128 -9522 11158 -9466
rect 11214 -9519 11282 -9466
rect 11338 -9513 11424 -9463
rect 11480 -9513 11568 -9459
rect 11338 -9515 11568 -9513
rect 11624 -9515 11694 -9459
rect 11338 -9519 11694 -9515
rect 11214 -9522 11694 -9519
rect 11128 -9574 11694 -9522
rect 11128 -9576 11421 -9574
rect 11128 -9581 11281 -9576
rect 11128 -9637 11154 -9581
rect 11210 -9632 11281 -9581
rect 11337 -9630 11421 -9576
rect 11477 -9578 11694 -9574
rect 11477 -9630 11562 -9578
rect 11337 -9632 11562 -9630
rect 11210 -9634 11562 -9632
rect 11618 -9634 11694 -9578
rect 11210 -9637 11694 -9634
rect 11128 -9656 11694 -9637
rect 19341 -9450 19907 -9411
rect 19341 -9456 19637 -9450
rect 19693 -9452 19907 -9450
rect 19341 -9459 19495 -9456
rect 19341 -9515 19371 -9459
rect 19427 -9512 19495 -9459
rect 19551 -9506 19637 -9456
rect 19693 -9506 19781 -9452
rect 19551 -9508 19781 -9506
rect 19837 -9508 19907 -9452
rect 19551 -9512 19907 -9508
rect 19427 -9515 19907 -9512
rect 19341 -9567 19907 -9515
rect 19341 -9569 19634 -9567
rect 19341 -9574 19494 -9569
rect 19341 -9630 19367 -9574
rect 19423 -9625 19494 -9574
rect 19550 -9623 19634 -9569
rect 19690 -9571 19907 -9567
rect 19690 -9623 19775 -9571
rect 19550 -9625 19775 -9623
rect 19423 -9627 19775 -9625
rect 19831 -9627 19907 -9571
rect 19423 -9630 19907 -9627
rect 26403 -9431 26969 -9392
rect 26403 -9437 26699 -9431
rect 26755 -9433 26969 -9431
rect 26403 -9440 26557 -9437
rect 26403 -9496 26433 -9440
rect 26489 -9493 26557 -9440
rect 26613 -9487 26699 -9437
rect 26755 -9487 26843 -9433
rect 26613 -9489 26843 -9487
rect 26899 -9489 26969 -9433
rect 26613 -9493 26969 -9489
rect 26489 -9496 26969 -9493
rect 26403 -9548 26969 -9496
rect 26403 -9550 26696 -9548
rect 26403 -9555 26556 -9550
rect 26403 -9611 26429 -9555
rect 26485 -9606 26556 -9555
rect 26612 -9604 26696 -9550
rect 26752 -9552 26969 -9548
rect 26752 -9604 26837 -9552
rect 26612 -9606 26837 -9604
rect 26485 -9608 26837 -9606
rect 26893 -9608 26969 -9552
rect 26485 -9611 26969 -9608
rect 26403 -9630 26969 -9611
rect 33208 -9429 33774 -9390
rect 33208 -9435 33504 -9429
rect 33560 -9431 33774 -9429
rect 33208 -9438 33362 -9435
rect 33208 -9494 33238 -9438
rect 33294 -9491 33362 -9438
rect 33418 -9485 33504 -9435
rect 33560 -9485 33648 -9431
rect 33418 -9487 33648 -9485
rect 33704 -9487 33774 -9431
rect 33418 -9491 33774 -9487
rect 33294 -9494 33774 -9491
rect 33208 -9546 33774 -9494
rect 33208 -9548 33501 -9546
rect 33208 -9553 33361 -9548
rect 33208 -9609 33234 -9553
rect 33290 -9604 33361 -9553
rect 33417 -9602 33501 -9548
rect 33557 -9550 33774 -9546
rect 33557 -9602 33642 -9550
rect 33417 -9604 33642 -9602
rect 33290 -9606 33642 -9604
rect 33698 -9606 33774 -9550
rect 33290 -9609 33774 -9606
rect 33208 -9628 33774 -9609
rect 19341 -9649 19907 -9630
rect 15100 -9880 15666 -9841
rect 15100 -9886 15396 -9880
rect 15452 -9882 15666 -9880
rect 15100 -9889 15254 -9886
rect 5214 -9962 5780 -9923
rect 5214 -9968 5510 -9962
rect 5566 -9964 5780 -9962
rect 5214 -9971 5368 -9968
rect 5214 -10027 5244 -9971
rect 5300 -10024 5368 -9971
rect 5424 -10018 5510 -9968
rect 5566 -10018 5654 -9964
rect 5424 -10020 5654 -10018
rect 5710 -10020 5780 -9964
rect 5424 -10024 5780 -10020
rect 5300 -10027 5780 -10024
rect 5214 -10079 5780 -10027
rect 15100 -9945 15130 -9889
rect 15186 -9942 15254 -9889
rect 15310 -9936 15396 -9886
rect 15452 -9936 15540 -9882
rect 15310 -9938 15540 -9936
rect 15596 -9938 15666 -9882
rect 15310 -9942 15666 -9938
rect 15186 -9945 15666 -9942
rect 15100 -9997 15666 -9945
rect 15100 -9999 15393 -9997
rect 15100 -10004 15253 -9999
rect 15100 -10060 15126 -10004
rect 15182 -10055 15253 -10004
rect 15309 -10053 15393 -9999
rect 15449 -10001 15666 -9997
rect 15449 -10053 15534 -10001
rect 15309 -10055 15534 -10053
rect 15182 -10057 15534 -10055
rect 15590 -10057 15666 -10001
rect 22631 -9850 23197 -9811
rect 22631 -9856 22927 -9850
rect 22983 -9852 23197 -9850
rect 22631 -9859 22785 -9856
rect 22631 -9915 22661 -9859
rect 22717 -9912 22785 -9859
rect 22841 -9906 22927 -9856
rect 22983 -9906 23071 -9852
rect 22841 -9908 23071 -9906
rect 23127 -9908 23197 -9852
rect 22841 -9912 23197 -9908
rect 22717 -9915 23197 -9912
rect 22631 -9967 23197 -9915
rect 22631 -9969 22924 -9967
rect 22631 -9974 22784 -9969
rect 22631 -10030 22657 -9974
rect 22713 -10025 22784 -9974
rect 22840 -10023 22924 -9969
rect 22980 -9971 23197 -9967
rect 22980 -10023 23065 -9971
rect 22840 -10025 23065 -10023
rect 22713 -10027 23065 -10025
rect 23121 -10027 23197 -9971
rect 22713 -10030 23197 -10027
rect 22631 -10049 23197 -10030
rect 15182 -10060 15666 -10057
rect 15100 -10079 15666 -10060
rect 5214 -10081 5507 -10079
rect 5214 -10086 5367 -10081
rect 5214 -10142 5240 -10086
rect 5296 -10137 5367 -10086
rect 5423 -10135 5507 -10081
rect 5563 -10083 5780 -10079
rect 5563 -10135 5648 -10083
rect 5423 -10137 5648 -10135
rect 5296 -10139 5648 -10137
rect 5704 -10139 5780 -10083
rect 5296 -10142 5780 -10139
rect 5214 -10161 5780 -10142
<< via2 >>
rect 22919 12081 22975 12083
rect 22777 12075 22833 12077
rect 22653 12072 22709 12074
rect 22653 12020 22655 12072
rect 22655 12020 22707 12072
rect 22707 12020 22709 12072
rect 22777 12023 22779 12075
rect 22779 12023 22831 12075
rect 22831 12023 22833 12075
rect 22919 12029 22921 12081
rect 22921 12029 22973 12081
rect 22973 12029 22975 12081
rect 22919 12027 22975 12029
rect 23063 12079 23119 12081
rect 23063 12027 23065 12079
rect 23065 12027 23117 12079
rect 23117 12027 23119 12079
rect 23063 12025 23119 12027
rect 22777 12021 22833 12023
rect 22653 12018 22709 12020
rect 5263 11965 5319 11967
rect 5121 11959 5177 11961
rect 4997 11956 5053 11958
rect 4997 11904 4999 11956
rect 4999 11904 5051 11956
rect 5051 11904 5053 11956
rect 5121 11907 5123 11959
rect 5123 11907 5175 11959
rect 5175 11907 5177 11959
rect 5263 11913 5265 11965
rect 5265 11913 5317 11965
rect 5317 11913 5319 11965
rect 5263 11911 5319 11913
rect 5407 11963 5463 11965
rect 5407 11911 5409 11963
rect 5409 11911 5461 11963
rect 5461 11911 5463 11963
rect 5407 11909 5463 11911
rect 5121 11905 5177 11907
rect 4997 11902 5053 11904
rect 5260 11848 5316 11850
rect 5120 11846 5176 11848
rect 4993 11841 5049 11843
rect 4993 11789 4995 11841
rect 4995 11789 5047 11841
rect 5047 11789 5049 11841
rect 5120 11794 5122 11846
rect 5122 11794 5174 11846
rect 5174 11794 5176 11846
rect 5260 11796 5262 11848
rect 5262 11796 5314 11848
rect 5314 11796 5316 11848
rect 5260 11794 5316 11796
rect 5401 11844 5457 11846
rect 5120 11792 5176 11794
rect 5401 11792 5403 11844
rect 5403 11792 5455 11844
rect 5455 11792 5457 11844
rect 5401 11790 5457 11792
rect 4993 11787 5049 11789
rect 15396 11955 15452 11957
rect 15254 11949 15310 11951
rect 15130 11946 15186 11948
rect 15130 11894 15132 11946
rect 15132 11894 15184 11946
rect 15184 11894 15186 11946
rect 15254 11897 15256 11949
rect 15256 11897 15308 11949
rect 15308 11897 15310 11949
rect 15396 11903 15398 11955
rect 15398 11903 15450 11955
rect 15450 11903 15452 11955
rect 15396 11901 15452 11903
rect 15540 11953 15596 11955
rect 15540 11901 15542 11953
rect 15542 11901 15594 11953
rect 15594 11901 15596 11953
rect 15540 11899 15596 11901
rect 15254 11895 15310 11897
rect 15130 11892 15186 11894
rect 22916 11964 22972 11966
rect 22776 11962 22832 11964
rect 22649 11957 22705 11959
rect 22649 11905 22651 11957
rect 22651 11905 22703 11957
rect 22703 11905 22705 11957
rect 22776 11910 22778 11962
rect 22778 11910 22830 11962
rect 22830 11910 22832 11962
rect 22916 11912 22918 11964
rect 22918 11912 22970 11964
rect 22970 11912 22972 11964
rect 22916 11910 22972 11912
rect 23057 11960 23113 11962
rect 22776 11908 22832 11910
rect 23057 11908 23059 11960
rect 23059 11908 23111 11960
rect 23111 11908 23113 11960
rect 23057 11906 23113 11908
rect 22649 11903 22705 11905
rect 15393 11838 15449 11840
rect 15253 11836 15309 11838
rect 15126 11831 15182 11833
rect 15126 11779 15128 11831
rect 15128 11779 15180 11831
rect 15180 11779 15182 11831
rect 15253 11784 15255 11836
rect 15255 11784 15307 11836
rect 15307 11784 15309 11836
rect 15393 11786 15395 11838
rect 15395 11786 15447 11838
rect 15447 11786 15449 11838
rect 15393 11784 15449 11786
rect 15534 11834 15590 11836
rect 15253 11782 15309 11784
rect 15534 11782 15536 11834
rect 15536 11782 15588 11834
rect 15588 11782 15590 11834
rect 15534 11780 15590 11782
rect 15126 11777 15182 11779
rect 33278 11762 33334 11764
rect 33136 11756 33192 11758
rect 11559 11744 11615 11746
rect 11417 11738 11473 11740
rect 11293 11735 11349 11737
rect 11293 11683 11295 11735
rect 11295 11683 11347 11735
rect 11347 11683 11349 11735
rect 11417 11686 11419 11738
rect 11419 11686 11471 11738
rect 11471 11686 11473 11738
rect 11559 11692 11561 11744
rect 11561 11692 11613 11744
rect 11613 11692 11615 11744
rect 11559 11690 11615 11692
rect 11703 11742 11759 11744
rect 11703 11690 11705 11742
rect 11705 11690 11757 11742
rect 11757 11690 11759 11742
rect 11703 11688 11759 11690
rect 11417 11684 11473 11686
rect 11293 11681 11349 11683
rect 1900 11631 1956 11633
rect 1758 11625 1814 11627
rect 1634 11622 1690 11624
rect 1634 11570 1636 11622
rect 1636 11570 1688 11622
rect 1688 11570 1690 11622
rect 1758 11573 1760 11625
rect 1760 11573 1812 11625
rect 1812 11573 1814 11625
rect 1900 11579 1902 11631
rect 1902 11579 1954 11631
rect 1954 11579 1956 11631
rect 1900 11577 1956 11579
rect 2044 11629 2100 11631
rect 2044 11577 2046 11629
rect 2046 11577 2098 11629
rect 2098 11577 2100 11629
rect 2044 11575 2100 11577
rect 1758 11571 1814 11573
rect 1634 11568 1690 11570
rect 11556 11627 11612 11629
rect 11416 11625 11472 11627
rect 11289 11620 11345 11622
rect 11289 11568 11291 11620
rect 11291 11568 11343 11620
rect 11343 11568 11345 11620
rect 11416 11573 11418 11625
rect 11418 11573 11470 11625
rect 11470 11573 11472 11625
rect 11556 11575 11558 11627
rect 11558 11575 11610 11627
rect 11610 11575 11612 11627
rect 11556 11573 11612 11575
rect 11697 11623 11753 11625
rect 11416 11571 11472 11573
rect 11697 11571 11699 11623
rect 11699 11571 11751 11623
rect 11751 11571 11753 11623
rect 11697 11569 11753 11571
rect 11289 11566 11345 11568
rect 19424 11708 19480 11710
rect 19282 11702 19338 11704
rect 19158 11699 19214 11701
rect 19158 11647 19160 11699
rect 19160 11647 19212 11699
rect 19212 11647 19214 11699
rect 19282 11650 19284 11702
rect 19284 11650 19336 11702
rect 19336 11650 19338 11702
rect 19424 11656 19426 11708
rect 19426 11656 19478 11708
rect 19478 11656 19480 11708
rect 19424 11654 19480 11656
rect 19568 11706 19624 11708
rect 19568 11654 19570 11706
rect 19570 11654 19622 11706
rect 19622 11654 19624 11706
rect 19568 11652 19624 11654
rect 19282 11648 19338 11650
rect 19158 11645 19214 11647
rect 19421 11591 19477 11593
rect 19281 11589 19337 11591
rect 1897 11514 1953 11516
rect 1757 11512 1813 11514
rect 1630 11507 1686 11509
rect 1630 11455 1632 11507
rect 1632 11455 1684 11507
rect 1684 11455 1686 11507
rect 1757 11460 1759 11512
rect 1759 11460 1811 11512
rect 1811 11460 1813 11512
rect 1897 11462 1899 11514
rect 1899 11462 1951 11514
rect 1951 11462 1953 11514
rect 1897 11460 1953 11462
rect 2038 11510 2094 11512
rect 1757 11458 1813 11460
rect 2038 11458 2040 11510
rect 2040 11458 2092 11510
rect 2092 11458 2094 11510
rect 2038 11456 2094 11458
rect 19154 11584 19210 11586
rect 19154 11532 19156 11584
rect 19156 11532 19208 11584
rect 19208 11532 19210 11584
rect 19281 11537 19283 11589
rect 19283 11537 19335 11589
rect 19335 11537 19337 11589
rect 19421 11539 19423 11591
rect 19423 11539 19475 11591
rect 19475 11539 19477 11591
rect 19421 11537 19477 11539
rect 19562 11587 19618 11589
rect 19281 11535 19337 11537
rect 19562 11535 19564 11587
rect 19564 11535 19616 11587
rect 19616 11535 19618 11587
rect 19562 11533 19618 11535
rect 19154 11530 19210 11532
rect 26405 11690 26461 11692
rect 26263 11684 26319 11686
rect 26139 11681 26195 11683
rect 26139 11629 26141 11681
rect 26141 11629 26193 11681
rect 26193 11629 26195 11681
rect 26263 11632 26265 11684
rect 26265 11632 26317 11684
rect 26317 11632 26319 11684
rect 26405 11638 26407 11690
rect 26407 11638 26459 11690
rect 26459 11638 26461 11690
rect 26405 11636 26461 11638
rect 26549 11688 26605 11690
rect 26549 11636 26551 11688
rect 26551 11636 26603 11688
rect 26603 11636 26605 11688
rect 26549 11634 26605 11636
rect 26263 11630 26319 11632
rect 26139 11627 26195 11629
rect 26402 11573 26458 11575
rect 26262 11571 26318 11573
rect 26135 11566 26191 11568
rect 26135 11514 26137 11566
rect 26137 11514 26189 11566
rect 26189 11514 26191 11566
rect 26262 11519 26264 11571
rect 26264 11519 26316 11571
rect 26316 11519 26318 11571
rect 26402 11521 26404 11573
rect 26404 11521 26456 11573
rect 26456 11521 26458 11573
rect 26402 11519 26458 11521
rect 26543 11569 26599 11571
rect 26262 11517 26318 11519
rect 26543 11517 26545 11569
rect 26545 11517 26597 11569
rect 26597 11517 26599 11569
rect 26543 11515 26599 11517
rect 33012 11753 33068 11755
rect 33012 11701 33014 11753
rect 33014 11701 33066 11753
rect 33066 11701 33068 11753
rect 33136 11704 33138 11756
rect 33138 11704 33190 11756
rect 33190 11704 33192 11756
rect 33278 11710 33280 11762
rect 33280 11710 33332 11762
rect 33332 11710 33334 11762
rect 33278 11708 33334 11710
rect 33422 11760 33478 11762
rect 33422 11708 33424 11760
rect 33424 11708 33476 11760
rect 33476 11708 33478 11760
rect 33422 11706 33478 11708
rect 33136 11702 33192 11704
rect 33012 11699 33068 11701
rect 33275 11645 33331 11647
rect 33135 11643 33191 11645
rect 33008 11638 33064 11640
rect 33008 11586 33010 11638
rect 33010 11586 33062 11638
rect 33062 11586 33064 11638
rect 33135 11591 33137 11643
rect 33137 11591 33189 11643
rect 33189 11591 33191 11643
rect 33275 11593 33277 11645
rect 33277 11593 33329 11645
rect 33329 11593 33331 11645
rect 33275 11591 33331 11593
rect 33416 11641 33472 11643
rect 33135 11589 33191 11591
rect 33416 11589 33418 11641
rect 33418 11589 33470 11641
rect 33470 11589 33472 11641
rect 33416 11587 33472 11589
rect 33008 11584 33064 11586
rect 26135 11512 26191 11514
rect 1630 11453 1686 11455
rect 18247 11268 18303 11324
rect 18463 11270 18519 11326
rect 5156 10570 5212 10572
rect 5156 10518 5158 10570
rect 5158 10518 5210 10570
rect 5210 10518 5212 10570
rect 5156 10516 5212 10518
rect 1703 9573 1759 9575
rect 1703 9521 1705 9573
rect 1705 9521 1757 9573
rect 1757 9521 1759 9573
rect 1703 9519 1759 9521
rect 1075 8721 1131 8777
rect 1076 8648 1132 8650
rect 1076 8596 1078 8648
rect 1078 8596 1130 8648
rect 1130 8596 1132 8648
rect 1076 8594 1132 8596
rect 9867 8718 9923 8774
rect 19521 8804 19577 8806
rect 19521 8752 19523 8804
rect 19523 8752 19575 8804
rect 19575 8752 19577 8804
rect 19521 8750 19577 8752
rect 9857 8654 9913 8657
rect 9857 8602 9902 8654
rect 9902 8602 9913 8654
rect 9857 8601 9913 8602
rect 10200 8542 10256 8544
rect 10200 8490 10202 8542
rect 10202 8490 10254 8542
rect 10254 8490 10256 8542
rect 10200 8488 10256 8490
rect 10340 8541 10396 8543
rect 10340 8489 10342 8541
rect 10342 8489 10394 8541
rect 10394 8489 10396 8541
rect 10340 8487 10396 8489
rect 10205 8430 10261 8432
rect 10205 8378 10207 8430
rect 10207 8378 10259 8430
rect 10259 8378 10261 8430
rect 10205 8376 10261 8378
rect 11530 8478 11586 8480
rect 11530 8426 11532 8478
rect 11532 8426 11584 8478
rect 11584 8426 11586 8478
rect 11530 8424 11586 8426
rect 26568 8415 26624 8417
rect 26568 8363 26570 8415
rect 26570 8363 26622 8415
rect 26622 8363 26624 8415
rect 26568 8361 26624 8363
rect 21698 8169 21754 8225
rect 21835 8168 21891 8224
rect 11731 8030 11787 8086
rect 11895 8032 11951 8088
rect 18190 8052 18246 8108
rect 18373 8053 18429 8109
rect 1683 7999 1739 8001
rect 1683 7947 1685 7999
rect 1685 7947 1737 7999
rect 1737 7947 1739 7999
rect 1683 7945 1739 7947
rect 10299 7846 10355 7848
rect 10299 7794 10301 7846
rect 10301 7794 10353 7846
rect 10353 7794 10355 7846
rect 10299 7792 10355 7794
rect 10469 7846 10525 7848
rect 10469 7794 10471 7846
rect 10471 7794 10523 7846
rect 10523 7794 10525 7846
rect 10469 7792 10525 7794
rect 11515 7897 11571 7899
rect 11515 7845 11517 7897
rect 11517 7845 11569 7897
rect 11569 7845 11571 7897
rect 11515 7843 11571 7845
rect 19469 7609 19525 7611
rect 19469 7557 19471 7609
rect 19471 7557 19523 7609
rect 19523 7557 19525 7609
rect 19469 7555 19525 7557
rect 7942 7139 7998 7141
rect 7942 7087 7943 7139
rect 7943 7087 7995 7139
rect 7995 7087 7998 7139
rect 7942 7085 7998 7087
rect 7949 6993 8005 6995
rect 7949 6941 7950 6993
rect 7950 6941 8002 6993
rect 8002 6941 8005 6993
rect 7949 6939 8005 6941
rect 18603 6000 18659 6056
rect 18726 6002 18782 6058
rect 18604 5886 18660 5942
rect 18725 5893 18781 5949
rect 15519 5734 15575 5736
rect 15519 5682 15521 5734
rect 15521 5682 15573 5734
rect 15573 5682 15575 5734
rect 15519 5680 15575 5682
rect 5151 5348 5207 5350
rect 5151 5296 5153 5348
rect 5153 5296 5205 5348
rect 5205 5296 5207 5348
rect 5151 5294 5207 5296
rect 22904 5677 22960 5733
rect 1424 2956 1480 3012
rect 3084 3009 3140 3011
rect 3084 2957 3085 3009
rect 3085 2957 3137 3009
rect 3137 2957 3140 3009
rect 3084 2955 3140 2957
rect 3374 3010 3430 3012
rect 3374 2958 3375 3010
rect 3375 2958 3427 3010
rect 3427 2958 3430 3010
rect 3374 2956 3430 2958
rect 1306 2877 1362 2933
rect 1425 2818 1481 2874
rect 9855 3431 9911 3435
rect 9855 3379 9903 3431
rect 9903 3379 9911 3431
rect 9854 3266 9910 3322
rect 19476 3612 19532 3614
rect 19476 3560 19478 3612
rect 19478 3560 19530 3612
rect 19530 3560 19532 3612
rect 19476 3558 19532 3560
rect 11322 3224 11378 3226
rect 11322 3172 11324 3224
rect 11324 3172 11376 3224
rect 11376 3172 11378 3224
rect 11322 3170 11378 3172
rect 11543 3219 11599 3221
rect 11543 3167 11545 3219
rect 11545 3167 11597 3219
rect 11597 3167 11599 3219
rect 11543 3165 11599 3167
rect 11738 3229 11794 3231
rect 11738 3177 11740 3229
rect 11740 3177 11792 3229
rect 11792 3177 11794 3229
rect 11738 3175 11794 3177
rect 1739 2803 1795 2805
rect 1739 2751 1741 2803
rect 1741 2751 1793 2803
rect 1793 2751 1795 2803
rect 1739 2749 1795 2751
rect 10095 2825 10151 2881
rect 10333 2826 10389 2882
rect 11496 2717 11552 2719
rect 11496 2665 11498 2717
rect 11498 2665 11550 2717
rect 11550 2665 11552 2717
rect 11496 2663 11552 2665
rect 11034 2316 11090 2318
rect 11034 2264 11036 2316
rect 11036 2264 11088 2316
rect 11088 2264 11090 2316
rect 11034 2262 11090 2264
rect 11039 2181 11095 2183
rect 11039 2129 11041 2181
rect 11041 2129 11093 2181
rect 11093 2129 11095 2181
rect 11039 2127 11095 2129
rect 7662 390 7718 393
rect 7662 338 7663 390
rect 7663 338 7715 390
rect 7715 338 7718 390
rect 7662 337 7718 338
rect 7817 391 7873 394
rect 7817 339 7818 391
rect 7818 339 7870 391
rect 7870 339 7873 391
rect 7817 338 7873 339
rect 4511 113 4567 115
rect 4511 61 4512 113
rect 4512 61 4564 113
rect 4564 61 4567 113
rect 4511 59 4567 61
rect 11260 96 11316 152
rect 11494 100 11550 156
rect 2367 -53 2423 -51
rect 2367 -105 2368 -53
rect 2368 -105 2420 -53
rect 2420 -105 2423 -53
rect 2978 -75 3034 -73
rect 2367 -107 2423 -105
rect 2554 -116 2610 -114
rect 2554 -168 2555 -116
rect 2555 -168 2607 -116
rect 2607 -168 2610 -116
rect 2554 -170 2610 -168
rect 2978 -127 2979 -75
rect 2979 -127 3031 -75
rect 3031 -127 3034 -75
rect 3182 -77 3238 -75
rect 2978 -129 3034 -127
rect 3182 -129 3183 -77
rect 3183 -129 3235 -77
rect 3235 -129 3238 -77
rect 13928 57 13984 113
rect 14138 58 14194 114
rect 15215 517 15271 519
rect 15215 465 15217 517
rect 15217 465 15269 517
rect 15269 465 15271 517
rect 15215 463 15271 465
rect 6036 13 6092 16
rect 6036 -39 6037 13
rect 6037 -39 6089 13
rect 6089 -39 6092 13
rect 6036 -40 6092 -39
rect 3182 -131 3238 -129
rect 6301 -87 6357 -31
rect 6495 -86 6551 -30
rect 22515 320 22571 376
rect 25831 2944 25887 3000
rect 25979 2944 26035 3000
rect 26136 2948 26192 3004
rect 26465 2687 26521 2689
rect 26465 2635 26467 2687
rect 26467 2635 26519 2687
rect 26519 2635 26521 2687
rect 26465 2633 26521 2635
rect 28948 1888 29004 1893
rect 28948 1837 28999 1888
rect 28999 1837 29004 1888
rect 29231 1887 29287 1892
rect 29231 1836 29282 1887
rect 29282 1836 29287 1887
rect 22690 318 22746 374
rect 14681 -89 14737 -33
rect 14884 -93 14940 -37
rect 533 -192 589 -190
rect 533 -244 534 -192
rect 534 -244 586 -192
rect 586 -244 589 -192
rect 533 -246 589 -244
rect 19491 -163 19547 -160
rect 19491 -215 19492 -163
rect 19492 -215 19544 -163
rect 19544 -215 19547 -163
rect 19491 -216 19547 -215
rect 1196 -285 1252 -229
rect 1348 -286 1404 -230
rect 23490 -137 23546 -136
rect 23490 -189 23493 -137
rect 23493 -189 23545 -137
rect 23545 -189 23546 -137
rect 23490 -192 23546 -189
rect 31710 2006 31766 2011
rect 31710 1955 31761 2006
rect 31761 1955 31766 2006
rect 529 -359 585 -357
rect 529 -411 530 -359
rect 530 -411 582 -359
rect 582 -411 585 -359
rect 4150 -375 4206 -373
rect 529 -413 585 -411
rect 3927 -379 3983 -377
rect 3927 -431 3928 -379
rect 3928 -431 3980 -379
rect 3980 -431 3983 -379
rect 4150 -427 4151 -375
rect 4151 -427 4203 -375
rect 4203 -427 4206 -375
rect 3927 -433 3983 -431
rect 4150 -429 4206 -427
rect 6044 -367 6100 -364
rect 6044 -419 6045 -367
rect 6045 -419 6097 -367
rect 6097 -419 6100 -367
rect 6044 -420 6100 -419
rect 23491 -306 23547 -305
rect 23491 -358 23494 -306
rect 23494 -358 23546 -306
rect 23546 -358 23547 -306
rect 23491 -361 23547 -358
rect 30480 -449 30536 -446
rect 30480 -501 30481 -449
rect 30481 -501 30533 -449
rect 30533 -501 30536 -449
rect 30480 -502 30536 -501
rect 30677 -442 30733 -439
rect 30677 -494 30678 -442
rect 30678 -494 30730 -442
rect 30730 -494 30733 -442
rect 30677 -495 30733 -494
rect 3823 -1209 3879 -1206
rect 3823 -1261 3824 -1209
rect 3824 -1261 3876 -1209
rect 3876 -1261 3879 -1209
rect 3823 -1262 3879 -1261
rect 6221 -1262 6277 -1259
rect 6221 -1314 6222 -1262
rect 6222 -1314 6274 -1262
rect 6274 -1314 6277 -1262
rect 6221 -1315 6277 -1314
rect 7426 -1205 7482 -1202
rect 7426 -1257 7427 -1205
rect 7427 -1257 7479 -1205
rect 7479 -1257 7482 -1205
rect 7426 -1258 7482 -1257
rect 9846 -1233 9902 -1230
rect 9846 -1285 9847 -1233
rect 9847 -1285 9899 -1233
rect 9899 -1285 9902 -1233
rect 9846 -1286 9902 -1285
rect 327 -1348 383 -1345
rect 327 -1400 328 -1348
rect 328 -1400 380 -1348
rect 380 -1400 383 -1348
rect 327 -1401 383 -1400
rect 2734 -1442 2790 -1439
rect 2734 -1494 2735 -1442
rect 2735 -1494 2787 -1442
rect 2787 -1494 2790 -1442
rect 2734 -1495 2790 -1494
rect 6226 -1431 6282 -1428
rect 6226 -1483 6227 -1431
rect 6227 -1483 6279 -1431
rect 6279 -1483 6282 -1431
rect 6226 -1484 6282 -1483
rect 334 -1532 390 -1529
rect 334 -1584 335 -1532
rect 335 -1584 387 -1532
rect 387 -1584 390 -1532
rect 334 -1585 390 -1584
rect 3819 -1515 3875 -1512
rect 3819 -1567 3820 -1515
rect 3820 -1567 3872 -1515
rect 3872 -1567 3875 -1515
rect 3819 -1568 3875 -1567
rect 7418 -1455 7474 -1452
rect 7418 -1507 7419 -1455
rect 7419 -1507 7471 -1455
rect 7471 -1507 7474 -1455
rect 7418 -1508 7474 -1507
rect 14901 -1652 14957 -1596
rect 1775 -2430 1831 -2428
rect 1775 -2482 1777 -2430
rect 1777 -2482 1829 -2430
rect 1829 -2482 1831 -2430
rect 1775 -2484 1831 -2482
rect 21886 -1649 21942 -1648
rect 21886 -1701 21890 -1649
rect 21890 -1701 21942 -1649
rect 21886 -1704 21942 -1701
rect 22328 -1650 22384 -1649
rect 22328 -1702 22331 -1650
rect 22331 -1702 22383 -1650
rect 22383 -1702 22384 -1650
rect 22328 -1705 22384 -1702
rect 14900 -1813 14956 -1757
rect 4355 -2387 4411 -2385
rect 4355 -2439 4356 -2387
rect 4356 -2439 4408 -2387
rect 4408 -2439 4411 -2387
rect 4355 -2441 4411 -2439
rect 3807 -2571 3863 -2568
rect 3807 -2623 3808 -2571
rect 3808 -2623 3860 -2571
rect 3860 -2623 3863 -2571
rect 3807 -2624 3863 -2623
rect 4067 -2573 4123 -2570
rect 4067 -2625 4068 -2573
rect 4068 -2625 4120 -2573
rect 4120 -2625 4123 -2573
rect 4067 -2626 4123 -2625
rect 498 -3288 554 -3285
rect 498 -3340 499 -3288
rect 499 -3340 551 -3288
rect 551 -3340 554 -3288
rect 498 -3341 554 -3340
rect 494 -3497 550 -3494
rect 494 -3549 495 -3497
rect 495 -3549 547 -3497
rect 547 -3549 550 -3497
rect 494 -3550 550 -3549
rect 776 -4368 832 -4365
rect 776 -4420 777 -4368
rect 777 -4420 829 -4368
rect 829 -4420 832 -4368
rect 776 -4421 832 -4420
rect 975 -4369 1031 -4366
rect 975 -4421 976 -4369
rect 976 -4421 1028 -4369
rect 1028 -4421 1031 -4369
rect 975 -4422 1031 -4421
rect 9706 -2542 9762 -2540
rect 9706 -2594 9707 -2542
rect 9707 -2594 9759 -2542
rect 9759 -2594 9762 -2542
rect 9706 -2596 9762 -2594
rect 9898 -2542 9954 -2540
rect 9898 -2594 9899 -2542
rect 9899 -2594 9951 -2542
rect 9951 -2594 9954 -2542
rect 9898 -2596 9954 -2594
rect 7291 -2971 7347 -2968
rect 7291 -3023 7292 -2971
rect 7292 -3023 7344 -2971
rect 7344 -3023 7347 -2971
rect 7291 -3024 7347 -3023
rect 7275 -3331 7331 -3328
rect 7275 -3383 7276 -3331
rect 7276 -3383 7328 -3331
rect 7328 -3383 7331 -3331
rect 7275 -3384 7331 -3383
rect 14760 -2773 14816 -2717
rect 14946 -2775 15002 -2719
rect 21784 -2662 21840 -2659
rect 21784 -2714 21785 -2662
rect 21785 -2714 21837 -2662
rect 21837 -2714 21840 -2662
rect 21784 -2715 21840 -2714
rect 21939 -2666 21995 -2663
rect 21939 -2718 21940 -2666
rect 21940 -2718 21992 -2666
rect 21992 -2718 21995 -2666
rect 21939 -2719 21995 -2718
rect 11603 -2798 11659 -2796
rect 11603 -2850 11605 -2798
rect 11605 -2850 11657 -2798
rect 11657 -2850 11659 -2798
rect 11603 -2852 11659 -2850
rect 17877 -2825 17933 -2824
rect 17877 -2877 17880 -2825
rect 17880 -2877 17932 -2825
rect 17932 -2877 17933 -2825
rect 17877 -2880 17933 -2877
rect 18135 -2825 18191 -2824
rect 18135 -2877 18138 -2825
rect 18138 -2877 18190 -2825
rect 18190 -2877 18191 -2825
rect 18135 -2880 18191 -2877
rect 22858 -1506 22914 -1450
rect 22855 -1677 22911 -1621
rect 31773 -436 31829 -433
rect 31773 -488 31774 -436
rect 31774 -488 31826 -436
rect 31826 -488 31829 -436
rect 31773 -489 31829 -488
rect 31959 -434 32015 -431
rect 31959 -486 31960 -434
rect 31960 -486 32012 -434
rect 32012 -486 32015 -434
rect 31959 -487 32015 -486
rect 11129 -3310 11185 -3307
rect 11129 -3362 11130 -3310
rect 11130 -3362 11182 -3310
rect 11182 -3362 11185 -3310
rect 11129 -3363 11185 -3362
rect 13363 -3304 13419 -3301
rect 13363 -3356 13364 -3304
rect 13364 -3356 13416 -3304
rect 13416 -3356 13419 -3304
rect 13363 -3357 13419 -3356
rect 13359 -3465 13415 -3462
rect 13359 -3517 13360 -3465
rect 13360 -3517 13412 -3465
rect 13412 -3517 13415 -3465
rect 13359 -3518 13415 -3517
rect 5576 -4202 5632 -4200
rect 5576 -4254 5578 -4202
rect 5578 -4254 5630 -4202
rect 5630 -4254 5632 -4202
rect 5576 -4256 5632 -4254
rect 15464 -4188 15520 -4186
rect 15464 -4240 15466 -4188
rect 15466 -4240 15518 -4188
rect 15518 -4240 15520 -4188
rect 15464 -4242 15520 -4240
rect 3623 -4523 3679 -4520
rect 3289 -4529 3345 -4526
rect 3289 -4581 3290 -4529
rect 3290 -4581 3342 -4529
rect 3342 -4581 3345 -4529
rect 3623 -4575 3624 -4523
rect 3624 -4575 3676 -4523
rect 3676 -4575 3679 -4523
rect 3623 -4576 3679 -4575
rect 3289 -4582 3345 -4581
rect 9810 -4533 9866 -4531
rect 316 -4672 372 -4669
rect 316 -4724 317 -4672
rect 317 -4724 369 -4672
rect 369 -4724 372 -4672
rect 316 -4725 372 -4724
rect 9573 -4542 9629 -4540
rect 9573 -4594 9574 -4542
rect 9574 -4594 9626 -4542
rect 9626 -4594 9629 -4542
rect 9810 -4585 9811 -4533
rect 9811 -4585 9863 -4533
rect 9863 -4585 9866 -4533
rect 9810 -4587 9866 -4585
rect 10408 -4542 10464 -4540
rect 9573 -4596 9629 -4594
rect 10408 -4594 10409 -4542
rect 10409 -4594 10461 -4542
rect 10461 -4594 10464 -4542
rect 10408 -4596 10464 -4594
rect 10655 -4542 10711 -4540
rect 10655 -4594 10656 -4542
rect 10656 -4594 10708 -4542
rect 10708 -4594 10711 -4542
rect 10655 -4596 10711 -4594
rect 314 -4829 370 -4826
rect 314 -4881 315 -4829
rect 315 -4881 367 -4829
rect 367 -4881 370 -4829
rect 314 -4882 370 -4881
rect 2372 -4839 2428 -4836
rect 2614 -4837 2670 -4834
rect -77 -5221 -21 -5218
rect -77 -5273 -76 -5221
rect -76 -5273 -24 -5221
rect -24 -5273 -21 -5221
rect -77 -5274 -21 -5273
rect -85 -5400 -29 -5397
rect -85 -5452 -84 -5400
rect -84 -5452 -32 -5400
rect -32 -5452 -29 -5400
rect -85 -5453 -29 -5452
rect 2372 -4891 2373 -4839
rect 2373 -4891 2425 -4839
rect 2425 -4891 2428 -4839
rect 2614 -4889 2615 -4837
rect 2615 -4889 2667 -4837
rect 2667 -4889 2670 -4837
rect 2614 -4890 2670 -4889
rect 2372 -4892 2428 -4891
rect 10667 -4691 10723 -4689
rect 10418 -4695 10474 -4693
rect 9824 -4706 9880 -4704
rect 9576 -4708 9632 -4706
rect 9576 -4760 9577 -4708
rect 9577 -4760 9629 -4708
rect 9629 -4760 9632 -4708
rect 9824 -4758 9825 -4706
rect 9825 -4758 9877 -4706
rect 9877 -4758 9880 -4706
rect 10418 -4747 10419 -4695
rect 10419 -4747 10471 -4695
rect 10471 -4747 10474 -4695
rect 10667 -4743 10668 -4691
rect 10668 -4743 10720 -4691
rect 10720 -4743 10723 -4691
rect 10667 -4745 10723 -4743
rect 10418 -4749 10474 -4747
rect 9824 -4760 9880 -4758
rect 9576 -4762 9632 -4760
rect 21030 -4928 21086 -4925
rect 21030 -4980 21031 -4928
rect 21031 -4980 21083 -4928
rect 21083 -4980 21086 -4928
rect 21030 -4981 21086 -4980
rect 21323 -4922 21379 -4919
rect 21323 -4974 21324 -4922
rect 21324 -4974 21376 -4922
rect 21376 -4974 21379 -4922
rect 21323 -4975 21379 -4974
rect 21905 -4957 21961 -4954
rect 21905 -5009 21906 -4957
rect 21906 -5009 21958 -4957
rect 21958 -5009 21961 -4957
rect 21905 -5010 21961 -5009
rect 22074 -4949 22130 -4946
rect 22074 -5001 22075 -4949
rect 22075 -5001 22127 -4949
rect 22127 -5001 22130 -4949
rect 22074 -5002 22130 -5001
rect 3688 -5479 3744 -5476
rect 3688 -5531 3689 -5479
rect 3689 -5531 3741 -5479
rect 3741 -5531 3744 -5479
rect 3688 -5532 3744 -5531
rect 2761 -5836 2817 -5833
rect 2761 -5888 2762 -5836
rect 2762 -5888 2814 -5836
rect 2814 -5888 2817 -5836
rect 2761 -5889 2817 -5888
rect 6252 -5824 6308 -5821
rect 6252 -5876 6253 -5824
rect 6253 -5876 6305 -5824
rect 6305 -5876 6308 -5824
rect 6252 -5877 6308 -5876
rect 7435 -5844 7491 -5841
rect 7435 -5896 7436 -5844
rect 7436 -5896 7488 -5844
rect 7488 -5896 7491 -5844
rect 7435 -5897 7491 -5896
rect 9826 -5855 9882 -5852
rect 9826 -5907 9827 -5855
rect 9827 -5907 9879 -5855
rect 9879 -5907 9882 -5855
rect 9826 -5908 9882 -5907
rect 2759 -6009 2815 -6006
rect 2759 -6061 2760 -6009
rect 2760 -6061 2812 -6009
rect 2812 -6061 2815 -6009
rect 2759 -6062 2815 -6061
rect 6250 -6000 6306 -5997
rect 6250 -6052 6251 -6000
rect 6251 -6052 6303 -6000
rect 6303 -6052 6306 -6000
rect 6250 -6053 6306 -6052
rect 7426 -6061 7482 -6058
rect 7426 -6113 7427 -6061
rect 7427 -6113 7479 -6061
rect 7479 -6113 7482 -6061
rect 7426 -6114 7482 -6113
rect 9825 -6036 9881 -6033
rect 9825 -6088 9826 -6036
rect 9826 -6088 9878 -6036
rect 9878 -6088 9881 -6036
rect 9825 -6089 9881 -6088
rect 928 -6937 984 -6934
rect 928 -6989 929 -6937
rect 929 -6989 981 -6937
rect 981 -6989 984 -6937
rect 928 -6990 984 -6989
rect 1147 -6940 1203 -6937
rect 1147 -6992 1148 -6940
rect 1148 -6992 1200 -6940
rect 1200 -6992 1203 -6940
rect 1147 -6993 1203 -6992
rect 11418 -7242 11474 -7240
rect 11418 -7294 11420 -7242
rect 11420 -7294 11472 -7242
rect 11472 -7294 11474 -7242
rect 11418 -7296 11474 -7294
rect 23380 -4954 23436 -4951
rect 23380 -5006 23381 -4954
rect 23381 -5006 23433 -4954
rect 23433 -5006 23436 -4954
rect 23380 -5007 23436 -5006
rect 23602 -4946 23658 -4943
rect 23602 -4998 23603 -4946
rect 23603 -4998 23655 -4946
rect 23655 -4998 23658 -4946
rect 23602 -4999 23658 -4998
rect 26717 -5997 26773 -5994
rect 26717 -6049 26718 -5997
rect 26718 -6049 26770 -5997
rect 26770 -6049 26773 -5997
rect 26717 -6050 26773 -6049
rect 27058 -5999 27114 -5996
rect 27058 -6051 27059 -5999
rect 27059 -6051 27111 -5999
rect 27111 -6051 27114 -5999
rect 27058 -6052 27114 -6051
rect 3784 -7763 3840 -7760
rect 3784 -7815 3785 -7763
rect 3785 -7815 3837 -7763
rect 3837 -7815 3840 -7763
rect 3784 -7816 3840 -7815
rect 6222 -7781 6278 -7778
rect 6222 -7833 6274 -7781
rect 6274 -7833 6278 -7781
rect 6222 -7834 6278 -7833
rect 9700 -7783 9756 -7780
rect 9700 -7835 9701 -7783
rect 9701 -7835 9753 -7783
rect 9753 -7835 9756 -7783
rect 9700 -7836 9756 -7835
rect 10943 -7785 10999 -7782
rect 10943 -7837 10944 -7785
rect 10944 -7837 10996 -7785
rect 10996 -7837 10999 -7785
rect 10943 -7838 10999 -7837
rect 13398 -7808 13454 -7805
rect 13398 -7860 13399 -7808
rect 13399 -7860 13451 -7808
rect 13451 -7860 13454 -7808
rect 13398 -7861 13454 -7860
rect 3779 -7945 3835 -7942
rect 3779 -7997 3780 -7945
rect 3780 -7997 3832 -7945
rect 3832 -7997 3835 -7945
rect 3779 -7998 3835 -7997
rect 6223 -7932 6279 -7930
rect 6223 -7984 6225 -7932
rect 6225 -7984 6277 -7932
rect 6277 -7984 6279 -7932
rect 6223 -7986 6279 -7984
rect 9704 -7948 9760 -7945
rect 9704 -8000 9705 -7948
rect 9705 -8000 9757 -7948
rect 9757 -8000 9760 -7948
rect 9704 -8001 9760 -8000
rect 10941 -8003 10997 -8000
rect 10941 -8055 10942 -8003
rect 10942 -8055 10994 -8003
rect 10994 -8055 10997 -8003
rect 10941 -8056 10997 -8055
rect 13396 -8023 13452 -8020
rect 13396 -8075 13397 -8023
rect 13397 -8075 13449 -8023
rect 13449 -8075 13452 -8023
rect 13396 -8076 13452 -8075
rect 318 -8116 374 -8113
rect 318 -8168 319 -8116
rect 319 -8168 371 -8116
rect 371 -8168 374 -8116
rect 318 -8169 374 -8168
rect 501 -8115 557 -8112
rect 501 -8167 502 -8115
rect 502 -8167 554 -8115
rect 554 -8167 557 -8115
rect 501 -8168 557 -8167
rect 2904 -8879 2960 -8823
rect 3151 -8879 3207 -8823
rect 645 -8928 701 -8925
rect 645 -8980 646 -8928
rect 646 -8980 698 -8928
rect 698 -8980 701 -8928
rect 645 -8981 701 -8980
rect 922 -8927 978 -8924
rect 922 -8979 923 -8927
rect 923 -8979 975 -8927
rect 975 -8979 978 -8927
rect 922 -8980 978 -8979
rect 2010 -9248 2066 -9246
rect 1859 -9254 1915 -9252
rect 1732 -9257 1788 -9255
rect 1615 -9259 1671 -9257
rect 1500 -9264 1556 -9262
rect 1500 -9316 1502 -9264
rect 1502 -9316 1554 -9264
rect 1554 -9316 1556 -9264
rect 1615 -9311 1617 -9259
rect 1617 -9311 1669 -9259
rect 1669 -9311 1671 -9259
rect 1732 -9309 1734 -9257
rect 1734 -9309 1786 -9257
rect 1786 -9309 1788 -9257
rect 1859 -9306 1861 -9254
rect 1861 -9306 1913 -9254
rect 1913 -9306 1915 -9254
rect 2010 -9300 2012 -9248
rect 2012 -9300 2064 -9248
rect 2064 -9300 2066 -9248
rect 2010 -9302 2066 -9300
rect 1859 -9308 1915 -9306
rect 1732 -9311 1788 -9309
rect 1615 -9313 1671 -9311
rect 1500 -9318 1556 -9316
rect 1627 -9382 1683 -9380
rect 1512 -9384 1568 -9382
rect 1512 -9436 1514 -9384
rect 1514 -9436 1566 -9384
rect 1566 -9436 1568 -9384
rect 1627 -9434 1629 -9382
rect 1629 -9434 1681 -9382
rect 1681 -9434 1683 -9382
rect 1627 -9436 1683 -9434
rect 1770 -9384 1826 -9382
rect 1770 -9436 1772 -9384
rect 1772 -9436 1824 -9384
rect 1824 -9436 1826 -9384
rect 1512 -9438 1568 -9436
rect 1770 -9438 1826 -9436
rect 1900 -9384 1956 -9382
rect 1900 -9436 1902 -9384
rect 1902 -9436 1954 -9384
rect 1954 -9436 1956 -9384
rect 1900 -9438 1956 -9436
rect 2024 -9386 2080 -9384
rect 2024 -9438 2026 -9386
rect 2026 -9438 2078 -9386
rect 2078 -9438 2080 -9386
rect 2024 -9440 2080 -9438
rect 11424 -9459 11480 -9457
rect 11282 -9465 11338 -9463
rect 11158 -9468 11214 -9466
rect 11158 -9520 11160 -9468
rect 11160 -9520 11212 -9468
rect 11212 -9520 11214 -9468
rect 11282 -9517 11284 -9465
rect 11284 -9517 11336 -9465
rect 11336 -9517 11338 -9465
rect 11424 -9511 11426 -9459
rect 11426 -9511 11478 -9459
rect 11478 -9511 11480 -9459
rect 11424 -9513 11480 -9511
rect 11568 -9461 11624 -9459
rect 11568 -9513 11570 -9461
rect 11570 -9513 11622 -9461
rect 11622 -9513 11624 -9461
rect 11568 -9515 11624 -9513
rect 11282 -9519 11338 -9517
rect 11158 -9522 11214 -9520
rect 11421 -9576 11477 -9574
rect 11281 -9578 11337 -9576
rect 11154 -9583 11210 -9581
rect 11154 -9635 11156 -9583
rect 11156 -9635 11208 -9583
rect 11208 -9635 11210 -9583
rect 11281 -9630 11283 -9578
rect 11283 -9630 11335 -9578
rect 11335 -9630 11337 -9578
rect 11421 -9628 11423 -9576
rect 11423 -9628 11475 -9576
rect 11475 -9628 11477 -9576
rect 11421 -9630 11477 -9628
rect 11562 -9580 11618 -9578
rect 11281 -9632 11337 -9630
rect 11562 -9632 11564 -9580
rect 11564 -9632 11616 -9580
rect 11616 -9632 11618 -9580
rect 11562 -9634 11618 -9632
rect 11154 -9637 11210 -9635
rect 19637 -9452 19693 -9450
rect 19495 -9458 19551 -9456
rect 19371 -9461 19427 -9459
rect 19371 -9513 19373 -9461
rect 19373 -9513 19425 -9461
rect 19425 -9513 19427 -9461
rect 19495 -9510 19497 -9458
rect 19497 -9510 19549 -9458
rect 19549 -9510 19551 -9458
rect 19637 -9504 19639 -9452
rect 19639 -9504 19691 -9452
rect 19691 -9504 19693 -9452
rect 19637 -9506 19693 -9504
rect 19781 -9454 19837 -9452
rect 19781 -9506 19783 -9454
rect 19783 -9506 19835 -9454
rect 19835 -9506 19837 -9454
rect 19781 -9508 19837 -9506
rect 19495 -9512 19551 -9510
rect 19371 -9515 19427 -9513
rect 19634 -9569 19690 -9567
rect 19494 -9571 19550 -9569
rect 19367 -9576 19423 -9574
rect 19367 -9628 19369 -9576
rect 19369 -9628 19421 -9576
rect 19421 -9628 19423 -9576
rect 19494 -9623 19496 -9571
rect 19496 -9623 19548 -9571
rect 19548 -9623 19550 -9571
rect 19634 -9621 19636 -9569
rect 19636 -9621 19688 -9569
rect 19688 -9621 19690 -9569
rect 19634 -9623 19690 -9621
rect 19775 -9573 19831 -9571
rect 19494 -9625 19550 -9623
rect 19775 -9625 19777 -9573
rect 19777 -9625 19829 -9573
rect 19829 -9625 19831 -9573
rect 19775 -9627 19831 -9625
rect 19367 -9630 19423 -9628
rect 26699 -9433 26755 -9431
rect 26557 -9439 26613 -9437
rect 26433 -9442 26489 -9440
rect 26433 -9494 26435 -9442
rect 26435 -9494 26487 -9442
rect 26487 -9494 26489 -9442
rect 26557 -9491 26559 -9439
rect 26559 -9491 26611 -9439
rect 26611 -9491 26613 -9439
rect 26699 -9485 26701 -9433
rect 26701 -9485 26753 -9433
rect 26753 -9485 26755 -9433
rect 26699 -9487 26755 -9485
rect 26843 -9435 26899 -9433
rect 26843 -9487 26845 -9435
rect 26845 -9487 26897 -9435
rect 26897 -9487 26899 -9435
rect 26843 -9489 26899 -9487
rect 26557 -9493 26613 -9491
rect 26433 -9496 26489 -9494
rect 26696 -9550 26752 -9548
rect 26556 -9552 26612 -9550
rect 26429 -9557 26485 -9555
rect 26429 -9609 26431 -9557
rect 26431 -9609 26483 -9557
rect 26483 -9609 26485 -9557
rect 26556 -9604 26558 -9552
rect 26558 -9604 26610 -9552
rect 26610 -9604 26612 -9552
rect 26696 -9602 26698 -9550
rect 26698 -9602 26750 -9550
rect 26750 -9602 26752 -9550
rect 26696 -9604 26752 -9602
rect 26837 -9554 26893 -9552
rect 26556 -9606 26612 -9604
rect 26837 -9606 26839 -9554
rect 26839 -9606 26891 -9554
rect 26891 -9606 26893 -9554
rect 26837 -9608 26893 -9606
rect 26429 -9611 26485 -9609
rect 33504 -9431 33560 -9429
rect 33362 -9437 33418 -9435
rect 33238 -9440 33294 -9438
rect 33238 -9492 33240 -9440
rect 33240 -9492 33292 -9440
rect 33292 -9492 33294 -9440
rect 33362 -9489 33364 -9437
rect 33364 -9489 33416 -9437
rect 33416 -9489 33418 -9437
rect 33504 -9483 33506 -9431
rect 33506 -9483 33558 -9431
rect 33558 -9483 33560 -9431
rect 33504 -9485 33560 -9483
rect 33648 -9433 33704 -9431
rect 33648 -9485 33650 -9433
rect 33650 -9485 33702 -9433
rect 33702 -9485 33704 -9433
rect 33648 -9487 33704 -9485
rect 33362 -9491 33418 -9489
rect 33238 -9494 33294 -9492
rect 33501 -9548 33557 -9546
rect 33361 -9550 33417 -9548
rect 33234 -9555 33290 -9553
rect 33234 -9607 33236 -9555
rect 33236 -9607 33288 -9555
rect 33288 -9607 33290 -9555
rect 33361 -9602 33363 -9550
rect 33363 -9602 33415 -9550
rect 33415 -9602 33417 -9550
rect 33501 -9600 33503 -9548
rect 33503 -9600 33555 -9548
rect 33555 -9600 33557 -9548
rect 33501 -9602 33557 -9600
rect 33642 -9552 33698 -9550
rect 33361 -9604 33417 -9602
rect 33642 -9604 33644 -9552
rect 33644 -9604 33696 -9552
rect 33696 -9604 33698 -9552
rect 33642 -9606 33698 -9604
rect 33234 -9609 33290 -9607
rect 15396 -9882 15452 -9880
rect 15254 -9888 15310 -9886
rect 5510 -9964 5566 -9962
rect 5368 -9970 5424 -9968
rect 5244 -9973 5300 -9971
rect 5244 -10025 5246 -9973
rect 5246 -10025 5298 -9973
rect 5298 -10025 5300 -9973
rect 5368 -10022 5370 -9970
rect 5370 -10022 5422 -9970
rect 5422 -10022 5424 -9970
rect 5510 -10016 5512 -9964
rect 5512 -10016 5564 -9964
rect 5564 -10016 5566 -9964
rect 5510 -10018 5566 -10016
rect 5654 -9966 5710 -9964
rect 5654 -10018 5656 -9966
rect 5656 -10018 5708 -9966
rect 5708 -10018 5710 -9966
rect 5654 -10020 5710 -10018
rect 5368 -10024 5424 -10022
rect 5244 -10027 5300 -10025
rect 15130 -9891 15186 -9889
rect 15130 -9943 15132 -9891
rect 15132 -9943 15184 -9891
rect 15184 -9943 15186 -9891
rect 15254 -9940 15256 -9888
rect 15256 -9940 15308 -9888
rect 15308 -9940 15310 -9888
rect 15396 -9934 15398 -9882
rect 15398 -9934 15450 -9882
rect 15450 -9934 15452 -9882
rect 15396 -9936 15452 -9934
rect 15540 -9884 15596 -9882
rect 15540 -9936 15542 -9884
rect 15542 -9936 15594 -9884
rect 15594 -9936 15596 -9884
rect 15540 -9938 15596 -9936
rect 15254 -9942 15310 -9940
rect 15130 -9945 15186 -9943
rect 15393 -9999 15449 -9997
rect 15253 -10001 15309 -9999
rect 15126 -10006 15182 -10004
rect 15126 -10058 15128 -10006
rect 15128 -10058 15180 -10006
rect 15180 -10058 15182 -10006
rect 15253 -10053 15255 -10001
rect 15255 -10053 15307 -10001
rect 15307 -10053 15309 -10001
rect 15393 -10051 15395 -9999
rect 15395 -10051 15447 -9999
rect 15447 -10051 15449 -9999
rect 15393 -10053 15449 -10051
rect 15534 -10003 15590 -10001
rect 15253 -10055 15309 -10053
rect 15534 -10055 15536 -10003
rect 15536 -10055 15588 -10003
rect 15588 -10055 15590 -10003
rect 15534 -10057 15590 -10055
rect 22927 -9852 22983 -9850
rect 22785 -9858 22841 -9856
rect 22661 -9861 22717 -9859
rect 22661 -9913 22663 -9861
rect 22663 -9913 22715 -9861
rect 22715 -9913 22717 -9861
rect 22785 -9910 22787 -9858
rect 22787 -9910 22839 -9858
rect 22839 -9910 22841 -9858
rect 22927 -9904 22929 -9852
rect 22929 -9904 22981 -9852
rect 22981 -9904 22983 -9852
rect 22927 -9906 22983 -9904
rect 23071 -9854 23127 -9852
rect 23071 -9906 23073 -9854
rect 23073 -9906 23125 -9854
rect 23125 -9906 23127 -9854
rect 23071 -9908 23127 -9906
rect 22785 -9912 22841 -9910
rect 22661 -9915 22717 -9913
rect 22924 -9969 22980 -9967
rect 22784 -9971 22840 -9969
rect 22657 -9976 22713 -9974
rect 22657 -10028 22659 -9976
rect 22659 -10028 22711 -9976
rect 22711 -10028 22713 -9976
rect 22784 -10023 22786 -9971
rect 22786 -10023 22838 -9971
rect 22838 -10023 22840 -9971
rect 22924 -10021 22926 -9969
rect 22926 -10021 22978 -9969
rect 22978 -10021 22980 -9969
rect 22924 -10023 22980 -10021
rect 23065 -9973 23121 -9971
rect 22784 -10025 22840 -10023
rect 23065 -10025 23067 -9973
rect 23067 -10025 23119 -9973
rect 23119 -10025 23121 -9973
rect 23065 -10027 23121 -10025
rect 22657 -10030 22713 -10028
rect 15126 -10060 15182 -10058
rect 5507 -10081 5563 -10079
rect 5367 -10083 5423 -10081
rect 5240 -10088 5296 -10086
rect 5240 -10140 5242 -10088
rect 5242 -10140 5294 -10088
rect 5294 -10140 5296 -10088
rect 5367 -10135 5369 -10083
rect 5369 -10135 5421 -10083
rect 5421 -10135 5423 -10083
rect 5507 -10133 5509 -10081
rect 5509 -10133 5561 -10081
rect 5561 -10133 5563 -10081
rect 5507 -10135 5563 -10133
rect 5648 -10085 5704 -10083
rect 5367 -10137 5423 -10135
rect 5648 -10137 5650 -10085
rect 5650 -10137 5702 -10085
rect 5702 -10137 5704 -10085
rect 5648 -10139 5704 -10137
rect 5240 -10142 5296 -10140
<< metal3 >>
rect -341 2215 -129 12493
rect 996 8777 1221 12749
rect 4967 11967 5533 12006
rect 4967 11961 5263 11967
rect 4967 11958 5121 11961
rect 4967 11902 4997 11958
rect 5053 11905 5121 11958
rect 5177 11911 5263 11961
rect 5319 11965 5533 11967
rect 5319 11911 5407 11965
rect 5177 11909 5407 11911
rect 5463 11909 5533 11965
rect 5177 11905 5533 11909
rect 5053 11902 5533 11905
rect 4967 11850 5533 11902
rect 4967 11848 5260 11850
rect 4967 11843 5120 11848
rect 4967 11787 4993 11843
rect 5049 11792 5120 11843
rect 5176 11794 5260 11848
rect 5316 11846 5533 11850
rect 5316 11794 5401 11846
rect 5176 11792 5401 11794
rect 5049 11790 5401 11792
rect 5457 11790 5533 11846
rect 5049 11787 5533 11790
rect 4967 11768 5533 11787
rect 1604 11633 2170 11672
rect 1604 11627 1900 11633
rect 1604 11624 1758 11627
rect 1604 11568 1634 11624
rect 1690 11571 1758 11624
rect 1814 11577 1900 11627
rect 1956 11631 2170 11633
rect 1956 11577 2044 11631
rect 1814 11575 2044 11577
rect 2100 11575 2170 11631
rect 1814 11571 2170 11575
rect 1690 11568 2170 11571
rect 1604 11516 2170 11568
rect 1604 11514 1897 11516
rect 1604 11509 1757 11514
rect 1604 11453 1630 11509
rect 1686 11458 1757 11509
rect 1813 11460 1897 11514
rect 1953 11512 2170 11516
rect 1953 11460 2038 11512
rect 1813 11458 2038 11460
rect 1686 11456 2038 11458
rect 2094 11456 2170 11512
rect 1686 11453 2170 11456
rect 1604 11434 2170 11453
rect 5140 10572 5228 10587
rect 5140 10516 5156 10572
rect 5212 10516 5228 10572
rect 5140 10499 5228 10516
rect 1654 9575 1814 9622
rect 1654 9519 1703 9575
rect 1759 9519 1814 9575
rect 1654 9483 1814 9519
rect 996 8721 1075 8777
rect 1131 8721 1221 8777
rect 9821 8774 9960 12103
rect 9821 8726 9867 8774
rect 996 8650 1221 8721
rect 996 8594 1076 8650
rect 1132 8594 1221 8650
rect 996 8391 1221 8594
rect 9843 8718 9867 8726
rect 9923 8726 9960 8774
rect 9923 8718 9935 8726
rect 9843 8657 9935 8718
rect 9843 8601 9857 8657
rect 9913 8601 9935 8657
rect 9843 8543 9935 8601
rect 10198 8563 10369 12087
rect 22623 12083 23189 12122
rect 22623 12077 22919 12083
rect 22623 12074 22777 12077
rect 22623 12018 22653 12074
rect 22709 12021 22777 12074
rect 22833 12027 22919 12077
rect 22975 12081 23189 12083
rect 22975 12027 23063 12081
rect 22833 12025 23063 12027
rect 23119 12025 23189 12081
rect 22833 12021 23189 12025
rect 22709 12018 23189 12021
rect 15100 11957 15666 11996
rect 15100 11951 15396 11957
rect 15100 11948 15254 11951
rect 15100 11892 15130 11948
rect 15186 11895 15254 11948
rect 15310 11901 15396 11951
rect 15452 11955 15666 11957
rect 15452 11901 15540 11955
rect 15310 11899 15540 11901
rect 15596 11899 15666 11955
rect 15310 11895 15666 11899
rect 15186 11892 15666 11895
rect 15100 11840 15666 11892
rect 22623 11966 23189 12018
rect 22623 11964 22916 11966
rect 22623 11959 22776 11964
rect 22623 11903 22649 11959
rect 22705 11908 22776 11959
rect 22832 11910 22916 11964
rect 22972 11962 23189 11966
rect 22972 11910 23057 11962
rect 22832 11908 23057 11910
rect 22705 11906 23057 11908
rect 23113 11906 23189 11962
rect 22705 11903 23189 11906
rect 15100 11838 15393 11840
rect 15100 11833 15253 11838
rect 11263 11746 11829 11785
rect 15100 11777 15126 11833
rect 15182 11782 15253 11833
rect 15309 11784 15393 11838
rect 15449 11836 15666 11840
rect 15449 11784 15534 11836
rect 15309 11782 15534 11784
rect 15182 11780 15534 11782
rect 15590 11780 15666 11836
rect 15182 11777 15666 11780
rect 15100 11758 15666 11777
rect 11263 11740 11559 11746
rect 11263 11737 11417 11740
rect 11263 11681 11293 11737
rect 11349 11684 11417 11737
rect 11473 11690 11559 11740
rect 11615 11744 11829 11746
rect 11615 11690 11703 11744
rect 11473 11688 11703 11690
rect 11759 11688 11829 11744
rect 11473 11684 11829 11688
rect 11349 11681 11829 11684
rect 11263 11629 11829 11681
rect 11263 11627 11556 11629
rect 11263 11622 11416 11627
rect 11263 11566 11289 11622
rect 11345 11571 11416 11622
rect 11472 11573 11556 11627
rect 11612 11625 11829 11629
rect 11612 11573 11697 11625
rect 11472 11571 11697 11573
rect 11345 11569 11697 11571
rect 11753 11569 11829 11625
rect 11345 11566 11829 11569
rect 11263 11547 11829 11566
rect 18502 11336 18580 11888
rect 22623 11884 23189 11903
rect 18237 11326 18580 11336
rect 18237 11324 18463 11326
rect 18237 11268 18247 11324
rect 18303 11270 18463 11324
rect 18519 11270 18580 11326
rect 18303 11268 18580 11270
rect 18237 11258 18580 11268
rect 10183 8544 10411 8563
rect 10183 8488 10200 8544
rect 10256 8543 10411 8544
rect 10256 8488 10340 8543
rect 10183 8487 10340 8488
rect 10396 8487 10411 8543
rect 10183 8432 10411 8487
rect 1053 8390 1151 8391
rect 10183 8376 10205 8432
rect 10261 8376 10411 8432
rect 11490 8480 11609 8504
rect 11490 8424 11530 8480
rect 11586 8424 11609 8480
rect 11490 8396 11609 8424
rect 10183 8332 10411 8376
rect 18502 8119 18580 11258
rect 18180 8109 18580 8119
rect 18180 8108 18373 8109
rect 11721 8088 11961 8098
rect 11721 8086 11895 8088
rect 1634 8001 1794 8048
rect 1634 7945 1683 8001
rect 1739 7945 1794 8001
rect 1634 7909 1794 7945
rect 4643 7971 7219 8032
rect 11721 8030 11731 8086
rect 11787 8032 11895 8086
rect 11951 8032 11961 8088
rect 18180 8052 18190 8108
rect 18246 8053 18373 8108
rect 18429 8053 18580 8109
rect 18246 8052 18580 8053
rect 18180 8041 18580 8052
rect 11787 8030 11961 8032
rect 11721 8020 11961 8030
rect 4643 5693 4704 7971
rect 7158 7580 7219 7971
rect 10271 7901 10607 7903
rect 10271 7848 10872 7901
rect 10271 7792 10299 7848
rect 10355 7792 10469 7848
rect 10525 7792 10872 7848
rect 11475 7899 11594 7923
rect 11475 7843 11515 7899
rect 11571 7843 11594 7899
rect 11475 7815 11594 7843
rect 10271 7743 10872 7792
rect 10271 7741 10607 7743
rect 7158 7519 8004 7580
rect 7943 7151 8004 7519
rect 7931 7141 8009 7151
rect 7931 7085 7942 7141
rect 7998 7085 8009 7141
rect 7931 7075 8009 7085
rect 7943 7005 8004 7075
rect 7938 6995 8016 7005
rect 7938 6939 7949 6995
rect 8005 6939 8016 6995
rect 7938 6929 8016 6939
rect 10714 6057 10872 7743
rect 9804 5899 10872 6057
rect 4643 5632 7225 5693
rect 5131 5350 5219 5364
rect 5131 5294 5151 5350
rect 5207 5294 5219 5350
rect 5131 5276 5219 5294
rect 7164 3174 7225 5632
rect 9804 3686 9962 5899
rect 9804 3435 9963 3686
rect 9804 3379 9855 3435
rect 9911 3379 9963 3435
rect 9804 3322 9963 3379
rect 9804 3266 9854 3322
rect 9910 3266 9963 3322
rect 9804 3235 9963 3266
rect 11725 3242 11794 8020
rect 18782 7799 18937 11882
rect 19128 11710 19694 11749
rect 19128 11704 19424 11710
rect 19128 11701 19282 11704
rect 19128 11645 19158 11701
rect 19214 11648 19282 11701
rect 19338 11654 19424 11704
rect 19480 11708 19694 11710
rect 19480 11654 19568 11708
rect 19338 11652 19568 11654
rect 19624 11652 19694 11708
rect 19338 11648 19694 11652
rect 19214 11645 19694 11648
rect 19128 11593 19694 11645
rect 19128 11591 19421 11593
rect 19128 11586 19281 11591
rect 19128 11530 19154 11586
rect 19210 11535 19281 11586
rect 19337 11537 19421 11591
rect 19477 11589 19694 11593
rect 19477 11537 19562 11589
rect 19337 11535 19562 11537
rect 19210 11533 19562 11535
rect 19618 11533 19694 11589
rect 19210 11530 19694 11533
rect 19128 11511 19694 11530
rect 19481 8806 19600 8830
rect 19481 8750 19521 8806
rect 19577 8750 19600 8806
rect 19481 8722 19600 8750
rect 21686 8226 21766 8236
rect 21823 8226 21903 8236
rect 21686 8225 21929 8226
rect 21686 8169 21698 8225
rect 21754 8224 21929 8225
rect 21754 8169 21835 8224
rect 21686 8168 21835 8169
rect 21891 8168 21929 8224
rect 21686 8167 21929 8168
rect 21686 8159 21903 8167
rect 18618 7644 18937 7799
rect 21697 8158 21903 8159
rect 18618 6136 18773 7644
rect 19429 7611 19548 7635
rect 19429 7555 19469 7611
rect 19525 7555 19548 7611
rect 19429 7527 19548 7555
rect 18585 6058 18796 6136
rect 18585 6056 18726 6058
rect 18585 6000 18603 6056
rect 18659 6002 18726 6056
rect 18782 6002 18796 6058
rect 18659 6000 18796 6002
rect 18585 5949 18796 6000
rect 18585 5942 18725 5949
rect 18585 5886 18604 5942
rect 18660 5893 18725 5942
rect 18781 5893 18796 5949
rect 18660 5886 18796 5893
rect 18585 5865 18796 5886
rect 15496 5736 15593 5762
rect 15496 5680 15519 5736
rect 15575 5680 15593 5736
rect 15496 5658 15593 5680
rect 19436 3614 19555 3638
rect 19436 3558 19476 3614
rect 19532 3558 19555 3614
rect 19436 3530 19555 3558
rect 2126 3113 7225 3174
rect 11296 3231 11806 3242
rect 11296 3226 11738 3231
rect 11296 3173 11322 3226
rect 11311 3170 11322 3173
rect 11378 3221 11738 3226
rect 11378 3173 11543 3221
rect 11378 3170 11390 3173
rect 11311 3159 11390 3170
rect 11532 3165 11543 3173
rect 11599 3175 11738 3221
rect 11794 3175 11806 3231
rect 11599 3173 11806 3175
rect 11599 3165 11611 3173
rect 11532 3154 11611 3165
rect 11727 3164 11806 3173
rect 1295 3012 1513 3024
rect 1295 2956 1424 3012
rect 1480 2956 1513 3012
rect 1295 2933 1513 2956
rect 1295 2877 1306 2933
rect 1362 2877 1513 2933
rect 1295 2874 1513 2877
rect 1295 2818 1425 2874
rect 1481 2818 1513 2874
rect 1295 2802 1513 2818
rect 1690 2805 1850 2852
rect 1363 2215 1490 2802
rect 1690 2749 1739 2805
rect 1795 2749 1850 2805
rect 1690 2713 1850 2749
rect -341 2088 1490 2215
rect -341 2045 -129 2088
rect 2126 -40 2187 3113
rect 21697 3074 21794 8158
rect 22892 5733 22976 5753
rect 22892 5677 22904 5733
rect 22960 5677 22976 5733
rect 22892 5669 22976 5677
rect 3073 3014 3151 3021
rect 3363 3014 3441 3022
rect 3054 3012 4712 3014
rect 3054 3011 3374 3012
rect 3054 2955 3084 3011
rect 3140 2956 3374 3011
rect 3430 2956 4712 3012
rect 3140 2955 4712 2956
rect 3054 2946 4712 2955
rect 3073 2945 3151 2946
rect 4644 391 4712 2946
rect 8267 2977 21794 3074
rect 25756 3021 25945 11975
rect 26109 11692 26675 11731
rect 26109 11686 26405 11692
rect 26109 11683 26263 11686
rect 26109 11627 26139 11683
rect 26195 11630 26263 11683
rect 26319 11636 26405 11686
rect 26461 11690 26675 11692
rect 26461 11636 26549 11690
rect 26319 11634 26549 11636
rect 26605 11634 26675 11690
rect 26319 11630 26675 11634
rect 26195 11627 26675 11630
rect 26109 11575 26675 11627
rect 26109 11573 26402 11575
rect 26109 11568 26262 11573
rect 26109 11512 26135 11568
rect 26191 11517 26262 11568
rect 26318 11519 26402 11573
rect 26458 11571 26675 11575
rect 26458 11519 26543 11571
rect 26318 11517 26543 11519
rect 26191 11515 26543 11517
rect 26599 11515 26675 11571
rect 26191 11512 26675 11515
rect 26109 11493 26675 11512
rect 26519 8417 26679 8472
rect 26519 8361 26568 8417
rect 26624 8361 26679 8417
rect 26519 8325 26679 8361
rect 29862 6993 30093 11969
rect 32982 11764 33548 11803
rect 32982 11758 33278 11764
rect 32982 11755 33136 11758
rect 32982 11699 33012 11755
rect 33068 11702 33136 11755
rect 33192 11708 33278 11758
rect 33334 11762 33548 11764
rect 33334 11708 33422 11762
rect 33192 11706 33422 11708
rect 33478 11706 33548 11762
rect 33192 11702 33548 11706
rect 33068 11699 33548 11702
rect 32982 11647 33548 11699
rect 32982 11645 33275 11647
rect 32982 11640 33135 11645
rect 32982 11584 33008 11640
rect 33064 11589 33135 11640
rect 33191 11591 33275 11645
rect 33331 11643 33548 11647
rect 33331 11591 33416 11643
rect 33191 11589 33416 11591
rect 33064 11587 33416 11589
rect 33472 11587 33548 11643
rect 33064 11584 33548 11587
rect 32982 11565 33548 11584
rect 25756 3004 26304 3021
rect 25756 3000 26136 3004
rect 7651 395 7730 404
rect 7806 395 7885 405
rect 6033 394 7885 395
rect 6033 393 7817 394
rect 4644 323 5941 391
rect 4500 125 4561 185
rect 4500 115 4578 125
rect 4500 59 4511 115
rect 4567 59 4578 115
rect 4500 49 4578 59
rect 2126 -133 2203 -40
rect 2356 -51 2434 -41
rect 2356 -61 2367 -51
rect 2354 -107 2367 -61
rect 2423 -61 2434 -51
rect 2423 -104 2601 -61
rect 2967 -70 3045 -63
rect 3171 -70 3249 -65
rect 2725 -73 3331 -70
rect 2423 -107 2621 -104
rect 2354 -114 2621 -107
rect 2354 -127 2554 -114
rect 522 -188 600 -180
rect -82 -190 600 -188
rect -82 -245 533 -190
rect -82 -4962 -25 -245
rect 475 -246 533 -245
rect 589 -246 600 -190
rect 475 -247 600 -246
rect 522 -256 600 -247
rect 906 -229 1417 -218
rect 527 -347 593 -256
rect 906 -285 1196 -229
rect 1252 -230 1417 -229
rect 1252 -285 1348 -230
rect 906 -286 1348 -285
rect 1404 -286 1417 -230
rect 906 -298 1417 -286
rect 518 -357 596 -347
rect 518 -413 529 -357
rect 585 -413 596 -357
rect 518 -423 596 -413
rect 906 -531 986 -298
rect 325 -611 986 -531
rect 325 -1334 405 -611
rect 316 -1345 405 -1334
rect 316 -1401 327 -1345
rect 383 -1401 405 -1345
rect 316 -1412 405 -1401
rect 325 -1518 405 -1412
rect 323 -1529 405 -1518
rect 323 -1585 334 -1529
rect 390 -1585 405 -1529
rect 323 -1596 405 -1585
rect 325 -2268 405 -1596
rect 309 -2316 405 -2268
rect 309 -4658 368 -2316
rect 1726 -2428 1886 -2381
rect 1726 -2484 1775 -2428
rect 1831 -2484 1886 -2428
rect 1726 -2520 1886 -2484
rect 2144 -2580 2203 -133
rect 2535 -170 2554 -127
rect 2610 -170 2621 -114
rect 2535 -180 2621 -170
rect 2725 -129 2978 -73
rect 3034 -75 3331 -73
rect 3034 -129 3182 -75
rect 2725 -131 3182 -129
rect 3238 -131 3331 -75
rect 2725 -135 3331 -131
rect 2535 -1761 2601 -180
rect 2725 -1428 2790 -135
rect 2967 -139 3045 -135
rect 3171 -141 3249 -135
rect 3805 -363 4215 -359
rect 3805 -373 4217 -363
rect 3805 -377 4150 -373
rect 3805 -433 3927 -377
rect 3983 -429 4150 -377
rect 4206 -429 4217 -373
rect 3983 -433 4217 -429
rect 3805 -439 4217 -433
rect 3805 -451 4215 -439
rect 3805 -1206 3897 -451
rect 3805 -1262 3823 -1206
rect 3879 -1262 3897 -1206
rect 2723 -1439 2802 -1428
rect 2723 -1495 2734 -1439
rect 2790 -1495 2802 -1439
rect 2723 -1506 2802 -1495
rect 2725 -1511 2790 -1506
rect 3805 -1512 3897 -1262
rect 3805 -1568 3819 -1512
rect 3875 -1568 3897 -1512
rect 3805 -1591 3897 -1568
rect 2535 -1827 4428 -1761
rect 496 -2639 2203 -2580
rect 496 -3274 555 -2639
rect 487 -3285 566 -3274
rect 487 -3341 498 -3285
rect 554 -3341 566 -3285
rect 487 -3352 566 -3341
rect 496 -3483 555 -3352
rect 483 -3494 562 -3483
rect 483 -3550 494 -3494
rect 550 -3550 562 -3494
rect 483 -3561 562 -3550
rect 496 -4366 555 -3561
rect 3511 -4301 3577 -1827
rect 4362 -2375 4428 -1827
rect 4344 -2385 4428 -2375
rect 4344 -2441 4355 -2385
rect 4411 -2441 4428 -2385
rect 4344 -2451 4428 -2441
rect 4362 -2464 4428 -2451
rect 3796 -2568 3875 -2557
rect 3796 -2573 3807 -2568
rect 765 -4365 844 -4354
rect 765 -4366 776 -4365
rect 496 -4421 776 -4366
rect 832 -4366 844 -4365
rect 964 -4366 1043 -4355
rect 832 -4421 975 -4366
rect 496 -4422 975 -4421
rect 1031 -4422 1043 -4366
rect 496 -4425 1043 -4422
rect 765 -4432 844 -4425
rect 964 -4433 1043 -4425
rect 2831 -4367 3577 -4301
rect 305 -4669 384 -4658
rect 305 -4725 316 -4669
rect 372 -4725 384 -4669
rect 305 -4736 384 -4725
rect 309 -4815 368 -4736
rect 303 -4826 382 -4815
rect 303 -4882 314 -4826
rect 370 -4882 382 -4826
rect 2361 -4836 2440 -4825
rect 2361 -4840 2372 -4836
rect 303 -4893 382 -4882
rect 2352 -4892 2372 -4840
rect 2428 -4840 2440 -4836
rect 2603 -4834 2682 -4823
rect 2603 -4840 2614 -4834
rect 2428 -4890 2614 -4840
rect 2670 -4840 2682 -4834
rect 2831 -4840 2897 -4367
rect 3511 -4370 3577 -4367
rect 3783 -2624 3807 -2573
rect 3863 -2573 3875 -2568
rect 4056 -2570 4135 -2559
rect 4056 -2573 4067 -2570
rect 3863 -2624 4067 -2573
rect 3783 -2626 4067 -2624
rect 4123 -2573 4135 -2570
rect 4502 -2573 4561 49
rect 4123 -2626 4561 -2573
rect 3783 -2632 4561 -2626
rect 3783 -2635 3875 -2632
rect 3783 -4334 3842 -2635
rect 4056 -2637 4135 -2632
rect 5554 -4200 5648 -4184
rect 5554 -4256 5576 -4200
rect 5632 -4256 5648 -4200
rect 5554 -4267 5648 -4256
rect 3783 -4393 5779 -4334
rect 3612 -4515 3691 -4509
rect 2980 -4520 4915 -4515
rect 2980 -4526 3623 -4520
rect 2980 -4581 3289 -4526
rect 3278 -4582 3289 -4581
rect 3345 -4576 3623 -4526
rect 3679 -4576 4915 -4520
rect 3345 -4581 4915 -4576
rect 3345 -4582 3357 -4581
rect 3278 -4593 3357 -4582
rect 3612 -4587 3691 -4581
rect 2670 -4890 2897 -4840
rect 2428 -4892 2897 -4890
rect 2352 -4906 2897 -4892
rect -82 -5019 3750 -4962
rect -88 -5209 -9 -5207
rect -103 -5218 -9 -5209
rect -103 -5274 -77 -5218
rect -21 -5274 -9 -5218
rect -103 -5285 -9 -5274
rect -103 -5397 -11 -5285
rect -103 -5453 -85 -5397
rect -29 -5453 -11 -5397
rect -103 -8091 -11 -5453
rect 3693 -5465 3750 -5019
rect 3677 -5476 3756 -5465
rect 3677 -5532 3688 -5476
rect 3744 -5532 3756 -5476
rect 3677 -5543 3756 -5532
rect 2751 -5756 4475 -5690
rect 2751 -5822 2817 -5756
rect 2750 -5833 2829 -5822
rect 2750 -5889 2761 -5833
rect 2817 -5889 2829 -5833
rect 2750 -5900 2829 -5889
rect 2751 -5995 2817 -5900
rect 2748 -6006 2827 -5995
rect 2748 -6062 2759 -6006
rect 2815 -6062 2827 -6006
rect 2748 -6073 2827 -6062
rect 2751 -6093 2817 -6073
rect 4409 -6281 4475 -5756
rect 4849 -5857 4915 -4581
rect 4849 -5923 5624 -5857
rect 5558 -6281 5624 -5923
rect 4409 -6347 5624 -6281
rect 5720 -6711 5779 -4393
rect 5873 -4549 5941 323
rect 6033 337 7662 393
rect 7718 338 7817 393
rect 7873 338 7885 394
rect 7718 337 7885 338
rect 6033 335 7885 337
rect 6033 27 6093 335
rect 7651 326 7730 335
rect 7806 327 7885 335
rect 6025 16 6104 27
rect 6025 -40 6036 16
rect 6092 -40 6104 16
rect 6247 -21 6574 -19
rect 6025 -51 6104 -40
rect 6221 -30 6574 -21
rect 6221 -31 6495 -30
rect 6033 -353 6093 -51
rect 6221 -87 6301 -31
rect 6357 -86 6495 -31
rect 6551 -86 6574 -30
rect 6357 -87 6574 -86
rect 6221 -108 6574 -87
rect 6033 -364 6112 -353
rect 6033 -420 6044 -364
rect 6100 -420 6112 -364
rect 6033 -431 6112 -420
rect 6033 -2263 6093 -431
rect 6221 -1248 6280 -108
rect 8267 -360 8364 2977
rect 25756 2955 25831 3000
rect 25807 2944 25831 2955
rect 25887 2944 25979 3000
rect 26035 2948 26136 3000
rect 26192 2948 26304 3004
rect 26035 2944 26304 2948
rect 25807 2929 26304 2944
rect 9964 2882 10911 2894
rect 9964 2881 10333 2882
rect 9964 2825 10095 2881
rect 10151 2826 10333 2881
rect 10389 2826 10911 2882
rect 10151 2825 10911 2826
rect 9964 2812 10911 2825
rect 10829 -232 10911 2812
rect 11456 2719 11575 2743
rect 11456 2663 11496 2719
rect 11552 2663 11575 2719
rect 11456 2635 11575 2663
rect 26416 2689 26576 2744
rect 26416 2633 26465 2689
rect 26521 2633 26576 2689
rect 26416 2597 26576 2633
rect 11023 2318 11102 2329
rect 11023 2262 11034 2318
rect 11090 2262 11102 2318
rect 11023 2251 11102 2262
rect 11032 2194 11094 2251
rect 11028 2190 11107 2194
rect 7393 -457 8364 -360
rect 9639 -314 10911 -232
rect 10992 2183 11107 2190
rect 10992 2127 11039 2183
rect 11095 2127 11107 2183
rect 10992 2116 11107 2127
rect 7393 -1191 7490 -457
rect 9639 -499 9721 -314
rect 10992 -403 11054 2116
rect 15199 519 15283 533
rect 15199 463 15215 519
rect 15271 463 15283 519
rect 15199 447 15283 463
rect 11526 385 22753 387
rect 11526 376 22758 385
rect 11526 320 22515 376
rect 22571 374 22758 376
rect 22571 320 22690 374
rect 11526 318 22690 320
rect 22746 318 22758 374
rect 11526 308 22758 318
rect 23071 344 23128 2350
rect 31692 2011 31786 2029
rect 31692 2001 31710 2011
rect 30395 1955 31710 2001
rect 31766 2001 31786 2011
rect 31766 1955 31792 2001
rect 30395 1924 31792 1955
rect 29168 1923 31792 1924
rect 28898 1909 31792 1923
rect 28898 1893 30487 1909
rect 28898 1837 28948 1893
rect 29004 1892 30487 1893
rect 29004 1837 29231 1892
rect 28898 1836 29231 1837
rect 29287 1836 30487 1892
rect 28898 1832 30487 1836
rect 28898 1821 29204 1832
rect 11526 302 22753 308
rect 11526 198 11611 302
rect 23071 287 23537 344
rect 11221 156 11611 198
rect 11221 152 11494 156
rect 11221 113 11260 152
rect 11249 96 11260 113
rect 11316 113 11494 152
rect 11316 96 11328 113
rect 11249 86 11328 96
rect 11483 100 11494 113
rect 11550 113 11611 156
rect 13873 114 17681 125
rect 13873 113 14138 114
rect 11550 100 11562 113
rect 11483 90 11562 100
rect 13873 57 13928 113
rect 13984 58 14138 113
rect 14194 58 17681 114
rect 13984 57 17681 58
rect 13873 45 17681 57
rect 14670 -33 14749 -22
rect 14670 -35 14681 -33
rect 9839 -465 11054 -403
rect 7393 -1202 7494 -1191
rect 6210 -1259 6289 -1248
rect 6210 -1315 6221 -1259
rect 6277 -1315 6289 -1259
rect 6210 -1326 6289 -1315
rect 7393 -1258 7426 -1202
rect 7482 -1258 7494 -1202
rect 7393 -1269 7494 -1258
rect 6221 -1417 6280 -1326
rect 6215 -1428 6294 -1417
rect 6215 -1484 6226 -1428
rect 6282 -1484 6294 -1428
rect 6215 -1495 6294 -1484
rect 7393 -1452 7490 -1269
rect 7393 -1508 7418 -1452
rect 7474 -1508 7490 -1452
rect 9646 -1436 9713 -499
rect 9845 -1219 9906 -465
rect 9835 -1230 9914 -1219
rect 9835 -1286 9846 -1230
rect 9902 -1286 9914 -1230
rect 9835 -1297 9914 -1286
rect 9646 -1503 10022 -1436
rect 7393 -1519 7490 -1508
rect 7413 -1831 7472 -1519
rect 7413 -1890 8328 -1831
rect 6033 -2323 7350 -2263
rect 7287 -2957 7347 -2323
rect 7280 -2968 7359 -2957
rect 7280 -3024 7291 -2968
rect 7347 -3024 7359 -2968
rect 7280 -3035 7359 -3024
rect 7287 -3317 7347 -3035
rect 8269 -3066 8328 -1890
rect 9955 -2528 10022 -1503
rect 9697 -2530 10022 -2528
rect 9695 -2540 10022 -2530
rect 9695 -2596 9706 -2540
rect 9762 -2596 9898 -2540
rect 9954 -2596 10022 -2540
rect 9695 -2604 10022 -2596
rect 9695 -2606 9773 -2604
rect 9887 -2606 9965 -2604
rect 8266 -3125 10094 -3066
rect 7264 -3328 7347 -3317
rect 7264 -3384 7275 -3328
rect 7331 -3384 7347 -3328
rect 7264 -3393 7347 -3384
rect 7264 -3395 7343 -3393
rect 9751 -4521 9891 -4515
rect 9546 -4531 9891 -4521
rect 9546 -4540 9810 -4531
rect 9546 -4549 9573 -4540
rect 5873 -4596 9573 -4549
rect 9629 -4587 9810 -4540
rect 9866 -4571 9891 -4531
rect 9866 -4587 9889 -4571
rect 9629 -4596 9889 -4587
rect 5873 -4617 9889 -4596
rect 5873 -6642 5941 -4617
rect 6244 -4704 9904 -4692
rect 6244 -4706 9824 -4704
rect 6244 -4762 9576 -4706
rect 9632 -4760 9824 -4706
rect 9880 -4760 9904 -4704
rect 9632 -4762 9904 -4760
rect 6244 -4767 9904 -4762
rect 6244 -5810 6318 -4767
rect 9565 -4772 9643 -4767
rect 9813 -4770 9891 -4767
rect 10035 -4991 10094 -3125
rect 10992 -4232 11054 -465
rect 14593 -89 14681 -35
rect 14737 -35 14749 -33
rect 14873 -35 14952 -26
rect 14737 -37 14952 -35
rect 14737 -89 14884 -37
rect 14593 -93 14884 -89
rect 14940 -93 14952 -37
rect 14593 -102 14952 -93
rect 14593 -1543 14660 -102
rect 14873 -103 14952 -102
rect 14593 -1585 14956 -1543
rect 14593 -1596 14969 -1585
rect 14593 -1610 14901 -1596
rect 14889 -1652 14901 -1610
rect 14957 -1652 14969 -1596
rect 14889 -1662 14969 -1652
rect 14889 -1746 14956 -1662
rect 14889 -1757 14968 -1746
rect 14889 -1813 14900 -1757
rect 14956 -1813 14968 -1757
rect 14889 -1823 14968 -1813
rect 17601 -2272 17681 45
rect 23480 3 23537 287
rect 19477 -54 23537 3
rect 19477 -149 19534 -54
rect 23480 -125 23537 -54
rect 23480 -136 23559 -125
rect 19477 -160 19559 -149
rect 19477 -216 19491 -160
rect 19547 -216 19559 -160
rect 19477 -227 19559 -216
rect 23480 -192 23490 -136
rect 23546 -192 23559 -136
rect 23480 -202 23559 -192
rect 19477 -262 19534 -227
rect 23480 -294 23537 -202
rect 23480 -305 23560 -294
rect 23480 -361 23491 -305
rect 23547 -324 23560 -305
rect 23547 -361 23726 -324
rect 23480 -381 23726 -361
rect 31762 -424 31841 -422
rect 31948 -424 32027 -420
rect 30473 -431 32035 -424
rect 30473 -433 31959 -431
rect 30473 -435 31773 -433
rect 30469 -439 31773 -435
rect 30469 -446 30677 -439
rect 30469 -502 30480 -446
rect 30536 -495 30677 -446
rect 30733 -489 31773 -439
rect 31829 -487 31959 -433
rect 32015 -487 32035 -431
rect 31829 -489 32035 -487
rect 30733 -495 32035 -489
rect 30536 -502 32035 -495
rect 30469 -511 32035 -502
rect 30469 -513 30548 -511
rect 22854 -1450 22919 -1427
rect 22854 -1506 22858 -1450
rect 22914 -1506 22919 -1450
rect 22854 -1621 22919 -1506
rect 22854 -1645 22855 -1621
rect 21857 -1648 22855 -1645
rect 21857 -1704 21886 -1648
rect 21942 -1649 22855 -1648
rect 21942 -1704 22328 -1649
rect 21857 -1705 22328 -1704
rect 22384 -1677 22855 -1649
rect 22911 -1677 22919 -1621
rect 22384 -1705 22919 -1677
rect 21857 -1710 22919 -1705
rect 17601 -2352 18532 -2272
rect 11150 -2648 16501 -2589
rect 11150 -3296 11209 -2648
rect 14749 -2717 14828 -2706
rect 14749 -2720 14760 -2717
rect 14700 -2721 14760 -2720
rect 11563 -2796 11682 -2772
rect 11563 -2852 11603 -2796
rect 11659 -2852 11682 -2796
rect 11563 -2880 11682 -2852
rect 14432 -2773 14760 -2721
rect 14816 -2720 14828 -2717
rect 14935 -2719 15014 -2708
rect 14935 -2720 14946 -2719
rect 14816 -2773 14946 -2720
rect 14432 -2775 14946 -2773
rect 15002 -2775 15014 -2719
rect 14432 -2780 15014 -2775
rect 13352 -3294 13431 -3290
rect 11118 -3307 11209 -3296
rect 11118 -3363 11129 -3307
rect 11185 -3363 11209 -3307
rect 11118 -3374 11209 -3363
rect 11150 -3689 11209 -3374
rect 13338 -3301 13436 -3294
rect 13338 -3357 13363 -3301
rect 13419 -3357 13436 -3301
rect 13338 -3462 13436 -3357
rect 13338 -3518 13359 -3462
rect 13415 -3518 13436 -3462
rect 10219 -4294 11054 -4232
rect 10219 -4947 10281 -4294
rect 13338 -4479 13436 -3518
rect 10370 -4540 13436 -4479
rect 10370 -4577 10408 -4540
rect 10397 -4596 10408 -4577
rect 10464 -4577 10655 -4540
rect 10464 -4596 10475 -4577
rect 10397 -4606 10475 -4596
rect 10644 -4596 10655 -4577
rect 10711 -4577 13436 -4540
rect 10711 -4596 10722 -4577
rect 10644 -4606 10722 -4596
rect 10407 -4693 10485 -4683
rect 10407 -4698 10418 -4693
rect 10376 -4749 10418 -4698
rect 10474 -4698 10485 -4693
rect 10656 -4689 10734 -4679
rect 10656 -4698 10667 -4689
rect 10474 -4745 10667 -4698
rect 10723 -4698 10734 -4689
rect 14432 -4698 14491 -2780
rect 14700 -2781 15014 -2780
rect 14749 -2783 14828 -2781
rect 14935 -2785 15014 -2781
rect 16442 -2806 16501 -2648
rect 17740 -2806 17799 -2805
rect 16442 -2824 18284 -2806
rect 16442 -2865 17877 -2824
rect 15441 -4186 15541 -4171
rect 15441 -4242 15464 -4186
rect 15520 -4242 15541 -4186
rect 15441 -4262 15541 -4242
rect 17740 -4280 17799 -2865
rect 17867 -2880 17877 -2865
rect 17933 -2865 18135 -2824
rect 17933 -2880 17946 -2865
rect 17867 -2890 17946 -2880
rect 18125 -2880 18135 -2865
rect 18191 -2865 18284 -2824
rect 18191 -2880 18204 -2865
rect 18125 -2890 18204 -2880
rect 18452 -2947 18532 -2352
rect 21773 -2656 21852 -2648
rect 21928 -2656 22007 -2652
rect 10723 -4745 14491 -4698
rect 10474 -4749 14491 -4745
rect 10376 -4757 14491 -4749
rect 16470 -4339 17799 -4280
rect 17884 -3021 18532 -2947
rect 21760 -2659 22229 -2656
rect 21760 -2715 21784 -2659
rect 21840 -2663 22229 -2659
rect 21840 -2715 21939 -2663
rect 21760 -2719 21939 -2715
rect 21995 -2719 22229 -2663
rect 21760 -2733 22229 -2719
rect 21760 -2999 21837 -2733
rect 10407 -4759 10485 -4757
rect 7397 -5050 10094 -4991
rect 6241 -5821 6320 -5810
rect 6241 -5877 6252 -5821
rect 6308 -5877 6320 -5821
rect 6241 -5888 6320 -5877
rect 7397 -5830 7456 -5050
rect 10218 -5134 10281 -4947
rect 9822 -5197 10281 -5134
rect 14745 -4918 14804 -4917
rect 16470 -4918 16529 -4339
rect 17884 -4437 17964 -3021
rect 18452 -3026 18532 -3021
rect 14745 -4977 16529 -4918
rect 16634 -4517 17964 -4437
rect 20975 -3076 21837 -2999
rect 7397 -5841 7503 -5830
rect 9822 -5841 9885 -5197
rect 6244 -5986 6318 -5888
rect 6239 -5997 6318 -5986
rect 6239 -6053 6250 -5997
rect 6306 -6053 6318 -5997
rect 6239 -6064 6318 -6053
rect 6244 -6086 6318 -6064
rect 7397 -5897 7435 -5841
rect 7491 -5897 7503 -5841
rect 7397 -5908 7503 -5897
rect 9815 -5852 9894 -5841
rect 9815 -5908 9826 -5852
rect 9882 -5908 9894 -5852
rect 7397 -6047 7456 -5908
rect 9815 -5919 9894 -5908
rect 9822 -6022 9885 -5919
rect 9814 -6033 9893 -6022
rect 7397 -6058 7494 -6047
rect 7397 -6114 7426 -6058
rect 7482 -6114 7494 -6058
rect 9814 -6089 9825 -6033
rect 9881 -6089 9893 -6033
rect 9814 -6100 9893 -6089
rect 7397 -6125 7494 -6114
rect 7397 -6140 7456 -6125
rect 5873 -6710 13451 -6642
rect 3779 -6770 5779 -6711
rect 916 -6934 1255 -6915
rect 916 -6990 928 -6934
rect 984 -6937 1255 -6934
rect 984 -6990 1147 -6937
rect 916 -6993 1147 -6990
rect 1203 -6993 1255 -6937
rect 916 -6995 1255 -6993
rect 917 -7001 1056 -6995
rect -103 -8112 596 -8091
rect -103 -8113 501 -8112
rect -103 -8169 318 -8113
rect 374 -8168 501 -8113
rect 557 -8168 596 -8112
rect 374 -8169 596 -8168
rect -103 -8183 596 -8169
rect 976 -8913 1056 -7001
rect 1136 -7004 1215 -6995
rect 3779 -7749 3838 -6770
rect 5720 -6784 5779 -6770
rect 11378 -7240 11497 -7216
rect 11378 -7296 11418 -7240
rect 11474 -7296 11497 -7240
rect 11378 -7324 11497 -7296
rect 3773 -7760 3852 -7749
rect 3773 -7816 3784 -7760
rect 3840 -7816 3852 -7760
rect 6215 -7767 6274 -7766
rect 3773 -7827 3852 -7816
rect 6209 -7778 6291 -7767
rect 3779 -7931 3838 -7827
rect 6209 -7834 6222 -7778
rect 6278 -7834 6291 -7778
rect 6209 -7844 6291 -7834
rect 9689 -7780 9768 -7769
rect 10946 -7771 11005 -7761
rect 9689 -7836 9700 -7780
rect 9756 -7836 9768 -7780
rect 6215 -7919 6274 -7844
rect 9689 -7847 9768 -7836
rect 10932 -7782 11011 -7771
rect 10932 -7838 10943 -7782
rect 10999 -7838 11011 -7782
rect 6210 -7930 6292 -7919
rect 3768 -7942 3847 -7931
rect 3768 -7998 3779 -7942
rect 3835 -7998 3847 -7942
rect 6210 -7986 6223 -7930
rect 6279 -7986 6292 -7930
rect 9697 -7934 9761 -7847
rect 10932 -7849 11011 -7838
rect 13383 -7794 13451 -6710
rect 13383 -7805 13466 -7794
rect 6210 -7996 6292 -7986
rect 9693 -7945 9772 -7934
rect 3768 -8009 3847 -7998
rect 3779 -8102 3838 -8009
rect 2891 -8820 2973 -8812
rect 3138 -8820 3220 -8812
rect 6215 -8820 6274 -7996
rect 9693 -8001 9704 -7945
rect 9760 -8001 9772 -7945
rect 10946 -7989 11005 -7849
rect 13383 -7861 13398 -7805
rect 13454 -7861 13466 -7805
rect 13383 -7872 13466 -7861
rect 9693 -8012 9772 -8001
rect 10930 -8000 11009 -7989
rect 2889 -8823 6274 -8820
rect 2889 -8879 2904 -8823
rect 2960 -8879 3151 -8823
rect 3207 -8879 6274 -8823
rect 9697 -8767 9761 -8012
rect 10930 -8056 10941 -8000
rect 10997 -8056 11009 -8000
rect 10930 -8067 11009 -8056
rect 13383 -8009 13451 -7872
rect 13383 -8020 13464 -8009
rect 10946 -8604 11005 -8067
rect 13383 -8076 13396 -8020
rect 13452 -8076 13464 -8020
rect 13383 -8087 13464 -8076
rect 13383 -8181 13451 -8087
rect 14745 -8604 14804 -4977
rect 16634 -5687 16714 -4517
rect 20975 -4913 21052 -3076
rect 22854 -4442 22919 -1710
rect 26504 -4438 26617 -4403
rect 26504 -4442 26528 -4438
rect 22854 -4494 26528 -4442
rect 26584 -4442 26617 -4438
rect 27040 -4442 27105 -4441
rect 26584 -4494 27124 -4442
rect 22854 -4507 27124 -4494
rect 21312 -4913 21391 -4908
rect 20975 -4919 21395 -4913
rect 20975 -4925 21323 -4919
rect 20975 -4981 21030 -4925
rect 21086 -4975 21323 -4925
rect 21379 -4975 21395 -4919
rect 22063 -4936 22142 -4935
rect 23591 -4936 23670 -4932
rect 21899 -4943 23670 -4936
rect 21086 -4981 21395 -4975
rect 20975 -4990 21395 -4981
rect 21894 -4946 23602 -4943
rect 21894 -4954 22074 -4946
rect 21019 -4992 21098 -4990
rect 21894 -5010 21905 -4954
rect 21961 -5002 22074 -4954
rect 22130 -4951 23602 -4946
rect 22130 -5002 23380 -4951
rect 21961 -5007 23380 -5002
rect 23436 -4999 23602 -4951
rect 23658 -4999 23670 -4943
rect 23436 -5007 23670 -4999
rect 21961 -5010 23670 -5007
rect 21894 -5013 23657 -5010
rect 21894 -5021 21973 -5013
rect 23369 -5018 23448 -5013
rect 16634 -5767 17596 -5687
rect 17516 -7552 17596 -5767
rect 26706 -5994 26785 -5983
rect 26706 -5999 26717 -5994
rect 26688 -6050 26717 -5999
rect 26773 -5999 26785 -5994
rect 27040 -5985 27105 -4507
rect 27040 -5996 27126 -5985
rect 27040 -5999 27058 -5996
rect 26773 -6050 27058 -5999
rect 26688 -6052 27058 -6050
rect 27114 -6052 27126 -5996
rect 26688 -6063 27126 -6052
rect 26688 -6064 27105 -6063
rect 10946 -8663 14804 -8604
rect 15488 -7632 17596 -7552
rect 15488 -8767 15568 -7632
rect 9697 -8847 15568 -8767
rect 2891 -8889 2973 -8879
rect 3138 -8889 3220 -8879
rect 634 -8917 713 -8914
rect 911 -8917 1056 -8913
rect 626 -8924 1056 -8917
rect 626 -8925 922 -8924
rect 626 -8981 645 -8925
rect 701 -8980 922 -8925
rect 978 -8980 1056 -8924
rect 701 -8981 1056 -8980
rect 626 -8997 1056 -8981
rect 1480 -9246 2100 -9240
rect 1480 -9252 2010 -9246
rect 1480 -9255 1859 -9252
rect 1480 -9257 1732 -9255
rect 1480 -9262 1615 -9257
rect 1480 -9318 1500 -9262
rect 1556 -9313 1615 -9262
rect 1671 -9311 1732 -9257
rect 1788 -9308 1859 -9255
rect 1915 -9302 2010 -9252
rect 2066 -9302 2100 -9246
rect 1915 -9308 2100 -9302
rect 1788 -9311 2100 -9308
rect 1671 -9313 2100 -9311
rect 1556 -9318 2100 -9313
rect 1480 -9380 2100 -9318
rect 1480 -9382 1627 -9380
rect 1480 -9438 1512 -9382
rect 1568 -9436 1627 -9382
rect 1683 -9382 2100 -9380
rect 1683 -9436 1770 -9382
rect 1568 -9438 1770 -9436
rect 1826 -9438 1900 -9382
rect 1956 -9384 2100 -9382
rect 1956 -9438 2024 -9384
rect 1480 -9440 2024 -9438
rect 2080 -9440 2100 -9384
rect 1480 -9460 2100 -9440
rect 11128 -9457 11694 -9418
rect 11128 -9463 11424 -9457
rect 11128 -9466 11282 -9463
rect 11128 -9522 11158 -9466
rect 11214 -9519 11282 -9466
rect 11338 -9513 11424 -9463
rect 11480 -9459 11694 -9457
rect 11480 -9513 11568 -9459
rect 11338 -9515 11568 -9513
rect 11624 -9515 11694 -9459
rect 11338 -9519 11694 -9515
rect 11214 -9522 11694 -9519
rect 11128 -9574 11694 -9522
rect 11128 -9576 11421 -9574
rect 11128 -9581 11281 -9576
rect 11128 -9637 11154 -9581
rect 11210 -9632 11281 -9581
rect 11337 -9630 11421 -9576
rect 11477 -9578 11694 -9574
rect 11477 -9630 11562 -9578
rect 11337 -9632 11562 -9630
rect 11210 -9634 11562 -9632
rect 11618 -9634 11694 -9578
rect 11210 -9637 11694 -9634
rect 11128 -9656 11694 -9637
rect 19341 -9450 19907 -9411
rect 19341 -9456 19637 -9450
rect 19341 -9459 19495 -9456
rect 19341 -9515 19371 -9459
rect 19427 -9512 19495 -9459
rect 19551 -9506 19637 -9456
rect 19693 -9452 19907 -9450
rect 19693 -9506 19781 -9452
rect 19551 -9508 19781 -9506
rect 19837 -9508 19907 -9452
rect 19551 -9512 19907 -9508
rect 19427 -9515 19907 -9512
rect 19341 -9567 19907 -9515
rect 19341 -9569 19634 -9567
rect 19341 -9574 19494 -9569
rect 19341 -9630 19367 -9574
rect 19423 -9625 19494 -9574
rect 19550 -9623 19634 -9569
rect 19690 -9571 19907 -9567
rect 19690 -9623 19775 -9571
rect 19550 -9625 19775 -9623
rect 19423 -9627 19775 -9625
rect 19831 -9627 19907 -9571
rect 19423 -9630 19907 -9627
rect 26403 -9431 26969 -9392
rect 26403 -9437 26699 -9431
rect 26403 -9440 26557 -9437
rect 26403 -9496 26433 -9440
rect 26489 -9493 26557 -9440
rect 26613 -9487 26699 -9437
rect 26755 -9433 26969 -9431
rect 26755 -9487 26843 -9433
rect 26613 -9489 26843 -9487
rect 26899 -9489 26969 -9433
rect 26613 -9493 26969 -9489
rect 26489 -9496 26969 -9493
rect 26403 -9548 26969 -9496
rect 26403 -9550 26696 -9548
rect 26403 -9555 26556 -9550
rect 26403 -9611 26429 -9555
rect 26485 -9606 26556 -9555
rect 26612 -9604 26696 -9550
rect 26752 -9552 26969 -9548
rect 26752 -9604 26837 -9552
rect 26612 -9606 26837 -9604
rect 26485 -9608 26837 -9606
rect 26893 -9608 26969 -9552
rect 26485 -9611 26969 -9608
rect 26403 -9630 26969 -9611
rect 33208 -9429 33774 -9390
rect 33208 -9435 33504 -9429
rect 33208 -9438 33362 -9435
rect 33208 -9494 33238 -9438
rect 33294 -9491 33362 -9438
rect 33418 -9485 33504 -9435
rect 33560 -9431 33774 -9429
rect 33560 -9485 33648 -9431
rect 33418 -9487 33648 -9485
rect 33704 -9487 33774 -9431
rect 33418 -9491 33774 -9487
rect 33294 -9494 33774 -9491
rect 33208 -9546 33774 -9494
rect 33208 -9548 33501 -9546
rect 33208 -9553 33361 -9548
rect 33208 -9609 33234 -9553
rect 33290 -9604 33361 -9553
rect 33417 -9602 33501 -9548
rect 33557 -9550 33774 -9546
rect 33557 -9602 33642 -9550
rect 33417 -9604 33642 -9602
rect 33290 -9606 33642 -9604
rect 33698 -9606 33774 -9550
rect 33290 -9609 33774 -9606
rect 33208 -9628 33774 -9609
rect 19341 -9649 19907 -9630
rect 15100 -9880 15666 -9841
rect 15100 -9886 15396 -9880
rect 15100 -9889 15254 -9886
rect 5214 -9962 5780 -9923
rect 5214 -9968 5510 -9962
rect 5214 -9971 5368 -9968
rect 5214 -10027 5244 -9971
rect 5300 -10024 5368 -9971
rect 5424 -10018 5510 -9968
rect 5566 -9964 5780 -9962
rect 5566 -10018 5654 -9964
rect 5424 -10020 5654 -10018
rect 5710 -10020 5780 -9964
rect 5424 -10024 5780 -10020
rect 5300 -10027 5780 -10024
rect 5214 -10079 5780 -10027
rect 15100 -9945 15130 -9889
rect 15186 -9942 15254 -9889
rect 15310 -9936 15396 -9886
rect 15452 -9882 15666 -9880
rect 15452 -9936 15540 -9882
rect 15310 -9938 15540 -9936
rect 15596 -9938 15666 -9882
rect 15310 -9942 15666 -9938
rect 15186 -9945 15666 -9942
rect 15100 -9997 15666 -9945
rect 15100 -9999 15393 -9997
rect 15100 -10004 15253 -9999
rect 15100 -10060 15126 -10004
rect 15182 -10055 15253 -10004
rect 15309 -10053 15393 -9999
rect 15449 -10001 15666 -9997
rect 15449 -10053 15534 -10001
rect 15309 -10055 15534 -10053
rect 15182 -10057 15534 -10055
rect 15590 -10057 15666 -10001
rect 22631 -9850 23197 -9811
rect 22631 -9856 22927 -9850
rect 22631 -9859 22785 -9856
rect 22631 -9915 22661 -9859
rect 22717 -9912 22785 -9859
rect 22841 -9906 22927 -9856
rect 22983 -9852 23197 -9850
rect 22983 -9906 23071 -9852
rect 22841 -9908 23071 -9906
rect 23127 -9908 23197 -9852
rect 22841 -9912 23197 -9908
rect 22717 -9915 23197 -9912
rect 22631 -9967 23197 -9915
rect 22631 -9969 22924 -9967
rect 22631 -9974 22784 -9969
rect 22631 -10030 22657 -9974
rect 22713 -10025 22784 -9974
rect 22840 -10023 22924 -9969
rect 22980 -9971 23197 -9967
rect 22980 -10023 23065 -9971
rect 22840 -10025 23065 -10023
rect 22713 -10027 23065 -10025
rect 23121 -10027 23197 -9971
rect 22713 -10030 23197 -10027
rect 22631 -10049 23197 -10030
rect 15182 -10060 15666 -10057
rect 15100 -10079 15666 -10060
rect 5214 -10081 5507 -10079
rect 5214 -10086 5367 -10081
rect 5214 -10142 5240 -10086
rect 5296 -10137 5367 -10086
rect 5423 -10135 5507 -10081
rect 5563 -10083 5780 -10079
rect 5563 -10135 5648 -10083
rect 5423 -10137 5648 -10135
rect 5296 -10139 5648 -10137
rect 5704 -10139 5780 -10083
rect 5296 -10142 5780 -10139
rect 5214 -10161 5780 -10142
<< via3 >>
rect 4997 11902 5053 11958
rect 5121 11905 5177 11961
rect 5263 11911 5319 11967
rect 5407 11909 5463 11965
rect 4993 11787 5049 11843
rect 5120 11792 5176 11848
rect 5260 11794 5316 11850
rect 5401 11790 5457 11846
rect 1634 11568 1690 11624
rect 1758 11571 1814 11627
rect 1900 11577 1956 11633
rect 2044 11575 2100 11631
rect 1630 11453 1686 11509
rect 1757 11458 1813 11514
rect 1897 11460 1953 11516
rect 2038 11456 2094 11512
rect 5156 10516 5212 10572
rect 1703 9519 1759 9575
rect 22653 12018 22709 12074
rect 22777 12021 22833 12077
rect 22919 12027 22975 12083
rect 23063 12025 23119 12081
rect 15130 11892 15186 11948
rect 15254 11895 15310 11951
rect 15396 11901 15452 11957
rect 15540 11899 15596 11955
rect 22649 11903 22705 11959
rect 22776 11908 22832 11964
rect 22916 11910 22972 11966
rect 23057 11906 23113 11962
rect 15126 11777 15182 11833
rect 15253 11782 15309 11838
rect 15393 11784 15449 11840
rect 15534 11780 15590 11836
rect 11293 11681 11349 11737
rect 11417 11684 11473 11740
rect 11559 11690 11615 11746
rect 11703 11688 11759 11744
rect 11289 11566 11345 11622
rect 11416 11571 11472 11627
rect 11556 11573 11612 11629
rect 11697 11569 11753 11625
rect 11530 8424 11586 8480
rect 1683 7945 1739 8001
rect 11515 7843 11571 7899
rect 5151 5294 5207 5350
rect 19158 11645 19214 11701
rect 19282 11648 19338 11704
rect 19424 11654 19480 11710
rect 19568 11652 19624 11708
rect 19154 11530 19210 11586
rect 19281 11535 19337 11591
rect 19421 11537 19477 11593
rect 19562 11533 19618 11589
rect 19521 8750 19577 8806
rect 19469 7555 19525 7611
rect 15519 5680 15575 5736
rect 19476 3558 19532 3614
rect 1739 2749 1795 2805
rect 22904 5677 22960 5733
rect 26139 11627 26195 11683
rect 26263 11630 26319 11686
rect 26405 11636 26461 11692
rect 26549 11634 26605 11690
rect 26135 11512 26191 11568
rect 26262 11517 26318 11573
rect 26402 11519 26458 11575
rect 26543 11515 26599 11571
rect 26568 8361 26624 8417
rect 33012 11699 33068 11755
rect 33136 11702 33192 11758
rect 33278 11708 33334 11764
rect 33422 11706 33478 11762
rect 33008 11584 33064 11640
rect 33135 11589 33191 11645
rect 33275 11591 33331 11647
rect 33416 11587 33472 11643
rect 1775 -2484 1831 -2428
rect 5576 -4256 5632 -4200
rect 11496 2663 11552 2719
rect 26465 2633 26521 2689
rect 15215 463 15271 519
rect 11603 -2852 11659 -2796
rect 15464 -4242 15520 -4186
rect 11418 -7296 11474 -7240
rect 26528 -4494 26584 -4438
rect 1500 -9318 1556 -9262
rect 1615 -9313 1671 -9257
rect 1732 -9311 1788 -9255
rect 1859 -9308 1915 -9252
rect 2010 -9302 2066 -9246
rect 1512 -9438 1568 -9382
rect 1627 -9436 1683 -9380
rect 1770 -9438 1826 -9382
rect 1900 -9438 1956 -9382
rect 2024 -9440 2080 -9384
rect 11158 -9522 11214 -9466
rect 11282 -9519 11338 -9463
rect 11424 -9513 11480 -9457
rect 11568 -9515 11624 -9459
rect 11154 -9637 11210 -9581
rect 11281 -9632 11337 -9576
rect 11421 -9630 11477 -9574
rect 11562 -9634 11618 -9578
rect 19371 -9515 19427 -9459
rect 19495 -9512 19551 -9456
rect 19637 -9506 19693 -9450
rect 19781 -9508 19837 -9452
rect 19367 -9630 19423 -9574
rect 19494 -9625 19550 -9569
rect 19634 -9623 19690 -9567
rect 19775 -9627 19831 -9571
rect 26433 -9496 26489 -9440
rect 26557 -9493 26613 -9437
rect 26699 -9487 26755 -9431
rect 26843 -9489 26899 -9433
rect 26429 -9611 26485 -9555
rect 26556 -9606 26612 -9550
rect 26696 -9604 26752 -9548
rect 26837 -9608 26893 -9552
rect 33238 -9494 33294 -9438
rect 33362 -9491 33418 -9435
rect 33504 -9485 33560 -9429
rect 33648 -9487 33704 -9431
rect 33234 -9609 33290 -9553
rect 33361 -9604 33417 -9548
rect 33501 -9602 33557 -9546
rect 33642 -9606 33698 -9550
rect 5244 -10027 5300 -9971
rect 5368 -10024 5424 -9968
rect 5510 -10018 5566 -9962
rect 5654 -10020 5710 -9964
rect 15130 -9945 15186 -9889
rect 15254 -9942 15310 -9886
rect 15396 -9936 15452 -9880
rect 15540 -9938 15596 -9882
rect 15126 -10060 15182 -10004
rect 15253 -10055 15309 -9999
rect 15393 -10053 15449 -9997
rect 15534 -10057 15590 -10001
rect 22661 -9915 22717 -9859
rect 22785 -9912 22841 -9856
rect 22927 -9906 22983 -9850
rect 23071 -9908 23127 -9852
rect 22657 -10030 22713 -9974
rect 22784 -10025 22840 -9969
rect 22924 -10023 22980 -9967
rect 23065 -10027 23121 -9971
rect 5240 -10142 5296 -10086
rect 5367 -10137 5423 -10081
rect 5507 -10135 5563 -10079
rect 5648 -10139 5704 -10083
<< metal4 >>
rect 4975 12195 23146 12672
rect 4975 12011 5452 12195
rect 4975 12006 5529 12011
rect 4967 11967 5533 12006
rect 15139 12001 15616 12195
rect 22669 12127 23146 12195
rect 22669 12122 23185 12127
rect 22623 12083 23189 12122
rect 22623 12077 22919 12083
rect 22623 12074 22777 12077
rect 22623 12018 22653 12074
rect 22709 12021 22777 12074
rect 22833 12027 22919 12077
rect 22975 12081 23189 12083
rect 22975 12027 23063 12081
rect 22833 12025 23063 12027
rect 23119 12025 23189 12081
rect 22833 12021 23189 12025
rect 22709 12018 23189 12021
rect 22623 12010 23189 12018
rect 15139 11996 15662 12001
rect 4967 11961 5263 11967
rect 4967 11958 5121 11961
rect 4967 11902 4997 11958
rect 5053 11905 5121 11958
rect 5177 11911 5263 11961
rect 5319 11965 5533 11967
rect 5319 11911 5407 11965
rect 5177 11909 5407 11911
rect 5463 11909 5533 11965
rect 5177 11905 5533 11909
rect 5053 11902 5533 11905
rect 4967 11850 5533 11902
rect 4967 11848 5260 11850
rect 4967 11843 5120 11848
rect 4967 11787 4993 11843
rect 5049 11792 5120 11843
rect 5176 11794 5260 11848
rect 5316 11846 5533 11850
rect 5316 11794 5401 11846
rect 5176 11792 5401 11794
rect 5049 11790 5401 11792
rect 5457 11790 5533 11846
rect 5049 11787 5533 11790
rect 4967 11768 5533 11787
rect 15100 11957 15666 11996
rect 15100 11951 15396 11957
rect 15100 11948 15254 11951
rect 15100 11892 15130 11948
rect 15186 11895 15254 11948
rect 15310 11901 15396 11951
rect 15452 11955 15666 11957
rect 15452 11901 15540 11955
rect 15310 11899 15540 11901
rect 15596 11899 15666 11955
rect 15310 11895 15666 11899
rect 15186 11892 15666 11895
rect 15100 11840 15666 11892
rect 22623 11966 23190 12010
rect 22623 11964 22916 11966
rect 22623 11959 22776 11964
rect 22623 11903 22649 11959
rect 22705 11908 22776 11959
rect 22832 11910 22916 11964
rect 22972 11962 23190 11966
rect 22972 11910 23057 11962
rect 22832 11908 23057 11910
rect 22705 11906 23057 11908
rect 23113 11906 23190 11962
rect 22705 11903 23190 11906
rect 22623 11884 23190 11903
rect 15100 11838 15393 11840
rect 15100 11833 15253 11838
rect 1604 11633 2170 11672
rect 1604 11627 1900 11633
rect 1604 11624 1758 11627
rect 1604 11568 1634 11624
rect 1690 11571 1758 11624
rect 1814 11577 1900 11627
rect 1956 11631 2170 11633
rect 1956 11577 2044 11631
rect 1814 11575 2044 11577
rect 2100 11575 2170 11631
rect 1814 11571 2170 11575
rect 1690 11568 2170 11571
rect 1604 11517 2170 11568
rect 1593 11516 2170 11517
rect 1593 11514 1897 11516
rect 1593 11509 1757 11514
rect 1593 11453 1630 11509
rect 1686 11458 1757 11509
rect 1813 11460 1897 11514
rect 1953 11512 2170 11516
rect 1953 11460 2038 11512
rect 1813 11458 2038 11460
rect 1686 11456 2038 11458
rect 2094 11456 2170 11512
rect 1686 11453 2170 11456
rect 1593 11434 2170 11453
rect 1593 9575 2072 11434
rect 1593 9519 1703 9575
rect 1759 9519 2072 9575
rect 1593 8001 2072 9519
rect 1593 7945 1683 8001
rect 1739 7945 2072 8001
rect 1593 5410 2072 7945
rect 4975 10572 5452 11768
rect 11263 11746 11829 11785
rect 15100 11777 15126 11833
rect 15182 11782 15253 11833
rect 15309 11784 15393 11838
rect 15449 11836 15666 11840
rect 15449 11784 15534 11836
rect 15309 11782 15534 11784
rect 15182 11780 15534 11782
rect 15590 11780 15666 11836
rect 15182 11777 15666 11780
rect 15100 11758 15666 11777
rect 11263 11740 11559 11746
rect 11263 11737 11417 11740
rect 11263 11681 11293 11737
rect 11349 11684 11417 11737
rect 11473 11690 11559 11740
rect 11615 11744 11829 11746
rect 11615 11690 11703 11744
rect 11473 11688 11703 11690
rect 11759 11688 11829 11744
rect 11473 11684 11829 11688
rect 11349 11681 11829 11684
rect 11263 11629 11829 11681
rect 11263 11627 11556 11629
rect 11263 11622 11416 11627
rect 11263 11614 11289 11622
rect 4975 10516 5156 10572
rect 5212 10516 5452 10572
rect 4975 5350 5452 10516
rect 4975 5294 5151 5350
rect 5207 5294 5452 5350
rect 1593 2805 2072 5280
rect 1593 2749 1739 2805
rect 1795 2749 2072 2805
rect 1593 -2428 2072 2749
rect 1593 -2484 1775 -2428
rect 1831 -2484 2072 -2428
rect 1593 -9240 2072 -2484
rect 4975 -4173 5452 5294
rect 11261 11566 11289 11614
rect 11345 11571 11416 11622
rect 11472 11573 11556 11627
rect 11612 11625 11829 11629
rect 11612 11573 11697 11625
rect 11472 11571 11697 11573
rect 11345 11569 11697 11571
rect 11753 11569 11829 11625
rect 11345 11566 11829 11569
rect 11261 11547 11829 11566
rect 11261 8480 11690 11547
rect 11261 8424 11530 8480
rect 11586 8424 11690 8480
rect 11261 7899 11690 8424
rect 11261 7843 11515 7899
rect 11571 7843 11690 7899
rect 11261 2719 11690 7843
rect 11261 2663 11496 2719
rect 11552 2663 11690 2719
rect 11261 -2753 11690 2663
rect 15139 5736 15616 11758
rect 19128 11710 19694 11749
rect 19128 11704 19424 11710
rect 19128 11701 19282 11704
rect 19128 11645 19158 11701
rect 19214 11648 19282 11701
rect 19338 11654 19424 11704
rect 19480 11708 19694 11710
rect 19480 11654 19568 11708
rect 19338 11652 19568 11654
rect 19624 11652 19694 11708
rect 19338 11648 19694 11652
rect 19214 11645 19694 11648
rect 19128 11636 19694 11645
rect 19128 11593 19716 11636
rect 22669 11626 23190 11884
rect 32982 11764 33548 11803
rect 32982 11758 33278 11764
rect 32982 11755 33136 11758
rect 19128 11591 19421 11593
rect 19128 11586 19281 11591
rect 19128 11530 19154 11586
rect 19210 11535 19281 11586
rect 19337 11537 19421 11591
rect 19477 11589 19716 11593
rect 19477 11537 19562 11589
rect 19337 11535 19562 11537
rect 19210 11533 19562 11535
rect 19618 11533 19716 11589
rect 19210 11530 19716 11533
rect 19128 11511 19716 11530
rect 15139 5680 15519 5736
rect 15575 5680 15616 5736
rect 15139 519 15616 5680
rect 15139 463 15215 519
rect 15271 463 15616 519
rect 11261 -2796 11705 -2753
rect 11261 -2852 11603 -2796
rect 11659 -2852 11705 -2796
rect 11261 -2904 11705 -2852
rect 4975 -4200 5660 -4173
rect 4975 -4256 5576 -4200
rect 5632 -4256 5660 -4200
rect 4975 -4284 5660 -4256
rect 1480 -9246 2100 -9240
rect 1480 -9252 2010 -9246
rect 1480 -9255 1859 -9252
rect 1480 -9257 1732 -9255
rect 1480 -9262 1615 -9257
rect 1480 -9318 1500 -9262
rect 1556 -9313 1615 -9262
rect 1671 -9311 1732 -9257
rect 1788 -9308 1859 -9255
rect 1915 -9302 2010 -9252
rect 2066 -9302 2100 -9246
rect 1915 -9308 2100 -9302
rect 1788 -9311 2100 -9308
rect 1671 -9313 2100 -9311
rect 1556 -9318 2100 -9313
rect 1480 -9380 2100 -9318
rect 1480 -9382 1627 -9380
rect 1480 -9438 1512 -9382
rect 1568 -9436 1627 -9382
rect 1683 -9382 2100 -9380
rect 1683 -9436 1770 -9382
rect 1568 -9438 1770 -9436
rect 1826 -9438 1900 -9382
rect 1956 -9384 2100 -9382
rect 1956 -9438 2024 -9384
rect 1480 -9440 2024 -9438
rect 2080 -9440 2100 -9384
rect 1480 -9460 2100 -9440
rect 4975 -9737 5452 -4284
rect 11261 -7240 11690 -2904
rect 11261 -7296 11418 -7240
rect 11474 -7296 11690 -7240
rect 11261 -9418 11690 -7296
rect 15139 -4186 15616 463
rect 15139 -4242 15464 -4186
rect 15520 -4242 15616 -4186
rect 11128 -9457 11694 -9418
rect 11128 -9463 11424 -9457
rect 11128 -9466 11282 -9463
rect 11128 -9522 11158 -9466
rect 11214 -9519 11282 -9466
rect 11338 -9513 11424 -9463
rect 11480 -9459 11694 -9457
rect 11480 -9513 11568 -9459
rect 11338 -9515 11568 -9513
rect 11624 -9515 11694 -9459
rect 11338 -9519 11694 -9515
rect 11214 -9522 11694 -9519
rect 11128 -9574 11694 -9522
rect 11128 -9576 11421 -9574
rect 11128 -9581 11281 -9576
rect 11128 -9637 11154 -9581
rect 11210 -9632 11281 -9581
rect 11337 -9630 11421 -9576
rect 11477 -9578 11694 -9574
rect 11477 -9630 11562 -9578
rect 11337 -9632 11562 -9630
rect 11210 -9634 11562 -9632
rect 11618 -9634 11694 -9578
rect 11210 -9637 11694 -9634
rect 11128 -9656 11694 -9637
rect 4975 -9817 5782 -9737
rect 15139 -9817 15616 -4242
rect 19287 8806 19716 11511
rect 19287 8750 19521 8806
rect 19577 8750 19716 8806
rect 19287 7611 19716 8750
rect 19287 7555 19469 7611
rect 19525 7555 19716 7611
rect 19287 3614 19716 7555
rect 19287 3558 19476 3614
rect 19532 3558 19716 3614
rect 19287 -9411 19716 3558
rect 22713 5733 23190 11626
rect 26109 11692 26675 11731
rect 26109 11686 26405 11692
rect 26109 11683 26263 11686
rect 26109 11627 26139 11683
rect 26195 11630 26263 11683
rect 26319 11636 26405 11686
rect 26461 11690 26675 11692
rect 26461 11636 26549 11690
rect 26319 11634 26549 11636
rect 26605 11675 26675 11690
rect 32982 11699 33012 11755
rect 33068 11702 33136 11755
rect 33192 11708 33278 11758
rect 33334 11762 33548 11764
rect 33334 11708 33422 11762
rect 33192 11706 33422 11708
rect 33478 11722 33548 11762
rect 33478 11706 33736 11722
rect 33192 11702 33736 11706
rect 33068 11699 33736 11702
rect 26605 11634 26820 11675
rect 26319 11630 26820 11634
rect 26195 11627 26820 11630
rect 26109 11575 26820 11627
rect 26109 11573 26402 11575
rect 26109 11568 26262 11573
rect 26109 11512 26135 11568
rect 26191 11517 26262 11568
rect 26318 11519 26402 11573
rect 26458 11571 26820 11575
rect 26458 11519 26543 11571
rect 26318 11517 26543 11519
rect 26191 11515 26543 11517
rect 26599 11515 26820 11571
rect 32982 11647 33736 11699
rect 32982 11645 33275 11647
rect 32982 11640 33135 11645
rect 32982 11584 33008 11640
rect 33064 11589 33135 11640
rect 33191 11591 33275 11645
rect 33331 11643 33736 11647
rect 33331 11591 33416 11643
rect 33191 11589 33416 11591
rect 33064 11587 33416 11589
rect 33472 11587 33736 11643
rect 33064 11584 33736 11587
rect 32982 11565 33736 11584
rect 26191 11512 26820 11515
rect 26109 11493 26820 11512
rect 22713 5677 22904 5733
rect 22960 5677 23190 5733
rect 19287 -9449 19907 -9411
rect 19341 -9450 19907 -9449
rect 19341 -9456 19637 -9450
rect 19341 -9459 19495 -9456
rect 19341 -9515 19371 -9459
rect 19427 -9512 19495 -9459
rect 19551 -9506 19637 -9456
rect 19693 -9452 19907 -9450
rect 19693 -9506 19781 -9452
rect 19551 -9508 19781 -9506
rect 19837 -9508 19907 -9452
rect 19551 -9512 19907 -9508
rect 19427 -9515 19907 -9512
rect 19341 -9567 19907 -9515
rect 19341 -9569 19634 -9567
rect 19341 -9574 19494 -9569
rect 19341 -9630 19367 -9574
rect 19423 -9625 19494 -9574
rect 19550 -9623 19634 -9569
rect 19690 -9571 19907 -9567
rect 19690 -9623 19775 -9571
rect 19550 -9625 19775 -9623
rect 19423 -9627 19775 -9625
rect 19831 -9627 19907 -9571
rect 19423 -9630 19907 -9627
rect 19341 -9649 19907 -9630
rect 22713 -9806 23190 5677
rect 26391 8417 26820 11493
rect 26391 8361 26568 8417
rect 26624 8361 26820 8417
rect 26391 2689 26820 8361
rect 26391 2633 26465 2689
rect 26521 2633 26820 2689
rect 26391 -4438 26820 2633
rect 26391 -4494 26528 -4438
rect 26584 -4494 26820 -4438
rect 26391 -9392 26820 -4494
rect 33273 -9390 33736 11565
rect 26391 -9410 26969 -9392
rect 26403 -9431 26969 -9410
rect 26403 -9437 26699 -9431
rect 26403 -9440 26557 -9437
rect 26403 -9496 26433 -9440
rect 26489 -9493 26557 -9440
rect 26613 -9487 26699 -9437
rect 26755 -9433 26969 -9431
rect 26755 -9487 26843 -9433
rect 26613 -9489 26843 -9487
rect 26899 -9489 26969 -9433
rect 26613 -9493 26969 -9489
rect 26489 -9496 26969 -9493
rect 26403 -9548 26969 -9496
rect 26403 -9550 26696 -9548
rect 26403 -9555 26556 -9550
rect 26403 -9611 26429 -9555
rect 26485 -9606 26556 -9555
rect 26612 -9604 26696 -9550
rect 26752 -9552 26969 -9548
rect 26752 -9604 26837 -9552
rect 26612 -9606 26837 -9604
rect 26485 -9608 26837 -9606
rect 26893 -9608 26969 -9552
rect 26485 -9611 26969 -9608
rect 26403 -9630 26969 -9611
rect 33208 -9429 33774 -9390
rect 33208 -9435 33504 -9429
rect 33208 -9438 33362 -9435
rect 33208 -9494 33238 -9438
rect 33294 -9491 33362 -9438
rect 33418 -9485 33504 -9435
rect 33560 -9431 33774 -9429
rect 33560 -9485 33648 -9431
rect 33418 -9487 33648 -9485
rect 33704 -9487 33774 -9431
rect 33418 -9491 33774 -9487
rect 33294 -9494 33774 -9491
rect 33208 -9546 33774 -9494
rect 33208 -9548 33501 -9546
rect 33208 -9553 33361 -9548
rect 33208 -9609 33234 -9553
rect 33290 -9604 33361 -9553
rect 33417 -9602 33501 -9548
rect 33557 -9550 33774 -9546
rect 33557 -9602 33642 -9550
rect 33417 -9604 33642 -9602
rect 33290 -9606 33642 -9604
rect 33698 -9606 33774 -9550
rect 33290 -9609 33774 -9606
rect 33208 -9628 33774 -9609
rect 22713 -9811 23193 -9806
rect 22631 -9817 23197 -9811
rect 4975 -9850 23244 -9817
rect 4975 -9856 22927 -9850
rect 4975 -9859 22785 -9856
rect 4975 -9880 22661 -9859
rect 4975 -9886 15396 -9880
rect 4975 -9889 15254 -9886
rect 4975 -9945 15130 -9889
rect 15186 -9942 15254 -9889
rect 15310 -9936 15396 -9886
rect 15452 -9882 22661 -9880
rect 15452 -9936 15540 -9882
rect 15310 -9938 15540 -9936
rect 15596 -9915 22661 -9882
rect 22717 -9912 22785 -9859
rect 22841 -9906 22927 -9856
rect 22983 -9852 23244 -9850
rect 22983 -9906 23071 -9852
rect 22841 -9908 23071 -9906
rect 23127 -9908 23244 -9852
rect 22841 -9912 23244 -9908
rect 22717 -9915 23244 -9912
rect 15596 -9938 23244 -9915
rect 15310 -9942 23244 -9938
rect 15186 -9945 23244 -9942
rect 4975 -9962 23244 -9945
rect 4975 -9968 5510 -9962
rect 4975 -9971 5368 -9968
rect 4975 -10027 5244 -9971
rect 5300 -10024 5368 -9971
rect 5424 -10018 5510 -9968
rect 5566 -9964 23244 -9962
rect 5566 -10018 5654 -9964
rect 5424 -10020 5654 -10018
rect 5710 -9967 23244 -9964
rect 5710 -9969 22924 -9967
rect 5710 -9974 22784 -9969
rect 5710 -9997 22657 -9974
rect 5710 -9999 15393 -9997
rect 5710 -10004 15253 -9999
rect 5710 -10020 15126 -10004
rect 5424 -10024 15126 -10020
rect 5300 -10027 15126 -10024
rect 4975 -10060 15126 -10027
rect 15182 -10055 15253 -10004
rect 15309 -10053 15393 -9999
rect 15449 -10001 22657 -9997
rect 15449 -10053 15534 -10001
rect 15309 -10055 15534 -10053
rect 15182 -10057 15534 -10055
rect 15590 -10030 22657 -10001
rect 22713 -10025 22784 -9974
rect 22840 -10023 22924 -9969
rect 22980 -9971 23244 -9967
rect 22980 -10023 23065 -9971
rect 22840 -10025 23065 -10023
rect 22713 -10027 23065 -10025
rect 23121 -10027 23244 -9971
rect 22713 -10030 23244 -10027
rect 15590 -10057 23244 -10030
rect 15182 -10060 23244 -10057
rect 4975 -10079 23244 -10060
rect 4975 -10081 5507 -10079
rect 4975 -10086 5367 -10081
rect 4975 -10142 5240 -10086
rect 5296 -10137 5367 -10086
rect 5423 -10135 5507 -10081
rect 5563 -10083 23244 -10079
rect 5563 -10135 5648 -10083
rect 5423 -10137 5648 -10135
rect 5296 -10139 5648 -10137
rect 5704 -10084 23244 -10083
rect 5704 -10139 5782 -10084
rect 5296 -10142 5782 -10139
rect 4975 -10214 5782 -10142
use 7b_counter  7b_counter_0
timestamp 1713971515
transform 1 0 155 0 1 5517
box -155 -5517 33192 5581
use DFF_magic  DFF_magic_0
timestamp 1713971515
transform 1 0 25560 0 1 -2039
box -2075 -819 5510 1706
use divide_by_2  divide_by_2_0
timestamp 1713971633
transform 1 0 26748 0 1 -6541
box -2075 -819 5510 1759
use divide_by_2  divide_by_2_1
timestamp 1713971633
transform 1 0 32663 0 1 1452
box -2075 -819 5510 1759
use mux_magic  mux_magic_0
timestamp 1713277963
transform 1 0 33242 0 1 -1944
box -1637 -810 2187 1564
use OR_magic  OR_magic_1
timestamp 1713277963
transform 1 0 30279 0 1 4792
box 0 -1478 1136 611
use OR_magic  OR_magic_2
timestamp 1713277963
transform 1 0 23266 0 1 -5520
box 0 -1478 1136 611
use p2_gen_magic  p2_gen_magic_0
timestamp 1713971515
transform 1 0 315 0 1 -2358
box -265 -2108 22479 2062
use p3_gen_magic  p3_gen_magic_0
timestamp 1713971633
transform 1 0 315 0 1 -6856
box -265 -2148 22479 2078
<< labels >>
flabel metal1 s 22692 -1023 22692 -1023 0 FreeSans 750 0 0 0 P2
port 1 nsew
flabel metal1 s 22770 -937 22770 -937 0 FreeSans 750 0 0 0 P2
port 1 nsew
flabel metal1 s 35531 -1507 35531 -1507 0 FreeSans 750 0 0 0 OUT1
port 2 nsew
flabel metal1 s 33355 9801 33355 9801 0 FreeSans 750 0 0 0 VDD
port 3 nsew
flabel metal1 s 32299 -1851 32299 -1851 0 FreeSans 750 0 0 0 VSS
port 4 nsew
flabel metal1 s 24241 -358 24241 -358 0 FreeSans 750 0 0 0 CLK
port 5 nsew
flabel metal1 s 22530 9388 22530 9388 0 FreeSans 750 0 0 0 Q1
port 6 nsew
flabel metal1 s 15869 7770 15869 7770 0 FreeSans 750 0 0 0 D2_1
port 7 nsew
flabel metal1 s 13700 7760 13700 7760 0 FreeSans 750 0 0 0 D2_2
port 8 nsew
flabel metal1 s 6884 9750 6884 9750 0 FreeSans 750 0 0 0 Q2
port 9 nsew
flabel metal1 s 21770 1713 21770 1713 0 FreeSans 750 0 0 0 Q4
port 10 nsew
flabel metal1 s 28518 3285 28518 3285 0 FreeSans 750 0 0 0 D2_4
port 11 nsew
flabel metal1 s 22634 4559 22634 4559 0 FreeSans 750 0 0 0 Q3
port 12 nsew
flabel metal1 s 15859 2553 15859 2553 0 FreeSans 750 0 0 0 D2_3
port 13 nsew
flabel metal1 s 6893 4478 6893 4478 0 FreeSans 750 0 0 0 Q6
port 14 nsew
flabel metal1 s 13699 2548 13699 2548 0 FreeSans 750 0 0 0 D2_6
port 15 nsew
flabel metal1 s 7978 1275 7978 1275 0 FreeSans 750 0 0 0 Q5
port 16 nsew
flabel metal1 s 1170 3293 1170 3293 0 FreeSans 750 0 0 0 D2_5
port 17 nsew
flabel metal1 s 7836 6734 7836 6734 0 FreeSans 750 0 0 0 Q7
port 18 nsew
flabel metal1 s 1211 8502 1211 8502 0 FreeSans 750 0 0 0 D2_7
port 19 nsew
flabel metal1 s 174 9335 174 9335 0 FreeSans 750 0 0 0 LD
port 20 nsew
<< end >>
