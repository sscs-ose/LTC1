magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1591 -1045 1591 1045
<< metal1 >>
rect -591 39 591 45
rect -591 -39 -585 39
rect 585 -39 591 39
rect -591 -45 591 -39
<< via1 >>
rect -585 -39 585 39
<< metal2 >>
rect -591 39 591 45
rect -591 -39 -585 39
rect 585 -39 591 39
rect -591 -45 591 -39
<< end >>
