magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 2472 2444
<< mvnmos >>
rect 0 0 140 400
rect 244 0 384 400
<< mvndiff >>
rect -88 387 0 400
rect -88 341 -75 387
rect -29 341 0 387
rect -88 278 0 341
rect -88 232 -75 278
rect -29 232 0 278
rect -88 169 0 232
rect -88 123 -75 169
rect -29 123 0 169
rect -88 59 0 123
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 387 244 400
rect 140 341 169 387
rect 215 341 244 387
rect 140 278 244 341
rect 140 232 169 278
rect 215 232 244 278
rect 140 169 244 232
rect 140 123 169 169
rect 215 123 244 169
rect 140 59 244 123
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 387 472 400
rect 384 341 413 387
rect 459 341 472 387
rect 384 278 472 341
rect 384 232 413 278
rect 459 232 472 278
rect 384 169 472 232
rect 384 123 413 169
rect 459 123 472 169
rect 384 59 472 123
rect 384 13 413 59
rect 459 13 472 59
rect 384 0 472 13
<< mvndiffc >>
rect -75 341 -29 387
rect -75 232 -29 278
rect -75 123 -29 169
rect -75 13 -29 59
rect 169 341 215 387
rect 169 232 215 278
rect 169 123 215 169
rect 169 13 215 59
rect 413 341 459 387
rect 413 232 459 278
rect 413 123 459 169
rect 413 13 459 59
<< polysilicon >>
rect 0 400 140 444
rect 244 400 384 444
rect 0 -44 140 0
rect 244 -44 384 0
<< metal1 >>
rect -75 387 -29 400
rect -75 278 -29 341
rect -75 169 -29 232
rect -75 59 -29 123
rect -75 0 -29 13
rect 169 387 215 400
rect 169 278 215 341
rect 169 169 215 232
rect 169 59 215 123
rect 169 0 215 13
rect 413 387 459 400
rect 413 278 459 341
rect 413 169 459 232
rect 413 59 459 123
rect 413 0 459 13
<< labels >>
rlabel metal1 192 200 192 200 4 D
rlabel metal1 436 200 436 200 4 S
rlabel metal1 -52 200 -52 200 4 S
<< end >>
