magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2088 -2044 3204 2684
<< mvnmos >>
rect 0 0 140 640
rect 244 0 384 640
rect 488 0 628 640
rect 732 0 872 640
rect 976 0 1116 640
<< mvndiff >>
rect -88 627 0 640
rect -88 581 -75 627
rect -29 581 0 627
rect -88 514 0 581
rect -88 468 -75 514
rect -29 468 0 514
rect -88 401 0 468
rect -88 355 -75 401
rect -29 355 0 401
rect -88 287 0 355
rect -88 241 -75 287
rect -29 241 0 287
rect -88 173 0 241
rect -88 127 -75 173
rect -29 127 0 173
rect -88 59 0 127
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 140 627 244 640
rect 140 581 169 627
rect 215 581 244 627
rect 140 514 244 581
rect 140 468 169 514
rect 215 468 244 514
rect 140 401 244 468
rect 140 355 169 401
rect 215 355 244 401
rect 140 287 244 355
rect 140 241 169 287
rect 215 241 244 287
rect 140 173 244 241
rect 140 127 169 173
rect 215 127 244 173
rect 140 59 244 127
rect 140 13 169 59
rect 215 13 244 59
rect 140 0 244 13
rect 384 627 488 640
rect 384 581 413 627
rect 459 581 488 627
rect 384 514 488 581
rect 384 468 413 514
rect 459 468 488 514
rect 384 401 488 468
rect 384 355 413 401
rect 459 355 488 401
rect 384 287 488 355
rect 384 241 413 287
rect 459 241 488 287
rect 384 173 488 241
rect 384 127 413 173
rect 459 127 488 173
rect 384 59 488 127
rect 384 13 413 59
rect 459 13 488 59
rect 384 0 488 13
rect 628 627 732 640
rect 628 581 657 627
rect 703 581 732 627
rect 628 514 732 581
rect 628 468 657 514
rect 703 468 732 514
rect 628 401 732 468
rect 628 355 657 401
rect 703 355 732 401
rect 628 287 732 355
rect 628 241 657 287
rect 703 241 732 287
rect 628 173 732 241
rect 628 127 657 173
rect 703 127 732 173
rect 628 59 732 127
rect 628 13 657 59
rect 703 13 732 59
rect 628 0 732 13
rect 872 627 976 640
rect 872 581 901 627
rect 947 581 976 627
rect 872 514 976 581
rect 872 468 901 514
rect 947 468 976 514
rect 872 401 976 468
rect 872 355 901 401
rect 947 355 976 401
rect 872 287 976 355
rect 872 241 901 287
rect 947 241 976 287
rect 872 173 976 241
rect 872 127 901 173
rect 947 127 976 173
rect 872 59 976 127
rect 872 13 901 59
rect 947 13 976 59
rect 872 0 976 13
rect 1116 627 1204 640
rect 1116 581 1145 627
rect 1191 581 1204 627
rect 1116 514 1204 581
rect 1116 468 1145 514
rect 1191 468 1204 514
rect 1116 401 1204 468
rect 1116 355 1145 401
rect 1191 355 1204 401
rect 1116 287 1204 355
rect 1116 241 1145 287
rect 1191 241 1204 287
rect 1116 173 1204 241
rect 1116 127 1145 173
rect 1191 127 1204 173
rect 1116 59 1204 127
rect 1116 13 1145 59
rect 1191 13 1204 59
rect 1116 0 1204 13
<< mvndiffc >>
rect -75 581 -29 627
rect -75 468 -29 514
rect -75 355 -29 401
rect -75 241 -29 287
rect -75 127 -29 173
rect -75 13 -29 59
rect 169 581 215 627
rect 169 468 215 514
rect 169 355 215 401
rect 169 241 215 287
rect 169 127 215 173
rect 169 13 215 59
rect 413 581 459 627
rect 413 468 459 514
rect 413 355 459 401
rect 413 241 459 287
rect 413 127 459 173
rect 413 13 459 59
rect 657 581 703 627
rect 657 468 703 514
rect 657 355 703 401
rect 657 241 703 287
rect 657 127 703 173
rect 657 13 703 59
rect 901 581 947 627
rect 901 468 947 514
rect 901 355 947 401
rect 901 241 947 287
rect 901 127 947 173
rect 901 13 947 59
rect 1145 581 1191 627
rect 1145 468 1191 514
rect 1145 355 1191 401
rect 1145 241 1191 287
rect 1145 127 1191 173
rect 1145 13 1191 59
<< polysilicon >>
rect 0 640 140 684
rect 244 640 384 684
rect 488 640 628 684
rect 732 640 872 684
rect 976 640 1116 684
rect 0 -44 140 0
rect 244 -44 384 0
rect 488 -44 628 0
rect 732 -44 872 0
rect 976 -44 1116 0
<< metal1 >>
rect -75 627 -29 640
rect -75 514 -29 581
rect -75 401 -29 468
rect -75 287 -29 355
rect -75 173 -29 241
rect -75 59 -29 127
rect -75 0 -29 13
rect 169 627 215 640
rect 169 514 215 581
rect 169 401 215 468
rect 169 287 215 355
rect 169 173 215 241
rect 169 59 215 127
rect 169 0 215 13
rect 413 627 459 640
rect 413 514 459 581
rect 413 401 459 468
rect 413 287 459 355
rect 413 173 459 241
rect 413 59 459 127
rect 413 0 459 13
rect 657 627 703 640
rect 657 514 703 581
rect 657 401 703 468
rect 657 287 703 355
rect 657 173 703 241
rect 657 59 703 127
rect 657 0 703 13
rect 901 627 947 640
rect 901 514 947 581
rect 901 401 947 468
rect 901 287 947 355
rect 901 173 947 241
rect 901 59 947 127
rect 901 0 947 13
rect 1145 627 1191 640
rect 1145 514 1191 581
rect 1145 401 1191 468
rect 1145 287 1191 355
rect 1145 173 1191 241
rect 1145 59 1191 127
rect 1145 0 1191 13
<< labels >>
rlabel metal1 924 320 924 320 4 S
rlabel metal1 680 320 680 320 4 D
rlabel metal1 436 320 436 320 4 S
rlabel metal1 192 320 192 320 4 D
rlabel metal1 1168 320 1168 320 4 D
rlabel metal1 -52 320 -52 320 4 S
<< end >>
