magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1071 1019 1071
<< metal1 >>
rect -19 65 19 71
rect -19 -65 -13 65
rect 13 -65 19 65
rect -19 -71 19 -65
<< via1 >>
rect -13 -65 13 65
<< metal2 >>
rect -19 65 19 71
rect -19 -65 -13 65
rect 13 -65 19 65
rect -19 -71 19 -65
<< end >>
