magic
tech gf180mcuC
magscale 1 10
timestamp 1692614673
<< nwell >>
rect 0 -393 882 484
<< pwell >>
rect 0 -633 882 -435
<< nmos >>
rect 178 -559 234 -509
rect 346 -559 402 -509
rect 648 -559 704 -509
<< pmos >>
rect 178 136 234 186
rect 346 136 402 186
rect 648 136 704 186
rect 178 6 234 56
rect 346 6 402 56
rect 178 -127 234 -77
rect 346 -127 402 -77
rect 648 -127 704 -77
rect 178 -257 234 -207
rect 346 -257 402 -207
rect 648 -257 704 -207
<< ndiff >>
rect 86 -509 158 -498
rect 254 -509 326 -498
rect 422 -509 494 -498
rect 86 -511 178 -509
rect 86 -557 99 -511
rect 145 -557 178 -511
rect 86 -559 178 -557
rect 234 -511 346 -509
rect 234 -557 267 -511
rect 313 -557 346 -511
rect 234 -559 346 -557
rect 402 -511 494 -509
rect 402 -557 435 -511
rect 481 -557 494 -511
rect 402 -559 494 -557
rect 86 -570 158 -559
rect 254 -570 326 -559
rect 422 -570 494 -559
rect 556 -509 628 -498
rect 724 -509 796 -498
rect 556 -511 648 -509
rect 556 -557 569 -511
rect 615 -557 648 -511
rect 556 -559 648 -557
rect 704 -511 796 -509
rect 704 -557 737 -511
rect 783 -557 796 -511
rect 704 -559 796 -557
rect 556 -570 628 -559
rect 724 -570 796 -559
<< pdiff >>
rect 86 186 158 197
rect 254 186 326 197
rect 422 186 494 197
rect 86 184 178 186
rect 86 138 99 184
rect 145 138 178 184
rect 86 136 178 138
rect 234 184 346 186
rect 234 138 267 184
rect 313 138 346 184
rect 234 136 346 138
rect 402 184 494 186
rect 402 138 435 184
rect 481 138 494 184
rect 402 136 494 138
rect 86 125 158 136
rect 86 56 158 67
rect 254 125 326 136
rect 254 56 326 67
rect 422 125 494 136
rect 556 186 628 197
rect 724 186 796 197
rect 556 184 648 186
rect 556 138 569 184
rect 615 138 648 184
rect 556 136 648 138
rect 704 184 796 186
rect 704 138 737 184
rect 783 138 796 184
rect 704 136 796 138
rect 556 125 628 136
rect 724 125 796 136
rect 422 56 494 67
rect 86 54 178 56
rect 86 8 99 54
rect 145 8 178 54
rect 86 6 178 8
rect 234 54 346 56
rect 234 8 267 54
rect 313 8 346 54
rect 234 6 346 8
rect 402 54 494 56
rect 402 8 435 54
rect 481 8 494 54
rect 402 6 494 8
rect 86 -5 158 6
rect 86 -77 158 -66
rect 254 -5 326 6
rect 254 -77 326 -66
rect 422 -5 494 6
rect 422 -77 494 -66
rect 86 -79 178 -77
rect 86 -125 99 -79
rect 145 -125 178 -79
rect 86 -127 178 -125
rect 234 -79 346 -77
rect 234 -125 267 -79
rect 313 -125 346 -79
rect 234 -127 346 -125
rect 402 -79 494 -77
rect 402 -125 435 -79
rect 481 -125 494 -79
rect 402 -127 494 -125
rect 86 -138 158 -127
rect 86 -207 158 -196
rect 254 -138 326 -127
rect 254 -207 326 -196
rect 422 -138 494 -127
rect 556 -77 628 -66
rect 724 -77 796 -66
rect 556 -79 648 -77
rect 556 -125 569 -79
rect 615 -125 648 -79
rect 556 -127 648 -125
rect 704 -79 796 -77
rect 704 -125 737 -79
rect 783 -125 796 -79
rect 704 -127 796 -125
rect 556 -138 628 -127
rect 422 -207 494 -196
rect 86 -209 178 -207
rect 86 -255 99 -209
rect 145 -255 178 -209
rect 86 -257 178 -255
rect 234 -209 346 -207
rect 234 -255 267 -209
rect 313 -255 346 -209
rect 234 -257 346 -255
rect 402 -209 494 -207
rect 402 -255 435 -209
rect 481 -255 494 -209
rect 402 -257 494 -255
rect 86 -268 158 -257
rect 254 -268 326 -257
rect 422 -268 494 -257
rect 556 -207 628 -196
rect 724 -138 796 -127
rect 724 -207 796 -196
rect 556 -209 648 -207
rect 556 -255 569 -209
rect 615 -255 648 -209
rect 556 -257 648 -255
rect 704 -209 796 -207
rect 704 -255 737 -209
rect 783 -255 796 -209
rect 704 -257 796 -255
rect 556 -268 628 -257
rect 724 -268 796 -257
<< ndiffc >>
rect 99 -557 145 -511
rect 267 -557 313 -511
rect 435 -557 481 -511
rect 569 -557 615 -511
rect 737 -557 783 -511
<< pdiffc >>
rect 99 138 145 184
rect 267 138 313 184
rect 435 138 481 184
rect 569 138 615 184
rect 737 138 783 184
rect 99 8 145 54
rect 267 8 313 54
rect 435 8 481 54
rect 99 -125 145 -79
rect 267 -125 313 -79
rect 435 -125 481 -79
rect 569 -125 615 -79
rect 737 -125 783 -79
rect 99 -255 145 -209
rect 267 -255 313 -209
rect 435 -255 481 -209
rect 569 -255 615 -209
rect 737 -255 783 -209
<< psubdiff >>
rect 28 -683 854 -668
rect 28 -738 44 -683
rect 99 -738 167 -683
rect 222 -738 290 -683
rect 345 -738 413 -683
rect 468 -738 536 -683
rect 591 -738 659 -683
rect 714 -738 782 -683
rect 837 -738 854 -683
rect 28 -754 854 -738
<< nsubdiff >>
rect 28 441 854 456
rect 28 386 44 441
rect 99 386 167 441
rect 222 386 290 441
rect 345 386 413 441
rect 468 386 536 441
rect 591 386 659 441
rect 714 386 782 441
rect 837 386 854 441
rect 28 370 854 386
<< psubdiffcont >>
rect 44 -738 99 -683
rect 167 -738 222 -683
rect 290 -738 345 -683
rect 413 -738 468 -683
rect 536 -738 591 -683
rect 659 -738 714 -683
rect 782 -738 837 -683
<< nsubdiffcont >>
rect 44 386 99 441
rect 167 386 222 441
rect 290 386 345 441
rect 413 386 468 441
rect 536 386 591 441
rect 659 386 714 441
rect 782 386 837 441
<< polysilicon >>
rect 640 295 712 309
rect -31 274 41 283
rect -31 269 234 274
rect -31 223 -18 269
rect 28 223 234 269
rect 640 249 653 295
rect 699 249 712 295
rect 640 236 712 249
rect -31 218 234 223
rect -31 210 41 218
rect 178 186 234 218
rect 346 186 402 230
rect 178 56 234 136
rect 346 56 402 136
rect 648 186 704 236
rect 648 92 704 136
rect 178 -77 234 6
rect 346 -77 402 6
rect 178 -207 234 -127
rect 346 -207 402 -127
rect 648 -77 704 -33
rect 178 -509 234 -257
rect 346 -301 402 -257
rect 648 -207 704 -127
rect 311 -314 402 -301
rect 648 -302 704 -257
rect 311 -360 324 -314
rect 370 -360 402 -314
rect 311 -373 402 -360
rect 346 -509 402 -373
rect 607 -315 704 -302
rect 607 -361 620 -315
rect 666 -361 704 -315
rect 607 -374 704 -361
rect 178 -603 234 -559
rect 346 -603 402 -559
rect 648 -509 704 -374
rect 648 -603 704 -559
<< polycontact >>
rect -18 223 28 269
rect 653 249 699 295
rect 324 -360 370 -314
rect 620 -361 666 -315
<< metal1 >>
rect 14 441 868 470
rect 14 386 44 441
rect 99 386 167 441
rect 222 386 290 441
rect 345 386 413 441
rect 468 386 536 441
rect 591 386 659 441
rect 714 386 782 441
rect 837 386 868 441
rect 14 356 868 386
rect -31 269 41 283
rect -66 223 -18 269
rect 28 223 41 269
rect -31 210 41 223
rect 99 184 145 356
rect 653 309 699 356
rect 640 295 712 309
rect 569 249 653 295
rect 699 249 783 295
rect 569 236 783 249
rect 569 184 615 236
rect 737 184 783 236
rect 88 138 99 184
rect 145 138 156 184
rect 256 138 267 184
rect 313 138 324 184
rect 424 138 435 184
rect 481 138 492 184
rect 558 138 569 184
rect 615 138 626 184
rect 726 138 737 184
rect 783 138 794 184
rect 99 54 145 138
rect 267 54 313 138
rect 435 54 481 138
rect 88 8 99 54
rect 145 8 156 54
rect 256 8 267 54
rect 313 8 324 54
rect 424 8 435 54
rect 481 8 492 54
rect 99 -79 145 8
rect 267 -79 313 8
rect 435 -79 481 8
rect 569 -79 615 138
rect 737 -14 912 32
rect 737 -79 783 -14
rect 88 -125 99 -79
rect 145 -125 156 -79
rect 256 -125 267 -79
rect 313 -125 324 -79
rect 424 -125 435 -79
rect 481 -125 492 -79
rect 558 -125 569 -79
rect 615 -125 626 -79
rect 726 -125 737 -79
rect 783 -125 794 -79
rect 99 -209 145 -125
rect 267 -209 313 -125
rect 435 -209 481 -125
rect 569 -209 615 -125
rect 737 -209 783 -125
rect 88 -255 99 -209
rect 145 -255 156 -209
rect 256 -255 267 -209
rect 313 -255 324 -209
rect 424 -255 435 -209
rect 481 -255 492 -209
rect 558 -255 569 -209
rect 615 -255 626 -209
rect 726 -255 737 -209
rect 783 -255 794 -209
rect 311 -314 383 -301
rect -66 -360 324 -314
rect 370 -360 383 -314
rect 311 -373 383 -360
rect 435 -315 481 -255
rect 607 -315 679 -302
rect 435 -361 620 -315
rect 666 -361 679 -315
rect 435 -419 481 -361
rect 607 -374 679 -361
rect 99 -465 481 -419
rect 99 -511 145 -465
rect 435 -511 481 -465
rect 737 -511 783 -255
rect 88 -557 99 -511
rect 145 -557 156 -511
rect 256 -557 267 -511
rect 313 -557 324 -511
rect 424 -557 435 -511
rect 481 -557 492 -511
rect 558 -557 569 -511
rect 615 -557 626 -511
rect 726 -557 737 -511
rect 783 -557 794 -511
rect 267 -654 313 -557
rect 569 -654 615 -557
rect 14 -683 868 -654
rect 14 -738 44 -683
rect 99 -738 167 -683
rect 222 -738 290 -683
rect 345 -738 413 -683
rect 468 -738 536 -683
rect 591 -738 659 -683
rect 714 -738 782 -683
rect 837 -738 868 -683
rect 14 -768 868 -738
<< labels >>
flabel metal1 -63 244 -63 244 0 FreeSans 320 0 0 0 A
port 1 nsew
flabel metal1 -60 -333 -60 -333 0 FreeSans 320 0 0 0 B
port 2 nsew
flabel metal1 829 14 829 14 0 FreeSans 320 0 0 0 OUT
port 3 nsew
flabel nsubdiffcont 442 414 442 414 0 FreeSans 480 0 0 0 VDD
port 5 nsew
flabel psubdiffcont 442 -713 442 -713 0 FreeSans 480 0 0 0 VSS
port 7 nsew
<< end >>
