magic
tech gf180mcuC
magscale 1 10
timestamp 1694155625
<< nwell >>
rect -864 -957 864 957
<< nsubdiff >>
rect -840 920 840 933
rect -840 874 -724 920
rect 724 874 840 920
rect -840 861 840 874
rect -840 817 -768 861
rect -840 -817 -827 817
rect -781 -817 -768 817
rect 768 817 840 861
rect -840 -861 -768 -817
rect 768 -817 781 817
rect 827 -817 840 817
rect 768 -861 840 -817
rect -840 -874 840 -861
rect -840 -920 -724 -874
rect 724 -920 840 -874
rect -840 -933 840 -920
<< nsubdiffcont >>
rect -724 874 724 920
rect -827 -817 -781 817
rect 781 -817 827 817
rect -724 -920 724 -874
<< polysilicon >>
rect -680 760 -520 773
rect -680 714 -667 760
rect -533 714 -520 760
rect -680 670 -520 714
rect -680 -714 -520 -670
rect -680 -760 -667 -714
rect -533 -760 -520 -714
rect -680 -773 -520 -760
rect -440 760 -280 773
rect -440 714 -427 760
rect -293 714 -280 760
rect -440 670 -280 714
rect -440 -714 -280 -670
rect -440 -760 -427 -714
rect -293 -760 -280 -714
rect -440 -773 -280 -760
rect -200 760 -40 773
rect -200 714 -187 760
rect -53 714 -40 760
rect -200 670 -40 714
rect -200 -714 -40 -670
rect -200 -760 -187 -714
rect -53 -760 -40 -714
rect -200 -773 -40 -760
rect 40 760 200 773
rect 40 714 53 760
rect 187 714 200 760
rect 40 670 200 714
rect 40 -714 200 -670
rect 40 -760 53 -714
rect 187 -760 200 -714
rect 40 -773 200 -760
rect 280 760 440 773
rect 280 714 293 760
rect 427 714 440 760
rect 280 670 440 714
rect 280 -714 440 -670
rect 280 -760 293 -714
rect 427 -760 440 -714
rect 280 -773 440 -760
rect 520 760 680 773
rect 520 714 533 760
rect 667 714 680 760
rect 520 670 680 714
rect 520 -714 680 -670
rect 520 -760 533 -714
rect 667 -760 680 -714
rect 520 -773 680 -760
<< polycontact >>
rect -667 714 -533 760
rect -667 -760 -533 -714
rect -427 714 -293 760
rect -427 -760 -293 -714
rect -187 714 -53 760
rect -187 -760 -53 -714
rect 53 714 187 760
rect 53 -760 187 -714
rect 293 714 427 760
rect 293 -760 427 -714
rect 533 714 667 760
rect 533 -760 667 -714
<< ppolyres >>
rect -680 -670 -520 670
rect -440 -670 -280 670
rect -200 -670 -40 670
rect 40 -670 200 670
rect 280 -670 440 670
rect 520 -670 680 670
<< metal1 >>
rect -827 874 -724 920
rect 724 874 827 920
rect -827 817 -781 874
rect 781 817 827 874
rect -678 714 -667 760
rect -533 714 -522 760
rect -438 714 -427 760
rect -293 714 -282 760
rect -198 714 -187 760
rect -53 714 -42 760
rect 42 714 53 760
rect 187 714 198 760
rect 282 714 293 760
rect 427 714 438 760
rect 522 714 533 760
rect 667 714 678 760
rect -678 -760 -667 -714
rect -533 -760 -522 -714
rect -438 -760 -427 -714
rect -293 -760 -282 -714
rect -198 -760 -187 -714
rect -53 -760 -42 -714
rect 42 -760 53 -714
rect 187 -760 198 -714
rect 282 -760 293 -714
rect 427 -760 438 -714
rect 522 -760 533 -714
rect 667 -760 678 -714
rect -827 -874 -781 -817
rect 781 -874 827 -817
rect -827 -920 -724 -874
rect 724 -920 827 -874
<< properties >>
string FIXED_BBOX -804 -897 804 897
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 6.697 m 1 nx 6 wmin 0.80 lmin 1.00 rho 315 val 2.889k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1
<< end >>
