magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -7262 -2045 7262 2045
<< psubdiff >>
rect -5262 23 5262 45
rect -5262 -23 -5240 23
rect 5240 -23 5262 23
rect -5262 -45 5262 -23
<< psubdiffcont >>
rect -5240 -23 5240 23
<< metal1 >>
rect -5251 23 5251 34
rect -5251 -23 -5240 23
rect 5240 -23 5251 23
rect -5251 -34 5251 -23
<< end >>
