magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1745 -3560 1745 3560
<< metal3 >>
rect -745 2555 745 2560
rect -745 2527 -740 2555
rect -712 2527 -674 2555
rect -646 2527 -608 2555
rect -580 2527 -542 2555
rect -514 2527 -476 2555
rect -448 2527 -410 2555
rect -382 2527 -344 2555
rect -316 2527 -278 2555
rect -250 2527 -212 2555
rect -184 2527 -146 2555
rect -118 2527 -80 2555
rect -52 2527 -14 2555
rect 14 2527 52 2555
rect 80 2527 118 2555
rect 146 2527 184 2555
rect 212 2527 250 2555
rect 278 2527 316 2555
rect 344 2527 382 2555
rect 410 2527 448 2555
rect 476 2527 514 2555
rect 542 2527 580 2555
rect 608 2527 646 2555
rect 674 2527 712 2555
rect 740 2527 745 2555
rect -745 2489 745 2527
rect -745 2461 -740 2489
rect -712 2461 -674 2489
rect -646 2461 -608 2489
rect -580 2461 -542 2489
rect -514 2461 -476 2489
rect -448 2461 -410 2489
rect -382 2461 -344 2489
rect -316 2461 -278 2489
rect -250 2461 -212 2489
rect -184 2461 -146 2489
rect -118 2461 -80 2489
rect -52 2461 -14 2489
rect 14 2461 52 2489
rect 80 2461 118 2489
rect 146 2461 184 2489
rect 212 2461 250 2489
rect 278 2461 316 2489
rect 344 2461 382 2489
rect 410 2461 448 2489
rect 476 2461 514 2489
rect 542 2461 580 2489
rect 608 2461 646 2489
rect 674 2461 712 2489
rect 740 2461 745 2489
rect -745 2423 745 2461
rect -745 2395 -740 2423
rect -712 2395 -674 2423
rect -646 2395 -608 2423
rect -580 2395 -542 2423
rect -514 2395 -476 2423
rect -448 2395 -410 2423
rect -382 2395 -344 2423
rect -316 2395 -278 2423
rect -250 2395 -212 2423
rect -184 2395 -146 2423
rect -118 2395 -80 2423
rect -52 2395 -14 2423
rect 14 2395 52 2423
rect 80 2395 118 2423
rect 146 2395 184 2423
rect 212 2395 250 2423
rect 278 2395 316 2423
rect 344 2395 382 2423
rect 410 2395 448 2423
rect 476 2395 514 2423
rect 542 2395 580 2423
rect 608 2395 646 2423
rect 674 2395 712 2423
rect 740 2395 745 2423
rect -745 2357 745 2395
rect -745 2329 -740 2357
rect -712 2329 -674 2357
rect -646 2329 -608 2357
rect -580 2329 -542 2357
rect -514 2329 -476 2357
rect -448 2329 -410 2357
rect -382 2329 -344 2357
rect -316 2329 -278 2357
rect -250 2329 -212 2357
rect -184 2329 -146 2357
rect -118 2329 -80 2357
rect -52 2329 -14 2357
rect 14 2329 52 2357
rect 80 2329 118 2357
rect 146 2329 184 2357
rect 212 2329 250 2357
rect 278 2329 316 2357
rect 344 2329 382 2357
rect 410 2329 448 2357
rect 476 2329 514 2357
rect 542 2329 580 2357
rect 608 2329 646 2357
rect 674 2329 712 2357
rect 740 2329 745 2357
rect -745 2291 745 2329
rect -745 2263 -740 2291
rect -712 2263 -674 2291
rect -646 2263 -608 2291
rect -580 2263 -542 2291
rect -514 2263 -476 2291
rect -448 2263 -410 2291
rect -382 2263 -344 2291
rect -316 2263 -278 2291
rect -250 2263 -212 2291
rect -184 2263 -146 2291
rect -118 2263 -80 2291
rect -52 2263 -14 2291
rect 14 2263 52 2291
rect 80 2263 118 2291
rect 146 2263 184 2291
rect 212 2263 250 2291
rect 278 2263 316 2291
rect 344 2263 382 2291
rect 410 2263 448 2291
rect 476 2263 514 2291
rect 542 2263 580 2291
rect 608 2263 646 2291
rect 674 2263 712 2291
rect 740 2263 745 2291
rect -745 2225 745 2263
rect -745 2197 -740 2225
rect -712 2197 -674 2225
rect -646 2197 -608 2225
rect -580 2197 -542 2225
rect -514 2197 -476 2225
rect -448 2197 -410 2225
rect -382 2197 -344 2225
rect -316 2197 -278 2225
rect -250 2197 -212 2225
rect -184 2197 -146 2225
rect -118 2197 -80 2225
rect -52 2197 -14 2225
rect 14 2197 52 2225
rect 80 2197 118 2225
rect 146 2197 184 2225
rect 212 2197 250 2225
rect 278 2197 316 2225
rect 344 2197 382 2225
rect 410 2197 448 2225
rect 476 2197 514 2225
rect 542 2197 580 2225
rect 608 2197 646 2225
rect 674 2197 712 2225
rect 740 2197 745 2225
rect -745 2159 745 2197
rect -745 2131 -740 2159
rect -712 2131 -674 2159
rect -646 2131 -608 2159
rect -580 2131 -542 2159
rect -514 2131 -476 2159
rect -448 2131 -410 2159
rect -382 2131 -344 2159
rect -316 2131 -278 2159
rect -250 2131 -212 2159
rect -184 2131 -146 2159
rect -118 2131 -80 2159
rect -52 2131 -14 2159
rect 14 2131 52 2159
rect 80 2131 118 2159
rect 146 2131 184 2159
rect 212 2131 250 2159
rect 278 2131 316 2159
rect 344 2131 382 2159
rect 410 2131 448 2159
rect 476 2131 514 2159
rect 542 2131 580 2159
rect 608 2131 646 2159
rect 674 2131 712 2159
rect 740 2131 745 2159
rect -745 2093 745 2131
rect -745 2065 -740 2093
rect -712 2065 -674 2093
rect -646 2065 -608 2093
rect -580 2065 -542 2093
rect -514 2065 -476 2093
rect -448 2065 -410 2093
rect -382 2065 -344 2093
rect -316 2065 -278 2093
rect -250 2065 -212 2093
rect -184 2065 -146 2093
rect -118 2065 -80 2093
rect -52 2065 -14 2093
rect 14 2065 52 2093
rect 80 2065 118 2093
rect 146 2065 184 2093
rect 212 2065 250 2093
rect 278 2065 316 2093
rect 344 2065 382 2093
rect 410 2065 448 2093
rect 476 2065 514 2093
rect 542 2065 580 2093
rect 608 2065 646 2093
rect 674 2065 712 2093
rect 740 2065 745 2093
rect -745 2027 745 2065
rect -745 1999 -740 2027
rect -712 1999 -674 2027
rect -646 1999 -608 2027
rect -580 1999 -542 2027
rect -514 1999 -476 2027
rect -448 1999 -410 2027
rect -382 1999 -344 2027
rect -316 1999 -278 2027
rect -250 1999 -212 2027
rect -184 1999 -146 2027
rect -118 1999 -80 2027
rect -52 1999 -14 2027
rect 14 1999 52 2027
rect 80 1999 118 2027
rect 146 1999 184 2027
rect 212 1999 250 2027
rect 278 1999 316 2027
rect 344 1999 382 2027
rect 410 1999 448 2027
rect 476 1999 514 2027
rect 542 1999 580 2027
rect 608 1999 646 2027
rect 674 1999 712 2027
rect 740 1999 745 2027
rect -745 1961 745 1999
rect -745 1933 -740 1961
rect -712 1933 -674 1961
rect -646 1933 -608 1961
rect -580 1933 -542 1961
rect -514 1933 -476 1961
rect -448 1933 -410 1961
rect -382 1933 -344 1961
rect -316 1933 -278 1961
rect -250 1933 -212 1961
rect -184 1933 -146 1961
rect -118 1933 -80 1961
rect -52 1933 -14 1961
rect 14 1933 52 1961
rect 80 1933 118 1961
rect 146 1933 184 1961
rect 212 1933 250 1961
rect 278 1933 316 1961
rect 344 1933 382 1961
rect 410 1933 448 1961
rect 476 1933 514 1961
rect 542 1933 580 1961
rect 608 1933 646 1961
rect 674 1933 712 1961
rect 740 1933 745 1961
rect -745 1895 745 1933
rect -745 1867 -740 1895
rect -712 1867 -674 1895
rect -646 1867 -608 1895
rect -580 1867 -542 1895
rect -514 1867 -476 1895
rect -448 1867 -410 1895
rect -382 1867 -344 1895
rect -316 1867 -278 1895
rect -250 1867 -212 1895
rect -184 1867 -146 1895
rect -118 1867 -80 1895
rect -52 1867 -14 1895
rect 14 1867 52 1895
rect 80 1867 118 1895
rect 146 1867 184 1895
rect 212 1867 250 1895
rect 278 1867 316 1895
rect 344 1867 382 1895
rect 410 1867 448 1895
rect 476 1867 514 1895
rect 542 1867 580 1895
rect 608 1867 646 1895
rect 674 1867 712 1895
rect 740 1867 745 1895
rect -745 1829 745 1867
rect -745 1801 -740 1829
rect -712 1801 -674 1829
rect -646 1801 -608 1829
rect -580 1801 -542 1829
rect -514 1801 -476 1829
rect -448 1801 -410 1829
rect -382 1801 -344 1829
rect -316 1801 -278 1829
rect -250 1801 -212 1829
rect -184 1801 -146 1829
rect -118 1801 -80 1829
rect -52 1801 -14 1829
rect 14 1801 52 1829
rect 80 1801 118 1829
rect 146 1801 184 1829
rect 212 1801 250 1829
rect 278 1801 316 1829
rect 344 1801 382 1829
rect 410 1801 448 1829
rect 476 1801 514 1829
rect 542 1801 580 1829
rect 608 1801 646 1829
rect 674 1801 712 1829
rect 740 1801 745 1829
rect -745 1763 745 1801
rect -745 1735 -740 1763
rect -712 1735 -674 1763
rect -646 1735 -608 1763
rect -580 1735 -542 1763
rect -514 1735 -476 1763
rect -448 1735 -410 1763
rect -382 1735 -344 1763
rect -316 1735 -278 1763
rect -250 1735 -212 1763
rect -184 1735 -146 1763
rect -118 1735 -80 1763
rect -52 1735 -14 1763
rect 14 1735 52 1763
rect 80 1735 118 1763
rect 146 1735 184 1763
rect 212 1735 250 1763
rect 278 1735 316 1763
rect 344 1735 382 1763
rect 410 1735 448 1763
rect 476 1735 514 1763
rect 542 1735 580 1763
rect 608 1735 646 1763
rect 674 1735 712 1763
rect 740 1735 745 1763
rect -745 1697 745 1735
rect -745 1669 -740 1697
rect -712 1669 -674 1697
rect -646 1669 -608 1697
rect -580 1669 -542 1697
rect -514 1669 -476 1697
rect -448 1669 -410 1697
rect -382 1669 -344 1697
rect -316 1669 -278 1697
rect -250 1669 -212 1697
rect -184 1669 -146 1697
rect -118 1669 -80 1697
rect -52 1669 -14 1697
rect 14 1669 52 1697
rect 80 1669 118 1697
rect 146 1669 184 1697
rect 212 1669 250 1697
rect 278 1669 316 1697
rect 344 1669 382 1697
rect 410 1669 448 1697
rect 476 1669 514 1697
rect 542 1669 580 1697
rect 608 1669 646 1697
rect 674 1669 712 1697
rect 740 1669 745 1697
rect -745 1631 745 1669
rect -745 1603 -740 1631
rect -712 1603 -674 1631
rect -646 1603 -608 1631
rect -580 1603 -542 1631
rect -514 1603 -476 1631
rect -448 1603 -410 1631
rect -382 1603 -344 1631
rect -316 1603 -278 1631
rect -250 1603 -212 1631
rect -184 1603 -146 1631
rect -118 1603 -80 1631
rect -52 1603 -14 1631
rect 14 1603 52 1631
rect 80 1603 118 1631
rect 146 1603 184 1631
rect 212 1603 250 1631
rect 278 1603 316 1631
rect 344 1603 382 1631
rect 410 1603 448 1631
rect 476 1603 514 1631
rect 542 1603 580 1631
rect 608 1603 646 1631
rect 674 1603 712 1631
rect 740 1603 745 1631
rect -745 1565 745 1603
rect -745 1537 -740 1565
rect -712 1537 -674 1565
rect -646 1537 -608 1565
rect -580 1537 -542 1565
rect -514 1537 -476 1565
rect -448 1537 -410 1565
rect -382 1537 -344 1565
rect -316 1537 -278 1565
rect -250 1537 -212 1565
rect -184 1537 -146 1565
rect -118 1537 -80 1565
rect -52 1537 -14 1565
rect 14 1537 52 1565
rect 80 1537 118 1565
rect 146 1537 184 1565
rect 212 1537 250 1565
rect 278 1537 316 1565
rect 344 1537 382 1565
rect 410 1537 448 1565
rect 476 1537 514 1565
rect 542 1537 580 1565
rect 608 1537 646 1565
rect 674 1537 712 1565
rect 740 1537 745 1565
rect -745 1499 745 1537
rect -745 1471 -740 1499
rect -712 1471 -674 1499
rect -646 1471 -608 1499
rect -580 1471 -542 1499
rect -514 1471 -476 1499
rect -448 1471 -410 1499
rect -382 1471 -344 1499
rect -316 1471 -278 1499
rect -250 1471 -212 1499
rect -184 1471 -146 1499
rect -118 1471 -80 1499
rect -52 1471 -14 1499
rect 14 1471 52 1499
rect 80 1471 118 1499
rect 146 1471 184 1499
rect 212 1471 250 1499
rect 278 1471 316 1499
rect 344 1471 382 1499
rect 410 1471 448 1499
rect 476 1471 514 1499
rect 542 1471 580 1499
rect 608 1471 646 1499
rect 674 1471 712 1499
rect 740 1471 745 1499
rect -745 1433 745 1471
rect -745 1405 -740 1433
rect -712 1405 -674 1433
rect -646 1405 -608 1433
rect -580 1405 -542 1433
rect -514 1405 -476 1433
rect -448 1405 -410 1433
rect -382 1405 -344 1433
rect -316 1405 -278 1433
rect -250 1405 -212 1433
rect -184 1405 -146 1433
rect -118 1405 -80 1433
rect -52 1405 -14 1433
rect 14 1405 52 1433
rect 80 1405 118 1433
rect 146 1405 184 1433
rect 212 1405 250 1433
rect 278 1405 316 1433
rect 344 1405 382 1433
rect 410 1405 448 1433
rect 476 1405 514 1433
rect 542 1405 580 1433
rect 608 1405 646 1433
rect 674 1405 712 1433
rect 740 1405 745 1433
rect -745 1367 745 1405
rect -745 1339 -740 1367
rect -712 1339 -674 1367
rect -646 1339 -608 1367
rect -580 1339 -542 1367
rect -514 1339 -476 1367
rect -448 1339 -410 1367
rect -382 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 382 1367
rect 410 1339 448 1367
rect 476 1339 514 1367
rect 542 1339 580 1367
rect 608 1339 646 1367
rect 674 1339 712 1367
rect 740 1339 745 1367
rect -745 1301 745 1339
rect -745 1273 -740 1301
rect -712 1273 -674 1301
rect -646 1273 -608 1301
rect -580 1273 -542 1301
rect -514 1273 -476 1301
rect -448 1273 -410 1301
rect -382 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 382 1301
rect 410 1273 448 1301
rect 476 1273 514 1301
rect 542 1273 580 1301
rect 608 1273 646 1301
rect 674 1273 712 1301
rect 740 1273 745 1301
rect -745 1235 745 1273
rect -745 1207 -740 1235
rect -712 1207 -674 1235
rect -646 1207 -608 1235
rect -580 1207 -542 1235
rect -514 1207 -476 1235
rect -448 1207 -410 1235
rect -382 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 382 1235
rect 410 1207 448 1235
rect 476 1207 514 1235
rect 542 1207 580 1235
rect 608 1207 646 1235
rect 674 1207 712 1235
rect 740 1207 745 1235
rect -745 1169 745 1207
rect -745 1141 -740 1169
rect -712 1141 -674 1169
rect -646 1141 -608 1169
rect -580 1141 -542 1169
rect -514 1141 -476 1169
rect -448 1141 -410 1169
rect -382 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 382 1169
rect 410 1141 448 1169
rect 476 1141 514 1169
rect 542 1141 580 1169
rect 608 1141 646 1169
rect 674 1141 712 1169
rect 740 1141 745 1169
rect -745 1103 745 1141
rect -745 1075 -740 1103
rect -712 1075 -674 1103
rect -646 1075 -608 1103
rect -580 1075 -542 1103
rect -514 1075 -476 1103
rect -448 1075 -410 1103
rect -382 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 382 1103
rect 410 1075 448 1103
rect 476 1075 514 1103
rect 542 1075 580 1103
rect 608 1075 646 1103
rect 674 1075 712 1103
rect 740 1075 745 1103
rect -745 1037 745 1075
rect -745 1009 -740 1037
rect -712 1009 -674 1037
rect -646 1009 -608 1037
rect -580 1009 -542 1037
rect -514 1009 -476 1037
rect -448 1009 -410 1037
rect -382 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 382 1037
rect 410 1009 448 1037
rect 476 1009 514 1037
rect 542 1009 580 1037
rect 608 1009 646 1037
rect 674 1009 712 1037
rect 740 1009 745 1037
rect -745 971 745 1009
rect -745 943 -740 971
rect -712 943 -674 971
rect -646 943 -608 971
rect -580 943 -542 971
rect -514 943 -476 971
rect -448 943 -410 971
rect -382 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 382 971
rect 410 943 448 971
rect 476 943 514 971
rect 542 943 580 971
rect 608 943 646 971
rect 674 943 712 971
rect 740 943 745 971
rect -745 905 745 943
rect -745 877 -740 905
rect -712 877 -674 905
rect -646 877 -608 905
rect -580 877 -542 905
rect -514 877 -476 905
rect -448 877 -410 905
rect -382 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 382 905
rect 410 877 448 905
rect 476 877 514 905
rect 542 877 580 905
rect 608 877 646 905
rect 674 877 712 905
rect 740 877 745 905
rect -745 839 745 877
rect -745 811 -740 839
rect -712 811 -674 839
rect -646 811 -608 839
rect -580 811 -542 839
rect -514 811 -476 839
rect -448 811 -410 839
rect -382 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 382 839
rect 410 811 448 839
rect 476 811 514 839
rect 542 811 580 839
rect 608 811 646 839
rect 674 811 712 839
rect 740 811 745 839
rect -745 773 745 811
rect -745 745 -740 773
rect -712 745 -674 773
rect -646 745 -608 773
rect -580 745 -542 773
rect -514 745 -476 773
rect -448 745 -410 773
rect -382 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 382 773
rect 410 745 448 773
rect 476 745 514 773
rect 542 745 580 773
rect 608 745 646 773
rect 674 745 712 773
rect 740 745 745 773
rect -745 707 745 745
rect -745 679 -740 707
rect -712 679 -674 707
rect -646 679 -608 707
rect -580 679 -542 707
rect -514 679 -476 707
rect -448 679 -410 707
rect -382 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 382 707
rect 410 679 448 707
rect 476 679 514 707
rect 542 679 580 707
rect 608 679 646 707
rect 674 679 712 707
rect 740 679 745 707
rect -745 641 745 679
rect -745 613 -740 641
rect -712 613 -674 641
rect -646 613 -608 641
rect -580 613 -542 641
rect -514 613 -476 641
rect -448 613 -410 641
rect -382 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 382 641
rect 410 613 448 641
rect 476 613 514 641
rect 542 613 580 641
rect 608 613 646 641
rect 674 613 712 641
rect 740 613 745 641
rect -745 575 745 613
rect -745 547 -740 575
rect -712 547 -674 575
rect -646 547 -608 575
rect -580 547 -542 575
rect -514 547 -476 575
rect -448 547 -410 575
rect -382 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 382 575
rect 410 547 448 575
rect 476 547 514 575
rect 542 547 580 575
rect 608 547 646 575
rect 674 547 712 575
rect 740 547 745 575
rect -745 509 745 547
rect -745 481 -740 509
rect -712 481 -674 509
rect -646 481 -608 509
rect -580 481 -542 509
rect -514 481 -476 509
rect -448 481 -410 509
rect -382 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 382 509
rect 410 481 448 509
rect 476 481 514 509
rect 542 481 580 509
rect 608 481 646 509
rect 674 481 712 509
rect 740 481 745 509
rect -745 443 745 481
rect -745 415 -740 443
rect -712 415 -674 443
rect -646 415 -608 443
rect -580 415 -542 443
rect -514 415 -476 443
rect -448 415 -410 443
rect -382 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 382 443
rect 410 415 448 443
rect 476 415 514 443
rect 542 415 580 443
rect 608 415 646 443
rect 674 415 712 443
rect 740 415 745 443
rect -745 377 745 415
rect -745 349 -740 377
rect -712 349 -674 377
rect -646 349 -608 377
rect -580 349 -542 377
rect -514 349 -476 377
rect -448 349 -410 377
rect -382 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 382 377
rect 410 349 448 377
rect 476 349 514 377
rect 542 349 580 377
rect 608 349 646 377
rect 674 349 712 377
rect 740 349 745 377
rect -745 311 745 349
rect -745 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 745 311
rect -745 245 745 283
rect -745 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 745 245
rect -745 179 745 217
rect -745 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 745 179
rect -745 113 745 151
rect -745 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 745 113
rect -745 47 745 85
rect -745 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 745 47
rect -745 -19 745 19
rect -745 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 745 -19
rect -745 -85 745 -47
rect -745 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 745 -85
rect -745 -151 745 -113
rect -745 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 745 -151
rect -745 -217 745 -179
rect -745 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 745 -217
rect -745 -283 745 -245
rect -745 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 745 -283
rect -745 -349 745 -311
rect -745 -377 -740 -349
rect -712 -377 -674 -349
rect -646 -377 -608 -349
rect -580 -377 -542 -349
rect -514 -377 -476 -349
rect -448 -377 -410 -349
rect -382 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 382 -349
rect 410 -377 448 -349
rect 476 -377 514 -349
rect 542 -377 580 -349
rect 608 -377 646 -349
rect 674 -377 712 -349
rect 740 -377 745 -349
rect -745 -415 745 -377
rect -745 -443 -740 -415
rect -712 -443 -674 -415
rect -646 -443 -608 -415
rect -580 -443 -542 -415
rect -514 -443 -476 -415
rect -448 -443 -410 -415
rect -382 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 382 -415
rect 410 -443 448 -415
rect 476 -443 514 -415
rect 542 -443 580 -415
rect 608 -443 646 -415
rect 674 -443 712 -415
rect 740 -443 745 -415
rect -745 -481 745 -443
rect -745 -509 -740 -481
rect -712 -509 -674 -481
rect -646 -509 -608 -481
rect -580 -509 -542 -481
rect -514 -509 -476 -481
rect -448 -509 -410 -481
rect -382 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 382 -481
rect 410 -509 448 -481
rect 476 -509 514 -481
rect 542 -509 580 -481
rect 608 -509 646 -481
rect 674 -509 712 -481
rect 740 -509 745 -481
rect -745 -547 745 -509
rect -745 -575 -740 -547
rect -712 -575 -674 -547
rect -646 -575 -608 -547
rect -580 -575 -542 -547
rect -514 -575 -476 -547
rect -448 -575 -410 -547
rect -382 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 382 -547
rect 410 -575 448 -547
rect 476 -575 514 -547
rect 542 -575 580 -547
rect 608 -575 646 -547
rect 674 -575 712 -547
rect 740 -575 745 -547
rect -745 -613 745 -575
rect -745 -641 -740 -613
rect -712 -641 -674 -613
rect -646 -641 -608 -613
rect -580 -641 -542 -613
rect -514 -641 -476 -613
rect -448 -641 -410 -613
rect -382 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 382 -613
rect 410 -641 448 -613
rect 476 -641 514 -613
rect 542 -641 580 -613
rect 608 -641 646 -613
rect 674 -641 712 -613
rect 740 -641 745 -613
rect -745 -679 745 -641
rect -745 -707 -740 -679
rect -712 -707 -674 -679
rect -646 -707 -608 -679
rect -580 -707 -542 -679
rect -514 -707 -476 -679
rect -448 -707 -410 -679
rect -382 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 382 -679
rect 410 -707 448 -679
rect 476 -707 514 -679
rect 542 -707 580 -679
rect 608 -707 646 -679
rect 674 -707 712 -679
rect 740 -707 745 -679
rect -745 -745 745 -707
rect -745 -773 -740 -745
rect -712 -773 -674 -745
rect -646 -773 -608 -745
rect -580 -773 -542 -745
rect -514 -773 -476 -745
rect -448 -773 -410 -745
rect -382 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 382 -745
rect 410 -773 448 -745
rect 476 -773 514 -745
rect 542 -773 580 -745
rect 608 -773 646 -745
rect 674 -773 712 -745
rect 740 -773 745 -745
rect -745 -811 745 -773
rect -745 -839 -740 -811
rect -712 -839 -674 -811
rect -646 -839 -608 -811
rect -580 -839 -542 -811
rect -514 -839 -476 -811
rect -448 -839 -410 -811
rect -382 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 382 -811
rect 410 -839 448 -811
rect 476 -839 514 -811
rect 542 -839 580 -811
rect 608 -839 646 -811
rect 674 -839 712 -811
rect 740 -839 745 -811
rect -745 -877 745 -839
rect -745 -905 -740 -877
rect -712 -905 -674 -877
rect -646 -905 -608 -877
rect -580 -905 -542 -877
rect -514 -905 -476 -877
rect -448 -905 -410 -877
rect -382 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 382 -877
rect 410 -905 448 -877
rect 476 -905 514 -877
rect 542 -905 580 -877
rect 608 -905 646 -877
rect 674 -905 712 -877
rect 740 -905 745 -877
rect -745 -943 745 -905
rect -745 -971 -740 -943
rect -712 -971 -674 -943
rect -646 -971 -608 -943
rect -580 -971 -542 -943
rect -514 -971 -476 -943
rect -448 -971 -410 -943
rect -382 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 382 -943
rect 410 -971 448 -943
rect 476 -971 514 -943
rect 542 -971 580 -943
rect 608 -971 646 -943
rect 674 -971 712 -943
rect 740 -971 745 -943
rect -745 -1009 745 -971
rect -745 -1037 -740 -1009
rect -712 -1037 -674 -1009
rect -646 -1037 -608 -1009
rect -580 -1037 -542 -1009
rect -514 -1037 -476 -1009
rect -448 -1037 -410 -1009
rect -382 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 382 -1009
rect 410 -1037 448 -1009
rect 476 -1037 514 -1009
rect 542 -1037 580 -1009
rect 608 -1037 646 -1009
rect 674 -1037 712 -1009
rect 740 -1037 745 -1009
rect -745 -1075 745 -1037
rect -745 -1103 -740 -1075
rect -712 -1103 -674 -1075
rect -646 -1103 -608 -1075
rect -580 -1103 -542 -1075
rect -514 -1103 -476 -1075
rect -448 -1103 -410 -1075
rect -382 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 382 -1075
rect 410 -1103 448 -1075
rect 476 -1103 514 -1075
rect 542 -1103 580 -1075
rect 608 -1103 646 -1075
rect 674 -1103 712 -1075
rect 740 -1103 745 -1075
rect -745 -1141 745 -1103
rect -745 -1169 -740 -1141
rect -712 -1169 -674 -1141
rect -646 -1169 -608 -1141
rect -580 -1169 -542 -1141
rect -514 -1169 -476 -1141
rect -448 -1169 -410 -1141
rect -382 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 382 -1141
rect 410 -1169 448 -1141
rect 476 -1169 514 -1141
rect 542 -1169 580 -1141
rect 608 -1169 646 -1141
rect 674 -1169 712 -1141
rect 740 -1169 745 -1141
rect -745 -1207 745 -1169
rect -745 -1235 -740 -1207
rect -712 -1235 -674 -1207
rect -646 -1235 -608 -1207
rect -580 -1235 -542 -1207
rect -514 -1235 -476 -1207
rect -448 -1235 -410 -1207
rect -382 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 382 -1207
rect 410 -1235 448 -1207
rect 476 -1235 514 -1207
rect 542 -1235 580 -1207
rect 608 -1235 646 -1207
rect 674 -1235 712 -1207
rect 740 -1235 745 -1207
rect -745 -1273 745 -1235
rect -745 -1301 -740 -1273
rect -712 -1301 -674 -1273
rect -646 -1301 -608 -1273
rect -580 -1301 -542 -1273
rect -514 -1301 -476 -1273
rect -448 -1301 -410 -1273
rect -382 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 382 -1273
rect 410 -1301 448 -1273
rect 476 -1301 514 -1273
rect 542 -1301 580 -1273
rect 608 -1301 646 -1273
rect 674 -1301 712 -1273
rect 740 -1301 745 -1273
rect -745 -1339 745 -1301
rect -745 -1367 -740 -1339
rect -712 -1367 -674 -1339
rect -646 -1367 -608 -1339
rect -580 -1367 -542 -1339
rect -514 -1367 -476 -1339
rect -448 -1367 -410 -1339
rect -382 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 382 -1339
rect 410 -1367 448 -1339
rect 476 -1367 514 -1339
rect 542 -1367 580 -1339
rect 608 -1367 646 -1339
rect 674 -1367 712 -1339
rect 740 -1367 745 -1339
rect -745 -1405 745 -1367
rect -745 -1433 -740 -1405
rect -712 -1433 -674 -1405
rect -646 -1433 -608 -1405
rect -580 -1433 -542 -1405
rect -514 -1433 -476 -1405
rect -448 -1433 -410 -1405
rect -382 -1433 -344 -1405
rect -316 -1433 -278 -1405
rect -250 -1433 -212 -1405
rect -184 -1433 -146 -1405
rect -118 -1433 -80 -1405
rect -52 -1433 -14 -1405
rect 14 -1433 52 -1405
rect 80 -1433 118 -1405
rect 146 -1433 184 -1405
rect 212 -1433 250 -1405
rect 278 -1433 316 -1405
rect 344 -1433 382 -1405
rect 410 -1433 448 -1405
rect 476 -1433 514 -1405
rect 542 -1433 580 -1405
rect 608 -1433 646 -1405
rect 674 -1433 712 -1405
rect 740 -1433 745 -1405
rect -745 -1471 745 -1433
rect -745 -1499 -740 -1471
rect -712 -1499 -674 -1471
rect -646 -1499 -608 -1471
rect -580 -1499 -542 -1471
rect -514 -1499 -476 -1471
rect -448 -1499 -410 -1471
rect -382 -1499 -344 -1471
rect -316 -1499 -278 -1471
rect -250 -1499 -212 -1471
rect -184 -1499 -146 -1471
rect -118 -1499 -80 -1471
rect -52 -1499 -14 -1471
rect 14 -1499 52 -1471
rect 80 -1499 118 -1471
rect 146 -1499 184 -1471
rect 212 -1499 250 -1471
rect 278 -1499 316 -1471
rect 344 -1499 382 -1471
rect 410 -1499 448 -1471
rect 476 -1499 514 -1471
rect 542 -1499 580 -1471
rect 608 -1499 646 -1471
rect 674 -1499 712 -1471
rect 740 -1499 745 -1471
rect -745 -1537 745 -1499
rect -745 -1565 -740 -1537
rect -712 -1565 -674 -1537
rect -646 -1565 -608 -1537
rect -580 -1565 -542 -1537
rect -514 -1565 -476 -1537
rect -448 -1565 -410 -1537
rect -382 -1565 -344 -1537
rect -316 -1565 -278 -1537
rect -250 -1565 -212 -1537
rect -184 -1565 -146 -1537
rect -118 -1565 -80 -1537
rect -52 -1565 -14 -1537
rect 14 -1565 52 -1537
rect 80 -1565 118 -1537
rect 146 -1565 184 -1537
rect 212 -1565 250 -1537
rect 278 -1565 316 -1537
rect 344 -1565 382 -1537
rect 410 -1565 448 -1537
rect 476 -1565 514 -1537
rect 542 -1565 580 -1537
rect 608 -1565 646 -1537
rect 674 -1565 712 -1537
rect 740 -1565 745 -1537
rect -745 -1603 745 -1565
rect -745 -1631 -740 -1603
rect -712 -1631 -674 -1603
rect -646 -1631 -608 -1603
rect -580 -1631 -542 -1603
rect -514 -1631 -476 -1603
rect -448 -1631 -410 -1603
rect -382 -1631 -344 -1603
rect -316 -1631 -278 -1603
rect -250 -1631 -212 -1603
rect -184 -1631 -146 -1603
rect -118 -1631 -80 -1603
rect -52 -1631 -14 -1603
rect 14 -1631 52 -1603
rect 80 -1631 118 -1603
rect 146 -1631 184 -1603
rect 212 -1631 250 -1603
rect 278 -1631 316 -1603
rect 344 -1631 382 -1603
rect 410 -1631 448 -1603
rect 476 -1631 514 -1603
rect 542 -1631 580 -1603
rect 608 -1631 646 -1603
rect 674 -1631 712 -1603
rect 740 -1631 745 -1603
rect -745 -1669 745 -1631
rect -745 -1697 -740 -1669
rect -712 -1697 -674 -1669
rect -646 -1697 -608 -1669
rect -580 -1697 -542 -1669
rect -514 -1697 -476 -1669
rect -448 -1697 -410 -1669
rect -382 -1697 -344 -1669
rect -316 -1697 -278 -1669
rect -250 -1697 -212 -1669
rect -184 -1697 -146 -1669
rect -118 -1697 -80 -1669
rect -52 -1697 -14 -1669
rect 14 -1697 52 -1669
rect 80 -1697 118 -1669
rect 146 -1697 184 -1669
rect 212 -1697 250 -1669
rect 278 -1697 316 -1669
rect 344 -1697 382 -1669
rect 410 -1697 448 -1669
rect 476 -1697 514 -1669
rect 542 -1697 580 -1669
rect 608 -1697 646 -1669
rect 674 -1697 712 -1669
rect 740 -1697 745 -1669
rect -745 -1735 745 -1697
rect -745 -1763 -740 -1735
rect -712 -1763 -674 -1735
rect -646 -1763 -608 -1735
rect -580 -1763 -542 -1735
rect -514 -1763 -476 -1735
rect -448 -1763 -410 -1735
rect -382 -1763 -344 -1735
rect -316 -1763 -278 -1735
rect -250 -1763 -212 -1735
rect -184 -1763 -146 -1735
rect -118 -1763 -80 -1735
rect -52 -1763 -14 -1735
rect 14 -1763 52 -1735
rect 80 -1763 118 -1735
rect 146 -1763 184 -1735
rect 212 -1763 250 -1735
rect 278 -1763 316 -1735
rect 344 -1763 382 -1735
rect 410 -1763 448 -1735
rect 476 -1763 514 -1735
rect 542 -1763 580 -1735
rect 608 -1763 646 -1735
rect 674 -1763 712 -1735
rect 740 -1763 745 -1735
rect -745 -1801 745 -1763
rect -745 -1829 -740 -1801
rect -712 -1829 -674 -1801
rect -646 -1829 -608 -1801
rect -580 -1829 -542 -1801
rect -514 -1829 -476 -1801
rect -448 -1829 -410 -1801
rect -382 -1829 -344 -1801
rect -316 -1829 -278 -1801
rect -250 -1829 -212 -1801
rect -184 -1829 -146 -1801
rect -118 -1829 -80 -1801
rect -52 -1829 -14 -1801
rect 14 -1829 52 -1801
rect 80 -1829 118 -1801
rect 146 -1829 184 -1801
rect 212 -1829 250 -1801
rect 278 -1829 316 -1801
rect 344 -1829 382 -1801
rect 410 -1829 448 -1801
rect 476 -1829 514 -1801
rect 542 -1829 580 -1801
rect 608 -1829 646 -1801
rect 674 -1829 712 -1801
rect 740 -1829 745 -1801
rect -745 -1867 745 -1829
rect -745 -1895 -740 -1867
rect -712 -1895 -674 -1867
rect -646 -1895 -608 -1867
rect -580 -1895 -542 -1867
rect -514 -1895 -476 -1867
rect -448 -1895 -410 -1867
rect -382 -1895 -344 -1867
rect -316 -1895 -278 -1867
rect -250 -1895 -212 -1867
rect -184 -1895 -146 -1867
rect -118 -1895 -80 -1867
rect -52 -1895 -14 -1867
rect 14 -1895 52 -1867
rect 80 -1895 118 -1867
rect 146 -1895 184 -1867
rect 212 -1895 250 -1867
rect 278 -1895 316 -1867
rect 344 -1895 382 -1867
rect 410 -1895 448 -1867
rect 476 -1895 514 -1867
rect 542 -1895 580 -1867
rect 608 -1895 646 -1867
rect 674 -1895 712 -1867
rect 740 -1895 745 -1867
rect -745 -1933 745 -1895
rect -745 -1961 -740 -1933
rect -712 -1961 -674 -1933
rect -646 -1961 -608 -1933
rect -580 -1961 -542 -1933
rect -514 -1961 -476 -1933
rect -448 -1961 -410 -1933
rect -382 -1961 -344 -1933
rect -316 -1961 -278 -1933
rect -250 -1961 -212 -1933
rect -184 -1961 -146 -1933
rect -118 -1961 -80 -1933
rect -52 -1961 -14 -1933
rect 14 -1961 52 -1933
rect 80 -1961 118 -1933
rect 146 -1961 184 -1933
rect 212 -1961 250 -1933
rect 278 -1961 316 -1933
rect 344 -1961 382 -1933
rect 410 -1961 448 -1933
rect 476 -1961 514 -1933
rect 542 -1961 580 -1933
rect 608 -1961 646 -1933
rect 674 -1961 712 -1933
rect 740 -1961 745 -1933
rect -745 -1999 745 -1961
rect -745 -2027 -740 -1999
rect -712 -2027 -674 -1999
rect -646 -2027 -608 -1999
rect -580 -2027 -542 -1999
rect -514 -2027 -476 -1999
rect -448 -2027 -410 -1999
rect -382 -2027 -344 -1999
rect -316 -2027 -278 -1999
rect -250 -2027 -212 -1999
rect -184 -2027 -146 -1999
rect -118 -2027 -80 -1999
rect -52 -2027 -14 -1999
rect 14 -2027 52 -1999
rect 80 -2027 118 -1999
rect 146 -2027 184 -1999
rect 212 -2027 250 -1999
rect 278 -2027 316 -1999
rect 344 -2027 382 -1999
rect 410 -2027 448 -1999
rect 476 -2027 514 -1999
rect 542 -2027 580 -1999
rect 608 -2027 646 -1999
rect 674 -2027 712 -1999
rect 740 -2027 745 -1999
rect -745 -2065 745 -2027
rect -745 -2093 -740 -2065
rect -712 -2093 -674 -2065
rect -646 -2093 -608 -2065
rect -580 -2093 -542 -2065
rect -514 -2093 -476 -2065
rect -448 -2093 -410 -2065
rect -382 -2093 -344 -2065
rect -316 -2093 -278 -2065
rect -250 -2093 -212 -2065
rect -184 -2093 -146 -2065
rect -118 -2093 -80 -2065
rect -52 -2093 -14 -2065
rect 14 -2093 52 -2065
rect 80 -2093 118 -2065
rect 146 -2093 184 -2065
rect 212 -2093 250 -2065
rect 278 -2093 316 -2065
rect 344 -2093 382 -2065
rect 410 -2093 448 -2065
rect 476 -2093 514 -2065
rect 542 -2093 580 -2065
rect 608 -2093 646 -2065
rect 674 -2093 712 -2065
rect 740 -2093 745 -2065
rect -745 -2131 745 -2093
rect -745 -2159 -740 -2131
rect -712 -2159 -674 -2131
rect -646 -2159 -608 -2131
rect -580 -2159 -542 -2131
rect -514 -2159 -476 -2131
rect -448 -2159 -410 -2131
rect -382 -2159 -344 -2131
rect -316 -2159 -278 -2131
rect -250 -2159 -212 -2131
rect -184 -2159 -146 -2131
rect -118 -2159 -80 -2131
rect -52 -2159 -14 -2131
rect 14 -2159 52 -2131
rect 80 -2159 118 -2131
rect 146 -2159 184 -2131
rect 212 -2159 250 -2131
rect 278 -2159 316 -2131
rect 344 -2159 382 -2131
rect 410 -2159 448 -2131
rect 476 -2159 514 -2131
rect 542 -2159 580 -2131
rect 608 -2159 646 -2131
rect 674 -2159 712 -2131
rect 740 -2159 745 -2131
rect -745 -2197 745 -2159
rect -745 -2225 -740 -2197
rect -712 -2225 -674 -2197
rect -646 -2225 -608 -2197
rect -580 -2225 -542 -2197
rect -514 -2225 -476 -2197
rect -448 -2225 -410 -2197
rect -382 -2225 -344 -2197
rect -316 -2225 -278 -2197
rect -250 -2225 -212 -2197
rect -184 -2225 -146 -2197
rect -118 -2225 -80 -2197
rect -52 -2225 -14 -2197
rect 14 -2225 52 -2197
rect 80 -2225 118 -2197
rect 146 -2225 184 -2197
rect 212 -2225 250 -2197
rect 278 -2225 316 -2197
rect 344 -2225 382 -2197
rect 410 -2225 448 -2197
rect 476 -2225 514 -2197
rect 542 -2225 580 -2197
rect 608 -2225 646 -2197
rect 674 -2225 712 -2197
rect 740 -2225 745 -2197
rect -745 -2263 745 -2225
rect -745 -2291 -740 -2263
rect -712 -2291 -674 -2263
rect -646 -2291 -608 -2263
rect -580 -2291 -542 -2263
rect -514 -2291 -476 -2263
rect -448 -2291 -410 -2263
rect -382 -2291 -344 -2263
rect -316 -2291 -278 -2263
rect -250 -2291 -212 -2263
rect -184 -2291 -146 -2263
rect -118 -2291 -80 -2263
rect -52 -2291 -14 -2263
rect 14 -2291 52 -2263
rect 80 -2291 118 -2263
rect 146 -2291 184 -2263
rect 212 -2291 250 -2263
rect 278 -2291 316 -2263
rect 344 -2291 382 -2263
rect 410 -2291 448 -2263
rect 476 -2291 514 -2263
rect 542 -2291 580 -2263
rect 608 -2291 646 -2263
rect 674 -2291 712 -2263
rect 740 -2291 745 -2263
rect -745 -2329 745 -2291
rect -745 -2357 -740 -2329
rect -712 -2357 -674 -2329
rect -646 -2357 -608 -2329
rect -580 -2357 -542 -2329
rect -514 -2357 -476 -2329
rect -448 -2357 -410 -2329
rect -382 -2357 -344 -2329
rect -316 -2357 -278 -2329
rect -250 -2357 -212 -2329
rect -184 -2357 -146 -2329
rect -118 -2357 -80 -2329
rect -52 -2357 -14 -2329
rect 14 -2357 52 -2329
rect 80 -2357 118 -2329
rect 146 -2357 184 -2329
rect 212 -2357 250 -2329
rect 278 -2357 316 -2329
rect 344 -2357 382 -2329
rect 410 -2357 448 -2329
rect 476 -2357 514 -2329
rect 542 -2357 580 -2329
rect 608 -2357 646 -2329
rect 674 -2357 712 -2329
rect 740 -2357 745 -2329
rect -745 -2395 745 -2357
rect -745 -2423 -740 -2395
rect -712 -2423 -674 -2395
rect -646 -2423 -608 -2395
rect -580 -2423 -542 -2395
rect -514 -2423 -476 -2395
rect -448 -2423 -410 -2395
rect -382 -2423 -344 -2395
rect -316 -2423 -278 -2395
rect -250 -2423 -212 -2395
rect -184 -2423 -146 -2395
rect -118 -2423 -80 -2395
rect -52 -2423 -14 -2395
rect 14 -2423 52 -2395
rect 80 -2423 118 -2395
rect 146 -2423 184 -2395
rect 212 -2423 250 -2395
rect 278 -2423 316 -2395
rect 344 -2423 382 -2395
rect 410 -2423 448 -2395
rect 476 -2423 514 -2395
rect 542 -2423 580 -2395
rect 608 -2423 646 -2395
rect 674 -2423 712 -2395
rect 740 -2423 745 -2395
rect -745 -2461 745 -2423
rect -745 -2489 -740 -2461
rect -712 -2489 -674 -2461
rect -646 -2489 -608 -2461
rect -580 -2489 -542 -2461
rect -514 -2489 -476 -2461
rect -448 -2489 -410 -2461
rect -382 -2489 -344 -2461
rect -316 -2489 -278 -2461
rect -250 -2489 -212 -2461
rect -184 -2489 -146 -2461
rect -118 -2489 -80 -2461
rect -52 -2489 -14 -2461
rect 14 -2489 52 -2461
rect 80 -2489 118 -2461
rect 146 -2489 184 -2461
rect 212 -2489 250 -2461
rect 278 -2489 316 -2461
rect 344 -2489 382 -2461
rect 410 -2489 448 -2461
rect 476 -2489 514 -2461
rect 542 -2489 580 -2461
rect 608 -2489 646 -2461
rect 674 -2489 712 -2461
rect 740 -2489 745 -2461
rect -745 -2527 745 -2489
rect -745 -2555 -740 -2527
rect -712 -2555 -674 -2527
rect -646 -2555 -608 -2527
rect -580 -2555 -542 -2527
rect -514 -2555 -476 -2527
rect -448 -2555 -410 -2527
rect -382 -2555 -344 -2527
rect -316 -2555 -278 -2527
rect -250 -2555 -212 -2527
rect -184 -2555 -146 -2527
rect -118 -2555 -80 -2527
rect -52 -2555 -14 -2527
rect 14 -2555 52 -2527
rect 80 -2555 118 -2527
rect 146 -2555 184 -2527
rect 212 -2555 250 -2527
rect 278 -2555 316 -2527
rect 344 -2555 382 -2527
rect 410 -2555 448 -2527
rect 476 -2555 514 -2527
rect 542 -2555 580 -2527
rect 608 -2555 646 -2527
rect 674 -2555 712 -2527
rect 740 -2555 745 -2527
rect -745 -2560 745 -2555
<< via3 >>
rect -740 2527 -712 2555
rect -674 2527 -646 2555
rect -608 2527 -580 2555
rect -542 2527 -514 2555
rect -476 2527 -448 2555
rect -410 2527 -382 2555
rect -344 2527 -316 2555
rect -278 2527 -250 2555
rect -212 2527 -184 2555
rect -146 2527 -118 2555
rect -80 2527 -52 2555
rect -14 2527 14 2555
rect 52 2527 80 2555
rect 118 2527 146 2555
rect 184 2527 212 2555
rect 250 2527 278 2555
rect 316 2527 344 2555
rect 382 2527 410 2555
rect 448 2527 476 2555
rect 514 2527 542 2555
rect 580 2527 608 2555
rect 646 2527 674 2555
rect 712 2527 740 2555
rect -740 2461 -712 2489
rect -674 2461 -646 2489
rect -608 2461 -580 2489
rect -542 2461 -514 2489
rect -476 2461 -448 2489
rect -410 2461 -382 2489
rect -344 2461 -316 2489
rect -278 2461 -250 2489
rect -212 2461 -184 2489
rect -146 2461 -118 2489
rect -80 2461 -52 2489
rect -14 2461 14 2489
rect 52 2461 80 2489
rect 118 2461 146 2489
rect 184 2461 212 2489
rect 250 2461 278 2489
rect 316 2461 344 2489
rect 382 2461 410 2489
rect 448 2461 476 2489
rect 514 2461 542 2489
rect 580 2461 608 2489
rect 646 2461 674 2489
rect 712 2461 740 2489
rect -740 2395 -712 2423
rect -674 2395 -646 2423
rect -608 2395 -580 2423
rect -542 2395 -514 2423
rect -476 2395 -448 2423
rect -410 2395 -382 2423
rect -344 2395 -316 2423
rect -278 2395 -250 2423
rect -212 2395 -184 2423
rect -146 2395 -118 2423
rect -80 2395 -52 2423
rect -14 2395 14 2423
rect 52 2395 80 2423
rect 118 2395 146 2423
rect 184 2395 212 2423
rect 250 2395 278 2423
rect 316 2395 344 2423
rect 382 2395 410 2423
rect 448 2395 476 2423
rect 514 2395 542 2423
rect 580 2395 608 2423
rect 646 2395 674 2423
rect 712 2395 740 2423
rect -740 2329 -712 2357
rect -674 2329 -646 2357
rect -608 2329 -580 2357
rect -542 2329 -514 2357
rect -476 2329 -448 2357
rect -410 2329 -382 2357
rect -344 2329 -316 2357
rect -278 2329 -250 2357
rect -212 2329 -184 2357
rect -146 2329 -118 2357
rect -80 2329 -52 2357
rect -14 2329 14 2357
rect 52 2329 80 2357
rect 118 2329 146 2357
rect 184 2329 212 2357
rect 250 2329 278 2357
rect 316 2329 344 2357
rect 382 2329 410 2357
rect 448 2329 476 2357
rect 514 2329 542 2357
rect 580 2329 608 2357
rect 646 2329 674 2357
rect 712 2329 740 2357
rect -740 2263 -712 2291
rect -674 2263 -646 2291
rect -608 2263 -580 2291
rect -542 2263 -514 2291
rect -476 2263 -448 2291
rect -410 2263 -382 2291
rect -344 2263 -316 2291
rect -278 2263 -250 2291
rect -212 2263 -184 2291
rect -146 2263 -118 2291
rect -80 2263 -52 2291
rect -14 2263 14 2291
rect 52 2263 80 2291
rect 118 2263 146 2291
rect 184 2263 212 2291
rect 250 2263 278 2291
rect 316 2263 344 2291
rect 382 2263 410 2291
rect 448 2263 476 2291
rect 514 2263 542 2291
rect 580 2263 608 2291
rect 646 2263 674 2291
rect 712 2263 740 2291
rect -740 2197 -712 2225
rect -674 2197 -646 2225
rect -608 2197 -580 2225
rect -542 2197 -514 2225
rect -476 2197 -448 2225
rect -410 2197 -382 2225
rect -344 2197 -316 2225
rect -278 2197 -250 2225
rect -212 2197 -184 2225
rect -146 2197 -118 2225
rect -80 2197 -52 2225
rect -14 2197 14 2225
rect 52 2197 80 2225
rect 118 2197 146 2225
rect 184 2197 212 2225
rect 250 2197 278 2225
rect 316 2197 344 2225
rect 382 2197 410 2225
rect 448 2197 476 2225
rect 514 2197 542 2225
rect 580 2197 608 2225
rect 646 2197 674 2225
rect 712 2197 740 2225
rect -740 2131 -712 2159
rect -674 2131 -646 2159
rect -608 2131 -580 2159
rect -542 2131 -514 2159
rect -476 2131 -448 2159
rect -410 2131 -382 2159
rect -344 2131 -316 2159
rect -278 2131 -250 2159
rect -212 2131 -184 2159
rect -146 2131 -118 2159
rect -80 2131 -52 2159
rect -14 2131 14 2159
rect 52 2131 80 2159
rect 118 2131 146 2159
rect 184 2131 212 2159
rect 250 2131 278 2159
rect 316 2131 344 2159
rect 382 2131 410 2159
rect 448 2131 476 2159
rect 514 2131 542 2159
rect 580 2131 608 2159
rect 646 2131 674 2159
rect 712 2131 740 2159
rect -740 2065 -712 2093
rect -674 2065 -646 2093
rect -608 2065 -580 2093
rect -542 2065 -514 2093
rect -476 2065 -448 2093
rect -410 2065 -382 2093
rect -344 2065 -316 2093
rect -278 2065 -250 2093
rect -212 2065 -184 2093
rect -146 2065 -118 2093
rect -80 2065 -52 2093
rect -14 2065 14 2093
rect 52 2065 80 2093
rect 118 2065 146 2093
rect 184 2065 212 2093
rect 250 2065 278 2093
rect 316 2065 344 2093
rect 382 2065 410 2093
rect 448 2065 476 2093
rect 514 2065 542 2093
rect 580 2065 608 2093
rect 646 2065 674 2093
rect 712 2065 740 2093
rect -740 1999 -712 2027
rect -674 1999 -646 2027
rect -608 1999 -580 2027
rect -542 1999 -514 2027
rect -476 1999 -448 2027
rect -410 1999 -382 2027
rect -344 1999 -316 2027
rect -278 1999 -250 2027
rect -212 1999 -184 2027
rect -146 1999 -118 2027
rect -80 1999 -52 2027
rect -14 1999 14 2027
rect 52 1999 80 2027
rect 118 1999 146 2027
rect 184 1999 212 2027
rect 250 1999 278 2027
rect 316 1999 344 2027
rect 382 1999 410 2027
rect 448 1999 476 2027
rect 514 1999 542 2027
rect 580 1999 608 2027
rect 646 1999 674 2027
rect 712 1999 740 2027
rect -740 1933 -712 1961
rect -674 1933 -646 1961
rect -608 1933 -580 1961
rect -542 1933 -514 1961
rect -476 1933 -448 1961
rect -410 1933 -382 1961
rect -344 1933 -316 1961
rect -278 1933 -250 1961
rect -212 1933 -184 1961
rect -146 1933 -118 1961
rect -80 1933 -52 1961
rect -14 1933 14 1961
rect 52 1933 80 1961
rect 118 1933 146 1961
rect 184 1933 212 1961
rect 250 1933 278 1961
rect 316 1933 344 1961
rect 382 1933 410 1961
rect 448 1933 476 1961
rect 514 1933 542 1961
rect 580 1933 608 1961
rect 646 1933 674 1961
rect 712 1933 740 1961
rect -740 1867 -712 1895
rect -674 1867 -646 1895
rect -608 1867 -580 1895
rect -542 1867 -514 1895
rect -476 1867 -448 1895
rect -410 1867 -382 1895
rect -344 1867 -316 1895
rect -278 1867 -250 1895
rect -212 1867 -184 1895
rect -146 1867 -118 1895
rect -80 1867 -52 1895
rect -14 1867 14 1895
rect 52 1867 80 1895
rect 118 1867 146 1895
rect 184 1867 212 1895
rect 250 1867 278 1895
rect 316 1867 344 1895
rect 382 1867 410 1895
rect 448 1867 476 1895
rect 514 1867 542 1895
rect 580 1867 608 1895
rect 646 1867 674 1895
rect 712 1867 740 1895
rect -740 1801 -712 1829
rect -674 1801 -646 1829
rect -608 1801 -580 1829
rect -542 1801 -514 1829
rect -476 1801 -448 1829
rect -410 1801 -382 1829
rect -344 1801 -316 1829
rect -278 1801 -250 1829
rect -212 1801 -184 1829
rect -146 1801 -118 1829
rect -80 1801 -52 1829
rect -14 1801 14 1829
rect 52 1801 80 1829
rect 118 1801 146 1829
rect 184 1801 212 1829
rect 250 1801 278 1829
rect 316 1801 344 1829
rect 382 1801 410 1829
rect 448 1801 476 1829
rect 514 1801 542 1829
rect 580 1801 608 1829
rect 646 1801 674 1829
rect 712 1801 740 1829
rect -740 1735 -712 1763
rect -674 1735 -646 1763
rect -608 1735 -580 1763
rect -542 1735 -514 1763
rect -476 1735 -448 1763
rect -410 1735 -382 1763
rect -344 1735 -316 1763
rect -278 1735 -250 1763
rect -212 1735 -184 1763
rect -146 1735 -118 1763
rect -80 1735 -52 1763
rect -14 1735 14 1763
rect 52 1735 80 1763
rect 118 1735 146 1763
rect 184 1735 212 1763
rect 250 1735 278 1763
rect 316 1735 344 1763
rect 382 1735 410 1763
rect 448 1735 476 1763
rect 514 1735 542 1763
rect 580 1735 608 1763
rect 646 1735 674 1763
rect 712 1735 740 1763
rect -740 1669 -712 1697
rect -674 1669 -646 1697
rect -608 1669 -580 1697
rect -542 1669 -514 1697
rect -476 1669 -448 1697
rect -410 1669 -382 1697
rect -344 1669 -316 1697
rect -278 1669 -250 1697
rect -212 1669 -184 1697
rect -146 1669 -118 1697
rect -80 1669 -52 1697
rect -14 1669 14 1697
rect 52 1669 80 1697
rect 118 1669 146 1697
rect 184 1669 212 1697
rect 250 1669 278 1697
rect 316 1669 344 1697
rect 382 1669 410 1697
rect 448 1669 476 1697
rect 514 1669 542 1697
rect 580 1669 608 1697
rect 646 1669 674 1697
rect 712 1669 740 1697
rect -740 1603 -712 1631
rect -674 1603 -646 1631
rect -608 1603 -580 1631
rect -542 1603 -514 1631
rect -476 1603 -448 1631
rect -410 1603 -382 1631
rect -344 1603 -316 1631
rect -278 1603 -250 1631
rect -212 1603 -184 1631
rect -146 1603 -118 1631
rect -80 1603 -52 1631
rect -14 1603 14 1631
rect 52 1603 80 1631
rect 118 1603 146 1631
rect 184 1603 212 1631
rect 250 1603 278 1631
rect 316 1603 344 1631
rect 382 1603 410 1631
rect 448 1603 476 1631
rect 514 1603 542 1631
rect 580 1603 608 1631
rect 646 1603 674 1631
rect 712 1603 740 1631
rect -740 1537 -712 1565
rect -674 1537 -646 1565
rect -608 1537 -580 1565
rect -542 1537 -514 1565
rect -476 1537 -448 1565
rect -410 1537 -382 1565
rect -344 1537 -316 1565
rect -278 1537 -250 1565
rect -212 1537 -184 1565
rect -146 1537 -118 1565
rect -80 1537 -52 1565
rect -14 1537 14 1565
rect 52 1537 80 1565
rect 118 1537 146 1565
rect 184 1537 212 1565
rect 250 1537 278 1565
rect 316 1537 344 1565
rect 382 1537 410 1565
rect 448 1537 476 1565
rect 514 1537 542 1565
rect 580 1537 608 1565
rect 646 1537 674 1565
rect 712 1537 740 1565
rect -740 1471 -712 1499
rect -674 1471 -646 1499
rect -608 1471 -580 1499
rect -542 1471 -514 1499
rect -476 1471 -448 1499
rect -410 1471 -382 1499
rect -344 1471 -316 1499
rect -278 1471 -250 1499
rect -212 1471 -184 1499
rect -146 1471 -118 1499
rect -80 1471 -52 1499
rect -14 1471 14 1499
rect 52 1471 80 1499
rect 118 1471 146 1499
rect 184 1471 212 1499
rect 250 1471 278 1499
rect 316 1471 344 1499
rect 382 1471 410 1499
rect 448 1471 476 1499
rect 514 1471 542 1499
rect 580 1471 608 1499
rect 646 1471 674 1499
rect 712 1471 740 1499
rect -740 1405 -712 1433
rect -674 1405 -646 1433
rect -608 1405 -580 1433
rect -542 1405 -514 1433
rect -476 1405 -448 1433
rect -410 1405 -382 1433
rect -344 1405 -316 1433
rect -278 1405 -250 1433
rect -212 1405 -184 1433
rect -146 1405 -118 1433
rect -80 1405 -52 1433
rect -14 1405 14 1433
rect 52 1405 80 1433
rect 118 1405 146 1433
rect 184 1405 212 1433
rect 250 1405 278 1433
rect 316 1405 344 1433
rect 382 1405 410 1433
rect 448 1405 476 1433
rect 514 1405 542 1433
rect 580 1405 608 1433
rect 646 1405 674 1433
rect 712 1405 740 1433
rect -740 1339 -712 1367
rect -674 1339 -646 1367
rect -608 1339 -580 1367
rect -542 1339 -514 1367
rect -476 1339 -448 1367
rect -410 1339 -382 1367
rect -344 1339 -316 1367
rect -278 1339 -250 1367
rect -212 1339 -184 1367
rect -146 1339 -118 1367
rect -80 1339 -52 1367
rect -14 1339 14 1367
rect 52 1339 80 1367
rect 118 1339 146 1367
rect 184 1339 212 1367
rect 250 1339 278 1367
rect 316 1339 344 1367
rect 382 1339 410 1367
rect 448 1339 476 1367
rect 514 1339 542 1367
rect 580 1339 608 1367
rect 646 1339 674 1367
rect 712 1339 740 1367
rect -740 1273 -712 1301
rect -674 1273 -646 1301
rect -608 1273 -580 1301
rect -542 1273 -514 1301
rect -476 1273 -448 1301
rect -410 1273 -382 1301
rect -344 1273 -316 1301
rect -278 1273 -250 1301
rect -212 1273 -184 1301
rect -146 1273 -118 1301
rect -80 1273 -52 1301
rect -14 1273 14 1301
rect 52 1273 80 1301
rect 118 1273 146 1301
rect 184 1273 212 1301
rect 250 1273 278 1301
rect 316 1273 344 1301
rect 382 1273 410 1301
rect 448 1273 476 1301
rect 514 1273 542 1301
rect 580 1273 608 1301
rect 646 1273 674 1301
rect 712 1273 740 1301
rect -740 1207 -712 1235
rect -674 1207 -646 1235
rect -608 1207 -580 1235
rect -542 1207 -514 1235
rect -476 1207 -448 1235
rect -410 1207 -382 1235
rect -344 1207 -316 1235
rect -278 1207 -250 1235
rect -212 1207 -184 1235
rect -146 1207 -118 1235
rect -80 1207 -52 1235
rect -14 1207 14 1235
rect 52 1207 80 1235
rect 118 1207 146 1235
rect 184 1207 212 1235
rect 250 1207 278 1235
rect 316 1207 344 1235
rect 382 1207 410 1235
rect 448 1207 476 1235
rect 514 1207 542 1235
rect 580 1207 608 1235
rect 646 1207 674 1235
rect 712 1207 740 1235
rect -740 1141 -712 1169
rect -674 1141 -646 1169
rect -608 1141 -580 1169
rect -542 1141 -514 1169
rect -476 1141 -448 1169
rect -410 1141 -382 1169
rect -344 1141 -316 1169
rect -278 1141 -250 1169
rect -212 1141 -184 1169
rect -146 1141 -118 1169
rect -80 1141 -52 1169
rect -14 1141 14 1169
rect 52 1141 80 1169
rect 118 1141 146 1169
rect 184 1141 212 1169
rect 250 1141 278 1169
rect 316 1141 344 1169
rect 382 1141 410 1169
rect 448 1141 476 1169
rect 514 1141 542 1169
rect 580 1141 608 1169
rect 646 1141 674 1169
rect 712 1141 740 1169
rect -740 1075 -712 1103
rect -674 1075 -646 1103
rect -608 1075 -580 1103
rect -542 1075 -514 1103
rect -476 1075 -448 1103
rect -410 1075 -382 1103
rect -344 1075 -316 1103
rect -278 1075 -250 1103
rect -212 1075 -184 1103
rect -146 1075 -118 1103
rect -80 1075 -52 1103
rect -14 1075 14 1103
rect 52 1075 80 1103
rect 118 1075 146 1103
rect 184 1075 212 1103
rect 250 1075 278 1103
rect 316 1075 344 1103
rect 382 1075 410 1103
rect 448 1075 476 1103
rect 514 1075 542 1103
rect 580 1075 608 1103
rect 646 1075 674 1103
rect 712 1075 740 1103
rect -740 1009 -712 1037
rect -674 1009 -646 1037
rect -608 1009 -580 1037
rect -542 1009 -514 1037
rect -476 1009 -448 1037
rect -410 1009 -382 1037
rect -344 1009 -316 1037
rect -278 1009 -250 1037
rect -212 1009 -184 1037
rect -146 1009 -118 1037
rect -80 1009 -52 1037
rect -14 1009 14 1037
rect 52 1009 80 1037
rect 118 1009 146 1037
rect 184 1009 212 1037
rect 250 1009 278 1037
rect 316 1009 344 1037
rect 382 1009 410 1037
rect 448 1009 476 1037
rect 514 1009 542 1037
rect 580 1009 608 1037
rect 646 1009 674 1037
rect 712 1009 740 1037
rect -740 943 -712 971
rect -674 943 -646 971
rect -608 943 -580 971
rect -542 943 -514 971
rect -476 943 -448 971
rect -410 943 -382 971
rect -344 943 -316 971
rect -278 943 -250 971
rect -212 943 -184 971
rect -146 943 -118 971
rect -80 943 -52 971
rect -14 943 14 971
rect 52 943 80 971
rect 118 943 146 971
rect 184 943 212 971
rect 250 943 278 971
rect 316 943 344 971
rect 382 943 410 971
rect 448 943 476 971
rect 514 943 542 971
rect 580 943 608 971
rect 646 943 674 971
rect 712 943 740 971
rect -740 877 -712 905
rect -674 877 -646 905
rect -608 877 -580 905
rect -542 877 -514 905
rect -476 877 -448 905
rect -410 877 -382 905
rect -344 877 -316 905
rect -278 877 -250 905
rect -212 877 -184 905
rect -146 877 -118 905
rect -80 877 -52 905
rect -14 877 14 905
rect 52 877 80 905
rect 118 877 146 905
rect 184 877 212 905
rect 250 877 278 905
rect 316 877 344 905
rect 382 877 410 905
rect 448 877 476 905
rect 514 877 542 905
rect 580 877 608 905
rect 646 877 674 905
rect 712 877 740 905
rect -740 811 -712 839
rect -674 811 -646 839
rect -608 811 -580 839
rect -542 811 -514 839
rect -476 811 -448 839
rect -410 811 -382 839
rect -344 811 -316 839
rect -278 811 -250 839
rect -212 811 -184 839
rect -146 811 -118 839
rect -80 811 -52 839
rect -14 811 14 839
rect 52 811 80 839
rect 118 811 146 839
rect 184 811 212 839
rect 250 811 278 839
rect 316 811 344 839
rect 382 811 410 839
rect 448 811 476 839
rect 514 811 542 839
rect 580 811 608 839
rect 646 811 674 839
rect 712 811 740 839
rect -740 745 -712 773
rect -674 745 -646 773
rect -608 745 -580 773
rect -542 745 -514 773
rect -476 745 -448 773
rect -410 745 -382 773
rect -344 745 -316 773
rect -278 745 -250 773
rect -212 745 -184 773
rect -146 745 -118 773
rect -80 745 -52 773
rect -14 745 14 773
rect 52 745 80 773
rect 118 745 146 773
rect 184 745 212 773
rect 250 745 278 773
rect 316 745 344 773
rect 382 745 410 773
rect 448 745 476 773
rect 514 745 542 773
rect 580 745 608 773
rect 646 745 674 773
rect 712 745 740 773
rect -740 679 -712 707
rect -674 679 -646 707
rect -608 679 -580 707
rect -542 679 -514 707
rect -476 679 -448 707
rect -410 679 -382 707
rect -344 679 -316 707
rect -278 679 -250 707
rect -212 679 -184 707
rect -146 679 -118 707
rect -80 679 -52 707
rect -14 679 14 707
rect 52 679 80 707
rect 118 679 146 707
rect 184 679 212 707
rect 250 679 278 707
rect 316 679 344 707
rect 382 679 410 707
rect 448 679 476 707
rect 514 679 542 707
rect 580 679 608 707
rect 646 679 674 707
rect 712 679 740 707
rect -740 613 -712 641
rect -674 613 -646 641
rect -608 613 -580 641
rect -542 613 -514 641
rect -476 613 -448 641
rect -410 613 -382 641
rect -344 613 -316 641
rect -278 613 -250 641
rect -212 613 -184 641
rect -146 613 -118 641
rect -80 613 -52 641
rect -14 613 14 641
rect 52 613 80 641
rect 118 613 146 641
rect 184 613 212 641
rect 250 613 278 641
rect 316 613 344 641
rect 382 613 410 641
rect 448 613 476 641
rect 514 613 542 641
rect 580 613 608 641
rect 646 613 674 641
rect 712 613 740 641
rect -740 547 -712 575
rect -674 547 -646 575
rect -608 547 -580 575
rect -542 547 -514 575
rect -476 547 -448 575
rect -410 547 -382 575
rect -344 547 -316 575
rect -278 547 -250 575
rect -212 547 -184 575
rect -146 547 -118 575
rect -80 547 -52 575
rect -14 547 14 575
rect 52 547 80 575
rect 118 547 146 575
rect 184 547 212 575
rect 250 547 278 575
rect 316 547 344 575
rect 382 547 410 575
rect 448 547 476 575
rect 514 547 542 575
rect 580 547 608 575
rect 646 547 674 575
rect 712 547 740 575
rect -740 481 -712 509
rect -674 481 -646 509
rect -608 481 -580 509
rect -542 481 -514 509
rect -476 481 -448 509
rect -410 481 -382 509
rect -344 481 -316 509
rect -278 481 -250 509
rect -212 481 -184 509
rect -146 481 -118 509
rect -80 481 -52 509
rect -14 481 14 509
rect 52 481 80 509
rect 118 481 146 509
rect 184 481 212 509
rect 250 481 278 509
rect 316 481 344 509
rect 382 481 410 509
rect 448 481 476 509
rect 514 481 542 509
rect 580 481 608 509
rect 646 481 674 509
rect 712 481 740 509
rect -740 415 -712 443
rect -674 415 -646 443
rect -608 415 -580 443
rect -542 415 -514 443
rect -476 415 -448 443
rect -410 415 -382 443
rect -344 415 -316 443
rect -278 415 -250 443
rect -212 415 -184 443
rect -146 415 -118 443
rect -80 415 -52 443
rect -14 415 14 443
rect 52 415 80 443
rect 118 415 146 443
rect 184 415 212 443
rect 250 415 278 443
rect 316 415 344 443
rect 382 415 410 443
rect 448 415 476 443
rect 514 415 542 443
rect 580 415 608 443
rect 646 415 674 443
rect 712 415 740 443
rect -740 349 -712 377
rect -674 349 -646 377
rect -608 349 -580 377
rect -542 349 -514 377
rect -476 349 -448 377
rect -410 349 -382 377
rect -344 349 -316 377
rect -278 349 -250 377
rect -212 349 -184 377
rect -146 349 -118 377
rect -80 349 -52 377
rect -14 349 14 377
rect 52 349 80 377
rect 118 349 146 377
rect 184 349 212 377
rect 250 349 278 377
rect 316 349 344 377
rect 382 349 410 377
rect 448 349 476 377
rect 514 349 542 377
rect 580 349 608 377
rect 646 349 674 377
rect 712 349 740 377
rect -740 283 -712 311
rect -674 283 -646 311
rect -608 283 -580 311
rect -542 283 -514 311
rect -476 283 -448 311
rect -410 283 -382 311
rect -344 283 -316 311
rect -278 283 -250 311
rect -212 283 -184 311
rect -146 283 -118 311
rect -80 283 -52 311
rect -14 283 14 311
rect 52 283 80 311
rect 118 283 146 311
rect 184 283 212 311
rect 250 283 278 311
rect 316 283 344 311
rect 382 283 410 311
rect 448 283 476 311
rect 514 283 542 311
rect 580 283 608 311
rect 646 283 674 311
rect 712 283 740 311
rect -740 217 -712 245
rect -674 217 -646 245
rect -608 217 -580 245
rect -542 217 -514 245
rect -476 217 -448 245
rect -410 217 -382 245
rect -344 217 -316 245
rect -278 217 -250 245
rect -212 217 -184 245
rect -146 217 -118 245
rect -80 217 -52 245
rect -14 217 14 245
rect 52 217 80 245
rect 118 217 146 245
rect 184 217 212 245
rect 250 217 278 245
rect 316 217 344 245
rect 382 217 410 245
rect 448 217 476 245
rect 514 217 542 245
rect 580 217 608 245
rect 646 217 674 245
rect 712 217 740 245
rect -740 151 -712 179
rect -674 151 -646 179
rect -608 151 -580 179
rect -542 151 -514 179
rect -476 151 -448 179
rect -410 151 -382 179
rect -344 151 -316 179
rect -278 151 -250 179
rect -212 151 -184 179
rect -146 151 -118 179
rect -80 151 -52 179
rect -14 151 14 179
rect 52 151 80 179
rect 118 151 146 179
rect 184 151 212 179
rect 250 151 278 179
rect 316 151 344 179
rect 382 151 410 179
rect 448 151 476 179
rect 514 151 542 179
rect 580 151 608 179
rect 646 151 674 179
rect 712 151 740 179
rect -740 85 -712 113
rect -674 85 -646 113
rect -608 85 -580 113
rect -542 85 -514 113
rect -476 85 -448 113
rect -410 85 -382 113
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect 382 85 410 113
rect 448 85 476 113
rect 514 85 542 113
rect 580 85 608 113
rect 646 85 674 113
rect 712 85 740 113
rect -740 19 -712 47
rect -674 19 -646 47
rect -608 19 -580 47
rect -542 19 -514 47
rect -476 19 -448 47
rect -410 19 -382 47
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect 382 19 410 47
rect 448 19 476 47
rect 514 19 542 47
rect 580 19 608 47
rect 646 19 674 47
rect 712 19 740 47
rect -740 -47 -712 -19
rect -674 -47 -646 -19
rect -608 -47 -580 -19
rect -542 -47 -514 -19
rect -476 -47 -448 -19
rect -410 -47 -382 -19
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect 382 -47 410 -19
rect 448 -47 476 -19
rect 514 -47 542 -19
rect 580 -47 608 -19
rect 646 -47 674 -19
rect 712 -47 740 -19
rect -740 -113 -712 -85
rect -674 -113 -646 -85
rect -608 -113 -580 -85
rect -542 -113 -514 -85
rect -476 -113 -448 -85
rect -410 -113 -382 -85
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect 382 -113 410 -85
rect 448 -113 476 -85
rect 514 -113 542 -85
rect 580 -113 608 -85
rect 646 -113 674 -85
rect 712 -113 740 -85
rect -740 -179 -712 -151
rect -674 -179 -646 -151
rect -608 -179 -580 -151
rect -542 -179 -514 -151
rect -476 -179 -448 -151
rect -410 -179 -382 -151
rect -344 -179 -316 -151
rect -278 -179 -250 -151
rect -212 -179 -184 -151
rect -146 -179 -118 -151
rect -80 -179 -52 -151
rect -14 -179 14 -151
rect 52 -179 80 -151
rect 118 -179 146 -151
rect 184 -179 212 -151
rect 250 -179 278 -151
rect 316 -179 344 -151
rect 382 -179 410 -151
rect 448 -179 476 -151
rect 514 -179 542 -151
rect 580 -179 608 -151
rect 646 -179 674 -151
rect 712 -179 740 -151
rect -740 -245 -712 -217
rect -674 -245 -646 -217
rect -608 -245 -580 -217
rect -542 -245 -514 -217
rect -476 -245 -448 -217
rect -410 -245 -382 -217
rect -344 -245 -316 -217
rect -278 -245 -250 -217
rect -212 -245 -184 -217
rect -146 -245 -118 -217
rect -80 -245 -52 -217
rect -14 -245 14 -217
rect 52 -245 80 -217
rect 118 -245 146 -217
rect 184 -245 212 -217
rect 250 -245 278 -217
rect 316 -245 344 -217
rect 382 -245 410 -217
rect 448 -245 476 -217
rect 514 -245 542 -217
rect 580 -245 608 -217
rect 646 -245 674 -217
rect 712 -245 740 -217
rect -740 -311 -712 -283
rect -674 -311 -646 -283
rect -608 -311 -580 -283
rect -542 -311 -514 -283
rect -476 -311 -448 -283
rect -410 -311 -382 -283
rect -344 -311 -316 -283
rect -278 -311 -250 -283
rect -212 -311 -184 -283
rect -146 -311 -118 -283
rect -80 -311 -52 -283
rect -14 -311 14 -283
rect 52 -311 80 -283
rect 118 -311 146 -283
rect 184 -311 212 -283
rect 250 -311 278 -283
rect 316 -311 344 -283
rect 382 -311 410 -283
rect 448 -311 476 -283
rect 514 -311 542 -283
rect 580 -311 608 -283
rect 646 -311 674 -283
rect 712 -311 740 -283
rect -740 -377 -712 -349
rect -674 -377 -646 -349
rect -608 -377 -580 -349
rect -542 -377 -514 -349
rect -476 -377 -448 -349
rect -410 -377 -382 -349
rect -344 -377 -316 -349
rect -278 -377 -250 -349
rect -212 -377 -184 -349
rect -146 -377 -118 -349
rect -80 -377 -52 -349
rect -14 -377 14 -349
rect 52 -377 80 -349
rect 118 -377 146 -349
rect 184 -377 212 -349
rect 250 -377 278 -349
rect 316 -377 344 -349
rect 382 -377 410 -349
rect 448 -377 476 -349
rect 514 -377 542 -349
rect 580 -377 608 -349
rect 646 -377 674 -349
rect 712 -377 740 -349
rect -740 -443 -712 -415
rect -674 -443 -646 -415
rect -608 -443 -580 -415
rect -542 -443 -514 -415
rect -476 -443 -448 -415
rect -410 -443 -382 -415
rect -344 -443 -316 -415
rect -278 -443 -250 -415
rect -212 -443 -184 -415
rect -146 -443 -118 -415
rect -80 -443 -52 -415
rect -14 -443 14 -415
rect 52 -443 80 -415
rect 118 -443 146 -415
rect 184 -443 212 -415
rect 250 -443 278 -415
rect 316 -443 344 -415
rect 382 -443 410 -415
rect 448 -443 476 -415
rect 514 -443 542 -415
rect 580 -443 608 -415
rect 646 -443 674 -415
rect 712 -443 740 -415
rect -740 -509 -712 -481
rect -674 -509 -646 -481
rect -608 -509 -580 -481
rect -542 -509 -514 -481
rect -476 -509 -448 -481
rect -410 -509 -382 -481
rect -344 -509 -316 -481
rect -278 -509 -250 -481
rect -212 -509 -184 -481
rect -146 -509 -118 -481
rect -80 -509 -52 -481
rect -14 -509 14 -481
rect 52 -509 80 -481
rect 118 -509 146 -481
rect 184 -509 212 -481
rect 250 -509 278 -481
rect 316 -509 344 -481
rect 382 -509 410 -481
rect 448 -509 476 -481
rect 514 -509 542 -481
rect 580 -509 608 -481
rect 646 -509 674 -481
rect 712 -509 740 -481
rect -740 -575 -712 -547
rect -674 -575 -646 -547
rect -608 -575 -580 -547
rect -542 -575 -514 -547
rect -476 -575 -448 -547
rect -410 -575 -382 -547
rect -344 -575 -316 -547
rect -278 -575 -250 -547
rect -212 -575 -184 -547
rect -146 -575 -118 -547
rect -80 -575 -52 -547
rect -14 -575 14 -547
rect 52 -575 80 -547
rect 118 -575 146 -547
rect 184 -575 212 -547
rect 250 -575 278 -547
rect 316 -575 344 -547
rect 382 -575 410 -547
rect 448 -575 476 -547
rect 514 -575 542 -547
rect 580 -575 608 -547
rect 646 -575 674 -547
rect 712 -575 740 -547
rect -740 -641 -712 -613
rect -674 -641 -646 -613
rect -608 -641 -580 -613
rect -542 -641 -514 -613
rect -476 -641 -448 -613
rect -410 -641 -382 -613
rect -344 -641 -316 -613
rect -278 -641 -250 -613
rect -212 -641 -184 -613
rect -146 -641 -118 -613
rect -80 -641 -52 -613
rect -14 -641 14 -613
rect 52 -641 80 -613
rect 118 -641 146 -613
rect 184 -641 212 -613
rect 250 -641 278 -613
rect 316 -641 344 -613
rect 382 -641 410 -613
rect 448 -641 476 -613
rect 514 -641 542 -613
rect 580 -641 608 -613
rect 646 -641 674 -613
rect 712 -641 740 -613
rect -740 -707 -712 -679
rect -674 -707 -646 -679
rect -608 -707 -580 -679
rect -542 -707 -514 -679
rect -476 -707 -448 -679
rect -410 -707 -382 -679
rect -344 -707 -316 -679
rect -278 -707 -250 -679
rect -212 -707 -184 -679
rect -146 -707 -118 -679
rect -80 -707 -52 -679
rect -14 -707 14 -679
rect 52 -707 80 -679
rect 118 -707 146 -679
rect 184 -707 212 -679
rect 250 -707 278 -679
rect 316 -707 344 -679
rect 382 -707 410 -679
rect 448 -707 476 -679
rect 514 -707 542 -679
rect 580 -707 608 -679
rect 646 -707 674 -679
rect 712 -707 740 -679
rect -740 -773 -712 -745
rect -674 -773 -646 -745
rect -608 -773 -580 -745
rect -542 -773 -514 -745
rect -476 -773 -448 -745
rect -410 -773 -382 -745
rect -344 -773 -316 -745
rect -278 -773 -250 -745
rect -212 -773 -184 -745
rect -146 -773 -118 -745
rect -80 -773 -52 -745
rect -14 -773 14 -745
rect 52 -773 80 -745
rect 118 -773 146 -745
rect 184 -773 212 -745
rect 250 -773 278 -745
rect 316 -773 344 -745
rect 382 -773 410 -745
rect 448 -773 476 -745
rect 514 -773 542 -745
rect 580 -773 608 -745
rect 646 -773 674 -745
rect 712 -773 740 -745
rect -740 -839 -712 -811
rect -674 -839 -646 -811
rect -608 -839 -580 -811
rect -542 -839 -514 -811
rect -476 -839 -448 -811
rect -410 -839 -382 -811
rect -344 -839 -316 -811
rect -278 -839 -250 -811
rect -212 -839 -184 -811
rect -146 -839 -118 -811
rect -80 -839 -52 -811
rect -14 -839 14 -811
rect 52 -839 80 -811
rect 118 -839 146 -811
rect 184 -839 212 -811
rect 250 -839 278 -811
rect 316 -839 344 -811
rect 382 -839 410 -811
rect 448 -839 476 -811
rect 514 -839 542 -811
rect 580 -839 608 -811
rect 646 -839 674 -811
rect 712 -839 740 -811
rect -740 -905 -712 -877
rect -674 -905 -646 -877
rect -608 -905 -580 -877
rect -542 -905 -514 -877
rect -476 -905 -448 -877
rect -410 -905 -382 -877
rect -344 -905 -316 -877
rect -278 -905 -250 -877
rect -212 -905 -184 -877
rect -146 -905 -118 -877
rect -80 -905 -52 -877
rect -14 -905 14 -877
rect 52 -905 80 -877
rect 118 -905 146 -877
rect 184 -905 212 -877
rect 250 -905 278 -877
rect 316 -905 344 -877
rect 382 -905 410 -877
rect 448 -905 476 -877
rect 514 -905 542 -877
rect 580 -905 608 -877
rect 646 -905 674 -877
rect 712 -905 740 -877
rect -740 -971 -712 -943
rect -674 -971 -646 -943
rect -608 -971 -580 -943
rect -542 -971 -514 -943
rect -476 -971 -448 -943
rect -410 -971 -382 -943
rect -344 -971 -316 -943
rect -278 -971 -250 -943
rect -212 -971 -184 -943
rect -146 -971 -118 -943
rect -80 -971 -52 -943
rect -14 -971 14 -943
rect 52 -971 80 -943
rect 118 -971 146 -943
rect 184 -971 212 -943
rect 250 -971 278 -943
rect 316 -971 344 -943
rect 382 -971 410 -943
rect 448 -971 476 -943
rect 514 -971 542 -943
rect 580 -971 608 -943
rect 646 -971 674 -943
rect 712 -971 740 -943
rect -740 -1037 -712 -1009
rect -674 -1037 -646 -1009
rect -608 -1037 -580 -1009
rect -542 -1037 -514 -1009
rect -476 -1037 -448 -1009
rect -410 -1037 -382 -1009
rect -344 -1037 -316 -1009
rect -278 -1037 -250 -1009
rect -212 -1037 -184 -1009
rect -146 -1037 -118 -1009
rect -80 -1037 -52 -1009
rect -14 -1037 14 -1009
rect 52 -1037 80 -1009
rect 118 -1037 146 -1009
rect 184 -1037 212 -1009
rect 250 -1037 278 -1009
rect 316 -1037 344 -1009
rect 382 -1037 410 -1009
rect 448 -1037 476 -1009
rect 514 -1037 542 -1009
rect 580 -1037 608 -1009
rect 646 -1037 674 -1009
rect 712 -1037 740 -1009
rect -740 -1103 -712 -1075
rect -674 -1103 -646 -1075
rect -608 -1103 -580 -1075
rect -542 -1103 -514 -1075
rect -476 -1103 -448 -1075
rect -410 -1103 -382 -1075
rect -344 -1103 -316 -1075
rect -278 -1103 -250 -1075
rect -212 -1103 -184 -1075
rect -146 -1103 -118 -1075
rect -80 -1103 -52 -1075
rect -14 -1103 14 -1075
rect 52 -1103 80 -1075
rect 118 -1103 146 -1075
rect 184 -1103 212 -1075
rect 250 -1103 278 -1075
rect 316 -1103 344 -1075
rect 382 -1103 410 -1075
rect 448 -1103 476 -1075
rect 514 -1103 542 -1075
rect 580 -1103 608 -1075
rect 646 -1103 674 -1075
rect 712 -1103 740 -1075
rect -740 -1169 -712 -1141
rect -674 -1169 -646 -1141
rect -608 -1169 -580 -1141
rect -542 -1169 -514 -1141
rect -476 -1169 -448 -1141
rect -410 -1169 -382 -1141
rect -344 -1169 -316 -1141
rect -278 -1169 -250 -1141
rect -212 -1169 -184 -1141
rect -146 -1169 -118 -1141
rect -80 -1169 -52 -1141
rect -14 -1169 14 -1141
rect 52 -1169 80 -1141
rect 118 -1169 146 -1141
rect 184 -1169 212 -1141
rect 250 -1169 278 -1141
rect 316 -1169 344 -1141
rect 382 -1169 410 -1141
rect 448 -1169 476 -1141
rect 514 -1169 542 -1141
rect 580 -1169 608 -1141
rect 646 -1169 674 -1141
rect 712 -1169 740 -1141
rect -740 -1235 -712 -1207
rect -674 -1235 -646 -1207
rect -608 -1235 -580 -1207
rect -542 -1235 -514 -1207
rect -476 -1235 -448 -1207
rect -410 -1235 -382 -1207
rect -344 -1235 -316 -1207
rect -278 -1235 -250 -1207
rect -212 -1235 -184 -1207
rect -146 -1235 -118 -1207
rect -80 -1235 -52 -1207
rect -14 -1235 14 -1207
rect 52 -1235 80 -1207
rect 118 -1235 146 -1207
rect 184 -1235 212 -1207
rect 250 -1235 278 -1207
rect 316 -1235 344 -1207
rect 382 -1235 410 -1207
rect 448 -1235 476 -1207
rect 514 -1235 542 -1207
rect 580 -1235 608 -1207
rect 646 -1235 674 -1207
rect 712 -1235 740 -1207
rect -740 -1301 -712 -1273
rect -674 -1301 -646 -1273
rect -608 -1301 -580 -1273
rect -542 -1301 -514 -1273
rect -476 -1301 -448 -1273
rect -410 -1301 -382 -1273
rect -344 -1301 -316 -1273
rect -278 -1301 -250 -1273
rect -212 -1301 -184 -1273
rect -146 -1301 -118 -1273
rect -80 -1301 -52 -1273
rect -14 -1301 14 -1273
rect 52 -1301 80 -1273
rect 118 -1301 146 -1273
rect 184 -1301 212 -1273
rect 250 -1301 278 -1273
rect 316 -1301 344 -1273
rect 382 -1301 410 -1273
rect 448 -1301 476 -1273
rect 514 -1301 542 -1273
rect 580 -1301 608 -1273
rect 646 -1301 674 -1273
rect 712 -1301 740 -1273
rect -740 -1367 -712 -1339
rect -674 -1367 -646 -1339
rect -608 -1367 -580 -1339
rect -542 -1367 -514 -1339
rect -476 -1367 -448 -1339
rect -410 -1367 -382 -1339
rect -344 -1367 -316 -1339
rect -278 -1367 -250 -1339
rect -212 -1367 -184 -1339
rect -146 -1367 -118 -1339
rect -80 -1367 -52 -1339
rect -14 -1367 14 -1339
rect 52 -1367 80 -1339
rect 118 -1367 146 -1339
rect 184 -1367 212 -1339
rect 250 -1367 278 -1339
rect 316 -1367 344 -1339
rect 382 -1367 410 -1339
rect 448 -1367 476 -1339
rect 514 -1367 542 -1339
rect 580 -1367 608 -1339
rect 646 -1367 674 -1339
rect 712 -1367 740 -1339
rect -740 -1433 -712 -1405
rect -674 -1433 -646 -1405
rect -608 -1433 -580 -1405
rect -542 -1433 -514 -1405
rect -476 -1433 -448 -1405
rect -410 -1433 -382 -1405
rect -344 -1433 -316 -1405
rect -278 -1433 -250 -1405
rect -212 -1433 -184 -1405
rect -146 -1433 -118 -1405
rect -80 -1433 -52 -1405
rect -14 -1433 14 -1405
rect 52 -1433 80 -1405
rect 118 -1433 146 -1405
rect 184 -1433 212 -1405
rect 250 -1433 278 -1405
rect 316 -1433 344 -1405
rect 382 -1433 410 -1405
rect 448 -1433 476 -1405
rect 514 -1433 542 -1405
rect 580 -1433 608 -1405
rect 646 -1433 674 -1405
rect 712 -1433 740 -1405
rect -740 -1499 -712 -1471
rect -674 -1499 -646 -1471
rect -608 -1499 -580 -1471
rect -542 -1499 -514 -1471
rect -476 -1499 -448 -1471
rect -410 -1499 -382 -1471
rect -344 -1499 -316 -1471
rect -278 -1499 -250 -1471
rect -212 -1499 -184 -1471
rect -146 -1499 -118 -1471
rect -80 -1499 -52 -1471
rect -14 -1499 14 -1471
rect 52 -1499 80 -1471
rect 118 -1499 146 -1471
rect 184 -1499 212 -1471
rect 250 -1499 278 -1471
rect 316 -1499 344 -1471
rect 382 -1499 410 -1471
rect 448 -1499 476 -1471
rect 514 -1499 542 -1471
rect 580 -1499 608 -1471
rect 646 -1499 674 -1471
rect 712 -1499 740 -1471
rect -740 -1565 -712 -1537
rect -674 -1565 -646 -1537
rect -608 -1565 -580 -1537
rect -542 -1565 -514 -1537
rect -476 -1565 -448 -1537
rect -410 -1565 -382 -1537
rect -344 -1565 -316 -1537
rect -278 -1565 -250 -1537
rect -212 -1565 -184 -1537
rect -146 -1565 -118 -1537
rect -80 -1565 -52 -1537
rect -14 -1565 14 -1537
rect 52 -1565 80 -1537
rect 118 -1565 146 -1537
rect 184 -1565 212 -1537
rect 250 -1565 278 -1537
rect 316 -1565 344 -1537
rect 382 -1565 410 -1537
rect 448 -1565 476 -1537
rect 514 -1565 542 -1537
rect 580 -1565 608 -1537
rect 646 -1565 674 -1537
rect 712 -1565 740 -1537
rect -740 -1631 -712 -1603
rect -674 -1631 -646 -1603
rect -608 -1631 -580 -1603
rect -542 -1631 -514 -1603
rect -476 -1631 -448 -1603
rect -410 -1631 -382 -1603
rect -344 -1631 -316 -1603
rect -278 -1631 -250 -1603
rect -212 -1631 -184 -1603
rect -146 -1631 -118 -1603
rect -80 -1631 -52 -1603
rect -14 -1631 14 -1603
rect 52 -1631 80 -1603
rect 118 -1631 146 -1603
rect 184 -1631 212 -1603
rect 250 -1631 278 -1603
rect 316 -1631 344 -1603
rect 382 -1631 410 -1603
rect 448 -1631 476 -1603
rect 514 -1631 542 -1603
rect 580 -1631 608 -1603
rect 646 -1631 674 -1603
rect 712 -1631 740 -1603
rect -740 -1697 -712 -1669
rect -674 -1697 -646 -1669
rect -608 -1697 -580 -1669
rect -542 -1697 -514 -1669
rect -476 -1697 -448 -1669
rect -410 -1697 -382 -1669
rect -344 -1697 -316 -1669
rect -278 -1697 -250 -1669
rect -212 -1697 -184 -1669
rect -146 -1697 -118 -1669
rect -80 -1697 -52 -1669
rect -14 -1697 14 -1669
rect 52 -1697 80 -1669
rect 118 -1697 146 -1669
rect 184 -1697 212 -1669
rect 250 -1697 278 -1669
rect 316 -1697 344 -1669
rect 382 -1697 410 -1669
rect 448 -1697 476 -1669
rect 514 -1697 542 -1669
rect 580 -1697 608 -1669
rect 646 -1697 674 -1669
rect 712 -1697 740 -1669
rect -740 -1763 -712 -1735
rect -674 -1763 -646 -1735
rect -608 -1763 -580 -1735
rect -542 -1763 -514 -1735
rect -476 -1763 -448 -1735
rect -410 -1763 -382 -1735
rect -344 -1763 -316 -1735
rect -278 -1763 -250 -1735
rect -212 -1763 -184 -1735
rect -146 -1763 -118 -1735
rect -80 -1763 -52 -1735
rect -14 -1763 14 -1735
rect 52 -1763 80 -1735
rect 118 -1763 146 -1735
rect 184 -1763 212 -1735
rect 250 -1763 278 -1735
rect 316 -1763 344 -1735
rect 382 -1763 410 -1735
rect 448 -1763 476 -1735
rect 514 -1763 542 -1735
rect 580 -1763 608 -1735
rect 646 -1763 674 -1735
rect 712 -1763 740 -1735
rect -740 -1829 -712 -1801
rect -674 -1829 -646 -1801
rect -608 -1829 -580 -1801
rect -542 -1829 -514 -1801
rect -476 -1829 -448 -1801
rect -410 -1829 -382 -1801
rect -344 -1829 -316 -1801
rect -278 -1829 -250 -1801
rect -212 -1829 -184 -1801
rect -146 -1829 -118 -1801
rect -80 -1829 -52 -1801
rect -14 -1829 14 -1801
rect 52 -1829 80 -1801
rect 118 -1829 146 -1801
rect 184 -1829 212 -1801
rect 250 -1829 278 -1801
rect 316 -1829 344 -1801
rect 382 -1829 410 -1801
rect 448 -1829 476 -1801
rect 514 -1829 542 -1801
rect 580 -1829 608 -1801
rect 646 -1829 674 -1801
rect 712 -1829 740 -1801
rect -740 -1895 -712 -1867
rect -674 -1895 -646 -1867
rect -608 -1895 -580 -1867
rect -542 -1895 -514 -1867
rect -476 -1895 -448 -1867
rect -410 -1895 -382 -1867
rect -344 -1895 -316 -1867
rect -278 -1895 -250 -1867
rect -212 -1895 -184 -1867
rect -146 -1895 -118 -1867
rect -80 -1895 -52 -1867
rect -14 -1895 14 -1867
rect 52 -1895 80 -1867
rect 118 -1895 146 -1867
rect 184 -1895 212 -1867
rect 250 -1895 278 -1867
rect 316 -1895 344 -1867
rect 382 -1895 410 -1867
rect 448 -1895 476 -1867
rect 514 -1895 542 -1867
rect 580 -1895 608 -1867
rect 646 -1895 674 -1867
rect 712 -1895 740 -1867
rect -740 -1961 -712 -1933
rect -674 -1961 -646 -1933
rect -608 -1961 -580 -1933
rect -542 -1961 -514 -1933
rect -476 -1961 -448 -1933
rect -410 -1961 -382 -1933
rect -344 -1961 -316 -1933
rect -278 -1961 -250 -1933
rect -212 -1961 -184 -1933
rect -146 -1961 -118 -1933
rect -80 -1961 -52 -1933
rect -14 -1961 14 -1933
rect 52 -1961 80 -1933
rect 118 -1961 146 -1933
rect 184 -1961 212 -1933
rect 250 -1961 278 -1933
rect 316 -1961 344 -1933
rect 382 -1961 410 -1933
rect 448 -1961 476 -1933
rect 514 -1961 542 -1933
rect 580 -1961 608 -1933
rect 646 -1961 674 -1933
rect 712 -1961 740 -1933
rect -740 -2027 -712 -1999
rect -674 -2027 -646 -1999
rect -608 -2027 -580 -1999
rect -542 -2027 -514 -1999
rect -476 -2027 -448 -1999
rect -410 -2027 -382 -1999
rect -344 -2027 -316 -1999
rect -278 -2027 -250 -1999
rect -212 -2027 -184 -1999
rect -146 -2027 -118 -1999
rect -80 -2027 -52 -1999
rect -14 -2027 14 -1999
rect 52 -2027 80 -1999
rect 118 -2027 146 -1999
rect 184 -2027 212 -1999
rect 250 -2027 278 -1999
rect 316 -2027 344 -1999
rect 382 -2027 410 -1999
rect 448 -2027 476 -1999
rect 514 -2027 542 -1999
rect 580 -2027 608 -1999
rect 646 -2027 674 -1999
rect 712 -2027 740 -1999
rect -740 -2093 -712 -2065
rect -674 -2093 -646 -2065
rect -608 -2093 -580 -2065
rect -542 -2093 -514 -2065
rect -476 -2093 -448 -2065
rect -410 -2093 -382 -2065
rect -344 -2093 -316 -2065
rect -278 -2093 -250 -2065
rect -212 -2093 -184 -2065
rect -146 -2093 -118 -2065
rect -80 -2093 -52 -2065
rect -14 -2093 14 -2065
rect 52 -2093 80 -2065
rect 118 -2093 146 -2065
rect 184 -2093 212 -2065
rect 250 -2093 278 -2065
rect 316 -2093 344 -2065
rect 382 -2093 410 -2065
rect 448 -2093 476 -2065
rect 514 -2093 542 -2065
rect 580 -2093 608 -2065
rect 646 -2093 674 -2065
rect 712 -2093 740 -2065
rect -740 -2159 -712 -2131
rect -674 -2159 -646 -2131
rect -608 -2159 -580 -2131
rect -542 -2159 -514 -2131
rect -476 -2159 -448 -2131
rect -410 -2159 -382 -2131
rect -344 -2159 -316 -2131
rect -278 -2159 -250 -2131
rect -212 -2159 -184 -2131
rect -146 -2159 -118 -2131
rect -80 -2159 -52 -2131
rect -14 -2159 14 -2131
rect 52 -2159 80 -2131
rect 118 -2159 146 -2131
rect 184 -2159 212 -2131
rect 250 -2159 278 -2131
rect 316 -2159 344 -2131
rect 382 -2159 410 -2131
rect 448 -2159 476 -2131
rect 514 -2159 542 -2131
rect 580 -2159 608 -2131
rect 646 -2159 674 -2131
rect 712 -2159 740 -2131
rect -740 -2225 -712 -2197
rect -674 -2225 -646 -2197
rect -608 -2225 -580 -2197
rect -542 -2225 -514 -2197
rect -476 -2225 -448 -2197
rect -410 -2225 -382 -2197
rect -344 -2225 -316 -2197
rect -278 -2225 -250 -2197
rect -212 -2225 -184 -2197
rect -146 -2225 -118 -2197
rect -80 -2225 -52 -2197
rect -14 -2225 14 -2197
rect 52 -2225 80 -2197
rect 118 -2225 146 -2197
rect 184 -2225 212 -2197
rect 250 -2225 278 -2197
rect 316 -2225 344 -2197
rect 382 -2225 410 -2197
rect 448 -2225 476 -2197
rect 514 -2225 542 -2197
rect 580 -2225 608 -2197
rect 646 -2225 674 -2197
rect 712 -2225 740 -2197
rect -740 -2291 -712 -2263
rect -674 -2291 -646 -2263
rect -608 -2291 -580 -2263
rect -542 -2291 -514 -2263
rect -476 -2291 -448 -2263
rect -410 -2291 -382 -2263
rect -344 -2291 -316 -2263
rect -278 -2291 -250 -2263
rect -212 -2291 -184 -2263
rect -146 -2291 -118 -2263
rect -80 -2291 -52 -2263
rect -14 -2291 14 -2263
rect 52 -2291 80 -2263
rect 118 -2291 146 -2263
rect 184 -2291 212 -2263
rect 250 -2291 278 -2263
rect 316 -2291 344 -2263
rect 382 -2291 410 -2263
rect 448 -2291 476 -2263
rect 514 -2291 542 -2263
rect 580 -2291 608 -2263
rect 646 -2291 674 -2263
rect 712 -2291 740 -2263
rect -740 -2357 -712 -2329
rect -674 -2357 -646 -2329
rect -608 -2357 -580 -2329
rect -542 -2357 -514 -2329
rect -476 -2357 -448 -2329
rect -410 -2357 -382 -2329
rect -344 -2357 -316 -2329
rect -278 -2357 -250 -2329
rect -212 -2357 -184 -2329
rect -146 -2357 -118 -2329
rect -80 -2357 -52 -2329
rect -14 -2357 14 -2329
rect 52 -2357 80 -2329
rect 118 -2357 146 -2329
rect 184 -2357 212 -2329
rect 250 -2357 278 -2329
rect 316 -2357 344 -2329
rect 382 -2357 410 -2329
rect 448 -2357 476 -2329
rect 514 -2357 542 -2329
rect 580 -2357 608 -2329
rect 646 -2357 674 -2329
rect 712 -2357 740 -2329
rect -740 -2423 -712 -2395
rect -674 -2423 -646 -2395
rect -608 -2423 -580 -2395
rect -542 -2423 -514 -2395
rect -476 -2423 -448 -2395
rect -410 -2423 -382 -2395
rect -344 -2423 -316 -2395
rect -278 -2423 -250 -2395
rect -212 -2423 -184 -2395
rect -146 -2423 -118 -2395
rect -80 -2423 -52 -2395
rect -14 -2423 14 -2395
rect 52 -2423 80 -2395
rect 118 -2423 146 -2395
rect 184 -2423 212 -2395
rect 250 -2423 278 -2395
rect 316 -2423 344 -2395
rect 382 -2423 410 -2395
rect 448 -2423 476 -2395
rect 514 -2423 542 -2395
rect 580 -2423 608 -2395
rect 646 -2423 674 -2395
rect 712 -2423 740 -2395
rect -740 -2489 -712 -2461
rect -674 -2489 -646 -2461
rect -608 -2489 -580 -2461
rect -542 -2489 -514 -2461
rect -476 -2489 -448 -2461
rect -410 -2489 -382 -2461
rect -344 -2489 -316 -2461
rect -278 -2489 -250 -2461
rect -212 -2489 -184 -2461
rect -146 -2489 -118 -2461
rect -80 -2489 -52 -2461
rect -14 -2489 14 -2461
rect 52 -2489 80 -2461
rect 118 -2489 146 -2461
rect 184 -2489 212 -2461
rect 250 -2489 278 -2461
rect 316 -2489 344 -2461
rect 382 -2489 410 -2461
rect 448 -2489 476 -2461
rect 514 -2489 542 -2461
rect 580 -2489 608 -2461
rect 646 -2489 674 -2461
rect 712 -2489 740 -2461
rect -740 -2555 -712 -2527
rect -674 -2555 -646 -2527
rect -608 -2555 -580 -2527
rect -542 -2555 -514 -2527
rect -476 -2555 -448 -2527
rect -410 -2555 -382 -2527
rect -344 -2555 -316 -2527
rect -278 -2555 -250 -2527
rect -212 -2555 -184 -2527
rect -146 -2555 -118 -2527
rect -80 -2555 -52 -2527
rect -14 -2555 14 -2527
rect 52 -2555 80 -2527
rect 118 -2555 146 -2527
rect 184 -2555 212 -2527
rect 250 -2555 278 -2527
rect 316 -2555 344 -2527
rect 382 -2555 410 -2527
rect 448 -2555 476 -2527
rect 514 -2555 542 -2527
rect 580 -2555 608 -2527
rect 646 -2555 674 -2527
rect 712 -2555 740 -2527
<< metal4 >>
rect -745 2555 745 2560
rect -745 2527 -740 2555
rect -712 2527 -674 2555
rect -646 2527 -608 2555
rect -580 2527 -542 2555
rect -514 2527 -476 2555
rect -448 2527 -410 2555
rect -382 2527 -344 2555
rect -316 2527 -278 2555
rect -250 2527 -212 2555
rect -184 2527 -146 2555
rect -118 2527 -80 2555
rect -52 2527 -14 2555
rect 14 2527 52 2555
rect 80 2527 118 2555
rect 146 2527 184 2555
rect 212 2527 250 2555
rect 278 2527 316 2555
rect 344 2527 382 2555
rect 410 2527 448 2555
rect 476 2527 514 2555
rect 542 2527 580 2555
rect 608 2527 646 2555
rect 674 2527 712 2555
rect 740 2527 745 2555
rect -745 2489 745 2527
rect -745 2461 -740 2489
rect -712 2461 -674 2489
rect -646 2461 -608 2489
rect -580 2461 -542 2489
rect -514 2461 -476 2489
rect -448 2461 -410 2489
rect -382 2461 -344 2489
rect -316 2461 -278 2489
rect -250 2461 -212 2489
rect -184 2461 -146 2489
rect -118 2461 -80 2489
rect -52 2461 -14 2489
rect 14 2461 52 2489
rect 80 2461 118 2489
rect 146 2461 184 2489
rect 212 2461 250 2489
rect 278 2461 316 2489
rect 344 2461 382 2489
rect 410 2461 448 2489
rect 476 2461 514 2489
rect 542 2461 580 2489
rect 608 2461 646 2489
rect 674 2461 712 2489
rect 740 2461 745 2489
rect -745 2423 745 2461
rect -745 2395 -740 2423
rect -712 2395 -674 2423
rect -646 2395 -608 2423
rect -580 2395 -542 2423
rect -514 2395 -476 2423
rect -448 2395 -410 2423
rect -382 2395 -344 2423
rect -316 2395 -278 2423
rect -250 2395 -212 2423
rect -184 2395 -146 2423
rect -118 2395 -80 2423
rect -52 2395 -14 2423
rect 14 2395 52 2423
rect 80 2395 118 2423
rect 146 2395 184 2423
rect 212 2395 250 2423
rect 278 2395 316 2423
rect 344 2395 382 2423
rect 410 2395 448 2423
rect 476 2395 514 2423
rect 542 2395 580 2423
rect 608 2395 646 2423
rect 674 2395 712 2423
rect 740 2395 745 2423
rect -745 2357 745 2395
rect -745 2329 -740 2357
rect -712 2329 -674 2357
rect -646 2329 -608 2357
rect -580 2329 -542 2357
rect -514 2329 -476 2357
rect -448 2329 -410 2357
rect -382 2329 -344 2357
rect -316 2329 -278 2357
rect -250 2329 -212 2357
rect -184 2329 -146 2357
rect -118 2329 -80 2357
rect -52 2329 -14 2357
rect 14 2329 52 2357
rect 80 2329 118 2357
rect 146 2329 184 2357
rect 212 2329 250 2357
rect 278 2329 316 2357
rect 344 2329 382 2357
rect 410 2329 448 2357
rect 476 2329 514 2357
rect 542 2329 580 2357
rect 608 2329 646 2357
rect 674 2329 712 2357
rect 740 2329 745 2357
rect -745 2291 745 2329
rect -745 2263 -740 2291
rect -712 2263 -674 2291
rect -646 2263 -608 2291
rect -580 2263 -542 2291
rect -514 2263 -476 2291
rect -448 2263 -410 2291
rect -382 2263 -344 2291
rect -316 2263 -278 2291
rect -250 2263 -212 2291
rect -184 2263 -146 2291
rect -118 2263 -80 2291
rect -52 2263 -14 2291
rect 14 2263 52 2291
rect 80 2263 118 2291
rect 146 2263 184 2291
rect 212 2263 250 2291
rect 278 2263 316 2291
rect 344 2263 382 2291
rect 410 2263 448 2291
rect 476 2263 514 2291
rect 542 2263 580 2291
rect 608 2263 646 2291
rect 674 2263 712 2291
rect 740 2263 745 2291
rect -745 2225 745 2263
rect -745 2197 -740 2225
rect -712 2197 -674 2225
rect -646 2197 -608 2225
rect -580 2197 -542 2225
rect -514 2197 -476 2225
rect -448 2197 -410 2225
rect -382 2197 -344 2225
rect -316 2197 -278 2225
rect -250 2197 -212 2225
rect -184 2197 -146 2225
rect -118 2197 -80 2225
rect -52 2197 -14 2225
rect 14 2197 52 2225
rect 80 2197 118 2225
rect 146 2197 184 2225
rect 212 2197 250 2225
rect 278 2197 316 2225
rect 344 2197 382 2225
rect 410 2197 448 2225
rect 476 2197 514 2225
rect 542 2197 580 2225
rect 608 2197 646 2225
rect 674 2197 712 2225
rect 740 2197 745 2225
rect -745 2159 745 2197
rect -745 2131 -740 2159
rect -712 2131 -674 2159
rect -646 2131 -608 2159
rect -580 2131 -542 2159
rect -514 2131 -476 2159
rect -448 2131 -410 2159
rect -382 2131 -344 2159
rect -316 2131 -278 2159
rect -250 2131 -212 2159
rect -184 2131 -146 2159
rect -118 2131 -80 2159
rect -52 2131 -14 2159
rect 14 2131 52 2159
rect 80 2131 118 2159
rect 146 2131 184 2159
rect 212 2131 250 2159
rect 278 2131 316 2159
rect 344 2131 382 2159
rect 410 2131 448 2159
rect 476 2131 514 2159
rect 542 2131 580 2159
rect 608 2131 646 2159
rect 674 2131 712 2159
rect 740 2131 745 2159
rect -745 2093 745 2131
rect -745 2065 -740 2093
rect -712 2065 -674 2093
rect -646 2065 -608 2093
rect -580 2065 -542 2093
rect -514 2065 -476 2093
rect -448 2065 -410 2093
rect -382 2065 -344 2093
rect -316 2065 -278 2093
rect -250 2065 -212 2093
rect -184 2065 -146 2093
rect -118 2065 -80 2093
rect -52 2065 -14 2093
rect 14 2065 52 2093
rect 80 2065 118 2093
rect 146 2065 184 2093
rect 212 2065 250 2093
rect 278 2065 316 2093
rect 344 2065 382 2093
rect 410 2065 448 2093
rect 476 2065 514 2093
rect 542 2065 580 2093
rect 608 2065 646 2093
rect 674 2065 712 2093
rect 740 2065 745 2093
rect -745 2027 745 2065
rect -745 1999 -740 2027
rect -712 1999 -674 2027
rect -646 1999 -608 2027
rect -580 1999 -542 2027
rect -514 1999 -476 2027
rect -448 1999 -410 2027
rect -382 1999 -344 2027
rect -316 1999 -278 2027
rect -250 1999 -212 2027
rect -184 1999 -146 2027
rect -118 1999 -80 2027
rect -52 1999 -14 2027
rect 14 1999 52 2027
rect 80 1999 118 2027
rect 146 1999 184 2027
rect 212 1999 250 2027
rect 278 1999 316 2027
rect 344 1999 382 2027
rect 410 1999 448 2027
rect 476 1999 514 2027
rect 542 1999 580 2027
rect 608 1999 646 2027
rect 674 1999 712 2027
rect 740 1999 745 2027
rect -745 1961 745 1999
rect -745 1933 -740 1961
rect -712 1933 -674 1961
rect -646 1933 -608 1961
rect -580 1933 -542 1961
rect -514 1933 -476 1961
rect -448 1933 -410 1961
rect -382 1933 -344 1961
rect -316 1933 -278 1961
rect -250 1933 -212 1961
rect -184 1933 -146 1961
rect -118 1933 -80 1961
rect -52 1933 -14 1961
rect 14 1933 52 1961
rect 80 1933 118 1961
rect 146 1933 184 1961
rect 212 1933 250 1961
rect 278 1933 316 1961
rect 344 1933 382 1961
rect 410 1933 448 1961
rect 476 1933 514 1961
rect 542 1933 580 1961
rect 608 1933 646 1961
rect 674 1933 712 1961
rect 740 1933 745 1961
rect -745 1895 745 1933
rect -745 1867 -740 1895
rect -712 1867 -674 1895
rect -646 1867 -608 1895
rect -580 1867 -542 1895
rect -514 1867 -476 1895
rect -448 1867 -410 1895
rect -382 1867 -344 1895
rect -316 1867 -278 1895
rect -250 1867 -212 1895
rect -184 1867 -146 1895
rect -118 1867 -80 1895
rect -52 1867 -14 1895
rect 14 1867 52 1895
rect 80 1867 118 1895
rect 146 1867 184 1895
rect 212 1867 250 1895
rect 278 1867 316 1895
rect 344 1867 382 1895
rect 410 1867 448 1895
rect 476 1867 514 1895
rect 542 1867 580 1895
rect 608 1867 646 1895
rect 674 1867 712 1895
rect 740 1867 745 1895
rect -745 1829 745 1867
rect -745 1801 -740 1829
rect -712 1801 -674 1829
rect -646 1801 -608 1829
rect -580 1801 -542 1829
rect -514 1801 -476 1829
rect -448 1801 -410 1829
rect -382 1801 -344 1829
rect -316 1801 -278 1829
rect -250 1801 -212 1829
rect -184 1801 -146 1829
rect -118 1801 -80 1829
rect -52 1801 -14 1829
rect 14 1801 52 1829
rect 80 1801 118 1829
rect 146 1801 184 1829
rect 212 1801 250 1829
rect 278 1801 316 1829
rect 344 1801 382 1829
rect 410 1801 448 1829
rect 476 1801 514 1829
rect 542 1801 580 1829
rect 608 1801 646 1829
rect 674 1801 712 1829
rect 740 1801 745 1829
rect -745 1763 745 1801
rect -745 1735 -740 1763
rect -712 1735 -674 1763
rect -646 1735 -608 1763
rect -580 1735 -542 1763
rect -514 1735 -476 1763
rect -448 1735 -410 1763
rect -382 1735 -344 1763
rect -316 1735 -278 1763
rect -250 1735 -212 1763
rect -184 1735 -146 1763
rect -118 1735 -80 1763
rect -52 1735 -14 1763
rect 14 1735 52 1763
rect 80 1735 118 1763
rect 146 1735 184 1763
rect 212 1735 250 1763
rect 278 1735 316 1763
rect 344 1735 382 1763
rect 410 1735 448 1763
rect 476 1735 514 1763
rect 542 1735 580 1763
rect 608 1735 646 1763
rect 674 1735 712 1763
rect 740 1735 745 1763
rect -745 1697 745 1735
rect -745 1669 -740 1697
rect -712 1669 -674 1697
rect -646 1669 -608 1697
rect -580 1669 -542 1697
rect -514 1669 -476 1697
rect -448 1669 -410 1697
rect -382 1669 -344 1697
rect -316 1669 -278 1697
rect -250 1669 -212 1697
rect -184 1669 -146 1697
rect -118 1669 -80 1697
rect -52 1669 -14 1697
rect 14 1669 52 1697
rect 80 1669 118 1697
rect 146 1669 184 1697
rect 212 1669 250 1697
rect 278 1669 316 1697
rect 344 1669 382 1697
rect 410 1669 448 1697
rect 476 1669 514 1697
rect 542 1669 580 1697
rect 608 1669 646 1697
rect 674 1669 712 1697
rect 740 1669 745 1697
rect -745 1631 745 1669
rect -745 1603 -740 1631
rect -712 1603 -674 1631
rect -646 1603 -608 1631
rect -580 1603 -542 1631
rect -514 1603 -476 1631
rect -448 1603 -410 1631
rect -382 1603 -344 1631
rect -316 1603 -278 1631
rect -250 1603 -212 1631
rect -184 1603 -146 1631
rect -118 1603 -80 1631
rect -52 1603 -14 1631
rect 14 1603 52 1631
rect 80 1603 118 1631
rect 146 1603 184 1631
rect 212 1603 250 1631
rect 278 1603 316 1631
rect 344 1603 382 1631
rect 410 1603 448 1631
rect 476 1603 514 1631
rect 542 1603 580 1631
rect 608 1603 646 1631
rect 674 1603 712 1631
rect 740 1603 745 1631
rect -745 1565 745 1603
rect -745 1537 -740 1565
rect -712 1537 -674 1565
rect -646 1537 -608 1565
rect -580 1537 -542 1565
rect -514 1537 -476 1565
rect -448 1537 -410 1565
rect -382 1537 -344 1565
rect -316 1537 -278 1565
rect -250 1537 -212 1565
rect -184 1537 -146 1565
rect -118 1537 -80 1565
rect -52 1537 -14 1565
rect 14 1537 52 1565
rect 80 1537 118 1565
rect 146 1537 184 1565
rect 212 1537 250 1565
rect 278 1537 316 1565
rect 344 1537 382 1565
rect 410 1537 448 1565
rect 476 1537 514 1565
rect 542 1537 580 1565
rect 608 1537 646 1565
rect 674 1537 712 1565
rect 740 1537 745 1565
rect -745 1499 745 1537
rect -745 1471 -740 1499
rect -712 1471 -674 1499
rect -646 1471 -608 1499
rect -580 1471 -542 1499
rect -514 1471 -476 1499
rect -448 1471 -410 1499
rect -382 1471 -344 1499
rect -316 1471 -278 1499
rect -250 1471 -212 1499
rect -184 1471 -146 1499
rect -118 1471 -80 1499
rect -52 1471 -14 1499
rect 14 1471 52 1499
rect 80 1471 118 1499
rect 146 1471 184 1499
rect 212 1471 250 1499
rect 278 1471 316 1499
rect 344 1471 382 1499
rect 410 1471 448 1499
rect 476 1471 514 1499
rect 542 1471 580 1499
rect 608 1471 646 1499
rect 674 1471 712 1499
rect 740 1471 745 1499
rect -745 1433 745 1471
rect -745 1405 -740 1433
rect -712 1405 -674 1433
rect -646 1405 -608 1433
rect -580 1405 -542 1433
rect -514 1405 -476 1433
rect -448 1405 -410 1433
rect -382 1405 -344 1433
rect -316 1405 -278 1433
rect -250 1405 -212 1433
rect -184 1405 -146 1433
rect -118 1405 -80 1433
rect -52 1405 -14 1433
rect 14 1405 52 1433
rect 80 1405 118 1433
rect 146 1405 184 1433
rect 212 1405 250 1433
rect 278 1405 316 1433
rect 344 1405 382 1433
rect 410 1405 448 1433
rect 476 1405 514 1433
rect 542 1405 580 1433
rect 608 1405 646 1433
rect 674 1405 712 1433
rect 740 1405 745 1433
rect -745 1367 745 1405
rect -745 1339 -740 1367
rect -712 1339 -674 1367
rect -646 1339 -608 1367
rect -580 1339 -542 1367
rect -514 1339 -476 1367
rect -448 1339 -410 1367
rect -382 1339 -344 1367
rect -316 1339 -278 1367
rect -250 1339 -212 1367
rect -184 1339 -146 1367
rect -118 1339 -80 1367
rect -52 1339 -14 1367
rect 14 1339 52 1367
rect 80 1339 118 1367
rect 146 1339 184 1367
rect 212 1339 250 1367
rect 278 1339 316 1367
rect 344 1339 382 1367
rect 410 1339 448 1367
rect 476 1339 514 1367
rect 542 1339 580 1367
rect 608 1339 646 1367
rect 674 1339 712 1367
rect 740 1339 745 1367
rect -745 1301 745 1339
rect -745 1273 -740 1301
rect -712 1273 -674 1301
rect -646 1273 -608 1301
rect -580 1273 -542 1301
rect -514 1273 -476 1301
rect -448 1273 -410 1301
rect -382 1273 -344 1301
rect -316 1273 -278 1301
rect -250 1273 -212 1301
rect -184 1273 -146 1301
rect -118 1273 -80 1301
rect -52 1273 -14 1301
rect 14 1273 52 1301
rect 80 1273 118 1301
rect 146 1273 184 1301
rect 212 1273 250 1301
rect 278 1273 316 1301
rect 344 1273 382 1301
rect 410 1273 448 1301
rect 476 1273 514 1301
rect 542 1273 580 1301
rect 608 1273 646 1301
rect 674 1273 712 1301
rect 740 1273 745 1301
rect -745 1235 745 1273
rect -745 1207 -740 1235
rect -712 1207 -674 1235
rect -646 1207 -608 1235
rect -580 1207 -542 1235
rect -514 1207 -476 1235
rect -448 1207 -410 1235
rect -382 1207 -344 1235
rect -316 1207 -278 1235
rect -250 1207 -212 1235
rect -184 1207 -146 1235
rect -118 1207 -80 1235
rect -52 1207 -14 1235
rect 14 1207 52 1235
rect 80 1207 118 1235
rect 146 1207 184 1235
rect 212 1207 250 1235
rect 278 1207 316 1235
rect 344 1207 382 1235
rect 410 1207 448 1235
rect 476 1207 514 1235
rect 542 1207 580 1235
rect 608 1207 646 1235
rect 674 1207 712 1235
rect 740 1207 745 1235
rect -745 1169 745 1207
rect -745 1141 -740 1169
rect -712 1141 -674 1169
rect -646 1141 -608 1169
rect -580 1141 -542 1169
rect -514 1141 -476 1169
rect -448 1141 -410 1169
rect -382 1141 -344 1169
rect -316 1141 -278 1169
rect -250 1141 -212 1169
rect -184 1141 -146 1169
rect -118 1141 -80 1169
rect -52 1141 -14 1169
rect 14 1141 52 1169
rect 80 1141 118 1169
rect 146 1141 184 1169
rect 212 1141 250 1169
rect 278 1141 316 1169
rect 344 1141 382 1169
rect 410 1141 448 1169
rect 476 1141 514 1169
rect 542 1141 580 1169
rect 608 1141 646 1169
rect 674 1141 712 1169
rect 740 1141 745 1169
rect -745 1103 745 1141
rect -745 1075 -740 1103
rect -712 1075 -674 1103
rect -646 1075 -608 1103
rect -580 1075 -542 1103
rect -514 1075 -476 1103
rect -448 1075 -410 1103
rect -382 1075 -344 1103
rect -316 1075 -278 1103
rect -250 1075 -212 1103
rect -184 1075 -146 1103
rect -118 1075 -80 1103
rect -52 1075 -14 1103
rect 14 1075 52 1103
rect 80 1075 118 1103
rect 146 1075 184 1103
rect 212 1075 250 1103
rect 278 1075 316 1103
rect 344 1075 382 1103
rect 410 1075 448 1103
rect 476 1075 514 1103
rect 542 1075 580 1103
rect 608 1075 646 1103
rect 674 1075 712 1103
rect 740 1075 745 1103
rect -745 1037 745 1075
rect -745 1009 -740 1037
rect -712 1009 -674 1037
rect -646 1009 -608 1037
rect -580 1009 -542 1037
rect -514 1009 -476 1037
rect -448 1009 -410 1037
rect -382 1009 -344 1037
rect -316 1009 -278 1037
rect -250 1009 -212 1037
rect -184 1009 -146 1037
rect -118 1009 -80 1037
rect -52 1009 -14 1037
rect 14 1009 52 1037
rect 80 1009 118 1037
rect 146 1009 184 1037
rect 212 1009 250 1037
rect 278 1009 316 1037
rect 344 1009 382 1037
rect 410 1009 448 1037
rect 476 1009 514 1037
rect 542 1009 580 1037
rect 608 1009 646 1037
rect 674 1009 712 1037
rect 740 1009 745 1037
rect -745 971 745 1009
rect -745 943 -740 971
rect -712 943 -674 971
rect -646 943 -608 971
rect -580 943 -542 971
rect -514 943 -476 971
rect -448 943 -410 971
rect -382 943 -344 971
rect -316 943 -278 971
rect -250 943 -212 971
rect -184 943 -146 971
rect -118 943 -80 971
rect -52 943 -14 971
rect 14 943 52 971
rect 80 943 118 971
rect 146 943 184 971
rect 212 943 250 971
rect 278 943 316 971
rect 344 943 382 971
rect 410 943 448 971
rect 476 943 514 971
rect 542 943 580 971
rect 608 943 646 971
rect 674 943 712 971
rect 740 943 745 971
rect -745 905 745 943
rect -745 877 -740 905
rect -712 877 -674 905
rect -646 877 -608 905
rect -580 877 -542 905
rect -514 877 -476 905
rect -448 877 -410 905
rect -382 877 -344 905
rect -316 877 -278 905
rect -250 877 -212 905
rect -184 877 -146 905
rect -118 877 -80 905
rect -52 877 -14 905
rect 14 877 52 905
rect 80 877 118 905
rect 146 877 184 905
rect 212 877 250 905
rect 278 877 316 905
rect 344 877 382 905
rect 410 877 448 905
rect 476 877 514 905
rect 542 877 580 905
rect 608 877 646 905
rect 674 877 712 905
rect 740 877 745 905
rect -745 839 745 877
rect -745 811 -740 839
rect -712 811 -674 839
rect -646 811 -608 839
rect -580 811 -542 839
rect -514 811 -476 839
rect -448 811 -410 839
rect -382 811 -344 839
rect -316 811 -278 839
rect -250 811 -212 839
rect -184 811 -146 839
rect -118 811 -80 839
rect -52 811 -14 839
rect 14 811 52 839
rect 80 811 118 839
rect 146 811 184 839
rect 212 811 250 839
rect 278 811 316 839
rect 344 811 382 839
rect 410 811 448 839
rect 476 811 514 839
rect 542 811 580 839
rect 608 811 646 839
rect 674 811 712 839
rect 740 811 745 839
rect -745 773 745 811
rect -745 745 -740 773
rect -712 745 -674 773
rect -646 745 -608 773
rect -580 745 -542 773
rect -514 745 -476 773
rect -448 745 -410 773
rect -382 745 -344 773
rect -316 745 -278 773
rect -250 745 -212 773
rect -184 745 -146 773
rect -118 745 -80 773
rect -52 745 -14 773
rect 14 745 52 773
rect 80 745 118 773
rect 146 745 184 773
rect 212 745 250 773
rect 278 745 316 773
rect 344 745 382 773
rect 410 745 448 773
rect 476 745 514 773
rect 542 745 580 773
rect 608 745 646 773
rect 674 745 712 773
rect 740 745 745 773
rect -745 707 745 745
rect -745 679 -740 707
rect -712 679 -674 707
rect -646 679 -608 707
rect -580 679 -542 707
rect -514 679 -476 707
rect -448 679 -410 707
rect -382 679 -344 707
rect -316 679 -278 707
rect -250 679 -212 707
rect -184 679 -146 707
rect -118 679 -80 707
rect -52 679 -14 707
rect 14 679 52 707
rect 80 679 118 707
rect 146 679 184 707
rect 212 679 250 707
rect 278 679 316 707
rect 344 679 382 707
rect 410 679 448 707
rect 476 679 514 707
rect 542 679 580 707
rect 608 679 646 707
rect 674 679 712 707
rect 740 679 745 707
rect -745 641 745 679
rect -745 613 -740 641
rect -712 613 -674 641
rect -646 613 -608 641
rect -580 613 -542 641
rect -514 613 -476 641
rect -448 613 -410 641
rect -382 613 -344 641
rect -316 613 -278 641
rect -250 613 -212 641
rect -184 613 -146 641
rect -118 613 -80 641
rect -52 613 -14 641
rect 14 613 52 641
rect 80 613 118 641
rect 146 613 184 641
rect 212 613 250 641
rect 278 613 316 641
rect 344 613 382 641
rect 410 613 448 641
rect 476 613 514 641
rect 542 613 580 641
rect 608 613 646 641
rect 674 613 712 641
rect 740 613 745 641
rect -745 575 745 613
rect -745 547 -740 575
rect -712 547 -674 575
rect -646 547 -608 575
rect -580 547 -542 575
rect -514 547 -476 575
rect -448 547 -410 575
rect -382 547 -344 575
rect -316 547 -278 575
rect -250 547 -212 575
rect -184 547 -146 575
rect -118 547 -80 575
rect -52 547 -14 575
rect 14 547 52 575
rect 80 547 118 575
rect 146 547 184 575
rect 212 547 250 575
rect 278 547 316 575
rect 344 547 382 575
rect 410 547 448 575
rect 476 547 514 575
rect 542 547 580 575
rect 608 547 646 575
rect 674 547 712 575
rect 740 547 745 575
rect -745 509 745 547
rect -745 481 -740 509
rect -712 481 -674 509
rect -646 481 -608 509
rect -580 481 -542 509
rect -514 481 -476 509
rect -448 481 -410 509
rect -382 481 -344 509
rect -316 481 -278 509
rect -250 481 -212 509
rect -184 481 -146 509
rect -118 481 -80 509
rect -52 481 -14 509
rect 14 481 52 509
rect 80 481 118 509
rect 146 481 184 509
rect 212 481 250 509
rect 278 481 316 509
rect 344 481 382 509
rect 410 481 448 509
rect 476 481 514 509
rect 542 481 580 509
rect 608 481 646 509
rect 674 481 712 509
rect 740 481 745 509
rect -745 443 745 481
rect -745 415 -740 443
rect -712 415 -674 443
rect -646 415 -608 443
rect -580 415 -542 443
rect -514 415 -476 443
rect -448 415 -410 443
rect -382 415 -344 443
rect -316 415 -278 443
rect -250 415 -212 443
rect -184 415 -146 443
rect -118 415 -80 443
rect -52 415 -14 443
rect 14 415 52 443
rect 80 415 118 443
rect 146 415 184 443
rect 212 415 250 443
rect 278 415 316 443
rect 344 415 382 443
rect 410 415 448 443
rect 476 415 514 443
rect 542 415 580 443
rect 608 415 646 443
rect 674 415 712 443
rect 740 415 745 443
rect -745 377 745 415
rect -745 349 -740 377
rect -712 349 -674 377
rect -646 349 -608 377
rect -580 349 -542 377
rect -514 349 -476 377
rect -448 349 -410 377
rect -382 349 -344 377
rect -316 349 -278 377
rect -250 349 -212 377
rect -184 349 -146 377
rect -118 349 -80 377
rect -52 349 -14 377
rect 14 349 52 377
rect 80 349 118 377
rect 146 349 184 377
rect 212 349 250 377
rect 278 349 316 377
rect 344 349 382 377
rect 410 349 448 377
rect 476 349 514 377
rect 542 349 580 377
rect 608 349 646 377
rect 674 349 712 377
rect 740 349 745 377
rect -745 311 745 349
rect -745 283 -740 311
rect -712 283 -674 311
rect -646 283 -608 311
rect -580 283 -542 311
rect -514 283 -476 311
rect -448 283 -410 311
rect -382 283 -344 311
rect -316 283 -278 311
rect -250 283 -212 311
rect -184 283 -146 311
rect -118 283 -80 311
rect -52 283 -14 311
rect 14 283 52 311
rect 80 283 118 311
rect 146 283 184 311
rect 212 283 250 311
rect 278 283 316 311
rect 344 283 382 311
rect 410 283 448 311
rect 476 283 514 311
rect 542 283 580 311
rect 608 283 646 311
rect 674 283 712 311
rect 740 283 745 311
rect -745 245 745 283
rect -745 217 -740 245
rect -712 217 -674 245
rect -646 217 -608 245
rect -580 217 -542 245
rect -514 217 -476 245
rect -448 217 -410 245
rect -382 217 -344 245
rect -316 217 -278 245
rect -250 217 -212 245
rect -184 217 -146 245
rect -118 217 -80 245
rect -52 217 -14 245
rect 14 217 52 245
rect 80 217 118 245
rect 146 217 184 245
rect 212 217 250 245
rect 278 217 316 245
rect 344 217 382 245
rect 410 217 448 245
rect 476 217 514 245
rect 542 217 580 245
rect 608 217 646 245
rect 674 217 712 245
rect 740 217 745 245
rect -745 179 745 217
rect -745 151 -740 179
rect -712 151 -674 179
rect -646 151 -608 179
rect -580 151 -542 179
rect -514 151 -476 179
rect -448 151 -410 179
rect -382 151 -344 179
rect -316 151 -278 179
rect -250 151 -212 179
rect -184 151 -146 179
rect -118 151 -80 179
rect -52 151 -14 179
rect 14 151 52 179
rect 80 151 118 179
rect 146 151 184 179
rect 212 151 250 179
rect 278 151 316 179
rect 344 151 382 179
rect 410 151 448 179
rect 476 151 514 179
rect 542 151 580 179
rect 608 151 646 179
rect 674 151 712 179
rect 740 151 745 179
rect -745 113 745 151
rect -745 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 745 113
rect -745 47 745 85
rect -745 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 745 47
rect -745 -19 745 19
rect -745 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 745 -19
rect -745 -85 745 -47
rect -745 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 745 -85
rect -745 -151 745 -113
rect -745 -179 -740 -151
rect -712 -179 -674 -151
rect -646 -179 -608 -151
rect -580 -179 -542 -151
rect -514 -179 -476 -151
rect -448 -179 -410 -151
rect -382 -179 -344 -151
rect -316 -179 -278 -151
rect -250 -179 -212 -151
rect -184 -179 -146 -151
rect -118 -179 -80 -151
rect -52 -179 -14 -151
rect 14 -179 52 -151
rect 80 -179 118 -151
rect 146 -179 184 -151
rect 212 -179 250 -151
rect 278 -179 316 -151
rect 344 -179 382 -151
rect 410 -179 448 -151
rect 476 -179 514 -151
rect 542 -179 580 -151
rect 608 -179 646 -151
rect 674 -179 712 -151
rect 740 -179 745 -151
rect -745 -217 745 -179
rect -745 -245 -740 -217
rect -712 -245 -674 -217
rect -646 -245 -608 -217
rect -580 -245 -542 -217
rect -514 -245 -476 -217
rect -448 -245 -410 -217
rect -382 -245 -344 -217
rect -316 -245 -278 -217
rect -250 -245 -212 -217
rect -184 -245 -146 -217
rect -118 -245 -80 -217
rect -52 -245 -14 -217
rect 14 -245 52 -217
rect 80 -245 118 -217
rect 146 -245 184 -217
rect 212 -245 250 -217
rect 278 -245 316 -217
rect 344 -245 382 -217
rect 410 -245 448 -217
rect 476 -245 514 -217
rect 542 -245 580 -217
rect 608 -245 646 -217
rect 674 -245 712 -217
rect 740 -245 745 -217
rect -745 -283 745 -245
rect -745 -311 -740 -283
rect -712 -311 -674 -283
rect -646 -311 -608 -283
rect -580 -311 -542 -283
rect -514 -311 -476 -283
rect -448 -311 -410 -283
rect -382 -311 -344 -283
rect -316 -311 -278 -283
rect -250 -311 -212 -283
rect -184 -311 -146 -283
rect -118 -311 -80 -283
rect -52 -311 -14 -283
rect 14 -311 52 -283
rect 80 -311 118 -283
rect 146 -311 184 -283
rect 212 -311 250 -283
rect 278 -311 316 -283
rect 344 -311 382 -283
rect 410 -311 448 -283
rect 476 -311 514 -283
rect 542 -311 580 -283
rect 608 -311 646 -283
rect 674 -311 712 -283
rect 740 -311 745 -283
rect -745 -349 745 -311
rect -745 -377 -740 -349
rect -712 -377 -674 -349
rect -646 -377 -608 -349
rect -580 -377 -542 -349
rect -514 -377 -476 -349
rect -448 -377 -410 -349
rect -382 -377 -344 -349
rect -316 -377 -278 -349
rect -250 -377 -212 -349
rect -184 -377 -146 -349
rect -118 -377 -80 -349
rect -52 -377 -14 -349
rect 14 -377 52 -349
rect 80 -377 118 -349
rect 146 -377 184 -349
rect 212 -377 250 -349
rect 278 -377 316 -349
rect 344 -377 382 -349
rect 410 -377 448 -349
rect 476 -377 514 -349
rect 542 -377 580 -349
rect 608 -377 646 -349
rect 674 -377 712 -349
rect 740 -377 745 -349
rect -745 -415 745 -377
rect -745 -443 -740 -415
rect -712 -443 -674 -415
rect -646 -443 -608 -415
rect -580 -443 -542 -415
rect -514 -443 -476 -415
rect -448 -443 -410 -415
rect -382 -443 -344 -415
rect -316 -443 -278 -415
rect -250 -443 -212 -415
rect -184 -443 -146 -415
rect -118 -443 -80 -415
rect -52 -443 -14 -415
rect 14 -443 52 -415
rect 80 -443 118 -415
rect 146 -443 184 -415
rect 212 -443 250 -415
rect 278 -443 316 -415
rect 344 -443 382 -415
rect 410 -443 448 -415
rect 476 -443 514 -415
rect 542 -443 580 -415
rect 608 -443 646 -415
rect 674 -443 712 -415
rect 740 -443 745 -415
rect -745 -481 745 -443
rect -745 -509 -740 -481
rect -712 -509 -674 -481
rect -646 -509 -608 -481
rect -580 -509 -542 -481
rect -514 -509 -476 -481
rect -448 -509 -410 -481
rect -382 -509 -344 -481
rect -316 -509 -278 -481
rect -250 -509 -212 -481
rect -184 -509 -146 -481
rect -118 -509 -80 -481
rect -52 -509 -14 -481
rect 14 -509 52 -481
rect 80 -509 118 -481
rect 146 -509 184 -481
rect 212 -509 250 -481
rect 278 -509 316 -481
rect 344 -509 382 -481
rect 410 -509 448 -481
rect 476 -509 514 -481
rect 542 -509 580 -481
rect 608 -509 646 -481
rect 674 -509 712 -481
rect 740 -509 745 -481
rect -745 -547 745 -509
rect -745 -575 -740 -547
rect -712 -575 -674 -547
rect -646 -575 -608 -547
rect -580 -575 -542 -547
rect -514 -575 -476 -547
rect -448 -575 -410 -547
rect -382 -575 -344 -547
rect -316 -575 -278 -547
rect -250 -575 -212 -547
rect -184 -575 -146 -547
rect -118 -575 -80 -547
rect -52 -575 -14 -547
rect 14 -575 52 -547
rect 80 -575 118 -547
rect 146 -575 184 -547
rect 212 -575 250 -547
rect 278 -575 316 -547
rect 344 -575 382 -547
rect 410 -575 448 -547
rect 476 -575 514 -547
rect 542 -575 580 -547
rect 608 -575 646 -547
rect 674 -575 712 -547
rect 740 -575 745 -547
rect -745 -613 745 -575
rect -745 -641 -740 -613
rect -712 -641 -674 -613
rect -646 -641 -608 -613
rect -580 -641 -542 -613
rect -514 -641 -476 -613
rect -448 -641 -410 -613
rect -382 -641 -344 -613
rect -316 -641 -278 -613
rect -250 -641 -212 -613
rect -184 -641 -146 -613
rect -118 -641 -80 -613
rect -52 -641 -14 -613
rect 14 -641 52 -613
rect 80 -641 118 -613
rect 146 -641 184 -613
rect 212 -641 250 -613
rect 278 -641 316 -613
rect 344 -641 382 -613
rect 410 -641 448 -613
rect 476 -641 514 -613
rect 542 -641 580 -613
rect 608 -641 646 -613
rect 674 -641 712 -613
rect 740 -641 745 -613
rect -745 -679 745 -641
rect -745 -707 -740 -679
rect -712 -707 -674 -679
rect -646 -707 -608 -679
rect -580 -707 -542 -679
rect -514 -707 -476 -679
rect -448 -707 -410 -679
rect -382 -707 -344 -679
rect -316 -707 -278 -679
rect -250 -707 -212 -679
rect -184 -707 -146 -679
rect -118 -707 -80 -679
rect -52 -707 -14 -679
rect 14 -707 52 -679
rect 80 -707 118 -679
rect 146 -707 184 -679
rect 212 -707 250 -679
rect 278 -707 316 -679
rect 344 -707 382 -679
rect 410 -707 448 -679
rect 476 -707 514 -679
rect 542 -707 580 -679
rect 608 -707 646 -679
rect 674 -707 712 -679
rect 740 -707 745 -679
rect -745 -745 745 -707
rect -745 -773 -740 -745
rect -712 -773 -674 -745
rect -646 -773 -608 -745
rect -580 -773 -542 -745
rect -514 -773 -476 -745
rect -448 -773 -410 -745
rect -382 -773 -344 -745
rect -316 -773 -278 -745
rect -250 -773 -212 -745
rect -184 -773 -146 -745
rect -118 -773 -80 -745
rect -52 -773 -14 -745
rect 14 -773 52 -745
rect 80 -773 118 -745
rect 146 -773 184 -745
rect 212 -773 250 -745
rect 278 -773 316 -745
rect 344 -773 382 -745
rect 410 -773 448 -745
rect 476 -773 514 -745
rect 542 -773 580 -745
rect 608 -773 646 -745
rect 674 -773 712 -745
rect 740 -773 745 -745
rect -745 -811 745 -773
rect -745 -839 -740 -811
rect -712 -839 -674 -811
rect -646 -839 -608 -811
rect -580 -839 -542 -811
rect -514 -839 -476 -811
rect -448 -839 -410 -811
rect -382 -839 -344 -811
rect -316 -839 -278 -811
rect -250 -839 -212 -811
rect -184 -839 -146 -811
rect -118 -839 -80 -811
rect -52 -839 -14 -811
rect 14 -839 52 -811
rect 80 -839 118 -811
rect 146 -839 184 -811
rect 212 -839 250 -811
rect 278 -839 316 -811
rect 344 -839 382 -811
rect 410 -839 448 -811
rect 476 -839 514 -811
rect 542 -839 580 -811
rect 608 -839 646 -811
rect 674 -839 712 -811
rect 740 -839 745 -811
rect -745 -877 745 -839
rect -745 -905 -740 -877
rect -712 -905 -674 -877
rect -646 -905 -608 -877
rect -580 -905 -542 -877
rect -514 -905 -476 -877
rect -448 -905 -410 -877
rect -382 -905 -344 -877
rect -316 -905 -278 -877
rect -250 -905 -212 -877
rect -184 -905 -146 -877
rect -118 -905 -80 -877
rect -52 -905 -14 -877
rect 14 -905 52 -877
rect 80 -905 118 -877
rect 146 -905 184 -877
rect 212 -905 250 -877
rect 278 -905 316 -877
rect 344 -905 382 -877
rect 410 -905 448 -877
rect 476 -905 514 -877
rect 542 -905 580 -877
rect 608 -905 646 -877
rect 674 -905 712 -877
rect 740 -905 745 -877
rect -745 -943 745 -905
rect -745 -971 -740 -943
rect -712 -971 -674 -943
rect -646 -971 -608 -943
rect -580 -971 -542 -943
rect -514 -971 -476 -943
rect -448 -971 -410 -943
rect -382 -971 -344 -943
rect -316 -971 -278 -943
rect -250 -971 -212 -943
rect -184 -971 -146 -943
rect -118 -971 -80 -943
rect -52 -971 -14 -943
rect 14 -971 52 -943
rect 80 -971 118 -943
rect 146 -971 184 -943
rect 212 -971 250 -943
rect 278 -971 316 -943
rect 344 -971 382 -943
rect 410 -971 448 -943
rect 476 -971 514 -943
rect 542 -971 580 -943
rect 608 -971 646 -943
rect 674 -971 712 -943
rect 740 -971 745 -943
rect -745 -1009 745 -971
rect -745 -1037 -740 -1009
rect -712 -1037 -674 -1009
rect -646 -1037 -608 -1009
rect -580 -1037 -542 -1009
rect -514 -1037 -476 -1009
rect -448 -1037 -410 -1009
rect -382 -1037 -344 -1009
rect -316 -1037 -278 -1009
rect -250 -1037 -212 -1009
rect -184 -1037 -146 -1009
rect -118 -1037 -80 -1009
rect -52 -1037 -14 -1009
rect 14 -1037 52 -1009
rect 80 -1037 118 -1009
rect 146 -1037 184 -1009
rect 212 -1037 250 -1009
rect 278 -1037 316 -1009
rect 344 -1037 382 -1009
rect 410 -1037 448 -1009
rect 476 -1037 514 -1009
rect 542 -1037 580 -1009
rect 608 -1037 646 -1009
rect 674 -1037 712 -1009
rect 740 -1037 745 -1009
rect -745 -1075 745 -1037
rect -745 -1103 -740 -1075
rect -712 -1103 -674 -1075
rect -646 -1103 -608 -1075
rect -580 -1103 -542 -1075
rect -514 -1103 -476 -1075
rect -448 -1103 -410 -1075
rect -382 -1103 -344 -1075
rect -316 -1103 -278 -1075
rect -250 -1103 -212 -1075
rect -184 -1103 -146 -1075
rect -118 -1103 -80 -1075
rect -52 -1103 -14 -1075
rect 14 -1103 52 -1075
rect 80 -1103 118 -1075
rect 146 -1103 184 -1075
rect 212 -1103 250 -1075
rect 278 -1103 316 -1075
rect 344 -1103 382 -1075
rect 410 -1103 448 -1075
rect 476 -1103 514 -1075
rect 542 -1103 580 -1075
rect 608 -1103 646 -1075
rect 674 -1103 712 -1075
rect 740 -1103 745 -1075
rect -745 -1141 745 -1103
rect -745 -1169 -740 -1141
rect -712 -1169 -674 -1141
rect -646 -1169 -608 -1141
rect -580 -1169 -542 -1141
rect -514 -1169 -476 -1141
rect -448 -1169 -410 -1141
rect -382 -1169 -344 -1141
rect -316 -1169 -278 -1141
rect -250 -1169 -212 -1141
rect -184 -1169 -146 -1141
rect -118 -1169 -80 -1141
rect -52 -1169 -14 -1141
rect 14 -1169 52 -1141
rect 80 -1169 118 -1141
rect 146 -1169 184 -1141
rect 212 -1169 250 -1141
rect 278 -1169 316 -1141
rect 344 -1169 382 -1141
rect 410 -1169 448 -1141
rect 476 -1169 514 -1141
rect 542 -1169 580 -1141
rect 608 -1169 646 -1141
rect 674 -1169 712 -1141
rect 740 -1169 745 -1141
rect -745 -1207 745 -1169
rect -745 -1235 -740 -1207
rect -712 -1235 -674 -1207
rect -646 -1235 -608 -1207
rect -580 -1235 -542 -1207
rect -514 -1235 -476 -1207
rect -448 -1235 -410 -1207
rect -382 -1235 -344 -1207
rect -316 -1235 -278 -1207
rect -250 -1235 -212 -1207
rect -184 -1235 -146 -1207
rect -118 -1235 -80 -1207
rect -52 -1235 -14 -1207
rect 14 -1235 52 -1207
rect 80 -1235 118 -1207
rect 146 -1235 184 -1207
rect 212 -1235 250 -1207
rect 278 -1235 316 -1207
rect 344 -1235 382 -1207
rect 410 -1235 448 -1207
rect 476 -1235 514 -1207
rect 542 -1235 580 -1207
rect 608 -1235 646 -1207
rect 674 -1235 712 -1207
rect 740 -1235 745 -1207
rect -745 -1273 745 -1235
rect -745 -1301 -740 -1273
rect -712 -1301 -674 -1273
rect -646 -1301 -608 -1273
rect -580 -1301 -542 -1273
rect -514 -1301 -476 -1273
rect -448 -1301 -410 -1273
rect -382 -1301 -344 -1273
rect -316 -1301 -278 -1273
rect -250 -1301 -212 -1273
rect -184 -1301 -146 -1273
rect -118 -1301 -80 -1273
rect -52 -1301 -14 -1273
rect 14 -1301 52 -1273
rect 80 -1301 118 -1273
rect 146 -1301 184 -1273
rect 212 -1301 250 -1273
rect 278 -1301 316 -1273
rect 344 -1301 382 -1273
rect 410 -1301 448 -1273
rect 476 -1301 514 -1273
rect 542 -1301 580 -1273
rect 608 -1301 646 -1273
rect 674 -1301 712 -1273
rect 740 -1301 745 -1273
rect -745 -1339 745 -1301
rect -745 -1367 -740 -1339
rect -712 -1367 -674 -1339
rect -646 -1367 -608 -1339
rect -580 -1367 -542 -1339
rect -514 -1367 -476 -1339
rect -448 -1367 -410 -1339
rect -382 -1367 -344 -1339
rect -316 -1367 -278 -1339
rect -250 -1367 -212 -1339
rect -184 -1367 -146 -1339
rect -118 -1367 -80 -1339
rect -52 -1367 -14 -1339
rect 14 -1367 52 -1339
rect 80 -1367 118 -1339
rect 146 -1367 184 -1339
rect 212 -1367 250 -1339
rect 278 -1367 316 -1339
rect 344 -1367 382 -1339
rect 410 -1367 448 -1339
rect 476 -1367 514 -1339
rect 542 -1367 580 -1339
rect 608 -1367 646 -1339
rect 674 -1367 712 -1339
rect 740 -1367 745 -1339
rect -745 -1405 745 -1367
rect -745 -1433 -740 -1405
rect -712 -1433 -674 -1405
rect -646 -1433 -608 -1405
rect -580 -1433 -542 -1405
rect -514 -1433 -476 -1405
rect -448 -1433 -410 -1405
rect -382 -1433 -344 -1405
rect -316 -1433 -278 -1405
rect -250 -1433 -212 -1405
rect -184 -1433 -146 -1405
rect -118 -1433 -80 -1405
rect -52 -1433 -14 -1405
rect 14 -1433 52 -1405
rect 80 -1433 118 -1405
rect 146 -1433 184 -1405
rect 212 -1433 250 -1405
rect 278 -1433 316 -1405
rect 344 -1433 382 -1405
rect 410 -1433 448 -1405
rect 476 -1433 514 -1405
rect 542 -1433 580 -1405
rect 608 -1433 646 -1405
rect 674 -1433 712 -1405
rect 740 -1433 745 -1405
rect -745 -1471 745 -1433
rect -745 -1499 -740 -1471
rect -712 -1499 -674 -1471
rect -646 -1499 -608 -1471
rect -580 -1499 -542 -1471
rect -514 -1499 -476 -1471
rect -448 -1499 -410 -1471
rect -382 -1499 -344 -1471
rect -316 -1499 -278 -1471
rect -250 -1499 -212 -1471
rect -184 -1499 -146 -1471
rect -118 -1499 -80 -1471
rect -52 -1499 -14 -1471
rect 14 -1499 52 -1471
rect 80 -1499 118 -1471
rect 146 -1499 184 -1471
rect 212 -1499 250 -1471
rect 278 -1499 316 -1471
rect 344 -1499 382 -1471
rect 410 -1499 448 -1471
rect 476 -1499 514 -1471
rect 542 -1499 580 -1471
rect 608 -1499 646 -1471
rect 674 -1499 712 -1471
rect 740 -1499 745 -1471
rect -745 -1537 745 -1499
rect -745 -1565 -740 -1537
rect -712 -1565 -674 -1537
rect -646 -1565 -608 -1537
rect -580 -1565 -542 -1537
rect -514 -1565 -476 -1537
rect -448 -1565 -410 -1537
rect -382 -1565 -344 -1537
rect -316 -1565 -278 -1537
rect -250 -1565 -212 -1537
rect -184 -1565 -146 -1537
rect -118 -1565 -80 -1537
rect -52 -1565 -14 -1537
rect 14 -1565 52 -1537
rect 80 -1565 118 -1537
rect 146 -1565 184 -1537
rect 212 -1565 250 -1537
rect 278 -1565 316 -1537
rect 344 -1565 382 -1537
rect 410 -1565 448 -1537
rect 476 -1565 514 -1537
rect 542 -1565 580 -1537
rect 608 -1565 646 -1537
rect 674 -1565 712 -1537
rect 740 -1565 745 -1537
rect -745 -1603 745 -1565
rect -745 -1631 -740 -1603
rect -712 -1631 -674 -1603
rect -646 -1631 -608 -1603
rect -580 -1631 -542 -1603
rect -514 -1631 -476 -1603
rect -448 -1631 -410 -1603
rect -382 -1631 -344 -1603
rect -316 -1631 -278 -1603
rect -250 -1631 -212 -1603
rect -184 -1631 -146 -1603
rect -118 -1631 -80 -1603
rect -52 -1631 -14 -1603
rect 14 -1631 52 -1603
rect 80 -1631 118 -1603
rect 146 -1631 184 -1603
rect 212 -1631 250 -1603
rect 278 -1631 316 -1603
rect 344 -1631 382 -1603
rect 410 -1631 448 -1603
rect 476 -1631 514 -1603
rect 542 -1631 580 -1603
rect 608 -1631 646 -1603
rect 674 -1631 712 -1603
rect 740 -1631 745 -1603
rect -745 -1669 745 -1631
rect -745 -1697 -740 -1669
rect -712 -1697 -674 -1669
rect -646 -1697 -608 -1669
rect -580 -1697 -542 -1669
rect -514 -1697 -476 -1669
rect -448 -1697 -410 -1669
rect -382 -1697 -344 -1669
rect -316 -1697 -278 -1669
rect -250 -1697 -212 -1669
rect -184 -1697 -146 -1669
rect -118 -1697 -80 -1669
rect -52 -1697 -14 -1669
rect 14 -1697 52 -1669
rect 80 -1697 118 -1669
rect 146 -1697 184 -1669
rect 212 -1697 250 -1669
rect 278 -1697 316 -1669
rect 344 -1697 382 -1669
rect 410 -1697 448 -1669
rect 476 -1697 514 -1669
rect 542 -1697 580 -1669
rect 608 -1697 646 -1669
rect 674 -1697 712 -1669
rect 740 -1697 745 -1669
rect -745 -1735 745 -1697
rect -745 -1763 -740 -1735
rect -712 -1763 -674 -1735
rect -646 -1763 -608 -1735
rect -580 -1763 -542 -1735
rect -514 -1763 -476 -1735
rect -448 -1763 -410 -1735
rect -382 -1763 -344 -1735
rect -316 -1763 -278 -1735
rect -250 -1763 -212 -1735
rect -184 -1763 -146 -1735
rect -118 -1763 -80 -1735
rect -52 -1763 -14 -1735
rect 14 -1763 52 -1735
rect 80 -1763 118 -1735
rect 146 -1763 184 -1735
rect 212 -1763 250 -1735
rect 278 -1763 316 -1735
rect 344 -1763 382 -1735
rect 410 -1763 448 -1735
rect 476 -1763 514 -1735
rect 542 -1763 580 -1735
rect 608 -1763 646 -1735
rect 674 -1763 712 -1735
rect 740 -1763 745 -1735
rect -745 -1801 745 -1763
rect -745 -1829 -740 -1801
rect -712 -1829 -674 -1801
rect -646 -1829 -608 -1801
rect -580 -1829 -542 -1801
rect -514 -1829 -476 -1801
rect -448 -1829 -410 -1801
rect -382 -1829 -344 -1801
rect -316 -1829 -278 -1801
rect -250 -1829 -212 -1801
rect -184 -1829 -146 -1801
rect -118 -1829 -80 -1801
rect -52 -1829 -14 -1801
rect 14 -1829 52 -1801
rect 80 -1829 118 -1801
rect 146 -1829 184 -1801
rect 212 -1829 250 -1801
rect 278 -1829 316 -1801
rect 344 -1829 382 -1801
rect 410 -1829 448 -1801
rect 476 -1829 514 -1801
rect 542 -1829 580 -1801
rect 608 -1829 646 -1801
rect 674 -1829 712 -1801
rect 740 -1829 745 -1801
rect -745 -1867 745 -1829
rect -745 -1895 -740 -1867
rect -712 -1895 -674 -1867
rect -646 -1895 -608 -1867
rect -580 -1895 -542 -1867
rect -514 -1895 -476 -1867
rect -448 -1895 -410 -1867
rect -382 -1895 -344 -1867
rect -316 -1895 -278 -1867
rect -250 -1895 -212 -1867
rect -184 -1895 -146 -1867
rect -118 -1895 -80 -1867
rect -52 -1895 -14 -1867
rect 14 -1895 52 -1867
rect 80 -1895 118 -1867
rect 146 -1895 184 -1867
rect 212 -1895 250 -1867
rect 278 -1895 316 -1867
rect 344 -1895 382 -1867
rect 410 -1895 448 -1867
rect 476 -1895 514 -1867
rect 542 -1895 580 -1867
rect 608 -1895 646 -1867
rect 674 -1895 712 -1867
rect 740 -1895 745 -1867
rect -745 -1933 745 -1895
rect -745 -1961 -740 -1933
rect -712 -1961 -674 -1933
rect -646 -1961 -608 -1933
rect -580 -1961 -542 -1933
rect -514 -1961 -476 -1933
rect -448 -1961 -410 -1933
rect -382 -1961 -344 -1933
rect -316 -1961 -278 -1933
rect -250 -1961 -212 -1933
rect -184 -1961 -146 -1933
rect -118 -1961 -80 -1933
rect -52 -1961 -14 -1933
rect 14 -1961 52 -1933
rect 80 -1961 118 -1933
rect 146 -1961 184 -1933
rect 212 -1961 250 -1933
rect 278 -1961 316 -1933
rect 344 -1961 382 -1933
rect 410 -1961 448 -1933
rect 476 -1961 514 -1933
rect 542 -1961 580 -1933
rect 608 -1961 646 -1933
rect 674 -1961 712 -1933
rect 740 -1961 745 -1933
rect -745 -1999 745 -1961
rect -745 -2027 -740 -1999
rect -712 -2027 -674 -1999
rect -646 -2027 -608 -1999
rect -580 -2027 -542 -1999
rect -514 -2027 -476 -1999
rect -448 -2027 -410 -1999
rect -382 -2027 -344 -1999
rect -316 -2027 -278 -1999
rect -250 -2027 -212 -1999
rect -184 -2027 -146 -1999
rect -118 -2027 -80 -1999
rect -52 -2027 -14 -1999
rect 14 -2027 52 -1999
rect 80 -2027 118 -1999
rect 146 -2027 184 -1999
rect 212 -2027 250 -1999
rect 278 -2027 316 -1999
rect 344 -2027 382 -1999
rect 410 -2027 448 -1999
rect 476 -2027 514 -1999
rect 542 -2027 580 -1999
rect 608 -2027 646 -1999
rect 674 -2027 712 -1999
rect 740 -2027 745 -1999
rect -745 -2065 745 -2027
rect -745 -2093 -740 -2065
rect -712 -2093 -674 -2065
rect -646 -2093 -608 -2065
rect -580 -2093 -542 -2065
rect -514 -2093 -476 -2065
rect -448 -2093 -410 -2065
rect -382 -2093 -344 -2065
rect -316 -2093 -278 -2065
rect -250 -2093 -212 -2065
rect -184 -2093 -146 -2065
rect -118 -2093 -80 -2065
rect -52 -2093 -14 -2065
rect 14 -2093 52 -2065
rect 80 -2093 118 -2065
rect 146 -2093 184 -2065
rect 212 -2093 250 -2065
rect 278 -2093 316 -2065
rect 344 -2093 382 -2065
rect 410 -2093 448 -2065
rect 476 -2093 514 -2065
rect 542 -2093 580 -2065
rect 608 -2093 646 -2065
rect 674 -2093 712 -2065
rect 740 -2093 745 -2065
rect -745 -2131 745 -2093
rect -745 -2159 -740 -2131
rect -712 -2159 -674 -2131
rect -646 -2159 -608 -2131
rect -580 -2159 -542 -2131
rect -514 -2159 -476 -2131
rect -448 -2159 -410 -2131
rect -382 -2159 -344 -2131
rect -316 -2159 -278 -2131
rect -250 -2159 -212 -2131
rect -184 -2159 -146 -2131
rect -118 -2159 -80 -2131
rect -52 -2159 -14 -2131
rect 14 -2159 52 -2131
rect 80 -2159 118 -2131
rect 146 -2159 184 -2131
rect 212 -2159 250 -2131
rect 278 -2159 316 -2131
rect 344 -2159 382 -2131
rect 410 -2159 448 -2131
rect 476 -2159 514 -2131
rect 542 -2159 580 -2131
rect 608 -2159 646 -2131
rect 674 -2159 712 -2131
rect 740 -2159 745 -2131
rect -745 -2197 745 -2159
rect -745 -2225 -740 -2197
rect -712 -2225 -674 -2197
rect -646 -2225 -608 -2197
rect -580 -2225 -542 -2197
rect -514 -2225 -476 -2197
rect -448 -2225 -410 -2197
rect -382 -2225 -344 -2197
rect -316 -2225 -278 -2197
rect -250 -2225 -212 -2197
rect -184 -2225 -146 -2197
rect -118 -2225 -80 -2197
rect -52 -2225 -14 -2197
rect 14 -2225 52 -2197
rect 80 -2225 118 -2197
rect 146 -2225 184 -2197
rect 212 -2225 250 -2197
rect 278 -2225 316 -2197
rect 344 -2225 382 -2197
rect 410 -2225 448 -2197
rect 476 -2225 514 -2197
rect 542 -2225 580 -2197
rect 608 -2225 646 -2197
rect 674 -2225 712 -2197
rect 740 -2225 745 -2197
rect -745 -2263 745 -2225
rect -745 -2291 -740 -2263
rect -712 -2291 -674 -2263
rect -646 -2291 -608 -2263
rect -580 -2291 -542 -2263
rect -514 -2291 -476 -2263
rect -448 -2291 -410 -2263
rect -382 -2291 -344 -2263
rect -316 -2291 -278 -2263
rect -250 -2291 -212 -2263
rect -184 -2291 -146 -2263
rect -118 -2291 -80 -2263
rect -52 -2291 -14 -2263
rect 14 -2291 52 -2263
rect 80 -2291 118 -2263
rect 146 -2291 184 -2263
rect 212 -2291 250 -2263
rect 278 -2291 316 -2263
rect 344 -2291 382 -2263
rect 410 -2291 448 -2263
rect 476 -2291 514 -2263
rect 542 -2291 580 -2263
rect 608 -2291 646 -2263
rect 674 -2291 712 -2263
rect 740 -2291 745 -2263
rect -745 -2329 745 -2291
rect -745 -2357 -740 -2329
rect -712 -2357 -674 -2329
rect -646 -2357 -608 -2329
rect -580 -2357 -542 -2329
rect -514 -2357 -476 -2329
rect -448 -2357 -410 -2329
rect -382 -2357 -344 -2329
rect -316 -2357 -278 -2329
rect -250 -2357 -212 -2329
rect -184 -2357 -146 -2329
rect -118 -2357 -80 -2329
rect -52 -2357 -14 -2329
rect 14 -2357 52 -2329
rect 80 -2357 118 -2329
rect 146 -2357 184 -2329
rect 212 -2357 250 -2329
rect 278 -2357 316 -2329
rect 344 -2357 382 -2329
rect 410 -2357 448 -2329
rect 476 -2357 514 -2329
rect 542 -2357 580 -2329
rect 608 -2357 646 -2329
rect 674 -2357 712 -2329
rect 740 -2357 745 -2329
rect -745 -2395 745 -2357
rect -745 -2423 -740 -2395
rect -712 -2423 -674 -2395
rect -646 -2423 -608 -2395
rect -580 -2423 -542 -2395
rect -514 -2423 -476 -2395
rect -448 -2423 -410 -2395
rect -382 -2423 -344 -2395
rect -316 -2423 -278 -2395
rect -250 -2423 -212 -2395
rect -184 -2423 -146 -2395
rect -118 -2423 -80 -2395
rect -52 -2423 -14 -2395
rect 14 -2423 52 -2395
rect 80 -2423 118 -2395
rect 146 -2423 184 -2395
rect 212 -2423 250 -2395
rect 278 -2423 316 -2395
rect 344 -2423 382 -2395
rect 410 -2423 448 -2395
rect 476 -2423 514 -2395
rect 542 -2423 580 -2395
rect 608 -2423 646 -2395
rect 674 -2423 712 -2395
rect 740 -2423 745 -2395
rect -745 -2461 745 -2423
rect -745 -2489 -740 -2461
rect -712 -2489 -674 -2461
rect -646 -2489 -608 -2461
rect -580 -2489 -542 -2461
rect -514 -2489 -476 -2461
rect -448 -2489 -410 -2461
rect -382 -2489 -344 -2461
rect -316 -2489 -278 -2461
rect -250 -2489 -212 -2461
rect -184 -2489 -146 -2461
rect -118 -2489 -80 -2461
rect -52 -2489 -14 -2461
rect 14 -2489 52 -2461
rect 80 -2489 118 -2461
rect 146 -2489 184 -2461
rect 212 -2489 250 -2461
rect 278 -2489 316 -2461
rect 344 -2489 382 -2461
rect 410 -2489 448 -2461
rect 476 -2489 514 -2461
rect 542 -2489 580 -2461
rect 608 -2489 646 -2461
rect 674 -2489 712 -2461
rect 740 -2489 745 -2461
rect -745 -2527 745 -2489
rect -745 -2555 -740 -2527
rect -712 -2555 -674 -2527
rect -646 -2555 -608 -2527
rect -580 -2555 -542 -2527
rect -514 -2555 -476 -2527
rect -448 -2555 -410 -2527
rect -382 -2555 -344 -2527
rect -316 -2555 -278 -2527
rect -250 -2555 -212 -2527
rect -184 -2555 -146 -2527
rect -118 -2555 -80 -2527
rect -52 -2555 -14 -2527
rect 14 -2555 52 -2527
rect 80 -2555 118 -2527
rect 146 -2555 184 -2527
rect 212 -2555 250 -2527
rect 278 -2555 316 -2527
rect 344 -2555 382 -2527
rect 410 -2555 448 -2527
rect 476 -2555 514 -2527
rect 542 -2555 580 -2527
rect 608 -2555 646 -2527
rect 674 -2555 712 -2527
rect 740 -2555 745 -2527
rect -745 -2560 745 -2555
<< end >>
