magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1208 -1019 1208 1019
<< metal1 >>
rect -208 13 208 19
rect -208 -13 -202 13
rect -176 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 176 13
rect 202 -13 208 13
rect -208 -19 208 -13
<< via1 >>
rect -202 -13 -176 13
rect -148 -13 -122 13
rect -94 -13 -68 13
rect -40 -13 -14 13
rect 14 -13 40 13
rect 68 -13 94 13
rect 122 -13 148 13
rect 176 -13 202 13
<< metal2 >>
rect -208 13 208 19
rect -208 -13 -202 13
rect -176 -13 -148 13
rect -122 -13 -94 13
rect -68 -13 -40 13
rect -14 -13 14 13
rect 40 -13 68 13
rect 94 -13 122 13
rect 148 -13 176 13
rect 202 -13 208 13
rect -208 -19 208 -13
<< end >>
