* NGSPICE file created from MSB_Unit_Cell_flat.ext - technology: gf180mcuC

.subckt pex_MSB_Unit_Cell IOUT+ IOUT- VDD Ri-1 Ci Ri IM_T IM VSS 
X0 IOUT- Local_Enc_0.QB.t3 CM_MSB_V2_0.OUT.t66 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 CM_MSB_V2_0.OUT IM_T.t0 CM_MSB_V2_0.SD.t32 VSS.t39 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X2 IOUT+ Local_Enc_0.Q.t3 CM_MSB_V2_0.OUT.t150 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X3 VSS IM.t0 CM_MSB_V2_0.SD.t0 VSS.t13 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X4 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_6.B VDD.t27 VDD.t26 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X5 IOUT- Local_Enc_0.QB.t4 CM_MSB_V2_0.OUT.t65 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X6 IOUT+ Local_Enc_0.Q.t4 CM_MSB_V2_0.OUT.t151 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 CM_MSB_V2_0.OUT Local_Enc_0.Q.t5 IOUT+.t61 VSS.t44 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X8 IOUT- Local_Enc_0.QB.t5 CM_MSB_V2_0.OUT.t64 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 IOUT+ Local_Enc_0.Q.t6 CM_MSB_V2_0.OUT.t123 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X10 IOUT+ Local_Enc_0.Q.t7 CM_MSB_V2_0.OUT.t86 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X11 CM_MSB_V2_0.SD IM_T.t1 CM_MSB_V2_0.OUT.t85 VSS.t58 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X12 IOUT+ Local_Enc_0.Q.t8 CM_MSB_V2_0.OUT.t87 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X13 CM_MSB_V2_0.SD IM_T.t2 CM_MSB_V2_0.OUT.t0 VSS.t4 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X14 IOUT- Local_Enc_0.QB.t6 CM_MSB_V2_0.OUT.t63 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X15 CM_MSB_V2_0.OUT Local_Enc_0.QB.t7 IOUT-.t59 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X16 IOUT- Local_Enc_0.QB.t8 CM_MSB_V2_0.OUT.t62 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X17 CM_MSB_V2_0.OUT Local_Enc_0.QB.t9 IOUT-.t57 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X18 CM_MSB_V2_0.OUT Local_Enc_0.Q.t9 IOUT+.t57 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X19 CM_MSB_V2_0.SD IM_T.t3 CM_MSB_V2_0.OUT.t3 VSS.t9 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X20 CM_MSB_V2_0.OUT Local_Enc_0.Q.t10 IOUT+.t56 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X21 CM_MSB_V2_0.OUT Local_Enc_0.Q.t11 IOUT+.t55 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X22 CM_MSB_V2_0.OUT Local_Enc_0.Q.t12 IOUT+.t54 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X23 IOUT+ Local_Enc_0.Q.t13 CM_MSB_V2_0.OUT.t129 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X24 IOUT+ Local_Enc_0.Q.t14 CM_MSB_V2_0.OUT.t130 VSS.t40 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X25 CM_MSB_V2_0.OUT Local_Enc_0.Q.t15 IOUT+.t51 VSS.t46 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X26 CM_MSB_V2_0.OUT Local_Enc_0.QB.t10 IOUT-.t56 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X27 CM_MSB_V2_0.OUT Local_Enc_0.QB.t11 IOUT-.t55 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X28 IOUT- Local_Enc_0.QB.t12 CM_MSB_V2_0.OUT.t61 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X29 CM_MSB_V2_0.OUT IM_T.t4 CM_MSB_V2_0.SD.t28 VSS.t35 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X30 CM_MSB_V2_0.OUT Local_Enc_0.Q.t16 IOUT+.t50 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X31 CM_MSB_V2_0.OUT IM_T.t5 CM_MSB_V2_0.SD.t27 VSS.t21 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X32 IOUT+ Local_Enc_0.Q.t17 CM_MSB_V2_0.OUT.t88 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X33 CM_MSB_V2_0.OUT Local_Enc_0.Q.t18 IOUT+.t48 VSS.t44 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X34 VSS IM.t1 CM_MSB_V2_0.SD.t33 VSS.t6 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X35 CM_MSB_V2_0.SD IM_T.t6 CM_MSB_V2_0.OUT.t8 VSS.t14 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X36 IOUT+ Local_Enc_0.Q.t19 CM_MSB_V2_0.OUT.t120 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X37 CM_MSB_V2_0.OUT Local_Enc_0.QB.t13 IOUT-.t53 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X38 Local_Enc_0.Q Local_Enc_0.NAND_8.A a_n1035_4741# VSS.t3 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X39 CM_MSB_V2_0.OUT Local_Enc_0.Q.t20 IOUT+.t46 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X40 CM_MSB_V2_0.SD IM_T.t7 CM_MSB_V2_0.OUT.t16 VSS.t29 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X41 CM_MSB_V2_0.OUT IM_T.t8 CM_MSB_V2_0.SD.t24 VSS.t18 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X42 IOUT+ Local_Enc_0.Q.t21 CM_MSB_V2_0.OUT.t116 VSS.t40 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X43 a_n1035_4741# Local_Enc_0.QB.t14 VSS.t57 VSS.t56 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X44 IOUT+ Local_Enc_0.Q.t22 CM_MSB_V2_0.OUT.t117 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X45 CM_MSB_V2_0.OUT Local_Enc_0.QB.t15 IOUT-.t52 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X46 CM_MSB_V2_0.SD IM_T.t9 CM_MSB_V2_0.OUT.t103 VSS.t63 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X47 CM_MSB_V2_0.SD IM_T.t10 CM_MSB_V2_0.OUT.t102 VSS.t62 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X48 VSS IM.t2 CM_MSB_V2_0.SD.t62 VSS.t119 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X49 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_5.B VDD.t36 VDD.t35 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X50 IOUT- Local_Enc_0.QB.t16 CM_MSB_V2_0.OUT.t60 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X51 a_n1846_3765# Local_Enc_0.NAND_6.B VSS.t38 VSS.t37 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X52 IOUT+ Local_Enc_0.Q.t23 CM_MSB_V2_0.OUT.t132 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X53 CM_MSB_V2_0.SD IM.t3 VSS.t122 VSS.t20 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X54 IOUT+ Local_Enc_0.Q.t24 CM_MSB_V2_0.OUT.t133 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X55 IOUT+ Local_Enc_0.Q.t25 CM_MSB_V2_0.OUT.t104 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X56 CM_MSB_V2_0.OUT Local_Enc_0.QB.t17 IOUT-.t50 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X57 IOUT- Local_Enc_0.QB.t18 CM_MSB_V2_0.OUT.t59 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X58 IOUT- Local_Enc_0.QB.t19 CM_MSB_V2_0.OUT.t58 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X59 CM_MSB_V2_0.SD IM.t4 VSS.t69 VSS.t68 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X60 CM_MSB_V2_0.OUT Local_Enc_0.QB.t20 IOUT-.t47 VSS.t46 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X61 IOUT- Local_Enc_0.QB.t21 CM_MSB_V2_0.OUT.t57 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X62 CM_MSB_V2_0.SD IM.t5 VSS.t70 VSS.t10 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X63 CM_MSB_V2_0.OUT Local_Enc_0.Q.t26 IOUT+.t40 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X64 VDD Local_Enc_0.NAND_6.A Local_Enc_0.NAND_5.A VDD.t21 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X65 Local_Enc_0.NAND_6.B Ci.t0 VDD.t20 VDD.t19 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X66 VSS IM.t6 CM_MSB_V2_0.SD.t40 VSS.t11 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X67 CM_MSB_V2_0.OUT Local_Enc_0.Q.t27 IOUT+.t39 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X68 CM_MSB_V2_0.OUT Local_Enc_0.Q.t28 IOUT+.t38 VSS.t46 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X69 CM_MSB_V2_0.OUT IM_T.t11 CM_MSB_V2_0.SD.t21 VSS.t103 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X70 CM_MSB_V2_0.SD IM.t7 VSS.t82 VSS.t5 nfet_03v3 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X71 CM_MSB_V2_0.OUT Local_Enc_0.Q.t29 IOUT+.t37 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X72 CM_MSB_V2_0.OUT Local_Enc_0.QB.t22 IOUT-.t45 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X73 CM_MSB_V2_0.OUT Local_Enc_0.QB.t23 IOUT-.t44 VSS.t44 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X74 IOUT+ Local_Enc_0.Q.t30 CM_MSB_V2_0.OUT.t140 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X75 CM_MSB_V2_0.OUT Local_Enc_0.QB.t24 IOUT-.t43 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X76 CM_MSB_V2_0.OUT Local_Enc_0.QB.t25 IOUT-.t42 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X77 VDD Ci.t1 Local_Enc_0.NAND_6.B VDD.t28 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X78 CM_MSB_V2_0.OUT Local_Enc_0.Q.t31 IOUT+.t35 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X79 CM_MSB_V2_0.OUT Local_Enc_0.Q.t32 IOUT+.t34 VSS.t44 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X80 VSS IM.t8 CM_MSB_V2_0.SD.t60 VSS.t113 nfet_03v3 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
X81 IOUT+ Local_Enc_0.Q.t33 CM_MSB_V2_0.OUT.t96 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X82 VSS IM.t9 CM_MSB_V2_0.SD.t61 VSS.t116 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X83 IOUT+ Local_Enc_0.Q.t34 CM_MSB_V2_0.OUT.t97 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X84 CM_MSB_V2_0.OUT IM_T.t12 CM_MSB_V2_0.SD.t20 VSS.t73 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X85 CM_MSB_V2_0.SD IM_T.t13 CM_MSB_V2_0.OUT.t6 VSS.t12 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X86 CM_MSB_V2_0.OUT Local_Enc_0.QB.t26 IOUT-.t41 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X87 IOUT- Local_Enc_0.QB.t27 CM_MSB_V2_0.OUT.t56 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X88 IOUT- Local_Enc_0.QB.t28 CM_MSB_V2_0.OUT.t55 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X89 IOUT- Local_Enc_0.QB.t29 CM_MSB_V2_0.OUT.t54 VSS.t40 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X90 VSS IM.t10 CM_MSB_V2_0.SD.t52 VSS.t39 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X91 IOUT- Local_Enc_0.QB.t30 CM_MSB_V2_0.OUT.t53 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X92 CM_MSB_V2_0.OUT IM_T.t14 CM_MSB_V2_0.SD.t18 VSS.t13 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X93 IOUT+ Local_Enc_0.Q.t35 CM_MSB_V2_0.OUT.t131 VSS.t40 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X94 VDD Local_Enc_0.Q.t36 Local_Enc_0.QB.t1 VDD.t42 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X95 Local_Enc_0.QB Local_Enc_0.Q.t37 a_n1035_5712# VSS.t86 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X96 Local_Enc_0.NAND_6.A Ri.t0 VDD.t41 VDD.t40 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X97 a_n1035_5712# Local_Enc_0.NAND_4.B VSS.t65 VSS.t64 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X98 CM_MSB_V2_0.SD IM.t11 VSS.t102 VSS.t58 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X99 Local_Enc_0.QB Local_Enc_0.NAND_4.B VDD.t34 VDD.t33 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X100 IOUT- Local_Enc_0.QB.t31 CM_MSB_V2_0.OUT.t52 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X101 CM_MSB_V2_0.SD IM.t12 VSS.t111 VSS.t4 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X102 a_n1846_4741# Local_Enc_0.NAND_5.B VSS.t72 VSS.t71 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X103 IOUT- Local_Enc_0.QB.t32 CM_MSB_V2_0.OUT.t51 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X104 VDD Ri.t1 Local_Enc_0.NAND_6.A VDD.t37 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X105 CM_MSB_V2_0.OUT Local_Enc_0.Q.t38 IOUT+.t30 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X106 CM_MSB_V2_0.SD IM.t13 VSS.t112 VSS.t9 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X107 CM_MSB_V2_0.SD IM_T.t15 CM_MSB_V2_0.OUT.t10 VSS.t16 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X108 VSS IM.t14 CM_MSB_V2_0.SD.t51 VSS.t97 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X109 IOUT- Local_Enc_0.QB.t33 CM_MSB_V2_0.OUT.t50 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X110 CM_MSB_V2_0.OUT Local_Enc_0.QB.t34 IOUT-.t33 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X111 CM_MSB_V2_0.OUT Local_Enc_0.Q.t39 IOUT+.t29 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X112 CM_MSB_V2_0.SD IM_T.t16 CM_MSB_V2_0.OUT.t11 VSS.t17 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X113 CM_MSB_V2_0.OUT Local_Enc_0.QB.t35 IOUT-.t32 VSS.t46 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X114 VDD Local_Enc_0.NAND_5.A Local_Enc_0.NAND_8.A VDD.t11 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X115 CM_MSB_V2_0.OUT Local_Enc_0.Q.t40 IOUT+.t28 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X116 CM_MSB_V2_0.SD IM.t15 VSS.t94 VSS.t93 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X117 CM_MSB_V2_0.OUT Local_Enc_0.Q.t41 IOUT+.t27 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X118 CM_MSB_V2_0.OUT Local_Enc_0.Q.t42 IOUT+.t26 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X119 IOUT+ Local_Enc_0.Q.t43 CM_MSB_V2_0.OUT.t147 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X120 VSS IM.t16 CM_MSB_V2_0.SD.t50 VSS.t35 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X121 CM_MSB_V2_0.OUT Local_Enc_0.Q.t44 IOUT+.t24 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X122 CM_MSB_V2_0.OUT Local_Enc_0.Q.t45 IOUT+.t23 VSS.t46 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X123 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_6.A a_n1846_3765# VSS.t36 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X124 a_n2609_4741# Ci.t2 VSS.t32 VSS.t31 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X125 CM_MSB_V2_0.OUT IM_T.t17 CM_MSB_V2_0.SD.t15 VSS.t33 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X126 CM_MSB_V2_0.OUT Local_Enc_0.QB.t36 IOUT-.t31 VSS.t44 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X127 CM_MSB_V2_0.OUT Local_Enc_0.QB.t37 IOUT-.t30 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X128 CM_MSB_V2_0.SD IM_T.t18 CM_MSB_V2_0.OUT.t18 VSS.t34 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X129 IOUT- Local_Enc_0.QB.t38 CM_MSB_V2_0.OUT.t49 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X130 CM_MSB_V2_0.OUT IM_T.t19 CM_MSB_V2_0.SD.t13 VSS.t19 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X131 IOUT- Local_Enc_0.QB.t39 CM_MSB_V2_0.OUT.t48 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X132 IOUT+ Local_Enc_0.Q.t46 CM_MSB_V2_0.OUT.t144 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X133 CM_MSB_V2_0.OUT Local_Enc_0.Q.t47 IOUT+.t21 VSS.t44 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X134 Local_Enc_0.NAND_6.B Ci.t3 a_n2609_4741# VSS.t59 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X135 VSS IM.t17 CM_MSB_V2_0.SD.t56 VSS.t15 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X136 IOUT+ Local_Enc_0.Q.t48 CM_MSB_V2_0.OUT.t146 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X137 IOUT- Local_Enc_0.QB.t40 CM_MSB_V2_0.OUT.t47 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X138 IOUT+ Local_Enc_0.Q.t49 CM_MSB_V2_0.OUT.t118 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X139 CM_MSB_V2_0.OUT Local_Enc_0.QB.t41 IOUT-.t26 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X140 IOUT- Local_Enc_0.QB.t42 CM_MSB_V2_0.OUT.t46 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X141 IOUT- Local_Enc_0.QB.t43 CM_MSB_V2_0.OUT.t45 VSS.t40 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X142 IOUT- Local_Enc_0.QB.t44 CM_MSB_V2_0.OUT.t44 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X143 IOUT- Local_Enc_0.QB.t45 CM_MSB_V2_0.OUT.t43 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X144 CM_MSB_V2_0.SD IM.t18 VSS.t110 VSS.t62 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X145 CM_MSB_V2_0.OUT Local_Enc_0.Q.t50 IOUT+.t18 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X146 CM_MSB_V2_0.OUT Local_Enc_0.Q.t51 IOUT+.t17 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X147 CM_MSB_V2_0.OUT Local_Enc_0.Q.t52 IOUT+.t16 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X148 IOUT+ Local_Enc_0.Q.t53 CM_MSB_V2_0.OUT.t135 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X149 IOUT+ Local_Enc_0.Q.t54 CM_MSB_V2_0.OUT.t136 VSS.t40 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X150 CM_MSB_V2_0.SD IM_T.t20 CM_MSB_V2_0.OUT.t14 VSS.t20 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X151 a_n2609_3766# Ri.t2 VSS.t28 VSS.t27 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X152 a_n1846_5712# Local_Enc_0.NAND_1.B VSS.t26 VSS.t25 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X153 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_1.B VDD.t18 VDD.t17 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X154 CM_MSB_V2_0.SD IM_T.t21 CM_MSB_V2_0.OUT.t4 VSS.t10 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X155 Local_Enc_0.NAND_6.A Ri.t3 a_n2609_3766# VSS.t8 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X156 IOUT+ Local_Enc_0.Q.t55 CM_MSB_V2_0.OUT.t111 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X157 CM_MSB_V2_0.OUT IM_T.t22 CM_MSB_V2_0.SD.t10 VSS.t11 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X158 VSS IM.t19 CM_MSB_V2_0.SD.t54 VSS.t103 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X159 CM_MSB_V2_0.SD IM_T.t23 CM_MSB_V2_0.OUT.t1 VSS.t5 nfet_03v3 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X160 CM_MSB_V2_0.OUT Local_Enc_0.QB.t46 IOUT-.t21 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X161 CM_MSB_V2_0.OUT Local_Enc_0.QB.t47 IOUT-.t20 VSS.t46 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X162 CM_MSB_V2_0.OUT Local_Enc_0.QB.t48 IOUT-.t19 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X163 VSS IM.t20 CM_MSB_V2_0.SD.t55 VSS.t21 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X164 CM_MSB_V2_0.OUT IM_T.t24 CM_MSB_V2_0.SD.t8 VSS.t6 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X165 VDD Local_Enc_0.NAND_8.A Local_Enc_0.NAND_4.B VDD.t8 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X166 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_5.A a_n1846_4741# VSS.t7 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X167 CM_MSB_V2_0.SD IM.t21 VSS.t91 VSS.t14 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X168 CM_MSB_V2_0.OUT Local_Enc_0.Q.t56 IOUT+.t12 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X169 CM_MSB_V2_0.OUT Local_Enc_0.Q.t57 IOUT+.t11 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X170 CM_MSB_V2_0.OUT Local_Enc_0.QB.t49 IOUT-.t18 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X171 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_8.A VDD.t7 VDD.t6 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X172 Local_Enc_0.NAND_1.B Ri-1.t0 VDD.t25 VDD.t24 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X173 a_n2609_5712# Ri-1.t1 VSS.t61 VSS.t60 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X174 CM_MSB_V2_0.OUT Local_Enc_0.QB.t50 IOUT-.t17 VSS.t44 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X175 CM_MSB_V2_0.OUT IM_T.t25 CM_MSB_V2_0.SD.t7 VSS.t113 nfet_03v3 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
X176 IOUT+ Local_Enc_0.Q.t58 CM_MSB_V2_0.OUT.t95 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X177 CM_MSB_V2_0.OUT Local_Enc_0.QB.t51 IOUT-.t16 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X178 CM_MSB_V2_0.OUT Local_Enc_0.QB.t52 IOUT-.t15 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X179 IOUT- Local_Enc_0.QB.t53 CM_MSB_V2_0.OUT.t42 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X180 CM_MSB_V2_0.SD IM.t22 VSS.t92 VSS.t29 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X181 IOUT- Local_Enc_0.QB.t54 CM_MSB_V2_0.OUT.t41 VSS.t52 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X182 VDD Ri-1.t2 Local_Enc_0.NAND_1.B VDD.t0 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X183 Local_Enc_0.NAND_1.B Ri-1.t3 a_n2609_5712# VSS.t30 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X184 VSS IM.t23 CM_MSB_V2_0.SD.t45 VSS.t18 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X185 IOUT+ Local_Enc_0.Q.t59 CM_MSB_V2_0.OUT.t127 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X186 IOUT+ Local_Enc_0.Q.t60 CM_MSB_V2_0.OUT.t128 VSS.t53 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X187 CM_MSB_V2_0.SD IM.t24 VSS.t90 VSS.t63 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X188 IOUT+ Local_Enc_0.Q.t61 CM_MSB_V2_0.OUT.t100 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X189 CM_MSB_V2_0.OUT IM_T.t26 CM_MSB_V2_0.SD.t6 VSS.t119 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X190 IOUT+ Local_Enc_0.Q.t62 CM_MSB_V2_0.OUT.t149 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X191 IOUT+ Local_Enc_0.Q.t63 CM_MSB_V2_0.OUT.t137 VSS.t55 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X192 CM_MSB_V2_0.OUT Local_Enc_0.QB.t55 IOUT-.t12 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X193 IOUT- Local_Enc_0.QB.t56 CM_MSB_V2_0.OUT.t40 VSS.t50 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X194 IOUT- Local_Enc_0.QB.t57 CM_MSB_V2_0.OUT.t39 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X195 IOUT- Local_Enc_0.QB.t58 CM_MSB_V2_0.OUT.t38 VSS.t40 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X196 IOUT- Local_Enc_0.QB.t59 CM_MSB_V2_0.OUT.t37 VSS.t48 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X197 IOUT- Local_Enc_0.QB.t60 CM_MSB_V2_0.OUT.t36 VSS.t47 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X198 CM_MSB_V2_0.OUT Local_Enc_0.QB.t61 IOUT-.t6 VSS.t46 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X199 CM_MSB_V2_0.OUT Local_Enc_0.Q.t64 IOUT+.t4 VSS.t51 nfet_03v3 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X200 IOUT+ Local_Enc_0.Q.t65 CM_MSB_V2_0.OUT.t115 VSS.t49 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X201 CM_MSB_V2_0.SD IM_T.t27 CM_MSB_V2_0.OUT.t156 VSS.t68 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X202 CM_MSB_V2_0.OUT Local_Enc_0.QB.t62 IOUT-.t5 VSS.t45 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X203 CM_MSB_V2_0.OUT Local_Enc_0.QB.t63 IOUT-.t4 VSS.t44 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X204 CM_MSB_V2_0.SD IM.t25 VSS.t87 VSS.t16 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X205 CM_MSB_V2_0.OUT Local_Enc_0.QB.t64 IOUT-.t3 VSS.t43 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X206 CM_MSB_V2_0.OUT Local_Enc_0.Q.t66 IOUT+.t2 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X207 CM_MSB_V2_0.OUT IM_T.t28 CM_MSB_V2_0.SD.t4 VSS.t97 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X208 CM_MSB_V2_0.SD IM.t26 VSS.t77 VSS.t17 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X209 CM_MSB_V2_0.SD IM_T.t29 CM_MSB_V2_0.OUT.t158 VSS.t93 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X210 CM_MSB_V2_0.OUT Local_Enc_0.QB.t65 IOUT-.t2 VSS.t42 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X211 CM_MSB_V2_0.OUT Local_Enc_0.QB.t66 IOUT-.t1 VSS.t41 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X212 VSS IM.t27 CM_MSB_V2_0.SD.t39 VSS.t33 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X213 IOUT- Local_Enc_0.QB.t67 CM_MSB_V2_0.OUT.t35 VSS.t40 nfet_03v3 ad=0.264p pd=2.08u as=0.156p ps=1.12u w=0.6u l=0.5u
X214 VDD Local_Enc_0.NAND_8.A Local_Enc_0.Q.t1 VDD.t3 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X215 CM_MSB_V2_0.OUT Local_Enc_0.Q.t67 IOUT+.t1 VSS.t54 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X216 VSS IM.t28 CM_MSB_V2_0.SD.t42 VSS.t19 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X217 CM_MSB_V2_0.SD IM.t29 VSS.t85 VSS.t34 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X218 CM_MSB_V2_0.OUT Local_Enc_0.Q.t68 IOUT+.t0 VSS.t46 nfet_03v3 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X219 CM_MSB_V2_0.OUT IM_T.t30 CM_MSB_V2_0.SD.t2 VSS.t116 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X220 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_1.B a_n1846_5712# VSS.t24 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X221 Local_Enc_0.Q Local_Enc_0.QB.t68 VDD.t32 VDD.t31 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X222 CM_MSB_V2_0.OUT IM_T.t31 CM_MSB_V2_0.SD.t1 VSS.t15 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X223 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_8.A a_n1035_3765# VSS.t2 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X224 VDD Local_Enc_0.NAND_1.B Local_Enc_0.NAND_5.B VDD.t14 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X225 VSS IM.t30 CM_MSB_V2_0.SD.t36 VSS.t73 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X226 CM_MSB_V2_0.SD IM.t31 VSS.t76 VSS.t12 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X227 a_n1035_3765# Local_Enc_0.NAND_8.A VSS.t1 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 Local_Enc_0.QB.n1 Local_Enc_0.QB.t14 26.9784
R1 Local_Enc_0.QB.n17 Local_Enc_0.QB.t29 24.9712
R2 Local_Enc_0.QB.n32 Local_Enc_0.QB.t58 24.9712
R3 Local_Enc_0.QB.n47 Local_Enc_0.QB.t43 24.9712
R4 Local_Enc_0.QB.n2 Local_Enc_0.QB.t67 24.9712
R5 Local_Enc_0.QB.n62 Local_Enc_0.QB.n61 21.4076
R6 Local_Enc_0.QB.n0 Local_Enc_0.QB.n16 21.1997
R7 Local_Enc_0.QB.n0 Local_Enc_0.QB.n31 20.1581
R8 Local_Enc_0.QB.n62 Local_Enc_0.QB.n46 20.1567
R9 Local_Enc_0.QB.n19 Local_Enc_0.QB.t23 15.1115
R10 Local_Enc_0.QB.n20 Local_Enc_0.QB.t57 15.1115
R11 Local_Enc_0.QB.n23 Local_Enc_0.QB.t34 15.1115
R12 Local_Enc_0.QB.n24 Local_Enc_0.QB.t4 15.1115
R13 Local_Enc_0.QB.n27 Local_Enc_0.QB.t20 15.1115
R14 Local_Enc_0.QB.n28 Local_Enc_0.QB.t38 15.1115
R15 Local_Enc_0.QB.n34 Local_Enc_0.QB.t50 15.1115
R16 Local_Enc_0.QB.n35 Local_Enc_0.QB.t19 15.1115
R17 Local_Enc_0.QB.n38 Local_Enc_0.QB.t66 15.1115
R18 Local_Enc_0.QB.n39 Local_Enc_0.QB.t31 15.1115
R19 Local_Enc_0.QB.n42 Local_Enc_0.QB.t47 15.1115
R20 Local_Enc_0.QB.n43 Local_Enc_0.QB.t3 15.1115
R21 Local_Enc_0.QB.n49 Local_Enc_0.QB.t36 15.1115
R22 Local_Enc_0.QB.n50 Local_Enc_0.QB.t6 15.1115
R23 Local_Enc_0.QB.n53 Local_Enc_0.QB.t48 15.1115
R24 Local_Enc_0.QB.n54 Local_Enc_0.QB.t16 15.1115
R25 Local_Enc_0.QB.n57 Local_Enc_0.QB.t35 15.1115
R26 Local_Enc_0.QB.n58 Local_Enc_0.QB.t53 15.1115
R27 Local_Enc_0.QB.n4 Local_Enc_0.QB.t63 15.1115
R28 Local_Enc_0.QB.n5 Local_Enc_0.QB.t28 15.1115
R29 Local_Enc_0.QB.n8 Local_Enc_0.QB.t9 15.1115
R30 Local_Enc_0.QB.n9 Local_Enc_0.QB.t39 15.1115
R31 Local_Enc_0.QB.n12 Local_Enc_0.QB.t61 15.1115
R32 Local_Enc_0.QB.n13 Local_Enc_0.QB.t12 15.1115
R33 Local_Enc_0.QB.n1 Local_Enc_0.QB.t68 14.7248
R34 Local_Enc_0.QB.n17 Local_Enc_0.QB.t46 14.4545
R35 Local_Enc_0.QB.n18 Local_Enc_0.QB.t45 14.4545
R36 Local_Enc_0.QB.n21 Local_Enc_0.QB.t64 14.4545
R37 Local_Enc_0.QB.n22 Local_Enc_0.QB.t30 14.4545
R38 Local_Enc_0.QB.n25 Local_Enc_0.QB.t24 14.4545
R39 Local_Enc_0.QB.n26 Local_Enc_0.QB.t40 14.4545
R40 Local_Enc_0.QB.n29 Local_Enc_0.QB.t62 14.4545
R41 Local_Enc_0.QB.n30 Local_Enc_0.QB.t27 14.4545
R42 Local_Enc_0.QB.n32 Local_Enc_0.QB.t13 14.4545
R43 Local_Enc_0.QB.n33 Local_Enc_0.QB.t8 14.4545
R44 Local_Enc_0.QB.n36 Local_Enc_0.QB.t25 14.4545
R45 Local_Enc_0.QB.n37 Local_Enc_0.QB.t60 14.4545
R46 Local_Enc_0.QB.n40 Local_Enc_0.QB.t51 14.4545
R47 Local_Enc_0.QB.n41 Local_Enc_0.QB.t5 14.4545
R48 Local_Enc_0.QB.n44 Local_Enc_0.QB.t22 14.4545
R49 Local_Enc_0.QB.n45 Local_Enc_0.QB.t56 14.4545
R50 Local_Enc_0.QB.n47 Local_Enc_0.QB.t41 14.4545
R51 Local_Enc_0.QB.n48 Local_Enc_0.QB.t33 14.4545
R52 Local_Enc_0.QB.n51 Local_Enc_0.QB.t52 14.4545
R53 Local_Enc_0.QB.n52 Local_Enc_0.QB.t21 14.4545
R54 Local_Enc_0.QB.n55 Local_Enc_0.QB.t15 14.4545
R55 Local_Enc_0.QB.n56 Local_Enc_0.QB.t32 14.4545
R56 Local_Enc_0.QB.n59 Local_Enc_0.QB.t49 14.4545
R57 Local_Enc_0.QB.n60 Local_Enc_0.QB.t18 14.4545
R58 Local_Enc_0.QB.n2 Local_Enc_0.QB.t65 14.4545
R59 Local_Enc_0.QB.n3 Local_Enc_0.QB.t59 14.4545
R60 Local_Enc_0.QB.n6 Local_Enc_0.QB.t11 14.4545
R61 Local_Enc_0.QB.n7 Local_Enc_0.QB.t44 14.4545
R62 Local_Enc_0.QB.n10 Local_Enc_0.QB.t37 14.4545
R63 Local_Enc_0.QB.n11 Local_Enc_0.QB.t54 14.4545
R64 Local_Enc_0.QB.n14 Local_Enc_0.QB.t10 14.4545
R65 Local_Enc_0.QB.n15 Local_Enc_0.QB.t42 14.4545
R66 Local_Enc_0.QB.n31 Local_Enc_0.QB.n30 12.7802
R67 Local_Enc_0.QB.n46 Local_Enc_0.QB.n45 12.7802
R68 Local_Enc_0.QB.n61 Local_Enc_0.QB.n60 12.7802
R69 Local_Enc_0.QB.n16 Local_Enc_0.QB.n15 12.7802
R70 Local_Enc_0.QB.n31 Local_Enc_0.QB.t55 12.1915
R71 Local_Enc_0.QB.n46 Local_Enc_0.QB.t17 12.1915
R72 Local_Enc_0.QB.n61 Local_Enc_0.QB.t7 12.1915
R73 Local_Enc_0.QB.n16 Local_Enc_0.QB.t26 12.1915
R74 Local_Enc_0.QB.n18 Local_Enc_0.QB.n17 9.86024
R75 Local_Enc_0.QB.n19 Local_Enc_0.QB.n18 9.86024
R76 Local_Enc_0.QB.n20 Local_Enc_0.QB.n19 9.86024
R77 Local_Enc_0.QB.n21 Local_Enc_0.QB.n20 9.86024
R78 Local_Enc_0.QB.n22 Local_Enc_0.QB.n21 9.86024
R79 Local_Enc_0.QB.n23 Local_Enc_0.QB.n22 9.86024
R80 Local_Enc_0.QB.n24 Local_Enc_0.QB.n23 9.86024
R81 Local_Enc_0.QB.n25 Local_Enc_0.QB.n24 9.86024
R82 Local_Enc_0.QB.n26 Local_Enc_0.QB.n25 9.86024
R83 Local_Enc_0.QB.n27 Local_Enc_0.QB.n26 9.86024
R84 Local_Enc_0.QB.n28 Local_Enc_0.QB.n27 9.86024
R85 Local_Enc_0.QB.n29 Local_Enc_0.QB.n28 9.86024
R86 Local_Enc_0.QB.n30 Local_Enc_0.QB.n29 9.86024
R87 Local_Enc_0.QB.n33 Local_Enc_0.QB.n32 9.86024
R88 Local_Enc_0.QB.n34 Local_Enc_0.QB.n33 9.86024
R89 Local_Enc_0.QB.n35 Local_Enc_0.QB.n34 9.86024
R90 Local_Enc_0.QB.n36 Local_Enc_0.QB.n35 9.86024
R91 Local_Enc_0.QB.n37 Local_Enc_0.QB.n36 9.86024
R92 Local_Enc_0.QB.n38 Local_Enc_0.QB.n37 9.86024
R93 Local_Enc_0.QB.n39 Local_Enc_0.QB.n38 9.86024
R94 Local_Enc_0.QB.n40 Local_Enc_0.QB.n39 9.86024
R95 Local_Enc_0.QB.n41 Local_Enc_0.QB.n40 9.86024
R96 Local_Enc_0.QB.n42 Local_Enc_0.QB.n41 9.86024
R97 Local_Enc_0.QB.n43 Local_Enc_0.QB.n42 9.86024
R98 Local_Enc_0.QB.n44 Local_Enc_0.QB.n43 9.86024
R99 Local_Enc_0.QB.n45 Local_Enc_0.QB.n44 9.86024
R100 Local_Enc_0.QB.n48 Local_Enc_0.QB.n47 9.86024
R101 Local_Enc_0.QB.n49 Local_Enc_0.QB.n48 9.86024
R102 Local_Enc_0.QB.n50 Local_Enc_0.QB.n49 9.86024
R103 Local_Enc_0.QB.n51 Local_Enc_0.QB.n50 9.86024
R104 Local_Enc_0.QB.n52 Local_Enc_0.QB.n51 9.86024
R105 Local_Enc_0.QB.n53 Local_Enc_0.QB.n52 9.86024
R106 Local_Enc_0.QB.n54 Local_Enc_0.QB.n53 9.86024
R107 Local_Enc_0.QB.n55 Local_Enc_0.QB.n54 9.86024
R108 Local_Enc_0.QB.n56 Local_Enc_0.QB.n55 9.86024
R109 Local_Enc_0.QB.n57 Local_Enc_0.QB.n56 9.86024
R110 Local_Enc_0.QB.n58 Local_Enc_0.QB.n57 9.86024
R111 Local_Enc_0.QB.n59 Local_Enc_0.QB.n58 9.86024
R112 Local_Enc_0.QB.n60 Local_Enc_0.QB.n59 9.86024
R113 Local_Enc_0.QB.n3 Local_Enc_0.QB.n2 9.86024
R114 Local_Enc_0.QB.n4 Local_Enc_0.QB.n3 9.86024
R115 Local_Enc_0.QB.n5 Local_Enc_0.QB.n4 9.86024
R116 Local_Enc_0.QB.n6 Local_Enc_0.QB.n5 9.86024
R117 Local_Enc_0.QB.n7 Local_Enc_0.QB.n6 9.86024
R118 Local_Enc_0.QB.n8 Local_Enc_0.QB.n7 9.86024
R119 Local_Enc_0.QB.n9 Local_Enc_0.QB.n8 9.86024
R120 Local_Enc_0.QB.n10 Local_Enc_0.QB.n9 9.86024
R121 Local_Enc_0.QB.n11 Local_Enc_0.QB.n10 9.86024
R122 Local_Enc_0.QB.n12 Local_Enc_0.QB.n11 9.86024
R123 Local_Enc_0.QB.n13 Local_Enc_0.QB.n12 9.86024
R124 Local_Enc_0.QB.n14 Local_Enc_0.QB.n13 9.86024
R125 Local_Enc_0.QB.n15 Local_Enc_0.QB.n14 9.86024
R126 Local_Enc_0.QB.n63 Local_Enc_0.QB 8.0222
R127 Local_Enc_0.QB Local_Enc_0.QB.n1 4.18544
R128 Local_Enc_0.QB.t1 Local_Enc_0.QB.n64 3.6405
R129 Local_Enc_0.QB Local_Enc_0.QB.t1 3.08447
R130 Local_Enc_0.QB Local_Enc_0.QB.n63 2.66528
R131 Local_Enc_0.QB.n0 Local_Enc_0.QB.n62 1.23881
R132 Local_Enc_0.QB.n63 Local_Enc_0.QB.n0 1.033
R133 CM_MSB_V2_0.OUT.n228 CM_MSB_V2_0.OUT.t1 5.37963
R134 CM_MSB_V2_0.OUT CM_MSB_V2_0.OUT.n196 4.89917
R135 CM_MSB_V2_0.OUT.n243 CM_MSB_V2_0.OUT.n197 4.86963
R136 CM_MSB_V2_0.OUT.n46 CM_MSB_V2_0.OUT.n45 3.9342
R137 CM_MSB_V2_0.OUT.n38 CM_MSB_V2_0.OUT.n37 3.9339
R138 CM_MSB_V2_0.OUT.n133 CM_MSB_V2_0.OUT.n132 3.78102
R139 CM_MSB_V2_0.OUT.n228 CM_MSB_V2_0.OUT.n227 3.61615
R140 CM_MSB_V2_0.OUT.n230 CM_MSB_V2_0.OUT.n223 3.61615
R141 CM_MSB_V2_0.OUT.n232 CM_MSB_V2_0.OUT.n219 3.61615
R142 CM_MSB_V2_0.OUT.n234 CM_MSB_V2_0.OUT.n215 3.61615
R143 CM_MSB_V2_0.OUT.n236 CM_MSB_V2_0.OUT.n211 3.61615
R144 CM_MSB_V2_0.OUT.n238 CM_MSB_V2_0.OUT.n207 3.61615
R145 CM_MSB_V2_0.OUT.n240 CM_MSB_V2_0.OUT.n203 3.61615
R146 CM_MSB_V2_0.OUT.n242 CM_MSB_V2_0.OUT.n199 3.61615
R147 CM_MSB_V2_0.OUT.n32 CM_MSB_V2_0.OUT.n31 3.50723
R148 CM_MSB_V2_0.OUT.n12 CM_MSB_V2_0.OUT.n11 3.50723
R149 CM_MSB_V2_0.OUT.n22 CM_MSB_V2_0.OUT.n21 3.50723
R150 CM_MSB_V2_0.OUT.n33 CM_MSB_V2_0.OUT.n27 3.50518
R151 CM_MSB_V2_0.OUT.n13 CM_MSB_V2_0.OUT.n7 3.50518
R152 CM_MSB_V2_0.OUT.n23 CM_MSB_V2_0.OUT.n17 3.50518
R153 CM_MSB_V2_0.OUT.n46 CM_MSB_V2_0.OUT.n43 3.50518
R154 CM_MSB_V2_0.OUT.n241 CM_MSB_V2_0.OUT.n201 3.50463
R155 CM_MSB_V2_0.OUT.n239 CM_MSB_V2_0.OUT.n205 3.50463
R156 CM_MSB_V2_0.OUT.n237 CM_MSB_V2_0.OUT.n209 3.50463
R157 CM_MSB_V2_0.OUT.n235 CM_MSB_V2_0.OUT.n213 3.50463
R158 CM_MSB_V2_0.OUT.n233 CM_MSB_V2_0.OUT.n217 3.50463
R159 CM_MSB_V2_0.OUT.n231 CM_MSB_V2_0.OUT.n221 3.50463
R160 CM_MSB_V2_0.OUT.n229 CM_MSB_V2_0.OUT.n225 3.50463
R161 CM_MSB_V2_0.OUT.n183 CM_MSB_V2_0.OUT.n175 3.5031
R162 CM_MSB_V2_0.OUT.n143 CM_MSB_V2_0.OUT.n137 3.5031
R163 CM_MSB_V2_0.OUT.n142 CM_MSB_V2_0.OUT.n141 3.5031
R164 CM_MSB_V2_0.OUT.n153 CM_MSB_V2_0.OUT.n147 3.5031
R165 CM_MSB_V2_0.OUT.n152 CM_MSB_V2_0.OUT.n151 3.5031
R166 CM_MSB_V2_0.OUT.n38 CM_MSB_V2_0.OUT.n35 3.5031
R167 CM_MSB_V2_0.OUT.n180 CM_MSB_V2_0.OUT.n179 3.5031
R168 CM_MSB_V2_0.OUT.n143 CM_MSB_V2_0.OUT.n135 3.41897
R169 CM_MSB_V2_0.OUT.n142 CM_MSB_V2_0.OUT.n139 3.41897
R170 CM_MSB_V2_0.OUT.n153 CM_MSB_V2_0.OUT.n145 3.41897
R171 CM_MSB_V2_0.OUT.n152 CM_MSB_V2_0.OUT.n149 3.41897
R172 CM_MSB_V2_0.OUT.n32 CM_MSB_V2_0.OUT.n29 3.41897
R173 CM_MSB_V2_0.OUT.n33 CM_MSB_V2_0.OUT.n25 3.41897
R174 CM_MSB_V2_0.OUT.n12 CM_MSB_V2_0.OUT.n9 3.41897
R175 CM_MSB_V2_0.OUT.n13 CM_MSB_V2_0.OUT.n5 3.41897
R176 CM_MSB_V2_0.OUT.n22 CM_MSB_V2_0.OUT.n19 3.41897
R177 CM_MSB_V2_0.OUT.n23 CM_MSB_V2_0.OUT.n15 3.41897
R178 CM_MSB_V2_0.OUT.n180 CM_MSB_V2_0.OUT.n177 3.41897
R179 CM_MSB_V2_0.OUT.n183 CM_MSB_V2_0.OUT.n182 3.41897
R180 CM_MSB_V2_0.OUT.n196 CM_MSB_V2_0.OUT.n1 3.37397
R181 CM_MSB_V2_0.OUT.n195 CM_MSB_V2_0.OUT.n3 3.37397
R182 CM_MSB_V2_0.OUT.n133 CM_MSB_V2_0.OUT.n130 3.37397
R183 CM_MSB_V2_0.OUT.n50 CM_MSB_V2_0.OUT.n49 3.1505
R184 CM_MSB_V2_0.OUT.n53 CM_MSB_V2_0.OUT.n52 3.1505
R185 CM_MSB_V2_0.OUT.n57 CM_MSB_V2_0.OUT.n56 3.1505
R186 CM_MSB_V2_0.OUT.n60 CM_MSB_V2_0.OUT.n59 3.1505
R187 CM_MSB_V2_0.OUT.n64 CM_MSB_V2_0.OUT.n63 3.1505
R188 CM_MSB_V2_0.OUT.n67 CM_MSB_V2_0.OUT.n66 3.1505
R189 CM_MSB_V2_0.OUT.n71 CM_MSB_V2_0.OUT.n70 3.1505
R190 CM_MSB_V2_0.OUT.n74 CM_MSB_V2_0.OUT.n73 3.1505
R191 CM_MSB_V2_0.OUT.n80 CM_MSB_V2_0.OUT.n79 3.1505
R192 CM_MSB_V2_0.OUT.n77 CM_MSB_V2_0.OUT.n76 3.1505
R193 CM_MSB_V2_0.OUT.n87 CM_MSB_V2_0.OUT.n86 3.1505
R194 CM_MSB_V2_0.OUT.n84 CM_MSB_V2_0.OUT.n83 3.1505
R195 CM_MSB_V2_0.OUT.n94 CM_MSB_V2_0.OUT.n93 3.1505
R196 CM_MSB_V2_0.OUT.n91 CM_MSB_V2_0.OUT.n90 3.1505
R197 CM_MSB_V2_0.OUT.n101 CM_MSB_V2_0.OUT.n100 3.1505
R198 CM_MSB_V2_0.OUT.n98 CM_MSB_V2_0.OUT.n97 3.1505
R199 CM_MSB_V2_0.OUT.n107 CM_MSB_V2_0.OUT.n106 3.1505
R200 CM_MSB_V2_0.OUT.n104 CM_MSB_V2_0.OUT.n103 3.1505
R201 CM_MSB_V2_0.OUT.n114 CM_MSB_V2_0.OUT.n113 3.1505
R202 CM_MSB_V2_0.OUT.n111 CM_MSB_V2_0.OUT.n110 3.1505
R203 CM_MSB_V2_0.OUT.n121 CM_MSB_V2_0.OUT.n120 3.1505
R204 CM_MSB_V2_0.OUT.n118 CM_MSB_V2_0.OUT.n117 3.1505
R205 CM_MSB_V2_0.OUT.n128 CM_MSB_V2_0.OUT.n127 3.1505
R206 CM_MSB_V2_0.OUT.n125 CM_MSB_V2_0.OUT.n124 3.1505
R207 CM_MSB_V2_0.OUT.n159 CM_MSB_V2_0.OUT.n158 3.1505
R208 CM_MSB_V2_0.OUT.n156 CM_MSB_V2_0.OUT.n155 3.1505
R209 CM_MSB_V2_0.OUT.n166 CM_MSB_V2_0.OUT.n165 3.1505
R210 CM_MSB_V2_0.OUT.n163 CM_MSB_V2_0.OUT.n162 3.1505
R211 CM_MSB_V2_0.OUT.n173 CM_MSB_V2_0.OUT.n172 3.1505
R212 CM_MSB_V2_0.OUT.n170 CM_MSB_V2_0.OUT.n169 3.1505
R213 CM_MSB_V2_0.OUT.n190 CM_MSB_V2_0.OUT.n189 3.1505
R214 CM_MSB_V2_0.OUT.n187 CM_MSB_V2_0.OUT.n186 3.1505
R215 CM_MSB_V2_0.OUT.n175 CM_MSB_V2_0.OUT.t132 2.7305
R216 CM_MSB_V2_0.OUT.n175 CM_MSB_V2_0.OUT.n174 2.7305
R217 CM_MSB_V2_0.OUT.n186 CM_MSB_V2_0.OUT.t51 2.7305
R218 CM_MSB_V2_0.OUT.n186 CM_MSB_V2_0.OUT.n185 2.7305
R219 CM_MSB_V2_0.OUT.n189 CM_MSB_V2_0.OUT.t150 2.7305
R220 CM_MSB_V2_0.OUT.n189 CM_MSB_V2_0.OUT.n188 2.7305
R221 CM_MSB_V2_0.OUT.n169 CM_MSB_V2_0.OUT.t64 2.7305
R222 CM_MSB_V2_0.OUT.n169 CM_MSB_V2_0.OUT.n168 2.7305
R223 CM_MSB_V2_0.OUT.n172 CM_MSB_V2_0.OUT.t117 2.7305
R224 CM_MSB_V2_0.OUT.n172 CM_MSB_V2_0.OUT.n171 2.7305
R225 CM_MSB_V2_0.OUT.n162 CM_MSB_V2_0.OUT.t47 2.7305
R226 CM_MSB_V2_0.OUT.n162 CM_MSB_V2_0.OUT.n161 2.7305
R227 CM_MSB_V2_0.OUT.n165 CM_MSB_V2_0.OUT.t95 2.7305
R228 CM_MSB_V2_0.OUT.n165 CM_MSB_V2_0.OUT.n164 2.7305
R229 CM_MSB_V2_0.OUT.n155 CM_MSB_V2_0.OUT.t41 2.7305
R230 CM_MSB_V2_0.OUT.n155 CM_MSB_V2_0.OUT.n154 2.7305
R231 CM_MSB_V2_0.OUT.n158 CM_MSB_V2_0.OUT.t140 2.7305
R232 CM_MSB_V2_0.OUT.n158 CM_MSB_V2_0.OUT.n157 2.7305
R233 CM_MSB_V2_0.OUT.n137 CM_MSB_V2_0.OUT.t128 2.7305
R234 CM_MSB_V2_0.OUT.n137 CM_MSB_V2_0.OUT.n136 2.7305
R235 CM_MSB_V2_0.OUT.n135 CM_MSB_V2_0.OUT.t49 2.7305
R236 CM_MSB_V2_0.OUT.n135 CM_MSB_V2_0.OUT.n134 2.7305
R237 CM_MSB_V2_0.OUT.n141 CM_MSB_V2_0.OUT.t40 2.7305
R238 CM_MSB_V2_0.OUT.n141 CM_MSB_V2_0.OUT.n140 2.7305
R239 CM_MSB_V2_0.OUT.n139 CM_MSB_V2_0.OUT.t144 2.7305
R240 CM_MSB_V2_0.OUT.n139 CM_MSB_V2_0.OUT.n138 2.7305
R241 CM_MSB_V2_0.OUT.n147 CM_MSB_V2_0.OUT.t96 2.7305
R242 CM_MSB_V2_0.OUT.n147 CM_MSB_V2_0.OUT.n146 2.7305
R243 CM_MSB_V2_0.OUT.n145 CM_MSB_V2_0.OUT.t61 2.7305
R244 CM_MSB_V2_0.OUT.n145 CM_MSB_V2_0.OUT.n144 2.7305
R245 CM_MSB_V2_0.OUT.n151 CM_MSB_V2_0.OUT.t56 2.7305
R246 CM_MSB_V2_0.OUT.n151 CM_MSB_V2_0.OUT.n150 2.7305
R247 CM_MSB_V2_0.OUT.n149 CM_MSB_V2_0.OUT.t88 2.7305
R248 CM_MSB_V2_0.OUT.n149 CM_MSB_V2_0.OUT.n148 2.7305
R249 CM_MSB_V2_0.OUT.n37 CM_MSB_V2_0.OUT.t46 2.7305
R250 CM_MSB_V2_0.OUT.n37 CM_MSB_V2_0.OUT.n36 2.7305
R251 CM_MSB_V2_0.OUT.n35 CM_MSB_V2_0.OUT.t146 2.7305
R252 CM_MSB_V2_0.OUT.n35 CM_MSB_V2_0.OUT.n34 2.7305
R253 CM_MSB_V2_0.OUT.n1 CM_MSB_V2_0.OUT.t45 2.7305
R254 CM_MSB_V2_0.OUT.n1 CM_MSB_V2_0.OUT.n0 2.7305
R255 CM_MSB_V2_0.OUT.n3 CM_MSB_V2_0.OUT.t87 2.7305
R256 CM_MSB_V2_0.OUT.n3 CM_MSB_V2_0.OUT.n2 2.7305
R257 CM_MSB_V2_0.OUT.n124 CM_MSB_V2_0.OUT.t111 2.7305
R258 CM_MSB_V2_0.OUT.n124 CM_MSB_V2_0.OUT.n123 2.7305
R259 CM_MSB_V2_0.OUT.n127 CM_MSB_V2_0.OUT.t60 2.7305
R260 CM_MSB_V2_0.OUT.n127 CM_MSB_V2_0.OUT.n126 2.7305
R261 CM_MSB_V2_0.OUT.n117 CM_MSB_V2_0.OUT.t104 2.7305
R262 CM_MSB_V2_0.OUT.n117 CM_MSB_V2_0.OUT.n116 2.7305
R263 CM_MSB_V2_0.OUT.n120 CM_MSB_V2_0.OUT.t52 2.7305
R264 CM_MSB_V2_0.OUT.n120 CM_MSB_V2_0.OUT.n119 2.7305
R265 CM_MSB_V2_0.OUT.n110 CM_MSB_V2_0.OUT.t137 2.7305
R266 CM_MSB_V2_0.OUT.n110 CM_MSB_V2_0.OUT.n109 2.7305
R267 CM_MSB_V2_0.OUT.n113 CM_MSB_V2_0.OUT.t65 2.7305
R268 CM_MSB_V2_0.OUT.n113 CM_MSB_V2_0.OUT.n112 2.7305
R269 CM_MSB_V2_0.OUT.n103 CM_MSB_V2_0.OUT.t86 2.7305
R270 CM_MSB_V2_0.OUT.n103 CM_MSB_V2_0.OUT.n102 2.7305
R271 CM_MSB_V2_0.OUT.n106 CM_MSB_V2_0.OUT.t48 2.7305
R272 CM_MSB_V2_0.OUT.n106 CM_MSB_V2_0.OUT.n105 2.7305
R273 CM_MSB_V2_0.OUT.n97 CM_MSB_V2_0.OUT.t57 2.7305
R274 CM_MSB_V2_0.OUT.n97 CM_MSB_V2_0.OUT.n96 2.7305
R275 CM_MSB_V2_0.OUT.n100 CM_MSB_V2_0.OUT.t149 2.7305
R276 CM_MSB_V2_0.OUT.n100 CM_MSB_V2_0.OUT.n99 2.7305
R277 CM_MSB_V2_0.OUT.n90 CM_MSB_V2_0.OUT.t36 2.7305
R278 CM_MSB_V2_0.OUT.n90 CM_MSB_V2_0.OUT.n89 2.7305
R279 CM_MSB_V2_0.OUT.n93 CM_MSB_V2_0.OUT.t123 2.7305
R280 CM_MSB_V2_0.OUT.n93 CM_MSB_V2_0.OUT.n92 2.7305
R281 CM_MSB_V2_0.OUT.n83 CM_MSB_V2_0.OUT.t53 2.7305
R282 CM_MSB_V2_0.OUT.n83 CM_MSB_V2_0.OUT.n82 2.7305
R283 CM_MSB_V2_0.OUT.n86 CM_MSB_V2_0.OUT.t118 2.7305
R284 CM_MSB_V2_0.OUT.n86 CM_MSB_V2_0.OUT.n85 2.7305
R285 CM_MSB_V2_0.OUT.n76 CM_MSB_V2_0.OUT.t44 2.7305
R286 CM_MSB_V2_0.OUT.n76 CM_MSB_V2_0.OUT.n75 2.7305
R287 CM_MSB_V2_0.OUT.n79 CM_MSB_V2_0.OUT.t120 2.7305
R288 CM_MSB_V2_0.OUT.n79 CM_MSB_V2_0.OUT.n78 2.7305
R289 CM_MSB_V2_0.OUT.n31 CM_MSB_V2_0.OUT.t116 2.7305
R290 CM_MSB_V2_0.OUT.n31 CM_MSB_V2_0.OUT.n30 2.7305
R291 CM_MSB_V2_0.OUT.n29 CM_MSB_V2_0.OUT.t35 2.7305
R292 CM_MSB_V2_0.OUT.n29 CM_MSB_V2_0.OUT.n28 2.7305
R293 CM_MSB_V2_0.OUT.n27 CM_MSB_V2_0.OUT.t43 2.7305
R294 CM_MSB_V2_0.OUT.n27 CM_MSB_V2_0.OUT.n26 2.7305
R295 CM_MSB_V2_0.OUT.n25 CM_MSB_V2_0.OUT.t97 2.7305
R296 CM_MSB_V2_0.OUT.n25 CM_MSB_V2_0.OUT.n24 2.7305
R297 CM_MSB_V2_0.OUT.n73 CM_MSB_V2_0.OUT.t63 2.7305
R298 CM_MSB_V2_0.OUT.n73 CM_MSB_V2_0.OUT.n72 2.7305
R299 CM_MSB_V2_0.OUT.n70 CM_MSB_V2_0.OUT.t147 2.7305
R300 CM_MSB_V2_0.OUT.n70 CM_MSB_V2_0.OUT.n69 2.7305
R301 CM_MSB_V2_0.OUT.n66 CM_MSB_V2_0.OUT.t58 2.7305
R302 CM_MSB_V2_0.OUT.n66 CM_MSB_V2_0.OUT.n65 2.7305
R303 CM_MSB_V2_0.OUT.n63 CM_MSB_V2_0.OUT.t129 2.7305
R304 CM_MSB_V2_0.OUT.n63 CM_MSB_V2_0.OUT.n62 2.7305
R305 CM_MSB_V2_0.OUT.n59 CM_MSB_V2_0.OUT.t39 2.7305
R306 CM_MSB_V2_0.OUT.n59 CM_MSB_V2_0.OUT.n58 2.7305
R307 CM_MSB_V2_0.OUT.n56 CM_MSB_V2_0.OUT.t135 2.7305
R308 CM_MSB_V2_0.OUT.n56 CM_MSB_V2_0.OUT.n55 2.7305
R309 CM_MSB_V2_0.OUT.n52 CM_MSB_V2_0.OUT.t55 2.7305
R310 CM_MSB_V2_0.OUT.n52 CM_MSB_V2_0.OUT.n51 2.7305
R311 CM_MSB_V2_0.OUT.n49 CM_MSB_V2_0.OUT.t115 2.7305
R312 CM_MSB_V2_0.OUT.n49 CM_MSB_V2_0.OUT.n48 2.7305
R313 CM_MSB_V2_0.OUT.n11 CM_MSB_V2_0.OUT.t130 2.7305
R314 CM_MSB_V2_0.OUT.n11 CM_MSB_V2_0.OUT.n10 2.7305
R315 CM_MSB_V2_0.OUT.n9 CM_MSB_V2_0.OUT.t38 2.7305
R316 CM_MSB_V2_0.OUT.n9 CM_MSB_V2_0.OUT.n8 2.7305
R317 CM_MSB_V2_0.OUT.n7 CM_MSB_V2_0.OUT.t50 2.7305
R318 CM_MSB_V2_0.OUT.n7 CM_MSB_V2_0.OUT.n6 2.7305
R319 CM_MSB_V2_0.OUT.n5 CM_MSB_V2_0.OUT.t133 2.7305
R320 CM_MSB_V2_0.OUT.n5 CM_MSB_V2_0.OUT.n4 2.7305
R321 CM_MSB_V2_0.OUT.n21 CM_MSB_V2_0.OUT.t136 2.7305
R322 CM_MSB_V2_0.OUT.n21 CM_MSB_V2_0.OUT.n20 2.7305
R323 CM_MSB_V2_0.OUT.n19 CM_MSB_V2_0.OUT.t54 2.7305
R324 CM_MSB_V2_0.OUT.n19 CM_MSB_V2_0.OUT.n18 2.7305
R325 CM_MSB_V2_0.OUT.n17 CM_MSB_V2_0.OUT.t62 2.7305
R326 CM_MSB_V2_0.OUT.n17 CM_MSB_V2_0.OUT.n16 2.7305
R327 CM_MSB_V2_0.OUT.n15 CM_MSB_V2_0.OUT.t100 2.7305
R328 CM_MSB_V2_0.OUT.n15 CM_MSB_V2_0.OUT.n14 2.7305
R329 CM_MSB_V2_0.OUT.n43 CM_MSB_V2_0.OUT.t37 2.7305
R330 CM_MSB_V2_0.OUT.n43 CM_MSB_V2_0.OUT.n42 2.7305
R331 CM_MSB_V2_0.OUT.n45 CM_MSB_V2_0.OUT.t131 2.7305
R332 CM_MSB_V2_0.OUT.n45 CM_MSB_V2_0.OUT.n44 2.7305
R333 CM_MSB_V2_0.OUT.n130 CM_MSB_V2_0.OUT.t42 2.7305
R334 CM_MSB_V2_0.OUT.n130 CM_MSB_V2_0.OUT.n129 2.7305
R335 CM_MSB_V2_0.OUT.n132 CM_MSB_V2_0.OUT.t127 2.7305
R336 CM_MSB_V2_0.OUT.n132 CM_MSB_V2_0.OUT.n131 2.7305
R337 CM_MSB_V2_0.OUT.n179 CM_MSB_V2_0.OUT.t59 2.7305
R338 CM_MSB_V2_0.OUT.n179 CM_MSB_V2_0.OUT.n178 2.7305
R339 CM_MSB_V2_0.OUT.n177 CM_MSB_V2_0.OUT.t151 2.7305
R340 CM_MSB_V2_0.OUT.n177 CM_MSB_V2_0.OUT.n176 2.7305
R341 CM_MSB_V2_0.OUT.n182 CM_MSB_V2_0.OUT.t66 2.7305
R342 CM_MSB_V2_0.OUT.n182 CM_MSB_V2_0.OUT.n181 2.7305
R343 CM_MSB_V2_0.OUT.n201 CM_MSB_V2_0.OUT.t4 1.3655
R344 CM_MSB_V2_0.OUT.n201 CM_MSB_V2_0.OUT.n200 1.3655
R345 CM_MSB_V2_0.OUT.n205 CM_MSB_V2_0.OUT.t103 1.3655
R346 CM_MSB_V2_0.OUT.n205 CM_MSB_V2_0.OUT.n204 1.3655
R347 CM_MSB_V2_0.OUT.n209 CM_MSB_V2_0.OUT.t14 1.3655
R348 CM_MSB_V2_0.OUT.n209 CM_MSB_V2_0.OUT.n208 1.3655
R349 CM_MSB_V2_0.OUT.n213 CM_MSB_V2_0.OUT.t16 1.3655
R350 CM_MSB_V2_0.OUT.n213 CM_MSB_V2_0.OUT.n212 1.3655
R351 CM_MSB_V2_0.OUT.n217 CM_MSB_V2_0.OUT.t6 1.3655
R352 CM_MSB_V2_0.OUT.n217 CM_MSB_V2_0.OUT.n216 1.3655
R353 CM_MSB_V2_0.OUT.n221 CM_MSB_V2_0.OUT.t158 1.3655
R354 CM_MSB_V2_0.OUT.n221 CM_MSB_V2_0.OUT.n220 1.3655
R355 CM_MSB_V2_0.OUT.n225 CM_MSB_V2_0.OUT.t8 1.3655
R356 CM_MSB_V2_0.OUT.n225 CM_MSB_V2_0.OUT.n224 1.3655
R357 CM_MSB_V2_0.OUT.n227 CM_MSB_V2_0.OUT.t3 1.3655
R358 CM_MSB_V2_0.OUT.n227 CM_MSB_V2_0.OUT.n226 1.3655
R359 CM_MSB_V2_0.OUT.n223 CM_MSB_V2_0.OUT.t11 1.3655
R360 CM_MSB_V2_0.OUT.n223 CM_MSB_V2_0.OUT.n222 1.3655
R361 CM_MSB_V2_0.OUT.n219 CM_MSB_V2_0.OUT.t102 1.3655
R362 CM_MSB_V2_0.OUT.n219 CM_MSB_V2_0.OUT.n218 1.3655
R363 CM_MSB_V2_0.OUT.n215 CM_MSB_V2_0.OUT.t18 1.3655
R364 CM_MSB_V2_0.OUT.n215 CM_MSB_V2_0.OUT.n214 1.3655
R365 CM_MSB_V2_0.OUT.n211 CM_MSB_V2_0.OUT.t85 1.3655
R366 CM_MSB_V2_0.OUT.n211 CM_MSB_V2_0.OUT.n210 1.3655
R367 CM_MSB_V2_0.OUT.n207 CM_MSB_V2_0.OUT.t10 1.3655
R368 CM_MSB_V2_0.OUT.n207 CM_MSB_V2_0.OUT.n206 1.3655
R369 CM_MSB_V2_0.OUT.n203 CM_MSB_V2_0.OUT.t0 1.3655
R370 CM_MSB_V2_0.OUT.n203 CM_MSB_V2_0.OUT.n202 1.3655
R371 CM_MSB_V2_0.OUT.n199 CM_MSB_V2_0.OUT.t156 1.3655
R372 CM_MSB_V2_0.OUT.n199 CM_MSB_V2_0.OUT.n198 1.3655
R373 CM_MSB_V2_0.OUT.n143 CM_MSB_V2_0.OUT.n142 0.583357
R374 CM_MSB_V2_0.OUT.n153 CM_MSB_V2_0.OUT.n152 0.583357
R375 CM_MSB_V2_0.OUT.n33 CM_MSB_V2_0.OUT.n32 0.583357
R376 CM_MSB_V2_0.OUT.n13 CM_MSB_V2_0.OUT.n12 0.583357
R377 CM_MSB_V2_0.OUT.n23 CM_MSB_V2_0.OUT.n22 0.583357
R378 CM_MSB_V2_0.OUT.n183 CM_MSB_V2_0.OUT.n180 0.583357
R379 CM_MSB_V2_0.OUT.n54 CM_MSB_V2_0.OUT.n33 0.521929
R380 CM_MSB_V2_0.OUT.n68 CM_MSB_V2_0.OUT.n13 0.521929
R381 CM_MSB_V2_0.OUT.n61 CM_MSB_V2_0.OUT.n23 0.521929
R382 CM_MSB_V2_0.OUT.n167 CM_MSB_V2_0.OUT.n143 0.5105
R383 CM_MSB_V2_0.OUT.n160 CM_MSB_V2_0.OUT.n153 0.5105
R384 CM_MSB_V2_0.OUT.n243 CM_MSB_V2_0.OUT.n242 0.5105
R385 CM_MSB_V2_0.OUT.n242 CM_MSB_V2_0.OUT.n241 0.5105
R386 CM_MSB_V2_0.OUT.n241 CM_MSB_V2_0.OUT.n240 0.5105
R387 CM_MSB_V2_0.OUT.n240 CM_MSB_V2_0.OUT.n239 0.5105
R388 CM_MSB_V2_0.OUT.n239 CM_MSB_V2_0.OUT.n238 0.5105
R389 CM_MSB_V2_0.OUT.n238 CM_MSB_V2_0.OUT.n237 0.5105
R390 CM_MSB_V2_0.OUT.n237 CM_MSB_V2_0.OUT.n236 0.5105
R391 CM_MSB_V2_0.OUT.n236 CM_MSB_V2_0.OUT.n235 0.5105
R392 CM_MSB_V2_0.OUT.n235 CM_MSB_V2_0.OUT.n234 0.5105
R393 CM_MSB_V2_0.OUT.n234 CM_MSB_V2_0.OUT.n233 0.5105
R394 CM_MSB_V2_0.OUT.n233 CM_MSB_V2_0.OUT.n232 0.5105
R395 CM_MSB_V2_0.OUT.n232 CM_MSB_V2_0.OUT.n231 0.5105
R396 CM_MSB_V2_0.OUT.n231 CM_MSB_V2_0.OUT.n230 0.5105
R397 CM_MSB_V2_0.OUT.n230 CM_MSB_V2_0.OUT.n229 0.5105
R398 CM_MSB_V2_0.OUT.n229 CM_MSB_V2_0.OUT.n228 0.5105
R399 CM_MSB_V2_0.OUT.n184 CM_MSB_V2_0.OUT.n183 0.5105
R400 CM_MSB_V2_0.OUT.n193 CM_MSB_V2_0.OUT.n192 0.41094
R401 CM_MSB_V2_0.OUT.n195 CM_MSB_V2_0.OUT.n194 0.406984
R402 CM_MSB_V2_0.OUT.n192 CM_MSB_V2_0.OUT.n191 0.405005
R403 CM_MSB_V2_0.OUT.n196 CM_MSB_V2_0.OUT.n195 0.404016
R404 CM_MSB_V2_0.OUT.n53 CM_MSB_V2_0.OUT.n50 0.401049
R405 CM_MSB_V2_0.OUT.n60 CM_MSB_V2_0.OUT.n57 0.401049
R406 CM_MSB_V2_0.OUT.n67 CM_MSB_V2_0.OUT.n64 0.401049
R407 CM_MSB_V2_0.OUT.n74 CM_MSB_V2_0.OUT.n71 0.401049
R408 CM_MSB_V2_0.OUT.n80 CM_MSB_V2_0.OUT.n77 0.401049
R409 CM_MSB_V2_0.OUT.n87 CM_MSB_V2_0.OUT.n84 0.401049
R410 CM_MSB_V2_0.OUT.n94 CM_MSB_V2_0.OUT.n91 0.401049
R411 CM_MSB_V2_0.OUT.n101 CM_MSB_V2_0.OUT.n98 0.401049
R412 CM_MSB_V2_0.OUT.n107 CM_MSB_V2_0.OUT.n104 0.401049
R413 CM_MSB_V2_0.OUT.n114 CM_MSB_V2_0.OUT.n111 0.401049
R414 CM_MSB_V2_0.OUT.n121 CM_MSB_V2_0.OUT.n118 0.401049
R415 CM_MSB_V2_0.OUT.n128 CM_MSB_V2_0.OUT.n125 0.401049
R416 CM_MSB_V2_0.OUT.n159 CM_MSB_V2_0.OUT.n156 0.401049
R417 CM_MSB_V2_0.OUT.n166 CM_MSB_V2_0.OUT.n163 0.401049
R418 CM_MSB_V2_0.OUT.n173 CM_MSB_V2_0.OUT.n170 0.401049
R419 CM_MSB_V2_0.OUT.n190 CM_MSB_V2_0.OUT.n187 0.401049
R420 CM_MSB_V2_0.OUT.n194 CM_MSB_V2_0.OUT.n193 0.399071
R421 CM_MSB_V2_0.OUT.n191 CM_MSB_V2_0.OUT.n133 0.398082
R422 CM_MSB_V2_0.OUT.n47 CM_MSB_V2_0.OUT.n46 0.382477
R423 CM_MSB_V2_0.OUT.n39 CM_MSB_V2_0.OUT.n38 0.374105
R424 CM_MSB_V2_0.OUT.n41 CM_MSB_V2_0.OUT.n40 0.33957
R425 CM_MSB_V2_0.OUT CM_MSB_V2_0.OUT.n243 0.33675
R426 CM_MSB_V2_0.OUT.n40 CM_MSB_V2_0.OUT.n39 0.333291
R427 CM_MSB_V2_0.OUT.n47 CM_MSB_V2_0.OUT.n41 0.327012
R428 CM_MSB_V2_0.OUT.n50 CM_MSB_V2_0.OUT.n47 0.226984
R429 CM_MSB_V2_0.OUT.n57 CM_MSB_V2_0.OUT.n54 0.215115
R430 CM_MSB_V2_0.OUT.n64 CM_MSB_V2_0.OUT.n61 0.215115
R431 CM_MSB_V2_0.OUT.n71 CM_MSB_V2_0.OUT.n68 0.215115
R432 CM_MSB_V2_0.OUT.n84 CM_MSB_V2_0.OUT.n81 0.215115
R433 CM_MSB_V2_0.OUT.n91 CM_MSB_V2_0.OUT.n88 0.215115
R434 CM_MSB_V2_0.OUT.n98 CM_MSB_V2_0.OUT.n95 0.215115
R435 CM_MSB_V2_0.OUT.n111 CM_MSB_V2_0.OUT.n108 0.215115
R436 CM_MSB_V2_0.OUT.n118 CM_MSB_V2_0.OUT.n115 0.215115
R437 CM_MSB_V2_0.OUT.n125 CM_MSB_V2_0.OUT.n122 0.215115
R438 CM_MSB_V2_0.OUT.n163 CM_MSB_V2_0.OUT.n160 0.215115
R439 CM_MSB_V2_0.OUT.n170 CM_MSB_V2_0.OUT.n167 0.215115
R440 CM_MSB_V2_0.OUT.n187 CM_MSB_V2_0.OUT.n184 0.215115
R441 CM_MSB_V2_0.OUT.n54 CM_MSB_V2_0.OUT.n53 0.173577
R442 CM_MSB_V2_0.OUT.n61 CM_MSB_V2_0.OUT.n60 0.173577
R443 CM_MSB_V2_0.OUT.n68 CM_MSB_V2_0.OUT.n67 0.173577
R444 CM_MSB_V2_0.OUT.n81 CM_MSB_V2_0.OUT.n80 0.173577
R445 CM_MSB_V2_0.OUT.n88 CM_MSB_V2_0.OUT.n87 0.173577
R446 CM_MSB_V2_0.OUT.n95 CM_MSB_V2_0.OUT.n94 0.173577
R447 CM_MSB_V2_0.OUT.n108 CM_MSB_V2_0.OUT.n107 0.173577
R448 CM_MSB_V2_0.OUT.n115 CM_MSB_V2_0.OUT.n114 0.173577
R449 CM_MSB_V2_0.OUT.n122 CM_MSB_V2_0.OUT.n121 0.173577
R450 CM_MSB_V2_0.OUT.n160 CM_MSB_V2_0.OUT.n159 0.173577
R451 CM_MSB_V2_0.OUT.n167 CM_MSB_V2_0.OUT.n166 0.173577
R452 CM_MSB_V2_0.OUT.n184 CM_MSB_V2_0.OUT.n173 0.173577
R453 CM_MSB_V2_0.OUT.n194 CM_MSB_V2_0.OUT.n74 0.119181
R454 CM_MSB_V2_0.OUT.n193 CM_MSB_V2_0.OUT.n101 0.119181
R455 CM_MSB_V2_0.OUT.n192 CM_MSB_V2_0.OUT.n128 0.119181
R456 CM_MSB_V2_0.OUT.n191 CM_MSB_V2_0.OUT.n190 0.119181
R457 IOUT-.n89 IOUT-.t41 9.52957
R458 IOUT-.n18 IOUT-.t59 9.52957
R459 IOUT-.n41 IOUT-.t50 9.52957
R460 IOUT-.n65 IOUT-.t12 9.52957
R461 IOUT-.n93 IOUT-.n71 8.25388
R462 IOUT-.n22 IOUT-.n0 8.25388
R463 IOUT-.n45 IOUT-.n23 8.25388
R464 IOUT-.n69 IOUT-.n47 8.25388
R465 IOUT-.n78 IOUT-.n77 6.83298
R466 IOUT-.n7 IOUT-.n6 6.83298
R467 IOUT-.n30 IOUT-.n29 6.83298
R468 IOUT-.n54 IOUT-.n53 6.83298
R469 IOUT-.n82 IOUT-.n81 5.5481
R470 IOUT-.n79 IOUT-.n73 5.5481
R471 IOUT-.n78 IOUT-.n75 5.5481
R472 IOUT-.n11 IOUT-.n10 5.5481
R473 IOUT-.n8 IOUT-.n2 5.5481
R474 IOUT-.n7 IOUT-.n4 5.5481
R475 IOUT-.n34 IOUT-.n33 5.5481
R476 IOUT-.n31 IOUT-.n25 5.5481
R477 IOUT-.n30 IOUT-.n27 5.5481
R478 IOUT-.n58 IOUT-.n57 5.5481
R479 IOUT-.n55 IOUT-.n49 5.5481
R480 IOUT-.n54 IOUT-.n51 5.5481
R481 IOUT-.n89 IOUT-.n88 5.53001
R482 IOUT-.n18 IOUT-.n17 5.53001
R483 IOUT-.n41 IOUT-.n40 5.53001
R484 IOUT-.n65 IOUT-.n64 5.53001
R485 IOUT-.n90 IOUT-.n86 5.52516
R486 IOUT-.n19 IOUT-.n15 5.52516
R487 IOUT-.n42 IOUT-.n38 5.52516
R488 IOUT-.n66 IOUT-.n62 5.52516
R489 IOUT-.n91 IOUT-.n84 5.51961
R490 IOUT-.n20 IOUT-.n13 5.51961
R491 IOUT-.n43 IOUT-.n36 5.51961
R492 IOUT-.n67 IOUT-.n60 5.51961
R493 IOUT-.n84 IOUT-.t4 2.7305
R494 IOUT-.n84 IOUT-.n83 2.7305
R495 IOUT-.n86 IOUT-.t57 2.7305
R496 IOUT-.n86 IOUT-.n85 2.7305
R497 IOUT-.n88 IOUT-.t6 2.7305
R498 IOUT-.n88 IOUT-.n87 2.7305
R499 IOUT-.n81 IOUT-.t2 2.7305
R500 IOUT-.n81 IOUT-.n80 2.7305
R501 IOUT-.n73 IOUT-.t55 2.7305
R502 IOUT-.n73 IOUT-.n72 2.7305
R503 IOUT-.n75 IOUT-.t30 2.7305
R504 IOUT-.n75 IOUT-.n74 2.7305
R505 IOUT-.n77 IOUT-.t56 2.7305
R506 IOUT-.n77 IOUT-.n76 2.7305
R507 IOUT-.n13 IOUT-.t31 2.7305
R508 IOUT-.n13 IOUT-.n12 2.7305
R509 IOUT-.n15 IOUT-.t19 2.7305
R510 IOUT-.n15 IOUT-.n14 2.7305
R511 IOUT-.n17 IOUT-.t32 2.7305
R512 IOUT-.n17 IOUT-.n16 2.7305
R513 IOUT-.n10 IOUT-.t26 2.7305
R514 IOUT-.n10 IOUT-.n9 2.7305
R515 IOUT-.n2 IOUT-.t15 2.7305
R516 IOUT-.n2 IOUT-.n1 2.7305
R517 IOUT-.n4 IOUT-.t52 2.7305
R518 IOUT-.n4 IOUT-.n3 2.7305
R519 IOUT-.n6 IOUT-.t18 2.7305
R520 IOUT-.n6 IOUT-.n5 2.7305
R521 IOUT-.n36 IOUT-.t17 2.7305
R522 IOUT-.n36 IOUT-.n35 2.7305
R523 IOUT-.n38 IOUT-.t1 2.7305
R524 IOUT-.n38 IOUT-.n37 2.7305
R525 IOUT-.n40 IOUT-.t20 2.7305
R526 IOUT-.n40 IOUT-.n39 2.7305
R527 IOUT-.n33 IOUT-.t53 2.7305
R528 IOUT-.n33 IOUT-.n32 2.7305
R529 IOUT-.n25 IOUT-.t42 2.7305
R530 IOUT-.n25 IOUT-.n24 2.7305
R531 IOUT-.n27 IOUT-.t16 2.7305
R532 IOUT-.n27 IOUT-.n26 2.7305
R533 IOUT-.n29 IOUT-.t45 2.7305
R534 IOUT-.n29 IOUT-.n28 2.7305
R535 IOUT-.n60 IOUT-.t44 2.7305
R536 IOUT-.n60 IOUT-.n59 2.7305
R537 IOUT-.n62 IOUT-.t33 2.7305
R538 IOUT-.n62 IOUT-.n61 2.7305
R539 IOUT-.n64 IOUT-.t47 2.7305
R540 IOUT-.n64 IOUT-.n63 2.7305
R541 IOUT-.n57 IOUT-.t21 2.7305
R542 IOUT-.n57 IOUT-.n56 2.7305
R543 IOUT-.n49 IOUT-.t3 2.7305
R544 IOUT-.n49 IOUT-.n48 2.7305
R545 IOUT-.n51 IOUT-.t43 2.7305
R546 IOUT-.n51 IOUT-.n50 2.7305
R547 IOUT-.n53 IOUT-.t5 2.7305
R548 IOUT-.n53 IOUT-.n52 2.7305
R549 IOUT-.n46 IOUT-.n22 1.46638
R550 IOUT- IOUT-.n70 1.44371
R551 IOUT-.n91 IOUT-.n90 1.28037
R552 IOUT-.n20 IOUT-.n19 1.28037
R553 IOUT-.n43 IOUT-.n42 1.28037
R554 IOUT-.n67 IOUT-.n66 1.28037
R555 IOUT-.n79 IOUT-.n78 1.27854
R556 IOUT-.n8 IOUT-.n7 1.27854
R557 IOUT-.n31 IOUT-.n30 1.27854
R558 IOUT-.n55 IOUT-.n54 1.27854
R559 IOUT-.n82 IOUT-.n79 1.27492
R560 IOUT-.n11 IOUT-.n8 1.27492
R561 IOUT-.n34 IOUT-.n31 1.27492
R562 IOUT-.n58 IOUT-.n55 1.27492
R563 IOUT-.n90 IOUT-.n89 1.26834
R564 IOUT-.n19 IOUT-.n18 1.26834
R565 IOUT-.n42 IOUT-.n41 1.26834
R566 IOUT-.n66 IOUT-.n65 1.26834
R567 IOUT-.n70 IOUT-.n46 1.19621
R568 IOUT-.n93 IOUT-.n92 0.637571
R569 IOUT-.n22 IOUT-.n21 0.637571
R570 IOUT-.n45 IOUT-.n44 0.637571
R571 IOUT-.n69 IOUT-.n68 0.637571
R572 IOUT-.n92 IOUT-.n91 0.636636
R573 IOUT-.n21 IOUT-.n20 0.636636
R574 IOUT-.n44 IOUT-.n43 0.636636
R575 IOUT-.n68 IOUT-.n67 0.636636
R576 IOUT-.n92 IOUT-.n82 0.550143
R577 IOUT-.n21 IOUT-.n11 0.550143
R578 IOUT-.n44 IOUT-.n34 0.550143
R579 IOUT-.n68 IOUT-.n58 0.550143
R580 IOUT-.n46 IOUT-.n45 0.270661
R581 IOUT-.n70 IOUT-.n69 0.270661
R582 IOUT- IOUT-.n93 0.026375
R583 VSS.t60 VSS.n15 2763.56
R584 VSS.t31 VSS.n399 2739.78
R585 VSS.n12 VSS.n11 2723.91
R586 VSS.n390 VSS.n12 2381.26
R587 VSS.t64 VSS.n22 2298.26
R588 VSS.t56 VSS.n391 2273.61
R589 VSS.n14 VSS.t25 2129.07
R590 VSS.t30 VSS.n14 2122.02
R591 VSS.n398 VSS.t71 2106.22
R592 VSS.t59 VSS.n398 2102.28
R593 VSS.n390 VSS.t86 1424.08
R594 VSS.t3 VSS.n390 1408.8
R595 VSS.t86 VSS.n23 599.241
R596 VSS.n13 VSS.t24 599.241
R597 VSS.n16 VSS.t30 599.241
R598 VSS.n400 VSS.t59 594.087
R599 VSS.n392 VSS.t3 592.812
R600 VSS.n397 VSS.t7 592.812
R601 VSS.n23 VSS.t64 528.742
R602 VSS.t25 VSS.n13 528.742
R603 VSS.n16 VSS.t60 528.742
R604 VSS.n400 VSS.t31 524.194
R605 VSS.n392 VSS.t56 523.069
R606 VSS.t71 VSS.n397 523.069
R607 VSS.n422 VSS.t9 233.171
R608 VSS.n377 VSS.t39 214.006
R609 VSS.n3 VSS.t36 135.75
R610 VSS.n7 VSS.t27 119.779
R611 VSS.n376 VSS.t17 105.406
R612 VSS.t17 VSS.n31 102.212
R613 VSS.t2 VSS.t116 99.0177
R614 VSS.n370 VSS.t93 91.0324
R615 VSS.n411 VSS.t15 86.2413
R616 VSS.n419 VSS.t119 79.8531
R617 VSS.n416 VSS.t5 67.0767
R618 VSS.n428 VSS.t14 60.6885
R619 VSS.n204 VSS.t51 51.4643
R620 VSS.t5 VSS.n415 47.912
R621 VSS.n95 VSS.t21 45.4802
R622 VSS.n360 VSS.t12 43.0865
R623 VSS.n380 VSS.t13 41.5238
R624 VSS.n352 VSS.t34 38.2992
R625 VSS.n390 VSS.t62 38.2992
R626 VSS.n348 VSS.t11 35.9055
R627 VSS.n339 VSS.t33 31.1182
R628 VSS.t93 VSS.t0 28.7474
R629 VSS.n333 VSS.t58 28.7245
R630 VSS.n32 VSS.t2 25.5533
R631 VSS.n324 VSS.t20 23.9372
R632 VSS.n319 VSS.t6 21.5435
R633 VSS.t14 VSS.t37 20.7622
R634 VSS.n308 VSS.t73 16.7562
R635 VSS.n239 VSS.t43 15.5593
R636 VSS.n302 VSS.t63 14.3625
R637 VSS.n296 VSS.t19 11.9688
R638 VSS.n35 VSS.n33 11.2304
R639 VSS.n375 VSS.n35 11.2304
R640 VSS.n430 VSS.n412 11.2304
R641 VSS.n407 VSS.n405 11.2304
R642 VSS.t68 VSS.t40 9.57516
R643 VSS.t35 VSS.t42 9.57516
R644 VSS.t10 VSS.t48 9.57516
R645 VSS.t18 VSS.t44 9.57516
R646 VSS.n291 VSS.t4 9.57516
R647 VSS.t4 VSS.t49 9.57516
R648 VSS.t63 VSS.t47 9.57516
R649 VSS.t73 VSS.t41 9.57516
R650 VSS.t55 VSS.t16 9.57516
R651 VSS.t6 VSS.t54 9.57516
R652 VSS.t20 VSS.t52 9.57516
R653 VSS.t46 VSS.t97 9.57516
R654 VSS.t58 VSS.t53 9.57516
R655 VSS.t33 VSS.t45 9.57516
R656 VSS.n417 VSS.n416 8.98871
R657 VSS.n230 VSS.t55 8.37833
R658 VSS.t62 VSS.n389 8.37833
R659 VSS.n285 VSS.t18 7.1815
R660 VSS.n20 VSS.t65 6.65541
R661 VSS.n18 VSS.t26 6.65541
R662 VSS.n10 VSS.t61 6.65541
R663 VSS.n9 VSS.t28 6.65541
R664 VSS.n394 VSS.t57 6.65541
R665 VSS.n395 VSS.t72 6.65541
R666 VSS.n402 VSS.t32 6.65541
R667 VSS.n372 VSS.t1 6.65541
R668 VSS.n4 VSS.t38 6.65541
R669 VSS.n377 VSS.n376 6.38871
R670 VSS.n429 VSS.n428 6.38871
R671 VSS.t119 VSS.t8 6.38871
R672 VSS.n261 VSS.n260 6.21452
R673 VSS.n401 VSS.n400 5.2005
R674 VSS.n393 VSS.n392 5.2005
R675 VSS.n397 VSS.n396 5.2005
R676 VSS.n8 VSS.n7 5.2005
R677 VSS.n23 VSS.n21 5.2005
R678 VSS.n19 VSS.n13 5.2005
R679 VSS.n17 VSS.n16 5.2005
R680 VSS.n371 VSS.n370 5.2005
R681 VSS.n432 VSS.n3 5.2005
R682 VSS.n418 VSS.t82 5.13332
R683 VSS.n260 VSS.n184 5.10637
R684 VSS.n279 VSS.t10 4.78783
R685 VSS.n403 VSS.n10 3.81335
R686 VSS.n409 VSS.n6 3.78833
R687 VSS.n355 VSS.n100 3.78833
R688 VSS.n336 VSS.n102 3.78833
R689 VSS.n317 VSS.n104 3.78833
R690 VSS.n294 VSS.n106 3.78833
R691 VSS.n271 VSS.n108 3.78833
R692 VSS.n368 VSS.n37 3.78833
R693 VSS.n2 VSS.n1 3.78833
R694 VSS.n247 VSS.n186 3.74137
R695 VSS.n238 VSS.n188 3.74137
R696 VSS.n224 VSS.n190 3.74137
R697 VSS.n208 VSS.n192 3.74137
R698 VSS.n28 VSS.n27 3.74137
R699 VSS.n383 VSS.n30 3.74137
R700 VSS.n425 VSS.n414 3.74137
R701 VSS.n404 VSS.n403 3.68866
R702 VSS.n210 VSS.t29 3.591
R703 VSS.n211 VSS.t50 3.591
R704 VSS.n152 VSS.n151 2.64635
R705 VSS.n155 VSS.n154 2.64635
R706 VSS.n158 VSS.n157 2.64635
R707 VSS.n183 VSS.n111 2.60322
R708 VSS.n405 VSS.n404 2.6005
R709 VSS.n412 VSS.n410 2.6005
R710 VSS.n412 VSS.n411 2.6005
R711 VSS.n408 VSS.n407 2.6005
R712 VSS.n407 VSS.n406 2.6005
R713 VSS.n386 VSS.n385 2.6005
R714 VSS.n385 VSS.n384 2.6005
R715 VSS.n382 VSS.n381 2.6005
R716 VSS.n381 VSS.n380 2.6005
R717 VSS.n379 VSS.n378 2.6005
R718 VSS.n378 VSS.n377 2.6005
R719 VSS.n427 VSS.n426 2.6005
R720 VSS.n428 VSS.n427 2.6005
R721 VSS.n424 VSS.n423 2.6005
R722 VSS.n423 VSS.n422 2.6005
R723 VSS.n421 VSS.n420 2.6005
R724 VSS.n420 VSS.n419 2.6005
R725 VSS.n418 VSS.n417 2.6005
R726 VSS.n259 VSS.n258 2.6005
R727 VSS.n258 VSS.n257 2.6005
R728 VSS.n255 VSS.n254 2.6005
R729 VSS.n254 VSS.n253 2.6005
R730 VSS.n251 VSS.n250 2.6005
R731 VSS.n250 VSS.n249 2.6005
R732 VSS.n246 VSS.n245 2.6005
R733 VSS.n245 VSS.n244 2.6005
R734 VSS.n242 VSS.n241 2.6005
R735 VSS.n241 VSS.n240 2.6005
R736 VSS.n237 VSS.n236 2.6005
R737 VSS.n236 VSS.n235 2.6005
R738 VSS.n233 VSS.n232 2.6005
R739 VSS.n232 VSS.n231 2.6005
R740 VSS.n229 VSS.n228 2.6005
R741 VSS.n228 VSS.n227 2.6005
R742 VSS.n223 VSS.n222 2.6005
R743 VSS.n222 VSS.n221 2.6005
R744 VSS.n218 VSS.n217 2.6005
R745 VSS.n217 VSS.n216 2.6005
R746 VSS.n213 VSS.n212 2.6005
R747 VSS.n212 VSS.n211 2.6005
R748 VSS.n207 VSS.n206 2.6005
R749 VSS.n206 VSS.n205 2.6005
R750 VSS.n202 VSS.n201 2.6005
R751 VSS.n201 VSS.n200 2.6005
R752 VSS.n197 VSS.n196 2.6005
R753 VSS.n196 VSS.n195 2.6005
R754 VSS.n388 VSS.n387 2.6005
R755 VSS.n389 VSS.n388 2.6005
R756 VSS.n98 VSS.n97 2.6005
R757 VSS.n58 VSS.n57 2.6005
R758 VSS.n60 VSS.n59 2.6005
R759 VSS.n62 VSS.n61 2.6005
R760 VSS.n64 VSS.n63 2.6005
R761 VSS.n66 VSS.n65 2.6005
R762 VSS.n68 VSS.n67 2.6005
R763 VSS.n70 VSS.n69 2.6005
R764 VSS.n72 VSS.n71 2.6005
R765 VSS.n74 VSS.n73 2.6005
R766 VSS.n76 VSS.n75 2.6005
R767 VSS.n78 VSS.n77 2.6005
R768 VSS.n80 VSS.n79 2.6005
R769 VSS.n82 VSS.n81 2.6005
R770 VSS.n85 VSS.n84 2.6005
R771 VSS.n87 VSS.n86 2.6005
R772 VSS.n56 VSS.n55 2.6005
R773 VSS.n54 VSS.n53 2.6005
R774 VSS.n122 VSS.n121 2.6005
R775 VSS.n110 VSS.n109 2.6005
R776 VSS.n263 VSS.n262 2.6005
R777 VSS.t68 VSS.n268 2.6005
R778 VSS.n275 VSS.n274 2.6005
R779 VSS.n279 VSS.n278 2.6005
R780 VSS.n285 VSS.n284 2.6005
R781 VSS.n291 VSS.n290 2.6005
R782 VSS.n296 VSS.n295 2.6005
R783 VSS.n302 VSS.n301 2.6005
R784 VSS.n308 VSS.n307 2.6005
R785 VSS.n312 VSS.n311 2.6005
R786 VSS.n319 VSS.n318 2.6005
R787 VSS.n324 VSS.n323 2.6005
R788 VSS.n328 VSS.n327 2.6005
R789 VSS.n333 VSS.n332 2.6005
R790 VSS.n339 VSS.n338 2.6005
R791 VSS.n343 VSS.n342 2.6005
R792 VSS.n348 VSS.n347 2.6005
R793 VSS.n48 VSS.n47 2.6005
R794 VSS.n50 VSS.n49 2.6005
R795 VSS.n52 VSS.n51 2.6005
R796 VSS.n126 VSS.n125 2.6005
R797 VSS.n176 VSS.n175 2.6005
R798 VSS.n159 VSS.n158 2.6005
R799 VSS.n156 VSS.n155 2.6005
R800 VSS.n153 VSS.n152 2.6005
R801 VSS.n150 VSS.n149 2.6005
R802 VSS.n148 VSS.n147 2.6005
R803 VSS.n146 VSS.n145 2.6005
R804 VSS.n144 VSS.n143 2.6005
R805 VSS.n142 VSS.n141 2.6005
R806 VSS.n140 VSS.n139 2.6005
R807 VSS.n138 VSS.n137 2.6005
R808 VSS.n136 VSS.n135 2.6005
R809 VSS.n134 VSS.n133 2.6005
R810 VSS.n132 VSS.n131 2.6005
R811 VSS.n130 VSS.n129 2.6005
R812 VSS.n128 VSS.n127 2.6005
R813 VSS.n124 VSS.n123 2.6005
R814 VSS.n179 VSS.n178 2.6005
R815 VSS.n182 VSS.n181 2.6005
R816 VSS.n181 VSS.n180 2.6005
R817 VSS.n366 VSS.n365 2.6005
R818 VSS.n362 VSS.n361 2.6005
R819 VSS.n361 VSS.n360 2.6005
R820 VSS.n358 VSS.n357 2.6005
R821 VSS.n357 VSS.n356 2.6005
R822 VSS.n354 VSS.n353 2.6005
R823 VSS.n353 VSS.n352 2.6005
R824 VSS.n350 VSS.n349 2.6005
R825 VSS.n349 VSS.n348 2.6005
R826 VSS.n345 VSS.n344 2.6005
R827 VSS.n344 VSS.n343 2.6005
R828 VSS.n341 VSS.n340 2.6005
R829 VSS.n340 VSS.n339 2.6005
R830 VSS.n335 VSS.n334 2.6005
R831 VSS.n334 VSS.n333 2.6005
R832 VSS.n330 VSS.n329 2.6005
R833 VSS.n329 VSS.n328 2.6005
R834 VSS.n326 VSS.n325 2.6005
R835 VSS.n325 VSS.n324 2.6005
R836 VSS.n321 VSS.n320 2.6005
R837 VSS.n320 VSS.n319 2.6005
R838 VSS.n314 VSS.n313 2.6005
R839 VSS.n313 VSS.n312 2.6005
R840 VSS.n310 VSS.n309 2.6005
R841 VSS.n309 VSS.n308 2.6005
R842 VSS.n304 VSS.n303 2.6005
R843 VSS.n303 VSS.n302 2.6005
R844 VSS.n298 VSS.n297 2.6005
R845 VSS.n297 VSS.n296 2.6005
R846 VSS.n293 VSS.n292 2.6005
R847 VSS.n292 VSS.n291 2.6005
R848 VSS.n287 VSS.n286 2.6005
R849 VSS.n286 VSS.n285 2.6005
R850 VSS.n281 VSS.n280 2.6005
R851 VSS.n280 VSS.n279 2.6005
R852 VSS.n277 VSS.n276 2.6005
R853 VSS.n276 VSS.n275 2.6005
R854 VSS.n270 VSS.n269 2.6005
R855 VSS.n269 VSS.t68 2.6005
R856 VSS.n265 VSS.n264 2.6005
R857 VSS.n264 VSS.n263 2.6005
R858 VSS.n111 VSS.n110 2.6005
R859 VSS.n273 VSS.n272 2.6005
R860 VSS.n283 VSS.n282 2.6005
R861 VSS.n289 VSS.n288 2.6005
R862 VSS.n300 VSS.n299 2.6005
R863 VSS.n306 VSS.n305 2.6005
R864 VSS.n316 VSS.n315 2.6005
R865 VSS.n226 VSS.n225 2.6005
R866 VSS.n220 VSS.n219 2.6005
R867 VSS.n215 VSS.n214 2.6005
R868 VSS.n210 VSS.n209 2.6005
R869 VSS.n204 VSS.n203 2.6005
R870 VSS.n199 VSS.n198 2.6005
R871 VSS.n194 VSS.n193 2.6005
R872 VSS.n267 VSS.n266 2.6005
R873 VSS.n25 VSS.n24 2.6005
R874 VSS.n33 VSS.n32 2.6005
R875 VSS.n373 VSS.n35 2.6005
R876 VSS.n35 VSS.n34 2.6005
R877 VSS.n375 VSS.n374 2.6005
R878 VSS.n376 VSS.n375 2.6005
R879 VSS.n431 VSS.n430 2.6005
R880 VSS.n430 VSS.n429 2.6005
R881 VSS.n403 VSS.n402 2.53474
R882 VSS.n263 VSS.t113 2.39417
R883 VSS.n257 VSS.n256 2.39417
R884 VSS.n253 VSS.n252 2.39417
R885 VSS.n275 VSS.t35 2.39417
R886 VSS.n249 VSS.n248 2.39417
R887 VSS.n244 VSS.n243 2.39417
R888 VSS.n240 VSS.n239 2.39417
R889 VSS.n235 VSS.n234 2.39417
R890 VSS.n231 VSS.n230 2.39417
R891 VSS.n227 VSS.n226 2.39417
R892 VSS.n221 VSS.n220 2.39417
R893 VSS.n216 VSS.n215 2.39417
R894 VSS.n211 VSS.n210 2.39417
R895 VSS.n205 VSS.n204 2.39417
R896 VSS.n200 VSS.n199 2.39417
R897 VSS.n195 VSS.n194 2.39417
R898 VSS.n389 VSS.n25 2.39417
R899 VSS.n97 VSS.n96 1.75437
R900 VSS.n84 VSS.n83 1.75437
R901 VSS.n175 VSS.n174 1.50887
R902 VSS.n186 VSS.t70 1.3655
R903 VSS.n186 VSS.n185 1.3655
R904 VSS.n188 VSS.t90 1.3655
R905 VSS.n188 VSS.n187 1.3655
R906 VSS.n190 VSS.t122 1.3655
R907 VSS.n190 VSS.n189 1.3655
R908 VSS.n192 VSS.t92 1.3655
R909 VSS.n192 VSS.n191 1.3655
R910 VSS.n27 VSS.t76 1.3655
R911 VSS.n27 VSS.n26 1.3655
R912 VSS.n30 VSS.t94 1.3655
R913 VSS.n30 VSS.n29 1.3655
R914 VSS.n414 VSS.t91 1.3655
R915 VSS.n414 VSS.n413 1.3655
R916 VSS.n6 VSS.t112 1.3655
R917 VSS.n6 VSS.n5 1.3655
R918 VSS.n100 VSS.t85 1.3655
R919 VSS.n100 VSS.n99 1.3655
R920 VSS.n102 VSS.t102 1.3655
R921 VSS.n102 VSS.n101 1.3655
R922 VSS.n104 VSS.t87 1.3655
R923 VSS.n104 VSS.n103 1.3655
R924 VSS.n106 VSS.t111 1.3655
R925 VSS.n106 VSS.n105 1.3655
R926 VSS.n108 VSS.t69 1.3655
R927 VSS.n108 VSS.n107 1.3655
R928 VSS.n37 VSS.t110 1.3655
R929 VSS.n37 VSS.n36 1.3655
R930 VSS.n1 VSS.t77 1.3655
R931 VSS.n1 VSS.n0 1.3655
R932 VSS.n173 VSS.n160 1.27833
R933 VSS.n173 VSS.n161 1.27833
R934 VSS.n173 VSS.n162 1.27833
R935 VSS.n173 VSS.n163 1.27833
R936 VSS.n173 VSS.n164 1.27833
R937 VSS.n173 VSS.n165 1.27833
R938 VSS.n173 VSS.n166 1.27833
R939 VSS.n173 VSS.n167 1.27833
R940 VSS.n173 VSS.n168 1.27833
R941 VSS.n173 VSS.n169 1.27833
R942 VSS.n173 VSS.n170 1.27833
R943 VSS.n173 VSS.n171 1.27833
R944 VSS.n183 VSS.n182 1.2289
R945 VSS.n220 VSS.t46 1.19733
R946 VSS.n200 VSS.t103 1.19733
R947 VSS.n173 VSS.n172 0.729291
R948 VSS.n174 VSS.n173 0.729086
R949 VSS.n20 VSS 0.684889
R950 VSS VSS.n394 0.684889
R951 VSS.n18 VSS 0.620412
R952 VSS.n395 VSS 0.620412
R953 VSS.n96 VSS.n95 0.424314
R954 VSS.n95 VSS.n94 0.424314
R955 VSS.n95 VSS.n93 0.424314
R956 VSS.n95 VSS.n92 0.424314
R957 VSS.n95 VSS.n91 0.424314
R958 VSS.n95 VSS.n90 0.424314
R959 VSS.n95 VSS.n89 0.424314
R960 VSS.n95 VSS.n88 0.424314
R961 VSS.n176 VSS.n159 0.240099
R962 VSS.n159 VSS.n156 0.240099
R963 VSS.n156 VSS.n153 0.240099
R964 VSS.n153 VSS.n150 0.240099
R965 VSS.n150 VSS.n148 0.240099
R966 VSS.n148 VSS.n146 0.240099
R967 VSS.n146 VSS.n144 0.240099
R968 VSS.n144 VSS.n142 0.240099
R969 VSS.n142 VSS.n140 0.240099
R970 VSS.n140 VSS.n138 0.240099
R971 VSS.n138 VSS.n136 0.240099
R972 VSS.n136 VSS.n134 0.240099
R973 VSS.n134 VSS.n132 0.240099
R974 VSS.n132 VSS.n130 0.240099
R975 VSS.n130 VSS.n128 0.240099
R976 VSS.n128 VSS.n126 0.240099
R977 VSS.n58 VSS.n56 0.240099
R978 VSS.n60 VSS.n58 0.240099
R979 VSS.n62 VSS.n60 0.240099
R980 VSS.n64 VSS.n62 0.240099
R981 VSS.n66 VSS.n64 0.240099
R982 VSS.n68 VSS.n66 0.240099
R983 VSS.n70 VSS.n68 0.240099
R984 VSS.n72 VSS.n70 0.240099
R985 VSS.n74 VSS.n72 0.240099
R986 VSS.n76 VSS.n74 0.240099
R987 VSS.n78 VSS.n76 0.240099
R988 VSS.n80 VSS.n78 0.240099
R989 VSS.n82 VSS.n80 0.240099
R990 VSS.n85 VSS.n82 0.240099
R991 VSS.n87 VSS.n85 0.240099
R992 VSS.n98 VSS.n87 0.240099
R993 VSS.n124 VSS.n122 0.234957
R994 VSS.n122 VSS.n120 0.234957
R995 VSS.n120 VSS.n119 0.234957
R996 VSS.n119 VSS.n118 0.234957
R997 VSS.n118 VSS.n117 0.234957
R998 VSS.n117 VSS.n116 0.234957
R999 VSS.n116 VSS.n115 0.234957
R1000 VSS.n115 VSS.n114 0.234957
R1001 VSS.n114 VSS.n113 0.234957
R1002 VSS.n113 VSS.n112 0.234957
R1003 VSS.n39 VSS.n38 0.234957
R1004 VSS.n40 VSS.n39 0.234957
R1005 VSS.n41 VSS.n40 0.234957
R1006 VSS.n42 VSS.n41 0.234957
R1007 VSS.n43 VSS.n42 0.234957
R1008 VSS.n44 VSS.n43 0.234957
R1009 VSS.n45 VSS.n44 0.234957
R1010 VSS.n46 VSS.n45 0.234957
R1011 VSS.n48 VSS.n46 0.234957
R1012 VSS.n50 VSS.n48 0.234957
R1013 VSS.n52 VSS.n50 0.234957
R1014 VSS.n54 VSS.n52 0.234957
R1015 VSS.n182 VSS.n179 0.234957
R1016 VSS.n366 VSS.n98 0.220714
R1017 VSS.n56 VSS.n54 0.209695
R1018 VSS.n126 VSS.n124 0.199945
R1019 VSS.n179 VSS.n176 0.197176
R1020 VSS.n259 VSS.n255 0.144885
R1021 VSS.n255 VSS.n251 0.144885
R1022 VSS.n246 VSS.n242 0.144885
R1023 VSS.n237 VSS.n233 0.144885
R1024 VSS.n233 VSS.n229 0.144885
R1025 VSS.n223 VSS.n218 0.144885
R1026 VSS.n218 VSS.n213 0.144885
R1027 VSS.n207 VSS.n202 0.144885
R1028 VSS.n202 VSS.n197 0.144885
R1029 VSS.n387 VSS.n386 0.144885
R1030 VSS.n382 VSS.n379 0.144885
R1031 VSS.n424 VSS.n421 0.144885
R1032 VSS.n421 VSS.n418 0.144885
R1033 VSS.n21 VSS.n20 0.142847
R1034 VSS.n17 VSS.n10 0.142847
R1035 VSS.n394 VSS.n393 0.142847
R1036 VSS.n396 VSS.n395 0.142847
R1037 VSS.n402 VSS.n401 0.142847
R1038 VSS.n387 VSS.n28 0.141035
R1039 VSS VSS.n18 0.130908
R1040 VSS.n242 VSS.n238 0.125634
R1041 VSS.n247 VSS.n246 0.123709
R1042 VSS.n386 VSS.n383 0.108307
R1043 VSS.n365 VSS.n364 0.108192
R1044 VSS.n178 VSS.n177 0.108192
R1045 VSS.n208 VSS.n207 0.100607
R1046 VSS.n229 VSS.n224 0.0852059
R1047 VSS.n260 VSS.n259 0.0832807
R1048 VSS.n425 VSS.n424 0.0775053
R1049 VSS.n426 VSS.n425 0.0678797
R1050 VSS.n224 VSS.n223 0.0601791
R1051 VSS.n367 VSS.n366 0.055041
R1052 VSS.n410 VSS.n409 0.0549122
R1053 VSS VSS.n2 0.0523246
R1054 VSS.n213 VSS.n208 0.0447781
R1055 VSS.n281 VSS.n277 0.0390439
R1056 VSS.n314 VSS.n310 0.0390439
R1057 VSS.n330 VSS.n326 0.0390439
R1058 VSS.n345 VSS.n341 0.0390439
R1059 VSS.n369 VSS.n368 0.0388886
R1060 VSS.n383 VSS.n382 0.0370775
R1061 VSS.n374 VSS 0.0353367
R1062 VSS.n372 VSS.n371 0.0335569
R1063 VSS.n9 VSS.n8 0.0334787
R1064 VSS.n355 VSS.n354 0.0324914
R1065 VSS.n289 VSS.n287 0.0317206
R1066 VSS.n306 VSS.n304 0.0317206
R1067 VSS.n322 VSS.n321 0.0317206
R1068 VSS.n351 VSS.n350 0.0317206
R1069 VSS.n363 VSS.n362 0.0317206
R1070 VSS VSS.n4 0.0314242
R1071 VSS VSS.n373 0.0307574
R1072 VSS.n408 VSS 0.0307128
R1073 VSS.n336 VSS.n335 0.0294079
R1074 VSS.n431 VSS.n4 0.0292915
R1075 VSS.n270 VSS.n267 0.0270953
R1076 VSS.n287 VSS.n283 0.0270953
R1077 VSS.n304 VSS.n300 0.0270953
R1078 VSS.n335 VSS.n331 0.0270953
R1079 VSS.n350 VSS.n346 0.0270953
R1080 VSS.n362 VSS.n359 0.0270953
R1081 VSS.n368 VSS.n367 0.0260924
R1082 VSS.n265 VSS.n261 0.0253608
R1083 VSS.n294 VSS.n293 0.0232409
R1084 VSS.n251 VSS.n247 0.0216765
R1085 VSS.n271 VSS.n270 0.0201574
R1086 VSS.n238 VSS.n237 0.0197513
R1087 VSS.n373 VSS.n372 0.0167085
R1088 VSS.n298 VSS.n294 0.016303
R1089 VSS VSS.n369 0.0150024
R1090 VSS.n317 VSS.n316 0.0143758
R1091 VSS.n321 VSS.n317 0.0132195
R1092 VSS.n261 VSS.n183 0.0124649
R1093 VSS.n267 VSS.n265 0.0124486
R1094 VSS.n283 VSS.n281 0.0124486
R1095 VSS.n300 VSS.n298 0.0124486
R1096 VSS.n316 VSS.n314 0.0124486
R1097 VSS.n331 VSS.n330 0.0124486
R1098 VSS.n346 VSS.n345 0.0124486
R1099 VSS.n359 VSS.n358 0.0124486
R1100 VSS.n19 VSS 0.0124388
R1101 VSS.n273 VSS.n271 0.0120632
R1102 VSS.n409 VSS.n408 0.0107128
R1103 VSS.n374 VSS.n2 0.00817773
R1104 VSS.n277 VSS.n273 0.00782334
R1105 VSS.n293 VSS.n289 0.00782334
R1106 VSS.n310 VSS.n306 0.00782334
R1107 VSS.n326 VSS.n322 0.00782334
R1108 VSS.n341 VSS.n337 0.00782334
R1109 VSS.n354 VSS.n351 0.00782334
R1110 VSS.n366 VSS.n363 0.00782334
R1111 VSS.n358 VSS.n355 0.00705246
R1112 VSS.n410 VSS 0.00487385
R1113 VSS.n432 VSS.n431 0.0047654
R1114 VSS.n197 VSS.n28 0.00435027
R1115 VSS.n337 VSS.n336 0.00281263
R1116 VSS.n21 VSS 0.00141837
R1117 VSS VSS.n19 0.00141837
R1118 VSS VSS.n17 0.00141837
R1119 VSS.n393 VSS 0.00141837
R1120 VSS.n396 VSS 0.00141837
R1121 VSS.n401 VSS 0.00141837
R1122 VSS.n404 VSS.n9 0.000925532
R1123 VSS.n371 VSS 0.00071327
R1124 VSS VSS.n432 0.00071327
R1125 VSS.n8 VSS 0.000712766
R1126 IM_T.n1 IM_T.t25 84.5899
R1127 IM_T.n3 IM_T.n2 64.4419
R1128 IM_T.n5 IM_T.n4 64.4419
R1129 IM_T.n7 IM_T.n6 64.4419
R1130 IM_T.n9 IM_T.n8 64.4419
R1131 IM_T.n11 IM_T.n10 64.4419
R1132 IM_T.n13 IM_T.n12 64.4419
R1133 IM_T.n15 IM_T.n14 64.4419
R1134 IM_T.n18 IM_T.n17 63.3497
R1135 IM_T.n20 IM_T.n19 63.3497
R1136 IM_T.n22 IM_T.n21 63.3497
R1137 IM_T.n24 IM_T.n23 63.3497
R1138 IM_T.n26 IM_T.n25 63.3497
R1139 IM_T.n28 IM_T.n27 63.3497
R1140 IM_T.n30 IM_T.n29 63.3497
R1141 IM_T.n32 IM_T.n31 57.704
R1142 IM_T.n17 IM_T.t27 31.3373
R1143 IM_T.n16 IM_T.n15 31.1695
R1144 IM_T.n1 IM_T.t21 20.1485
R1145 IM_T.n2 IM_T.t8 20.1485
R1146 IM_T.n3 IM_T.t9 20.1485
R1147 IM_T.n4 IM_T.t12 20.1485
R1148 IM_T.n5 IM_T.t20 20.1485
R1149 IM_T.n6 IM_T.t28 20.1485
R1150 IM_T.n7 IM_T.t7 20.1485
R1151 IM_T.n8 IM_T.t22 20.1485
R1152 IM_T.n9 IM_T.t13 20.1485
R1153 IM_T.n10 IM_T.t5 20.1485
R1154 IM_T.n11 IM_T.t29 20.1485
R1155 IM_T.n12 IM_T.t14 20.1485
R1156 IM_T.n13 IM_T.t6 20.1485
R1157 IM_T.n14 IM_T.t31 20.1485
R1158 IM_T.n15 IM_T.t23 20.1485
R1159 IM_T.n17 IM_T.t4 18.4695
R1160 IM_T.n18 IM_T.t2 18.4695
R1161 IM_T.n19 IM_T.t19 18.4695
R1162 IM_T.n20 IM_T.t15 18.4695
R1163 IM_T.n21 IM_T.t24 18.4695
R1164 IM_T.n22 IM_T.t1 18.4695
R1165 IM_T.n23 IM_T.t17 18.4695
R1166 IM_T.n24 IM_T.t18 18.4695
R1167 IM_T.n25 IM_T.t11 18.4695
R1168 IM_T.n26 IM_T.t10 18.4695
R1169 IM_T.n27 IM_T.t30 18.4695
R1170 IM_T.n28 IM_T.t16 18.4695
R1171 IM_T.n29 IM_T.t0 18.4695
R1172 IM_T.n30 IM_T.t3 18.4695
R1173 IM_T.n31 IM_T.t26 18.4695
R1174 IM_T.n2 IM_T.n1 13.0902
R1175 IM_T.n4 IM_T.n3 13.0902
R1176 IM_T.n6 IM_T.n5 13.0902
R1177 IM_T.n8 IM_T.n7 13.0902
R1178 IM_T.n10 IM_T.n9 13.0902
R1179 IM_T.n12 IM_T.n11 13.0902
R1180 IM_T.n14 IM_T.n13 13.0902
R1181 IM_T.n19 IM_T.n18 12.8683
R1182 IM_T.n21 IM_T.n20 12.8683
R1183 IM_T.n23 IM_T.n22 12.8683
R1184 IM_T.n25 IM_T.n24 12.8683
R1185 IM_T.n27 IM_T.n26 12.8683
R1186 IM_T.n29 IM_T.n28 12.8683
R1187 IM_T.n31 IM_T.n30 12.8683
R1188 IM_T.n0 IM_T 4.52248
R1189 IM_T.n33 IM_T.n16 1.1293
R1190 IM_T.n33 IM_T.n32 0.0277093
R1191 IM_T.n16 IM_T.n0 0.0026666
R1192 IM_T IM_T.n33 0.00154651
R1193 CM_MSB_V2_0.SD.n3 CM_MSB_V2_0.SD.n76 4.5005
R1194 CM_MSB_V2_0.SD.n4 CM_MSB_V2_0.SD.n19 3.63741
R1195 CM_MSB_V2_0.SD.n48 CM_MSB_V2_0.SD.n47 3.28149
R1196 CM_MSB_V2_0.SD.n57 CM_MSB_V2_0.SD.n33 3.28101
R1197 CM_MSB_V2_0.SD.n0 CM_MSB_V2_0.SD.n24 3.27542
R1198 CM_MSB_V2_0.SD.n3 CM_MSB_V2_0.SD.n8 3.26817
R1199 CM_MSB_V2_0.SD.n98 CM_MSB_V2_0.SD.n82 3.258
R1200 CM_MSB_V2_0.SD.n50 CM_MSB_V2_0.SD.n40 3.25644
R1201 CM_MSB_V2_0.SD.n73 CM_MSB_V2_0.SD.n10 3.24511
R1202 CM_MSB_V2_0.SD.n92 CM_MSB_V2_0.SD.n89 3.23798
R1203 CM_MSB_V2_0.SD.n6 CM_MSB_V2_0.SD.n87 3.23061
R1204 CM_MSB_V2_0.SD.n2 CM_MSB_V2_0.SD.n17 3.2111
R1205 CM_MSB_V2_0.SD.n5 CM_MSB_V2_0.SD.n26 3.20644
R1206 CM_MSB_V2_0.SD.n60 CM_MSB_V2_0.SD.n28 3.20496
R1207 CM_MSB_V2_0.SD.n1 CM_MSB_V2_0.SD.n38 3.204
R1208 CM_MSB_V2_0.SD.n100 CM_MSB_V2_0.SD.n80 3.19428
R1209 CM_MSB_V2_0.SD.n105 CM_MSB_V2_0.SD.n78 3.16815
R1210 CM_MSB_V2_0.SD.n103 CM_MSB_V2_0.SD.n102 2.58749
R1211 CM_MSB_V2_0.SD.n72 CM_MSB_V2_0.SD.n12 2.5852
R1212 CM_MSB_V2_0.SD.n48 CM_MSB_V2_0.SD.n45 2.57457
R1213 CM_MSB_V2_0.SD.n92 CM_MSB_V2_0.SD.n91 2.56564
R1214 CM_MSB_V2_0.SD.n1 CM_MSB_V2_0.SD.n54 2.24976
R1215 CM_MSB_V2_0.SD.n65 CM_MSB_V2_0.SD.n64 2.24638
R1216 CM_MSB_V2_0.SD.n96 CM_MSB_V2_0.SD.n95 2.24631
R1217 CM_MSB_V2_0.SD.n70 CM_MSB_V2_0.SD.n69 2.24557
R1218 CM_MSB_V2_0.SD.n109 CM_MSB_V2_0.SD.n108 2.24508
R1219 CM_MSB_V2_0.SD.n59 CM_MSB_V2_0.SD.n31 1.49577
R1220 CM_MSB_V2_0.SD.n97 CM_MSB_V2_0.SD.n85 1.49564
R1221 CM_MSB_V2_0.SD.n2 CM_MSB_V2_0.SD.n15 1.49548
R1222 CM_MSB_V2_0.SD.n49 CM_MSB_V2_0.SD.n43 1.49542
R1223 CM_MSB_V2_0.SD.n0 CM_MSB_V2_0.SD.n22 1.49542
R1224 CM_MSB_V2_0.SD.n56 CM_MSB_V2_0.SD.n36 1.49542
R1225 CM_MSB_V2_0.SD.n102 CM_MSB_V2_0.SD.t0 1.47093
R1226 CM_MSB_V2_0.SD.n33 CM_MSB_V2_0.SD.t42 1.47081
R1227 CM_MSB_V2_0.SD.n8 CM_MSB_V2_0.SD.t27 1.4708
R1228 CM_MSB_V2_0.SD.n24 CM_MSB_V2_0.SD.t4 1.46022
R1229 CM_MSB_V2_0.SD.n12 CM_MSB_V2_0.SD.t21 1.4602
R1230 CM_MSB_V2_0.SD.n82 CM_MSB_V2_0.SD.t52 1.46017
R1231 CM_MSB_V2_0.SD.n40 CM_MSB_V2_0.SD.t50 1.46008
R1232 CM_MSB_V2_0.SD.n68 CM_MSB_V2_0.SD.n67 1.45967
R1233 CM_MSB_V2_0.SD.n53 CM_MSB_V2_0.SD.n52 1.45927
R1234 CM_MSB_V2_0.SD.n10 CM_MSB_V2_0.SD.n9 1.45919
R1235 CM_MSB_V2_0.SD.n63 CM_MSB_V2_0.SD.n62 1.45916
R1236 CM_MSB_V2_0.SD.n108 CM_MSB_V2_0.SD.n107 1.4476
R1237 CM_MSB_V2_0.SD.n75 CM_MSB_V2_0.SD.n74 1.44746
R1238 CM_MSB_V2_0.SD.n85 CM_MSB_V2_0.SD.n84 1.44692
R1239 CM_MSB_V2_0.SD.n22 CM_MSB_V2_0.SD.n21 1.44631
R1240 CM_MSB_V2_0.SD.n43 CM_MSB_V2_0.SD.n42 1.4456
R1241 CM_MSB_V2_0.SD.n36 CM_MSB_V2_0.SD.n35 1.44501
R1242 CM_MSB_V2_0.SD.n15 CM_MSB_V2_0.SD.n14 1.44371
R1243 CM_MSB_V2_0.SD.n31 CM_MSB_V2_0.SD.n30 1.44299
R1244 CM_MSB_V2_0.SD.n94 CM_MSB_V2_0.SD.t56 1.42418
R1245 CM_MSB_V2_0.SD.n47 CM_MSB_V2_0.SD.n46 1.41105
R1246 CM_MSB_V2_0.SD.n91 CM_MSB_V2_0.SD.t6 1.3655
R1247 CM_MSB_V2_0.SD.n91 CM_MSB_V2_0.SD.n90 1.3655
R1248 CM_MSB_V2_0.SD.n89 CM_MSB_V2_0.SD.t62 1.3655
R1249 CM_MSB_V2_0.SD.n89 CM_MSB_V2_0.SD.n88 1.3655
R1250 CM_MSB_V2_0.SD.n87 CM_MSB_V2_0.SD.t1 1.3655
R1251 CM_MSB_V2_0.SD.n87 CM_MSB_V2_0.SD.n86 1.3655
R1252 CM_MSB_V2_0.SD.n107 CM_MSB_V2_0.SD.t2 1.3655
R1253 CM_MSB_V2_0.SD.n107 CM_MSB_V2_0.SD.n106 1.3655
R1254 CM_MSB_V2_0.SD.n14 CM_MSB_V2_0.SD.t40 1.3655
R1255 CM_MSB_V2_0.SD.n14 CM_MSB_V2_0.SD.n13 1.3655
R1256 CM_MSB_V2_0.SD.n21 CM_MSB_V2_0.SD.t51 1.3655
R1257 CM_MSB_V2_0.SD.n21 CM_MSB_V2_0.SD.n20 1.3655
R1258 CM_MSB_V2_0.SD.n30 CM_MSB_V2_0.SD.t36 1.3655
R1259 CM_MSB_V2_0.SD.n30 CM_MSB_V2_0.SD.n29 1.3655
R1260 CM_MSB_V2_0.SD.n35 CM_MSB_V2_0.SD.t13 1.3655
R1261 CM_MSB_V2_0.SD.n35 CM_MSB_V2_0.SD.n34 1.3655
R1262 CM_MSB_V2_0.SD.n42 CM_MSB_V2_0.SD.t28 1.3655
R1263 CM_MSB_V2_0.SD.n42 CM_MSB_V2_0.SD.n41 1.3655
R1264 CM_MSB_V2_0.SD.n45 CM_MSB_V2_0.SD.t60 1.3655
R1265 CM_MSB_V2_0.SD.n45 CM_MSB_V2_0.SD.n44 1.3655
R1266 CM_MSB_V2_0.SD.n38 CM_MSB_V2_0.SD.t24 1.3655
R1267 CM_MSB_V2_0.SD.n38 CM_MSB_V2_0.SD.n37 1.3655
R1268 CM_MSB_V2_0.SD.n28 CM_MSB_V2_0.SD.t20 1.3655
R1269 CM_MSB_V2_0.SD.n28 CM_MSB_V2_0.SD.n27 1.3655
R1270 CM_MSB_V2_0.SD.n26 CM_MSB_V2_0.SD.t33 1.3655
R1271 CM_MSB_V2_0.SD.n26 CM_MSB_V2_0.SD.n25 1.3655
R1272 CM_MSB_V2_0.SD.n19 CM_MSB_V2_0.SD.t39 1.3655
R1273 CM_MSB_V2_0.SD.n19 CM_MSB_V2_0.SD.n18 1.3655
R1274 CM_MSB_V2_0.SD.n17 CM_MSB_V2_0.SD.t10 1.3655
R1275 CM_MSB_V2_0.SD.n17 CM_MSB_V2_0.SD.n16 1.3655
R1276 CM_MSB_V2_0.SD.n78 CM_MSB_V2_0.SD.t61 1.3655
R1277 CM_MSB_V2_0.SD.n78 CM_MSB_V2_0.SD.n77 1.3655
R1278 CM_MSB_V2_0.SD.n80 CM_MSB_V2_0.SD.t18 1.3655
R1279 CM_MSB_V2_0.SD.n80 CM_MSB_V2_0.SD.n79 1.3655
R1280 CM_MSB_V2_0.SD.n84 CM_MSB_V2_0.SD.t32 1.3655
R1281 CM_MSB_V2_0.SD.n84 CM_MSB_V2_0.SD.n83 1.3655
R1282 CM_MSB_V2_0.SD.n47 CM_MSB_V2_0.SD.t7 1.28824
R1283 CM_MSB_V2_0.SD.n94 CM_MSB_V2_0.SD.n93 1.2738
R1284 CM_MSB_V2_0.SD.n75 CM_MSB_V2_0.SD.t55 1.24719
R1285 CM_MSB_V2_0.SD.n63 CM_MSB_V2_0.SD.t8 1.23341
R1286 CM_MSB_V2_0.SD.n10 CM_MSB_V2_0.SD.t54 1.23339
R1287 CM_MSB_V2_0.SD.n53 CM_MSB_V2_0.SD.t45 1.23331
R1288 CM_MSB_V2_0.SD.n68 CM_MSB_V2_0.SD.t15 1.23295
R1289 CM_MSB_V2_0.SD.n40 CM_MSB_V2_0.SD.n39 1.23247
R1290 CM_MSB_V2_0.SD.n82 CM_MSB_V2_0.SD.n81 1.23239
R1291 CM_MSB_V2_0.SD.n12 CM_MSB_V2_0.SD.n11 1.23236
R1292 CM_MSB_V2_0.SD.n24 CM_MSB_V2_0.SD.n23 1.23234
R1293 CM_MSB_V2_0.SD.n8 CM_MSB_V2_0.SD.n7 1.21851
R1294 CM_MSB_V2_0.SD.n33 CM_MSB_V2_0.SD.n32 1.21849
R1295 CM_MSB_V2_0.SD.n102 CM_MSB_V2_0.SD.n101 1.21839
R1296 CM_MSB_V2_0.SD.n69 CM_MSB_V2_0.SD.n68 1.09468
R1297 CM_MSB_V2_0.SD.n54 CM_MSB_V2_0.SD.n53 1.09004
R1298 CM_MSB_V2_0.SD.n76 CM_MSB_V2_0.SD.n75 1.08925
R1299 CM_MSB_V2_0.SD.n64 CM_MSB_V2_0.SD.n63 1.08871
R1300 CM_MSB_V2_0.SD.n95 CM_MSB_V2_0.SD.n94 1.08617
R1301 CM_MSB_V2_0.SD.n3 CM_MSB_V2_0.SD.n73 0.605393
R1302 CM_MSB_V2_0.SD.n6 CM_MSB_V2_0.SD.n92 0.603024
R1303 CM_MSB_V2_0.SD.n4 CM_MSB_V2_0.SD.n0 0.590381
R1304 CM_MSB_V2_0.SD.n1 CM_MSB_V2_0.SD.n51 0.57793
R1305 CM_MSB_V2_0.SD.n100 CM_MSB_V2_0.SD.n99 0.571801
R1306 CM_MSB_V2_0.SD.n49 CM_MSB_V2_0.SD.n48 0.571708
R1307 CM_MSB_V2_0.SD.n5 CM_MSB_V2_0.SD.n61 0.570677
R1308 CM_MSB_V2_0.SD.n72 CM_MSB_V2_0.SD.n2 0.57026
R1309 CM_MSB_V2_0.SD.n104 CM_MSB_V2_0.SD.n103 0.56537
R1310 CM_MSB_V2_0.SD.n59 CM_MSB_V2_0.SD.n58 0.560195
R1311 CM_MSB_V2_0.SD.n97 CM_MSB_V2_0.SD.n96 0.559568
R1312 CM_MSB_V2_0.SD.n56 CM_MSB_V2_0.SD.n55 0.553694
R1313 CM_MSB_V2_0.SD.n110 CM_MSB_V2_0.SD.n109 0.551536
R1314 CM_MSB_V2_0.SD.n71 CM_MSB_V2_0.SD.n70 0.54879
R1315 CM_MSB_V2_0.SD.n66 CM_MSB_V2_0.SD.n65 0.545974
R1316 CM_MSB_V2_0.SD.n2 CM_MSB_V2_0.SD.n71 0.0345612
R1317 CM_MSB_V2_0.SD.n0 CM_MSB_V2_0.SD.n66 0.034267
R1318 CM_MSB_V2_0.SD.n55 CM_MSB_V2_0.SD.n1 0.0252294
R1319 CM_MSB_V2_0.SD.n58 CM_MSB_V2_0.SD.n57 0.0202802
R1320 CM_MSB_V2_0.SD.n51 CM_MSB_V2_0.SD.n50 0.0192912
R1321 CM_MSB_V2_0.SD.n99 CM_MSB_V2_0.SD.n98 0.0192912
R1322 CM_MSB_V2_0.SD.n96 CM_MSB_V2_0.SD.n6 0.0182881
R1323 CM_MSB_V2_0.SD.n61 CM_MSB_V2_0.SD.n60 0.0181289
R1324 CM_MSB_V2_0.SD.n70 CM_MSB_V2_0.SD.n4 0.0177869
R1325 CM_MSB_V2_0.SD.n50 CM_MSB_V2_0.SD.n49 0.0164699
R1326 CM_MSB_V2_0.SD.n98 CM_MSB_V2_0.SD.n97 0.0154775
R1327 CM_MSB_V2_0.SD CM_MSB_V2_0.SD.n110 0.0153352
R1328 CM_MSB_V2_0.SD.n65 CM_MSB_V2_0.SD.n5 0.0152801
R1329 CM_MSB_V2_0.SD.n60 CM_MSB_V2_0.SD.n59 0.0149378
R1330 CM_MSB_V2_0.SD.n57 CM_MSB_V2_0.SD.n56 0.0148219
R1331 CM_MSB_V2_0.SD.n105 CM_MSB_V2_0.SD.n104 0.0148149
R1332 CM_MSB_V2_0.SD.n73 CM_MSB_V2_0.SD.n72 0.0138281
R1333 CM_MSB_V2_0.SD.n109 CM_MSB_V2_0.SD.n105 0.0138259
R1334 CM_MSB_V2_0.SD.n103 CM_MSB_V2_0.SD.n100 0.0134986
R1335 CM_MSB_V2_0.SD CM_MSB_V2_0.SD.n3 0.0123681
R1336 Local_Enc_0.Q.n55 Local_Enc_0.Q.n54 74.7525
R1337 Local_Enc_0.Q.n57 Local_Enc_0.Q.n56 74.7525
R1338 Local_Enc_0.Q.n59 Local_Enc_0.Q.n58 74.7525
R1339 Local_Enc_0.Q.n15 Local_Enc_0.Q.t35 63.1408
R1340 Local_Enc_0.Q.n61 Local_Enc_0.Q.n60 60.196
R1341 Local_Enc_0.Q.n21 Local_Enc_0.Q.n20 50.8038
R1342 Local_Enc_0.Q.n17 Local_Enc_0.Q.n16 48.5408
R1343 Local_Enc_0.Q.n19 Local_Enc_0.Q.n18 48.5408
R1344 Local_Enc_0.Q.n64 Local_Enc_0.Q.t36 28.2228
R1345 Local_Enc_0.Q.n54 Local_Enc_0.Q.t16 28.1785
R1346 Local_Enc_0.Q.n0 Local_Enc_0.Q.t14 24.4602
R1347 Local_Enc_0.Q.n38 Local_Enc_0.Q.t54 24.4602
R1348 Local_Enc_0.Q.n22 Local_Enc_0.Q.t21 24.4602
R1349 Local_Enc_0.Q.n56 Local_Enc_0.Q.n55 15.1845
R1350 Local_Enc_0.Q.n58 Local_Enc_0.Q.n57 15.1845
R1351 Local_Enc_0.Q.n60 Local_Enc_0.Q.n59 15.1845
R1352 Local_Enc_0.Q.n2 Local_Enc_0.Q.t5 14.6005
R1353 Local_Enc_0.Q.n3 Local_Enc_0.Q.t43 14.6005
R1354 Local_Enc_0.Q.n6 Local_Enc_0.Q.t20 14.6005
R1355 Local_Enc_0.Q.n7 Local_Enc_0.Q.t55 14.6005
R1356 Local_Enc_0.Q.n10 Local_Enc_0.Q.t68 14.6005
R1357 Local_Enc_0.Q.n11 Local_Enc_0.Q.t23 14.6005
R1358 Local_Enc_0.Q.n40 Local_Enc_0.Q.t47 14.6005
R1359 Local_Enc_0.Q.n41 Local_Enc_0.Q.t13 14.6005
R1360 Local_Enc_0.Q.n44 Local_Enc_0.Q.t57 14.6005
R1361 Local_Enc_0.Q.n45 Local_Enc_0.Q.t25 14.6005
R1362 Local_Enc_0.Q.n48 Local_Enc_0.Q.t45 14.6005
R1363 Local_Enc_0.Q.n49 Local_Enc_0.Q.t60 14.6005
R1364 Local_Enc_0.Q.n24 Local_Enc_0.Q.t18 14.6005
R1365 Local_Enc_0.Q.n25 Local_Enc_0.Q.t53 14.6005
R1366 Local_Enc_0.Q.n28 Local_Enc_0.Q.t29 14.6005
R1367 Local_Enc_0.Q.n29 Local_Enc_0.Q.t63 14.6005
R1368 Local_Enc_0.Q.n32 Local_Enc_0.Q.t15 14.6005
R1369 Local_Enc_0.Q.n33 Local_Enc_0.Q.t33 14.6005
R1370 Local_Enc_0.Q.n15 Local_Enc_0.Q.t32 14.6005
R1371 Local_Enc_0.Q.n16 Local_Enc_0.Q.t65 14.6005
R1372 Local_Enc_0.Q.n17 Local_Enc_0.Q.t44 14.6005
R1373 Local_Enc_0.Q.n18 Local_Enc_0.Q.t7 14.6005
R1374 Local_Enc_0.Q.n19 Local_Enc_0.Q.t28 14.6005
R1375 Local_Enc_0.Q.n20 Local_Enc_0.Q.t48 14.6005
R1376 Local_Enc_0.Q.n64 Local_Enc_0.Q.t37 14.4701
R1377 Local_Enc_0.Q.n0 Local_Enc_0.Q.t31 14.0165
R1378 Local_Enc_0.Q.n1 Local_Enc_0.Q.t24 14.0165
R1379 Local_Enc_0.Q.n4 Local_Enc_0.Q.t42 14.0165
R1380 Local_Enc_0.Q.n5 Local_Enc_0.Q.t6 14.0165
R1381 Local_Enc_0.Q.n8 Local_Enc_0.Q.t67 14.0165
R1382 Local_Enc_0.Q.n9 Local_Enc_0.Q.t22 14.0165
R1383 Local_Enc_0.Q.n12 Local_Enc_0.Q.t39 14.0165
R1384 Local_Enc_0.Q.n13 Local_Enc_0.Q.t4 14.0165
R1385 Local_Enc_0.Q.n38 Local_Enc_0.Q.t66 14.0165
R1386 Local_Enc_0.Q.n39 Local_Enc_0.Q.t61 14.0165
R1387 Local_Enc_0.Q.n42 Local_Enc_0.Q.t12 14.0165
R1388 Local_Enc_0.Q.n43 Local_Enc_0.Q.t49 14.0165
R1389 Local_Enc_0.Q.n46 Local_Enc_0.Q.t41 14.0165
R1390 Local_Enc_0.Q.n47 Local_Enc_0.Q.t58 14.0165
R1391 Local_Enc_0.Q.n50 Local_Enc_0.Q.t9 14.0165
R1392 Local_Enc_0.Q.n51 Local_Enc_0.Q.t46 14.0165
R1393 Local_Enc_0.Q.n22 Local_Enc_0.Q.t38 14.0165
R1394 Local_Enc_0.Q.n23 Local_Enc_0.Q.t34 14.0165
R1395 Local_Enc_0.Q.n26 Local_Enc_0.Q.t52 14.0165
R1396 Local_Enc_0.Q.n27 Local_Enc_0.Q.t19 14.0165
R1397 Local_Enc_0.Q.n30 Local_Enc_0.Q.t11 14.0165
R1398 Local_Enc_0.Q.n31 Local_Enc_0.Q.t30 14.0165
R1399 Local_Enc_0.Q.n34 Local_Enc_0.Q.t50 14.0165
R1400 Local_Enc_0.Q.n35 Local_Enc_0.Q.t17 14.0165
R1401 Local_Enc_0.Q.n54 Local_Enc_0.Q.t8 12.9945
R1402 Local_Enc_0.Q.n55 Local_Enc_0.Q.t27 12.9945
R1403 Local_Enc_0.Q.n56 Local_Enc_0.Q.t62 12.9945
R1404 Local_Enc_0.Q.n57 Local_Enc_0.Q.t56 12.9945
R1405 Local_Enc_0.Q.n58 Local_Enc_0.Q.t3 12.9945
R1406 Local_Enc_0.Q.n59 Local_Enc_0.Q.t26 12.9945
R1407 Local_Enc_0.Q.n60 Local_Enc_0.Q.t59 12.9945
R1408 Local_Enc_0.Q.n14 Local_Enc_0.Q.t40 12.3375
R1409 Local_Enc_0.Q.n52 Local_Enc_0.Q.t10 12.3375
R1410 Local_Enc_0.Q.n36 Local_Enc_0.Q.t51 12.3375
R1411 Local_Enc_0.Q.n21 Local_Enc_0.Q.t64 12.3375
R1412 Local_Enc_0.Q.n14 Local_Enc_0.Q.n13 12.1232
R1413 Local_Enc_0.Q.n52 Local_Enc_0.Q.n51 12.1232
R1414 Local_Enc_0.Q.n36 Local_Enc_0.Q.n35 12.1232
R1415 Local_Enc_0.Q.n1 Local_Enc_0.Q.n0 9.86024
R1416 Local_Enc_0.Q.n2 Local_Enc_0.Q.n1 9.86024
R1417 Local_Enc_0.Q.n3 Local_Enc_0.Q.n2 9.86024
R1418 Local_Enc_0.Q.n4 Local_Enc_0.Q.n3 9.86024
R1419 Local_Enc_0.Q.n5 Local_Enc_0.Q.n4 9.86024
R1420 Local_Enc_0.Q.n6 Local_Enc_0.Q.n5 9.86024
R1421 Local_Enc_0.Q.n7 Local_Enc_0.Q.n6 9.86024
R1422 Local_Enc_0.Q.n8 Local_Enc_0.Q.n7 9.86024
R1423 Local_Enc_0.Q.n9 Local_Enc_0.Q.n8 9.86024
R1424 Local_Enc_0.Q.n10 Local_Enc_0.Q.n9 9.86024
R1425 Local_Enc_0.Q.n11 Local_Enc_0.Q.n10 9.86024
R1426 Local_Enc_0.Q.n12 Local_Enc_0.Q.n11 9.86024
R1427 Local_Enc_0.Q.n13 Local_Enc_0.Q.n12 9.86024
R1428 Local_Enc_0.Q.n39 Local_Enc_0.Q.n38 9.86024
R1429 Local_Enc_0.Q.n40 Local_Enc_0.Q.n39 9.86024
R1430 Local_Enc_0.Q.n41 Local_Enc_0.Q.n40 9.86024
R1431 Local_Enc_0.Q.n42 Local_Enc_0.Q.n41 9.86024
R1432 Local_Enc_0.Q.n43 Local_Enc_0.Q.n42 9.86024
R1433 Local_Enc_0.Q.n44 Local_Enc_0.Q.n43 9.86024
R1434 Local_Enc_0.Q.n45 Local_Enc_0.Q.n44 9.86024
R1435 Local_Enc_0.Q.n46 Local_Enc_0.Q.n45 9.86024
R1436 Local_Enc_0.Q.n47 Local_Enc_0.Q.n46 9.86024
R1437 Local_Enc_0.Q.n48 Local_Enc_0.Q.n47 9.86024
R1438 Local_Enc_0.Q.n49 Local_Enc_0.Q.n48 9.86024
R1439 Local_Enc_0.Q.n50 Local_Enc_0.Q.n49 9.86024
R1440 Local_Enc_0.Q.n51 Local_Enc_0.Q.n50 9.86024
R1441 Local_Enc_0.Q.n23 Local_Enc_0.Q.n22 9.86024
R1442 Local_Enc_0.Q.n24 Local_Enc_0.Q.n23 9.86024
R1443 Local_Enc_0.Q.n25 Local_Enc_0.Q.n24 9.86024
R1444 Local_Enc_0.Q.n26 Local_Enc_0.Q.n25 9.86024
R1445 Local_Enc_0.Q.n27 Local_Enc_0.Q.n26 9.86024
R1446 Local_Enc_0.Q.n28 Local_Enc_0.Q.n27 9.86024
R1447 Local_Enc_0.Q.n29 Local_Enc_0.Q.n28 9.86024
R1448 Local_Enc_0.Q.n30 Local_Enc_0.Q.n29 9.86024
R1449 Local_Enc_0.Q.n31 Local_Enc_0.Q.n30 9.86024
R1450 Local_Enc_0.Q.n32 Local_Enc_0.Q.n31 9.86024
R1451 Local_Enc_0.Q.n33 Local_Enc_0.Q.n32 9.86024
R1452 Local_Enc_0.Q.n34 Local_Enc_0.Q.n33 9.86024
R1453 Local_Enc_0.Q.n35 Local_Enc_0.Q.n34 9.86024
R1454 Local_Enc_0.Q.n16 Local_Enc_0.Q.n15 9.86024
R1455 Local_Enc_0.Q.n18 Local_Enc_0.Q.n17 9.86024
R1456 Local_Enc_0.Q.n20 Local_Enc_0.Q.n19 9.86024
R1457 Local_Enc_0.Q.n37 Local_Enc_0.Q.n21 9.72687
R1458 Local_Enc_0.Q.n53 Local_Enc_0.Q.n52 8.44029
R1459 Local_Enc_0.Q.n37 Local_Enc_0.Q.n36 8.44029
R1460 Local_Enc_0.Q Local_Enc_0.Q.n63 6.8765
R1461 Local_Enc_0.Q.n62 Local_Enc_0.Q.n14 6.14729
R1462 Local_Enc_0.Q.n67 Local_Enc_0.Q 6.04981
R1463 Local_Enc_0.Q Local_Enc_0.Q.n62 5.90026
R1464 Local_Enc_0.Q Local_Enc_0.Q.n64 4.53357
R1465 Local_Enc_0.Q.n66 Local_Enc_0.Q.t1 3.6405
R1466 Local_Enc_0.Q.n66 Local_Enc_0.Q.n65 3.6405
R1467 Local_Enc_0.Q.n67 Local_Enc_0.Q.n66 2.6005
R1468 Local_Enc_0.Q.n62 Local_Enc_0.Q.n61 2.2505
R1469 Local_Enc_0.Q.n53 Local_Enc_0.Q.n37 1.24534
R1470 Local_Enc_0.Q.n61 Local_Enc_0.Q.n53 1.24509
R1471 Local_Enc_0.Q Local_Enc_0.Q.n67 0.818982
R1472 IOUT+.n38 IOUT+.t17 9.53443
R1473 IOUT+.n61 IOUT+.t56 9.53443
R1474 IOUT+.n84 IOUT+.t28 9.53443
R1475 IOUT+.n14 IOUT+.t4 9.53443
R1476 IOUT+.n46 IOUT+.n24 6.13289
R1477 IOUT+.n92 IOUT+.n70 6.13289
R1478 IOUT+.n69 IOUT+.n47 6.08789
R1479 IOUT+.n22 IOUT+.n0 6.08789
R1480 IOUT+.n43 IOUT+.n42 5.91472
R1481 IOUT+.n66 IOUT+.n65 5.91472
R1482 IOUT+.n89 IOUT+.n88 5.91472
R1483 IOUT+.n19 IOUT+.n18 5.91472
R1484 IOUT+.n39 IOUT+.n32 5.84965
R1485 IOUT+.n62 IOUT+.n55 5.84965
R1486 IOUT+.n85 IOUT+.n78 5.84965
R1487 IOUT+.n15 IOUT+.n8 5.84965
R1488 IOUT+.n40 IOUT+.n30 5.54055
R1489 IOUT+.n63 IOUT+.n53 5.54055
R1490 IOUT+.n86 IOUT+.n76 5.54055
R1491 IOUT+.n16 IOUT+.n6 5.54055
R1492 IOUT+.n37 IOUT+.n36 4.38877
R1493 IOUT+.n60 IOUT+.n59 4.38877
R1494 IOUT+.n83 IOUT+.n82 4.38877
R1495 IOUT+.n13 IOUT+.n12 4.38877
R1496 IOUT+.n93 IOUT+.n92 4.07638
R1497 IOUT+.n45 IOUT+.n26 3.64354
R1498 IOUT+.n68 IOUT+.n49 3.64354
R1499 IOUT+.n91 IOUT+.n72 3.64354
R1500 IOUT+.n21 IOUT+.n2 3.64354
R1501 IOUT+.n44 IOUT+.n28 3.29178
R1502 IOUT+.n67 IOUT+.n51 3.29178
R1503 IOUT+.n90 IOUT+.n74 3.29178
R1504 IOUT+.n20 IOUT+.n4 3.29178
R1505 IOUT+.n37 IOUT+.n34 3.29055
R1506 IOUT+.n60 IOUT+.n57 3.29055
R1507 IOUT+.n83 IOUT+.n80 3.29055
R1508 IOUT+.n13 IOUT+.n10 3.29055
R1509 IOUT+.n44 IOUT+.n43 3.08985
R1510 IOUT+.n67 IOUT+.n66 3.08985
R1511 IOUT+.n90 IOUT+.n89 3.08985
R1512 IOUT+.n20 IOUT+.n19 3.08985
R1513 IOUT+.n93 IOUT+.n69 2.87254
R1514 IOUT+.n94 IOUT+.n46 2.83004
R1515 IOUT+.n42 IOUT+.t54 2.7305
R1516 IOUT+.n42 IOUT+.n41 2.7305
R1517 IOUT+.n30 IOUT+.t37 2.7305
R1518 IOUT+.n30 IOUT+.n29 2.7305
R1519 IOUT+.n32 IOUT+.t27 2.7305
R1520 IOUT+.n32 IOUT+.n31 2.7305
R1521 IOUT+.n34 IOUT+.t51 2.7305
R1522 IOUT+.n34 IOUT+.n33 2.7305
R1523 IOUT+.n36 IOUT+.t57 2.7305
R1524 IOUT+.n36 IOUT+.n35 2.7305
R1525 IOUT+.n28 IOUT+.t48 2.7305
R1526 IOUT+.n28 IOUT+.n27 2.7305
R1527 IOUT+.n26 IOUT+.t2 2.7305
R1528 IOUT+.n26 IOUT+.n25 2.7305
R1529 IOUT+.n65 IOUT+.t26 2.7305
R1530 IOUT+.n65 IOUT+.n64 2.7305
R1531 IOUT+.n53 IOUT+.t11 2.7305
R1532 IOUT+.n53 IOUT+.n52 2.7305
R1533 IOUT+.n55 IOUT+.t1 2.7305
R1534 IOUT+.n55 IOUT+.n54 2.7305
R1535 IOUT+.n57 IOUT+.t23 2.7305
R1536 IOUT+.n57 IOUT+.n56 2.7305
R1537 IOUT+.n59 IOUT+.t29 2.7305
R1538 IOUT+.n59 IOUT+.n58 2.7305
R1539 IOUT+.n51 IOUT+.t21 2.7305
R1540 IOUT+.n51 IOUT+.n50 2.7305
R1541 IOUT+.n49 IOUT+.t35 2.7305
R1542 IOUT+.n49 IOUT+.n48 2.7305
R1543 IOUT+.n88 IOUT+.t39 2.7305
R1544 IOUT+.n88 IOUT+.n87 2.7305
R1545 IOUT+.n76 IOUT+.t46 2.7305
R1546 IOUT+.n76 IOUT+.n75 2.7305
R1547 IOUT+.n78 IOUT+.t12 2.7305
R1548 IOUT+.n78 IOUT+.n77 2.7305
R1549 IOUT+.n80 IOUT+.t0 2.7305
R1550 IOUT+.n80 IOUT+.n79 2.7305
R1551 IOUT+.n82 IOUT+.t40 2.7305
R1552 IOUT+.n82 IOUT+.n81 2.7305
R1553 IOUT+.n74 IOUT+.t61 2.7305
R1554 IOUT+.n74 IOUT+.n73 2.7305
R1555 IOUT+.n72 IOUT+.t50 2.7305
R1556 IOUT+.n72 IOUT+.n71 2.7305
R1557 IOUT+.n18 IOUT+.t16 2.7305
R1558 IOUT+.n18 IOUT+.n17 2.7305
R1559 IOUT+.n6 IOUT+.t24 2.7305
R1560 IOUT+.n6 IOUT+.n5 2.7305
R1561 IOUT+.n8 IOUT+.t55 2.7305
R1562 IOUT+.n8 IOUT+.n7 2.7305
R1563 IOUT+.n10 IOUT+.t38 2.7305
R1564 IOUT+.n10 IOUT+.n9 2.7305
R1565 IOUT+.n12 IOUT+.t18 2.7305
R1566 IOUT+.n12 IOUT+.n11 2.7305
R1567 IOUT+.n4 IOUT+.t34 2.7305
R1568 IOUT+.n4 IOUT+.n3 2.7305
R1569 IOUT+.n2 IOUT+.t30 2.7305
R1570 IOUT+.n2 IOUT+.n1 2.7305
R1571 IOUT+ IOUT+.n23 2.25862
R1572 IOUT+.n38 IOUT+.n37 2.2505
R1573 IOUT+.n61 IOUT+.n60 2.2505
R1574 IOUT+.n84 IOUT+.n83 2.2505
R1575 IOUT+.n14 IOUT+.n13 2.2505
R1576 IOUT+ IOUT+.n94 1.24572
R1577 IOUT+.n94 IOUT+.n93 1.24325
R1578 IOUT+.n69 IOUT+.n68 0.797345
R1579 IOUT+.n22 IOUT+.n21 0.797304
R1580 IOUT+.n45 IOUT+.n44 0.76828
R1581 IOUT+.n68 IOUT+.n67 0.76828
R1582 IOUT+.n91 IOUT+.n90 0.76828
R1583 IOUT+.n21 IOUT+.n20 0.76828
R1584 IOUT+.n46 IOUT+.n45 0.755717
R1585 IOUT+.n92 IOUT+.n91 0.755717
R1586 IOUT+.n23 IOUT+.n22 0.618164
R1587 IOUT+.n39 IOUT+.n38 0.60021
R1588 IOUT+.n62 IOUT+.n61 0.60021
R1589 IOUT+.n85 IOUT+.n84 0.60021
R1590 IOUT+.n15 IOUT+.n14 0.60021
R1591 IOUT+.n40 IOUT+.n39 0.59455
R1592 IOUT+.n63 IOUT+.n62 0.59455
R1593 IOUT+.n86 IOUT+.n85 0.59455
R1594 IOUT+.n16 IOUT+.n15 0.59455
R1595 IOUT+.n43 IOUT+.n40 0.58347
R1596 IOUT+.n66 IOUT+.n63 0.58347
R1597 IOUT+.n89 IOUT+.n86 0.58347
R1598 IOUT+.n19 IOUT+.n16 0.58347
R1599 IM IM.n30 32.397
R1600 IM.n0 IM.t8 30.5343
R1601 IM.n0 IM.t4 18.1775
R1602 IM.n1 IM.t16 18.1775
R1603 IM.n4 IM.t12 18.1775
R1604 IM.n5 IM.t28 18.1775
R1605 IM.n8 IM.t25 18.1775
R1606 IM.n9 IM.t1 18.1775
R1607 IM.n12 IM.t11 18.1775
R1608 IM.n13 IM.t27 18.1775
R1609 IM.n16 IM.t29 18.1775
R1610 IM.n17 IM.t19 18.1775
R1611 IM.n20 IM.t18 18.1775
R1612 IM.n21 IM.t9 18.1775
R1613 IM.n24 IM.t26 18.1775
R1614 IM.n25 IM.t10 18.1775
R1615 IM.n28 IM.t13 18.1775
R1616 IM.n29 IM.t2 18.1775
R1617 IM.n2 IM.t5 17.6665
R1618 IM.n3 IM.t23 17.6665
R1619 IM.n6 IM.t24 17.6665
R1620 IM.n7 IM.t30 17.6665
R1621 IM.n10 IM.t3 17.6665
R1622 IM.n11 IM.t14 17.6665
R1623 IM.n14 IM.t22 17.6665
R1624 IM.n15 IM.t6 17.6665
R1625 IM.n18 IM.t31 17.6665
R1626 IM.n19 IM.t20 17.6665
R1627 IM.n22 IM.t15 17.6665
R1628 IM.n23 IM.t0 17.6665
R1629 IM.n26 IM.t21 17.6665
R1630 IM.n27 IM.t17 17.6665
R1631 IM.n30 IM.t7 17.6665
R1632 IM.n1 IM.n0 12.8683
R1633 IM.n2 IM.n1 12.8683
R1634 IM.n3 IM.n2 12.8683
R1635 IM.n4 IM.n3 12.8683
R1636 IM.n5 IM.n4 12.8683
R1637 IM.n6 IM.n5 12.8683
R1638 IM.n7 IM.n6 12.8683
R1639 IM.n8 IM.n7 12.8683
R1640 IM.n9 IM.n8 12.8683
R1641 IM.n10 IM.n9 12.8683
R1642 IM.n11 IM.n10 12.8683
R1643 IM.n12 IM.n11 12.8683
R1644 IM.n13 IM.n12 12.8683
R1645 IM.n14 IM.n13 12.8683
R1646 IM.n15 IM.n14 12.8683
R1647 IM.n16 IM.n15 12.8683
R1648 IM.n17 IM.n16 12.8683
R1649 IM.n18 IM.n17 12.8683
R1650 IM.n19 IM.n18 12.8683
R1651 IM.n20 IM.n19 12.8683
R1652 IM.n21 IM.n20 12.8683
R1653 IM.n22 IM.n21 12.8683
R1654 IM.n23 IM.n22 12.8683
R1655 IM.n24 IM.n23 12.8683
R1656 IM.n25 IM.n24 12.8683
R1657 IM.n26 IM.n25 12.8683
R1658 IM.n27 IM.n26 12.8683
R1659 IM.n28 IM.n27 12.8683
R1660 IM.n29 IM.n28 12.8683
R1661 IM.n30 IM.n29 12.8683
R1662 VDD.n24 VDD.t28 178.431
R1663 VDD.n20 VDD.t11 178.431
R1664 VDD.n16 VDD.t3 178.431
R1665 VDD.n38 VDD.t37 178.431
R1666 VDD.n34 VDD.t21 178.431
R1667 VDD.n30 VDD.t8 178.431
R1668 VDD.n11 VDD.t0 178.431
R1669 VDD.n7 VDD.t14 178.431
R1670 VDD.n3 VDD.t42 178.431
R1671 VDD.n24 VDD.t19 135.294
R1672 VDD.n20 VDD.t35 135.294
R1673 VDD.n16 VDD.t31 135.294
R1674 VDD.n38 VDD.t40 135.294
R1675 VDD.n34 VDD.t26 135.294
R1676 VDD.n30 VDD.t6 135.294
R1677 VDD.n11 VDD.t24 135.294
R1678 VDD.n7 VDD.t17 135.294
R1679 VDD.n3 VDD.t33 135.294
R1680 VDD.n17 VDD.n15 6.69527
R1681 VDD.n31 VDD.n29 6.69527
R1682 VDD.n4 VDD.n2 6.69527
R1683 VDD.n19 VDD.n14 6.59267
R1684 VDD.n23 VDD.n13 6.59267
R1685 VDD.n33 VDD.n28 6.59267
R1686 VDD.n37 VDD.n27 6.59267
R1687 VDD.n6 VDD.n1 6.59267
R1688 VDD.n10 VDD.n0 6.59267
R1689 VDD.n18 VDD.t32 6.55815
R1690 VDD.n22 VDD.t36 6.55815
R1691 VDD.n26 VDD.t20 6.55815
R1692 VDD.n32 VDD.t7 6.55815
R1693 VDD.n36 VDD.t27 6.55815
R1694 VDD.n40 VDD.t41 6.55815
R1695 VDD.n5 VDD.t34 6.55815
R1696 VDD.n9 VDD.t18 6.55815
R1697 VDD.n42 VDD.t25 6.55815
R1698 VDD.n17 VDD.n16 6.3005
R1699 VDD.n21 VDD.n20 6.3005
R1700 VDD.n25 VDD.n24 6.3005
R1701 VDD.n31 VDD.n30 6.3005
R1702 VDD.n35 VDD.n34 6.3005
R1703 VDD.n39 VDD.n38 6.3005
R1704 VDD.n4 VDD.n3 6.3005
R1705 VDD.n8 VDD.n7 6.3005
R1706 VDD.n12 VDD.n11 6.3005
R1707 VDD.n41 VDD.n40 3.87957
R1708 VDD VDD.n41 3.85281
R1709 VDD.n41 VDD.n26 2.58214
R1710 VDD.n19 VDD.n18 0.339604
R1711 VDD.n33 VDD.n32 0.339604
R1712 VDD.n6 VDD.n5 0.339604
R1713 VDD.n23 VDD.n22 0.302039
R1714 VDD.n37 VDD.n36 0.302039
R1715 VDD.n10 VDD.n9 0.302039
R1716 VDD.n21 VDD.n19 0.1031
R1717 VDD.n25 VDD.n23 0.1031
R1718 VDD.n35 VDD.n33 0.1031
R1719 VDD.n39 VDD.n37 0.1031
R1720 VDD.n8 VDD.n6 0.1031
R1721 VDD.n12 VDD.n10 0.1031
R1722 VDD.n42 VDD 0.0996385
R1723 VDD.n18 VDD 0.0893
R1724 VDD.n22 VDD 0.0893
R1725 VDD.n26 VDD 0.0893
R1726 VDD.n32 VDD 0.0893
R1727 VDD.n36 VDD 0.0893
R1728 VDD.n40 VDD 0.0893
R1729 VDD.n5 VDD 0.0893
R1730 VDD VDD.n42 0.0893
R1731 VDD.n9 VDD 0.0839
R1732 VDD VDD.n17 0.0017
R1733 VDD VDD.n21 0.0017
R1734 VDD VDD.n25 0.0017
R1735 VDD VDD.n31 0.0017
R1736 VDD VDD.n35 0.0017
R1737 VDD VDD.n39 0.0017
R1738 VDD VDD.n4 0.0017
R1739 VDD VDD.n8 0.0017
R1740 VDD VDD.n12 0.0017
R1741 Ci.n1 Ci.t1 28.2228
R1742 Ci.n0 Ci.t2 26.9784
R1743 Ci.n0 Ci.t0 14.7248
R1744 Ci.n1 Ci.t3 14.4701
R1745 Ci Ci.n1 4.53357
R1746 Ci.n3 Ci.n0 4.15413
R1747 Ci.n2 Ci 0.0963696
R1748 Ci.n2 Ci 0.0728913
R1749 Ci.n3 Ci.n2 0.00441304
R1750 Ci Ci.n3 0.00245652
R1751 Ri.n1 Ri.t1 28.2228
R1752 Ri.n0 Ri.t2 26.9784
R1753 Ri.n0 Ri.t0 14.7248
R1754 Ri.n1 Ri.t3 14.4701
R1755 Ri Ri.n1 4.53357
R1756 Ri Ri.n0 4.18544
R1757 Ri-1.n1 Ri-1.t2 28.2228
R1758 Ri-1.n0 Ri-1.t1 26.9784
R1759 Ri-1.n0 Ri-1.t0 14.7248
R1760 Ri-1.n1 Ri-1.t3 14.4701
R1761 Ri-1.n2 Ri-1.n1 4.50813
R1762 Ri-1 Ri-1.n0 4.18544
R1763 Ri-1.n3 Ri-1 0.086587
R1764 Ri-1.n3 Ri-1.n2 0.0787609
R1765 Ri-1 Ri-1.n3 0.0200652
R1766 Ri-1.n2 Ri-1 0.00636957
C0 Local_Enc_0.NAND_6.A Ci 1.17e-19
C1 Local_Enc_0.NAND_6.A VDD 0.358f
C2 Local_Enc_0.NAND_6.A Local_Enc_0.NAND_6.B 0.429f
C3 CM_MSB_V2_0.SD IOUT+ 0.00427f
C4 IM_T Local_Enc_0.NAND_6.A 0.00339f
C5 IOUT+ CM_MSB_V2_0.OUT 7.37f
C6 Local_Enc_0.NAND_5.B Local_Enc_0.QB 0.00682f
C7 CM_MSB_V2_0.SD CM_MSB_V2_0.OUT 4.67f
C8 VDD Local_Enc_0.NAND_1.B 0.628f
C9 Local_Enc_0.NAND_1.B Local_Enc_0.NAND_6.B 1.35e-19
C10 a_n1846_3765# Local_Enc_0.NAND_6.A 0.0812f
C11 Local_Enc_0.Q Local_Enc_0.NAND_1.B 0.004f
C12 Local_Enc_0.NAND_5.B a_n1846_4741# 0.0043f
C13 Local_Enc_0.NAND_5.B Ri-1 0.00973f
C14 Ri Local_Enc_0.NAND_6.A 0.233f
C15 Ci Local_Enc_0.NAND_8.A 8.53e-19
C16 VDD Local_Enc_0.NAND_8.A 0.864f
C17 Local_Enc_0.NAND_8.A Local_Enc_0.NAND_6.B 0.00405f
C18 Local_Enc_0.NAND_4.B a_n1035_5712# 0.00495f
C19 IM_T Local_Enc_0.NAND_8.A 0.0073f
C20 Local_Enc_0.QB Local_Enc_0.NAND_1.B 1.31e-19
C21 Local_Enc_0.Q Local_Enc_0.NAND_8.A 0.208f
C22 a_n1846_4741# Local_Enc_0.NAND_6.A 5.69e-20
C23 a_n1035_3765# Local_Enc_0.NAND_8.A 0.0852f
C24 Local_Enc_0.NAND_6.A CM_MSB_V2_0.SD 0.00198f
C25 Ri-1 Local_Enc_0.NAND_1.B 0.24f
C26 Local_Enc_0.QB Local_Enc_0.NAND_8.A 0.43f
C27 Ri Local_Enc_0.NAND_8.A 5.21e-19
C28 IM Local_Enc_0.NAND_8.A 3.24e-19
C29 a_n1035_4741# Local_Enc_0.NAND_8.A 0.0821f
C30 IOUT+ Local_Enc_0.NAND_8.A 7.56e-20
C31 a_n1846_4741# Local_Enc_0.NAND_8.A 0.045f
C32 CM_MSB_V2_0.SD Local_Enc_0.NAND_8.A 0.00473f
C33 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_1.B 0.344f
C34 CM_MSB_V2_0.OUT Local_Enc_0.NAND_8.A 1.41e-19
C35 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_5.A 0.00496f
C36 a_n1846_5712# Local_Enc_0.NAND_5.A 5.76e-20
C37 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_8.A 0.0646f
C38 Local_Enc_0.NAND_6.A Local_Enc_0.NAND_8.A 0.0124f
C39 IM_T IOUT- 0.0211f
C40 Local_Enc_0.NAND_4.B VDD 0.673f
C41 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_6.B 2.09e-20
C42 Local_Enc_0.NAND_1.B Local_Enc_0.NAND_8.A 1.18e-19
C43 IOUT- Local_Enc_0.Q 1.18f
C44 Local_Enc_0.NAND_4.B IM_T 0.00103f
C45 Local_Enc_0.NAND_4.B Local_Enc_0.Q 0.686f
C46 Local_Enc_0.NAND_4.B a_n1035_3765# 0.0419f
C47 a_n1035_5712# Local_Enc_0.Q 0.0961f
C48 a_n2609_5712# Ci 5.76e-20
C49 a_n2609_5712# VDD 8.42e-19
C50 IOUT- Local_Enc_0.QB 1.68f
C51 a_n1846_5712# Local_Enc_0.Q 6.06e-19
C52 IM IOUT- 0.0126f
C53 Local_Enc_0.NAND_4.B Local_Enc_0.QB 0.495f
C54 Local_Enc_0.NAND_4.B Ri 2.34e-22
C55 a_n1035_5712# Local_Enc_0.QB 0.0423f
C56 Local_Enc_0.NAND_4.B IM 1.99e-19
C57 IOUT+ IOUT- 7.98f
C58 Local_Enc_0.NAND_4.B a_n1035_4741# 0.00331f
C59 Local_Enc_0.NAND_4.B Ri-1 1.08e-19
C60 CM_MSB_V2_0.SD IOUT- 0.0307f
C61 IOUT- CM_MSB_V2_0.OUT 8.39f
C62 Local_Enc_0.NAND_4.B CM_MSB_V2_0.SD 0.00299f
C63 Local_Enc_0.NAND_4.B CM_MSB_V2_0.OUT 2.29e-19
C64 Ci Local_Enc_0.NAND_5.A 0.00321f
C65 VDD Local_Enc_0.NAND_5.A 0.503f
C66 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_6.B 0.232f
C67 IM_T Local_Enc_0.NAND_5.A 0.00438f
C68 a_n2609_5712# Ri-1 0.0852f
C69 Local_Enc_0.Q Local_Enc_0.NAND_5.A 2.28e-19
C70 a_n1035_3765# Local_Enc_0.NAND_5.A 1.88e-20
C71 a_n2609_4741# Local_Enc_0.NAND_5.A 2.15e-19
C72 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_5.B 0.026f
C73 a_n1846_3765# Local_Enc_0.NAND_5.A 0.0451f
C74 Local_Enc_0.NAND_5.B a_n1035_5712# 6.99e-20
C75 Local_Enc_0.QB Local_Enc_0.NAND_5.A 0.00927f
C76 Local_Enc_0.NAND_5.B a_n1846_5712# 0.0469f
C77 Ri Local_Enc_0.NAND_5.A 9.03e-19
C78 IM Local_Enc_0.NAND_5.A 0.00213f
C79 Local_Enc_0.NAND_5.B a_n2609_5712# 0.00175f
C80 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_6.A 1.31e-19
C81 a_n2609_3766# IM_T 2.11e-19
C82 a_n1846_4741# Local_Enc_0.NAND_5.A 0.0874f
C83 VDD Ci 0.378f
C84 Ci Local_Enc_0.NAND_6.B 0.235f
C85 CM_MSB_V2_0.SD Local_Enc_0.NAND_5.A 0.0153f
C86 CM_MSB_V2_0.OUT Local_Enc_0.NAND_5.A 0.00106f
C87 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_1.B 0.00819f
C88 VDD Local_Enc_0.NAND_6.B 0.618f
C89 IM_T VDD 0.0096f
C90 IM_T Local_Enc_0.NAND_6.B 0.00448f
C91 VDD Local_Enc_0.Q 0.588f
C92 a_n1846_5712# Local_Enc_0.NAND_1.B 0.0852f
C93 a_n2609_4741# Ci 0.0852f
C94 IM_T Local_Enc_0.Q 0.0573f
C95 IOUT- Local_Enc_0.NAND_8.A 1.62e-19
C96 a_n2609_4741# Local_Enc_0.NAND_6.B 0.0444f
C97 a_n1035_3765# IM_T 2.11e-19
C98 IM_T a_n2609_4741# 1.47e-20
C99 a_n2609_3766# Ri 0.0852f
C100 a_n1846_3765# Local_Enc_0.NAND_6.B 0.00403f
C101 a_n2609_5712# Local_Enc_0.NAND_1.B 0.0419f
C102 Local_Enc_0.NAND_4.B Local_Enc_0.NAND_8.A 0.345f
C103 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_5.A 0.316f
C104 a_n1035_3765# Local_Enc_0.Q 1.23e-19
C105 a_n1846_3765# IM_T 2.11e-19
C106 Local_Enc_0.QB Ci 5.92e-19
C107 a_n1035_5712# Local_Enc_0.NAND_8.A 5.76e-20
C108 VDD Local_Enc_0.QB 0.639f
C109 Local_Enc_0.QB Local_Enc_0.NAND_6.B 4.6e-19
C110 Ri Ci 0.00475f
C111 IM_T Local_Enc_0.QB 0.00321f
C112 Ri VDD 0.364f
C113 Ri Local_Enc_0.NAND_6.B 0.0132f
C114 IM Local_Enc_0.NAND_6.B 0.00136f
C115 IM_T Ri 0.00518f
C116 Local_Enc_0.Q Local_Enc_0.QB 5.71f
C117 IM_T IM 1.99f
C118 a_n1035_3765# Local_Enc_0.QB 3.34e-19
C119 a_n2609_3766# CM_MSB_V2_0.SD 4.2e-19
C120 Local_Enc_0.NAND_6.A Local_Enc_0.NAND_5.A 0.216f
C121 IM Local_Enc_0.Q 7.41e-19
C122 IM_T a_n1035_4741# 1.47e-20
C123 a_n1035_3765# Ri 3.42e-22
C124 Ri-1 Ci 0.00479f
C125 VDD Ri-1 0.389f
C126 a_n2609_4741# Ri 5.71e-20
C127 a_n1846_4741# Local_Enc_0.NAND_6.B 2.79e-20
C128 Ri-1 Local_Enc_0.NAND_6.B 1.18e-19
C129 a_n1035_4741# Local_Enc_0.Q 0.043f
C130 IM_T IOUT+ 0.00188f
C131 IM_T a_n1846_4741# 1.47e-20
C132 a_n1846_3765# Ri 1.61e-21
C133 CM_MSB_V2_0.SD VDD 0.00235f
C134 CM_MSB_V2_0.SD Local_Enc_0.NAND_6.B 0.00526f
C135 CM_MSB_V2_0.OUT Local_Enc_0.NAND_6.B 1.93e-19
C136 IOUT+ Local_Enc_0.Q 1.2f
C137 Local_Enc_0.NAND_1.B Local_Enc_0.NAND_5.A 0.00251f
C138 IM_T CM_MSB_V2_0.SD 1f
C139 IM_T CM_MSB_V2_0.OUT 0.762f
C140 IM Local_Enc_0.QB 7.5e-19
C141 CM_MSB_V2_0.SD Local_Enc_0.Q 0.00613f
C142 Local_Enc_0.Q CM_MSB_V2_0.OUT 4.21f
C143 a_n1035_3765# CM_MSB_V2_0.SD 3.62e-19
C144 a_n1035_4741# Local_Enc_0.QB 0.0055f
C145 a_n1846_3765# CM_MSB_V2_0.SD 3.72e-19
C146 IOUT+ Local_Enc_0.QB 1.83f
C147 Local_Enc_0.NAND_5.B Ci 0.0105f
C148 Local_Enc_0.NAND_5.B VDD 0.864f
C149 Local_Enc_0.NAND_5.B Local_Enc_0.NAND_6.B 0.0342f
C150 Local_Enc_0.NAND_5.A Local_Enc_0.NAND_8.A 0.333f
C151 IM IOUT+ 8.52e-21
C152 CM_MSB_V2_0.SD Local_Enc_0.QB 0.00262f
C153 Local_Enc_0.QB CM_MSB_V2_0.OUT 2.71f
C154 a_n2609_3766# Local_Enc_0.NAND_6.A 0.0419f
C155 Local_Enc_0.NAND_5.B Local_Enc_0.Q 0.0478f
C156 Ri CM_MSB_V2_0.SD 9.7e-19
C157 IM CM_MSB_V2_0.SD 0.916f
C158 IM CM_MSB_V2_0.OUT 1.33f
C159 IOUT- VSS 2.91f
C160 IOUT+ VSS 3.17f
C161 CM_MSB_V2_0.SD VSS 5.44f
C162 IM VSS 8.13f
C163 IM_T VSS 14.9f
C164 a_n1035_3765# VSS 0.0983f
C165 a_n1846_3765# VSS 0.0986f
C166 a_n2609_3766# VSS 0.0998f
C167 Local_Enc_0.NAND_6.A VSS 0.56f
C168 Ri VSS 0.635f
C169 a_n1035_4741# VSS 0.0983f
C170 a_n1846_4741# VSS 0.0983f
C171 a_n2609_4741# VSS 0.0997f
C172 Local_Enc_0.NAND_6.B VSS 0.669f
C173 Local_Enc_0.NAND_8.A VSS 1.42f
C174 Local_Enc_0.NAND_5.A VSS 0.674f
C175 Ci VSS 0.628f
C176 a_n1035_5712# VSS 0.0983f
C177 a_n1846_5712# VSS 0.0983f
C178 a_n2609_5712# VSS 0.0983f
C179 Local_Enc_0.NAND_5.B VSS 0.697f
C180 Local_Enc_0.NAND_4.B VSS 0.67f
C181 Local_Enc_0.NAND_1.B VSS 0.754f
C182 Ri-1 VSS 0.613f
C183 CM_MSB_V2_0.OUT VSS 9.61f
C184 Local_Enc_0.QB VSS 18.3f
C185 Local_Enc_0.Q VSS 20.1f
C186 VDD VSS 14f
C187 IOUT+.n0 VSS 0.0568f
C188 IOUT+.t30 VSS 0.024f
C189 IOUT+.n1 VSS 0.024f
C190 IOUT+.n2 VSS 0.0568f
C191 IOUT+.t34 VSS 0.024f
C192 IOUT+.n3 VSS 0.024f
C193 IOUT+.n4 VSS 0.0495f
C194 IOUT+.t24 VSS 0.024f
C195 IOUT+.n5 VSS 0.024f
C196 IOUT+.n6 VSS 0.0831f
C197 IOUT+.t55 VSS 0.024f
C198 IOUT+.n7 VSS 0.024f
C199 IOUT+.n8 VSS 0.109f
C200 IOUT+.t38 VSS 0.024f
C201 IOUT+.n9 VSS 0.024f
C202 IOUT+.n10 VSS 0.0495f
C203 IOUT+.t18 VSS 0.024f
C204 IOUT+.n11 VSS 0.024f
C205 IOUT+.n12 VSS 0.0874f
C206 IOUT+.n13 VSS 0.307f
C207 IOUT+.t4 VSS 0.124f
C208 IOUT+.n14 VSS 0.516f
C209 IOUT+.n15 VSS 0.319f
C210 IOUT+.n16 VSS 0.227f
C211 IOUT+.t16 VSS 0.024f
C212 IOUT+.n17 VSS 0.024f
C213 IOUT+.n18 VSS 0.108f
C214 IOUT+.n19 VSS 0.399f
C215 IOUT+.n20 VSS 0.191f
C216 IOUT+.n21 VSS 0.244f
C217 IOUT+.n22 VSS 0.211f
C218 IOUT+.n23 VSS 0.0957f
C219 IOUT+.n24 VSS 0.0575f
C220 IOUT+.t2 VSS 0.024f
C221 IOUT+.n25 VSS 0.024f
C222 IOUT+.n26 VSS 0.0568f
C223 IOUT+.t48 VSS 0.024f
C224 IOUT+.n27 VSS 0.024f
C225 IOUT+.n28 VSS 0.0495f
C226 IOUT+.t37 VSS 0.024f
C227 IOUT+.n29 VSS 0.024f
C228 IOUT+.n30 VSS 0.0831f
C229 IOUT+.t27 VSS 0.024f
C230 IOUT+.n31 VSS 0.024f
C231 IOUT+.n32 VSS 0.109f
C232 IOUT+.t51 VSS 0.024f
C233 IOUT+.n33 VSS 0.024f
C234 IOUT+.n34 VSS 0.0495f
C235 IOUT+.t57 VSS 0.024f
C236 IOUT+.n35 VSS 0.024f
C237 IOUT+.n36 VSS 0.0874f
C238 IOUT+.n37 VSS 0.307f
C239 IOUT+.t17 VSS 0.124f
C240 IOUT+.n38 VSS 0.516f
C241 IOUT+.n39 VSS 0.319f
C242 IOUT+.n40 VSS 0.227f
C243 IOUT+.t54 VSS 0.024f
C244 IOUT+.n41 VSS 0.024f
C245 IOUT+.n42 VSS 0.108f
C246 IOUT+.n43 VSS 0.399f
C247 IOUT+.n44 VSS 0.191f
C248 IOUT+.n45 VSS 0.24f
C249 IOUT+.n46 VSS 0.292f
C250 IOUT+.n47 VSS 0.0568f
C251 IOUT+.t35 VSS 0.024f
C252 IOUT+.n48 VSS 0.024f
C253 IOUT+.n49 VSS 0.0568f
C254 IOUT+.t21 VSS 0.024f
C255 IOUT+.n50 VSS 0.024f
C256 IOUT+.n51 VSS 0.0495f
C257 IOUT+.t11 VSS 0.024f
C258 IOUT+.n52 VSS 0.024f
C259 IOUT+.n53 VSS 0.0831f
C260 IOUT+.t1 VSS 0.024f
C261 IOUT+.n54 VSS 0.024f
C262 IOUT+.n55 VSS 0.109f
C263 IOUT+.t23 VSS 0.024f
C264 IOUT+.n56 VSS 0.024f
C265 IOUT+.n57 VSS 0.0495f
C266 IOUT+.t29 VSS 0.024f
C267 IOUT+.n58 VSS 0.024f
C268 IOUT+.n59 VSS 0.0874f
C269 IOUT+.n60 VSS 0.307f
C270 IOUT+.t56 VSS 0.124f
C271 IOUT+.n61 VSS 0.516f
C272 IOUT+.n62 VSS 0.319f
C273 IOUT+.n63 VSS 0.227f
C274 IOUT+.t26 VSS 0.024f
C275 IOUT+.n64 VSS 0.024f
C276 IOUT+.n65 VSS 0.108f
C277 IOUT+.n66 VSS 0.399f
C278 IOUT+.n67 VSS 0.191f
C279 IOUT+.n68 VSS 0.244f
C280 IOUT+.n69 VSS 0.286f
C281 IOUT+.n70 VSS 0.0575f
C282 IOUT+.t50 VSS 0.024f
C283 IOUT+.n71 VSS 0.024f
C284 IOUT+.n72 VSS 0.0568f
C285 IOUT+.t61 VSS 0.024f
C286 IOUT+.n73 VSS 0.024f
C287 IOUT+.n74 VSS 0.0495f
C288 IOUT+.t46 VSS 0.024f
C289 IOUT+.n75 VSS 0.024f
C290 IOUT+.n76 VSS 0.0831f
C291 IOUT+.t12 VSS 0.024f
C292 IOUT+.n77 VSS 0.024f
C293 IOUT+.n78 VSS 0.109f
C294 IOUT+.t0 VSS 0.024f
C295 IOUT+.n79 VSS 0.024f
C296 IOUT+.n80 VSS 0.0495f
C297 IOUT+.t40 VSS 0.024f
C298 IOUT+.n81 VSS 0.024f
C299 IOUT+.n82 VSS 0.0874f
C300 IOUT+.n83 VSS 0.307f
C301 IOUT+.t28 VSS 0.124f
C302 IOUT+.n84 VSS 0.516f
C303 IOUT+.n85 VSS 0.319f
C304 IOUT+.n86 VSS 0.227f
C305 IOUT+.t39 VSS 0.024f
C306 IOUT+.n87 VSS 0.024f
C307 IOUT+.n88 VSS 0.108f
C308 IOUT+.n89 VSS 0.399f
C309 IOUT+.n90 VSS 0.191f
C310 IOUT+.n91 VSS 0.24f
C311 IOUT+.n92 VSS 0.36f
C312 IOUT+.n93 VSS 0.533f
C313 IOUT+.n94 VSS 0.377f
C314 Local_Enc_0.Q.t14 VSS 0.0669f
C315 Local_Enc_0.Q.t31 VSS 0.0398f
C316 Local_Enc_0.Q.n0 VSS 0.114f
C317 Local_Enc_0.Q.t24 VSS 0.0398f
C318 Local_Enc_0.Q.n1 VSS 0.0761f
C319 Local_Enc_0.Q.t5 VSS 0.0412f
C320 Local_Enc_0.Q.n2 VSS 0.0779f
C321 Local_Enc_0.Q.t43 VSS 0.0412f
C322 Local_Enc_0.Q.n3 VSS 0.0779f
C323 Local_Enc_0.Q.t42 VSS 0.0398f
C324 Local_Enc_0.Q.n4 VSS 0.0761f
C325 Local_Enc_0.Q.t6 VSS 0.0398f
C326 Local_Enc_0.Q.n5 VSS 0.0761f
C327 Local_Enc_0.Q.t20 VSS 0.0412f
C328 Local_Enc_0.Q.n6 VSS 0.0779f
C329 Local_Enc_0.Q.t55 VSS 0.0412f
C330 Local_Enc_0.Q.n7 VSS 0.0779f
C331 Local_Enc_0.Q.t67 VSS 0.0398f
C332 Local_Enc_0.Q.n8 VSS 0.0761f
C333 Local_Enc_0.Q.t22 VSS 0.0398f
C334 Local_Enc_0.Q.n9 VSS 0.0761f
C335 Local_Enc_0.Q.t68 VSS 0.0412f
C336 Local_Enc_0.Q.n10 VSS 0.0779f
C337 Local_Enc_0.Q.t23 VSS 0.0412f
C338 Local_Enc_0.Q.n11 VSS 0.0779f
C339 Local_Enc_0.Q.t39 VSS 0.0398f
C340 Local_Enc_0.Q.n12 VSS 0.0761f
C341 Local_Enc_0.Q.t4 VSS 0.0398f
C342 Local_Enc_0.Q.n13 VSS 0.0824f
C343 Local_Enc_0.Q.t40 VSS 0.0357f
C344 Local_Enc_0.Q.n14 VSS 0.0765f
C345 Local_Enc_0.Q.t35 VSS 0.133f
C346 Local_Enc_0.Q.t32 VSS 0.0412f
C347 Local_Enc_0.Q.n15 VSS 0.161f
C348 Local_Enc_0.Q.t65 VSS 0.0412f
C349 Local_Enc_0.Q.n16 VSS 0.134f
C350 Local_Enc_0.Q.t44 VSS 0.0412f
C351 Local_Enc_0.Q.n17 VSS 0.134f
C352 Local_Enc_0.Q.t7 VSS 0.0412f
C353 Local_Enc_0.Q.n18 VSS 0.134f
C354 Local_Enc_0.Q.t28 VSS 0.0412f
C355 Local_Enc_0.Q.n19 VSS 0.134f
C356 Local_Enc_0.Q.t48 VSS 0.0412f
C357 Local_Enc_0.Q.n20 VSS 0.138f
C358 Local_Enc_0.Q.t64 VSS 0.0357f
C359 Local_Enc_0.Q.n21 VSS 0.169f
C360 Local_Enc_0.Q.t21 VSS 0.0669f
C361 Local_Enc_0.Q.t38 VSS 0.0398f
C362 Local_Enc_0.Q.n22 VSS 0.114f
C363 Local_Enc_0.Q.t34 VSS 0.0398f
C364 Local_Enc_0.Q.n23 VSS 0.0761f
C365 Local_Enc_0.Q.t18 VSS 0.0412f
C366 Local_Enc_0.Q.n24 VSS 0.0779f
C367 Local_Enc_0.Q.t53 VSS 0.0412f
C368 Local_Enc_0.Q.n25 VSS 0.0779f
C369 Local_Enc_0.Q.t52 VSS 0.0398f
C370 Local_Enc_0.Q.n26 VSS 0.0761f
C371 Local_Enc_0.Q.t19 VSS 0.0398f
C372 Local_Enc_0.Q.n27 VSS 0.0761f
C373 Local_Enc_0.Q.t29 VSS 0.0412f
C374 Local_Enc_0.Q.n28 VSS 0.0779f
C375 Local_Enc_0.Q.t63 VSS 0.0412f
C376 Local_Enc_0.Q.n29 VSS 0.0779f
C377 Local_Enc_0.Q.t11 VSS 0.0398f
C378 Local_Enc_0.Q.n30 VSS 0.0761f
C379 Local_Enc_0.Q.t30 VSS 0.0398f
C380 Local_Enc_0.Q.n31 VSS 0.0761f
C381 Local_Enc_0.Q.t15 VSS 0.0412f
C382 Local_Enc_0.Q.n32 VSS 0.0779f
C383 Local_Enc_0.Q.t33 VSS 0.0412f
C384 Local_Enc_0.Q.n33 VSS 0.0779f
C385 Local_Enc_0.Q.t50 VSS 0.0398f
C386 Local_Enc_0.Q.n34 VSS 0.0761f
C387 Local_Enc_0.Q.t17 VSS 0.0398f
C388 Local_Enc_0.Q.n35 VSS 0.0824f
C389 Local_Enc_0.Q.t51 VSS 0.0357f
C390 Local_Enc_0.Q.n36 VSS 0.0942f
C391 Local_Enc_0.Q.n37 VSS 0.333f
C392 Local_Enc_0.Q.t54 VSS 0.0669f
C393 Local_Enc_0.Q.t66 VSS 0.0398f
C394 Local_Enc_0.Q.n38 VSS 0.114f
C395 Local_Enc_0.Q.t61 VSS 0.0398f
C396 Local_Enc_0.Q.n39 VSS 0.0761f
C397 Local_Enc_0.Q.t47 VSS 0.0412f
C398 Local_Enc_0.Q.n40 VSS 0.0779f
C399 Local_Enc_0.Q.t13 VSS 0.0412f
C400 Local_Enc_0.Q.n41 VSS 0.0779f
C401 Local_Enc_0.Q.t12 VSS 0.0398f
C402 Local_Enc_0.Q.n42 VSS 0.0761f
C403 Local_Enc_0.Q.t49 VSS 0.0398f
C404 Local_Enc_0.Q.n43 VSS 0.0761f
C405 Local_Enc_0.Q.t57 VSS 0.0412f
C406 Local_Enc_0.Q.n44 VSS 0.0779f
C407 Local_Enc_0.Q.t25 VSS 0.0412f
C408 Local_Enc_0.Q.n45 VSS 0.0779f
C409 Local_Enc_0.Q.t41 VSS 0.0398f
C410 Local_Enc_0.Q.n46 VSS 0.0761f
C411 Local_Enc_0.Q.t58 VSS 0.0398f
C412 Local_Enc_0.Q.n47 VSS 0.0761f
C413 Local_Enc_0.Q.t45 VSS 0.0412f
C414 Local_Enc_0.Q.n48 VSS 0.0779f
C415 Local_Enc_0.Q.t60 VSS 0.0412f
C416 Local_Enc_0.Q.n49 VSS 0.0779f
C417 Local_Enc_0.Q.t9 VSS 0.0398f
C418 Local_Enc_0.Q.n50 VSS 0.0761f
C419 Local_Enc_0.Q.t46 VSS 0.0398f
C420 Local_Enc_0.Q.n51 VSS 0.0824f
C421 Local_Enc_0.Q.t10 VSS 0.0357f
C422 Local_Enc_0.Q.n52 VSS 0.0942f
C423 Local_Enc_0.Q.n53 VSS 0.212f
C424 Local_Enc_0.Q.t16 VSS 0.0641f
C425 Local_Enc_0.Q.t8 VSS 0.0373f
C426 Local_Enc_0.Q.n54 VSS 0.118f
C427 Local_Enc_0.Q.t27 VSS 0.0373f
C428 Local_Enc_0.Q.n55 VSS 0.0952f
C429 Local_Enc_0.Q.t62 VSS 0.0373f
C430 Local_Enc_0.Q.n56 VSS 0.0952f
C431 Local_Enc_0.Q.t56 VSS 0.0373f
C432 Local_Enc_0.Q.n57 VSS 0.0952f
C433 Local_Enc_0.Q.t3 VSS 0.0373f
C434 Local_Enc_0.Q.n58 VSS 0.0952f
C435 Local_Enc_0.Q.t26 VSS 0.0373f
C436 Local_Enc_0.Q.n59 VSS 0.0952f
C437 Local_Enc_0.Q.t59 VSS 0.0373f
C438 Local_Enc_0.Q.n60 VSS 0.0913f
C439 Local_Enc_0.Q.n61 VSS 0.336f
C440 Local_Enc_0.Q.n62 VSS 0.213f
C441 Local_Enc_0.Q.n63 VSS 0.0225f
C442 Local_Enc_0.Q.t36 VSS 0.0234f
C443 Local_Enc_0.Q.t37 VSS 0.0134f
C444 Local_Enc_0.Q.n64 VSS 0.0611f
C445 Local_Enc_0.Q.t1 VSS 0.00924f
C446 Local_Enc_0.Q.n65 VSS 0.00924f
C447 Local_Enc_0.Q.n66 VSS 0.0185f
C448 Local_Enc_0.Q.n67 VSS 0.158f
C449 CM_MSB_V2_0.SD.n0 VSS 0.101f
C450 CM_MSB_V2_0.SD.n1 VSS 0.103f
C451 CM_MSB_V2_0.SD.n2 VSS 0.104f
C452 CM_MSB_V2_0.SD.n3 VSS 0.0988f
C453 CM_MSB_V2_0.SD.n4 VSS 0.103f
C454 CM_MSB_V2_0.SD.n5 VSS 0.105f
C455 CM_MSB_V2_0.SD.n6 VSS 0.104f
C456 CM_MSB_V2_0.SD.n7 VSS 0.0127f
C457 CM_MSB_V2_0.SD.t27 VSS 0.0151f
C458 CM_MSB_V2_0.SD.n8 VSS 0.0561f
C459 CM_MSB_V2_0.SD.t54 VSS 0.0128f
C460 CM_MSB_V2_0.SD.n9 VSS 0.0149f
C461 CM_MSB_V2_0.SD.n10 VSS 0.0557f
C462 CM_MSB_V2_0.SD.t21 VSS 0.015f
C463 CM_MSB_V2_0.SD.n11 VSS 0.0128f
C464 CM_MSB_V2_0.SD.n12 VSS 0.0452f
C465 CM_MSB_V2_0.SD.t40 VSS 0.0136f
C466 CM_MSB_V2_0.SD.n13 VSS 0.0136f
C467 CM_MSB_V2_0.SD.n14 VSS 0.0276f
C468 CM_MSB_V2_0.SD.n15 VSS 0.0312f
C469 CM_MSB_V2_0.SD.t10 VSS 0.0136f
C470 CM_MSB_V2_0.SD.n16 VSS 0.0136f
C471 CM_MSB_V2_0.SD.n17 VSS 0.0532f
C472 CM_MSB_V2_0.SD.t39 VSS 0.0136f
C473 CM_MSB_V2_0.SD.n18 VSS 0.0136f
C474 CM_MSB_V2_0.SD.n19 VSS 0.0541f
C475 CM_MSB_V2_0.SD.t51 VSS 0.0136f
C476 CM_MSB_V2_0.SD.n20 VSS 0.0136f
C477 CM_MSB_V2_0.SD.n21 VSS 0.0276f
C478 CM_MSB_V2_0.SD.n22 VSS 0.0312f
C479 CM_MSB_V2_0.SD.t4 VSS 0.015f
C480 CM_MSB_V2_0.SD.n23 VSS 0.0128f
C481 CM_MSB_V2_0.SD.n24 VSS 0.0563f
C482 CM_MSB_V2_0.SD.t33 VSS 0.0136f
C483 CM_MSB_V2_0.SD.n25 VSS 0.0136f
C484 CM_MSB_V2_0.SD.n26 VSS 0.053f
C485 CM_MSB_V2_0.SD.t20 VSS 0.0136f
C486 CM_MSB_V2_0.SD.n27 VSS 0.0136f
C487 CM_MSB_V2_0.SD.n28 VSS 0.053f
C488 CM_MSB_V2_0.SD.t36 VSS 0.0136f
C489 CM_MSB_V2_0.SD.n29 VSS 0.0136f
C490 CM_MSB_V2_0.SD.n30 VSS 0.0276f
C491 CM_MSB_V2_0.SD.n31 VSS 0.0312f
C492 CM_MSB_V2_0.SD.n32 VSS 0.0127f
C493 CM_MSB_V2_0.SD.t42 VSS 0.0151f
C494 CM_MSB_V2_0.SD.n33 VSS 0.0563f
C495 CM_MSB_V2_0.SD.t13 VSS 0.0136f
C496 CM_MSB_V2_0.SD.n34 VSS 0.0136f
C497 CM_MSB_V2_0.SD.n35 VSS 0.0276f
C498 CM_MSB_V2_0.SD.n36 VSS 0.0312f
C499 CM_MSB_V2_0.SD.t24 VSS 0.0136f
C500 CM_MSB_V2_0.SD.n37 VSS 0.0136f
C501 CM_MSB_V2_0.SD.n38 VSS 0.0529f
C502 CM_MSB_V2_0.SD.t50 VSS 0.0149f
C503 CM_MSB_V2_0.SD.n39 VSS 0.0128f
C504 CM_MSB_V2_0.SD.n40 VSS 0.0559f
C505 CM_MSB_V2_0.SD.t28 VSS 0.0136f
C506 CM_MSB_V2_0.SD.n41 VSS 0.0136f
C507 CM_MSB_V2_0.SD.n42 VSS 0.0276f
C508 CM_MSB_V2_0.SD.n43 VSS 0.0312f
C509 CM_MSB_V2_0.SD.t60 VSS 0.0136f
C510 CM_MSB_V2_0.SD.n44 VSS 0.0136f
C511 CM_MSB_V2_0.SD.n45 VSS 0.0413f
C512 CM_MSB_V2_0.SD.t7 VSS 0.0133f
C513 CM_MSB_V2_0.SD.n46 VSS 0.0144f
C514 CM_MSB_V2_0.SD.n47 VSS 0.0567f
C515 CM_MSB_V2_0.SD.n48 VSS 0.125f
C516 CM_MSB_V2_0.SD.n49 VSS 0.0272f
C517 CM_MSB_V2_0.SD.n50 VSS 0.0724f
C518 CM_MSB_V2_0.SD.n51 VSS 0.0268f
C519 CM_MSB_V2_0.SD.t45 VSS 0.0128f
C520 CM_MSB_V2_0.SD.n52 VSS 0.0149f
C521 CM_MSB_V2_0.SD.n53 VSS 0.0271f
C522 CM_MSB_V2_0.SD.n54 VSS 0.0312f
C523 CM_MSB_V2_0.SD.n55 VSS 0.0258f
C524 CM_MSB_V2_0.SD.n56 VSS 0.0263f
C525 CM_MSB_V2_0.SD.n57 VSS 0.0737f
C526 CM_MSB_V2_0.SD.n58 VSS 0.0262f
C527 CM_MSB_V2_0.SD.n59 VSS 0.0273f
C528 CM_MSB_V2_0.SD.n60 VSS 0.077f
C529 CM_MSB_V2_0.SD.n61 VSS 0.0269f
C530 CM_MSB_V2_0.SD.n62 VSS 0.0149f
C531 CM_MSB_V2_0.SD.t8 VSS 0.0128f
C532 CM_MSB_V2_0.SD.n63 VSS 0.0271f
C533 CM_MSB_V2_0.SD.n64 VSS 0.0312f
C534 CM_MSB_V2_0.SD.n65 VSS 0.027f
C535 CM_MSB_V2_0.SD.n66 VSS 0.026f
C536 CM_MSB_V2_0.SD.t15 VSS 0.0128f
C537 CM_MSB_V2_0.SD.n67 VSS 0.015f
C538 CM_MSB_V2_0.SD.n68 VSS 0.0273f
C539 CM_MSB_V2_0.SD.n69 VSS 0.0312f
C540 CM_MSB_V2_0.SD.n70 VSS 0.0256f
C541 CM_MSB_V2_0.SD.n71 VSS 0.0263f
C542 CM_MSB_V2_0.SD.n72 VSS 0.0402f
C543 CM_MSB_V2_0.SD.n73 VSS 0.0979f
C544 CM_MSB_V2_0.SD.t55 VSS 0.0129f
C545 CM_MSB_V2_0.SD.n74 VSS 0.0148f
C546 CM_MSB_V2_0.SD.n75 VSS 0.0272f
C547 CM_MSB_V2_0.SD.n76 VSS 0.0312f
C548 CM_MSB_V2_0.SD.t61 VSS 0.0136f
C549 CM_MSB_V2_0.SD.n77 VSS 0.0136f
C550 CM_MSB_V2_0.SD.n78 VSS 0.0522f
C551 CM_MSB_V2_0.SD.t18 VSS 0.0136f
C552 CM_MSB_V2_0.SD.n79 VSS 0.0136f
C553 CM_MSB_V2_0.SD.n80 VSS 0.0527f
C554 CM_MSB_V2_0.SD.t52 VSS 0.015f
C555 CM_MSB_V2_0.SD.n81 VSS 0.0128f
C556 CM_MSB_V2_0.SD.n82 VSS 0.0558f
C557 CM_MSB_V2_0.SD.t32 VSS 0.0136f
C558 CM_MSB_V2_0.SD.n83 VSS 0.0136f
C559 CM_MSB_V2_0.SD.n84 VSS 0.0277f
C560 CM_MSB_V2_0.SD.n85 VSS 0.0311f
C561 CM_MSB_V2_0.SD.t1 VSS 0.0136f
C562 CM_MSB_V2_0.SD.n86 VSS 0.0136f
C563 CM_MSB_V2_0.SD.n87 VSS 0.0535f
C564 CM_MSB_V2_0.SD.t62 VSS 0.0136f
C565 CM_MSB_V2_0.SD.n88 VSS 0.0136f
C566 CM_MSB_V2_0.SD.n89 VSS 0.0538f
C567 CM_MSB_V2_0.SD.t6 VSS 0.0136f
C568 CM_MSB_V2_0.SD.n90 VSS 0.0136f
C569 CM_MSB_V2_0.SD.n91 VSS 0.0412f
C570 CM_MSB_V2_0.SD.n92 VSS 0.129f
C571 CM_MSB_V2_0.SD.t56 VSS 0.0146f
C572 CM_MSB_V2_0.SD.n93 VSS 0.0132f
C573 CM_MSB_V2_0.SD.n94 VSS 0.0272f
C574 CM_MSB_V2_0.SD.n95 VSS 0.0312f
C575 CM_MSB_V2_0.SD.n96 VSS 0.027f
C576 CM_MSB_V2_0.SD.n97 VSS 0.0264f
C577 CM_MSB_V2_0.SD.n98 VSS 0.0723f
C578 CM_MSB_V2_0.SD.n99 VSS 0.0267f
C579 CM_MSB_V2_0.SD.n100 VSS 0.101f
C580 CM_MSB_V2_0.SD.n101 VSS 0.0127f
C581 CM_MSB_V2_0.SD.t0 VSS 0.0151f
C582 CM_MSB_V2_0.SD.n102 VSS 0.0451f
C583 CM_MSB_V2_0.SD.n103 VSS 0.0398f
C584 CM_MSB_V2_0.SD.n104 VSS 0.0263f
C585 CM_MSB_V2_0.SD.n105 VSS 0.0752f
C586 CM_MSB_V2_0.SD.t2 VSS 0.0136f
C587 CM_MSB_V2_0.SD.n106 VSS 0.0136f
C588 CM_MSB_V2_0.SD.n107 VSS 0.0277f
C589 CM_MSB_V2_0.SD.n108 VSS 0.0311f
C590 CM_MSB_V2_0.SD.n109 VSS 0.0252f
C591 CM_MSB_V2_0.SD.n110 VSS 0.0258f
C592 IOUT-.n0 VSS 0.0744f
C593 IOUT-.t15 VSS 0.0209f
C594 IOUT-.n1 VSS 0.0209f
C595 IOUT-.n2 VSS 0.0733f
C596 IOUT-.t52 VSS 0.0209f
C597 IOUT-.n3 VSS 0.0209f
C598 IOUT-.n4 VSS 0.0733f
C599 IOUT-.t18 VSS 0.0209f
C600 IOUT-.n5 VSS 0.0209f
C601 IOUT-.n6 VSS 0.115f
C602 IOUT-.n7 VSS 0.543f
C603 IOUT-.n8 VSS 0.361f
C604 IOUT-.t26 VSS 0.0209f
C605 IOUT-.n9 VSS 0.0209f
C606 IOUT-.n10 VSS 0.0733f
C607 IOUT-.n11 VSS 0.287f
C608 IOUT-.t31 VSS 0.0209f
C609 IOUT-.n12 VSS 0.0209f
C610 IOUT-.n13 VSS 0.072f
C611 IOUT-.t19 VSS 0.0209f
C612 IOUT-.n14 VSS 0.0209f
C613 IOUT-.n15 VSS 0.073f
C614 IOUT-.t32 VSS 0.0209f
C615 IOUT-.n16 VSS 0.0209f
C616 IOUT-.n17 VSS 0.0717f
C617 IOUT-.t59 VSS 0.127f
C618 IOUT-.n18 VSS 0.553f
C619 IOUT-.n19 VSS 0.362f
C620 IOUT-.n20 VSS 0.286f
C621 IOUT-.n21 VSS 0.214f
C622 IOUT-.n22 VSS 0.345f
C623 IOUT-.n23 VSS 0.0744f
C624 IOUT-.t42 VSS 0.0209f
C625 IOUT-.n24 VSS 0.0209f
C626 IOUT-.n25 VSS 0.0733f
C627 IOUT-.t16 VSS 0.0209f
C628 IOUT-.n26 VSS 0.0209f
C629 IOUT-.n27 VSS 0.0733f
C630 IOUT-.t45 VSS 0.0209f
C631 IOUT-.n28 VSS 0.0209f
C632 IOUT-.n29 VSS 0.115f
C633 IOUT-.n30 VSS 0.543f
C634 IOUT-.n31 VSS 0.361f
C635 IOUT-.t53 VSS 0.0209f
C636 IOUT-.n32 VSS 0.0209f
C637 IOUT-.n33 VSS 0.0733f
C638 IOUT-.n34 VSS 0.287f
C639 IOUT-.t17 VSS 0.0209f
C640 IOUT-.n35 VSS 0.0209f
C641 IOUT-.n36 VSS 0.072f
C642 IOUT-.t1 VSS 0.0209f
C643 IOUT-.n37 VSS 0.0209f
C644 IOUT-.n38 VSS 0.073f
C645 IOUT-.t20 VSS 0.0209f
C646 IOUT-.n39 VSS 0.0209f
C647 IOUT-.n40 VSS 0.0717f
C648 IOUT-.t50 VSS 0.127f
C649 IOUT-.n41 VSS 0.553f
C650 IOUT-.n42 VSS 0.362f
C651 IOUT-.n43 VSS 0.286f
C652 IOUT-.n44 VSS 0.214f
C653 IOUT-.n45 VSS 0.196f
C654 IOUT-.n46 VSS 0.356f
C655 IOUT-.n47 VSS 0.0744f
C656 IOUT-.t3 VSS 0.0209f
C657 IOUT-.n48 VSS 0.0209f
C658 IOUT-.n49 VSS 0.0733f
C659 IOUT-.t43 VSS 0.0209f
C660 IOUT-.n50 VSS 0.0209f
C661 IOUT-.n51 VSS 0.0733f
C662 IOUT-.t5 VSS 0.0209f
C663 IOUT-.n52 VSS 0.0209f
C664 IOUT-.n53 VSS 0.115f
C665 IOUT-.n54 VSS 0.543f
C666 IOUT-.n55 VSS 0.361f
C667 IOUT-.t21 VSS 0.0209f
C668 IOUT-.n56 VSS 0.0209f
C669 IOUT-.n57 VSS 0.0733f
C670 IOUT-.n58 VSS 0.287f
C671 IOUT-.t44 VSS 0.0209f
C672 IOUT-.n59 VSS 0.0209f
C673 IOUT-.n60 VSS 0.072f
C674 IOUT-.t33 VSS 0.0209f
C675 IOUT-.n61 VSS 0.0209f
C676 IOUT-.n62 VSS 0.073f
C677 IOUT-.t47 VSS 0.0209f
C678 IOUT-.n63 VSS 0.0209f
C679 IOUT-.n64 VSS 0.0717f
C680 IOUT-.t12 VSS 0.127f
C681 IOUT-.n65 VSS 0.553f
C682 IOUT-.n66 VSS 0.362f
C683 IOUT-.n67 VSS 0.286f
C684 IOUT-.n68 VSS 0.214f
C685 IOUT-.n69 VSS 0.196f
C686 IOUT-.n70 VSS 0.353f
C687 IOUT-.n71 VSS 0.0744f
C688 IOUT-.t55 VSS 0.0209f
C689 IOUT-.n72 VSS 0.0209f
C690 IOUT-.n73 VSS 0.0733f
C691 IOUT-.t30 VSS 0.0209f
C692 IOUT-.n74 VSS 0.0209f
C693 IOUT-.n75 VSS 0.0733f
C694 IOUT-.t56 VSS 0.0209f
C695 IOUT-.n76 VSS 0.0209f
C696 IOUT-.n77 VSS 0.115f
C697 IOUT-.n78 VSS 0.543f
C698 IOUT-.n79 VSS 0.361f
C699 IOUT-.t2 VSS 0.0209f
C700 IOUT-.n80 VSS 0.0209f
C701 IOUT-.n81 VSS 0.0733f
C702 IOUT-.n82 VSS 0.287f
C703 IOUT-.t4 VSS 0.0209f
C704 IOUT-.n83 VSS 0.0209f
C705 IOUT-.n84 VSS 0.072f
C706 IOUT-.t57 VSS 0.0209f
C707 IOUT-.n85 VSS 0.0209f
C708 IOUT-.n86 VSS 0.073f
C709 IOUT-.t6 VSS 0.0209f
C710 IOUT-.n87 VSS 0.0209f
C711 IOUT-.n88 VSS 0.0717f
C712 IOUT-.t41 VSS 0.127f
C713 IOUT-.n89 VSS 0.553f
C714 IOUT-.n90 VSS 0.362f
C715 IOUT-.n91 VSS 0.286f
C716 IOUT-.n92 VSS 0.214f
C717 IOUT-.n93 VSS 0.16f
C718 CM_MSB_V2_0.OUT.t45 VSS 0.0182f
C719 CM_MSB_V2_0.OUT.n0 VSS 0.0182f
C720 CM_MSB_V2_0.OUT.n1 VSS 0.0387f
C721 CM_MSB_V2_0.OUT.t87 VSS 0.0182f
C722 CM_MSB_V2_0.OUT.n2 VSS 0.0182f
C723 CM_MSB_V2_0.OUT.n3 VSS 0.0387f
C724 CM_MSB_V2_0.OUT.t133 VSS 0.0182f
C725 CM_MSB_V2_0.OUT.n4 VSS 0.0182f
C726 CM_MSB_V2_0.OUT.n5 VSS 0.0394f
C727 CM_MSB_V2_0.OUT.t50 VSS 0.0182f
C728 CM_MSB_V2_0.OUT.n6 VSS 0.0182f
C729 CM_MSB_V2_0.OUT.n7 VSS 0.0408f
C730 CM_MSB_V2_0.OUT.t38 VSS 0.0182f
C731 CM_MSB_V2_0.OUT.n8 VSS 0.0182f
C732 CM_MSB_V2_0.OUT.n9 VSS 0.0394f
C733 CM_MSB_V2_0.OUT.t130 VSS 0.0182f
C734 CM_MSB_V2_0.OUT.n10 VSS 0.0182f
C735 CM_MSB_V2_0.OUT.n11 VSS 0.0407f
C736 CM_MSB_V2_0.OUT.n12 VSS 0.203f
C737 CM_MSB_V2_0.OUT.n13 VSS 0.26f
C738 CM_MSB_V2_0.OUT.t100 VSS 0.0182f
C739 CM_MSB_V2_0.OUT.n14 VSS 0.0182f
C740 CM_MSB_V2_0.OUT.n15 VSS 0.0394f
C741 CM_MSB_V2_0.OUT.t62 VSS 0.0182f
C742 CM_MSB_V2_0.OUT.n16 VSS 0.0182f
C743 CM_MSB_V2_0.OUT.n17 VSS 0.0408f
C744 CM_MSB_V2_0.OUT.t54 VSS 0.0182f
C745 CM_MSB_V2_0.OUT.n18 VSS 0.0182f
C746 CM_MSB_V2_0.OUT.n19 VSS 0.0394f
C747 CM_MSB_V2_0.OUT.t136 VSS 0.0182f
C748 CM_MSB_V2_0.OUT.n20 VSS 0.0182f
C749 CM_MSB_V2_0.OUT.n21 VSS 0.0407f
C750 CM_MSB_V2_0.OUT.n22 VSS 0.203f
C751 CM_MSB_V2_0.OUT.n23 VSS 0.26f
C752 CM_MSB_V2_0.OUT.t97 VSS 0.0182f
C753 CM_MSB_V2_0.OUT.n24 VSS 0.0182f
C754 CM_MSB_V2_0.OUT.n25 VSS 0.0394f
C755 CM_MSB_V2_0.OUT.t43 VSS 0.0182f
C756 CM_MSB_V2_0.OUT.n26 VSS 0.0182f
C757 CM_MSB_V2_0.OUT.n27 VSS 0.0408f
C758 CM_MSB_V2_0.OUT.t35 VSS 0.0182f
C759 CM_MSB_V2_0.OUT.n28 VSS 0.0182f
C760 CM_MSB_V2_0.OUT.n29 VSS 0.0394f
C761 CM_MSB_V2_0.OUT.t116 VSS 0.0182f
C762 CM_MSB_V2_0.OUT.n30 VSS 0.0182f
C763 CM_MSB_V2_0.OUT.n31 VSS 0.0407f
C764 CM_MSB_V2_0.OUT.n32 VSS 0.203f
C765 CM_MSB_V2_0.OUT.n33 VSS 0.26f
C766 CM_MSB_V2_0.OUT.t146 VSS 0.0182f
C767 CM_MSB_V2_0.OUT.n34 VSS 0.0182f
C768 CM_MSB_V2_0.OUT.n35 VSS 0.0408f
C769 CM_MSB_V2_0.OUT.t46 VSS 0.0182f
C770 CM_MSB_V2_0.OUT.n36 VSS 0.0182f
C771 CM_MSB_V2_0.OUT.n37 VSS 0.06f
C772 CM_MSB_V2_0.OUT.n38 VSS 0.413f
C773 CM_MSB_V2_0.OUT.n39 VSS 0.253f
C774 CM_MSB_V2_0.OUT.n40 VSS 0.244f
C775 CM_MSB_V2_0.OUT.n41 VSS 0.243f
C776 CM_MSB_V2_0.OUT.t37 VSS 0.0182f
C777 CM_MSB_V2_0.OUT.n42 VSS 0.0182f
C778 CM_MSB_V2_0.OUT.n43 VSS 0.0408f
C779 CM_MSB_V2_0.OUT.t131 VSS 0.0182f
C780 CM_MSB_V2_0.OUT.n44 VSS 0.0182f
C781 CM_MSB_V2_0.OUT.n45 VSS 0.0597f
C782 CM_MSB_V2_0.OUT.n46 VSS 0.414f
C783 CM_MSB_V2_0.OUT.n47 VSS 0.253f
C784 CM_MSB_V2_0.OUT.t115 VSS 0.0182f
C785 CM_MSB_V2_0.OUT.n48 VSS 0.0182f
C786 CM_MSB_V2_0.OUT.n49 VSS 0.0363f
C787 CM_MSB_V2_0.OUT.n50 VSS 0.168f
C788 CM_MSB_V2_0.OUT.t55 VSS 0.0182f
C789 CM_MSB_V2_0.OUT.n51 VSS 0.0182f
C790 CM_MSB_V2_0.OUT.n52 VSS 0.0363f
C791 CM_MSB_V2_0.OUT.n53 VSS 0.154f
C792 CM_MSB_V2_0.OUT.n54 VSS 0.228f
C793 CM_MSB_V2_0.OUT.t135 VSS 0.0182f
C794 CM_MSB_V2_0.OUT.n55 VSS 0.0182f
C795 CM_MSB_V2_0.OUT.n56 VSS 0.0363f
C796 CM_MSB_V2_0.OUT.n57 VSS 0.165f
C797 CM_MSB_V2_0.OUT.t39 VSS 0.0182f
C798 CM_MSB_V2_0.OUT.n58 VSS 0.0182f
C799 CM_MSB_V2_0.OUT.n59 VSS 0.0363f
C800 CM_MSB_V2_0.OUT.n60 VSS 0.154f
C801 CM_MSB_V2_0.OUT.n61 VSS 0.228f
C802 CM_MSB_V2_0.OUT.t129 VSS 0.0182f
C803 CM_MSB_V2_0.OUT.n62 VSS 0.0182f
C804 CM_MSB_V2_0.OUT.n63 VSS 0.0363f
C805 CM_MSB_V2_0.OUT.n64 VSS 0.165f
C806 CM_MSB_V2_0.OUT.t58 VSS 0.0182f
C807 CM_MSB_V2_0.OUT.n65 VSS 0.0182f
C808 CM_MSB_V2_0.OUT.n66 VSS 0.0363f
C809 CM_MSB_V2_0.OUT.n67 VSS 0.154f
C810 CM_MSB_V2_0.OUT.n68 VSS 0.228f
C811 CM_MSB_V2_0.OUT.t147 VSS 0.0182f
C812 CM_MSB_V2_0.OUT.n69 VSS 0.0182f
C813 CM_MSB_V2_0.OUT.n70 VSS 0.0363f
C814 CM_MSB_V2_0.OUT.n71 VSS 0.165f
C815 CM_MSB_V2_0.OUT.t63 VSS 0.0182f
C816 CM_MSB_V2_0.OUT.n72 VSS 0.0182f
C817 CM_MSB_V2_0.OUT.n73 VSS 0.0363f
C818 CM_MSB_V2_0.OUT.n74 VSS 0.139f
C819 CM_MSB_V2_0.OUT.t44 VSS 0.0182f
C820 CM_MSB_V2_0.OUT.n75 VSS 0.0182f
C821 CM_MSB_V2_0.OUT.n76 VSS 0.0363f
C822 CM_MSB_V2_0.OUT.n77 VSS 0.168f
C823 CM_MSB_V2_0.OUT.t120 VSS 0.0182f
C824 CM_MSB_V2_0.OUT.n78 VSS 0.0182f
C825 CM_MSB_V2_0.OUT.n79 VSS 0.0363f
C826 CM_MSB_V2_0.OUT.n80 VSS 0.154f
C827 CM_MSB_V2_0.OUT.n81 VSS 0.221f
C828 CM_MSB_V2_0.OUT.t53 VSS 0.0182f
C829 CM_MSB_V2_0.OUT.n82 VSS 0.0182f
C830 CM_MSB_V2_0.OUT.n83 VSS 0.0363f
C831 CM_MSB_V2_0.OUT.n84 VSS 0.165f
C832 CM_MSB_V2_0.OUT.t118 VSS 0.0182f
C833 CM_MSB_V2_0.OUT.n85 VSS 0.0182f
C834 CM_MSB_V2_0.OUT.n86 VSS 0.0363f
C835 CM_MSB_V2_0.OUT.n87 VSS 0.154f
C836 CM_MSB_V2_0.OUT.n88 VSS 0.221f
C837 CM_MSB_V2_0.OUT.t36 VSS 0.0182f
C838 CM_MSB_V2_0.OUT.n89 VSS 0.0182f
C839 CM_MSB_V2_0.OUT.n90 VSS 0.0363f
C840 CM_MSB_V2_0.OUT.n91 VSS 0.165f
C841 CM_MSB_V2_0.OUT.t123 VSS 0.0182f
C842 CM_MSB_V2_0.OUT.n92 VSS 0.0182f
C843 CM_MSB_V2_0.OUT.n93 VSS 0.0363f
C844 CM_MSB_V2_0.OUT.n94 VSS 0.154f
C845 CM_MSB_V2_0.OUT.n95 VSS 0.221f
C846 CM_MSB_V2_0.OUT.t57 VSS 0.0182f
C847 CM_MSB_V2_0.OUT.n96 VSS 0.0182f
C848 CM_MSB_V2_0.OUT.n97 VSS 0.0363f
C849 CM_MSB_V2_0.OUT.n98 VSS 0.165f
C850 CM_MSB_V2_0.OUT.t149 VSS 0.0182f
C851 CM_MSB_V2_0.OUT.n99 VSS 0.0182f
C852 CM_MSB_V2_0.OUT.n100 VSS 0.0363f
C853 CM_MSB_V2_0.OUT.n101 VSS 0.139f
C854 CM_MSB_V2_0.OUT.t86 VSS 0.0182f
C855 CM_MSB_V2_0.OUT.n102 VSS 0.0182f
C856 CM_MSB_V2_0.OUT.n103 VSS 0.0363f
C857 CM_MSB_V2_0.OUT.n104 VSS 0.168f
C858 CM_MSB_V2_0.OUT.t48 VSS 0.0182f
C859 CM_MSB_V2_0.OUT.n105 VSS 0.0182f
C860 CM_MSB_V2_0.OUT.n106 VSS 0.0363f
C861 CM_MSB_V2_0.OUT.n107 VSS 0.154f
C862 CM_MSB_V2_0.OUT.n108 VSS 0.222f
C863 CM_MSB_V2_0.OUT.t137 VSS 0.0182f
C864 CM_MSB_V2_0.OUT.n109 VSS 0.0182f
C865 CM_MSB_V2_0.OUT.n110 VSS 0.0363f
C866 CM_MSB_V2_0.OUT.n111 VSS 0.165f
C867 CM_MSB_V2_0.OUT.t65 VSS 0.0182f
C868 CM_MSB_V2_0.OUT.n112 VSS 0.0182f
C869 CM_MSB_V2_0.OUT.n113 VSS 0.0363f
C870 CM_MSB_V2_0.OUT.n114 VSS 0.154f
C871 CM_MSB_V2_0.OUT.n115 VSS 0.222f
C872 CM_MSB_V2_0.OUT.t104 VSS 0.0182f
C873 CM_MSB_V2_0.OUT.n116 VSS 0.0182f
C874 CM_MSB_V2_0.OUT.n117 VSS 0.0363f
C875 CM_MSB_V2_0.OUT.n118 VSS 0.165f
C876 CM_MSB_V2_0.OUT.t52 VSS 0.0182f
C877 CM_MSB_V2_0.OUT.n119 VSS 0.0182f
C878 CM_MSB_V2_0.OUT.n120 VSS 0.0363f
C879 CM_MSB_V2_0.OUT.n121 VSS 0.154f
C880 CM_MSB_V2_0.OUT.n122 VSS 0.222f
C881 CM_MSB_V2_0.OUT.t111 VSS 0.0182f
C882 CM_MSB_V2_0.OUT.n123 VSS 0.0182f
C883 CM_MSB_V2_0.OUT.n124 VSS 0.0363f
C884 CM_MSB_V2_0.OUT.n125 VSS 0.165f
C885 CM_MSB_V2_0.OUT.t60 VSS 0.0182f
C886 CM_MSB_V2_0.OUT.n126 VSS 0.0182f
C887 CM_MSB_V2_0.OUT.n127 VSS 0.0363f
C888 CM_MSB_V2_0.OUT.n128 VSS 0.139f
C889 CM_MSB_V2_0.OUT.t42 VSS 0.0182f
C890 CM_MSB_V2_0.OUT.n129 VSS 0.0182f
C891 CM_MSB_V2_0.OUT.n130 VSS 0.0387f
C892 CM_MSB_V2_0.OUT.t127 VSS 0.0182f
C893 CM_MSB_V2_0.OUT.n131 VSS 0.0182f
C894 CM_MSB_V2_0.OUT.n132 VSS 0.0567f
C895 CM_MSB_V2_0.OUT.n133 VSS 0.414f
C896 CM_MSB_V2_0.OUT.t49 VSS 0.0182f
C897 CM_MSB_V2_0.OUT.n134 VSS 0.0182f
C898 CM_MSB_V2_0.OUT.n135 VSS 0.0394f
C899 CM_MSB_V2_0.OUT.t128 VSS 0.0182f
C900 CM_MSB_V2_0.OUT.n136 VSS 0.0182f
C901 CM_MSB_V2_0.OUT.n137 VSS 0.0408f
C902 CM_MSB_V2_0.OUT.t144 VSS 0.0182f
C903 CM_MSB_V2_0.OUT.n138 VSS 0.0182f
C904 CM_MSB_V2_0.OUT.n139 VSS 0.0394f
C905 CM_MSB_V2_0.OUT.t40 VSS 0.0182f
C906 CM_MSB_V2_0.OUT.n140 VSS 0.0182f
C907 CM_MSB_V2_0.OUT.n141 VSS 0.0408f
C908 CM_MSB_V2_0.OUT.n142 VSS 0.202f
C909 CM_MSB_V2_0.OUT.n143 VSS 0.259f
C910 CM_MSB_V2_0.OUT.t61 VSS 0.0182f
C911 CM_MSB_V2_0.OUT.n144 VSS 0.0182f
C912 CM_MSB_V2_0.OUT.n145 VSS 0.0394f
C913 CM_MSB_V2_0.OUT.t96 VSS 0.0182f
C914 CM_MSB_V2_0.OUT.n146 VSS 0.0182f
C915 CM_MSB_V2_0.OUT.n147 VSS 0.0408f
C916 CM_MSB_V2_0.OUT.t88 VSS 0.0182f
C917 CM_MSB_V2_0.OUT.n148 VSS 0.0182f
C918 CM_MSB_V2_0.OUT.n149 VSS 0.0394f
C919 CM_MSB_V2_0.OUT.t56 VSS 0.0182f
C920 CM_MSB_V2_0.OUT.n150 VSS 0.0182f
C921 CM_MSB_V2_0.OUT.n151 VSS 0.0408f
C922 CM_MSB_V2_0.OUT.n152 VSS 0.202f
C923 CM_MSB_V2_0.OUT.n153 VSS 0.259f
C924 CM_MSB_V2_0.OUT.t41 VSS 0.0182f
C925 CM_MSB_V2_0.OUT.n154 VSS 0.0182f
C926 CM_MSB_V2_0.OUT.n155 VSS 0.0363f
C927 CM_MSB_V2_0.OUT.n156 VSS 0.168f
C928 CM_MSB_V2_0.OUT.t140 VSS 0.0182f
C929 CM_MSB_V2_0.OUT.n157 VSS 0.0182f
C930 CM_MSB_V2_0.OUT.n158 VSS 0.0363f
C931 CM_MSB_V2_0.OUT.n159 VSS 0.154f
C932 CM_MSB_V2_0.OUT.n160 VSS 0.228f
C933 CM_MSB_V2_0.OUT.t47 VSS 0.0182f
C934 CM_MSB_V2_0.OUT.n161 VSS 0.0182f
C935 CM_MSB_V2_0.OUT.n162 VSS 0.0363f
C936 CM_MSB_V2_0.OUT.n163 VSS 0.165f
C937 CM_MSB_V2_0.OUT.t95 VSS 0.0182f
C938 CM_MSB_V2_0.OUT.n164 VSS 0.0182f
C939 CM_MSB_V2_0.OUT.n165 VSS 0.0363f
C940 CM_MSB_V2_0.OUT.n166 VSS 0.154f
C941 CM_MSB_V2_0.OUT.n167 VSS 0.228f
C942 CM_MSB_V2_0.OUT.t64 VSS 0.0182f
C943 CM_MSB_V2_0.OUT.n168 VSS 0.0182f
C944 CM_MSB_V2_0.OUT.n169 VSS 0.0363f
C945 CM_MSB_V2_0.OUT.n170 VSS 0.165f
C946 CM_MSB_V2_0.OUT.t117 VSS 0.0182f
C947 CM_MSB_V2_0.OUT.n171 VSS 0.0182f
C948 CM_MSB_V2_0.OUT.n172 VSS 0.0363f
C949 CM_MSB_V2_0.OUT.n173 VSS 0.154f
C950 CM_MSB_V2_0.OUT.t132 VSS 0.0182f
C951 CM_MSB_V2_0.OUT.n174 VSS 0.0182f
C952 CM_MSB_V2_0.OUT.n175 VSS 0.0408f
C953 CM_MSB_V2_0.OUT.t151 VSS 0.0182f
C954 CM_MSB_V2_0.OUT.n176 VSS 0.0182f
C955 CM_MSB_V2_0.OUT.n177 VSS 0.0394f
C956 CM_MSB_V2_0.OUT.t59 VSS 0.0182f
C957 CM_MSB_V2_0.OUT.n178 VSS 0.0182f
C958 CM_MSB_V2_0.OUT.n179 VSS 0.0408f
C959 CM_MSB_V2_0.OUT.n180 VSS 0.202f
C960 CM_MSB_V2_0.OUT.t66 VSS 0.0182f
C961 CM_MSB_V2_0.OUT.n181 VSS 0.0182f
C962 CM_MSB_V2_0.OUT.n182 VSS 0.0394f
C963 CM_MSB_V2_0.OUT.n183 VSS 0.259f
C964 CM_MSB_V2_0.OUT.n184 VSS 0.228f
C965 CM_MSB_V2_0.OUT.t51 VSS 0.0182f
C966 CM_MSB_V2_0.OUT.n185 VSS 0.0182f
C967 CM_MSB_V2_0.OUT.n186 VSS 0.0363f
C968 CM_MSB_V2_0.OUT.n187 VSS 0.165f
C969 CM_MSB_V2_0.OUT.t150 VSS 0.0182f
C970 CM_MSB_V2_0.OUT.n188 VSS 0.0182f
C971 CM_MSB_V2_0.OUT.n189 VSS 0.0363f
C972 CM_MSB_V2_0.OUT.n190 VSS 0.139f
C973 CM_MSB_V2_0.OUT.n191 VSS 0.247f
C974 CM_MSB_V2_0.OUT.n192 VSS 0.25f
C975 CM_MSB_V2_0.OUT.n193 VSS 0.249f
C976 CM_MSB_V2_0.OUT.n194 VSS 0.248f
C977 CM_MSB_V2_0.OUT.n195 VSS 0.266f
C978 CM_MSB_V2_0.OUT.n196 VSS 1.24f
C979 CM_MSB_V2_0.OUT.n197 VSS 0.103f
C980 CM_MSB_V2_0.OUT.t156 VSS 0.0363f
C981 CM_MSB_V2_0.OUT.n198 VSS 0.0363f
C982 CM_MSB_V2_0.OUT.n199 VSS 0.0809f
C983 CM_MSB_V2_0.OUT.t4 VSS 0.0363f
C984 CM_MSB_V2_0.OUT.n200 VSS 0.0363f
C985 CM_MSB_V2_0.OUT.n201 VSS 0.0783f
C986 CM_MSB_V2_0.OUT.t0 VSS 0.0363f
C987 CM_MSB_V2_0.OUT.n202 VSS 0.0363f
C988 CM_MSB_V2_0.OUT.n203 VSS 0.0809f
C989 CM_MSB_V2_0.OUT.t103 VSS 0.0363f
C990 CM_MSB_V2_0.OUT.n204 VSS 0.0363f
C991 CM_MSB_V2_0.OUT.n205 VSS 0.0783f
C992 CM_MSB_V2_0.OUT.t10 VSS 0.0363f
C993 CM_MSB_V2_0.OUT.n206 VSS 0.0363f
C994 CM_MSB_V2_0.OUT.n207 VSS 0.0809f
C995 CM_MSB_V2_0.OUT.t14 VSS 0.0363f
C996 CM_MSB_V2_0.OUT.n208 VSS 0.0363f
C997 CM_MSB_V2_0.OUT.n209 VSS 0.0783f
C998 CM_MSB_V2_0.OUT.t85 VSS 0.0363f
C999 CM_MSB_V2_0.OUT.n210 VSS 0.0363f
C1000 CM_MSB_V2_0.OUT.n211 VSS 0.0809f
C1001 CM_MSB_V2_0.OUT.t16 VSS 0.0363f
C1002 CM_MSB_V2_0.OUT.n212 VSS 0.0363f
C1003 CM_MSB_V2_0.OUT.n213 VSS 0.0783f
C1004 CM_MSB_V2_0.OUT.t18 VSS 0.0363f
C1005 CM_MSB_V2_0.OUT.n214 VSS 0.0363f
C1006 CM_MSB_V2_0.OUT.n215 VSS 0.0809f
C1007 CM_MSB_V2_0.OUT.t6 VSS 0.0363f
C1008 CM_MSB_V2_0.OUT.n216 VSS 0.0363f
C1009 CM_MSB_V2_0.OUT.n217 VSS 0.0783f
C1010 CM_MSB_V2_0.OUT.t102 VSS 0.0363f
C1011 CM_MSB_V2_0.OUT.n218 VSS 0.0363f
C1012 CM_MSB_V2_0.OUT.n219 VSS 0.0809f
C1013 CM_MSB_V2_0.OUT.t158 VSS 0.0363f
C1014 CM_MSB_V2_0.OUT.n220 VSS 0.0363f
C1015 CM_MSB_V2_0.OUT.n221 VSS 0.0783f
C1016 CM_MSB_V2_0.OUT.t11 VSS 0.0363f
C1017 CM_MSB_V2_0.OUT.n222 VSS 0.0363f
C1018 CM_MSB_V2_0.OUT.n223 VSS 0.0809f
C1019 CM_MSB_V2_0.OUT.t8 VSS 0.0363f
C1020 CM_MSB_V2_0.OUT.n224 VSS 0.0363f
C1021 CM_MSB_V2_0.OUT.n225 VSS 0.0783f
C1022 CM_MSB_V2_0.OUT.t3 VSS 0.0363f
C1023 CM_MSB_V2_0.OUT.n226 VSS 0.0363f
C1024 CM_MSB_V2_0.OUT.n227 VSS 0.0809f
C1025 CM_MSB_V2_0.OUT.t1 VSS 0.121f
C1026 CM_MSB_V2_0.OUT.n228 VSS 0.435f
C1027 CM_MSB_V2_0.OUT.n229 VSS 0.246f
C1028 CM_MSB_V2_0.OUT.n230 VSS 0.258f
C1029 CM_MSB_V2_0.OUT.n231 VSS 0.246f
C1030 CM_MSB_V2_0.OUT.n232 VSS 0.258f
C1031 CM_MSB_V2_0.OUT.n233 VSS 0.246f
C1032 CM_MSB_V2_0.OUT.n234 VSS 0.258f
C1033 CM_MSB_V2_0.OUT.n235 VSS 0.246f
C1034 CM_MSB_V2_0.OUT.n236 VSS 0.258f
C1035 CM_MSB_V2_0.OUT.n237 VSS 0.246f
C1036 CM_MSB_V2_0.OUT.n238 VSS 0.258f
C1037 CM_MSB_V2_0.OUT.n239 VSS 0.246f
C1038 CM_MSB_V2_0.OUT.n240 VSS 0.258f
C1039 CM_MSB_V2_0.OUT.n241 VSS 0.246f
C1040 CM_MSB_V2_0.OUT.n242 VSS 0.258f
C1041 CM_MSB_V2_0.OUT.n243 VSS 0.242f
C1042 Local_Enc_0.QB.n0 VSS 0.409f
C1043 Local_Enc_0.QB.t68 VSS 0.0123f
C1044 Local_Enc_0.QB.t14 VSS 0.02f
C1045 Local_Enc_0.QB.n1 VSS 0.0569f
C1046 Local_Enc_0.QB.t67 VSS 0.0603f
C1047 Local_Enc_0.QB.t65 VSS 0.0362f
C1048 Local_Enc_0.QB.n2 VSS 0.103f
C1049 Local_Enc_0.QB.t59 VSS 0.0362f
C1050 Local_Enc_0.QB.n3 VSS 0.0684f
C1051 Local_Enc_0.QB.t63 VSS 0.0376f
C1052 Local_Enc_0.QB.n4 VSS 0.0701f
C1053 Local_Enc_0.QB.t28 VSS 0.0376f
C1054 Local_Enc_0.QB.n5 VSS 0.0701f
C1055 Local_Enc_0.QB.t11 VSS 0.0362f
C1056 Local_Enc_0.QB.n6 VSS 0.0684f
C1057 Local_Enc_0.QB.t44 VSS 0.0362f
C1058 Local_Enc_0.QB.n7 VSS 0.0684f
C1059 Local_Enc_0.QB.t9 VSS 0.0376f
C1060 Local_Enc_0.QB.n8 VSS 0.0701f
C1061 Local_Enc_0.QB.t39 VSS 0.0376f
C1062 Local_Enc_0.QB.n9 VSS 0.0701f
C1063 Local_Enc_0.QB.t37 VSS 0.0362f
C1064 Local_Enc_0.QB.n10 VSS 0.0684f
C1065 Local_Enc_0.QB.t54 VSS 0.0362f
C1066 Local_Enc_0.QB.n11 VSS 0.0684f
C1067 Local_Enc_0.QB.t61 VSS 0.0376f
C1068 Local_Enc_0.QB.n12 VSS 0.0701f
C1069 Local_Enc_0.QB.t12 VSS 0.0376f
C1070 Local_Enc_0.QB.n13 VSS 0.0701f
C1071 Local_Enc_0.QB.t10 VSS 0.0362f
C1072 Local_Enc_0.QB.n14 VSS 0.0684f
C1073 Local_Enc_0.QB.t42 VSS 0.0362f
C1074 Local_Enc_0.QB.n15 VSS 0.0755f
C1075 Local_Enc_0.QB.t26 VSS 0.0313f
C1076 Local_Enc_0.QB.n16 VSS 0.0976f
C1077 Local_Enc_0.QB.t29 VSS 0.0603f
C1078 Local_Enc_0.QB.t46 VSS 0.0362f
C1079 Local_Enc_0.QB.n17 VSS 0.103f
C1080 Local_Enc_0.QB.t45 VSS 0.0362f
C1081 Local_Enc_0.QB.n18 VSS 0.0684f
C1082 Local_Enc_0.QB.t23 VSS 0.0376f
C1083 Local_Enc_0.QB.n19 VSS 0.0701f
C1084 Local_Enc_0.QB.t57 VSS 0.0376f
C1085 Local_Enc_0.QB.n20 VSS 0.0701f
C1086 Local_Enc_0.QB.t64 VSS 0.0362f
C1087 Local_Enc_0.QB.n21 VSS 0.0684f
C1088 Local_Enc_0.QB.t30 VSS 0.0362f
C1089 Local_Enc_0.QB.n22 VSS 0.0684f
C1090 Local_Enc_0.QB.t34 VSS 0.0376f
C1091 Local_Enc_0.QB.n23 VSS 0.0701f
C1092 Local_Enc_0.QB.t4 VSS 0.0376f
C1093 Local_Enc_0.QB.n24 VSS 0.0701f
C1094 Local_Enc_0.QB.t24 VSS 0.0362f
C1095 Local_Enc_0.QB.n25 VSS 0.0684f
C1096 Local_Enc_0.QB.t40 VSS 0.0362f
C1097 Local_Enc_0.QB.n26 VSS 0.0684f
C1098 Local_Enc_0.QB.t20 VSS 0.0376f
C1099 Local_Enc_0.QB.n27 VSS 0.0701f
C1100 Local_Enc_0.QB.t38 VSS 0.0376f
C1101 Local_Enc_0.QB.n28 VSS 0.0701f
C1102 Local_Enc_0.QB.t62 VSS 0.0362f
C1103 Local_Enc_0.QB.n29 VSS 0.0684f
C1104 Local_Enc_0.QB.t27 VSS 0.0362f
C1105 Local_Enc_0.QB.n30 VSS 0.0755f
C1106 Local_Enc_0.QB.t55 VSS 0.0313f
C1107 Local_Enc_0.QB.n31 VSS 0.0917f
C1108 Local_Enc_0.QB.t58 VSS 0.0603f
C1109 Local_Enc_0.QB.t13 VSS 0.0362f
C1110 Local_Enc_0.QB.n32 VSS 0.103f
C1111 Local_Enc_0.QB.t8 VSS 0.0362f
C1112 Local_Enc_0.QB.n33 VSS 0.0684f
C1113 Local_Enc_0.QB.t50 VSS 0.0376f
C1114 Local_Enc_0.QB.n34 VSS 0.0701f
C1115 Local_Enc_0.QB.t19 VSS 0.0376f
C1116 Local_Enc_0.QB.n35 VSS 0.0701f
C1117 Local_Enc_0.QB.t25 VSS 0.0362f
C1118 Local_Enc_0.QB.n36 VSS 0.0684f
C1119 Local_Enc_0.QB.t60 VSS 0.0362f
C1120 Local_Enc_0.QB.n37 VSS 0.0684f
C1121 Local_Enc_0.QB.t66 VSS 0.0376f
C1122 Local_Enc_0.QB.n38 VSS 0.0701f
C1123 Local_Enc_0.QB.t31 VSS 0.0376f
C1124 Local_Enc_0.QB.n39 VSS 0.0701f
C1125 Local_Enc_0.QB.t51 VSS 0.0362f
C1126 Local_Enc_0.QB.n40 VSS 0.0684f
C1127 Local_Enc_0.QB.t5 VSS 0.0362f
C1128 Local_Enc_0.QB.n41 VSS 0.0684f
C1129 Local_Enc_0.QB.t47 VSS 0.0376f
C1130 Local_Enc_0.QB.n42 VSS 0.0701f
C1131 Local_Enc_0.QB.t3 VSS 0.0376f
C1132 Local_Enc_0.QB.n43 VSS 0.0701f
C1133 Local_Enc_0.QB.t22 VSS 0.0362f
C1134 Local_Enc_0.QB.n44 VSS 0.0684f
C1135 Local_Enc_0.QB.t56 VSS 0.0362f
C1136 Local_Enc_0.QB.n45 VSS 0.0755f
C1137 Local_Enc_0.QB.t17 VSS 0.0313f
C1138 Local_Enc_0.QB.n46 VSS 0.0917f
C1139 Local_Enc_0.QB.t43 VSS 0.0603f
C1140 Local_Enc_0.QB.t41 VSS 0.0362f
C1141 Local_Enc_0.QB.n47 VSS 0.103f
C1142 Local_Enc_0.QB.t33 VSS 0.0362f
C1143 Local_Enc_0.QB.n48 VSS 0.0684f
C1144 Local_Enc_0.QB.t36 VSS 0.0376f
C1145 Local_Enc_0.QB.n49 VSS 0.0701f
C1146 Local_Enc_0.QB.t6 VSS 0.0376f
C1147 Local_Enc_0.QB.n50 VSS 0.0701f
C1148 Local_Enc_0.QB.t52 VSS 0.0362f
C1149 Local_Enc_0.QB.n51 VSS 0.0684f
C1150 Local_Enc_0.QB.t21 VSS 0.0362f
C1151 Local_Enc_0.QB.n52 VSS 0.0684f
C1152 Local_Enc_0.QB.t48 VSS 0.0376f
C1153 Local_Enc_0.QB.n53 VSS 0.0701f
C1154 Local_Enc_0.QB.t16 VSS 0.0376f
C1155 Local_Enc_0.QB.n54 VSS 0.0701f
C1156 Local_Enc_0.QB.t15 VSS 0.0362f
C1157 Local_Enc_0.QB.n55 VSS 0.0684f
C1158 Local_Enc_0.QB.t32 VSS 0.0362f
C1159 Local_Enc_0.QB.n56 VSS 0.0684f
C1160 Local_Enc_0.QB.t35 VSS 0.0376f
C1161 Local_Enc_0.QB.n57 VSS 0.0701f
C1162 Local_Enc_0.QB.t53 VSS 0.0376f
C1163 Local_Enc_0.QB.n58 VSS 0.0701f
C1164 Local_Enc_0.QB.t49 VSS 0.0362f
C1165 Local_Enc_0.QB.n59 VSS 0.0684f
C1166 Local_Enc_0.QB.t18 VSS 0.0362f
C1167 Local_Enc_0.QB.n60 VSS 0.0755f
C1168 Local_Enc_0.QB.t7 VSS 0.0313f
C1169 Local_Enc_0.QB.n61 VSS 0.101f
C1170 Local_Enc_0.QB.n62 VSS 0.37f
C1171 Local_Enc_0.QB.n63 VSS 0.289f
C1172 Local_Enc_0.QB.n64 VSS 0.00819f
C1173 Local_Enc_0.QB.t1 VSS 0.0289f
.ends

