magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1205 -1794 1205 1794
<< metal2 >>
rect -205 789 205 794
rect -205 761 -200 789
rect -172 761 -138 789
rect -110 761 -76 789
rect -48 761 -14 789
rect 14 761 48 789
rect 76 761 110 789
rect 138 761 172 789
rect 200 761 205 789
rect -205 727 205 761
rect -205 699 -200 727
rect -172 699 -138 727
rect -110 699 -76 727
rect -48 699 -14 727
rect 14 699 48 727
rect 76 699 110 727
rect 138 699 172 727
rect 200 699 205 727
rect -205 665 205 699
rect -205 637 -200 665
rect -172 637 -138 665
rect -110 637 -76 665
rect -48 637 -14 665
rect 14 637 48 665
rect 76 637 110 665
rect 138 637 172 665
rect 200 637 205 665
rect -205 603 205 637
rect -205 575 -200 603
rect -172 575 -138 603
rect -110 575 -76 603
rect -48 575 -14 603
rect 14 575 48 603
rect 76 575 110 603
rect 138 575 172 603
rect 200 575 205 603
rect -205 541 205 575
rect -205 513 -200 541
rect -172 513 -138 541
rect -110 513 -76 541
rect -48 513 -14 541
rect 14 513 48 541
rect 76 513 110 541
rect 138 513 172 541
rect 200 513 205 541
rect -205 479 205 513
rect -205 451 -200 479
rect -172 451 -138 479
rect -110 451 -76 479
rect -48 451 -14 479
rect 14 451 48 479
rect 76 451 110 479
rect 138 451 172 479
rect 200 451 205 479
rect -205 417 205 451
rect -205 389 -200 417
rect -172 389 -138 417
rect -110 389 -76 417
rect -48 389 -14 417
rect 14 389 48 417
rect 76 389 110 417
rect 138 389 172 417
rect 200 389 205 417
rect -205 355 205 389
rect -205 327 -200 355
rect -172 327 -138 355
rect -110 327 -76 355
rect -48 327 -14 355
rect 14 327 48 355
rect 76 327 110 355
rect 138 327 172 355
rect 200 327 205 355
rect -205 293 205 327
rect -205 265 -200 293
rect -172 265 -138 293
rect -110 265 -76 293
rect -48 265 -14 293
rect 14 265 48 293
rect 76 265 110 293
rect 138 265 172 293
rect 200 265 205 293
rect -205 231 205 265
rect -205 203 -200 231
rect -172 203 -138 231
rect -110 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 110 231
rect 138 203 172 231
rect 200 203 205 231
rect -205 169 205 203
rect -205 141 -200 169
rect -172 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 172 169
rect 200 141 205 169
rect -205 107 205 141
rect -205 79 -200 107
rect -172 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 172 107
rect 200 79 205 107
rect -205 45 205 79
rect -205 17 -200 45
rect -172 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 172 45
rect 200 17 205 45
rect -205 -17 205 17
rect -205 -45 -200 -17
rect -172 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 172 -17
rect 200 -45 205 -17
rect -205 -79 205 -45
rect -205 -107 -200 -79
rect -172 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 172 -79
rect 200 -107 205 -79
rect -205 -141 205 -107
rect -205 -169 -200 -141
rect -172 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 172 -141
rect 200 -169 205 -141
rect -205 -203 205 -169
rect -205 -231 -200 -203
rect -172 -231 -138 -203
rect -110 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 110 -203
rect 138 -231 172 -203
rect 200 -231 205 -203
rect -205 -265 205 -231
rect -205 -293 -200 -265
rect -172 -293 -138 -265
rect -110 -293 -76 -265
rect -48 -293 -14 -265
rect 14 -293 48 -265
rect 76 -293 110 -265
rect 138 -293 172 -265
rect 200 -293 205 -265
rect -205 -327 205 -293
rect -205 -355 -200 -327
rect -172 -355 -138 -327
rect -110 -355 -76 -327
rect -48 -355 -14 -327
rect 14 -355 48 -327
rect 76 -355 110 -327
rect 138 -355 172 -327
rect 200 -355 205 -327
rect -205 -389 205 -355
rect -205 -417 -200 -389
rect -172 -417 -138 -389
rect -110 -417 -76 -389
rect -48 -417 -14 -389
rect 14 -417 48 -389
rect 76 -417 110 -389
rect 138 -417 172 -389
rect 200 -417 205 -389
rect -205 -451 205 -417
rect -205 -479 -200 -451
rect -172 -479 -138 -451
rect -110 -479 -76 -451
rect -48 -479 -14 -451
rect 14 -479 48 -451
rect 76 -479 110 -451
rect 138 -479 172 -451
rect 200 -479 205 -451
rect -205 -513 205 -479
rect -205 -541 -200 -513
rect -172 -541 -138 -513
rect -110 -541 -76 -513
rect -48 -541 -14 -513
rect 14 -541 48 -513
rect 76 -541 110 -513
rect 138 -541 172 -513
rect 200 -541 205 -513
rect -205 -575 205 -541
rect -205 -603 -200 -575
rect -172 -603 -138 -575
rect -110 -603 -76 -575
rect -48 -603 -14 -575
rect 14 -603 48 -575
rect 76 -603 110 -575
rect 138 -603 172 -575
rect 200 -603 205 -575
rect -205 -637 205 -603
rect -205 -665 -200 -637
rect -172 -665 -138 -637
rect -110 -665 -76 -637
rect -48 -665 -14 -637
rect 14 -665 48 -637
rect 76 -665 110 -637
rect 138 -665 172 -637
rect 200 -665 205 -637
rect -205 -699 205 -665
rect -205 -727 -200 -699
rect -172 -727 -138 -699
rect -110 -727 -76 -699
rect -48 -727 -14 -699
rect 14 -727 48 -699
rect 76 -727 110 -699
rect 138 -727 172 -699
rect 200 -727 205 -699
rect -205 -761 205 -727
rect -205 -789 -200 -761
rect -172 -789 -138 -761
rect -110 -789 -76 -761
rect -48 -789 -14 -761
rect 14 -789 48 -761
rect 76 -789 110 -761
rect 138 -789 172 -761
rect 200 -789 205 -761
rect -205 -794 205 -789
<< via2 >>
rect -200 761 -172 789
rect -138 761 -110 789
rect -76 761 -48 789
rect -14 761 14 789
rect 48 761 76 789
rect 110 761 138 789
rect 172 761 200 789
rect -200 699 -172 727
rect -138 699 -110 727
rect -76 699 -48 727
rect -14 699 14 727
rect 48 699 76 727
rect 110 699 138 727
rect 172 699 200 727
rect -200 637 -172 665
rect -138 637 -110 665
rect -76 637 -48 665
rect -14 637 14 665
rect 48 637 76 665
rect 110 637 138 665
rect 172 637 200 665
rect -200 575 -172 603
rect -138 575 -110 603
rect -76 575 -48 603
rect -14 575 14 603
rect 48 575 76 603
rect 110 575 138 603
rect 172 575 200 603
rect -200 513 -172 541
rect -138 513 -110 541
rect -76 513 -48 541
rect -14 513 14 541
rect 48 513 76 541
rect 110 513 138 541
rect 172 513 200 541
rect -200 451 -172 479
rect -138 451 -110 479
rect -76 451 -48 479
rect -14 451 14 479
rect 48 451 76 479
rect 110 451 138 479
rect 172 451 200 479
rect -200 389 -172 417
rect -138 389 -110 417
rect -76 389 -48 417
rect -14 389 14 417
rect 48 389 76 417
rect 110 389 138 417
rect 172 389 200 417
rect -200 327 -172 355
rect -138 327 -110 355
rect -76 327 -48 355
rect -14 327 14 355
rect 48 327 76 355
rect 110 327 138 355
rect 172 327 200 355
rect -200 265 -172 293
rect -138 265 -110 293
rect -76 265 -48 293
rect -14 265 14 293
rect 48 265 76 293
rect 110 265 138 293
rect 172 265 200 293
rect -200 203 -172 231
rect -138 203 -110 231
rect -76 203 -48 231
rect -14 203 14 231
rect 48 203 76 231
rect 110 203 138 231
rect 172 203 200 231
rect -200 141 -172 169
rect -138 141 -110 169
rect -76 141 -48 169
rect -14 141 14 169
rect 48 141 76 169
rect 110 141 138 169
rect 172 141 200 169
rect -200 79 -172 107
rect -138 79 -110 107
rect -76 79 -48 107
rect -14 79 14 107
rect 48 79 76 107
rect 110 79 138 107
rect 172 79 200 107
rect -200 17 -172 45
rect -138 17 -110 45
rect -76 17 -48 45
rect -14 17 14 45
rect 48 17 76 45
rect 110 17 138 45
rect 172 17 200 45
rect -200 -45 -172 -17
rect -138 -45 -110 -17
rect -76 -45 -48 -17
rect -14 -45 14 -17
rect 48 -45 76 -17
rect 110 -45 138 -17
rect 172 -45 200 -17
rect -200 -107 -172 -79
rect -138 -107 -110 -79
rect -76 -107 -48 -79
rect -14 -107 14 -79
rect 48 -107 76 -79
rect 110 -107 138 -79
rect 172 -107 200 -79
rect -200 -169 -172 -141
rect -138 -169 -110 -141
rect -76 -169 -48 -141
rect -14 -169 14 -141
rect 48 -169 76 -141
rect 110 -169 138 -141
rect 172 -169 200 -141
rect -200 -231 -172 -203
rect -138 -231 -110 -203
rect -76 -231 -48 -203
rect -14 -231 14 -203
rect 48 -231 76 -203
rect 110 -231 138 -203
rect 172 -231 200 -203
rect -200 -293 -172 -265
rect -138 -293 -110 -265
rect -76 -293 -48 -265
rect -14 -293 14 -265
rect 48 -293 76 -265
rect 110 -293 138 -265
rect 172 -293 200 -265
rect -200 -355 -172 -327
rect -138 -355 -110 -327
rect -76 -355 -48 -327
rect -14 -355 14 -327
rect 48 -355 76 -327
rect 110 -355 138 -327
rect 172 -355 200 -327
rect -200 -417 -172 -389
rect -138 -417 -110 -389
rect -76 -417 -48 -389
rect -14 -417 14 -389
rect 48 -417 76 -389
rect 110 -417 138 -389
rect 172 -417 200 -389
rect -200 -479 -172 -451
rect -138 -479 -110 -451
rect -76 -479 -48 -451
rect -14 -479 14 -451
rect 48 -479 76 -451
rect 110 -479 138 -451
rect 172 -479 200 -451
rect -200 -541 -172 -513
rect -138 -541 -110 -513
rect -76 -541 -48 -513
rect -14 -541 14 -513
rect 48 -541 76 -513
rect 110 -541 138 -513
rect 172 -541 200 -513
rect -200 -603 -172 -575
rect -138 -603 -110 -575
rect -76 -603 -48 -575
rect -14 -603 14 -575
rect 48 -603 76 -575
rect 110 -603 138 -575
rect 172 -603 200 -575
rect -200 -665 -172 -637
rect -138 -665 -110 -637
rect -76 -665 -48 -637
rect -14 -665 14 -637
rect 48 -665 76 -637
rect 110 -665 138 -637
rect 172 -665 200 -637
rect -200 -727 -172 -699
rect -138 -727 -110 -699
rect -76 -727 -48 -699
rect -14 -727 14 -699
rect 48 -727 76 -699
rect 110 -727 138 -699
rect 172 -727 200 -699
rect -200 -789 -172 -761
rect -138 -789 -110 -761
rect -76 -789 -48 -761
rect -14 -789 14 -761
rect 48 -789 76 -761
rect 110 -789 138 -761
rect 172 -789 200 -761
<< metal3 >>
rect -205 789 205 794
rect -205 761 -200 789
rect -172 761 -138 789
rect -110 761 -76 789
rect -48 761 -14 789
rect 14 761 48 789
rect 76 761 110 789
rect 138 761 172 789
rect 200 761 205 789
rect -205 727 205 761
rect -205 699 -200 727
rect -172 699 -138 727
rect -110 699 -76 727
rect -48 699 -14 727
rect 14 699 48 727
rect 76 699 110 727
rect 138 699 172 727
rect 200 699 205 727
rect -205 665 205 699
rect -205 637 -200 665
rect -172 637 -138 665
rect -110 637 -76 665
rect -48 637 -14 665
rect 14 637 48 665
rect 76 637 110 665
rect 138 637 172 665
rect 200 637 205 665
rect -205 603 205 637
rect -205 575 -200 603
rect -172 575 -138 603
rect -110 575 -76 603
rect -48 575 -14 603
rect 14 575 48 603
rect 76 575 110 603
rect 138 575 172 603
rect 200 575 205 603
rect -205 541 205 575
rect -205 513 -200 541
rect -172 513 -138 541
rect -110 513 -76 541
rect -48 513 -14 541
rect 14 513 48 541
rect 76 513 110 541
rect 138 513 172 541
rect 200 513 205 541
rect -205 479 205 513
rect -205 451 -200 479
rect -172 451 -138 479
rect -110 451 -76 479
rect -48 451 -14 479
rect 14 451 48 479
rect 76 451 110 479
rect 138 451 172 479
rect 200 451 205 479
rect -205 417 205 451
rect -205 389 -200 417
rect -172 389 -138 417
rect -110 389 -76 417
rect -48 389 -14 417
rect 14 389 48 417
rect 76 389 110 417
rect 138 389 172 417
rect 200 389 205 417
rect -205 355 205 389
rect -205 327 -200 355
rect -172 327 -138 355
rect -110 327 -76 355
rect -48 327 -14 355
rect 14 327 48 355
rect 76 327 110 355
rect 138 327 172 355
rect 200 327 205 355
rect -205 293 205 327
rect -205 265 -200 293
rect -172 265 -138 293
rect -110 265 -76 293
rect -48 265 -14 293
rect 14 265 48 293
rect 76 265 110 293
rect 138 265 172 293
rect 200 265 205 293
rect -205 231 205 265
rect -205 203 -200 231
rect -172 203 -138 231
rect -110 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 110 231
rect 138 203 172 231
rect 200 203 205 231
rect -205 169 205 203
rect -205 141 -200 169
rect -172 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 172 169
rect 200 141 205 169
rect -205 107 205 141
rect -205 79 -200 107
rect -172 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 172 107
rect 200 79 205 107
rect -205 45 205 79
rect -205 17 -200 45
rect -172 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 172 45
rect 200 17 205 45
rect -205 -17 205 17
rect -205 -45 -200 -17
rect -172 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 172 -17
rect 200 -45 205 -17
rect -205 -79 205 -45
rect -205 -107 -200 -79
rect -172 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 172 -79
rect 200 -107 205 -79
rect -205 -141 205 -107
rect -205 -169 -200 -141
rect -172 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 172 -141
rect 200 -169 205 -141
rect -205 -203 205 -169
rect -205 -231 -200 -203
rect -172 -231 -138 -203
rect -110 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 110 -203
rect 138 -231 172 -203
rect 200 -231 205 -203
rect -205 -265 205 -231
rect -205 -293 -200 -265
rect -172 -293 -138 -265
rect -110 -293 -76 -265
rect -48 -293 -14 -265
rect 14 -293 48 -265
rect 76 -293 110 -265
rect 138 -293 172 -265
rect 200 -293 205 -265
rect -205 -327 205 -293
rect -205 -355 -200 -327
rect -172 -355 -138 -327
rect -110 -355 -76 -327
rect -48 -355 -14 -327
rect 14 -355 48 -327
rect 76 -355 110 -327
rect 138 -355 172 -327
rect 200 -355 205 -327
rect -205 -389 205 -355
rect -205 -417 -200 -389
rect -172 -417 -138 -389
rect -110 -417 -76 -389
rect -48 -417 -14 -389
rect 14 -417 48 -389
rect 76 -417 110 -389
rect 138 -417 172 -389
rect 200 -417 205 -389
rect -205 -451 205 -417
rect -205 -479 -200 -451
rect -172 -479 -138 -451
rect -110 -479 -76 -451
rect -48 -479 -14 -451
rect 14 -479 48 -451
rect 76 -479 110 -451
rect 138 -479 172 -451
rect 200 -479 205 -451
rect -205 -513 205 -479
rect -205 -541 -200 -513
rect -172 -541 -138 -513
rect -110 -541 -76 -513
rect -48 -541 -14 -513
rect 14 -541 48 -513
rect 76 -541 110 -513
rect 138 -541 172 -513
rect 200 -541 205 -513
rect -205 -575 205 -541
rect -205 -603 -200 -575
rect -172 -603 -138 -575
rect -110 -603 -76 -575
rect -48 -603 -14 -575
rect 14 -603 48 -575
rect 76 -603 110 -575
rect 138 -603 172 -575
rect 200 -603 205 -575
rect -205 -637 205 -603
rect -205 -665 -200 -637
rect -172 -665 -138 -637
rect -110 -665 -76 -637
rect -48 -665 -14 -637
rect 14 -665 48 -637
rect 76 -665 110 -637
rect 138 -665 172 -637
rect 200 -665 205 -637
rect -205 -699 205 -665
rect -205 -727 -200 -699
rect -172 -727 -138 -699
rect -110 -727 -76 -699
rect -48 -727 -14 -699
rect 14 -727 48 -699
rect 76 -727 110 -699
rect 138 -727 172 -699
rect 200 -727 205 -699
rect -205 -761 205 -727
rect -205 -789 -200 -761
rect -172 -789 -138 -761
rect -110 -789 -76 -761
rect -48 -789 -14 -761
rect 14 -789 48 -761
rect 76 -789 110 -761
rect 138 -789 172 -761
rect 200 -789 205 -761
rect -205 -794 205 -789
<< end >>
