* NGSPICE file created from RES_74k.ext - technology: gf180mcuD

.subckt ppolyf_u_DTYK2C a_n1010_n2224# a_n1010_n362# a_n1310_n2846# a_n2210_2744#
+ a_n1610_n1396# a_1390_1294# a_490_1916# a_n1610_n568# a_1690_1088# a_1090_2122#
+ a_n1610_n2018# a_2290_n1190# a_n710_1916# a_190_n2846# a_2290_1294# a_n2210_n1396#
+ a_n2510_n568# a_490_n1396# a_n710_n1190# a_n110_2744# a_n1310_1294# a_n2210_n2018#
+ a_490_n2018# a_1390_n1190# a_n1610_1088# a_n1010_2122# a_190_n568# a_1690_1916#
+ a_n1010_n2846# a_2290_466# a_n2510_466# a_n1310_n1396# a_1990_260# a_n2210_1294#
+ a_n410_n568# a_n2510_1088# a_1090_2744# a_n1310_n2018# a_1690_466# a_n1910_466#
+ a_790_n362# a_1990_n2224# a_n2210_260# a_190_n1396# a_n410_n1190# a_190_1088# a_n1610_1916#
+ a_n110_1294# a_1390_n568# a_1390_260# a_n1610_260# a_190_n2018# a_1090_n1190# a_n410_1088#
+ a_n1010_2744# a_1090_466# a_n1310_466# a_n2510_1916# a_n1010_n1396# a_2290_n568#
+ a_1990_n362# a_n1010_n2018# a_1090_1294# a_790_2122# a_n1310_n568# a_190_1916# a_n1010_260#
+ a_1390_1088# a_1690_n2224# a_1990_n2846# a_790_260# a_n110_n1190# a_n410_1916# a_n710_466#
+ a_490_466# a_n2210_n568# a_n1910_n362# a_2290_1088# a_2290_n2224# a_n1010_1294#
+ a_n1310_1088# a_n410_260# a_1990_2122# a_n710_n2224# a_190_260# a_1390_1916# a_n110_n568#
+ a_n110_466# a_790_2744# a_1390_n2224# a_1690_n2846# a_n2210_1088# a_1990_n1396#
+ a_490_n362# a_2290_1916# a_n1910_2122# a_n1310_1916# a_1990_n2018# a_n710_n362#
+ a_2290_n2846# a_1090_n568# a_n1910_n1190# a_n110_1088# a_n410_n2224# a_1990_2744#
+ a_n710_n2846# a_n2210_1916# a_790_1294# a_1090_n2224# a_1390_n2846# a_n2510_n1190#
+ a_1690_n362# a_790_n1190# a_490_2122# a_1690_n1396# a_n1010_n568# a_1090_1088# a_n710_2122#
+ a_n110_1916# a_n1910_2744# a_1690_n2018# a_2290_n1396# a_n1610_n1190# a_n1610_n362#
+ a_n110_n2224# a_n410_n2846# a_1990_1294# a_n710_n1396# a_2290_n2018# a_n1010_1088#
+ a_1690_2122# a_1090_n2846# a_n2210_n1190# a_1090_1916# a_490_n1190# a_n2510_n362#
+ a_490_2744# a_n710_n2018# a_1390_n1396# a_1990_466# a_n710_2744# a_1390_n2018# a_n1910_1294#
+ a_2290_260# a_190_n362# a_n2510_260# a_n1610_2122# a_n1310_n1190# a_n410_n362# a_n1010_1916#
+ a_790_n568# a_n110_n2846# a_1690_260# a_n2210_466# a_n410_n1396# a_n1910_260# a_1690_2744#
+ a_1390_466# a_n2510_2122# a_190_n1190# a_n1610_466# a_n410_n2018# a_1090_n1396#
+ a_n1910_n2224# a_490_1294# a_1390_n362# a_790_1088# a_1090_n2018# a_n710_1294# a_190_2122#
+ a_1090_260# a_1990_n568# a_n1310_260# a_n410_2122# a_n1010_n1190# a_n1610_2744#
+ a_n2510_n2224# a_2290_n362# a_790_n2224# a_n1010_466# a_n110_n1396# a_790_466# a_n1310_n362#
+ a_n2510_2744# a_1690_1294# a_n110_n2018# a_n1910_n568# a_1990_1088# a_790_1916#
+ a_n1910_n2846# a_n1610_n2224# a_n710_260# a_1390_2122# a_490_260# a_n2210_n362#
+ a_190_2744# a_n410_466# a_190_466# a_2290_2122# a_n410_2744# a_n2510_n2846# a_n2210_n2224#
+ a_n1610_1294# a_490_n2224# a_790_n2846# a_n1910_1088# a_n1310_2122# a_490_n568#
+ a_n110_n362# a_n110_260# a_1990_1916# a_1990_n1190# a_n710_n568# a_n2510_1294# a_n1610_n2846#
+ a_n1310_n2224# a_1390_2744# a_n2210_2122# a_n1910_n1396# a_190_1294# a_n1910_n2018#
+ a_1090_n362# a_490_1088# a_n1910_1916# a_n2210_n2846# a_n410_1294# a_2290_2744#
+ a_190_n2224# a_490_n2846# a_1690_n568# a_790_n1396# a_n2510_n1396# a_n710_1088#
+ a_n110_2122# a_n1310_2744# a_n2510_n2018# a_790_n2018# a_1690_n1190#
X0 a_2290_1088# a_2290_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X1 a_n1010_1916# a_n1010_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X2 a_n1610_n568# a_n1610_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X3 a_n2210_n2224# a_n2210_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X4 a_n1310_2744# a_n1310_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X5 a_1690_n2224# a_1690_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X6 a_790_n2224# a_790_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X7 a_n2210_n1396# a_n2210_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X8 a_1690_n1396# a_1690_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X9 a_1690_1088# a_1690_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X10 a_790_n1396# a_790_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X11 a_2290_1916# a_2290_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X12 a_n110_n2224# a_n110_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X13 a_n2510_n568# a_n2510_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X14 a_1990_n568# a_1990_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X15 a_790_260# a_790_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X16 a_n110_n1396# a_n110_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X17 a_n410_260# a_n410_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X18 a_n410_n568# a_n410_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X19 a_490_1916# a_490_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X20 a_790_2744# a_790_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X21 a_n2210_260# a_n2210_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X22 a_1990_260# a_1990_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X23 a_n110_1916# a_n110_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X24 a_1990_1088# a_1990_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X25 a_n410_2744# a_n410_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X26 a_n2210_2744# a_n2210_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X27 a_1690_1916# a_1690_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X28 a_1990_2744# a_1990_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X29 a_n1010_n2224# a_n1010_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X30 a_n1010_n1396# a_n1010_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X31 a_n1610_260# a_n1610_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X32 a_n1310_n568# a_n1310_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X33 a_n1310_1916# a_n1310_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X34 a_n1610_2744# a_n1610_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X35 a_1390_n2224# a_1390_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X36 a_490_n2224# a_490_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X37 a_1390_n1396# a_1390_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X38 a_490_n1396# a_490_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X39 a_1090_260# a_1090_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X40 a_n2210_n568# a_n2210_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X41 a_1690_n568# a_1690_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X42 a_790_n568# a_790_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X43 a_1090_2744# a_1090_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X44 a_2290_n2224# a_2290_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X45 a_n710_260# a_n710_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X46 a_2290_n1396# a_2290_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X47 a_790_1916# a_790_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X48 a_n110_n568# a_n110_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X49 a_n2510_260# a_n2510_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X50 a_n1910_n2224# a_n1910_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X51 a_n410_1916# a_n410_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X52 a_n710_2744# a_n710_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X53 a_n1910_n1396# a_n1910_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X54 a_n110_1088# a_n110_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X55 a_n2210_1916# a_n2210_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X56 a_n2510_2744# a_n2510_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X57 a_1990_1916# a_1990_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X58 a_190_1088# a_190_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X59 a_n710_n2224# a_n710_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X60 a_n1910_260# a_n1910_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X61 a_n410_1088# a_n410_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X62 a_n710_n1396# a_n710_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X63 a_190_260# a_190_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X64 a_n1010_n568# a_n1010_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X65 a_n1610_1916# a_n1610_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X66 a_490_1088# a_490_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X67 a_n1910_2744# a_n1910_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X68 a_1090_n2224# a_1090_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X69 a_190_n2224# a_190_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X70 a_190_2744# a_190_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X71 a_1090_n1396# a_1090_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X72 a_190_n1396# a_190_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X73 a_1390_260# a_1390_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X74 a_1390_n568# a_1390_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X75 a_1090_1916# a_1090_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X76 a_490_n568# a_490_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X77 a_n710_1088# a_n710_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X78 a_1390_2744# a_1390_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X79 a_790_1088# a_790_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X80 a_n1010_1088# a_n1010_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X81 a_n1610_n2224# a_n1610_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X82 a_n710_1916# a_n710_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X83 a_n1610_n1396# a_n1610_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X84 a_2290_n568# a_2290_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X85 a_n2510_1916# a_n2510_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X86 a_n1010_260# a_n1010_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X87 a_n1910_n568# a_n1910_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X88 a_n1010_2744# a_n1010_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X89 a_1990_n2224# a_1990_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X90 a_n2510_n2224# a_n2510_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X91 a_2290_260# a_2290_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X92 a_n1310_1088# a_n1310_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X93 a_n2510_n1396# a_n2510_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X94 a_1990_n1396# a_1990_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X95 a_n410_n2224# a_n410_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X96 a_2290_2744# a_2290_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X97 a_n410_n1396# a_n410_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X98 a_490_260# a_490_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X99 a_n1910_1916# a_n1910_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X100 a_n2210_1088# a_n2210_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X101 a_n110_260# a_n110_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X102 a_n710_n568# a_n710_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X103 a_1090_1088# a_1090_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X104 a_190_1916# a_190_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X105 a_490_2744# a_490_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X106 a_1690_260# a_1690_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X107 a_n1610_1088# a_n1610_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X108 a_n110_2744# a_n110_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X109 a_1090_n568# a_1090_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X110 a_1390_1916# a_1390_1294# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X111 a_190_n568# a_190_n1190# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X112 a_1690_2744# a_1690_2122# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X113 a_n2510_1088# a_n2510_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X114 a_1390_1088# a_1390_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X115 a_n1310_n2224# a_n1310_n2846# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X116 a_n1310_n1396# a_n1310_n2018# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X117 a_n1910_1088# a_n1910_466# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
X118 a_n1310_260# a_n1310_n362# w_n2726_n3062# ppolyf_u r_width=1.1u r_length=2.6u
.ends

.subckt RES_74k P M
Xppolyf_u_DTYK2C_0 m1_4088_n925# m1_5588_1559# m1_4088_n925# m1_4088_n925# m1_4688_555#
+ m1_7988_3215# m1_7088_3867# m1_4988_1383# m1_7988_3039# m1_4088_n925# m1_4988_n97#
+ m1_4088_n925# m1_5888_3867# m1_4088_n925# m1_4088_n925# a_4386_614# m1_4088_n925#
+ m1_7088_555# m1_5888_731# m1_4088_n925# m1_4988_3215# m1_4388_n97# m1_6788_n97#
+ m1_7688_731# m1_4988_3039# m1_4088_n925# m1_6788_1383# m1_8288_3867# m1_4088_n925#
+ m1_4088_n925# m1_4088_n925# m1_5288_555# m1_8288_2211# m1_4388_3215# m1_6188_1383#
+ m1_4088_n925# m1_4088_n925# m1_4988_n97# m1_8288_2387# m1_4688_2387# m1_7388_1559#
+ m1_4088_n925# a_4386_2270# m1_6488_555# m1_5888_731# m1_6788_3039# m1_4688_3867#
+ m1_6188_3215# m1_7988_1383# m1_7688_2211# m1_4688_2211# m1_6788_n97# m1_7688_731#
+ m1_6188_3039# m1_4088_n925# m1_7688_2387# m1_5288_2387# m1_4088_n925# m1_5288_555#
+ m1_4088_n925# a_8586_1442# m1_5588_n97# m1_7388_3215# m1_4088_n925# m1_4988_1383#
+ m1_6488_3867# m1_5288_2211# m1_7988_3039# m1_4088_n925# m1_4088_n925# m1_7088_2211#
+ m1_6488_731# m1_5888_3867# m1_5888_2387# m1_7088_2387# m1_4388_1383# m1_4388_1559#
+ m1_4088_n925# m1_4088_n925# m1_5588_3215# m1_4988_3039# m1_5888_2211# m1_4088_n925#
+ m1_4088_n925# m1_6488_2211# m1_7688_3867# m1_6188_1383# m1_6488_2387# m1_4088_n925#
+ m1_4088_n925# m1_4088_n925# m1_4388_3039# m1_8288_555# m1_6788_1559# m1_4088_n925#
+ m1_4088_n925# m1_5288_3867# M m1_5588_1559# m1_4088_n925# m1_7388_1383# m1_4688_731#
+ m1_6188_3039# m1_4088_n925# m1_4088_n925# m1_4088_n925# P m1_7388_3215# m1_4088_n925#
+ m1_4088_n925# m1_4088_n925# m1_7988_1559# m1_7088_731# m1_4088_n925# m1_8288_555#
+ m1_5588_1383# m1_7388_3039# m1_4088_n925# m1_6488_3867# m1_4088_n925# m1_7988_n97#
+ m1_4088_n925# m1_4688_731# m1_4988_1559# m1_4088_n925# m1_4088_n925# a_8586_3098#
+ m1_5888_555# m1_4088_n925# m1_5588_3039# m1_4088_n925# m1_4088_n925# a_4386_614#
+ m1_7688_3867# m1_7088_731# m1_4088_n925# m1_4088_n925# m1_5588_n97# m1_7688_555#
+ m1_8288_2387# m1_4088_n925# m1_7988_n97# m1_4388_3215# m1_4088_n925# m1_6788_1559#
+ m1_4088_n925# m1_4088_n925# m1_5288_731# m1_6188_1559# m1_5288_3867# m1_7388_1383#
+ m1_4088_n925# m1_8288_2211# a_4386_2270# m1_5888_555# m1_4688_2211# m1_4088_n925#
+ m1_7688_2387# m1_4088_n925# m1_6488_731# m1_4688_2387# m1_6188_n97# m1_7688_555#
+ m1_4088_n925# m1_6788_3215# m1_7988_1559# m1_7388_3039# m1_7388_n97# m1_5588_3215#
+ m1_4088_n925# m1_7688_2211# a_8586_1442# m1_5288_2211# m1_4088_n925# m1_5288_731#
+ m1_4088_n925# m1_4088_n925# m1_4088_n925# m1_4088_n925# m1_5288_2387# m1_6488_555#
+ m1_7088_2387# m1_4988_1559# m1_4088_n925# m1_7988_3215# m1_6188_n97# m1_4388_1383#
+ a_8586_3098# m1_7088_3867# m1_4088_n925# m1_4088_n925# m1_5888_2211# m1_4088_n925#
+ m1_7088_2211# m1_4388_1559# m1_4088_n925# m1_5888_2387# m1_6488_2387# m1_4088_n925#
+ m1_4088_n925# m1_4088_n925# m1_4088_n925# m1_4988_3215# m1_4088_n925# m1_4088_n925#
+ m1_4388_3039# m1_4088_n925# m1_6788_1383# m1_6188_1559# m1_6488_2211# m1_8288_3867#
+ m1_8288_731# m1_5588_1383# m1_4088_n925# m1_4088_n925# m1_4088_n925# m1_4088_n925#
+ m1_4088_n925# m1_4688_555# m1_6788_3215# m1_4388_n97# m1_7388_1559# m1_6788_3039#
+ m1_4688_3867# m1_4088_n925# m1_6188_3215# m1_4088_n925# m1_4088_n925# m1_4088_n925#
+ m1_7988_1383# m1_7088_555# m1_4088_n925# m1_5588_3039# m1_4088_n925# m1_4088_n925#
+ m1_4088_n925# m1_7388_n97# m1_8288_731# ppolyf_u_DTYK2C
.ends

