** sch_path: /home/shahid/Videos/AWG_MUX/mux/1x8_MUX/xschem/PEX_1x8_TB.sch
**.subckt PEX_1x8_TB
V4 VSS GND 0
.save i(v4)
V5 VDD VSS 3.3
.save i(v5)
V2 A0 VSS 50m
.save i(v2)
V3 A1 VSS 100m
.save i(v3)
V6 A2 VSS 200m
.save i(v6)
V7 A3 VSS 300m
.save i(v7)
V8 A4 VSS 400m
.save i(v8)
V9 A5 VSS 500m
.save i(v9)
V10 A6 VSS 600m
.save i(v10)
V11 A7 VSS 700m
.save i(v11)
V12 net1 VSS (pulse(0 3.3 0 10p 10p 4u 8u))
.save i(v12)
V13 net2 VSS (pulse(0 3.3 0 10p 10p 2u 4u))
.save i(v13)
V14 net3 VSS (pulse(0 3.3 0 10p 10p 1u 2u))
.save i(v14)
V1 ENA VSS 3.3
.save i(v1)
V15 S2 VSS 3
.save i(v15)
V16 S1 VSS 3
.save i(v16)
V17 S0 VSS 3
.save i(v17)
C1 net4 net5 1p m=1
x1 VDD Vout VSS A0 A1 A2 A3 A4 A5 A6 A7 S0 S1 S2 ENA pex_MUX_1x8
R1 Vout VSS 10k m=1
**** begin user architecture code

.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical



.include pex_MUX_1x8.spice
.control
*set color0=white
*set color1=black
save all

tran 1u 16u
plot v(S0) v(S1) v(S2)
plot v(A0) v(A1) v(A2)
Plot v(Vout)

.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
