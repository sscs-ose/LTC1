* NGSPICE file created from resistor_PGA_flat.ext - technology: gf180mcuC

.subckt resistor_PGA_flat
X0 a_7116_765.t0 a_6476_105.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X1 a_5836_1123.t1 a_7116_n857.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X2 a_6476_105.t0 a_6156_n197.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X3 a_5516_1123.t1 a_5836_n197.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X4 a_5516_n555.t1 a_5516_n857.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X5 a_6156_1425.t0 a_6476_1123.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X6 a_6476_463.t1 a_7116_n197.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X7 a_6796_n555.t1 a_5836_n857.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X8 a_6156_765.t1 a_5516_105.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X9 a_5516_765.t0 a_5516_463.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X10 a_6476_1123.t0 a_6796_463.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X11 a_5516_463.t0 a_6156_n197.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X12 a_5516_105.t0 a_5516_n197.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X13 a_5836_1425.t0 a_5836_1123.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X14 a_6156_1425.t1 a_6156_1123.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X15 a_6476_n555.t0 a_6156_n857.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X16 a_6796_105.t0 a_5836_n197.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X17 a_7116_1425.t0 a_6796_1123.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X18 a_6156_765.t0 a_6476_463.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X19 a_5516_1425.t0 a_5516_1123.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X20 a_6796_n555.t0 a_6796_1123.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X21 a_5516_n555.t0 a_5836_n857.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X22 a_5836_463.t1 a_6156_n857.t1 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
X23 a_5836_765.t0 a_5836_463.t0 w_5332_n1041# ppolyf_u r_width=1.2u r_length=1u
R0 a_6476_105.t0 a_6476_105.t1 10.6182
R1 a_5836_1123.t0 a_5836_1123.t1 12.2906
R2 a_6156_n197.t0 a_6156_n197.t1 12.3428
R3 a_5516_1123.t0 a_5516_1123.t1 8.82204
R4 a_5836_n197.t0 a_5836_n197.t1 13.0784
R5 a_5516_n555.t0 a_5516_n555.t1 12.3428
R6 a_6156_1425.t0 a_6156_1425.t1 12.3428
R7 a_6476_1123.t0 a_6476_1123.t1 12.5114
R8 a_6476_463.t0 a_6476_463.t1 8.27632
R9 a_6796_n555.t0 a_6796_n555.t1 11.5186
R10 a_5836_n857.t0 a_5836_n857.t1 12.8783
R11 a_6156_765.t0 a_6156_765.t1 12.3428
R12 a_5516_105.t0 a_5516_105.t1 12.7742
R13 a_5516_463.t0 a_5516_463.t1 8.39738
R14 a_6156_n857.t0 a_6156_n857.t1 12.3428
R15 a_6796_1123.t0 a_6796_1123.t1 12.3428
R16 a_5836_463.t0 a_5836_463.t1 10.6249
C0 m1_4783_490# m1_4778_733# 0.116f
C1 w_5332_n1041# m1_4778_733# 0.00303f
C2 w_5332_n1041# m1_4783_490# 0.00701f
C3 w_5332_n1041# m1_4677_n319# 0.00496f
C4 m1_4677_n319# VSUBS 0.0992f $ **FLOATING
C5 m1_4783_490# VSUBS 0.239f $ **FLOATING
C6 m1_4778_733# VSUBS 0.159f $ **FLOATING
C7 w_5332_n1041# VSUBS 18.2f
.ends

