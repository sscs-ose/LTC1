magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1247 -1551 1247 1551
<< metal1 >>
rect -247 545 247 551
rect -247 519 -241 545
rect -215 519 -165 545
rect -139 519 -89 545
rect -63 519 -13 545
rect 13 519 63 545
rect 89 519 139 545
rect 165 519 215 545
rect 241 519 247 545
rect -247 469 247 519
rect -247 443 -241 469
rect -215 443 -165 469
rect -139 443 -89 469
rect -63 443 -13 469
rect 13 443 63 469
rect 89 443 139 469
rect 165 443 215 469
rect 241 443 247 469
rect -247 393 247 443
rect -247 367 -241 393
rect -215 367 -165 393
rect -139 367 -89 393
rect -63 367 -13 393
rect 13 367 63 393
rect 89 367 139 393
rect 165 367 215 393
rect 241 367 247 393
rect -247 317 247 367
rect -247 291 -241 317
rect -215 291 -165 317
rect -139 291 -89 317
rect -63 291 -13 317
rect 13 291 63 317
rect 89 291 139 317
rect 165 291 215 317
rect 241 291 247 317
rect -247 241 247 291
rect -247 215 -241 241
rect -215 215 -165 241
rect -139 215 -89 241
rect -63 215 -13 241
rect 13 215 63 241
rect 89 215 139 241
rect 165 215 215 241
rect 241 215 247 241
rect -247 165 247 215
rect -247 139 -241 165
rect -215 139 -165 165
rect -139 139 -89 165
rect -63 139 -13 165
rect 13 139 63 165
rect 89 139 139 165
rect 165 139 215 165
rect 241 139 247 165
rect -247 89 247 139
rect -247 63 -241 89
rect -215 63 -165 89
rect -139 63 -89 89
rect -63 63 -13 89
rect 13 63 63 89
rect 89 63 139 89
rect 165 63 215 89
rect 241 63 247 89
rect -247 13 247 63
rect -247 -13 -241 13
rect -215 -13 -165 13
rect -139 -13 -89 13
rect -63 -13 -13 13
rect 13 -13 63 13
rect 89 -13 139 13
rect 165 -13 215 13
rect 241 -13 247 13
rect -247 -63 247 -13
rect -247 -89 -241 -63
rect -215 -89 -165 -63
rect -139 -89 -89 -63
rect -63 -89 -13 -63
rect 13 -89 63 -63
rect 89 -89 139 -63
rect 165 -89 215 -63
rect 241 -89 247 -63
rect -247 -139 247 -89
rect -247 -165 -241 -139
rect -215 -165 -165 -139
rect -139 -165 -89 -139
rect -63 -165 -13 -139
rect 13 -165 63 -139
rect 89 -165 139 -139
rect 165 -165 215 -139
rect 241 -165 247 -139
rect -247 -215 247 -165
rect -247 -241 -241 -215
rect -215 -241 -165 -215
rect -139 -241 -89 -215
rect -63 -241 -13 -215
rect 13 -241 63 -215
rect 89 -241 139 -215
rect 165 -241 215 -215
rect 241 -241 247 -215
rect -247 -291 247 -241
rect -247 -317 -241 -291
rect -215 -317 -165 -291
rect -139 -317 -89 -291
rect -63 -317 -13 -291
rect 13 -317 63 -291
rect 89 -317 139 -291
rect 165 -317 215 -291
rect 241 -317 247 -291
rect -247 -367 247 -317
rect -247 -393 -241 -367
rect -215 -393 -165 -367
rect -139 -393 -89 -367
rect -63 -393 -13 -367
rect 13 -393 63 -367
rect 89 -393 139 -367
rect 165 -393 215 -367
rect 241 -393 247 -367
rect -247 -443 247 -393
rect -247 -469 -241 -443
rect -215 -469 -165 -443
rect -139 -469 -89 -443
rect -63 -469 -13 -443
rect 13 -469 63 -443
rect 89 -469 139 -443
rect 165 -469 215 -443
rect 241 -469 247 -443
rect -247 -519 247 -469
rect -247 -545 -241 -519
rect -215 -545 -165 -519
rect -139 -545 -89 -519
rect -63 -545 -13 -519
rect 13 -545 63 -519
rect 89 -545 139 -519
rect 165 -545 215 -519
rect 241 -545 247 -519
rect -247 -551 247 -545
<< via1 >>
rect -241 519 -215 545
rect -165 519 -139 545
rect -89 519 -63 545
rect -13 519 13 545
rect 63 519 89 545
rect 139 519 165 545
rect 215 519 241 545
rect -241 443 -215 469
rect -165 443 -139 469
rect -89 443 -63 469
rect -13 443 13 469
rect 63 443 89 469
rect 139 443 165 469
rect 215 443 241 469
rect -241 367 -215 393
rect -165 367 -139 393
rect -89 367 -63 393
rect -13 367 13 393
rect 63 367 89 393
rect 139 367 165 393
rect 215 367 241 393
rect -241 291 -215 317
rect -165 291 -139 317
rect -89 291 -63 317
rect -13 291 13 317
rect 63 291 89 317
rect 139 291 165 317
rect 215 291 241 317
rect -241 215 -215 241
rect -165 215 -139 241
rect -89 215 -63 241
rect -13 215 13 241
rect 63 215 89 241
rect 139 215 165 241
rect 215 215 241 241
rect -241 139 -215 165
rect -165 139 -139 165
rect -89 139 -63 165
rect -13 139 13 165
rect 63 139 89 165
rect 139 139 165 165
rect 215 139 241 165
rect -241 63 -215 89
rect -165 63 -139 89
rect -89 63 -63 89
rect -13 63 13 89
rect 63 63 89 89
rect 139 63 165 89
rect 215 63 241 89
rect -241 -13 -215 13
rect -165 -13 -139 13
rect -89 -13 -63 13
rect -13 -13 13 13
rect 63 -13 89 13
rect 139 -13 165 13
rect 215 -13 241 13
rect -241 -89 -215 -63
rect -165 -89 -139 -63
rect -89 -89 -63 -63
rect -13 -89 13 -63
rect 63 -89 89 -63
rect 139 -89 165 -63
rect 215 -89 241 -63
rect -241 -165 -215 -139
rect -165 -165 -139 -139
rect -89 -165 -63 -139
rect -13 -165 13 -139
rect 63 -165 89 -139
rect 139 -165 165 -139
rect 215 -165 241 -139
rect -241 -241 -215 -215
rect -165 -241 -139 -215
rect -89 -241 -63 -215
rect -13 -241 13 -215
rect 63 -241 89 -215
rect 139 -241 165 -215
rect 215 -241 241 -215
rect -241 -317 -215 -291
rect -165 -317 -139 -291
rect -89 -317 -63 -291
rect -13 -317 13 -291
rect 63 -317 89 -291
rect 139 -317 165 -291
rect 215 -317 241 -291
rect -241 -393 -215 -367
rect -165 -393 -139 -367
rect -89 -393 -63 -367
rect -13 -393 13 -367
rect 63 -393 89 -367
rect 139 -393 165 -367
rect 215 -393 241 -367
rect -241 -469 -215 -443
rect -165 -469 -139 -443
rect -89 -469 -63 -443
rect -13 -469 13 -443
rect 63 -469 89 -443
rect 139 -469 165 -443
rect 215 -469 241 -443
rect -241 -545 -215 -519
rect -165 -545 -139 -519
rect -89 -545 -63 -519
rect -13 -545 13 -519
rect 63 -545 89 -519
rect 139 -545 165 -519
rect 215 -545 241 -519
<< metal2 >>
rect -247 545 247 551
rect -247 519 -241 545
rect -215 519 -165 545
rect -139 519 -89 545
rect -63 519 -13 545
rect 13 519 63 545
rect 89 519 139 545
rect 165 519 215 545
rect 241 519 247 545
rect -247 469 247 519
rect -247 443 -241 469
rect -215 443 -165 469
rect -139 443 -89 469
rect -63 443 -13 469
rect 13 443 63 469
rect 89 443 139 469
rect 165 443 215 469
rect 241 443 247 469
rect -247 393 247 443
rect -247 367 -241 393
rect -215 367 -165 393
rect -139 367 -89 393
rect -63 367 -13 393
rect 13 367 63 393
rect 89 367 139 393
rect 165 367 215 393
rect 241 367 247 393
rect -247 317 247 367
rect -247 291 -241 317
rect -215 291 -165 317
rect -139 291 -89 317
rect -63 291 -13 317
rect 13 291 63 317
rect 89 291 139 317
rect 165 291 215 317
rect 241 291 247 317
rect -247 241 247 291
rect -247 215 -241 241
rect -215 215 -165 241
rect -139 215 -89 241
rect -63 215 -13 241
rect 13 215 63 241
rect 89 215 139 241
rect 165 215 215 241
rect 241 215 247 241
rect -247 165 247 215
rect -247 139 -241 165
rect -215 139 -165 165
rect -139 139 -89 165
rect -63 139 -13 165
rect 13 139 63 165
rect 89 139 139 165
rect 165 139 215 165
rect 241 139 247 165
rect -247 89 247 139
rect -247 63 -241 89
rect -215 63 -165 89
rect -139 63 -89 89
rect -63 63 -13 89
rect 13 63 63 89
rect 89 63 139 89
rect 165 63 215 89
rect 241 63 247 89
rect -247 13 247 63
rect -247 -13 -241 13
rect -215 -13 -165 13
rect -139 -13 -89 13
rect -63 -13 -13 13
rect 13 -13 63 13
rect 89 -13 139 13
rect 165 -13 215 13
rect 241 -13 247 13
rect -247 -63 247 -13
rect -247 -89 -241 -63
rect -215 -89 -165 -63
rect -139 -89 -89 -63
rect -63 -89 -13 -63
rect 13 -89 63 -63
rect 89 -89 139 -63
rect 165 -89 215 -63
rect 241 -89 247 -63
rect -247 -139 247 -89
rect -247 -165 -241 -139
rect -215 -165 -165 -139
rect -139 -165 -89 -139
rect -63 -165 -13 -139
rect 13 -165 63 -139
rect 89 -165 139 -139
rect 165 -165 215 -139
rect 241 -165 247 -139
rect -247 -215 247 -165
rect -247 -241 -241 -215
rect -215 -241 -165 -215
rect -139 -241 -89 -215
rect -63 -241 -13 -215
rect 13 -241 63 -215
rect 89 -241 139 -215
rect 165 -241 215 -215
rect 241 -241 247 -215
rect -247 -291 247 -241
rect -247 -317 -241 -291
rect -215 -317 -165 -291
rect -139 -317 -89 -291
rect -63 -317 -13 -291
rect 13 -317 63 -291
rect 89 -317 139 -291
rect 165 -317 215 -291
rect 241 -317 247 -291
rect -247 -367 247 -317
rect -247 -393 -241 -367
rect -215 -393 -165 -367
rect -139 -393 -89 -367
rect -63 -393 -13 -367
rect 13 -393 63 -367
rect 89 -393 139 -367
rect 165 -393 215 -367
rect 241 -393 247 -367
rect -247 -443 247 -393
rect -247 -469 -241 -443
rect -215 -469 -165 -443
rect -139 -469 -89 -443
rect -63 -469 -13 -443
rect 13 -469 63 -443
rect 89 -469 139 -443
rect 165 -469 215 -443
rect 241 -469 247 -443
rect -247 -519 247 -469
rect -247 -545 -241 -519
rect -215 -545 -165 -519
rect -139 -545 -89 -519
rect -63 -545 -13 -519
rect 13 -545 63 -519
rect 89 -545 139 -519
rect 165 -545 215 -519
rect 241 -545 247 -519
rect -247 -551 247 -545
<< end >>
