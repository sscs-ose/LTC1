magic
tech gf180mcuC
magscale 1 10
timestamp 1699883071
<< nwell >>
rect 0 737 884 868
<< psubdiff >>
rect 265 -33 619 -20
rect 265 -79 278 -33
rect 324 -79 372 -33
rect 418 -79 466 -33
rect 512 -79 560 -33
rect 606 -79 619 -33
rect 265 -92 619 -79
<< nsubdiff >>
rect 30 822 854 835
rect 30 776 43 822
rect 89 776 137 822
rect 183 776 231 822
rect 277 776 325 822
rect 371 776 419 822
rect 465 776 513 822
rect 559 776 607 822
rect 653 776 701 822
rect 747 776 795 822
rect 841 776 854 822
rect 30 763 854 776
<< psubdiffcont >>
rect 278 -79 324 -33
rect 372 -79 418 -33
rect 466 -79 512 -33
rect 560 -79 606 -33
<< nsubdiffcont >>
rect 43 776 89 822
rect 137 776 183 822
rect 231 776 277 822
rect 325 776 371 822
rect 419 776 465 822
rect 513 776 559 822
rect 607 776 653 822
rect 701 776 747 822
rect 795 776 841 822
<< polysilicon >>
rect 174 268 230 446
rect 155 260 230 268
rect 334 260 390 440
rect 155 255 390 260
rect 155 209 168 255
rect 214 209 390 255
rect 155 204 390 209
rect 155 196 227 204
rect 334 162 390 204
rect 494 343 550 440
rect 654 343 710 446
rect 494 287 714 343
rect 494 162 550 287
rect 658 230 714 287
rect 762 230 834 238
rect 658 225 834 230
rect 658 178 775 225
rect 821 178 834 225
rect 658 174 834 178
rect 762 165 834 174
<< polycontact >>
rect 168 209 214 255
rect 775 178 821 225
<< metal1 >>
rect 0 822 884 855
rect 0 776 43 822
rect 89 776 137 822
rect 183 776 231 822
rect 277 776 325 822
rect 371 776 419 822
rect 465 776 513 822
rect 559 776 607 822
rect 653 776 701 822
rect 747 776 795 822
rect 841 776 884 822
rect 0 743 884 776
rect 259 576 305 743
rect 419 651 785 697
rect 419 576 465 651
rect 739 578 785 651
rect 99 363 145 470
rect 419 363 465 464
rect 99 317 465 363
rect 579 363 625 478
rect 579 317 713 363
rect 157 255 225 266
rect 579 258 625 317
rect 113 209 168 255
rect 214 209 225 255
rect 157 198 225 209
rect 419 212 625 258
rect 764 225 832 236
rect 419 137 465 212
rect 764 178 775 225
rect 821 178 902 225
rect 764 167 832 178
rect 259 0 305 98
rect 579 0 625 98
rect 222 -33 662 0
rect 222 -79 278 -33
rect 324 -79 372 -33
rect 418 -79 466 -33
rect 512 -79 560 -33
rect 606 -79 662 -33
rect 222 -112 662 -79
use nmos_3p3_GGGST2#0  nmos_3p3_GGGST2_0
timestamp 1691670445
transform 1 0 522 0 1 118
box -140 -118 140 118
use nmos_3p3_GGGST2#0  nmos_3p3_GGGST2_1
timestamp 1691670445
transform 1 0 362 0 1 118
box -140 -118 140 118
use pmos_3p3_MEVUAR  pmos_3p3_MEVUAR_0 ~/GF180Projects/Tapeout/Magic/Logic_Gates/OR_2_Input
timestamp 1692335619
transform 1 0 602 0 1 507
box -282 -230 282 230
use pmos_3p3_MEVUAR  pmos_3p3_MEVUAR_1
timestamp 1692335619
transform 1 0 282 0 1 507
box -282 -230 282 230
<< labels >>
flabel metal1 437 -56 437 -56 0 FreeSans 320 0 0 0 VSS
port 7 nsew
flabel nsubdiffcont 442 799 442 799 0 FreeSans 320 0 0 0 VDD
port 6 nsew
flabel metal1 123 232 123 232 0 FreeSans 320 0 0 0 A
port 0 nsew
flabel metal1 888 202 888 202 0 FreeSans 320 0 0 0 B
port 1 nsew
flabel metal1 681 340 681 340 0 FreeSans 320 0 0 0 OUT
port 4 nsew
flabel metal1 282 341 282 341 0 FreeSans 320 0 0 0 SD1
port 10 nsew
<< end >>
