* NGSPICE file created from VCO_mag_flat.ext - technology: gf180mcuC

.subckt VCO_mag_flat OUTB OUT VCONT EN VSS VDD
X0 VDD a_2201_n2780.t12 a_510_n1078# VDD.t101 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X1 VDD GF_INV16_1.IN OUTB.t5 VDD.t173 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X2 a_510_2660# a_2201_958.t12 VDD.t184 VDD.t161 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X3 Delay_Cell_mag_2.IN Delay_Cell_mag_2.INB VDD.t40 VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X4 GF_INV1_1.OUT Delay_Cell_mag_1.IN VDD.t183 VDD.t182 pfet_03v3 ad=0.165p pd=1.64u as=0.165p ps=1.64u w=0.35u l=0.35u
X5 a_6953_2661# Delay_Cell_mag_1.IN Delay_Cell_mag_1.IN VDD.t113 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X6 VDD Delay_Cell_mag_2.OUT.t16 Delay_Cell_mag_2.OUTB.t7 VDD.t47 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X7 OUTB GF_INV16_1.IN VSS.t103 VSS.t102 nfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X8 VDD GF_INV16_1.IN OUTB.t4 VDD.t170 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.35u
X9 a_6953_2661# Delay_Cell_mag_1.INB.t6 Delay_Cell_mag_1.INB.t7 VDD.t120 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X10 Delay_Cell_mag_0.OUT Delay_Cell_mag_0.IN a_7148_n3320# VSS.t17 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X11 VDD Delay_Cell_mag_0.OUTB.t16 Delay_Cell_mag_0.OUT VDD.t124 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X12 VDD Delay_Cell_mag_2.OUT.t17 Delay_Cell_mag_0.INB VDD.t74 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X13 a_705_418# Delay_Cell_mag_1.INB.t16 Delay_Cell_mag_2.IN.t6 VSS.t20 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X14 VDD a_2201_958.t13 a_510_2660# VDD.t105 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X15 VDD Delay_Cell_mag_2.IN.t16 Delay_Cell_mag_2.INB VDD.t38 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X16 Delay_Cell_mag_1.IN Delay_Cell_mag_0.OUT a_7148_419# VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X17 OUTB GF_INV16_1.IN VSS.t101 VSS.t100 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X18 Delay_Cell_mag_2.INB Delay_Cell_mag_1.IN a_705_418# VSS.t108 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X19 VSS VCONT.t2 a_2201_958.t10 VSS.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X20 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.OUTB.t10 a_6953_n1078# VDD.t131 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X21 a_7148_419# Delay_Cell_mag_0.OUTB.t18 Delay_Cell_mag_1.INB.t14 VSS.t114 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X22 a_7148_n3320# Delay_Cell_mag_0.INB Delay_Cell_mag_0.OUTB.t3 VSS.t3 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X23 OUT GF_INV16_2.IN VSS.t30 VSS.t29 nfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X24 Delay_Cell_mag_2.IN Delay_Cell_mag_2.IN.t14 a_510_2660# VDD.t39 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X25 GF_INV1_0.OUT Delay_Cell_mag_1.INB.t17 VDD.t63 VDD.t62 pfet_03v3 ad=0.165p pd=1.64u as=0.165p ps=1.64u w=0.35u l=0.35u
X26 VSS GF_INV1_1.OUT GF_INV16_1.IN VSS.t54 nfet_03v3 ad=0.308p pd=2.28u as=0.182p ps=1.22u w=0.7u l=0.35u
X27 Delay_Cell_mag_0.IN Delay_Cell_mag_2.OUTB.t16 VDD.t86 VDD.t85 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X28 VDD a_8644_959.t6 a_8644_959.t7 VDD.t134 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X29 Delay_Cell_mag_2.OUTB Delay_Cell_mag_2.OUTB.t14 a_510_n1078# VDD.t87 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X30 Delay_Cell_mag_0.IN Delay_Cell_mag_2.OUTB.t18 VDD.t14 VDD.t13 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X31 a_6953_n1078# a_8644_n2780.t13 VDD.t12 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X32 a_705_n3320# EN.t0 VSS.t51 VSS.t50 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X33 Delay_Cell_mag_0.OUT Delay_Cell_mag_0.OUT a_6953_n1078# VDD.t133 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X34 a_705_418# a_705_418# a_705_418# VSS.t9 nfet_03v3 ad=0.44p pd=2.88u as=4p ps=24u w=1u l=0.56u
X35 a_7148_419# a_7148_419# a_7148_419# VSS.t34 nfet_03v3 ad=0.26p pd=1.52u as=4p ps=24u w=1u l=0.56u
X36 a_510_2660# Delay_Cell_mag_2.INB Delay_Cell_mag_2.INB VDD.t38 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X37 a_705_n3320# Delay_Cell_mag_2.IN.t18 Delay_Cell_mag_2.OUT.t15 VSS.t50 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X38 a_510_n1078# Delay_Cell_mag_2.OUTB.t12 Delay_Cell_mag_2.OUTB.t13 VDD.t55 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X39 a_7148_n3320# a_7148_n3320# a_7148_n3320# VSS.t19 nfet_03v3 ad=0.44p pd=2.88u as=4p ps=24u w=1u l=0.56u
X40 GF_INV16_1.IN GF_INV1_1.OUT VDD.t143 VDD.t142 pfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X41 VSS VCONT.t3 a_2201_n2780.t10 VSS.t7 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X42 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.OUT VDD.t132 VDD.t131 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X43 VDD Delay_Cell_mag_2.OUTB.t19 Delay_Cell_mag_0.IN VDD.t5 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X44 a_6953_n1078# Delay_Cell_mag_0.OUT Delay_Cell_mag_0.OUT VDD.t77 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X45 GF_INV16_1.IN GF_INV1_1.OUT VSS.t53 VSS.t52 nfet_03v3 ad=0.182p pd=1.22u as=0.308p ps=2.28u w=0.7u l=0.35u
X46 VDD GF_INV1_0.OUT GF_INV16_2.IN VDD.t152 pfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X47 a_6953_2661# a_8644_959.t14 VDD.t135 VDD.t134 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X48 Delay_Cell_mag_1.INB Delay_Cell_mag_1.IN VDD.t181 VDD.t43 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X49 Delay_Cell_mag_2.OUTB Delay_Cell_mag_2.OUT.t18 VDD.t88 VDD.t87 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X50 a_7148_419# Delay_Cell_mag_0.OUT Delay_Cell_mag_1.IN VSS.t40 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X51 VDD a_8644_n2780.t7 a_8644_n2780.t8 VDD.t11 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X52 Delay_Cell_mag_2.OUTB Delay_Cell_mag_2.INB a_705_n3320# VSS.t7 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X53 Delay_Cell_mag_0.OUT Delay_Cell_mag_0.OUTB.t19 VDD.t187 VDD.t133 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X54 a_705_418# a_705_418# a_705_418# VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.56u
X55 VDD a_2201_958.t6 a_2201_958.t7 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X56 VDD a_8644_959.t15 a_6953_2661# VDD.t116 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X57 Delay_Cell_mag_1.INB Delay_Cell_mag_0.OUTB.t20 a_7148_419# VSS.t31 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X58 VDD a_2201_n2780.t14 a_510_n1078# VDD.t97 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X59 VDD Delay_Cell_mag_2.OUT.t19 Delay_Cell_mag_0.INB VDD.t50 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X60 VSS VCONT.t5 a_8644_959.t10 VSS.t41 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X61 a_705_418# Delay_Cell_mag_1.IN Delay_Cell_mag_2.INB VSS.t44 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X62 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.OUTB.t8 a_6953_n1078# VDD.t129 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X63 VDD a_8644_959.t16 a_6953_2661# VDD.t145 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X64 VDD Delay_Cell_mag_1.IN Delay_Cell_mag_1.INB.t12 VDD.t42 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X65 GF_INV1_1.OUT Delay_Cell_mag_1.IN VSS.t107 VSS.t106 nfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.35u
X66 VDD Delay_Cell_mag_2.OUT.t20 Delay_Cell_mag_2.OUTB.t5 VDD.t55 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X67 VDD GF_INV16_2.IN OUT.t3 VDD.t71 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X68 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.IN.t19 a_705_n3320# VSS.t113 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X69 VDD Delay_Cell_mag_0.OUTB.t22 Delay_Cell_mag_0.OUT VDD.t77 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X70 VDD GF_INV16_2.IN OUT.t2 VDD.t68 pfet_03v3 ad=1.23p pd=6.48u as=0.728p ps=3.32u w=2.8u l=0.35u
X71 Delay_Cell_mag_1.INB Delay_Cell_mag_1.INB.t4 a_6953_2661# VDD.t43 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X72 a_705_n3320# Delay_Cell_mag_2.INB Delay_Cell_mag_2.OUTB.t2 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X73 a_510_2660# a_2201_958.t15 VDD.t84 VDD.t83 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X74 Delay_Cell_mag_2.INB Delay_Cell_mag_2.IN.t20 VDD.t16 VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X75 VSS VCONT.t8 a_8644_959.t9 VSS.t34 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X76 Delay_Cell_mag_0.IN Delay_Cell_mag_2.OUTB.t20 VSS.t124 VSS.t123 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X77 Delay_Cell_mag_0.INB Delay_Cell_mag_2.OUT.t21 VSS.t66 VSS.t65 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X78 Delay_Cell_mag_0.INB Delay_Cell_mag_2.OUT.t22 VSS.t64 VSS.t63 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X79 OUT GF_INV16_2.IN VSS.t28 VSS.t27 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X80 Delay_Cell_mag_0.IN Delay_Cell_mag_2.OUTB.t21 VSS.t122 VSS.t121 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.35u
X81 a_7148_n3320# Delay_Cell_mag_0.INB Delay_Cell_mag_0.OUTB.t2 VSS.t2 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X82 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.IN.t21 a_705_n3320# VSS.t112 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X83 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.OUT VDD.t130 VDD.t129 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X84 GF_INV1_0.OUT Delay_Cell_mag_1.INB.t19 VSS.t11 VSS.t10 nfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.35u
X85 a_6953_2661# Delay_Cell_mag_1.INB.t2 Delay_Cell_mag_1.INB.t3 VDD.t42 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X86 a_705_n3320# a_705_n3320# a_705_n3320# VSS.t36 nfet_03v3 ad=0.44p pd=2.88u as=4p ps=24u w=1u l=0.56u
X87 VSS GF_INV16_1.IN OUTB.t7 VSS.t97 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X88 a_705_418# Delay_Cell_mag_1.INB.t20 Delay_Cell_mag_2.IN.t4 VSS.t12 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X89 Delay_Cell_mag_2.OUTB Delay_Cell_mag_2.OUTB.t10 a_510_n1078# VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X90 VDD a_2201_958.t16 a_510_2660# VDD.t8 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X91 Delay_Cell_mag_0.OUT Delay_Cell_mag_0.OUT a_6953_n1078# VDD.t128 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X92 a_7148_419# Delay_Cell_mag_0.OUTB.t23 Delay_Cell_mag_1.INB.t9 VSS.t32 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X93 VSS GF_INV16_1.IN OUTB.t6 VSS.t94 nfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X94 Delay_Cell_mag_2.IN Delay_Cell_mag_1.INB.t21 a_705_418# VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X95 VDD Delay_Cell_mag_2.IN.t22 Delay_Cell_mag_2.INB VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X96 VDD Delay_Cell_mag_2.OUTB.t23 Delay_Cell_mag_0.IN VDD.t26 pfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.35u
X97 a_510_n1078# Delay_Cell_mag_2.OUT.t9 Delay_Cell_mag_2.OUT.t10 VDD.t59 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X98 VSS VCONT.t10 a_2201_958.t8 VSS.t8 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X99 a_510_n1078# a_2201_n2780.t16 VDD.t96 VDD.t93 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X100 VSS Delay_Cell_mag_2.OUTB.t24 Delay_Cell_mag_0.IN VSS.t118 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X101 VSS Delay_Cell_mag_2.OUT.t23 Delay_Cell_mag_0.INB VSS.t60 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.35u
X102 Delay_Cell_mag_2.INB Delay_Cell_mag_2.INB a_510_2660# VDD.t15 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X103 VDD Delay_Cell_mag_1.INB.t22 Delay_Cell_mag_1.IN VDD.t44 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X104 a_7148_n3320# Delay_Cell_mag_0.IN Delay_Cell_mag_0.OUT VSS.t16 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X105 a_6953_n1078# Delay_Cell_mag_0.OUTB.t6 Delay_Cell_mag_0.OUTB.t7 VDD.t125 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X106 a_705_418# EN.t1 VSS.t45 VSS.t44 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X107 VSS VCONT.t11 a_2201_n2780.t8 VSS.t35 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X108 VSS EN.t2 a_7148_n3320# VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X109 Delay_Cell_mag_2.OUTB Delay_Cell_mag_2.OUT.t24 VDD.t108 VDD.t17 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X110 a_705_n3320# a_705_n3320# a_705_n3320# VSS.t35 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.56u
X111 Delay_Cell_mag_1.IN Delay_Cell_mag_1.INB.t23 VDD.t110 VDD.t109 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X112 Delay_Cell_mag_0.OUT Delay_Cell_mag_0.OUTB.t24 VDD.t193 VDD.t128 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X113 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.INB a_7148_n3320# VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X114 a_510_2660# Delay_Cell_mag_2.INB Delay_Cell_mag_2.INB VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X115 VDD GF_INV1_1.OUT GF_INV16_1.IN VDD.t139 pfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X116 GF_INV16_2.IN GF_INV1_0.OUT VDD.t151 VDD.t150 pfet_03v3 ad=0.364p pd=1.92u as=0.616p ps=3.68u w=1.4u l=0.35u
X117 VDD Delay_Cell_mag_2.OUTB.t25 Delay_Cell_mag_2.OUT.t2 VDD.t59 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X118 a_510_n1078# Delay_Cell_mag_2.OUT.t7 Delay_Cell_mag_2.OUT.t8 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X119 OUTB GF_INV16_1.IN VDD.t169 VDD.t168 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.35u
X120 VDD a_8644_n2780.t14 a_6953_n1078# VDD.t23 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X121 Delay_Cell_mag_1.IN Delay_Cell_mag_1.INB.t24 VDD.t112 VDD.t111 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X122 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.OUT.t5 a_510_n1078# VDD.t159 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X123 VDD a_2201_n2780.t2 a_2201_n2780.t3 VDD.t93 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X124 Delay_Cell_mag_2.IN Delay_Cell_mag_2.INB VDD.t37 VDD.t36 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X125 a_6953_2661# Delay_Cell_mag_1.IN Delay_Cell_mag_1.IN VDD.t44 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X126 Delay_Cell_mag_1.INB Delay_Cell_mag_1.IN VDD.t178 VDD.t41 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X127 VDD Delay_Cell_mag_0.OUT Delay_Cell_mag_0.OUTB.t13 VDD.t125 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X128 OUTB GF_INV16_1.IN VDD.t167 VDD.t166 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
X129 VDD Delay_Cell_mag_2.INB Delay_Cell_mag_2.IN.t1 VDD.t33 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X130 a_6953_n1078# a_8644_n2780.t15 VDD.t144 VDD.t80 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X131 Delay_Cell_mag_1.IN Delay_Cell_mag_0.OUT a_7148_419# VSS.t39 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X132 VSS GF_INV1_0.OUT GF_INV16_2.IN VSS.t82 nfet_03v3 ad=0.308p pd=2.28u as=0.182p ps=1.22u w=0.7u l=0.35u
X133 VSS EN.t3 a_705_n3320# VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X134 OUT GF_INV16_2.IN VDD.t67 VDD.t66 pfet_03v3 ad=0.728p pd=3.32u as=1.23p ps=6.48u w=2.8u l=0.35u
X135 VDD Delay_Cell_mag_2.INB Delay_Cell_mag_2.IN.t0 VDD.t30 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X136 Delay_Cell_mag_1.IN Delay_Cell_mag_1.IN a_6953_2661# VDD.t109 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X137 a_7148_419# EN.t4 VSS.t76 VSS.t32 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X138 VSS EN.t5 a_705_418# VSS.t13 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X139 a_7148_419# a_7148_419# a_7148_419# VSS.t33 nfet_03v3 ad=0.44p pd=2.88u as=0 ps=0 w=1u l=0.56u
X140 VDD Delay_Cell_mag_2.OUTB.t26 Delay_Cell_mag_2.OUT.t0 VDD.t18 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X141 Delay_Cell_mag_2.OUTB Delay_Cell_mag_2.INB a_705_n3320# VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X142 Delay_Cell_mag_1.IN Delay_Cell_mag_1.IN a_6953_2661# VDD.t111 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X143 Delay_Cell_mag_2.INB Delay_Cell_mag_1.IN a_705_418# VSS.t105 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X144 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.OUTB.t27 VDD.t160 VDD.t159 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X145 Delay_Cell_mag_0.OUT Delay_Cell_mag_0.IN a_7148_n3320# VSS.t15 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X146 Delay_Cell_mag_2.IN Delay_Cell_mag_2.IN.t12 a_510_2660# VDD.t36 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X147 Delay_Cell_mag_1.INB Delay_Cell_mag_1.INB.t0 a_6953_2661# VDD.t41 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X148 VSS Delay_Cell_mag_2.OUTB.t28 Delay_Cell_mag_0.IN VSS.t115 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X149 VSS Delay_Cell_mag_2.OUT.t26 Delay_Cell_mag_0.INB VSS.t57 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.35u
X150 VSS GF_INV16_2.IN OUT.t5 VSS.t24 nfet_03v3 ad=0.364p pd=1.92u as=0.364p ps=1.92u w=1.4u l=0.35u
X151 a_7148_n3320# EN.t6 VSS.t79 VSS.t14 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X152 a_510_2660# Delay_Cell_mag_2.IN.t10 Delay_Cell_mag_2.IN.t11 VDD.t33 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X153 a_705_n3320# Delay_Cell_mag_2.INB Delay_Cell_mag_2.OUTB.t0 VSS.t4 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X154 VSS GF_INV16_2.IN OUT.t4 VSS.t21 nfet_03v3 ad=0.616p pd=3.68u as=0.364p ps=1.92u w=1.4u l=0.35u
X155 Delay_Cell_mag_2.INB Delay_Cell_mag_2.IN.t24 VDD.t58 VDD.t29 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X156 VSS VCONT.t14 a_8644_n2780.t11 VSS.t18 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X157 VDD a_8644_n2780.t3 a_8644_n2780.t4 VDD.t80 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X158 a_7148_n3320# Delay_Cell_mag_0.IN Delay_Cell_mag_0.OUT VSS.t14 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X159 a_510_2660# Delay_Cell_mag_2.IN.t8 Delay_Cell_mag_2.IN.t9 VDD.t30 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X160 a_510_n1078# a_2201_n2780.t17 VDD.t92 VDD.t89 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X161 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.OUT.t3 a_510_n1078# VDD.t21 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X162 a_7148_n3320# a_7148_n3320# a_7148_n3320# VSS.t18 nfet_03v3 ad=0.26p pd=1.52u as=0 ps=0 w=1u l=0.56u
X163 a_6953_n1078# Delay_Cell_mag_0.OUTB.t4 Delay_Cell_mag_0.OUTB.t5 VDD.t121 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X164 GF_INV16_2.IN GF_INV1_0.OUT VSS.t81 VSS.t80 nfet_03v3 ad=0.182p pd=1.22u as=0.308p ps=2.28u w=0.7u l=0.35u
X165 VDD a_8644_959.t0 a_8644_959.t1 VDD.t155 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X166 VSS VCONT.t15 a_8644_n2780.t2 VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X167 a_7148_419# Delay_Cell_mag_0.OUT Delay_Cell_mag_1.IN VSS.t38 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X168 Delay_Cell_mag_2.IN Delay_Cell_mag_1.INB.t26 a_705_418# VSS.t37 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X169 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.INB a_7148_n3320# VSS.t0 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X170 a_705_n3320# Delay_Cell_mag_2.IN.t25 Delay_Cell_mag_2.OUT.t12 VSS.t111 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X171 Delay_Cell_mag_1.INB Delay_Cell_mag_0.OUTB.t25 a_7148_419# VSS.t125 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X172 VDD a_2201_958.t2 a_2201_958.t3 VDD.t161 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X173 VDD Delay_Cell_mag_1.INB.t27 Delay_Cell_mag_1.IN VDD.t113 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X174 VDD a_8644_n2780.t17 a_6953_n1078# VDD.t148 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X175 a_705_418# Delay_Cell_mag_1.IN Delay_Cell_mag_2.INB VSS.t104 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X176 Delay_Cell_mag_2.INB Delay_Cell_mag_2.INB a_510_2660# VDD.t29 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.56u
X177 VSS EN.t7 a_7148_419# VSS.t39 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X178 a_510_n1078# Delay_Cell_mag_2.OUTB.t8 Delay_Cell_mag_2.OUTB.t9 VDD.t47 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X179 VDD Delay_Cell_mag_1.IN Delay_Cell_mag_1.INB.t10 VDD.t120 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X180 a_6953_n1078# Delay_Cell_mag_0.OUT Delay_Cell_mag_0.OUT VDD.t124 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X181 VDD a_2201_n2780.t0 a_2201_n2780.t1 VDD.t89 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X182 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.OUTB.t29 VDD.t22 VDD.t21 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X183 Delay_Cell_mag_0.INB Delay_Cell_mag_2.OUT.t28 VDD.t4 VDD.t3 pfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.35u
X184 Delay_Cell_mag_0.INB Delay_Cell_mag_2.OUT.t29 VDD.t165 VDD.t164 pfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.35u
X185 VDD Delay_Cell_mag_0.OUT Delay_Cell_mag_0.OUTB.t12 VDD.t121 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.56u
X186 a_6953_2661# a_8644_959.t17 VDD.t156 VDD.t155 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.56u
X187 OUT GF_INV16_2.IN VDD.t65 VDD.t64 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.35u
R0 a_2201_n2780.t0 a_2201_n2780.n4 22.8782
R1 a_2201_n2780.n5 a_2201_n2780.t0 22.4219
R2 a_2201_n2780.n2 a_2201_n2780.t12 22.2916
R3 a_2201_n2780.n4 a_2201_n2780.n3 14.0791
R4 a_2201_n2780.n3 a_2201_n2780.n2 14.0791
R5 a_2201_n2780.n6 a_2201_n2780.n5 14.0791
R6 a_2201_n2780.n1 a_2201_n2780.t6 11.3416
R7 a_2201_n2780.n5 a_2201_n2780.t4 8.34336
R8 a_2201_n2780.n6 a_2201_n2780.t2 8.34336
R9 a_2201_n2780.n4 a_2201_n2780.t17 8.213
R10 a_2201_n2780.n3 a_2201_n2780.t14 8.213
R11 a_2201_n2780.n2 a_2201_n2780.t16 8.213
R12 a_2201_n2780.n0 a_2201_n2780.n6 8.17193
R13 a_2201_n2780.n0 a_2201_n2780.n1 4.0005
R14 a_2201_n2780.n0 a_2201_n2780.n8 3.63045
R15 a_2201_n2780.n17 a_2201_n2780.n0 2.89398
R16 a_2201_n2780.n13 a_2201_n2780.n10 2.26392
R17 a_2201_n2780.n8 a_2201_n2780.t1 1.8205
R18 a_2201_n2780.n8 a_2201_n2780.n7 1.8205
R19 a_2201_n2780.t3 a_2201_n2780.n17 1.8205
R20 a_2201_n2780.n17 a_2201_n2780.n16 1.8205
R21 a_2201_n2780.n10 a_2201_n2780.t10 1.6385
R22 a_2201_n2780.n10 a_2201_n2780.n9 1.6385
R23 a_2201_n2780.n12 a_2201_n2780.t8 1.6385
R24 a_2201_n2780.n12 a_2201_n2780.n11 1.6385
R25 a_2201_n2780.n1 a_2201_n2780.n15 1.62996
R26 a_2201_n2780.n13 a_2201_n2780.n12 1.4936
R27 a_2201_n2780.n0 a_2201_n2780.n14 1.37554
R28 a_2201_n2780.n14 a_2201_n2780.n13 1.18673
R29 VDD.n260 VDD.t62 335.682
R30 VDD.n208 VDD.t182 335.682
R31 VDD.n52 VDD.t26 179.427
R32 VDD.n481 VDD.t50 179.427
R33 VDD.n63 VDD.t5 112.441
R34 VDD.n487 VDD.t74 112.441
R35 VDD.n65 VDD.t85 52.6321
R36 VDD.n485 VDD.t3 52.6321
R37 VDD.n190 VDD.t64 46.3367
R38 VDD.n243 VDD.t166 46.3367
R39 VDD.n324 VDD.t155 42.1692
R40 VDD.n434 VDD.t80 42.1692
R41 VDD.n502 VDD.t89 42.1692
R42 VDD.n686 VDD.t161 42.1692
R43 VDD.n265 VDD.t150 39.8225
R44 VDD.n213 VDD.t142 39.8225
R45 VDD.n321 VDD.t116 35.5427
R46 VDD.n437 VDD.t148 35.5427
R47 VDD.n505 VDD.t97 35.5427
R48 VDD.n683 VDD.t105 35.5427
R49 VDD.n193 VDD.t68 32.3281
R50 VDD.n246 VDD.t170 32.3281
R51 VDD.n291 VDD.t41 30.7234
R52 VDD.n467 VDD.t133 30.7234
R53 VDD.n535 VDD.t159 30.7234
R54 VDD.n653 VDD.t29 30.7234
R55 VDD.n318 VDD.t134 28.9162
R56 VDD.n440 VDD.t11 28.9162
R57 VDD.n508 VDD.t93 28.9162
R58 VDD.n680 VDD.t83 28.9162
R59 VDD.n294 VDD.t42 24.0969
R60 VDD.n464 VDD.t124 24.0969
R61 VDD.n532 VDD.t59 24.0969
R62 VDD.n656 VDD.t0 24.0969
R63 VDD.n56 VDD.t13 23.9239
R64 VDD.n493 VDD.t164 23.9239
R65 VDD.n315 VDD.t145 22.2897
R66 VDD.n443 VDD.t23 22.2897
R67 VDD.n511 VDD.t101 22.2897
R68 VDD.n677 VDD.t8 22.2897
R69 VDD.n297 VDD.t43 17.4704
R70 VDD.n461 VDD.t128 17.4704
R71 VDD.n529 VDD.t21 17.4704
R72 VDD.n659 VDD.t15 17.4704
R73 VDD.n177 VDD.t66 16.8707
R74 VDD.n230 VDD.t168 16.8707
R75 VDD.n183 VDD.t71 16.1643
R76 VDD.n236 VDD.t173 16.1643
R77 VDD.n312 VDD.t44 15.6632
R78 VDD.n446 VDD.t121 15.6632
R79 VDD.n514 VDD.t55 15.6632
R80 VDD.n674 VDD.t33 15.6632
R81 VDD.n300 VDD.t120 10.8439
R82 VDD.n458 VDD.t77 10.8439
R83 VDD.n526 VDD.t18 10.8439
R84 VDD.n662 VDD.t38 10.8439
R85 VDD.n265 VDD.n264 9.93878
R86 VDD.n213 VDD.n212 9.93878
R87 VDD.n271 VDD.t152 9.6712
R88 VDD.n219 VDD.t139 9.6712
R89 VDD.n309 VDD.t109 9.03664
R90 VDD.n449 VDD.t129 9.03664
R91 VDD.n517 VDD.t17 9.03664
R92 VDD.n671 VDD.t36 9.03664
R93 VDD.n66 VDD.n64 8.70445
R94 VDD.n488 VDD.n486 8.70445
R95 VDD.n258 VDD.t63 8.26313
R96 VDD.n206 VDD.t183 8.26313
R97 VDD.n184 VDD.n182 8.15819
R98 VDD.n237 VDD.n235 8.15819
R99 VDD.n649 VDD.n590 7.10822
R100 VDD.n483 VDD.n480 6.66125
R101 VDD.n58 VDD.t14 6.58259
R102 VDD.n69 VDD.n51 6.49073
R103 VDD.n496 VDD.t165 6.48786
R104 VDD.n198 VDD.n197 6.3005
R105 VDD.n197 VDD.n196 6.3005
R106 VDD.n477 VDD.n69 6.07717
R107 VDD.n202 VDD.n201 5.38954
R108 VDD.n332 VDD.n331 4.85019
R109 VDD.n285 VDD.n284 4.5005
R110 VDD.n330 VDD.n151 4.5005
R111 VDD.n74 VDD.n73 4.5005
R112 VDD.n498 VDD.n497 4.46272
R113 VDD.n264 VDD.t151 4.3192
R114 VDD.n275 VDD.n263 4.3192
R115 VDD.n212 VDD.t143 4.3192
R116 VDD.n223 VDD.n211 4.3192
R117 VDD.n262 VDD.n261 4.29708
R118 VDD.n210 VDD.n209 4.29333
R119 VDD.n303 VDD.t111 4.21737
R120 VDD.n455 VDD.t131 4.21737
R121 VDD.n523 VDD.t87 4.21737
R122 VDD.n665 VDD.t39 4.21737
R123 VDD.n252 VDD.n251 3.94094
R124 VDD.n176 VDD.t67 3.92746
R125 VDD.n203 VDD.n173 3.92746
R126 VDD.n229 VDD.t169 3.92746
R127 VDD.n96 VDD.n95 3.9192
R128 VDD.n406 VDD.n405 3.9192
R129 VDD.n25 VDD.n24 3.9192
R130 VDD.n724 VDD.n723 3.9192
R131 VDD.n77 VDD.t178 3.80738
R132 VDD.n387 VDD.t187 3.80738
R133 VDD.n6 VDD.t160 3.80738
R134 VDD.n705 VDD.t58 3.80738
R135 VDD.n55 VDD.t86 3.6405
R136 VDD.n55 VDD.n54 3.6405
R137 VDD.n479 VDD.t4 3.6405
R138 VDD.n479 VDD.n478 3.6405
R139 VDD.n186 VDD.n175 3.27746
R140 VDD.n239 VDD.n228 3.27746
R141 VDD.n259 VDD.n258 3.19668
R142 VDD.n207 VDD.n206 3.19668
R143 VDD.n68 VDD.n53 3.1505
R144 VDD.n53 VDD.n52 3.1505
R145 VDD.n58 VDD.n57 3.1505
R146 VDD.n57 VDD.n56 3.1505
R147 VDD.n67 VDD.n66 3.1505
R148 VDD.n66 VDD.n65 3.1505
R149 VDD.n64 VDD.n62 3.1505
R150 VDD.n64 VDD.n63 3.1505
R151 VDD.n61 VDD.n60 3.1505
R152 VDD.n60 VDD.n59 3.1505
R153 VDD.n486 VDD.n484 3.1505
R154 VDD.n486 VDD.n485 3.1505
R155 VDD.n495 VDD.n494 3.1505
R156 VDD.n494 VDD.n493 3.1505
R157 VDD.n492 VDD.n491 3.1505
R158 VDD.n491 VDD.n490 3.1505
R159 VDD.n489 VDD.n488 3.1505
R160 VDD.n488 VDD.n487 3.1505
R161 VDD.n483 VDD.n482 3.1505
R162 VDD.n482 VDD.n481 3.1505
R163 VDD.n257 VDD.n256 3.1505
R164 VDD.n260 VDD.n259 3.1505
R165 VDD.n270 VDD.n269 3.1505
R166 VDD.n269 VDD.n268 3.1505
R167 VDD.n267 VDD.n266 3.1505
R168 VDD.n273 VDD.n272 3.1505
R169 VDD.n195 VDD.n194 3.1505
R170 VDD.n194 VDD.n193 3.1505
R171 VDD.n192 VDD.n191 3.1505
R172 VDD.n191 VDD.n190 3.1505
R173 VDD.n189 VDD.n188 3.1505
R174 VDD.n188 VDD.n187 3.1505
R175 VDD.n185 VDD.n184 3.1505
R176 VDD.n184 VDD.n183 3.1505
R177 VDD.n182 VDD.n180 3.1505
R178 VDD.n182 VDD.n181 3.1505
R179 VDD.n179 VDD.n178 3.1505
R180 VDD.n248 VDD.n247 3.1505
R181 VDD.n247 VDD.n246 3.1505
R182 VDD.n245 VDD.n244 3.1505
R183 VDD.n244 VDD.n243 3.1505
R184 VDD.n242 VDD.n241 3.1505
R185 VDD.n241 VDD.n240 3.1505
R186 VDD.n238 VDD.n237 3.1505
R187 VDD.n237 VDD.n236 3.1505
R188 VDD.n235 VDD.n233 3.1505
R189 VDD.n235 VDD.n234 3.1505
R190 VDD.n232 VDD.n231 3.1505
R191 VDD.n218 VDD.n217 3.1505
R192 VDD.n217 VDD.n216 3.1505
R193 VDD.n215 VDD.n214 3.1505
R194 VDD.n221 VDD.n220 3.1505
R195 VDD.n208 VDD.n207 3.1505
R196 VDD.n205 VDD.n204 3.1505
R197 VDD.n327 VDD.n153 3.1505
R198 VDD.n153 VDD.n152 3.1505
R199 VDD.n326 VDD.n325 3.1505
R200 VDD.n325 VDD.n324 3.1505
R201 VDD.n323 VDD.n322 3.1505
R202 VDD.n322 VDD.n321 3.1505
R203 VDD.n320 VDD.n319 3.1505
R204 VDD.n319 VDD.n318 3.1505
R205 VDD.n317 VDD.n316 3.1505
R206 VDD.n316 VDD.n315 3.1505
R207 VDD.n314 VDD.n313 3.1505
R208 VDD.n313 VDD.n312 3.1505
R209 VDD.n311 VDD.n310 3.1505
R210 VDD.n310 VDD.n309 3.1505
R211 VDD.n308 VDD.n307 3.1505
R212 VDD.n307 VDD.n306 3.1505
R213 VDD.n305 VDD.n304 3.1505
R214 VDD.n304 VDD.n303 3.1505
R215 VDD.n302 VDD.n301 3.1505
R216 VDD.n301 VDD.n300 3.1505
R217 VDD.n299 VDD.n298 3.1505
R218 VDD.n298 VDD.n297 3.1505
R219 VDD.n296 VDD.n295 3.1505
R220 VDD.n295 VDD.n294 3.1505
R221 VDD.n293 VDD.n292 3.1505
R222 VDD.n292 VDD.n291 3.1505
R223 VDD.n290 VDD.n289 3.1505
R224 VDD.n289 VDD.n288 3.1505
R225 VDD.n155 VDD.n154 3.1505
R226 VDD.n158 VDD.n157 3.1505
R227 VDD.n160 VDD.n159 3.1505
R228 VDD.n163 VDD.n162 3.1505
R229 VDD.n165 VDD.n164 3.1505
R230 VDD.n168 VDD.n167 3.1505
R231 VDD.n172 VDD.n171 3.1505
R232 VDD.n125 VDD.n124 3.1505
R233 VDD.n123 VDD.n122 3.1505
R234 VDD.n121 VDD.n120 3.1505
R235 VDD.n119 VDD.n118 3.1505
R236 VDD.n117 VDD.n116 3.1505
R237 VDD.n115 VDD.n114 3.1505
R238 VDD.n113 VDD.n112 3.1505
R239 VDD.n111 VDD.n110 3.1505
R240 VDD.n109 VDD.n108 3.1505
R241 VDD.n107 VDD.n106 3.1505
R242 VDD.n105 VDD.n104 3.1505
R243 VDD.n103 VDD.n102 3.1505
R244 VDD.n101 VDD.n100 3.1505
R245 VDD.n99 VDD.n98 3.1505
R246 VDD.n143 VDD.n142 3.1505
R247 VDD.n140 VDD.n139 3.1505
R248 VDD.n136 VDD.n135 3.1505
R249 VDD.n133 VDD.n132 3.1505
R250 VDD.n130 VDD.n129 3.1505
R251 VDD.n147 VDD.n146 3.1505
R252 VDD.n128 VDD.n127 3.1505
R253 VDD.n334 VDD.n333 3.1505
R254 VDD.n336 VDD.n335 3.1505
R255 VDD.n338 VDD.n337 3.1505
R256 VDD.n340 VDD.n339 3.1505
R257 VDD.n342 VDD.n341 3.1505
R258 VDD.n344 VDD.n343 3.1505
R259 VDD.n346 VDD.n345 3.1505
R260 VDD.n348 VDD.n347 3.1505
R261 VDD.n350 VDD.n349 3.1505
R262 VDD.n352 VDD.n351 3.1505
R263 VDD.n354 VDD.n353 3.1505
R264 VDD.n356 VDD.n355 3.1505
R265 VDD.n358 VDD.n357 3.1505
R266 VDD.n360 VDD.n359 3.1505
R267 VDD.n424 VDD.n423 3.1505
R268 VDD.n421 VDD.n420 3.1505
R269 VDD.n417 VDD.n416 3.1505
R270 VDD.n414 VDD.n413 3.1505
R271 VDD.n412 VDD.n411 3.1505
R272 VDD.n426 VDD.n425 3.1505
R273 VDD.n430 VDD.n429 3.1505
R274 VDD.n432 VDD.n431 3.1505
R275 VDD.n433 VDD.n432 3.1505
R276 VDD.n436 VDD.n435 3.1505
R277 VDD.n435 VDD.n434 3.1505
R278 VDD.n439 VDD.n438 3.1505
R279 VDD.n438 VDD.n437 3.1505
R280 VDD.n442 VDD.n441 3.1505
R281 VDD.n441 VDD.n440 3.1505
R282 VDD.n445 VDD.n444 3.1505
R283 VDD.n444 VDD.n443 3.1505
R284 VDD.n448 VDD.n447 3.1505
R285 VDD.n447 VDD.n446 3.1505
R286 VDD.n451 VDD.n450 3.1505
R287 VDD.n450 VDD.n449 3.1505
R288 VDD.n454 VDD.n453 3.1505
R289 VDD.n453 VDD.n452 3.1505
R290 VDD.n457 VDD.n456 3.1505
R291 VDD.n456 VDD.n455 3.1505
R292 VDD.n460 VDD.n459 3.1505
R293 VDD.n459 VDD.n458 3.1505
R294 VDD.n463 VDD.n462 3.1505
R295 VDD.n462 VDD.n461 3.1505
R296 VDD.n466 VDD.n465 3.1505
R297 VDD.n465 VDD.n464 3.1505
R298 VDD.n469 VDD.n468 3.1505
R299 VDD.n468 VDD.n467 3.1505
R300 VDD.n472 VDD.n471 3.1505
R301 VDD.n471 VDD.n470 3.1505
R302 VDD.n363 VDD.n362 3.1505
R303 VDD.n365 VDD.n364 3.1505
R304 VDD.n368 VDD.n367 3.1505
R305 VDD.n370 VDD.n369 3.1505
R306 VDD.n373 VDD.n372 3.1505
R307 VDD.n375 VDD.n374 3.1505
R308 VDD.n379 VDD.n378 3.1505
R309 VDD.n570 VDD.n541 3.1505
R310 VDD.n585 VDD.n584 3.1505
R311 VDD.n583 VDD.n582 3.1505
R312 VDD.n580 VDD.n579 3.1505
R313 VDD.n578 VDD.n577 3.1505
R314 VDD.n575 VDD.n574 3.1505
R315 VDD.n573 VDD.n572 3.1505
R316 VDD.n589 VDD.n588 3.1505
R317 VDD.n543 VDD.n542 3.1505
R318 VDD.n545 VDD.n544 3.1505
R319 VDD.n547 VDD.n546 3.1505
R320 VDD.n549 VDD.n548 3.1505
R321 VDD.n551 VDD.n550 3.1505
R322 VDD.n553 VDD.n552 3.1505
R323 VDD.n555 VDD.n554 3.1505
R324 VDD.n557 VDD.n556 3.1505
R325 VDD.n559 VDD.n558 3.1505
R326 VDD.n561 VDD.n560 3.1505
R327 VDD.n563 VDD.n562 3.1505
R328 VDD.n565 VDD.n564 3.1505
R329 VDD.n567 VDD.n566 3.1505
R330 VDD.n569 VDD.n568 3.1505
R331 VDD.n31 VDD.n30 3.1505
R332 VDD.n33 VDD.n32 3.1505
R333 VDD.n36 VDD.n35 3.1505
R334 VDD.n40 VDD.n39 3.1505
R335 VDD.n43 VDD.n42 3.1505
R336 VDD.n46 VDD.n45 3.1505
R337 VDD.n28 VDD.n27 3.1505
R338 VDD.n50 VDD.n49 3.1505
R339 VDD.n501 VDD.n500 3.1505
R340 VDD.n500 VDD.n499 3.1505
R341 VDD.n504 VDD.n503 3.1505
R342 VDD.n503 VDD.n502 3.1505
R343 VDD.n507 VDD.n506 3.1505
R344 VDD.n506 VDD.n505 3.1505
R345 VDD.n510 VDD.n509 3.1505
R346 VDD.n509 VDD.n508 3.1505
R347 VDD.n513 VDD.n512 3.1505
R348 VDD.n512 VDD.n511 3.1505
R349 VDD.n516 VDD.n515 3.1505
R350 VDD.n515 VDD.n514 3.1505
R351 VDD.n519 VDD.n518 3.1505
R352 VDD.n518 VDD.n517 3.1505
R353 VDD.n522 VDD.n521 3.1505
R354 VDD.n521 VDD.n520 3.1505
R355 VDD.n525 VDD.n524 3.1505
R356 VDD.n524 VDD.n523 3.1505
R357 VDD.n528 VDD.n527 3.1505
R358 VDD.n527 VDD.n526 3.1505
R359 VDD.n531 VDD.n530 3.1505
R360 VDD.n530 VDD.n529 3.1505
R361 VDD.n534 VDD.n533 3.1505
R362 VDD.n533 VDD.n532 3.1505
R363 VDD.n537 VDD.n536 3.1505
R364 VDD.n536 VDD.n535 3.1505
R365 VDD.n540 VDD.n539 3.1505
R366 VDD.n539 VDD.n538 3.1505
R367 VDD.n648 VDD.n647 3.1505
R368 VDD.n634 VDD.n633 3.1505
R369 VDD.n637 VDD.n636 3.1505
R370 VDD.n639 VDD.n638 3.1505
R371 VDD.n642 VDD.n641 3.1505
R372 VDD.n644 VDD.n643 3.1505
R373 VDD.n632 VDD.n631 3.1505
R374 VDD.n629 VDD.n628 3.1505
R375 VDD.n690 VDD.n689 3.1505
R376 VDD.n688 VDD.n687 3.1505
R377 VDD.n687 VDD.n686 3.1505
R378 VDD.n685 VDD.n684 3.1505
R379 VDD.n684 VDD.n683 3.1505
R380 VDD.n682 VDD.n681 3.1505
R381 VDD.n681 VDD.n680 3.1505
R382 VDD.n679 VDD.n678 3.1505
R383 VDD.n678 VDD.n677 3.1505
R384 VDD.n676 VDD.n675 3.1505
R385 VDD.n675 VDD.n674 3.1505
R386 VDD.n673 VDD.n672 3.1505
R387 VDD.n672 VDD.n671 3.1505
R388 VDD.n670 VDD.n669 3.1505
R389 VDD.n669 VDD.n668 3.1505
R390 VDD.n667 VDD.n666 3.1505
R391 VDD.n666 VDD.n665 3.1505
R392 VDD.n664 VDD.n663 3.1505
R393 VDD.n663 VDD.n662 3.1505
R394 VDD.n661 VDD.n660 3.1505
R395 VDD.n660 VDD.n659 3.1505
R396 VDD.n658 VDD.n657 3.1505
R397 VDD.n657 VDD.n656 3.1505
R398 VDD.n655 VDD.n654 3.1505
R399 VDD.n654 VDD.n653 3.1505
R400 VDD.n652 VDD.n651 3.1505
R401 VDD.n651 VDD.n650 3.1505
R402 VDD.n696 VDD.n695 3.1505
R403 VDD.n698 VDD.n697 3.1505
R404 VDD.n701 VDD.n700 3.1505
R405 VDD.n3 VDD.n2 3.1505
R406 VDD.n593 VDD.n592 3.1505
R407 VDD.n595 VDD.n594 3.1505
R408 VDD.n692 VDD.n691 3.1505
R409 VDD.n598 VDD.n597 3.1505
R410 VDD.n627 VDD.n626 3.1505
R411 VDD.n625 VDD.n624 3.1505
R412 VDD.n623 VDD.n622 3.1505
R413 VDD.n621 VDD.n620 3.1505
R414 VDD.n619 VDD.n618 3.1505
R415 VDD.n617 VDD.n616 3.1505
R416 VDD.n615 VDD.n614 3.1505
R417 VDD.n613 VDD.n612 3.1505
R418 VDD.n611 VDD.n610 3.1505
R419 VDD.n609 VDD.n608 3.1505
R420 VDD.n607 VDD.n606 3.1505
R421 VDD.n605 VDD.n604 3.1505
R422 VDD.n603 VDD.n602 3.1505
R423 VDD.n601 VDD.n600 3.1505
R424 VDD.n600 VDD.n599 3.1505
R425 VDD.n96 VDD.n93 3.07111
R426 VDD.n406 VDD.n403 3.07111
R427 VDD.n25 VDD.n22 3.07111
R428 VDD.n724 VDD.n721 3.07111
R429 VDD.n132 VDD.n131 3.001
R430 VDD.n135 VDD.n134 3.001
R431 VDD.n139 VDD.n138 3.001
R432 VDD.n416 VDD.n415 3.001
R433 VDD.n420 VDD.n419 3.001
R434 VDD.n45 VDD.n44 3.001
R435 VDD.n42 VDD.n41 3.001
R436 VDD.n39 VDD.n38 3.001
R437 VDD.n35 VDD.n34 3.001
R438 VDD.n592 VDD.n591 3.001
R439 VDD.n2 VDD.n0 3.001
R440 VDD.n2 VDD.n1 3.001
R441 VDD.n700 VDD.n699 3.001
R442 VDD.n254 VDD.n253 2.96108
R443 VDD.n477 VDD.n476 2.86102
R444 VDD VDD.n55 2.82941
R445 VDD VDD.n479 2.82941
R446 VDD.n91 VDD.n90 2.64616
R447 VDD.n401 VDD.n400 2.64616
R448 VDD.n20 VDD.n19 2.64616
R449 VDD.n719 VDD.n718 2.64616
R450 VDD.n475 VDD.n384 2.6255
R451 VDD.n278 VDD.n262 2.46744
R452 VDD.n306 VDD.t113 2.41014
R453 VDD.n452 VDD.t125 2.41014
R454 VDD.n520 VDD.t47 2.41014
R455 VDD.n668 VDD.t30 2.41014
R456 VDD.n497 VDD.n496 2.25606
R457 VDD.n157 VDD.n156 2.03336
R458 VDD.n429 VDD.n428 2.03336
R459 VDD.n162 VDD.n161 2.03326
R460 VDD.n167 VDD.n166 2.03326
R461 VDD.n372 VDD.n371 2.03326
R462 VDD.n378 VDD.n377 2.03326
R463 VDD.n588 VDD.n587 2.03326
R464 VDD.n582 VDD.n581 2.03326
R465 VDD.n577 VDD.n576 2.03326
R466 VDD.n572 VDD.n571 2.03326
R467 VDD.n647 VDD.n646 2.03326
R468 VDD.n641 VDD.n640 2.03326
R469 VDD.n636 VDD.n635 2.03326
R470 VDD.n631 VDD.n630 2.03326
R471 VDD.n226 VDD.n210 2.02931
R472 VDD.n146 VDD.n145 1.88586
R473 VDD.n171 VDD.n170 1.87058
R474 VDD.n250 VDD.n249 1.85344
R475 VDD.n93 VDD.t156 1.8205
R476 VDD.n93 VDD.n92 1.8205
R477 VDD.n95 VDD.t135 1.8205
R478 VDD.n95 VDD.n94 1.8205
R479 VDD.n76 VDD.t181 1.8205
R480 VDD.n76 VDD.n75 1.8205
R481 VDD.n79 VDD.t112 1.8205
R482 VDD.n79 VDD.n78 1.8205
R483 VDD.n82 VDD.t110 1.8205
R484 VDD.n82 VDD.n81 1.8205
R485 VDD.n85 VDD.t190 1.8205
R486 VDD.n85 VDD.n84 1.8205
R487 VDD.n88 VDD.t136 1.8205
R488 VDD.n88 VDD.n87 1.8205
R489 VDD.n403 VDD.t144 1.8205
R490 VDD.n403 VDD.n402 1.8205
R491 VDD.n405 VDD.t12 1.8205
R492 VDD.n405 VDD.n404 1.8205
R493 VDD.n386 VDD.t193 1.8205
R494 VDD.n386 VDD.n385 1.8205
R495 VDD.n389 VDD.t132 1.8205
R496 VDD.n389 VDD.n388 1.8205
R497 VDD.n392 VDD.t130 1.8205
R498 VDD.n392 VDD.n391 1.8205
R499 VDD.n395 VDD.t194 1.8205
R500 VDD.n395 VDD.n394 1.8205
R501 VDD.n398 VDD.t149 1.8205
R502 VDD.n398 VDD.n397 1.8205
R503 VDD.n22 VDD.t92 1.8205
R504 VDD.n22 VDD.n21 1.8205
R505 VDD.n24 VDD.t96 1.8205
R506 VDD.n24 VDD.n23 1.8205
R507 VDD.n5 VDD.t22 1.8205
R508 VDD.n5 VDD.n4 1.8205
R509 VDD.n8 VDD.t88 1.8205
R510 VDD.n8 VDD.n7 1.8205
R511 VDD.n11 VDD.t108 1.8205
R512 VDD.n11 VDD.n10 1.8205
R513 VDD.n14 VDD.t102 1.8205
R514 VDD.n14 VDD.n13 1.8205
R515 VDD.n17 VDD.t98 1.8205
R516 VDD.n17 VDD.n16 1.8205
R517 VDD.n721 VDD.t184 1.8205
R518 VDD.n721 VDD.n720 1.8205
R519 VDD.n723 VDD.t84 1.8205
R520 VDD.n723 VDD.n722 1.8205
R521 VDD.n704 VDD.t16 1.8205
R522 VDD.n704 VDD.n703 1.8205
R523 VDD.n707 VDD.t40 1.8205
R524 VDD.n707 VDD.n706 1.8205
R525 VDD.n710 VDD.t37 1.8205
R526 VDD.n710 VDD.n709 1.8205
R527 VDD.n713 VDD.t119 1.8205
R528 VDD.n713 VDD.n712 1.8205
R529 VDD.n716 VDD.t195 1.8205
R530 VDD.n716 VDD.n715 1.8205
R531 VDD.n127 VDD.n126 1.72716
R532 VDD.n411 VDD.n410 1.72716
R533 VDD.n49 VDD.n48 1.72716
R534 VDD.n597 VDD.n596 1.72716
R535 VDD.n142 VDD.n141 1.72703
R536 VDD.n362 VDD.n361 1.72703
R537 VDD.n367 VDD.n366 1.72703
R538 VDD.n423 VDD.n422 1.72703
R539 VDD.n30 VDD.n29 1.72703
R540 VDD.n695 VDD.n694 1.72703
R541 VDD.n280 VDD.n279 1.60323
R542 VDD.n255 VDD.n203 1.52757
R543 VDD.n253 VDD.n252 1.43172
R544 VDD.n77 VDD.n76 1.42427
R545 VDD.n80 VDD.n79 1.42427
R546 VDD.n83 VDD.n82 1.42427
R547 VDD.n86 VDD.n85 1.42427
R548 VDD.n89 VDD.n88 1.42427
R549 VDD.n387 VDD.n386 1.42427
R550 VDD.n390 VDD.n389 1.42427
R551 VDD.n393 VDD.n392 1.42427
R552 VDD.n396 VDD.n395 1.42427
R553 VDD.n399 VDD.n398 1.42427
R554 VDD.n6 VDD.n5 1.42427
R555 VDD.n9 VDD.n8 1.42427
R556 VDD.n12 VDD.n11 1.42427
R557 VDD.n15 VDD.n14 1.42427
R558 VDD.n18 VDD.n17 1.42427
R559 VDD.n705 VDD.n704 1.42427
R560 VDD.n708 VDD.n707 1.42427
R561 VDD.n711 VDD.n710 1.42427
R562 VDD.n714 VDD.n713 1.42427
R563 VDD.n717 VDD.n716 1.42427
R564 VDD.n253 VDD.n226 1.34003
R565 VDD.n384 VDD.n382 1.31777
R566 VDD.n279 VDD.n255 1.30655
R567 VDD.n384 VDD.n383 1.27368
R568 VDD.n497 VDD.n477 1.18161
R569 VDD.n91 VDD.n89 1.16194
R570 VDD.n401 VDD.n399 1.16194
R571 VDD.n20 VDD.n18 1.16194
R572 VDD.n719 VDD.n717 1.16194
R573 VDD.n149 VDD.n148 1.08868
R574 VDD.n48 VDD.n47 0.950516
R575 VDD.n694 VDD.n693 0.950315
R576 VDD.n73 VDD.n72 0.916864
R577 VDD.n277 VDD.n276 0.898937
R578 VDD.n225 VDD.n224 0.898718
R579 VDD.n282 VDD.n281 0.859591
R580 VDD.n170 VDD.n169 0.754483
R581 VDD.n145 VDD.n144 0.745201
R582 VDD.n175 VDD.t65 0.6505
R583 VDD.n175 VDD.n174 0.6505
R584 VDD.n228 VDD.t167 0.6505
R585 VDD.n228 VDD.n227 0.6505
R586 VDD.n80 VDD.n77 0.562605
R587 VDD.n83 VDD.n80 0.562605
R588 VDD.n86 VDD.n83 0.562605
R589 VDD.n89 VDD.n86 0.562605
R590 VDD.n390 VDD.n387 0.562605
R591 VDD.n393 VDD.n390 0.562605
R592 VDD.n396 VDD.n393 0.562605
R593 VDD.n399 VDD.n396 0.562605
R594 VDD.n9 VDD.n6 0.562605
R595 VDD.n12 VDD.n9 0.562605
R596 VDD.n15 VDD.n12 0.562605
R597 VDD.n18 VDD.n15 0.562605
R598 VDD.n708 VDD.n705 0.562605
R599 VDD.n711 VDD.n708 0.562605
R600 VDD.n714 VDD.n711 0.562605
R601 VDD.n717 VDD.n714 0.562605
R602 VDD.n428 VDD.n427 0.560113
R603 VDD.n377 VDD.n376 0.559871
R604 VDD.n587 VDD.n586 0.559871
R605 VDD.n646 VDD.n645 0.559871
R606 VDD.n261 VDD.n260 0.526923
R607 VDD.n209 VDD.n208 0.526923
R608 VDD.n97 VDD.n96 0.418343
R609 VDD.n407 VDD.n406 0.418343
R610 VDD.n26 VDD.n25 0.418343
R611 VDD.n725 VDD.n724 0.418343
R612 VDD.n97 VDD.n91 0.41547
R613 VDD.n407 VDD.n401 0.41547
R614 VDD.n26 VDD.n20 0.41547
R615 VDD.n725 VDD.n719 0.41547
R616 VDD.n278 VDD.n277 0.348354
R617 VDD.n284 VDD.n283 0.286864
R618 VDD.n226 VDD.n225 0.272998
R619 VDD.n201 VDD.n200 0.2719
R620 VDD.n283 VDD.n282 0.229591
R621 VDD.n150 VDD.n149 0.229591
R622 VDD.n71 VDD.n70 0.222053
R623 VDD.n72 VDD.n71 0.222053
R624 VDD.n178 VDD.n177 0.209658
R625 VDD.n231 VDD.n230 0.209419
R626 VDD.n327 VDD.n326 0.185
R627 VDD.n326 VDD.n323 0.185
R628 VDD.n323 VDD.n320 0.185
R629 VDD.n320 VDD.n317 0.185
R630 VDD.n317 VDD.n314 0.185
R631 VDD.n314 VDD.n311 0.185
R632 VDD.n311 VDD.n308 0.185
R633 VDD.n308 VDD.n305 0.185
R634 VDD.n305 VDD.n302 0.185
R635 VDD.n302 VDD.n299 0.185
R636 VDD.n299 VDD.n296 0.185
R637 VDD.n296 VDD.n293 0.185
R638 VDD.n293 VDD.n290 0.185
R639 VDD.n125 VDD.n123 0.185
R640 VDD.n123 VDD.n121 0.185
R641 VDD.n121 VDD.n119 0.185
R642 VDD.n119 VDD.n117 0.185
R643 VDD.n117 VDD.n115 0.185
R644 VDD.n115 VDD.n113 0.185
R645 VDD.n113 VDD.n111 0.185
R646 VDD.n111 VDD.n109 0.185
R647 VDD.n109 VDD.n107 0.185
R648 VDD.n107 VDD.n105 0.185
R649 VDD.n105 VDD.n103 0.185
R650 VDD.n103 VDD.n101 0.185
R651 VDD.n101 VDD.n99 0.185
R652 VDD.n336 VDD.n334 0.185
R653 VDD.n338 VDD.n336 0.185
R654 VDD.n340 VDD.n338 0.185
R655 VDD.n342 VDD.n340 0.185
R656 VDD.n344 VDD.n342 0.185
R657 VDD.n346 VDD.n344 0.185
R658 VDD.n348 VDD.n346 0.185
R659 VDD.n350 VDD.n348 0.185
R660 VDD.n352 VDD.n350 0.185
R661 VDD.n354 VDD.n352 0.185
R662 VDD.n356 VDD.n354 0.185
R663 VDD.n358 VDD.n356 0.185
R664 VDD.n360 VDD.n358 0.185
R665 VDD.n436 VDD.n433 0.185
R666 VDD.n439 VDD.n436 0.185
R667 VDD.n442 VDD.n439 0.185
R668 VDD.n445 VDD.n442 0.185
R669 VDD.n448 VDD.n445 0.185
R670 VDD.n451 VDD.n448 0.185
R671 VDD.n454 VDD.n451 0.185
R672 VDD.n457 VDD.n454 0.185
R673 VDD.n460 VDD.n457 0.185
R674 VDD.n463 VDD.n460 0.185
R675 VDD.n466 VDD.n463 0.185
R676 VDD.n469 VDD.n466 0.185
R677 VDD.n472 VDD.n469 0.185
R678 VDD.n545 VDD.n543 0.185
R679 VDD.n547 VDD.n545 0.185
R680 VDD.n549 VDD.n547 0.185
R681 VDD.n551 VDD.n549 0.185
R682 VDD.n553 VDD.n551 0.185
R683 VDD.n555 VDD.n553 0.185
R684 VDD.n557 VDD.n555 0.185
R685 VDD.n559 VDD.n557 0.185
R686 VDD.n561 VDD.n559 0.185
R687 VDD.n563 VDD.n561 0.185
R688 VDD.n565 VDD.n563 0.185
R689 VDD.n567 VDD.n565 0.185
R690 VDD.n569 VDD.n567 0.185
R691 VDD.n504 VDD.n501 0.185
R692 VDD.n507 VDD.n504 0.185
R693 VDD.n510 VDD.n507 0.185
R694 VDD.n513 VDD.n510 0.185
R695 VDD.n516 VDD.n513 0.185
R696 VDD.n519 VDD.n516 0.185
R697 VDD.n522 VDD.n519 0.185
R698 VDD.n525 VDD.n522 0.185
R699 VDD.n528 VDD.n525 0.185
R700 VDD.n531 VDD.n528 0.185
R701 VDD.n534 VDD.n531 0.185
R702 VDD.n537 VDD.n534 0.185
R703 VDD.n540 VDD.n537 0.185
R704 VDD.n690 VDD.n688 0.185
R705 VDD.n688 VDD.n685 0.185
R706 VDD.n685 VDD.n682 0.185
R707 VDD.n682 VDD.n679 0.185
R708 VDD.n679 VDD.n676 0.185
R709 VDD.n676 VDD.n673 0.185
R710 VDD.n673 VDD.n670 0.185
R711 VDD.n670 VDD.n667 0.185
R712 VDD.n667 VDD.n664 0.185
R713 VDD.n664 VDD.n661 0.185
R714 VDD.n661 VDD.n658 0.185
R715 VDD.n658 VDD.n655 0.185
R716 VDD.n655 VDD.n652 0.185
R717 VDD.n605 VDD.n603 0.185
R718 VDD.n607 VDD.n605 0.185
R719 VDD.n609 VDD.n607 0.185
R720 VDD.n611 VDD.n609 0.185
R721 VDD.n613 VDD.n611 0.185
R722 VDD.n615 VDD.n613 0.185
R723 VDD.n617 VDD.n615 0.185
R724 VDD.n619 VDD.n617 0.185
R725 VDD.n621 VDD.n619 0.185
R726 VDD.n623 VDD.n621 0.185
R727 VDD.n625 VDD.n623 0.185
R728 VDD.n627 VDD.n625 0.185
R729 VDD.n363 VDD.n360 0.172236
R730 VDD.n629 VDD.n627 0.172236
R731 VDD.n69 VDD.n68 0.171026
R732 VDD.n158 VDD.n155 0.164136
R733 VDD.n160 VDD.n158 0.164136
R734 VDD.n163 VDD.n160 0.164136
R735 VDD.n165 VDD.n163 0.164136
R736 VDD.n168 VDD.n165 0.164136
R737 VDD.n172 VDD.n168 0.164136
R738 VDD.n130 VDD.n128 0.164136
R739 VDD.n133 VDD.n130 0.164136
R740 VDD.n136 VDD.n133 0.164136
R741 VDD.n143 VDD.n140 0.164136
R742 VDD.n147 VDD.n143 0.164136
R743 VDD.n414 VDD.n412 0.164136
R744 VDD.n417 VDD.n414 0.164136
R745 VDD.n424 VDD.n421 0.164136
R746 VDD.n426 VDD.n424 0.164136
R747 VDD.n430 VDD.n426 0.164136
R748 VDD.n365 VDD.n363 0.164136
R749 VDD.n368 VDD.n365 0.164136
R750 VDD.n370 VDD.n368 0.164136
R751 VDD.n373 VDD.n370 0.164136
R752 VDD.n375 VDD.n373 0.164136
R753 VDD.n379 VDD.n375 0.164136
R754 VDD.n589 VDD.n585 0.164136
R755 VDD.n585 VDD.n583 0.164136
R756 VDD.n583 VDD.n580 0.164136
R757 VDD.n580 VDD.n578 0.164136
R758 VDD.n578 VDD.n575 0.164136
R759 VDD.n575 VDD.n573 0.164136
R760 VDD.n573 VDD.n570 0.164136
R761 VDD.n50 VDD.n46 0.164136
R762 VDD.n46 VDD.n43 0.164136
R763 VDD.n43 VDD.n40 0.164136
R764 VDD.n36 VDD.n33 0.164136
R765 VDD.n33 VDD.n31 0.164136
R766 VDD.n31 VDD.n28 0.164136
R767 VDD.n632 VDD.n629 0.164136
R768 VDD.n634 VDD.n632 0.164136
R769 VDD.n637 VDD.n634 0.164136
R770 VDD.n639 VDD.n637 0.164136
R771 VDD.n642 VDD.n639 0.164136
R772 VDD.n644 VDD.n642 0.164136
R773 VDD.n648 VDD.n644 0.164136
R774 VDD.n598 VDD.n595 0.164136
R775 VDD.n595 VDD.n593 0.164136
R776 VDD.n593 VDD.n3 0.164136
R777 VDD.n701 VDD.n698 0.164136
R778 VDD.n698 VDD.n696 0.164136
R779 VDD.n696 VDD.n692 0.164136
R780 VDD.n140 VDD.n137 0.161682
R781 VDD.n421 VDD.n418 0.161682
R782 VDD.n37 VDD.n36 0.161682
R783 VDD.n702 VDD.n701 0.161682
R784 VDD.n331 VDD.n147 0.159829
R785 VDD.n412 VDD.n409 0.157591
R786 VDD.n280 VDD.n172 0.155743
R787 VDD.n128 VDD.n125 0.151536
R788 VDD.n601 VDD.n598 0.151536
R789 VDD.n68 VDD.n67 0.143789
R790 VDD.n484 VDD.n483 0.143789
R791 VDD.n210 VDD.n205 0.140912
R792 VDD.n570 VDD.n569 0.137873
R793 VDD.n473 VDD.n472 0.137055
R794 VDD.n476 VDD.n379 0.136132
R795 VDD.n290 VDD.n287 0.1346
R796 VDD.n262 VDD.n257 0.134192
R797 VDD.n137 VDD 0.130885
R798 VDD.n418 VDD 0.130885
R799 VDD.n37 VDD 0.130885
R800 VDD VDD.n702 0.130885
R801 VDD.n334 VDD.n332 0.130485
R802 VDD.n62 VDD.n61 0.127211
R803 VDD.n492 VDD.n489 0.127211
R804 VDD.n272 VDD.n271 0.12598
R805 VDD.n220 VDD.n219 0.12598
R806 VDD.n266 VDD.n265 0.125861
R807 VDD.n214 VDD.n213 0.125861
R808 VDD.n61 VDD.n58 0.123658
R809 VDD.n495 VDD.n492 0.123658
R810 VDD.n433 VDD.n430 0.117173
R811 VDD.n692 VDD.n690 0.117173
R812 VDD.n195 VDD.n192 0.117038
R813 VDD.n192 VDD.n189 0.117038
R814 VDD.n180 VDD.n179 0.117038
R815 VDD.n250 VDD.n248 0.117038
R816 VDD.n248 VDD.n245 0.117038
R817 VDD.n245 VDD.n242 0.117038
R818 VDD.n233 VDD.n232 0.117038
R819 VDD.n328 VDD.n327 0.1139
R820 VDD.n198 VDD.n195 0.1055
R821 VDD.n273 VDD.n270 0.102773
R822 VDD.n270 VDD.n267 0.102773
R823 VDD.n221 VDD.n218 0.102773
R824 VDD.n218 VDD.n215 0.102773
R825 VDD.n603 VDD 0.0968
R826 VDD.n496 VDD.n495 0.0952368
R827 VDD.n590 VDD.n589 0.0921364
R828 VDD VDD.n601 0.0887
R829 VDD.n179 VDD.n176 0.0858846
R830 VDD.n232 VDD.n229 0.0858846
R831 VDD.n186 VDD.n185 0.0835769
R832 VDD.n239 VDD.n238 0.0835769
R833 VDD.n501 VDD.n498 0.0815
R834 VDD.n590 VDD.n540 0.0806
R835 VDD.n652 VDD.n649 0.0788
R836 VDD.n222 VDD.n221 0.0782273
R837 VDD.n67 VDD 0.0774737
R838 VDD.n484 VDD 0.0774737
R839 VDD.n274 VDD.n273 0.0772045
R840 VDD VDD.n257 0.0715526
R841 VDD VDD.n205 0.0715526
R842 VDD.n185 VDD 0.0708846
R843 VDD.n238 VDD 0.0708846
R844 VDD.n498 VDD.n50 0.0705364
R845 VDD.n649 VDD.n648 0.0595727
R846 VDD.n151 VDD.n150 0.0577727
R847 VDD.n267 VDD 0.0526591
R848 VDD.n215 VDD 0.0526591
R849 VDD.n62 VDD 0.0478684
R850 VDD.n489 VDD 0.0478684
R851 VDD.n180 VDD 0.0466538
R852 VDD.n233 VDD 0.0466538
R853 VDD.n279 VDD.n278 0.0423605
R854 VDD VDD.n97 0.0374231
R855 VDD VDD.n407 0.0374231
R856 VDD VDD.n26 0.0374231
R857 VDD VDD.n725 0.0374231
R858 VDD.n189 VDD.n186 0.0339615
R859 VDD.n242 VDD.n239 0.0339615
R860 VDD.n381 VDD.n380 0.0295068
R861 VDD.n382 VDD.n381 0.0295068
R862 VDD.n258 VDD 0.0253684
R863 VDD.n206 VDD 0.0253684
R864 VDD.n475 VDD.n474 0.0193182
R865 VDD.n276 VDD.n275 0.0178864
R866 VDD.n224 VDD.n223 0.0178864
R867 VDD.n202 VDD.n199 0.0178077
R868 VDD.n264 VDD 0.0148182
R869 VDD.n212 VDD 0.0148182
R870 VDD.n199 VDD.n198 0.0120385
R871 VDD.n476 VDD.n475 0.011585
R872 VDD.n332 VDD.n74 0.0103779
R873 VDD.n255 VDD.n254 0.0099186
R874 VDD.n275 VDD.n274 0.00868182
R875 VDD.n223 VDD.n222 0.00765909
R876 VDD.n252 VDD.n250 0.00742767
R877 VDD.n409 VDD.n408 0.00704545
R878 VDD.n285 VDD.n280 0.00672312
R879 VDD.n331 VDD.n330 0.00590945
R880 VDD.n286 VDD.n285 0.00459091
R881 VDD.n287 VDD.n286 0.00377273
R882 VDD.n329 VDD.n328 0.00377273
R883 VDD.n137 VDD.n136 0.00295455
R884 VDD.n418 VDD.n417 0.00295455
R885 VDD.n40 VDD.n37 0.00295455
R886 VDD.n702 VDD.n3 0.00295455
R887 VDD.n203 VDD.n202 0.00165385
R888 VDD.n330 VDD.n329 0.00131818
R889 VDD.n474 VDD.n473 0.00131818
R890 OUTB.n9 OUTB.n3 3.58485
R891 OUTB.n8 OUTB.n7 3.58485
R892 OUTB.n9 OUTB.n1 3.32833
R893 OUTB.n8 OUTB.n5 3.32833
R894 OUTB.n3 OUTB.t6 1.1705
R895 OUTB.n3 OUTB.n2 1.1705
R896 OUTB.n7 OUTB.t7 1.1705
R897 OUTB.n7 OUTB.n6 1.1705
R898 OUTB.n9 OUTB.n8 0.68137
R899 OUTB.n1 OUTB.t4 0.6505
R900 OUTB.n1 OUTB.n0 0.6505
R901 OUTB.n5 OUTB.t5 0.6505
R902 OUTB.n5 OUTB.n4 0.6505
R903 OUTB OUTB.n9 0.297728
R904 a_2201_958.t2 a_2201_958.n5 22.8782
R905 a_2201_958.n6 a_2201_958.t2 22.4219
R906 a_2201_958.n3 a_2201_958.t16 22.2916
R907 a_2201_958.n5 a_2201_958.n4 14.0791
R908 a_2201_958.n4 a_2201_958.n3 14.0791
R909 a_2201_958.n7 a_2201_958.n6 14.0791
R910 a_2201_958.n2 a_2201_958.t4 11.3416
R911 a_2201_958.n6 a_2201_958.t0 8.34336
R912 a_2201_958.n7 a_2201_958.t6 8.34336
R913 a_2201_958.n5 a_2201_958.t12 8.213
R914 a_2201_958.n4 a_2201_958.t13 8.213
R915 a_2201_958.n3 a_2201_958.t15 8.213
R916 a_2201_958.n0 a_2201_958.n7 8.17193
R917 a_2201_958.n1 a_2201_958.n2 4.0005
R918 a_2201_958.n0 a_2201_958.n9 3.63045
R919 a_2201_958.n18 a_2201_958.n1 2.89398
R920 a_2201_958.n14 a_2201_958.n11 2.26392
R921 a_2201_958.n9 a_2201_958.t3 1.8205
R922 a_2201_958.n9 a_2201_958.n8 1.8205
R923 a_2201_958.t7 a_2201_958.n18 1.8205
R924 a_2201_958.n18 a_2201_958.n17 1.8205
R925 a_2201_958.n11 a_2201_958.t10 1.6385
R926 a_2201_958.n11 a_2201_958.n10 1.6385
R927 a_2201_958.n13 a_2201_958.t8 1.6385
R928 a_2201_958.n13 a_2201_958.n12 1.6385
R929 a_2201_958.n2 a_2201_958.n16 1.62996
R930 a_2201_958.n14 a_2201_958.n13 1.4936
R931 a_2201_958.n1 a_2201_958.n15 1.22554
R932 a_2201_958.n15 a_2201_958.n14 1.18673
R933 a_2201_958.n1 a_2201_958.n0 0.1505
R934 Delay_Cell_mag_2.IN.n20 Delay_Cell_mag_2.IN.t16 22.2916
R935 Delay_Cell_mag_2.IN.n4 Delay_Cell_mag_2.IN.t14 22.1612
R936 Delay_Cell_mag_2.IN.n23 Delay_Cell_mag_2.IN.t19 21.774
R937 Delay_Cell_mag_2.IN.t16 Delay_Cell_mag_2.IN.n19 17.311
R938 Delay_Cell_mag_2.IN.n6 Delay_Cell_mag_2.IN.t10 15.1219
R939 Delay_Cell_mag_2.IN.n21 Delay_Cell_mag_2.IN.n20 14.0791
R940 Delay_Cell_mag_2.IN.n22 Delay_Cell_mag_2.IN.n21 14.0791
R941 Delay_Cell_mag_2.IN.n5 Delay_Cell_mag_2.IN.n4 14.0791
R942 Delay_Cell_mag_2.IN.n24 Delay_Cell_mag_2.IN.n23 12.7222
R943 Delay_Cell_mag_2.IN.n25 Delay_Cell_mag_2.IN.t18 11.9934
R944 Delay_Cell_mag_2.IN.n25 Delay_Cell_mag_2.IN.n24 9.78115
R945 Delay_Cell_mag_2.IN.n20 Delay_Cell_mag_2.IN.t20 8.213
R946 Delay_Cell_mag_2.IN.n21 Delay_Cell_mag_2.IN.t22 8.213
R947 Delay_Cell_mag_2.IN.n22 Delay_Cell_mag_2.IN.t24 8.213
R948 Delay_Cell_mag_2.IN.n5 Delay_Cell_mag_2.IN.t12 8.08264
R949 Delay_Cell_mag_2.IN.n4 Delay_Cell_mag_2.IN.t8 8.08264
R950 Delay_Cell_mag_2.IN.n6 Delay_Cell_mag_2.IN.n5 7.03979
R951 Delay_Cell_mag_2.IN.n23 Delay_Cell_mag_2.IN.t25 6.51836
R952 Delay_Cell_mag_2.IN.n24 Delay_Cell_mag_2.IN.t21 6.51836
R953 Delay_Cell_mag_2.IN.n14 Delay_Cell_mag_2.IN.n13 4.70398
R954 Delay_Cell_mag_2.IN.n15 Delay_Cell_mag_2.IN.n14 4.4843
R955 Delay_Cell_mag_2.IN.n7 Delay_Cell_mag_2.IN.n6 4.0005
R956 Delay_Cell_mag_2.IN.n19 Delay_Cell_mag_2.IN.n1 3.3342
R957 Delay_Cell_mag_2.IN.n14 Delay_Cell_mag_2.IN.n11 3.1505
R958 Delay_Cell_mag_2.IN.n7 Delay_Cell_mag_2.IN.n3 2.94411
R959 Delay_Cell_mag_2.IN.n19 Delay_Cell_mag_2.IN.n18 2.9292
R960 Delay_Cell_mag_2.IN Delay_Cell_mag_2.IN.n22 2.69696
R961 Delay_Cell_mag_2.IN.n15 Delay_Cell_mag_2.IN.n9 2.6005
R962 Delay_Cell_mag_2.IN Delay_Cell_mag_2.IN.n25 2.10481
R963 Delay_Cell_mag_2.IN.n1 Delay_Cell_mag_2.IN.t9 1.8205
R964 Delay_Cell_mag_2.IN.n1 Delay_Cell_mag_2.IN.n0 1.8205
R965 Delay_Cell_mag_2.IN.n9 Delay_Cell_mag_2.IN.t1 1.8205
R966 Delay_Cell_mag_2.IN.n9 Delay_Cell_mag_2.IN.n8 1.8205
R967 Delay_Cell_mag_2.IN.n3 Delay_Cell_mag_2.IN.t11 1.8205
R968 Delay_Cell_mag_2.IN.n3 Delay_Cell_mag_2.IN.n2 1.8205
R969 Delay_Cell_mag_2.IN.n18 Delay_Cell_mag_2.IN.t0 1.8205
R970 Delay_Cell_mag_2.IN.n18 Delay_Cell_mag_2.IN.n17 1.8205
R971 Delay_Cell_mag_2.IN.n11 Delay_Cell_mag_2.IN.t4 1.6385
R972 Delay_Cell_mag_2.IN.n11 Delay_Cell_mag_2.IN.n10 1.6385
R973 Delay_Cell_mag_2.IN.n13 Delay_Cell_mag_2.IN.t6 1.6385
R974 Delay_Cell_mag_2.IN.n13 Delay_Cell_mag_2.IN.n12 1.6385
R975 Delay_Cell_mag_2.IN.n19 Delay_Cell_mag_2.IN.n16 0.845717
R976 Delay_Cell_mag_2.IN.n16 Delay_Cell_mag_2.IN.n7 0.335065
R977 Delay_Cell_mag_2.IN.n16 Delay_Cell_mag_2.IN.n15 0.329196
R978 a_8644_n2780.t3 a_8644_n2780.n5 22.8782
R979 a_8644_n2780.n6 a_8644_n2780.t3 22.4219
R980 a_8644_n2780.n3 a_8644_n2780.t14 22.2916
R981 a_8644_n2780.n5 a_8644_n2780.n4 14.0791
R982 a_8644_n2780.n4 a_8644_n2780.n3 14.0791
R983 a_8644_n2780.n7 a_8644_n2780.n6 14.0791
R984 a_8644_n2780.n1 a_8644_n2780.t5 11.3416
R985 a_8644_n2780.n6 a_8644_n2780.t9 8.34336
R986 a_8644_n2780.n7 a_8644_n2780.t7 8.34336
R987 a_8644_n2780.n5 a_8644_n2780.t15 8.213
R988 a_8644_n2780.n4 a_8644_n2780.t17 8.213
R989 a_8644_n2780.n3 a_8644_n2780.t13 8.213
R990 a_8644_n2780.n2 a_8644_n2780.n7 8.17193
R991 a_8644_n2780.n0 a_8644_n2780.n1 4.0005
R992 a_8644_n2780.n17 a_8644_n2780.n2 3.63045
R993 a_8644_n2780.n0 a_8644_n2780.n9 2.89398
R994 a_8644_n2780.n14 a_8644_n2780.n11 2.26392
R995 a_8644_n2780.n9 a_8644_n2780.t8 1.8205
R996 a_8644_n2780.n9 a_8644_n2780.n8 1.8205
R997 a_8644_n2780.n17 a_8644_n2780.t4 1.8205
R998 a_8644_n2780.n18 a_8644_n2780.n17 1.8205
R999 a_8644_n2780.n11 a_8644_n2780.t2 1.6385
R1000 a_8644_n2780.n11 a_8644_n2780.n10 1.6385
R1001 a_8644_n2780.n13 a_8644_n2780.t11 1.6385
R1002 a_8644_n2780.n13 a_8644_n2780.n12 1.6385
R1003 a_8644_n2780.n1 a_8644_n2780.n16 1.62996
R1004 a_8644_n2780.n14 a_8644_n2780.n13 1.4936
R1005 a_8644_n2780.n0 a_8644_n2780.n15 1.22554
R1006 a_8644_n2780.n15 a_8644_n2780.n14 1.18673
R1007 a_8644_n2780.n2 a_8644_n2780.n0 0.1505
R1008 Delay_Cell_mag_2.OUT.n13 Delay_Cell_mag_2.OUT.t20 22.3568
R1009 Delay_Cell_mag_2.OUT.n2 Delay_Cell_mag_2.OUT.t7 22.096
R1010 Delay_Cell_mag_2.OUT.n12 Delay_Cell_mag_2.OUT.t18 19.4889
R1011 Delay_Cell_mag_2.OUT.n25 Delay_Cell_mag_2.OUT.t26 19.1891
R1012 Delay_Cell_mag_2.OUT.n26 Delay_Cell_mag_2.OUT.t21 19.1891
R1013 Delay_Cell_mag_2.OUT.n27 Delay_Cell_mag_2.OUT.t23 19.1891
R1014 Delay_Cell_mag_2.OUT.n28 Delay_Cell_mag_2.OUT.t22 18.6676
R1015 Delay_Cell_mag_2.OUT.n26 Delay_Cell_mag_2.OUT.n25 16.9365
R1016 Delay_Cell_mag_2.OUT.n27 Delay_Cell_mag_2.OUT.n26 16.9365
R1017 Delay_Cell_mag_2.OUT.n28 Delay_Cell_mag_2.OUT.n27 16.6457
R1018 Delay_Cell_mag_2.OUT.n3 Delay_Cell_mag_2.OUT.n2 14.0791
R1019 Delay_Cell_mag_2.OUT.n4 Delay_Cell_mag_2.OUT.n3 14.0791
R1020 Delay_Cell_mag_2.OUT.n25 Delay_Cell_mag_2.OUT.t19 11.6805
R1021 Delay_Cell_mag_2.OUT.n26 Delay_Cell_mag_2.OUT.t28 11.6805
R1022 Delay_Cell_mag_2.OUT.n27 Delay_Cell_mag_2.OUT.t17 11.6805
R1023 Delay_Cell_mag_2.OUT.n28 Delay_Cell_mag_2.OUT.t29 11.4719
R1024 Delay_Cell_mag_2.OUT.n14 Delay_Cell_mag_2.OUT.n13 9.33211
R1025 Delay_Cell_mag_2.OUT.n13 Delay_Cell_mag_2.OUT.t24 8.27818
R1026 Delay_Cell_mag_2.OUT.n11 Delay_Cell_mag_2.OUT.t16 8.27818
R1027 Delay_Cell_mag_2.OUT.n2 Delay_Cell_mag_2.OUT.t3 8.01746
R1028 Delay_Cell_mag_2.OUT.n3 Delay_Cell_mag_2.OUT.t9 8.01746
R1029 Delay_Cell_mag_2.OUT.n4 Delay_Cell_mag_2.OUT.t5 8.01746
R1030 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.OUT.n28 7.18457
R1031 Delay_Cell_mag_2.OUT.n0 Delay_Cell_mag_2.OUT 5.23607
R1032 Delay_Cell_mag_2.OUT.n19 Delay_Cell_mag_2.OUT.n18 4.67659
R1033 Delay_Cell_mag_2.OUT.n1 Delay_Cell_mag_2.OUT.n19 3.51328
R1034 Delay_Cell_mag_2.OUT.n24 Delay_Cell_mag_2.OUT.n6 3.20507
R1035 Delay_Cell_mag_2.OUT.n19 Delay_Cell_mag_2.OUT.n16 3.1505
R1036 Delay_Cell_mag_2.OUT.n21 Delay_Cell_mag_2.OUT.n8 3.02311
R1037 Delay_Cell_mag_2.OUT.n24 Delay_Cell_mag_2.OUT.n23 2.98985
R1038 Delay_Cell_mag_2.OUT.n12 Delay_Cell_mag_2.OUT.n11 2.86836
R1039 Delay_Cell_mag_2.OUT.n0 Delay_Cell_mag_2.OUT.n4 2.6373
R1040 Delay_Cell_mag_2.OUT.n20 Delay_Cell_mag_2.OUT.n10 2.6005
R1041 Delay_Cell_mag_2.OUT.n1 Delay_Cell_mag_2.OUT.n12 2.11815
R1042 Delay_Cell_mag_2.OUT.n6 Delay_Cell_mag_2.OUT.t2 1.8205
R1043 Delay_Cell_mag_2.OUT.n6 Delay_Cell_mag_2.OUT.n5 1.8205
R1044 Delay_Cell_mag_2.OUT.n10 Delay_Cell_mag_2.OUT.t0 1.8205
R1045 Delay_Cell_mag_2.OUT.n10 Delay_Cell_mag_2.OUT.n9 1.8205
R1046 Delay_Cell_mag_2.OUT.n8 Delay_Cell_mag_2.OUT.t8 1.8205
R1047 Delay_Cell_mag_2.OUT.n8 Delay_Cell_mag_2.OUT.n7 1.8205
R1048 Delay_Cell_mag_2.OUT.n23 Delay_Cell_mag_2.OUT.t10 1.8205
R1049 Delay_Cell_mag_2.OUT.n23 Delay_Cell_mag_2.OUT.n22 1.8205
R1050 Delay_Cell_mag_2.OUT.n16 Delay_Cell_mag_2.OUT.t15 1.6385
R1051 Delay_Cell_mag_2.OUT.n16 Delay_Cell_mag_2.OUT.n15 1.6385
R1052 Delay_Cell_mag_2.OUT.n18 Delay_Cell_mag_2.OUT.t12 1.6385
R1053 Delay_Cell_mag_2.OUT.n18 Delay_Cell_mag_2.OUT.n17 1.6385
R1054 Delay_Cell_mag_2.OUT.n1 Delay_Cell_mag_2.OUT.n14 1.50108
R1055 Delay_Cell_mag_2.OUT.n20 Delay_Cell_mag_2.OUT.n1 1.32596
R1056 Delay_Cell_mag_2.OUT.n24 Delay_Cell_mag_2.OUT.n21 0.826273
R1057 Delay_Cell_mag_2.OUT.n21 Delay_Cell_mag_2.OUT.n20 0.640283
R1058 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.OUT.n0 0.156737
R1059 Delay_Cell_mag_2.OUT.n0 Delay_Cell_mag_2.OUT.n24 0.128582
R1060 Delay_Cell_mag_2.OUTB.n20 Delay_Cell_mag_2.OUTB.t26 22.2916
R1061 Delay_Cell_mag_2.OUTB.n4 Delay_Cell_mag_2.OUTB.t14 22.1612
R1062 Delay_Cell_mag_2.OUTB.n23 Delay_Cell_mag_2.OUTB.t28 19.1891
R1063 Delay_Cell_mag_2.OUTB.n24 Delay_Cell_mag_2.OUTB.t20 19.1891
R1064 Delay_Cell_mag_2.OUTB.n25 Delay_Cell_mag_2.OUTB.t24 19.1891
R1065 Delay_Cell_mag_2.OUTB.n26 Delay_Cell_mag_2.OUTB.t21 18.6676
R1066 Delay_Cell_mag_2.OUTB.t26 Delay_Cell_mag_2.OUTB.n19 17.311
R1067 Delay_Cell_mag_2.OUTB.n24 Delay_Cell_mag_2.OUTB.n23 16.9365
R1068 Delay_Cell_mag_2.OUTB.n25 Delay_Cell_mag_2.OUTB.n24 16.9365
R1069 Delay_Cell_mag_2.OUTB.n26 Delay_Cell_mag_2.OUTB.n25 16.6457
R1070 Delay_Cell_mag_2.OUTB.n6 Delay_Cell_mag_2.OUTB.t12 15.1219
R1071 Delay_Cell_mag_2.OUTB.n21 Delay_Cell_mag_2.OUTB.n20 14.0791
R1072 Delay_Cell_mag_2.OUTB.n22 Delay_Cell_mag_2.OUTB.n21 14.0791
R1073 Delay_Cell_mag_2.OUTB.n5 Delay_Cell_mag_2.OUTB.n4 14.0791
R1074 Delay_Cell_mag_2.OUTB.n23 Delay_Cell_mag_2.OUTB.t23 11.6805
R1075 Delay_Cell_mag_2.OUTB.n24 Delay_Cell_mag_2.OUTB.t16 11.6805
R1076 Delay_Cell_mag_2.OUTB.n25 Delay_Cell_mag_2.OUTB.t19 11.6805
R1077 Delay_Cell_mag_2.OUTB.n26 Delay_Cell_mag_2.OUTB.t18 11.4719
R1078 Delay_Cell_mag_2.OUTB.n20 Delay_Cell_mag_2.OUTB.t29 8.213
R1079 Delay_Cell_mag_2.OUTB.n21 Delay_Cell_mag_2.OUTB.t25 8.213
R1080 Delay_Cell_mag_2.OUTB.n22 Delay_Cell_mag_2.OUTB.t27 8.213
R1081 Delay_Cell_mag_2.OUTB.n5 Delay_Cell_mag_2.OUTB.t10 8.08264
R1082 Delay_Cell_mag_2.OUTB.n4 Delay_Cell_mag_2.OUTB.t8 8.08264
R1083 Delay_Cell_mag_2.OUTB Delay_Cell_mag_2.OUTB.n26 7.24687
R1084 Delay_Cell_mag_2.OUTB.n6 Delay_Cell_mag_2.OUTB.n5 7.03979
R1085 Delay_Cell_mag_2.OUTB.n14 Delay_Cell_mag_2.OUTB.n13 4.70398
R1086 Delay_Cell_mag_2.OUTB.n15 Delay_Cell_mag_2.OUTB.n14 4.4843
R1087 Delay_Cell_mag_2.OUTB.n7 Delay_Cell_mag_2.OUTB.n6 4.0005
R1088 Delay_Cell_mag_2.OUTB.n19 Delay_Cell_mag_2.OUTB.n1 3.3342
R1089 Delay_Cell_mag_2.OUTB.n14 Delay_Cell_mag_2.OUTB.n11 3.1505
R1090 Delay_Cell_mag_2.OUTB.n7 Delay_Cell_mag_2.OUTB.n3 2.94411
R1091 Delay_Cell_mag_2.OUTB.n19 Delay_Cell_mag_2.OUTB.n18 2.9292
R1092 Delay_Cell_mag_2.OUTB Delay_Cell_mag_2.OUTB.n22 2.70347
R1093 Delay_Cell_mag_2.OUTB.n15 Delay_Cell_mag_2.OUTB.n9 2.6005
R1094 Delay_Cell_mag_2.OUTB.n1 Delay_Cell_mag_2.OUTB.t9 1.8205
R1095 Delay_Cell_mag_2.OUTB.n1 Delay_Cell_mag_2.OUTB.n0 1.8205
R1096 Delay_Cell_mag_2.OUTB.n9 Delay_Cell_mag_2.OUTB.t5 1.8205
R1097 Delay_Cell_mag_2.OUTB.n9 Delay_Cell_mag_2.OUTB.n8 1.8205
R1098 Delay_Cell_mag_2.OUTB.n3 Delay_Cell_mag_2.OUTB.t13 1.8205
R1099 Delay_Cell_mag_2.OUTB.n3 Delay_Cell_mag_2.OUTB.n2 1.8205
R1100 Delay_Cell_mag_2.OUTB.n18 Delay_Cell_mag_2.OUTB.t7 1.8205
R1101 Delay_Cell_mag_2.OUTB.n18 Delay_Cell_mag_2.OUTB.n17 1.8205
R1102 Delay_Cell_mag_2.OUTB.n11 Delay_Cell_mag_2.OUTB.t2 1.6385
R1103 Delay_Cell_mag_2.OUTB.n11 Delay_Cell_mag_2.OUTB.n10 1.6385
R1104 Delay_Cell_mag_2.OUTB.n13 Delay_Cell_mag_2.OUTB.t0 1.6385
R1105 Delay_Cell_mag_2.OUTB.n13 Delay_Cell_mag_2.OUTB.n12 1.6385
R1106 Delay_Cell_mag_2.OUTB.n19 Delay_Cell_mag_2.OUTB.n16 0.845717
R1107 Delay_Cell_mag_2.OUTB.n16 Delay_Cell_mag_2.OUTB.n7 0.335065
R1108 Delay_Cell_mag_2.OUTB.n16 Delay_Cell_mag_2.OUTB.n15 0.329196
R1109 VSS.n1731 VSS.t106 1075.7
R1110 VSS.n216 VSS.n215 513.072
R1111 VSS.n1618 VSS.n1617 391.741
R1112 VSS.n280 VSS.n279 372.031
R1113 VSS.n1698 VSS.n1697 302.113
R1114 VSS.n669 VSS.n668 254.78
R1115 VSS.n1726 VSS.t10 230.024
R1116 VSS.n1732 VSS.n1731 226.314
R1117 VSS.n1565 VSS.t52 218.702
R1118 VSS.n24 VSS.n23 218.161
R1119 VSS.n4 VSS.n3 198.471
R1120 VSS.n757 VSS.n756 172.927
R1121 VSS.n131 VSS.t82 167.84
R1122 VSS.n859 VSS.n858 159.599
R1123 VSS.n451 VSS.n450 149.141
R1124 VSS.n1415 VSS.n1414 147.409
R1125 VSS.n414 VSS.t18 144.998
R1126 VSS.n659 VSS.t35 144.998
R1127 VSS.n740 VSS.n739 134.505
R1128 VSS.n1317 VSS.t54 132.238
R1129 VSS.n417 VSS.t2 122.213
R1130 VSS.n656 VSS.t4 122.213
R1131 VSS.n1493 VSS.n1492 112.555
R1132 VSS.n267 VSS.n266 100.873
R1133 VSS.n420 VSS.t0 99.4269
R1134 VSS.n653 VSS.t7 99.4269
R1135 VSS.n1056 VSS.t57 93.7031
R1136 VSS.n468 VSS.t63 93.7031
R1137 VSS.n423 VSS.t3 76.6417
R1138 VSS.n650 VSS.t6 76.6417
R1139 VSS.n1345 VSS.n1344 76.2916
R1140 VSS.n108 VSS.n107 73.1516
R1141 VSS.n504 VSS.t121 64.3569
R1142 VSS.n514 VSS.t115 61.1391
R1143 VSS.n441 VSS.t19 60.0706
R1144 VSS.n632 VSS.t36 60.0706
R1145 VSS.n426 VSS.t1 53.8565
R1146 VSS.n647 VSS.t5 53.8565
R1147 VSS.n1208 VSS.n1207 53.2307
R1148 VSS.n730 VSS.t8 51.6126
R1149 VSS.n330 VSS.t34 51.5878
R1150 VSS.n963 VSS.t102 51.2592
R1151 VSS.n398 VSS.n397 45.5709
R1152 VSS.n815 VSS.t9 45.3566
R1153 VSS.n1197 VSS.t27 45.3448
R1154 VSS.n1483 VSS.t33 45.3348
R1155 VSS.n1190 VSS.n1189 45.1394
R1156 VSS.n1014 VSS.t94 45.1394
R1157 VSS.n1099 VSS.n1098 39.3568
R1158 VSS.n438 VSS.t15 37.2854
R1159 VSS.n635 VSS.t113 37.2854
R1160 VSS.n1335 VSS.t80 35.603
R1161 VSS.n727 VSS.t20 34.4086
R1162 VSS.n1434 VSS.n1433 34.392
R1163 VSS.n333 VSS.t40 34.392
R1164 VSS.n429 VSS.t14 31.0712
R1165 VSS.n644 VSS.t50 31.0712
R1166 VSS.n872 VSS.n871 29.7166
R1167 VSS.n1059 VSS.t65 29.5908
R1168 VSS.n471 VSS.t60 29.5908
R1169 VSS.n1203 VSS.t21 29.5728
R1170 VSS.n818 VSS.t105 28.1526
R1171 VSS.n1480 VSS.t125 28.139
R1172 VSS.n1256 VSS.n1255 25.5911
R1173 VSS.n827 VSS.t44 23.4606
R1174 VSS.n1471 VSS.t32 23.4493
R1175 VSS.n507 VSS.t118 22.5253
R1176 VSS.n999 VSS.t29 20.5182
R1177 VSS.n107 VSS.n106 20.3448
R1178 VSS.n511 VSS.t123 19.3074
R1179 VSS.n724 VSS.t37 17.2045
R1180 VSS.n719 VSS.t13 17.2045
R1181 VSS.n336 VSS.t41 17.1963
R1182 VSS.n341 VSS.t39 17.1963
R1183 VSS.n953 VSS.n952 16.7582
R1184 VSS.n435 VSS.t16 14.5002
R1185 VSS.n638 VSS.t111 14.5002
R1186 VSS.n821 VSS.t104 10.9485
R1187 VSS.n1477 VSS.t114 10.9433
R1188 VSS.n971 VSS.n970 10.8437
R1189 VSS.n432 VSS.t17 8.28603
R1190 VSS.n641 VSS.t112 8.28603
R1191 VSS.n824 VSS.t108 6.25652
R1192 VSS.n1474 VSS.t31 6.25351
R1193 VSS.n463 VSS.n462 5.99763
R1194 VSS.n297 VSS.n296 5.99763
R1195 VSS.n782 VSS.n781 5.99763
R1196 VSS.n599 VSS.n598 5.99763
R1197 VSS.n1568 VSS.t53 5.80213
R1198 VSS.n124 VSS.t81 5.80213
R1199 VSS.n1558 VSS.n90 5.80209
R1200 VSS.n134 VSS.n96 5.80209
R1201 VSS VSS.t107 5.6909
R1202 VSS VSS.t11 5.6909
R1203 VSS.n517 VSS.n501 5.15437
R1204 VSS.n1055 VSS.n1039 5.15437
R1205 VSS VSS.t122 5.11524
R1206 VSS VSS.t64 5.11524
R1207 VSS.n465 VSS.t79 5.0898
R1208 VSS.n299 VSS.t76 5.0898
R1209 VSS.n784 VSS.t45 5.0898
R1210 VSS.n601 VSS.t51 5.0898
R1211 VSS.n1206 VSS.n1179 4.79593
R1212 VSS.n1185 VSS.t30 4.79593
R1213 VSS.n1284 VSS.n1280 4.79593
R1214 VSS.n969 VSS.t103 4.79593
R1215 VSS VSS.n1181 3.60246
R1216 VSS VSS.n951 3.60246
R1217 VSS.n510 VSS.n503 3.51637
R1218 VSS.n1062 VSS.n1038 3.51637
R1219 VSS.n463 VSS.n461 3.51441
R1220 VSS.n464 VSS.n459 3.51441
R1221 VSS.n297 VSS.n295 3.51441
R1222 VSS.n298 VSS.n293 3.51441
R1223 VSS.n782 VSS.n780 3.51441
R1224 VSS.n783 VSS.n778 3.51441
R1225 VSS.n599 VSS.n597 3.51441
R1226 VSS.n600 VSS.n595 3.51441
R1227 VSS.n1025 VSS.n1024 3.00849
R1228 VSS.n1028 VSS.n1027 3.00849
R1229 VSS.n490 VSS.n489 3.00849
R1230 VSS.n960 VSS.t97 2.95773
R1231 VSS.n1193 VSS.t24 2.95773
R1232 VSS.n743 VSS.n674 2.60693
R1233 VSS.n74 VSS.n4 2.60693
R1234 VSS.n217 VSS.n216 2.60693
R1235 VSS.n320 VSS.n301 2.60693
R1236 VSS.n1364 VSS.n1363 2.60371
R1237 VSS.n907 VSS.n870 2.60371
R1238 VSS.n527 VSS.n526 2.60371
R1239 VSS.n1606 VSS.n86 2.60343
R1240 VSS.n1524 VSS.n92 2.60343
R1241 VSS.n1101 VSS.n1100 2.60243
R1242 VSS.n874 VSS.n873 2.60243
R1243 VSS.n1078 VSS.n587 2.60179
R1244 VSS.n854 VSS.n770 2.60179
R1245 VSS.n1446 VSS.n1439 2.60179
R1246 VSS.n404 VSS.n403 2.60179
R1247 VSS.n1572 VSS.n89 2.60148
R1248 VSS.n120 VSS.n119 2.60148
R1249 VSS.n1667 VSS.n1666 2.6005
R1250 VSS.n1674 VSS.n1673 2.6005
R1251 VSS.n1670 VSS.n1669 2.6005
R1252 VSS.n1636 VSS.n1635 2.6005
R1253 VSS.n1635 VSS.n1634 2.6005
R1254 VSS.n1633 VSS.n1632 2.6005
R1255 VSS.n1632 VSS.n1631 2.6005
R1256 VSS.n1630 VSS.n1629 2.6005
R1257 VSS.n1629 VSS.n1628 2.6005
R1258 VSS.n1627 VSS.n1626 2.6005
R1259 VSS.n1626 VSS.n1625 2.6005
R1260 VSS.n1639 VSS.n1638 2.6005
R1261 VSS.n1638 VSS.n1637 2.6005
R1262 VSS.n1642 VSS.n1641 2.6005
R1263 VSS.n1641 VSS.n1640 2.6005
R1264 VSS.n1646 VSS.n1645 2.6005
R1265 VSS.n1645 VSS.n1644 2.6005
R1266 VSS.n1664 VSS.n1663 2.6005
R1267 VSS.n1660 VSS.n1659 2.6005
R1268 VSS.n1103 VSS.n1102 2.6005
R1269 VSS.n1105 VSS.n1104 2.6005
R1270 VSS.n1107 VSS.n1106 2.6005
R1271 VSS.n1109 VSS.n1108 2.6005
R1272 VSS.n1111 VSS.n1110 2.6005
R1273 VSS.n1113 VSS.n1112 2.6005
R1274 VSS.n1115 VSS.n1114 2.6005
R1275 VSS.n1117 VSS.n1116 2.6005
R1276 VSS.n1119 VSS.n1118 2.6005
R1277 VSS.n1121 VSS.n1120 2.6005
R1278 VSS.n1123 VSS.n1122 2.6005
R1279 VSS.n1125 VSS.n1124 2.6005
R1280 VSS.n1127 VSS.n1126 2.6005
R1281 VSS.n1129 VSS.n1128 2.6005
R1282 VSS.n1131 VSS.n1130 2.6005
R1283 VSS.n1133 VSS.n1132 2.6005
R1284 VSS.n694 VSS.n675 2.6005
R1285 VSS.n742 VSS.n741 2.6005
R1286 VSS.n741 VSS.n740 2.6005
R1287 VSS.n738 VSS.n737 2.6005
R1288 VSS.n737 VSS.n736 2.6005
R1289 VSS.n735 VSS.n734 2.6005
R1290 VSS.n734 VSS.n733 2.6005
R1291 VSS.n732 VSS.n731 2.6005
R1292 VSS.n731 VSS.n730 2.6005
R1293 VSS.n729 VSS.n728 2.6005
R1294 VSS.n728 VSS.n727 2.6005
R1295 VSS.n726 VSS.n725 2.6005
R1296 VSS.n725 VSS.n724 2.6005
R1297 VSS.n723 VSS.n722 2.6005
R1298 VSS.n722 VSS.t12 2.6005
R1299 VSS.n721 VSS.n720 2.6005
R1300 VSS.n720 VSS.n719 2.6005
R1301 VSS.n718 VSS.n717 2.6005
R1302 VSS.n717 VSS.n716 2.6005
R1303 VSS.n715 VSS.n714 2.6005
R1304 VSS.n714 VSS.n713 2.6005
R1305 VSS.n712 VSS.n711 2.6005
R1306 VSS.n711 VSS.n710 2.6005
R1307 VSS.n709 VSS.n708 2.6005
R1308 VSS.n708 VSS.n707 2.6005
R1309 VSS.n706 VSS.n705 2.6005
R1310 VSS.n705 VSS.n704 2.6005
R1311 VSS.n703 VSS.n702 2.6005
R1312 VSS.n702 VSS.n701 2.6005
R1313 VSS.n700 VSS.n699 2.6005
R1314 VSS.n699 VSS.n698 2.6005
R1315 VSS.n697 VSS.n696 2.6005
R1316 VSS.n696 VSS.n695 2.6005
R1317 VSS.n693 VSS.n692 2.6005
R1318 VSS.n692 VSS.n691 2.6005
R1319 VSS.n690 VSS.n689 2.6005
R1320 VSS.n689 VSS.n688 2.6005
R1321 VSS.n687 VSS.n686 2.6005
R1322 VSS.n686 VSS.n685 2.6005
R1323 VSS.n684 VSS.n683 2.6005
R1324 VSS.n683 VSS.n682 2.6005
R1325 VSS.n681 VSS.n680 2.6005
R1326 VSS.n680 VSS.n679 2.6005
R1327 VSS.n678 VSS.n677 2.6005
R1328 VSS.n677 VSS.n676 2.6005
R1329 VSS.n590 VSS.n589 2.6005
R1330 VSS.n589 VSS.n588 2.6005
R1331 VSS.n593 VSS.n592 2.6005
R1332 VSS.n592 VSS.n591 2.6005
R1333 VSS.n618 VSS.n617 2.6005
R1334 VSS.n614 VSS.n613 2.6005
R1335 VSS.n612 VSS.n611 2.6005
R1336 VSS.n608 VSS.n607 2.6005
R1337 VSS.n606 VSS.n605 2.6005
R1338 VSS.n603 VSS.n602 2.6005
R1339 VSS.n1100 VSS.n1099 2.6005
R1340 VSS.n624 VSS.n623 2.6005
R1341 VSS.n671 VSS.n670 2.6005
R1342 VSS.n670 VSS.n669 2.6005
R1343 VSS.n667 VSS.n666 2.6005
R1344 VSS.n666 VSS.n665 2.6005
R1345 VSS.n664 VSS.n663 2.6005
R1346 VSS.n663 VSS.n662 2.6005
R1347 VSS.n661 VSS.n660 2.6005
R1348 VSS.n660 VSS.n659 2.6005
R1349 VSS.n658 VSS.n657 2.6005
R1350 VSS.n657 VSS.n656 2.6005
R1351 VSS.n655 VSS.n654 2.6005
R1352 VSS.n654 VSS.n653 2.6005
R1353 VSS.n652 VSS.n651 2.6005
R1354 VSS.n651 VSS.n650 2.6005
R1355 VSS.n649 VSS.n648 2.6005
R1356 VSS.n648 VSS.n647 2.6005
R1357 VSS.n646 VSS.n645 2.6005
R1358 VSS.n645 VSS.n644 2.6005
R1359 VSS.n643 VSS.n642 2.6005
R1360 VSS.n642 VSS.n641 2.6005
R1361 VSS.n640 VSS.n639 2.6005
R1362 VSS.n639 VSS.n638 2.6005
R1363 VSS.n637 VSS.n636 2.6005
R1364 VSS.n636 VSS.n635 2.6005
R1365 VSS.n634 VSS.n633 2.6005
R1366 VSS.n633 VSS.n632 2.6005
R1367 VSS.n631 VSS.n630 2.6005
R1368 VSS.n630 VSS.n629 2.6005
R1369 VSS.n628 VSS.n627 2.6005
R1370 VSS.n627 VSS.n626 2.6005
R1371 VSS.n625 VSS.n624 2.6005
R1372 VSS.n622 VSS.n621 2.6005
R1373 VSS.n1054 VSS.n1053 2.6005
R1374 VSS.n1053 VSS.n1052 2.6005
R1375 VSS.n1058 VSS.n1057 2.6005
R1376 VSS.n1057 VSS.n1056 2.6005
R1377 VSS.n1061 VSS.n1060 2.6005
R1378 VSS.n1060 VSS.n1059 2.6005
R1379 VSS.n1065 VSS.n1064 2.6005
R1380 VSS.n1064 VSS.n1063 2.6005
R1381 VSS.n1068 VSS.n1067 2.6005
R1382 VSS.n1067 VSS.n1066 2.6005
R1383 VSS.n1072 VSS.n1071 2.6005
R1384 VSS.n1071 VSS.n1070 2.6005
R1385 VSS.n480 VSS.n467 2.6005
R1386 VSS.n467 VSS.n466 2.6005
R1387 VSS.n479 VSS.n478 2.6005
R1388 VSS.n478 VSS.n477 2.6005
R1389 VSS.n476 VSS.n475 2.6005
R1390 VSS.n475 VSS.n474 2.6005
R1391 VSS.n473 VSS.n472 2.6005
R1392 VSS.n472 VSS.n471 2.6005
R1393 VSS.n470 VSS.n469 2.6005
R1394 VSS.n469 VSS.n468 2.6005
R1395 VSS.n564 VSS.n563 2.6005
R1396 VSS.n563 VSS.n562 2.6005
R1397 VSS.n580 VSS.n579 2.6005
R1398 VSS.n520 VSS.n519 2.6005
R1399 VSS.n519 VSS.n518 2.6005
R1400 VSS.n516 VSS.n515 2.6005
R1401 VSS.n515 VSS.n514 2.6005
R1402 VSS.n513 VSS.n512 2.6005
R1403 VSS.n512 VSS.n511 2.6005
R1404 VSS.n509 VSS.n508 2.6005
R1405 VSS.n508 VSS.n507 2.6005
R1406 VSS.n506 VSS.n505 2.6005
R1407 VSS.n505 VSS.n504 2.6005
R1408 VSS.n581 VSS.n580 2.6005
R1409 VSS.n583 VSS.n582 2.6005
R1410 VSS.n566 VSS.n565 2.6005
R1411 VSS.n568 VSS.n567 2.6005
R1412 VSS.n570 VSS.n569 2.6005
R1413 VSS.n572 VSS.n571 2.6005
R1414 VSS.n574 VSS.n573 2.6005
R1415 VSS.n577 VSS.n576 2.6005
R1416 VSS.n1036 VSS.n1035 2.6005
R1417 VSS.n1029 VSS.n1028 2.6005
R1418 VSS.n1026 VSS.n1025 2.6005
R1419 VSS.n1023 VSS.n1022 2.6005
R1420 VSS.n1021 VSS.n1020 2.6005
R1421 VSS.n1019 VSS.n1018 2.6005
R1422 VSS.n1075 VSS.n1074 2.6005
R1423 VSS.n1074 VSS.n1073 2.6005
R1424 VSS.n1087 VSS.n1086 2.6005
R1425 VSS.n1086 VSS.n1085 2.6005
R1426 VSS.n1084 VSS.n1083 2.6005
R1427 VSS.n1083 VSS.n1082 2.6005
R1428 VSS.n1081 VSS.n1080 2.6005
R1429 VSS.n1080 VSS.n1079 2.6005
R1430 VSS.n746 VSS.n745 2.6005
R1431 VSS.n745 VSS.n744 2.6005
R1432 VSS.n674 VSS.n673 2.6005
R1433 VSS.n749 VSS.n748 2.6005
R1434 VSS.n748 VSS.n747 2.6005
R1435 VSS.n993 VSS.n992 2.6005
R1436 VSS.n992 VSS.n991 2.6005
R1437 VSS.n990 VSS.n989 2.6005
R1438 VSS.n989 VSS.n988 2.6005
R1439 VSS.n987 VSS.n986 2.6005
R1440 VSS.n986 VSS.n985 2.6005
R1441 VSS.n984 VSS.n983 2.6005
R1442 VSS.n983 VSS.n982 2.6005
R1443 VSS.n981 VSS.n980 2.6005
R1444 VSS.n980 VSS.n979 2.6005
R1445 VSS.n996 VSS.n995 2.6005
R1446 VSS.n995 VSS.n994 2.6005
R1447 VSS.n587 VSS.n586 2.6005
R1448 VSS.n1090 VSS.n1089 2.6005
R1449 VSS.n1089 VSS.n1088 2.6005
R1450 VSS.n1094 VSS.n1093 2.6005
R1451 VSS.n1093 VSS.n1092 2.6005
R1452 VSS.n1137 VSS.n1136 2.6005
R1453 VSS.n1097 VSS.n1096 2.6005
R1454 VSS.n1096 VSS.n1095 2.6005
R1455 VSS.n913 VSS.n912 2.6005
R1456 VSS.n912 VSS.n911 2.6005
R1457 VSS.n864 VSS.n863 2.6005
R1458 VSS.n863 VSS.n862 2.6005
R1459 VSS.n861 VSS.n860 2.6005
R1460 VSS.n860 VSS.n859 2.6005
R1461 VSS.n857 VSS.n856 2.6005
R1462 VSS.n856 VSS.n855 2.6005
R1463 VSS.n867 VSS.n866 2.6005
R1464 VSS.n866 VSS.n865 2.6005
R1465 VSS.n910 VSS.n909 2.6005
R1466 VSS.n909 VSS.n908 2.6005
R1467 VSS.n906 VSS.n905 2.6005
R1468 VSS.n904 VSS.n903 2.6005
R1469 VSS.n902 VSS.n901 2.6005
R1470 VSS.n900 VSS.n899 2.6005
R1471 VSS.n898 VSS.n897 2.6005
R1472 VSS.n896 VSS.n895 2.6005
R1473 VSS.n894 VSS.n893 2.6005
R1474 VSS.n892 VSS.n891 2.6005
R1475 VSS.n890 VSS.n889 2.6005
R1476 VSS.n888 VSS.n887 2.6005
R1477 VSS.n886 VSS.n885 2.6005
R1478 VSS.n884 VSS.n883 2.6005
R1479 VSS.n882 VSS.n881 2.6005
R1480 VSS.n880 VSS.n879 2.6005
R1481 VSS.n878 VSS.n877 2.6005
R1482 VSS.n876 VSS.n875 2.6005
R1483 VSS.n870 VSS.n869 2.6005
R1484 VSS.n73 VSS.n72 2.6005
R1485 VSS.n72 VSS.n71 2.6005
R1486 VSS.n70 VSS.n69 2.6005
R1487 VSS.n69 VSS.n68 2.6005
R1488 VSS.n67 VSS.n66 2.6005
R1489 VSS.n66 VSS.n65 2.6005
R1490 VSS.n64 VSS.n63 2.6005
R1491 VSS.n63 VSS.n62 2.6005
R1492 VSS.n61 VSS.n60 2.6005
R1493 VSS.n60 VSS.n59 2.6005
R1494 VSS.n58 VSS.n57 2.6005
R1495 VSS.n57 VSS.n56 2.6005
R1496 VSS.n55 VSS.n54 2.6005
R1497 VSS.n54 VSS.n53 2.6005
R1498 VSS.n52 VSS.n51 2.6005
R1499 VSS.n51 VSS.n50 2.6005
R1500 VSS.n49 VSS.n48 2.6005
R1501 VSS.n48 VSS.n47 2.6005
R1502 VSS.n46 VSS.n45 2.6005
R1503 VSS.n45 VSS.n44 2.6005
R1504 VSS.n43 VSS.n42 2.6005
R1505 VSS.n42 VSS.n41 2.6005
R1506 VSS.n40 VSS.n39 2.6005
R1507 VSS.n39 VSS.n38 2.6005
R1508 VSS.n37 VSS.n36 2.6005
R1509 VSS.n36 VSS.n35 2.6005
R1510 VSS.n34 VSS.n33 2.6005
R1511 VSS.n33 VSS.n32 2.6005
R1512 VSS.n31 VSS.n30 2.6005
R1513 VSS.n30 VSS.n29 2.6005
R1514 VSS.n28 VSS.n27 2.6005
R1515 VSS.n27 VSS.n26 2.6005
R1516 VSS.n25 VSS.n24 2.6005
R1517 VSS.n19 VSS.n18 2.6005
R1518 VSS.n18 VSS.n17 2.6005
R1519 VSS.n16 VSS.n15 2.6005
R1520 VSS.n15 VSS.n14 2.6005
R1521 VSS.n13 VSS.n12 2.6005
R1522 VSS.n12 VSS.n11 2.6005
R1523 VSS.n10 VSS.n9 2.6005
R1524 VSS.n9 VSS.n8 2.6005
R1525 VSS.n7 VSS.n6 2.6005
R1526 VSS.n6 VSS.n5 2.6005
R1527 VSS.n773 VSS.n772 2.6005
R1528 VSS.n772 VSS.n771 2.6005
R1529 VSS.n776 VSS.n775 2.6005
R1530 VSS.n775 VSS.n774 2.6005
R1531 VSS.n22 VSS.n21 2.6005
R1532 VSS.n21 VSS.n20 2.6005
R1533 VSS.n801 VSS.n800 2.6005
R1534 VSS.n797 VSS.n796 2.6005
R1535 VSS.n795 VSS.n794 2.6005
R1536 VSS.n791 VSS.n790 2.6005
R1537 VSS.n789 VSS.n788 2.6005
R1538 VSS.n786 VSS.n785 2.6005
R1539 VSS.n873 VSS.n872 2.6005
R1540 VSS.n853 VSS.n852 2.6005
R1541 VSS.n852 VSS.n851 2.6005
R1542 VSS.n850 VSS.n849 2.6005
R1543 VSS.n849 VSS.n848 2.6005
R1544 VSS.n847 VSS.n846 2.6005
R1545 VSS.n846 VSS.n845 2.6005
R1546 VSS.n844 VSS.n843 2.6005
R1547 VSS.n843 VSS.n842 2.6005
R1548 VSS.n841 VSS.n840 2.6005
R1549 VSS.n840 VSS.n839 2.6005
R1550 VSS.n838 VSS.n837 2.6005
R1551 VSS.n837 VSS.n836 2.6005
R1552 VSS.n835 VSS.n834 2.6005
R1553 VSS.n834 VSS.n833 2.6005
R1554 VSS.n832 VSS.n831 2.6005
R1555 VSS.n831 VSS.n830 2.6005
R1556 VSS.n829 VSS.n828 2.6005
R1557 VSS.n828 VSS.n827 2.6005
R1558 VSS.n826 VSS.n825 2.6005
R1559 VSS.n825 VSS.n824 2.6005
R1560 VSS.n823 VSS.n822 2.6005
R1561 VSS.n822 VSS.n821 2.6005
R1562 VSS.n820 VSS.n819 2.6005
R1563 VSS.n819 VSS.n818 2.6005
R1564 VSS.n817 VSS.n816 2.6005
R1565 VSS.n816 VSS.n815 2.6005
R1566 VSS.n814 VSS.n813 2.6005
R1567 VSS.n813 VSS.n812 2.6005
R1568 VSS.n811 VSS.n810 2.6005
R1569 VSS.n810 VSS.n809 2.6005
R1570 VSS.n808 VSS.n807 2.6005
R1571 VSS.n807 VSS.n806 2.6005
R1572 VSS.n805 VSS.n804 2.6005
R1573 VSS.n770 VSS.n769 2.6005
R1574 VSS.n83 VSS.n82 2.6005
R1575 VSS.n82 VSS.n81 2.6005
R1576 VSS.n1620 VSS.n1619 2.6005
R1577 VSS.n1619 VSS.n1618 2.6005
R1578 VSS.n1616 VSS.n1615 2.6005
R1579 VSS.n1615 VSS.n1614 2.6005
R1580 VSS.n1613 VSS.n1612 2.6005
R1581 VSS.n1612 VSS.n1611 2.6005
R1582 VSS.n1610 VSS.n1609 2.6005
R1583 VSS.n1609 VSS.n1608 2.6005
R1584 VSS.n1623 VSS.n1622 2.6005
R1585 VSS.n1622 VSS.n1621 2.6005
R1586 VSS.n80 VSS.n79 2.6005
R1587 VSS.n79 VSS.n78 2.6005
R1588 VSS.n77 VSS.n76 2.6005
R1589 VSS.n76 VSS.n75 2.6005
R1590 VSS.n86 VSS.n85 2.6005
R1591 VSS.n1590 VSS.n1589 2.6005
R1592 VSS.n1589 VSS.n1588 2.6005
R1593 VSS.n1587 VSS.n1586 2.6005
R1594 VSS.n1586 VSS.n1585 2.6005
R1595 VSS.n1584 VSS.n1583 2.6005
R1596 VSS.n1583 VSS.n1582 2.6005
R1597 VSS.n1581 VSS.n1580 2.6005
R1598 VSS.n1580 VSS.n1579 2.6005
R1599 VSS.n1578 VSS.n1577 2.6005
R1600 VSS.n1577 VSS.n1576 2.6005
R1601 VSS.n1575 VSS.n1574 2.6005
R1602 VSS.n1574 VSS.n1573 2.6005
R1603 VSS.n1593 VSS.n1592 2.6005
R1604 VSS.n1592 VSS.n1591 2.6005
R1605 VSS.n89 VSS.n88 2.6005
R1606 VSS.n1596 VSS.n1595 2.6005
R1607 VSS.n1598 VSS.n1597 2.6005
R1608 VSS.n1602 VSS.n1601 2.6005
R1609 VSS.n1604 VSS.n1603 2.6005
R1610 VSS.n1511 VSS.n1510 2.6005
R1611 VSS.n1509 VSS.n1508 2.6005
R1612 VSS.n161 VSS.n160 2.6005
R1613 VSS.n160 VSS.n159 2.6005
R1614 VSS.n158 VSS.n157 2.6005
R1615 VSS.n157 VSS.n156 2.6005
R1616 VSS.n155 VSS.n154 2.6005
R1617 VSS.n154 VSS.n153 2.6005
R1618 VSS.n152 VSS.n151 2.6005
R1619 VSS.n151 VSS.n150 2.6005
R1620 VSS.n149 VSS.n148 2.6005
R1621 VSS.n148 VSS.n147 2.6005
R1622 VSS.n146 VSS.n145 2.6005
R1623 VSS.n145 VSS.n144 2.6005
R1624 VSS.n143 VSS.n142 2.6005
R1625 VSS.n142 VSS.n141 2.6005
R1626 VSS.n140 VSS.n139 2.6005
R1627 VSS.n139 VSS.n138 2.6005
R1628 VSS.n1350 VSS.n1349 2.6005
R1629 VSS.n1356 VSS.n1355 2.6005
R1630 VSS.n1352 VSS.n1351 2.6005
R1631 VSS.n1549 VSS.n1548 2.6005
R1632 VSS.n1551 VSS.n1550 2.6005
R1633 VSS.n1557 VSS.n1556 2.6005
R1634 VSS.n1556 VSS.n1555 2.6005
R1635 VSS.n1561 VSS.n1560 2.6005
R1636 VSS.n1560 VSS.n1559 2.6005
R1637 VSS.n1564 VSS.n1563 2.6005
R1638 VSS.n1563 VSS.n1562 2.6005
R1639 VSS.n1567 VSS.n1566 2.6005
R1640 VSS.n1566 VSS.n1565 2.6005
R1641 VSS.n1571 VSS.n1570 2.6005
R1642 VSS.n1570 VSS.n1569 2.6005
R1643 VSS.n1554 VSS.n1553 2.6005
R1644 VSS.n114 VSS.n113 2.6005
R1645 VSS.n116 VSS.n115 2.6005
R1646 VSS.n137 VSS.n136 2.6005
R1647 VSS.n136 VSS.n135 2.6005
R1648 VSS.n133 VSS.n132 2.6005
R1649 VSS.n132 VSS.n131 2.6005
R1650 VSS.n130 VSS.n129 2.6005
R1651 VSS.n129 VSS.n128 2.6005
R1652 VSS.n127 VSS.n126 2.6005
R1653 VSS.n126 VSS.n125 2.6005
R1654 VSS.n123 VSS.n122 2.6005
R1655 VSS.n122 VSS.n121 2.6005
R1656 VSS.n119 VSS.n118 2.6005
R1657 VSS.n1330 VSS.n1329 2.6005
R1658 VSS.n1329 VSS.n1328 2.6005
R1659 VSS.n1347 VSS.n1346 2.6005
R1660 VSS.n1346 VSS.n1345 2.6005
R1661 VSS.n1343 VSS.n1342 2.6005
R1662 VSS.n1342 VSS.n1341 2.6005
R1663 VSS.n1340 VSS.n1339 2.6005
R1664 VSS.n1339 VSS.n1338 2.6005
R1665 VSS.n1337 VSS.n1336 2.6005
R1666 VSS.n1336 VSS.n1335 2.6005
R1667 VSS.n1334 VSS.n1333 2.6005
R1668 VSS.n1333 VSS.n1332 2.6005
R1669 VSS.n1533 VSS.n1532 2.6005
R1670 VSS.n1532 VSS.n1531 2.6005
R1671 VSS.n1536 VSS.n1535 2.6005
R1672 VSS.n1535 VSS.n1534 2.6005
R1673 VSS.n1539 VSS.n1538 2.6005
R1674 VSS.n1538 VSS.n1537 2.6005
R1675 VSS.n1542 VSS.n1541 2.6005
R1676 VSS.n1541 VSS.n1540 2.6005
R1677 VSS.n1545 VSS.n1544 2.6005
R1678 VSS.n1544 VSS.n1543 2.6005
R1679 VSS.n99 VSS.n98 2.6005
R1680 VSS.n98 VSS.n97 2.6005
R1681 VSS.n102 VSS.n101 2.6005
R1682 VSS.n101 VSS.n100 2.6005
R1683 VSS.n105 VSS.n104 2.6005
R1684 VSS.n104 VSS.n103 2.6005
R1685 VSS.n110 VSS.n109 2.6005
R1686 VSS.n109 VSS.n108 2.6005
R1687 VSS.n95 VSS.n94 2.6005
R1688 VSS.n94 VSS.n93 2.6005
R1689 VSS.n1529 VSS.n1528 2.6005
R1690 VSS.n1526 VSS.n1525 2.6005
R1691 VSS.n1515 VSS.n1514 2.6005
R1692 VSS.n1517 VSS.n1516 2.6005
R1693 VSS.n1520 VSS.n1519 2.6005
R1694 VSS.n1522 VSS.n1521 2.6005
R1695 VSS.n1686 VSS.n1685 2.6005
R1696 VSS.n1685 VSS.n1684 2.6005
R1697 VSS.n1683 VSS.n1682 2.6005
R1698 VSS.n1682 VSS.n1681 2.6005
R1699 VSS.n1676 VSS.n1675 2.6005
R1700 VSS.n1680 VSS.n1679 2.6005
R1701 VSS.n1695 VSS.n1694 2.6005
R1702 VSS.n1694 VSS.n1693 2.6005
R1703 VSS.n1692 VSS.n1691 2.6005
R1704 VSS.n1691 VSS.n1690 2.6005
R1705 VSS.n1689 VSS.n1688 2.6005
R1706 VSS.n1688 VSS.n1687 2.6005
R1707 VSS.n1700 VSS.n1699 2.6005
R1708 VSS.n1699 VSS.n1698 2.6005
R1709 VSS.n1658 VSS.n1657 2.6005
R1710 VSS.n1657 VSS.n1656 2.6005
R1711 VSS.n1655 VSS.n1654 2.6005
R1712 VSS.n1654 VSS.n1653 2.6005
R1713 VSS.n1652 VSS.n1651 2.6005
R1714 VSS.n1651 VSS.n1650 2.6005
R1715 VSS.n1649 VSS.n1648 2.6005
R1716 VSS.n1648 VSS.n1647 2.6005
R1717 VSS.n1713 VSS.n1712 2.6005
R1718 VSS.n1712 VSS.n1711 2.6005
R1719 VSS.n1719 VSS.n1718 2.6005
R1720 VSS.n1718 VSS.n1717 2.6005
R1721 VSS.n1722 VSS.n1721 2.6005
R1722 VSS.n1721 VSS.n1720 2.6005
R1723 VSS.n1725 VSS.n1724 2.6005
R1724 VSS.n1724 VSS.n1723 2.6005
R1725 VSS.n1728 VSS.n1727 2.6005
R1726 VSS.n1727 VSS.n1726 2.6005
R1727 VSS.n1716 VSS.n1715 2.6005
R1728 VSS.n1715 VSS.n1714 2.6005
R1729 VSS.n1730 VSS.n1729 2.6005
R1730 VSS.n168 VSS.n167 2.6005
R1731 VSS.n164 VSS.n163 2.6005
R1732 VSS.n1 VSS.n0 2.6005
R1733 VSS.n1738 VSS.n1737 2.6005
R1734 VSS.n1735 VSS.n1734 2.6005
R1735 VSS.n185 VSS.n184 2.6005
R1736 VSS.n184 VSS.n183 2.6005
R1737 VSS.n182 VSS.n181 2.6005
R1738 VSS.n181 VSS.n180 2.6005
R1739 VSS.n179 VSS.n178 2.6005
R1740 VSS.n178 VSS.n177 2.6005
R1741 VSS.n176 VSS.n175 2.6005
R1742 VSS.n175 VSS.n174 2.6005
R1743 VSS.n173 VSS.n172 2.6005
R1744 VSS.n172 VSS.n171 2.6005
R1745 VSS.n170 VSS.n169 2.6005
R1746 VSS.n195 VSS.n194 2.6005
R1747 VSS.n190 VSS.n189 2.6005
R1748 VSS.n188 VSS.n187 2.6005
R1749 VSS.n187 VSS.n186 2.6005
R1750 VSS.n1703 VSS.n1702 2.6005
R1751 VSS.n1702 VSS.n1701 2.6005
R1752 VSS.n1706 VSS.n1705 2.6005
R1753 VSS.n1705 VSS.n1704 2.6005
R1754 VSS.n1709 VSS.n1708 2.6005
R1755 VSS.n1708 VSS.n1707 2.6005
R1756 VSS.n220 VSS.n219 2.6005
R1757 VSS.n219 VSS.n218 2.6005
R1758 VSS.n223 VSS.n222 2.6005
R1759 VSS.n222 VSS.n221 2.6005
R1760 VSS.n226 VSS.n225 2.6005
R1761 VSS.n225 VSS.n224 2.6005
R1762 VSS.n229 VSS.n228 2.6005
R1763 VSS.n228 VSS.n227 2.6005
R1764 VSS.n232 VSS.n231 2.6005
R1765 VSS.n231 VSS.n230 2.6005
R1766 VSS.n235 VSS.n234 2.6005
R1767 VSS.n234 VSS.n233 2.6005
R1768 VSS.n238 VSS.n237 2.6005
R1769 VSS.n237 VSS.n236 2.6005
R1770 VSS.n241 VSS.n240 2.6005
R1771 VSS.n240 VSS.n239 2.6005
R1772 VSS.n244 VSS.n243 2.6005
R1773 VSS.n243 VSS.n242 2.6005
R1774 VSS.n247 VSS.n246 2.6005
R1775 VSS.n246 VSS.n245 2.6005
R1776 VSS.n250 VSS.n249 2.6005
R1777 VSS.n249 VSS.n248 2.6005
R1778 VSS.n253 VSS.n252 2.6005
R1779 VSS.n252 VSS.n251 2.6005
R1780 VSS.n256 VSS.n255 2.6005
R1781 VSS.n255 VSS.n254 2.6005
R1782 VSS.n259 VSS.n258 2.6005
R1783 VSS.n258 VSS.n257 2.6005
R1784 VSS.n262 VSS.n261 2.6005
R1785 VSS.n261 VSS.n260 2.6005
R1786 VSS.n265 VSS.n264 2.6005
R1787 VSS.n264 VSS.n263 2.6005
R1788 VSS.n1442 VSS.n1441 2.6005
R1789 VSS.n1441 VSS.n1440 2.6005
R1790 VSS.n198 VSS.n197 2.6005
R1791 VSS.n197 VSS.n196 2.6005
R1792 VSS.n201 VSS.n200 2.6005
R1793 VSS.n200 VSS.n199 2.6005
R1794 VSS.n204 VSS.n203 2.6005
R1795 VSS.n203 VSS.n202 2.6005
R1796 VSS.n207 VSS.n206 2.6005
R1797 VSS.n206 VSS.n205 2.6005
R1798 VSS.n210 VSS.n209 2.6005
R1799 VSS.n209 VSS.n208 2.6005
R1800 VSS.n213 VSS.n212 2.6005
R1801 VSS.n212 VSS.n211 2.6005
R1802 VSS.n1445 VSS.n1444 2.6005
R1803 VSS.n1444 VSS.n1443 2.6005
R1804 VSS.n1449 VSS.n1448 2.6005
R1805 VSS.n1448 VSS.n1447 2.6005
R1806 VSS.n1452 VSS.n1451 2.6005
R1807 VSS.n1451 VSS.n1450 2.6005
R1808 VSS.n1455 VSS.n1454 2.6005
R1809 VSS.n1454 VSS.n1453 2.6005
R1810 VSS.n1458 VSS.n1457 2.6005
R1811 VSS.n1457 VSS.n1456 2.6005
R1812 VSS.n1461 VSS.n1460 2.6005
R1813 VSS.n1460 VSS.n1459 2.6005
R1814 VSS.n1464 VSS.n1463 2.6005
R1815 VSS.n1463 VSS.n1462 2.6005
R1816 VSS.n1467 VSS.n1466 2.6005
R1817 VSS.n1466 VSS.n1465 2.6005
R1818 VSS.n1470 VSS.n1469 2.6005
R1819 VSS.n1469 VSS.n1468 2.6005
R1820 VSS.n1473 VSS.n1472 2.6005
R1821 VSS.n1472 VSS.n1471 2.6005
R1822 VSS.n1476 VSS.n1475 2.6005
R1823 VSS.n1475 VSS.n1474 2.6005
R1824 VSS.n1479 VSS.n1478 2.6005
R1825 VSS.n1478 VSS.n1477 2.6005
R1826 VSS.n1482 VSS.n1481 2.6005
R1827 VSS.n1481 VSS.n1480 2.6005
R1828 VSS.n1485 VSS.n1484 2.6005
R1829 VSS.n1484 VSS.n1483 2.6005
R1830 VSS.n1488 VSS.n1487 2.6005
R1831 VSS.n1487 VSS.n1486 2.6005
R1832 VSS.n1491 VSS.n1490 2.6005
R1833 VSS.n1490 VSS.n1489 2.6005
R1834 VSS.n1495 VSS.n1494 2.6005
R1835 VSS.n1494 VSS.n1493 2.6005
R1836 VSS.n1437 VSS.n1436 2.6005
R1837 VSS.n1432 VSS.n1431 2.6005
R1838 VSS.n1430 VSS.n1429 2.6005
R1839 VSS.n1427 VSS.n1426 2.6005
R1840 VSS.n1425 VSS.n1424 2.6005
R1841 VSS.n1422 VSS.n1421 2.6005
R1842 VSS.n1366 VSS.n1365 2.6005
R1843 VSS.n1368 VSS.n1367 2.6005
R1844 VSS.n1370 VSS.n1369 2.6005
R1845 VSS.n1372 VSS.n1371 2.6005
R1846 VSS.n1374 VSS.n1373 2.6005
R1847 VSS.n1376 VSS.n1375 2.6005
R1848 VSS.n1378 VSS.n1377 2.6005
R1849 VSS.n1380 VSS.n1379 2.6005
R1850 VSS.n1382 VSS.n1381 2.6005
R1851 VSS.n1384 VSS.n1383 2.6005
R1852 VSS.n1386 VSS.n1385 2.6005
R1853 VSS.n1388 VSS.n1387 2.6005
R1854 VSS.n1390 VSS.n1389 2.6005
R1855 VSS.n1392 VSS.n1391 2.6005
R1856 VSS.n1394 VSS.n1393 2.6005
R1857 VSS.n1396 VSS.n1395 2.6005
R1858 VSS.n1363 VSS.n1362 2.6005
R1859 VSS.n1417 VSS.n1416 2.6005
R1860 VSS.n1416 VSS.n1415 2.6005
R1861 VSS.n1413 VSS.n1412 2.6005
R1862 VSS.n1412 VSS.n1411 2.6005
R1863 VSS.n1409 VSS.n1408 2.6005
R1864 VSS.n1408 VSS.n1407 2.6005
R1865 VSS.n1359 VSS.n1358 2.6005
R1866 VSS.n1358 VSS.n1357 2.6005
R1867 VSS.n1241 VSS.n1240 2.6005
R1868 VSS.n1240 VSS.n1239 2.6005
R1869 VSS.n1405 VSS.n1404 2.6005
R1870 VSS.n1404 VSS.n1403 2.6005
R1871 VSS.n1420 VSS.n1419 2.6005
R1872 VSS.n1419 VSS.n1418 2.6005
R1873 VSS.n1499 VSS.n1498 2.6005
R1874 VSS.n1498 VSS.n1497 2.6005
R1875 VSS.n1503 VSS.n1502 2.6005
R1876 VSS.n1502 VSS.n1501 2.6005
R1877 VSS.n291 VSS.n290 2.6005
R1878 VSS.n290 VSS.n289 2.6005
R1879 VSS.n288 VSS.n287 2.6005
R1880 VSS.n287 VSS.n286 2.6005
R1881 VSS.n285 VSS.n284 2.6005
R1882 VSS.n284 VSS.n283 2.6005
R1883 VSS.n282 VSS.n281 2.6005
R1884 VSS.n281 VSS.n280 2.6005
R1885 VSS.n278 VSS.n277 2.6005
R1886 VSS.n277 VSS.n276 2.6005
R1887 VSS.n268 VSS.n267 2.6005
R1888 VSS.n271 VSS.n270 2.6005
R1889 VSS.n270 VSS.n269 2.6005
R1890 VSS.n274 VSS.n273 2.6005
R1891 VSS.n273 VSS.n272 2.6005
R1892 VSS.n1238 VSS.n1237 2.6005
R1893 VSS.n1237 VSS.n1236 2.6005
R1894 VSS.n1235 VSS.n1234 2.6005
R1895 VSS.n1234 VSS.n1233 2.6005
R1896 VSS.n1232 VSS.n1231 2.6005
R1897 VSS.n1231 VSS.n1230 2.6005
R1898 VSS.n1229 VSS.n1228 2.6005
R1899 VSS.n1228 VSS.n1227 2.6005
R1900 VSS.n1226 VSS.n1225 2.6005
R1901 VSS.n1225 VSS.n1224 2.6005
R1902 VSS.n1223 VSS.n1222 2.6005
R1903 VSS.n1222 VSS.n1221 2.6005
R1904 VSS.n1220 VSS.n1219 2.6005
R1905 VSS.n1219 VSS.n1218 2.6005
R1906 VSS.n1217 VSS.n1216 2.6005
R1907 VSS.n1216 VSS.n1215 2.6005
R1908 VSS.n1214 VSS.n1213 2.6005
R1909 VSS.n1213 VSS.n1212 2.6005
R1910 VSS.n1402 VSS.n1401 2.6005
R1911 VSS.n1401 VSS.n1400 2.6005
R1912 VSS.n1399 VSS.n1398 2.6005
R1913 VSS.n1398 VSS.n1397 2.6005
R1914 VSS.n498 VSS.n497 2.6005
R1915 VSS.n491 VSS.n490 2.6005
R1916 VSS.n488 VSS.n487 2.6005
R1917 VSS.n486 VSS.n485 2.6005
R1918 VSS.n483 VSS.n482 2.6005
R1919 VSS.n482 VSS.n481 2.6005
R1920 VSS.n500 VSS.n499 2.6005
R1921 VSS.n523 VSS.n522 2.6005
R1922 VSS.n522 VSS.n521 2.6005
R1923 VSS.n998 VSS.n997 2.6005
R1924 VSS.n1041 VSS.n1040 2.6005
R1925 VSS.n1043 VSS.n1042 2.6005
R1926 VSS.n1045 VSS.n1044 2.6005
R1927 VSS.n1047 VSS.n1046 2.6005
R1928 VSS.n1049 VSS.n1048 2.6005
R1929 VSS.n1051 VSS.n1050 2.6005
R1930 VSS.n1254 VSS.n1253 2.6005
R1931 VSS.n1250 VSS.n1249 2.6005
R1932 VSS.n1248 VSS.n1247 2.6005
R1933 VSS.n1001 VSS.n1000 2.6005
R1934 VSS.n1000 VSS.n999 2.6005
R1935 VSS.n1004 VSS.n1003 2.6005
R1936 VSS.n1003 VSS.n1002 2.6005
R1937 VSS.n1007 VSS.n1006 2.6005
R1938 VSS.n1006 VSS.n1005 2.6005
R1939 VSS.n1010 VSS.n1009 2.6005
R1940 VSS.n1009 VSS.n1008 2.6005
R1941 VSS.n1013 VSS.n1012 2.6005
R1942 VSS.n1012 VSS.n1011 2.6005
R1943 VSS.n1016 VSS.n1015 2.6005
R1944 VSS.n1015 VSS.n1014 2.6005
R1945 VSS.n1273 VSS.n1272 2.6005
R1946 VSS.n1272 VSS.n1271 2.6005
R1947 VSS.n1270 VSS.n1269 2.6005
R1948 VSS.n1269 VSS.n1268 2.6005
R1949 VSS.n1267 VSS.n1266 2.6005
R1950 VSS.n1266 VSS.n1265 2.6005
R1951 VSS.n1264 VSS.n1263 2.6005
R1952 VSS.n1263 VSS.n1262 2.6005
R1953 VSS.n1261 VSS.n1260 2.6005
R1954 VSS.n1260 VSS.n1259 2.6005
R1955 VSS.n1258 VSS.n1257 2.6005
R1956 VSS.n1257 VSS.n1256 2.6005
R1957 VSS.n1276 VSS.n1275 2.6005
R1958 VSS.n1275 VSS.n1274 2.6005
R1959 VSS.n1316 VSS.n1278 2.6005
R1960 VSS.n1278 VSS.n1277 2.6005
R1961 VSS.n1293 VSS.n1292 2.6005
R1962 VSS.n1297 VSS.n1296 2.6005
R1963 VSS.n1300 VSS.n1299 2.6005
R1964 VSS.n1299 VSS.n1298 2.6005
R1965 VSS.n1303 VSS.n1302 2.6005
R1966 VSS.n1302 VSS.n1301 2.6005
R1967 VSS.n1306 VSS.n1305 2.6005
R1968 VSS.n1305 VSS.n1304 2.6005
R1969 VSS.n1309 VSS.n1308 2.6005
R1970 VSS.n1308 VSS.n1307 2.6005
R1971 VSS.n1312 VSS.n1311 2.6005
R1972 VSS.n1311 VSS.n1310 2.6005
R1973 VSS.n1315 VSS.n1314 2.6005
R1974 VSS.n1314 VSS.n1313 2.6005
R1975 VSS.n1291 VSS.n1290 2.6005
R1976 VSS.n918 VSS.n917 2.6005
R1977 VSS.n917 VSS.n916 2.6005
R1978 VSS.n1325 VSS.n1324 2.6005
R1979 VSS.n1324 VSS.n1323 2.6005
R1980 VSS.n1322 VSS.n1321 2.6005
R1981 VSS.n1321 VSS.n1320 2.6005
R1982 VSS.n1319 VSS.n1318 2.6005
R1983 VSS.n1318 VSS.n1317 2.6005
R1984 VSS.n752 VSS.n751 2.6005
R1985 VSS.n751 VSS.n750 2.6005
R1986 VSS.n755 VSS.n754 2.6005
R1987 VSS.n754 VSS.n753 2.6005
R1988 VSS.n759 VSS.n758 2.6005
R1989 VSS.n758 VSS.n757 2.6005
R1990 VSS.n761 VSS.n760 2.6005
R1991 VSS.n765 VSS.n764 2.6005
R1992 VSS.n767 VSS.n766 2.6005
R1993 VSS.n925 VSS.n924 2.6005
R1994 VSS.n924 VSS.n923 2.6005
R1995 VSS.n928 VSS.n927 2.6005
R1996 VSS.n927 VSS.n926 2.6005
R1997 VSS.n931 VSS.n930 2.6005
R1998 VSS.n930 VSS.n929 2.6005
R1999 VSS.n934 VSS.n933 2.6005
R2000 VSS.n933 VSS.n932 2.6005
R2001 VSS.n937 VSS.n936 2.6005
R2002 VSS.n936 VSS.n935 2.6005
R2003 VSS.n940 VSS.n939 2.6005
R2004 VSS.n939 VSS.n938 2.6005
R2005 VSS.n943 VSS.n942 2.6005
R2006 VSS.n942 VSS.n941 2.6005
R2007 VSS.n946 VSS.n945 2.6005
R2008 VSS.n945 VSS.n944 2.6005
R2009 VSS.n949 VSS.n948 2.6005
R2010 VSS.n948 VSS.n947 2.6005
R2011 VSS.n922 VSS.n921 2.6005
R2012 VSS.n921 VSS.n920 2.6005
R2013 VSS.n1288 VSS.n1279 2.6005
R2014 VSS.n1211 VSS.n1178 2.6005
R2015 VSS.n1178 VSS.n1177 2.6005
R2016 VSS.n1210 VSS.n1209 2.6005
R2017 VSS.n1209 VSS.n1208 2.6005
R2018 VSS.n1205 VSS.n1204 2.6005
R2019 VSS.n1204 VSS.n1203 2.6005
R2020 VSS.n1202 VSS.n1201 2.6005
R2021 VSS.n1201 VSS.n1200 2.6005
R2022 VSS.n1199 VSS.n1198 2.6005
R2023 VSS.n1198 VSS.n1197 2.6005
R2024 VSS.n1195 VSS.n1194 2.6005
R2025 VSS.n1194 VSS.n1193 2.6005
R2026 VSS.n1192 VSS.n1191 2.6005
R2027 VSS.n1191 VSS.n1190 2.6005
R2028 VSS.n1188 VSS.n1187 2.6005
R2029 VSS.n1187 VSS.n1186 2.6005
R2030 VSS.n1184 VSS.n1183 2.6005
R2031 VSS.n1183 VSS.n1182 2.6005
R2032 VSS.n1244 VSS.n1243 2.6005
R2033 VSS.n1243 VSS.n1242 2.6005
R2034 VSS.n1287 VSS.n1286 2.6005
R2035 VSS.n1286 VSS.n1285 2.6005
R2036 VSS.n1283 VSS.n1282 2.6005
R2037 VSS.n1282 VSS.n1281 2.6005
R2038 VSS.n955 VSS.n954 2.6005
R2039 VSS.n954 VSS.n953 2.6005
R2040 VSS.n958 VSS.n957 2.6005
R2041 VSS.n957 VSS.n956 2.6005
R2042 VSS.n962 VSS.n961 2.6005
R2043 VSS.n961 VSS.n960 2.6005
R2044 VSS.n965 VSS.n964 2.6005
R2045 VSS.n964 VSS.n963 2.6005
R2046 VSS.n968 VSS.n967 2.6005
R2047 VSS.n967 VSS.n966 2.6005
R2048 VSS.n973 VSS.n972 2.6005
R2049 VSS.n972 VSS.n971 2.6005
R2050 VSS.n976 VSS.n975 2.6005
R2051 VSS.n975 VSS.n974 2.6005
R2052 VSS.n1175 VSS.n378 2.6005
R2053 VSS.n378 VSS.n377 2.6005
R2054 VSS.n1162 VSS.n1161 2.6005
R2055 VSS.n1161 VSS.n1160 2.6005
R2056 VSS.n1165 VSS.n1164 2.6005
R2057 VSS.n1164 VSS.n1163 2.6005
R2058 VSS.n1168 VSS.n1167 2.6005
R2059 VSS.n1167 VSS.n1166 2.6005
R2060 VSS.n1171 VSS.n1170 2.6005
R2061 VSS.n1170 VSS.n1169 2.6005
R2062 VSS.n1174 VSS.n1173 2.6005
R2063 VSS.n1173 VSS.n1172 2.6005
R2064 VSS.n373 VSS.n372 2.6005
R2065 VSS.n372 VSS.n371 2.6005
R2066 VSS.n376 VSS.n375 2.6005
R2067 VSS.n375 VSS.n374 2.6005
R2068 VSS.n370 VSS.n369 2.6005
R2069 VSS.n369 VSS.n368 2.6005
R2070 VSS.n323 VSS.n322 2.6005
R2071 VSS.n322 VSS.n321 2.6005
R2072 VSS.n326 VSS.n325 2.6005
R2073 VSS.n325 VSS.n324 2.6005
R2074 VSS.n329 VSS.n328 2.6005
R2075 VSS.n328 VSS.n327 2.6005
R2076 VSS.n332 VSS.n331 2.6005
R2077 VSS.n331 VSS.n330 2.6005
R2078 VSS.n335 VSS.n334 2.6005
R2079 VSS.n334 VSS.n333 2.6005
R2080 VSS.n338 VSS.n337 2.6005
R2081 VSS.n337 VSS.n336 2.6005
R2082 VSS.n340 VSS.n339 2.6005
R2083 VSS.n339 VSS.t38 2.6005
R2084 VSS.n343 VSS.n342 2.6005
R2085 VSS.n342 VSS.n341 2.6005
R2086 VSS.n346 VSS.n345 2.6005
R2087 VSS.n345 VSS.n344 2.6005
R2088 VSS.n349 VSS.n348 2.6005
R2089 VSS.n348 VSS.n347 2.6005
R2090 VSS.n352 VSS.n351 2.6005
R2091 VSS.n351 VSS.n350 2.6005
R2092 VSS.n355 VSS.n354 2.6005
R2093 VSS.n354 VSS.n353 2.6005
R2094 VSS.n358 VSS.n357 2.6005
R2095 VSS.n357 VSS.n356 2.6005
R2096 VSS.n361 VSS.n360 2.6005
R2097 VSS.n360 VSS.n359 2.6005
R2098 VSS.n364 VSS.n363 2.6005
R2099 VSS.n363 VSS.n362 2.6005
R2100 VSS.n367 VSS.n366 2.6005
R2101 VSS.n366 VSS.n365 2.6005
R2102 VSS.n381 VSS.n380 2.6005
R2103 VSS.n380 VSS.n379 2.6005
R2104 VSS.n304 VSS.n303 2.6005
R2105 VSS.n303 VSS.n302 2.6005
R2106 VSS.n307 VSS.n306 2.6005
R2107 VSS.n306 VSS.n305 2.6005
R2108 VSS.n310 VSS.n309 2.6005
R2109 VSS.n309 VSS.n308 2.6005
R2110 VSS.n313 VSS.n312 2.6005
R2111 VSS.n312 VSS.n311 2.6005
R2112 VSS.n316 VSS.n315 2.6005
R2113 VSS.n315 VSS.n314 2.6005
R2114 VSS.n319 VSS.n318 2.6005
R2115 VSS.n318 VSS.n317 2.6005
R2116 VSS.n384 VSS.n383 2.6005
R2117 VSS.n383 VSS.n382 2.6005
R2118 VSS.n401 VSS.n400 2.6005
R2119 VSS.n396 VSS.n395 2.6005
R2120 VSS.n394 VSS.n393 2.6005
R2121 VSS.n391 VSS.n390 2.6005
R2122 VSS.n389 VSS.n388 2.6005
R2123 VSS.n386 VSS.n385 2.6005
R2124 VSS.n407 VSS.n406 2.6005
R2125 VSS.n406 VSS.n405 2.6005
R2126 VSS.n410 VSS.n409 2.6005
R2127 VSS.n409 VSS.n408 2.6005
R2128 VSS.n413 VSS.n412 2.6005
R2129 VSS.n412 VSS.n411 2.6005
R2130 VSS.n416 VSS.n415 2.6005
R2131 VSS.n415 VSS.n414 2.6005
R2132 VSS.n419 VSS.n418 2.6005
R2133 VSS.n418 VSS.n417 2.6005
R2134 VSS.n422 VSS.n421 2.6005
R2135 VSS.n421 VSS.n420 2.6005
R2136 VSS.n425 VSS.n424 2.6005
R2137 VSS.n424 VSS.n423 2.6005
R2138 VSS.n428 VSS.n427 2.6005
R2139 VSS.n427 VSS.n426 2.6005
R2140 VSS.n431 VSS.n430 2.6005
R2141 VSS.n430 VSS.n429 2.6005
R2142 VSS.n434 VSS.n433 2.6005
R2143 VSS.n433 VSS.n432 2.6005
R2144 VSS.n437 VSS.n436 2.6005
R2145 VSS.n436 VSS.n435 2.6005
R2146 VSS.n440 VSS.n439 2.6005
R2147 VSS.n439 VSS.n438 2.6005
R2148 VSS.n443 VSS.n442 2.6005
R2149 VSS.n442 VSS.n441 2.6005
R2150 VSS.n446 VSS.n445 2.6005
R2151 VSS.n445 VSS.n444 2.6005
R2152 VSS.n449 VSS.n448 2.6005
R2153 VSS.n448 VSS.n447 2.6005
R2154 VSS.n453 VSS.n452 2.6005
R2155 VSS.n452 VSS.n451 2.6005
R2156 VSS.n457 VSS.n456 2.6005
R2157 VSS.n456 VSS.n455 2.6005
R2158 VSS.n1155 VSS.n1154 2.6005
R2159 VSS.n1154 VSS.n1153 2.6005
R2160 VSS.n1152 VSS.n1151 2.6005
R2161 VSS.n1151 VSS.n1150 2.6005
R2162 VSS.n1148 VSS.n1147 2.6005
R2163 VSS.n1147 VSS.n1146 2.6005
R2164 VSS.n1144 VSS.n1143 2.6005
R2165 VSS.n1143 VSS.n1142 2.6005
R2166 VSS.n1141 VSS.n1140 2.6005
R2167 VSS.n1158 VSS.n1157 2.6005
R2168 VSS.n1157 VSS.n1156 2.6005
R2169 VSS.n529 VSS.n528 2.6005
R2170 VSS.n531 VSS.n530 2.6005
R2171 VSS.n533 VSS.n532 2.6005
R2172 VSS.n535 VSS.n534 2.6005
R2173 VSS.n537 VSS.n536 2.6005
R2174 VSS.n539 VSS.n538 2.6005
R2175 VSS.n541 VSS.n540 2.6005
R2176 VSS.n543 VSS.n542 2.6005
R2177 VSS.n545 VSS.n544 2.6005
R2178 VSS.n547 VSS.n546 2.6005
R2179 VSS.n549 VSS.n548 2.6005
R2180 VSS.n551 VSS.n550 2.6005
R2181 VSS.n553 VSS.n552 2.6005
R2182 VSS.n555 VSS.n554 2.6005
R2183 VSS.n557 VSS.n556 2.6005
R2184 VSS.n559 VSS.n558 2.6005
R2185 VSS.n561 VSS.n560 2.6005
R2186 VSS.n1033 VSS.t100 1.97199
R2187 VSS.n576 VSS.n575 1.90335
R2188 VSS.n113 VSS.n112 1.72783
R2189 VSS.n617 VSS.n616 1.7266
R2190 VSS.n611 VSS.n610 1.7266
R2191 VSS.n605 VSS.n604 1.7266
R2192 VSS.n800 VSS.n799 1.7266
R2193 VSS.n794 VSS.n793 1.7266
R2194 VSS.n788 VSS.n787 1.7266
R2195 VSS.n400 VSS.n399 1.7266
R2196 VSS.n393 VSS.n392 1.7266
R2197 VSS.n388 VSS.n387 1.7266
R2198 VSS.n1436 VSS.n1435 1.72592
R2199 VSS.n1429 VSS.n1428 1.72592
R2200 VSS.n1424 VSS.n1423 1.72592
R2201 VSS.n1528 VSS.n1527 1.69565
R2202 VSS.n1514 VSS.n1513 1.69565
R2203 VSS.n1508 VSS.n1507 1.69507
R2204 VSS.n1519 VSS.n1518 1.69497
R2205 VSS.n485 VSS.n484 1.68203
R2206 VSS.n497 VSS.n496 1.68193
R2207 VSS.n1035 VSS.n1034 1.67823
R2208 VSS.n461 VSS.t73 1.6385
R2209 VSS.n461 VSS.n460 1.6385
R2210 VSS.n459 VSS.t90 1.6385
R2211 VSS.n459 VSS.n458 1.6385
R2212 VSS.n295 VSS.t67 1.6385
R2213 VSS.n295 VSS.n294 1.6385
R2214 VSS.n293 VSS.t91 1.6385
R2215 VSS.n293 VSS.n292 1.6385
R2216 VSS.n780 VSS.t87 1.6385
R2217 VSS.n780 VSS.n779 1.6385
R2218 VSS.n778 VSS.t126 1.6385
R2219 VSS.n778 VSS.n777 1.6385
R2220 VSS.n503 VSS.t124 1.6385
R2221 VSS.n503 VSS.n502 1.6385
R2222 VSS.n597 VSS.t127 1.6385
R2223 VSS.n597 VSS.n596 1.6385
R2224 VSS.n595 VSS.t72 1.6385
R2225 VSS.n595 VSS.n594 1.6385
R2226 VSS.n1038 VSS.t66 1.6385
R2227 VSS.n1038 VSS.n1037 1.6385
R2228 VSS.n1296 VSS.n1295 1.62633
R2229 VSS.n1663 VSS.n1662 1.55471
R2230 VSS.n1734 VSS.n1733 1.55416
R2231 VSS.n194 VSS.n193 1.54032
R2232 VSS.n764 VSS.n763 1.53476
R2233 VSS.n1673 VSS.n1672 1.53464
R2234 VSS.n1666 VSS.n1665 1.53464
R2235 VSS.n163 VSS.n162 1.53464
R2236 VSS.n1737 VSS.n1736 1.53464
R2237 VSS.n1018 VSS.n1017 1.50072
R2238 VSS.n1548 VSS.n1547 1.4928
R2239 VSS VSS.n465 1.46704
R2240 VSS VSS.n299 1.46704
R2241 VSS VSS.n784 1.46704
R2242 VSS VSS.n601 1.46704
R2243 VSS.n167 VSS.n166 1.45083
R2244 VSS.n1679 VSS.n1678 1.4503
R2245 VSS.n1595 VSS.n1594 1.44361
R2246 VSS.n1601 VSS.n1600 1.44361
R2247 VSS.n1253 VSS.n1252 1.36965
R2248 VSS.n1247 VSS.n1246 1.36965
R2249 VSS.n1290 VSS.n1289 1.28498
R2250 VSS.n1355 VSS.n1354 1.27366
R2251 VSS.n1349 VSS.n1348 1.27366
R2252 VSS.n1553 VSS.n1552 1.25894
R2253 VSS.n1181 VSS.t28 1.1705
R2254 VSS.n1181 VSS.n1180 1.1705
R2255 VSS.n951 VSS.t101 1.1705
R2256 VSS.n951 VSS.n950 1.1705
R2257 VSS.n1033 VSS.n1032 1.09725
R2258 VSS.n1138 VSS 1.03013
R2259 VSS VSS.n1137 0.940271
R2260 VSS.n1145 VSS.n524 0.938847
R2261 VSS.n1077 VSS.n1076 0.929805
R2262 VSS.n1091 VSS.n584 0.91886
R2263 VSS.n1354 VSS.n1353 0.885896
R2264 VSS.n464 VSS.n463 0.845717
R2265 VSS.n298 VSS.n297 0.845717
R2266 VSS.n783 VSS.n782 0.845717
R2267 VSS.n600 VSS.n599 0.845717
R2268 VSS.n465 VSS.n464 0.827256
R2269 VSS.n299 VSS.n298 0.827256
R2270 VSS.n784 VSS.n783 0.827256
R2271 VSS.n601 VSS.n600 0.827256
R2272 VSS.n1252 VSS.n1251 0.8219
R2273 VSS.n1600 VSS.n1599 0.772592
R2274 VSS.n1547 VSS.n1546 0.739798
R2275 VSS.n1672 VSS.n1671 0.711907
R2276 VSS.n275 VSS.n195 0.669389
R2277 VSS.n1034 VSS.n1033 0.616183
R2278 VSS.n496 VSS.n495 0.613712
R2279 VSS.n495 VSS.n494 0.613712
R2280 VSS.n495 VSS.n493 0.613712
R2281 VSS.n1643 VSS.n1624 0.606056
R2282 VSS.n1505 VSS.n1504 0.580006
R2283 VSS.n1678 VSS.n1677 0.576657
R2284 VSS.n166 VSS.n165 0.576657
R2285 VSS.n763 VSS.n762 0.53442
R2286 VSS.n193 VSS.n192 0.531916
R2287 VSS.n1662 VSS.n1661 0.52472
R2288 VSS.n1733 VSS.n1732 0.52472
R2289 VSS.n1607 VSS.n1606 0.5185
R2290 VSS.n301 VSS.n300 0.5005
R2291 VSS.n216 VSS.n214 0.5005
R2292 VSS.n674 VSS.n672 0.5005
R2293 VSS.n4 VSS.n2 0.5005
R2294 VSS.n1295 VSS.n1294 0.488634
R2295 VSS.n1507 VSS.n1506 0.454258
R2296 VSS.n1513 VSS.n1512 0.454258
R2297 VSS.n616 VSS.n615 0.438783
R2298 VSS.n799 VSS.n798 0.438783
R2299 VSS.n399 VSS.n398 0.438783
R2300 VSS.n1435 VSS.n1434 0.43854
R2301 VSS.n112 VSS.n111 0.438169
R2302 VSS.n1033 VSS.n1031 0.428289
R2303 VSS.n495 VSS.n492 0.349863
R2304 VSS.n1033 VSS.n1030 0.348521
R2305 VSS.n92 VSS.n91 0.304848
R2306 VSS.n86 VSS.n84 0.304848
R2307 VSS.n526 VSS.n525 0.2505
R2308 VSS.n1363 VSS.n1361 0.2505
R2309 VSS.n1136 VSS.n1135 0.2505
R2310 VSS.n870 VSS.n868 0.2505
R2311 VSS.n1149 VSS 0.224346
R2312 VSS.n1410 VSS 0.224346
R2313 VSS.n792 VSS 0.224346
R2314 VSS.n609 VSS 0.224346
R2315 VSS.n1043 VSS.n1041 0.183918
R2316 VSS.n1045 VSS.n1043 0.183918
R2317 VSS.n1047 VSS.n1045 0.183918
R2318 VSS.n1023 VSS.n1021 0.183918
R2319 VSS.n1026 VSS.n1023 0.183918
R2320 VSS.n1029 VSS.n1026 0.183918
R2321 VSS.n488 VSS.n486 0.183918
R2322 VSS.n491 VSS.n488 0.183918
R2323 VSS.n498 VSS.n491 0.183918
R2324 VSS.n570 VSS.n568 0.183918
R2325 VSS.n572 VSS.n570 0.183918
R2326 VSS.n574 VSS.n572 0.183918
R2327 VSS.n1049 VSS.n1047 0.182778
R2328 VSS.n1036 VSS.n1029 0.182778
R2329 VSS.n500 VSS.n498 0.182778
R2330 VSS.n577 VSS.n574 0.182778
R2331 VSS.n1001 VSS.n998 0.177207
R2332 VSS.n1004 VSS.n1001 0.177207
R2333 VSS.n1007 VSS.n1004 0.177207
R2334 VSS.n1010 VSS.n1007 0.177207
R2335 VSS.n1013 VSS.n1010 0.177207
R2336 VSS.n1016 VSS.n1013 0.177207
R2337 VSS.n1019 VSS.n1016 0.177207
R2338 VSS.n1054 VSS.n1051 0.177207
R2339 VSS.n1061 VSS.n1058 0.177207
R2340 VSS.n1068 VSS.n1065 0.177207
R2341 VSS.n1075 VSS.n1072 0.177207
R2342 VSS.n483 VSS.n480 0.177207
R2343 VSS.n480 VSS.n479 0.177207
R2344 VSS.n479 VSS.n476 0.177207
R2345 VSS.n476 VSS.n473 0.177207
R2346 VSS.n473 VSS.n470 0.177207
R2347 VSS.n566 VSS.n564 0.177207
R2348 VSS.n523 VSS.n520 0.177207
R2349 VSS.n516 VSS.n513 0.177207
R2350 VSS.n509 VSS.n506 0.177207
R2351 VSS.n583 VSS.n581 0.177207
R2352 VSS.n1730 VSS.n1728 0.155256
R2353 VSS.n1695 VSS.n1692 0.1505
R2354 VSS.n1692 VSS.n1689 0.1505
R2355 VSS.n1689 VSS.n1686 0.1505
R2356 VSS.n1686 VSS.n1683 0.1505
R2357 VSS.n1683 VSS.n1680 0.1505
R2358 VSS.n185 VSS.n182 0.1505
R2359 VSS.n182 VSS.n179 0.1505
R2360 VSS.n179 VSS.n176 0.1505
R2361 VSS.n176 VSS.n173 0.1505
R2362 VSS.n173 VSS.n170 0.1505
R2363 VSS.n1366 VSS.n1364 0.149643
R2364 VSS.n1134 VSS.n1133 0.149643
R2365 VSS.n1078 VSS.n671 0.149643
R2366 VSS.n907 VSS.n906 0.149643
R2367 VSS.n854 VSS.n853 0.149643
R2368 VSS.n1449 VSS.n1446 0.149643
R2369 VSS.n407 VSS.n404 0.149643
R2370 VSS.n529 VSS.n527 0.149643
R2371 VSS.n1642 VSS.n1639 0.148671
R2372 VSS.n1639 VSS.n1636 0.148671
R2373 VSS.n1636 VSS.n1633 0.148671
R2374 VSS.n1633 VSS.n1630 0.148671
R2375 VSS.n1630 VSS.n1627 0.148671
R2376 VSS.n1716 VSS.n1713 0.148671
R2377 VSS.n1719 VSS.n1716 0.148671
R2378 VSS.n1722 VSS.n1719 0.148671
R2379 VSS.n1725 VSS.n1722 0.148671
R2380 VSS.n1728 VSS.n1725 0.148671
R2381 VSS.n697 VSS.n694 0.147071
R2382 VSS.n28 VSS.n25 0.147071
R2383 VSS.n268 VSS.n265 0.147071
R2384 VSS.n370 VSS.n367 0.147071
R2385 VSS.n1676 VSS.n1674 0.144731
R2386 VSS.n1674 VSS.n1670 0.144731
R2387 VSS.n1667 VSS.n1664 0.144731
R2388 VSS.n168 VSS.n164 0.144731
R2389 VSS.n164 VSS.n1 0.144731
R2390 VSS.n1738 VSS.n1735 0.144731
R2391 VSS.n1658 VSS.n1655 0.139389
R2392 VSS.n1655 VSS.n1652 0.139389
R2393 VSS.n1652 VSS.n1649 0.139389
R2394 VSS.n1649 VSS.n1646 0.139389
R2395 VSS.n190 VSS.n188 0.139389
R2396 VSS.n1706 VSS.n1703 0.139389
R2397 VSS.n1709 VSS.n1706 0.139389
R2398 VSS.n486 VSS.n483 0.139362
R2399 VSS.n1696 VSS.n1658 0.138278
R2400 VSS.n191 VSS.n190 0.138278
R2401 VSS.n1021 VSS.n1019 0.137167
R2402 VSS.n568 VSS.n566 0.137167
R2403 VSS.n1536 VSS.n1533 0.1355
R2404 VSS.n1539 VSS.n1536 0.1355
R2405 VSS.n1542 VSS.n1539 0.1355
R2406 VSS.n1545 VSS.n1542 0.1355
R2407 VSS.n1549 VSS.n1545 0.1355
R2408 VSS.n1551 VSS.n1549 0.1355
R2409 VSS.n161 VSS.n158 0.1355
R2410 VSS.n158 VSS.n155 0.1355
R2411 VSS.n155 VSS.n152 0.1355
R2412 VSS.n152 VSS.n149 0.1355
R2413 VSS.n149 VSS.n146 0.1355
R2414 VSS.n146 VSS.n143 0.1355
R2415 VSS.n1211 VSS.n1176 0.132808
R2416 VSS.n1593 VSS.n1590 0.132565
R2417 VSS.n1590 VSS.n1587 0.132565
R2418 VSS.n1587 VSS.n1584 0.132565
R2419 VSS.n1584 VSS.n1581 0.132565
R2420 VSS.n1581 VSS.n1578 0.132565
R2421 VSS.n1578 VSS.n1575 0.132565
R2422 VSS.n99 VSS.n95 0.132565
R2423 VSS.n102 VSS.n99 0.132565
R2424 VSS.n105 VSS.n102 0.132565
R2425 VSS.n110 VSS.n105 0.132565
R2426 VSS.n114 VSS.n110 0.132565
R2427 VSS.n116 VSS.n114 0.132565
R2428 VSS.n1406 VSS.n1360 0.132449
R2429 VSS.n1437 VSS.n1432 0.132286
R2430 VSS.n1432 VSS.n1430 0.132286
R2431 VSS.n1430 VSS.n1427 0.132286
R2432 VSS.n1427 VSS.n1425 0.132286
R2433 VSS.n1425 VSS.n1422 0.132286
R2434 VSS.n1368 VSS.n1366 0.132286
R2435 VSS.n1370 VSS.n1368 0.132286
R2436 VSS.n1372 VSS.n1370 0.132286
R2437 VSS.n1374 VSS.n1372 0.132286
R2438 VSS.n1376 VSS.n1374 0.132286
R2439 VSS.n1378 VSS.n1376 0.132286
R2440 VSS.n1380 VSS.n1378 0.132286
R2441 VSS.n1382 VSS.n1380 0.132286
R2442 VSS.n1384 VSS.n1382 0.132286
R2443 VSS.n1386 VSS.n1384 0.132286
R2444 VSS.n1388 VSS.n1386 0.132286
R2445 VSS.n1390 VSS.n1388 0.132286
R2446 VSS.n1392 VSS.n1390 0.132286
R2447 VSS.n1394 VSS.n1392 0.132286
R2448 VSS.n1396 VSS.n1394 0.132286
R2449 VSS.n1084 VSS.n1081 0.132286
R2450 VSS.n1087 VSS.n1084 0.132286
R2451 VSS.n1090 VSS.n1087 0.132286
R2452 VSS.n1097 VSS.n1094 0.132286
R2453 VSS.n1133 VSS.n1131 0.132286
R2454 VSS.n1131 VSS.n1129 0.132286
R2455 VSS.n1129 VSS.n1127 0.132286
R2456 VSS.n1127 VSS.n1125 0.132286
R2457 VSS.n1125 VSS.n1123 0.132286
R2458 VSS.n1123 VSS.n1121 0.132286
R2459 VSS.n1121 VSS.n1119 0.132286
R2460 VSS.n1119 VSS.n1117 0.132286
R2461 VSS.n1117 VSS.n1115 0.132286
R2462 VSS.n1115 VSS.n1113 0.132286
R2463 VSS.n1113 VSS.n1111 0.132286
R2464 VSS.n1111 VSS.n1109 0.132286
R2465 VSS.n1109 VSS.n1107 0.132286
R2466 VSS.n1107 VSS.n1105 0.132286
R2467 VSS.n1105 VSS.n1103 0.132286
R2468 VSS.n742 VSS.n738 0.132286
R2469 VSS.n738 VSS.n735 0.132286
R2470 VSS.n735 VSS.n732 0.132286
R2471 VSS.n732 VSS.n729 0.132286
R2472 VSS.n729 VSS.n726 0.132286
R2473 VSS.n726 VSS.n723 0.132286
R2474 VSS.n723 VSS.n721 0.132286
R2475 VSS.n721 VSS.n718 0.132286
R2476 VSS.n718 VSS.n715 0.132286
R2477 VSS.n715 VSS.n712 0.132286
R2478 VSS.n712 VSS.n709 0.132286
R2479 VSS.n709 VSS.n706 0.132286
R2480 VSS.n706 VSS.n703 0.132286
R2481 VSS.n703 VSS.n700 0.132286
R2482 VSS.n700 VSS.n697 0.132286
R2483 VSS.n693 VSS.n690 0.132286
R2484 VSS.n690 VSS.n687 0.132286
R2485 VSS.n687 VSS.n684 0.132286
R2486 VSS.n684 VSS.n681 0.132286
R2487 VSS.n681 VSS.n678 0.132286
R2488 VSS.n593 VSS.n590 0.132286
R2489 VSS.n618 VSS.n614 0.132286
R2490 VSS.n614 VSS.n612 0.132286
R2491 VSS.n608 VSS.n606 0.132286
R2492 VSS.n606 VSS.n603 0.132286
R2493 VSS.n671 VSS.n667 0.132286
R2494 VSS.n667 VSS.n664 0.132286
R2495 VSS.n664 VSS.n661 0.132286
R2496 VSS.n661 VSS.n658 0.132286
R2497 VSS.n658 VSS.n655 0.132286
R2498 VSS.n655 VSS.n652 0.132286
R2499 VSS.n652 VSS.n649 0.132286
R2500 VSS.n649 VSS.n646 0.132286
R2501 VSS.n646 VSS.n643 0.132286
R2502 VSS.n643 VSS.n640 0.132286
R2503 VSS.n640 VSS.n637 0.132286
R2504 VSS.n637 VSS.n634 0.132286
R2505 VSS.n634 VSS.n631 0.132286
R2506 VSS.n631 VSS.n628 0.132286
R2507 VSS.n628 VSS.n625 0.132286
R2508 VSS.n749 VSS.n746 0.132286
R2509 VSS.n984 VSS.n981 0.132286
R2510 VSS.n987 VSS.n984 0.132286
R2511 VSS.n990 VSS.n987 0.132286
R2512 VSS.n993 VSS.n990 0.132286
R2513 VSS.n996 VSS.n993 0.132286
R2514 VSS.n906 VSS.n904 0.132286
R2515 VSS.n904 VSS.n902 0.132286
R2516 VSS.n902 VSS.n900 0.132286
R2517 VSS.n900 VSS.n898 0.132286
R2518 VSS.n898 VSS.n896 0.132286
R2519 VSS.n896 VSS.n894 0.132286
R2520 VSS.n894 VSS.n892 0.132286
R2521 VSS.n892 VSS.n890 0.132286
R2522 VSS.n890 VSS.n888 0.132286
R2523 VSS.n888 VSS.n886 0.132286
R2524 VSS.n886 VSS.n884 0.132286
R2525 VSS.n884 VSS.n882 0.132286
R2526 VSS.n882 VSS.n880 0.132286
R2527 VSS.n880 VSS.n878 0.132286
R2528 VSS.n878 VSS.n876 0.132286
R2529 VSS.n861 VSS.n857 0.132286
R2530 VSS.n864 VSS.n861 0.132286
R2531 VSS.n867 VSS.n864 0.132286
R2532 VSS.n913 VSS.n910 0.132286
R2533 VSS.n73 VSS.n70 0.132286
R2534 VSS.n70 VSS.n67 0.132286
R2535 VSS.n67 VSS.n64 0.132286
R2536 VSS.n64 VSS.n61 0.132286
R2537 VSS.n61 VSS.n58 0.132286
R2538 VSS.n58 VSS.n55 0.132286
R2539 VSS.n55 VSS.n52 0.132286
R2540 VSS.n52 VSS.n49 0.132286
R2541 VSS.n49 VSS.n46 0.132286
R2542 VSS.n46 VSS.n43 0.132286
R2543 VSS.n43 VSS.n40 0.132286
R2544 VSS.n40 VSS.n37 0.132286
R2545 VSS.n37 VSS.n34 0.132286
R2546 VSS.n34 VSS.n31 0.132286
R2547 VSS.n31 VSS.n28 0.132286
R2548 VSS.n22 VSS.n19 0.132286
R2549 VSS.n19 VSS.n16 0.132286
R2550 VSS.n16 VSS.n13 0.132286
R2551 VSS.n13 VSS.n10 0.132286
R2552 VSS.n10 VSS.n7 0.132286
R2553 VSS.n776 VSS.n773 0.132286
R2554 VSS.n801 VSS.n797 0.132286
R2555 VSS.n797 VSS.n795 0.132286
R2556 VSS.n791 VSS.n789 0.132286
R2557 VSS.n789 VSS.n786 0.132286
R2558 VSS.n853 VSS.n850 0.132286
R2559 VSS.n850 VSS.n847 0.132286
R2560 VSS.n847 VSS.n844 0.132286
R2561 VSS.n844 VSS.n841 0.132286
R2562 VSS.n841 VSS.n838 0.132286
R2563 VSS.n838 VSS.n835 0.132286
R2564 VSS.n835 VSS.n832 0.132286
R2565 VSS.n832 VSS.n829 0.132286
R2566 VSS.n829 VSS.n826 0.132286
R2567 VSS.n826 VSS.n823 0.132286
R2568 VSS.n823 VSS.n820 0.132286
R2569 VSS.n820 VSS.n817 0.132286
R2570 VSS.n817 VSS.n814 0.132286
R2571 VSS.n814 VSS.n811 0.132286
R2572 VSS.n811 VSS.n808 0.132286
R2573 VSS.n80 VSS.n77 0.132286
R2574 VSS.n1623 VSS.n1620 0.132286
R2575 VSS.n1620 VSS.n1616 0.132286
R2576 VSS.n1616 VSS.n1613 0.132286
R2577 VSS.n1613 VSS.n1610 0.132286
R2578 VSS.n274 VSS.n271 0.132286
R2579 VSS.n282 VSS.n278 0.132286
R2580 VSS.n285 VSS.n282 0.132286
R2581 VSS.n288 VSS.n285 0.132286
R2582 VSS.n291 VSS.n288 0.132286
R2583 VSS.n1420 VSS.n1417 0.132286
R2584 VSS.n1417 VSS.n1413 0.132286
R2585 VSS.n1405 VSS.n1402 0.132286
R2586 VSS.n1452 VSS.n1449 0.132286
R2587 VSS.n1455 VSS.n1452 0.132286
R2588 VSS.n1458 VSS.n1455 0.132286
R2589 VSS.n1461 VSS.n1458 0.132286
R2590 VSS.n1464 VSS.n1461 0.132286
R2591 VSS.n1467 VSS.n1464 0.132286
R2592 VSS.n1470 VSS.n1467 0.132286
R2593 VSS.n1473 VSS.n1470 0.132286
R2594 VSS.n1476 VSS.n1473 0.132286
R2595 VSS.n1479 VSS.n1476 0.132286
R2596 VSS.n1482 VSS.n1479 0.132286
R2597 VSS.n1485 VSS.n1482 0.132286
R2598 VSS.n1488 VSS.n1485 0.132286
R2599 VSS.n1491 VSS.n1488 0.132286
R2600 VSS.n1495 VSS.n1491 0.132286
R2601 VSS.n213 VSS.n210 0.132286
R2602 VSS.n210 VSS.n207 0.132286
R2603 VSS.n207 VSS.n204 0.132286
R2604 VSS.n204 VSS.n201 0.132286
R2605 VSS.n201 VSS.n198 0.132286
R2606 VSS.n1445 VSS.n1442 0.132286
R2607 VSS.n223 VSS.n220 0.132286
R2608 VSS.n226 VSS.n223 0.132286
R2609 VSS.n229 VSS.n226 0.132286
R2610 VSS.n232 VSS.n229 0.132286
R2611 VSS.n235 VSS.n232 0.132286
R2612 VSS.n238 VSS.n235 0.132286
R2613 VSS.n241 VSS.n238 0.132286
R2614 VSS.n244 VSS.n241 0.132286
R2615 VSS.n247 VSS.n244 0.132286
R2616 VSS.n250 VSS.n247 0.132286
R2617 VSS.n253 VSS.n250 0.132286
R2618 VSS.n256 VSS.n253 0.132286
R2619 VSS.n259 VSS.n256 0.132286
R2620 VSS.n262 VSS.n259 0.132286
R2621 VSS.n265 VSS.n262 0.132286
R2622 VSS.n376 VSS.n373 0.132286
R2623 VSS.n1175 VSS.n1174 0.132286
R2624 VSS.n1174 VSS.n1171 0.132286
R2625 VSS.n1171 VSS.n1168 0.132286
R2626 VSS.n1168 VSS.n1165 0.132286
R2627 VSS.n1165 VSS.n1162 0.132286
R2628 VSS.n326 VSS.n323 0.132286
R2629 VSS.n329 VSS.n326 0.132286
R2630 VSS.n332 VSS.n329 0.132286
R2631 VSS.n335 VSS.n332 0.132286
R2632 VSS.n338 VSS.n335 0.132286
R2633 VSS.n340 VSS.n338 0.132286
R2634 VSS.n343 VSS.n340 0.132286
R2635 VSS.n346 VSS.n343 0.132286
R2636 VSS.n349 VSS.n346 0.132286
R2637 VSS.n352 VSS.n349 0.132286
R2638 VSS.n355 VSS.n352 0.132286
R2639 VSS.n358 VSS.n355 0.132286
R2640 VSS.n361 VSS.n358 0.132286
R2641 VSS.n364 VSS.n361 0.132286
R2642 VSS.n367 VSS.n364 0.132286
R2643 VSS.n319 VSS.n316 0.132286
R2644 VSS.n316 VSS.n313 0.132286
R2645 VSS.n313 VSS.n310 0.132286
R2646 VSS.n310 VSS.n307 0.132286
R2647 VSS.n307 VSS.n304 0.132286
R2648 VSS.n384 VSS.n381 0.132286
R2649 VSS.n401 VSS.n396 0.132286
R2650 VSS.n396 VSS.n394 0.132286
R2651 VSS.n394 VSS.n391 0.132286
R2652 VSS.n391 VSS.n389 0.132286
R2653 VSS.n389 VSS.n386 0.132286
R2654 VSS.n410 VSS.n407 0.132286
R2655 VSS.n413 VSS.n410 0.132286
R2656 VSS.n416 VSS.n413 0.132286
R2657 VSS.n419 VSS.n416 0.132286
R2658 VSS.n422 VSS.n419 0.132286
R2659 VSS.n425 VSS.n422 0.132286
R2660 VSS.n428 VSS.n425 0.132286
R2661 VSS.n431 VSS.n428 0.132286
R2662 VSS.n434 VSS.n431 0.132286
R2663 VSS.n437 VSS.n434 0.132286
R2664 VSS.n440 VSS.n437 0.132286
R2665 VSS.n443 VSS.n440 0.132286
R2666 VSS.n446 VSS.n443 0.132286
R2667 VSS.n449 VSS.n446 0.132286
R2668 VSS.n453 VSS.n449 0.132286
R2669 VSS.n1158 VSS.n1155 0.132286
R2670 VSS.n1155 VSS.n1152 0.132286
R2671 VSS.n1144 VSS.n1141 0.132286
R2672 VSS.n531 VSS.n529 0.132286
R2673 VSS.n533 VSS.n531 0.132286
R2674 VSS.n535 VSS.n533 0.132286
R2675 VSS.n537 VSS.n535 0.132286
R2676 VSS.n539 VSS.n537 0.132286
R2677 VSS.n541 VSS.n539 0.132286
R2678 VSS.n543 VSS.n541 0.132286
R2679 VSS.n545 VSS.n543 0.132286
R2680 VSS.n547 VSS.n545 0.132286
R2681 VSS.n549 VSS.n547 0.132286
R2682 VSS.n551 VSS.n549 0.132286
R2683 VSS.n553 VSS.n551 0.132286
R2684 VSS.n555 VSS.n553 0.132286
R2685 VSS.n557 VSS.n555 0.132286
R2686 VSS.n559 VSS.n557 0.132286
R2687 VSS.n1605 VSS.n1593 0.128652
R2688 VSS.n1523 VSS.n95 0.128652
R2689 VSS.n1331 VSS.n1276 0.127656
R2690 VSS.n922 VSS.n919 0.127656
R2691 VSS.n743 VSS.n742 0.125857
R2692 VSS.n74 VSS.n73 0.125857
R2693 VSS.n220 VSS.n217 0.125857
R2694 VSS.n323 VSS.n320 0.125857
R2695 VSS.n1557 VSS.n1554 0.1255
R2696 VSS.n1564 VSS.n1561 0.1255
R2697 VSS.n140 VSS.n137 0.1255
R2698 VSS.n133 VSS.n130 0.1255
R2699 VSS.n1330 VSS.n1326 0.125187
R2700 VSS.n1529 VSS.n1526 0.124126
R2701 VSS.n1598 VSS.n1596 0.124126
R2702 VSS.n1602 VSS.n1598 0.124126
R2703 VSS.n1604 VSS.n1602 0.124126
R2704 VSS.n1511 VSS.n1509 0.124126
R2705 VSS.n1515 VSS.n1511 0.124126
R2706 VSS.n1517 VSS.n1515 0.124126
R2707 VSS.n1520 VSS.n1517 0.124126
R2708 VSS.n1522 VSS.n1520 0.124126
R2709 VSS.n609 VSS.n608 0.123929
R2710 VSS.n792 VSS.n791 0.123929
R2711 VSS.n1410 VSS.n1409 0.123929
R2712 VSS.n1149 VSS.n1148 0.123929
R2713 VSS.n625 VSS.n622 0.123286
R2714 VSS.n808 VSS.n805 0.123286
R2715 VSS.n1499 VSS.n1495 0.123286
R2716 VSS.n457 VSS.n453 0.123286
R2717 VSS.n1399 VSS.n1396 0.122
R2718 VSS.n561 VSS.n559 0.122
R2719 VSS.n1360 VSS.n1241 0.12105
R2720 VSS.n1326 VSS.n1316 0.12105
R2721 VSS.n1329 VSS.n1327 0.120158
R2722 VSS.n917 VSS.n915 0.120158
R2723 VSS.n1211 VSS.n1210 0.119731
R2724 VSS.n1288 VSS.n1287 0.119731
R2725 VSS.n978 VSS.n977 0.118962
R2726 VSS.n1334 VSS.n1331 0.117958
R2727 VSS.n919 VSS.n767 0.117958
R2728 VSS.n1069 VSS.n1068 0.117939
R2729 VSS.n1668 VSS 0.117309
R2730 VSS VSS.n1739 0.117309
R2731 VSS.n918 VSS.n914 0.117084
R2732 VSS.n1058 VSS.n1055 0.116841
R2733 VSS.n517 VSS.n516 0.116841
R2734 VSS.n1696 VSS.n1695 0.114944
R2735 VSS.n191 VSS.n185 0.113833
R2736 VSS.n1670 VSS.n1668 0.112423
R2737 VSS.n1739 VSS.n1 0.112423
R2738 VSS.n1276 VSS.n1273 0.111968
R2739 VSS.n1273 VSS.n1270 0.111968
R2740 VSS.n1270 VSS.n1267 0.111968
R2741 VSS.n1267 VSS.n1264 0.111968
R2742 VSS.n1264 VSS.n1261 0.111968
R2743 VSS.n1261 VSS.n1258 0.111968
R2744 VSS.n1258 VSS.n1254 0.111968
R2745 VSS.n1254 VSS.n1250 0.111968
R2746 VSS.n1250 VSS.n1248 0.111968
R2747 VSS.n1241 VSS.n1238 0.111968
R2748 VSS.n1238 VSS.n1235 0.111968
R2749 VSS.n1235 VSS.n1232 0.111968
R2750 VSS.n1232 VSS.n1229 0.111968
R2751 VSS.n1229 VSS.n1226 0.111968
R2752 VSS.n1226 VSS.n1223 0.111968
R2753 VSS.n1223 VSS.n1220 0.111968
R2754 VSS.n1220 VSS.n1217 0.111968
R2755 VSS.n1217 VSS.n1214 0.111968
R2756 VSS.n1316 VSS.n1315 0.111968
R2757 VSS.n1315 VSS.n1312 0.111968
R2758 VSS.n1312 VSS.n1309 0.111968
R2759 VSS.n1309 VSS.n1306 0.111968
R2760 VSS.n1306 VSS.n1303 0.111968
R2761 VSS.n1303 VSS.n1300 0.111968
R2762 VSS.n1300 VSS.n1297 0.111968
R2763 VSS.n1297 VSS.n1293 0.111968
R2764 VSS.n1293 VSS.n1291 0.111968
R2765 VSS.n925 VSS.n922 0.111968
R2766 VSS.n928 VSS.n925 0.111968
R2767 VSS.n931 VSS.n928 0.111968
R2768 VSS.n934 VSS.n931 0.111968
R2769 VSS.n937 VSS.n934 0.111968
R2770 VSS.n940 VSS.n937 0.111968
R2771 VSS.n943 VSS.n940 0.111968
R2772 VSS.n946 VSS.n943 0.111968
R2773 VSS.n949 VSS.n946 0.111968
R2774 VSS.n1710 VSS.n1700 0.107167
R2775 VSS.n978 VSS.n749 0.105286
R2776 VSS.n1176 VSS.n376 0.105286
R2777 VSS.n619 VSS.n593 0.102071
R2778 VSS.n802 VSS.n776 0.102071
R2779 VSS.n854 VSS.n83 0.102071
R2780 VSS.n1503 VSS.n1500 0.102071
R2781 VSS.n1446 VSS.n1445 0.102071
R2782 VSS.n1162 VSS.n1159 0.102071
R2783 VSS.n404 VSS.n384 0.102071
R2784 VSS.n1530 VSS.n1524 0.101005
R2785 VSS.n403 VSS.n402 0.1005
R2786 VSS.n456 VSS.n454 0.1005
R2787 VSS.n1439 VSS.n1438 0.1005
R2788 VSS.n1498 VSS.n1496 0.1005
R2789 VSS.n587 VSS.n585 0.1005
R2790 VSS.n621 VSS.n620 0.1005
R2791 VSS.n770 VSS.n768 0.1005
R2792 VSS.n804 VSS.n803 0.1005
R2793 VSS.n1664 VSS.n1660 0.0996745
R2794 VSS.n1735 VSS.n1730 0.0996745
R2795 VSS.n1575 VSS.n1572 0.0983261
R2796 VSS.n120 VSS.n116 0.0983261
R2797 VSS.n1205 VSS.n1202 0.0966538
R2798 VSS.n1202 VSS.n1199 0.0966538
R2799 VSS.n1195 VSS.n1192 0.0966538
R2800 VSS.n1192 VSS.n1188 0.0966538
R2801 VSS.n958 VSS.n955 0.0966538
R2802 VSS.n965 VSS.n962 0.0966538
R2803 VSS.n968 VSS.n965 0.0966538
R2804 VSS.n976 VSS.n973 0.0966538
R2805 VSS.n694 VSS.n693 0.0962857
R2806 VSS.n25 VSS.n22 0.0962857
R2807 VSS.n271 VSS.n268 0.0962857
R2808 VSS.n373 VSS.n370 0.0962857
R2809 VSS.n1359 VSS.n1356 0.095839
R2810 VSS.n1356 VSS.n1352 0.095839
R2811 VSS.n1352 VSS.n1350 0.095839
R2812 VSS.n1350 VSS.n1347 0.095839
R2813 VSS.n1347 VSS.n1343 0.095839
R2814 VSS.n1343 VSS.n1340 0.095839
R2815 VSS.n1340 VSS.n1337 0.095839
R2816 VSS.n1337 VSS.n1334 0.095839
R2817 VSS.n1325 VSS.n1322 0.095839
R2818 VSS.n1322 VSS.n1319 0.095839
R2819 VSS.n755 VSS.n752 0.095839
R2820 VSS.n759 VSS.n755 0.095839
R2821 VSS.n761 VSS.n759 0.095839
R2822 VSS.n765 VSS.n761 0.095839
R2823 VSS.n767 VSS.n765 0.095839
R2824 VSS.n275 VSS.n274 0.0956429
R2825 VSS.n746 VSS.n743 0.095
R2826 VSS.n77 VSS.n74 0.095
R2827 VSS.n1624 VSS.n80 0.095
R2828 VSS.n217 VSS.n213 0.095
R2829 VSS.n320 VSS.n319 0.095
R2830 VSS.n1554 VSS.n1551 0.0945
R2831 VSS.n143 VSS.n140 0.0945
R2832 VSS.n1062 VSS.n1061 0.0894024
R2833 VSS.n513 VSS.n510 0.0894024
R2834 VSS.n1065 VSS.n1062 0.0883049
R2835 VSS.n510 VSS.n509 0.0883049
R2836 VSS.n1185 VSS.n1184 0.0858846
R2837 VSS.n973 VSS.n969 0.0858846
R2838 VSS.n1680 VSS.n1676 0.084688
R2839 VSS.n170 VSS.n168 0.084688
R2840 VSS.n1078 VSS.n1077 0.0827857
R2841 VSS.n1402 VSS.n1399 0.0821429
R2842 VSS.n1646 VSS.n1643 0.0816111
R2843 VSS.n1710 VSS.n1709 0.0816111
R2844 VSS.n1571 VSS.n1568 0.0815
R2845 VSS.n124 VSS.n123 0.0815
R2846 VSS.n1605 VSS.n1604 0.0806099
R2847 VSS.n1523 VSS.n1522 0.0806099
R2848 VSS.n1572 VSS.n1571 0.0805
R2849 VSS.n123 VSS.n120 0.0805
R2850 VSS.n1094 VSS.n1091 0.0795714
R2851 VSS.n1134 VSS.n1097 0.0795714
R2852 VSS.n1103 VSS.n1101 0.0795714
R2853 VSS.n876 VSS.n874 0.0795714
R2854 VSS.n910 VSS.n907 0.0795714
R2855 VSS.n1145 VSS.n1144 0.0795714
R2856 VSS.n1141 VSS.n1138 0.0795714
R2857 VSS.n119 VSS.n117 0.076587
R2858 VSS.n89 VSS.n87 0.076587
R2859 VSS.n914 VSS.n913 0.0757143
R2860 VSS.n1406 VSS.n1405 0.0750714
R2861 VSS.n1446 VSS.n1437 0.0725
R2862 VSS.n1081 VSS.n1078 0.0725
R2863 VSS.n619 VSS.n618 0.0725
R2864 VSS.n857 VSS.n854 0.0725
R2865 VSS.n802 VSS.n801 0.0725
R2866 VSS.n1558 VSS.n1557 0.0725
R2867 VSS.n137 VSS.n134 0.0725
R2868 VSS.n1500 VSS.n1420 0.0725
R2869 VSS.n404 VSS.n401 0.0725
R2870 VSS.n1159 VSS.n1158 0.0725
R2871 VSS.n1607 VSS.n83 0.0692857
R2872 VSS.n1051 VSS.n1049 0.0687711
R2873 VSS.n1504 VSS.n1503 0.0686429
R2874 VSS.n1076 VSS.n1036 0.066576
R2875 VSS.n524 VSS.n500 0.066576
R2876 VSS.n584 VSS.n577 0.066576
R2877 VSS.n1214 VSS.n1211 0.0657294
R2878 VSS.n1291 VSS.n1288 0.0657294
R2879 VSS.n1567 VSS 0.0655
R2880 VSS VSS.n127 0.0655
R2881 VSS.n1196 VSS.n1195 0.0651154
R2882 VSS.n962 VSS.n959 0.0651154
R2883 VSS.n1504 VSS.n291 0.0641429
R2884 VSS.n1610 VSS.n1607 0.0635
R2885 VSS.n1055 VSS.n1054 0.0608659
R2886 VSS.n520 VSS.n517 0.0608659
R2887 VSS VSS.n1564 0.0605
R2888 VSS.n130 VSS 0.0605
R2889 VSS.n1072 VSS.n1069 0.0597683
R2890 VSS.n581 VSS.n578 0.0597683
R2891 VSS.n1248 VSS.n1245 0.0591239
R2892 VSS.n977 VSS.n949 0.0591239
R2893 VSS.n1409 VSS.n1406 0.0577143
R2894 VSS.n914 VSS.n867 0.0570714
R2895 VSS.n1561 VSS.n1558 0.0535
R2896 VSS.n134 VSS.n133 0.0535
R2897 VSS.n1091 VSS.n1090 0.0532143
R2898 VSS.n1148 VSS.n1145 0.0532143
R2899 VSS.n1210 VSS.n1206 0.0528077
R2900 VSS.n1287 VSS.n1284 0.0528077
R2901 VSS.n1533 VSS.n1530 0.0525
R2902 VSS.n1505 VSS.n161 0.0525
R2903 VSS.n1568 VSS.n1567 0.0445
R2904 VSS.n127 VSS.n124 0.0445
R2905 VSS.n1206 VSS.n1205 0.0443462
R2906 VSS.n1284 VSS.n1283 0.0443462
R2907 VSS.n578 VSS 0.0396304
R2908 VSS.n1069 VSS 0.0396304
R2909 VSS.n1624 VSS.n1623 0.0377857
R2910 VSS.n278 VSS.n275 0.0371429
R2911 VSS.n1668 VSS.n1667 0.0328077
R2912 VSS.n1739 VSS.n1738 0.0328077
R2913 VSS.n1199 VSS.n1196 0.0320385
R2914 VSS.n959 VSS.n958 0.0320385
R2915 VSS.n981 VSS.n978 0.0275
R2916 VSS.n1176 VSS.n1175 0.0275
R2917 VSS.n1196 VSS 0.0239783
R2918 VSS.n959 VSS 0.0239783
R2919 VSS.n1077 VSS.n996 0.0197857
R2920 VSS.n1140 VSS.n1139 0.0129258
R2921 VSS.n1188 VSS.n1185 0.0112692
R2922 VSS.n969 VSS.n968 0.0112692
R2923 VSS.n612 VSS.n609 0.00885714
R2924 VSS.n795 VSS.n792 0.00885714
R2925 VSS.n1413 VSS.n1410 0.00885714
R2926 VSS.n1152 VSS.n1149 0.00885714
R2927 VSS.n1530 VSS.n1529 0.00445604
R2928 VSS.n1509 VSS.n1505 0.00445604
R2929 VSS.n1137 VSS.n1134 0.00371429
R2930 VSS.n1138 VSS.n561 0.00307143
R2931 VSS.n1643 VSS.n1642 0.00269512
R2932 VSS.n1076 VSS.n1075 0.00269512
R2933 VSS.n524 VSS.n523 0.00269512
R2934 VSS.n584 VSS.n583 0.00269512
R2935 VSS.n1360 VSS.n1359 0.00202542
R2936 VSS.n1331 VSS.n1330 0.00202542
R2937 VSS.n1326 VSS.n1325 0.00202542
R2938 VSS.n919 VSS.n918 0.00202542
R2939 VSS.n622 VSS.n619 0.00178571
R2940 VSS.n805 VSS.n802 0.00178571
R2941 VSS.n1500 VSS.n1499 0.00178571
R2942 VSS.n1159 VSS.n457 0.00178571
R2943 VSS.n1700 VSS.n1696 0.00161111
R2944 VSS.n195 VSS.n191 0.00161111
R2945 VSS.n1713 VSS.n1710 0.00159756
R2946 VSS.n1606 VSS.n1605 0.00147826
R2947 VSS.n1524 VSS.n1523 0.00147826
R2948 VSS.n1245 VSS.n1244 0.00126923
R2949 VSS.n977 VSS.n976 0.00126923
R2950 Delay_Cell_mag_1.INB.n13 Delay_Cell_mag_1.INB.t22 22.3568
R2951 Delay_Cell_mag_1.INB.n2 Delay_Cell_mag_1.INB.t6 22.096
R2952 Delay_Cell_mag_1.INB.n25 Delay_Cell_mag_1.INB.t21 21.8182
R2953 Delay_Cell_mag_1.INB.n12 Delay_Cell_mag_1.INB.t24 19.4889
R2954 Delay_Cell_mag_1.INB.n28 Delay_Cell_mag_1.INB.t19 17.2487
R2955 Delay_Cell_mag_1.INB.n3 Delay_Cell_mag_1.INB.n2 14.0791
R2956 Delay_Cell_mag_1.INB.n4 Delay_Cell_mag_1.INB.n3 14.0791
R2957 Delay_Cell_mag_1.INB.n26 Delay_Cell_mag_1.INB.n25 12.6801
R2958 Delay_Cell_mag_1.INB.n28 Delay_Cell_mag_1.INB.t17 12.2493
R2959 Delay_Cell_mag_1.INB.n27 Delay_Cell_mag_1.INB.t16 12.0585
R2960 Delay_Cell_mag_1.INB.n27 Delay_Cell_mag_1.INB.n26 9.76014
R2961 Delay_Cell_mag_1.INB.n14 Delay_Cell_mag_1.INB.n13 9.33211
R2962 Delay_Cell_mag_1.INB.n13 Delay_Cell_mag_1.INB.t23 8.27818
R2963 Delay_Cell_mag_1.INB.n11 Delay_Cell_mag_1.INB.t27 8.27818
R2964 Delay_Cell_mag_1.INB.n2 Delay_Cell_mag_1.INB.t4 8.01746
R2965 Delay_Cell_mag_1.INB.n3 Delay_Cell_mag_1.INB.t2 8.01746
R2966 Delay_Cell_mag_1.INB.n4 Delay_Cell_mag_1.INB.t0 8.01746
R2967 Delay_Cell_mag_1.INB.n25 Delay_Cell_mag_1.INB.t20 6.51836
R2968 Delay_Cell_mag_1.INB.n26 Delay_Cell_mag_1.INB.t26 6.51836
R2969 Delay_Cell_mag_1.INB.n19 Delay_Cell_mag_1.INB.n18 4.67659
R2970 Delay_Cell_mag_1.INB.n29 Delay_Cell_mag_1.INB 4.34457
R2971 Delay_Cell_mag_1.INB Delay_Cell_mag_1.INB.n28 4.1467
R2972 Delay_Cell_mag_1.INB.n29 Delay_Cell_mag_1.INB 4.06926
R2973 Delay_Cell_mag_1.INB.n0 Delay_Cell_mag_1.INB.n19 3.51328
R2974 Delay_Cell_mag_1.INB.n24 Delay_Cell_mag_1.INB.n8 3.20507
R2975 Delay_Cell_mag_1.INB.n19 Delay_Cell_mag_1.INB.n16 3.1505
R2976 Delay_Cell_mag_1.INB.n23 Delay_Cell_mag_1.INB.n22 3.02311
R2977 Delay_Cell_mag_1.INB.n24 Delay_Cell_mag_1.INB.n6 2.98985
R2978 Delay_Cell_mag_1.INB.n12 Delay_Cell_mag_1.INB.n11 2.86836
R2979 Delay_Cell_mag_1.INB.n1 Delay_Cell_mag_1.INB.n4 2.63789
R2980 Delay_Cell_mag_1.INB.n20 Delay_Cell_mag_1.INB.n10 2.6005
R2981 Delay_Cell_mag_1.INB Delay_Cell_mag_1.INB.n27 2.55586
R2982 Delay_Cell_mag_1.INB.n1 Delay_Cell_mag_1.INB.n29 2.17974
R2983 Delay_Cell_mag_1.INB.n0 Delay_Cell_mag_1.INB.n12 2.11815
R2984 Delay_Cell_mag_1.INB.n10 Delay_Cell_mag_1.INB.t10 1.8205
R2985 Delay_Cell_mag_1.INB.n10 Delay_Cell_mag_1.INB.n9 1.8205
R2986 Delay_Cell_mag_1.INB.n8 Delay_Cell_mag_1.INB.t12 1.8205
R2987 Delay_Cell_mag_1.INB.n8 Delay_Cell_mag_1.INB.n7 1.8205
R2988 Delay_Cell_mag_1.INB.n6 Delay_Cell_mag_1.INB.t3 1.8205
R2989 Delay_Cell_mag_1.INB.n6 Delay_Cell_mag_1.INB.n5 1.8205
R2990 Delay_Cell_mag_1.INB.n22 Delay_Cell_mag_1.INB.t7 1.8205
R2991 Delay_Cell_mag_1.INB.n22 Delay_Cell_mag_1.INB.n21 1.8205
R2992 Delay_Cell_mag_1.INB.n16 Delay_Cell_mag_1.INB.t9 1.6385
R2993 Delay_Cell_mag_1.INB.n16 Delay_Cell_mag_1.INB.n15 1.6385
R2994 Delay_Cell_mag_1.INB.n18 Delay_Cell_mag_1.INB.t14 1.6385
R2995 Delay_Cell_mag_1.INB.n18 Delay_Cell_mag_1.INB.n17 1.6385
R2996 Delay_Cell_mag_1.INB.n0 Delay_Cell_mag_1.INB.n14 1.50108
R2997 Delay_Cell_mag_1.INB.n20 Delay_Cell_mag_1.INB.n0 1.32596
R2998 Delay_Cell_mag_1.INB.n24 Delay_Cell_mag_1.INB.n23 0.826273
R2999 Delay_Cell_mag_1.INB.n23 Delay_Cell_mag_1.INB.n20 0.640283
R3000 Delay_Cell_mag_1.INB Delay_Cell_mag_1.INB.n1 0.16328
R3001 Delay_Cell_mag_1.INB.n1 Delay_Cell_mag_1.INB.n24 0.123037
R3002 Delay_Cell_mag_0.OUTB.n23 Delay_Cell_mag_0.OUTB.t22 22.2916
R3003 Delay_Cell_mag_0.OUTB.n7 Delay_Cell_mag_0.OUTB.t10 22.1612
R3004 Delay_Cell_mag_0.OUTB.n0 Delay_Cell_mag_0.OUTB.t25 21.774
R3005 Delay_Cell_mag_0.OUTB.t22 Delay_Cell_mag_0.OUTB.n22 17.311
R3006 Delay_Cell_mag_0.OUTB.n9 Delay_Cell_mag_0.OUTB.t4 15.1219
R3007 Delay_Cell_mag_0.OUTB.n24 Delay_Cell_mag_0.OUTB.n23 14.0791
R3008 Delay_Cell_mag_0.OUTB.n25 Delay_Cell_mag_0.OUTB.n24 14.0791
R3009 Delay_Cell_mag_0.OUTB.n8 Delay_Cell_mag_0.OUTB.n7 14.0791
R3010 Delay_Cell_mag_0.OUTB.n1 Delay_Cell_mag_0.OUTB.n0 12.7222
R3011 Delay_Cell_mag_0.OUTB.n2 Delay_Cell_mag_0.OUTB.t23 11.6444
R3012 Delay_Cell_mag_0.OUTB.n2 Delay_Cell_mag_0.OUTB.n1 10.0261
R3013 Delay_Cell_mag_0.OUTB.n23 Delay_Cell_mag_0.OUTB.t24 8.213
R3014 Delay_Cell_mag_0.OUTB.n24 Delay_Cell_mag_0.OUTB.t16 8.213
R3015 Delay_Cell_mag_0.OUTB.n25 Delay_Cell_mag_0.OUTB.t19 8.213
R3016 Delay_Cell_mag_0.OUTB.n8 Delay_Cell_mag_0.OUTB.t8 8.08264
R3017 Delay_Cell_mag_0.OUTB.n7 Delay_Cell_mag_0.OUTB.t6 8.08264
R3018 Delay_Cell_mag_0.OUTB.n9 Delay_Cell_mag_0.OUTB.n8 7.03979
R3019 Delay_Cell_mag_0.OUTB.n0 Delay_Cell_mag_0.OUTB.t18 6.51836
R3020 Delay_Cell_mag_0.OUTB.n1 Delay_Cell_mag_0.OUTB.t20 6.51836
R3021 Delay_Cell_mag_0.OUTB.n17 Delay_Cell_mag_0.OUTB.n16 4.70398
R3022 Delay_Cell_mag_0.OUTB.n18 Delay_Cell_mag_0.OUTB.n17 4.4843
R3023 Delay_Cell_mag_0.OUTB.n10 Delay_Cell_mag_0.OUTB.n9 4.0005
R3024 Delay_Cell_mag_0.OUTB.n22 Delay_Cell_mag_0.OUTB.n21 3.3342
R3025 Delay_Cell_mag_0.OUTB.n17 Delay_Cell_mag_0.OUTB.n14 3.1505
R3026 Delay_Cell_mag_0.OUTB.n10 Delay_Cell_mag_0.OUTB.n6 2.94411
R3027 Delay_Cell_mag_0.OUTB.n22 Delay_Cell_mag_0.OUTB.n4 2.9292
R3028 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.OUTB.n25 2.70614
R3029 Delay_Cell_mag_0.OUTB.n18 Delay_Cell_mag_0.OUTB.n12 2.6005
R3030 Delay_Cell_mag_0.OUTB.n4 Delay_Cell_mag_0.OUTB.t13 1.8205
R3031 Delay_Cell_mag_0.OUTB.n4 Delay_Cell_mag_0.OUTB.n3 1.8205
R3032 Delay_Cell_mag_0.OUTB.n12 Delay_Cell_mag_0.OUTB.t12 1.8205
R3033 Delay_Cell_mag_0.OUTB.n12 Delay_Cell_mag_0.OUTB.n11 1.8205
R3034 Delay_Cell_mag_0.OUTB.n6 Delay_Cell_mag_0.OUTB.t5 1.8205
R3035 Delay_Cell_mag_0.OUTB.n6 Delay_Cell_mag_0.OUTB.n5 1.8205
R3036 Delay_Cell_mag_0.OUTB.n21 Delay_Cell_mag_0.OUTB.t7 1.8205
R3037 Delay_Cell_mag_0.OUTB.n21 Delay_Cell_mag_0.OUTB.n20 1.8205
R3038 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.OUTB.n2 1.77023
R3039 Delay_Cell_mag_0.OUTB.n14 Delay_Cell_mag_0.OUTB.t3 1.6385
R3040 Delay_Cell_mag_0.OUTB.n14 Delay_Cell_mag_0.OUTB.n13 1.6385
R3041 Delay_Cell_mag_0.OUTB.n16 Delay_Cell_mag_0.OUTB.t2 1.6385
R3042 Delay_Cell_mag_0.OUTB.n16 Delay_Cell_mag_0.OUTB.n15 1.6385
R3043 Delay_Cell_mag_0.OUTB.n22 Delay_Cell_mag_0.OUTB.n19 0.845717
R3044 Delay_Cell_mag_0.OUTB.n19 Delay_Cell_mag_0.OUTB.n10 0.335065
R3045 Delay_Cell_mag_0.OUTB.n19 Delay_Cell_mag_0.OUTB.n18 0.329196
R3046 VCONT.n0 VCONT.t12 21.8873
R3047 VCONT.n6 VCONT.t0 21.8873
R3048 VCONT.n3 VCONT.t6 21.8873
R3049 VCONT.n12 VCONT.t1 21.8873
R3050 VCONT.n1 VCONT.n0 12.5576
R3051 VCONT.n7 VCONT.n6 12.5576
R3052 VCONT.n4 VCONT.n3 12.5576
R3053 VCONT.n13 VCONT.n12 12.5576
R3054 VCONT.n2 VCONT.t10 12.1889
R3055 VCONT.n8 VCONT.t14 12.1889
R3056 VCONT.n5 VCONT.t11 12.1889
R3057 VCONT.n14 VCONT.t8 12.1889
R3058 VCONT.n2 VCONT.n1 9.69888
R3059 VCONT.n8 VCONT.n7 9.69888
R3060 VCONT.n5 VCONT.n4 9.69888
R3061 VCONT.n14 VCONT.n13 9.69888
R3062 VCONT.n10 VCONT 9.20341
R3063 VCONT.n9 VCONT 8.99233
R3064 VCONT.n0 VCONT.t2 6.51836
R3065 VCONT.n1 VCONT.t4 6.51836
R3066 VCONT.n6 VCONT.t15 6.51836
R3067 VCONT.n7 VCONT.t7 6.51836
R3068 VCONT.n3 VCONT.t3 6.51836
R3069 VCONT.n4 VCONT.t13 6.51836
R3070 VCONT.n12 VCONT.t5 6.51836
R3071 VCONT.n13 VCONT.t9 6.51836
R3072 VCONT.n9 VCONT 4.75244
R3073 VCONT VCONT.n2 4.63297
R3074 VCONT VCONT.n8 4.63297
R3075 VCONT VCONT.n5 4.63297
R3076 VCONT VCONT.n14 4.63297
R3077 VCONT.n11 VCONT.n10 4.5005
R3078 VCONT.n10 VCONT.n9 2.30392
R3079 VCONT.n11 VCONT 0.244813
R3080 VCONT VCONT.n11 0.0469095
R3081 a_8644_959.t0 a_8644_959.n5 22.8782
R3082 a_8644_959.n6 a_8644_959.t0 22.4219
R3083 a_8644_959.n3 a_8644_959.t16 22.2916
R3084 a_8644_959.n5 a_8644_959.n4 14.0791
R3085 a_8644_959.n4 a_8644_959.n3 14.0791
R3086 a_8644_959.n7 a_8644_959.n6 14.0791
R3087 a_8644_959.n2 a_8644_959.t2 11.3416
R3088 a_8644_959.n6 a_8644_959.t4 8.34336
R3089 a_8644_959.n7 a_8644_959.t6 8.34336
R3090 a_8644_959.n5 a_8644_959.t17 8.213
R3091 a_8644_959.n4 a_8644_959.t15 8.213
R3092 a_8644_959.n3 a_8644_959.t14 8.213
R3093 a_8644_959.n0 a_8644_959.n7 8.17193
R3094 a_8644_959.n1 a_8644_959.n2 4.0005
R3095 a_8644_959.n0 a_8644_959.n9 3.63045
R3096 a_8644_959.n18 a_8644_959.n1 2.89398
R3097 a_8644_959.n14 a_8644_959.n11 2.26392
R3098 a_8644_959.n9 a_8644_959.t1 1.8205
R3099 a_8644_959.n9 a_8644_959.n8 1.8205
R3100 a_8644_959.t7 a_8644_959.n18 1.8205
R3101 a_8644_959.n18 a_8644_959.n17 1.8205
R3102 a_8644_959.n11 a_8644_959.t10 1.6385
R3103 a_8644_959.n11 a_8644_959.n10 1.6385
R3104 a_8644_959.n13 a_8644_959.t9 1.6385
R3105 a_8644_959.n13 a_8644_959.n12 1.6385
R3106 a_8644_959.n2 a_8644_959.n16 1.62996
R3107 a_8644_959.n14 a_8644_959.n13 1.4936
R3108 a_8644_959.n1 a_8644_959.n15 1.22554
R3109 a_8644_959.n15 a_8644_959.n14 1.18673
R3110 a_8644_959.n1 a_8644_959.n0 0.1505
R3111 OUT.n9 OUT.n3 3.58485
R3112 OUT.n8 OUT.n7 3.58485
R3113 OUT.n9 OUT.n1 3.32833
R3114 OUT.n8 OUT.n5 3.32833
R3115 OUT.n3 OUT.t4 1.1705
R3116 OUT.n3 OUT.n2 1.1705
R3117 OUT.n7 OUT.t5 1.1705
R3118 OUT.n7 OUT.n6 1.1705
R3119 OUT.n9 OUT.n8 0.68137
R3120 OUT.n1 OUT.t2 0.6505
R3121 OUT.n1 OUT.n0 0.6505
R3122 OUT.n5 OUT.t3 0.6505
R3123 OUT.n5 OUT.n4 0.6505
R3124 OUT OUT.n9 0.297891
R3125 EN EN.n2 60.8984
R3126 EN EN.n3 60.8974
R3127 EN EN.n1 60.897
R3128 EN EN.n0 60.8619
R3129 EN.n0 EN.t5 22.6826
R3130 EN.n1 EN.t7 22.6826
R3131 EN.n2 EN.t3 22.6826
R3132 EN.n3 EN.t2 22.6826
R3133 EN.n4 EN 9.24918
R3134 EN.n5 EN 9.00634
R3135 EN.n0 EN.t1 8.60407
R3136 EN.n1 EN.t4 8.60407
R3137 EN.n2 EN.t0 8.60407
R3138 EN.n3 EN.t6 8.60407
R3139 EN.n6 EN.n5 4.72867
R3140 EN.n4 EN 4.52738
R3141 EN.n5 EN.n4 2.26677
R3142 EN.n6 EN 0.1555
R3143 EN EN.n6 0.0196667
C0 GF_INV16_2.IN Delay_Cell_mag_0.INB 8.2e-19
C1 Delay_Cell_mag_1.IN a_705_418# 0.337f
C2 a_510_2660# VCONT 7.89e-19
C3 GF_INV16_1.IN OUTB 0.273f
C4 Delay_Cell_mag_2.INB a_510_2660# 0.542f
C5 a_705_418# EN 0.497f
C6 VCONT OUTB 0.00171f
C7 a_705_418# VDD 0.154f
C8 Delay_Cell_mag_2.OUT Delay_Cell_mag_2.OUTB 2.47f
C9 Delay_Cell_mag_2.OUT Delay_Cell_mag_0.IN 1.85e-19
C10 GF_INV1_0.OUT OUT 2.76e-19
C11 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.IN 0.0384f
C12 Delay_Cell_mag_2.IN Delay_Cell_mag_2.OUT 0.379f
C13 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.OUT 1.6f
C14 Delay_Cell_mag_2.OUT a_705_n3320# 0.487f
C15 Delay_Cell_mag_2.OUTB a_510_n1078# 0.422f
C16 Delay_Cell_mag_2.IN a_510_n1078# 0.0324f
C17 GF_INV16_2.IN EN 0.178f
C18 Delay_Cell_mag_1.INB GF_INV1_0.OUT 0.156f
C19 Delay_Cell_mag_0.OUTB a_6953_n1078# 0.455f
C20 GF_INV16_2.IN VDD 1.89f
C21 Delay_Cell_mag_0.IN a_7148_n3320# 0.61f
C22 Delay_Cell_mag_2.OUTB Delay_Cell_mag_0.INB 0.0121f
C23 Delay_Cell_mag_0.INB Delay_Cell_mag_0.IN 0.899f
C24 Delay_Cell_mag_0.OUT a_7148_n3320# 0.487f
C25 VCONT OUT 0.00147f
C26 Delay_Cell_mag_0.OUT Delay_Cell_mag_0.INB 0.00336f
C27 Delay_Cell_mag_1.IN a_7148_419# 0.4f
C28 Delay_Cell_mag_2.OUT OUTB 7.36e-20
C29 a_7148_419# EN 0.202f
C30 a_7148_419# VDD 0.101f
C31 Delay_Cell_mag_1.IN a_6953_2661# 0.454f
C32 Delay_Cell_mag_1.INB GF_INV16_1.IN 5.46e-19
C33 Delay_Cell_mag_1.INB VCONT 0.317f
C34 a_6953_2661# EN 8.31e-20
C35 a_6953_2661# VDD 1.13f
C36 Delay_Cell_mag_2.INB Delay_Cell_mag_1.INB 0.00447f
C37 Delay_Cell_mag_1.IN Delay_Cell_mag_2.OUTB 0.00793f
C38 Delay_Cell_mag_1.IN Delay_Cell_mag_0.OUT 0.257f
C39 Delay_Cell_mag_2.OUTB EN 0.43f
C40 Delay_Cell_mag_2.OUTB VDD 5.03f
C41 Delay_Cell_mag_0.IN EN 0.279f
C42 Delay_Cell_mag_2.IN Delay_Cell_mag_1.IN 0.0362f
C43 Delay_Cell_mag_0.IN VDD 0.513f
C44 Delay_Cell_mag_0.OUT EN 0.0623f
C45 Delay_Cell_mag_0.OUT VDD 3.34f
C46 Delay_Cell_mag_2.IN EN 0.289f
C47 Delay_Cell_mag_2.IN VDD 4.54f
C48 a_705_n3320# EN 0.405f
C49 a_705_n3320# VDD 0.054f
C50 Delay_Cell_mag_0.OUTB OUT 0.00979f
C51 GF_INV1_0.OUT GF_INV16_1.IN 0.00101f
C52 GF_INV1_0.OUT VCONT 0.107f
C53 a_6953_n1078# EN 8.31e-20
C54 a_6953_n1078# VDD 1.13f
C55 Delay_Cell_mag_1.INB Delay_Cell_mag_2.OUT 6.54e-20
C56 Delay_Cell_mag_1.INB Delay_Cell_mag_0.OUTB 0.316f
C57 a_510_2660# EN 1.82e-19
C58 a_510_2660# VDD 1.12f
C59 Delay_Cell_mag_1.INB a_510_n1078# 1.77e-19
C60 GF_INV16_1.IN VCONT 0.0252f
C61 EN OUTB 0.00986f
C62 VDD OUTB 1.02f
C63 Delay_Cell_mag_2.INB VCONT 0.0215f
C64 GF_INV1_1.OUT OUTB 2.64e-19
C65 EN OUT 0.00949f
C66 VDD OUT 1.13f
C67 GF_INV16_2.IN a_7148_419# 7.82e-20
C68 a_705_418# Delay_Cell_mag_2.OUTB 5.63e-19
C69 GF_INV16_1.IN Delay_Cell_mag_2.OUT 0.00213f
C70 Delay_Cell_mag_2.OUT VCONT 0.0362f
C71 Delay_Cell_mag_1.IN Delay_Cell_mag_1.INB 3.11f
C72 Delay_Cell_mag_2.INB Delay_Cell_mag_2.OUT 0.00326f
C73 Delay_Cell_mag_0.OUTB VCONT 0.214f
C74 Delay_Cell_mag_2.IN a_705_418# 0.404f
C75 Delay_Cell_mag_1.INB EN 0.209f
C76 Delay_Cell_mag_1.INB VDD 4.09f
C77 a_510_n1078# VCONT 7.78e-19
C78 Delay_Cell_mag_2.INB a_510_n1078# 7.46e-19
C79 a_7148_n3320# VCONT 0.0688f
C80 GF_INV16_2.IN Delay_Cell_mag_0.OUT 1.68e-19
C81 Delay_Cell_mag_0.INB VCONT 0.159f
C82 GF_INV1_1.OUT Delay_Cell_mag_1.INB 0.00154f
C83 Delay_Cell_mag_1.IN GF_INV1_0.OUT 0.00842f
C84 GF_INV1_0.OUT EN 0.0349f
C85 GF_INV1_0.OUT VDD 1.16f
C86 a_7148_419# Delay_Cell_mag_0.OUT 0.324f
C87 Delay_Cell_mag_2.OUT Delay_Cell_mag_0.OUTB 3.07e-20
C88 Delay_Cell_mag_2.OUT a_510_n1078# 1.31f
C89 a_7148_419# a_6953_n1078# 0.00736f
C90 Delay_Cell_mag_1.IN GF_INV16_1.IN 0.252f
C91 Delay_Cell_mag_1.IN VCONT 0.359f
C92 GF_INV16_2.IN OUTB 2.26e-19
C93 GF_INV1_1.OUT GF_INV1_0.OUT 0.00589f
C94 Delay_Cell_mag_2.INB Delay_Cell_mag_1.IN 0.245f
C95 GF_INV16_1.IN EN 0.184f
C96 EN VCONT 1.24f
C97 Delay_Cell_mag_2.OUTB Delay_Cell_mag_0.IN 0.253f
C98 GF_INV16_1.IN VDD 1.6f
C99 VDD VCONT 1.96f
C100 Delay_Cell_mag_2.OUT Delay_Cell_mag_0.INB 0.256f
C101 Delay_Cell_mag_2.INB EN 0.233f
C102 Delay_Cell_mag_0.OUTB a_7148_n3320# 0.4f
C103 Delay_Cell_mag_0.OUT Delay_Cell_mag_0.IN 0.314f
C104 Delay_Cell_mag_2.INB VDD 3.16f
C105 Delay_Cell_mag_2.IN Delay_Cell_mag_2.OUTB 0.269f
C106 Delay_Cell_mag_0.OUTB Delay_Cell_mag_0.INB 0.266f
C107 Delay_Cell_mag_2.OUTB a_705_n3320# 0.4f
C108 Delay_Cell_mag_2.IN a_705_n3320# 0.679f
C109 Delay_Cell_mag_1.INB a_705_418# 0.37f
C110 Delay_Cell_mag_0.OUT a_6953_n1078# 0.699f
C111 GF_INV1_1.OUT GF_INV16_1.IN 0.219f
C112 GF_INV1_1.OUT VCONT 0.146f
C113 Delay_Cell_mag_0.INB a_7148_n3320# 0.354f
C114 GF_INV16_2.IN OUT 0.27f
C115 Delay_Cell_mag_1.IN Delay_Cell_mag_2.OUT 0.00529f
C116 Delay_Cell_mag_1.IN Delay_Cell_mag_0.OUTB 0.04f
C117 Delay_Cell_mag_2.OUT EN 0.3f
C118 Delay_Cell_mag_2.IN a_510_2660# 0.454f
C119 Delay_Cell_mag_2.OUT VDD 4.23f
C120 Delay_Cell_mag_0.OUTB EN 0.0662f
C121 Delay_Cell_mag_1.INB GF_INV16_2.IN 3.07e-19
C122 Delay_Cell_mag_0.OUTB VDD 3.64f
C123 Delay_Cell_mag_1.IN a_510_n1078# 0.0927f
C124 a_510_n1078# EN 0.0879f
C125 a_510_n1078# VDD 0.846f
C126 Delay_Cell_mag_1.INB a_7148_419# 0.487f
C127 a_7148_n3320# EN 0.201f
C128 a_7148_n3320# VDD 0.0541f
C129 Delay_Cell_mag_0.INB EN 0.11f
C130 Delay_Cell_mag_0.INB VDD 0.795f
C131 Delay_Cell_mag_1.INB a_6953_2661# 0.566f
C132 GF_INV1_0.OUT GF_INV16_2.IN 0.228f
C133 a_705_418# GF_INV16_1.IN 4.81e-20
C134 a_705_418# VCONT 0.035f
C135 Delay_Cell_mag_2.INB a_705_418# 0.499f
C136 Delay_Cell_mag_1.INB Delay_Cell_mag_2.OUTB 0.00334f
C137 Delay_Cell_mag_1.INB Delay_Cell_mag_0.OUT 0.00336f
C138 Delay_Cell_mag_2.IN Delay_Cell_mag_1.INB 0.266f
C139 Delay_Cell_mag_1.IN EN 0.275f
C140 Delay_Cell_mag_1.IN VDD 4.35f
C141 GF_INV16_1.IN GF_INV16_2.IN 0.0054f
C142 GF_INV16_2.IN VCONT 0.0245f
C143 VDD EN 1.11f
C144 a_705_418# Delay_Cell_mag_2.OUT 0.00249f
C145 a_7148_419# VCONT 0.155f
C146 a_510_2660# Delay_Cell_mag_1.INB 0.0406f
C147 Delay_Cell_mag_1.IN GF_INV1_1.OUT 0.348f
C148 a_6953_2661# VCONT 0.0055f
C149 GF_INV1_1.OUT EN 0.0419f
C150 GF_INV1_1.OUT VDD 0.888f
C151 a_705_418# a_510_n1078# 0.0321f
C152 GF_INV16_1.IN Delay_Cell_mag_2.OUTB 0.00108f
C153 GF_INV16_2.IN Delay_Cell_mag_2.OUT 3.48e-19
C154 Delay_Cell_mag_2.OUTB VCONT 0.167f
C155 Delay_Cell_mag_0.IN VCONT 0.0304f
C156 GF_INV16_2.IN Delay_Cell_mag_0.OUTB 0.0163f
C157 Delay_Cell_mag_2.INB Delay_Cell_mag_2.OUTB 0.263f
C158 Delay_Cell_mag_0.OUT VCONT 0.222f
C159 Delay_Cell_mag_2.IN GF_INV16_1.IN 7.74e-23
C160 Delay_Cell_mag_2.IN VCONT 0.0301f
C161 a_705_n3320# VCONT 0.0346f
C162 Delay_Cell_mag_2.INB Delay_Cell_mag_2.IN 3.03f
C163 Delay_Cell_mag_2.INB a_705_n3320# 0.347f
C164 a_6953_n1078# VCONT 0.104f
C165 a_7148_419# Delay_Cell_mag_0.OUTB 0.584f
.ends

