magic
tech gf180mcuC
magscale 1 10
timestamp 1692086575
<< error_p >>
rect -258 -23 -247 23
rect -34 -23 -23 23
rect 190 -23 201 23
<< pwell >>
rect -284 -100 284 100
<< nmos >>
rect -168 -28 -56 28
rect 56 -28 168 28
<< ndiff >>
rect -260 28 -188 36
rect -36 28 36 36
rect 188 28 260 36
rect -260 23 -168 28
rect -260 -23 -247 23
rect -201 -23 -168 23
rect -260 -28 -168 -23
rect -56 23 56 28
rect -56 -23 -23 23
rect 23 -23 56 23
rect -56 -28 56 -23
rect 168 23 260 28
rect 168 -23 201 23
rect 247 -23 260 23
rect 168 -28 260 -23
rect -260 -36 -188 -28
rect -36 -36 36 -28
rect 188 -36 260 -28
<< ndiffc >>
rect -247 -23 -201 23
rect -23 -23 23 23
rect 201 -23 247 23
<< polysilicon >>
rect -168 28 -56 72
rect 56 28 168 72
rect -168 -72 -56 -28
rect 56 -72 168 -28
<< metal1 >>
rect -258 -23 -247 23
rect -201 -23 -190 23
rect -34 -23 -23 23
rect 23 -23 34 23
rect 190 -23 201 23
rect 247 -23 258 23
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 0.28 l 0.56 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
