magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2045 -8202 2045 8202
<< psubdiff >>
rect -45 6180 45 6202
rect -45 -6180 -23 6180
rect 23 -6180 45 6180
rect -45 -6202 45 -6180
<< psubdiffcont >>
rect -23 -6180 23 6180
<< metal1 >>
rect -34 6180 34 6191
rect -34 -6180 -23 6180
rect 23 -6180 34 6180
rect -34 -6191 34 -6180
<< end >>
