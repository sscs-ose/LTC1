magic
tech gf180mcuC
magscale 1 10
timestamp 1693309239
<< psubdiff >>
rect -3951 2798 -3758 2822
rect -3951 2639 -3926 2798
rect -3782 2639 -3758 2798
rect -3951 2613 -3758 2639
rect -3701 2798 -3508 2822
rect -3701 2639 -3676 2798
rect -3532 2639 -3508 2798
rect -3701 2613 -3508 2639
rect -3451 2798 -3258 2822
rect -3451 2639 -3426 2798
rect -3282 2639 -3258 2798
rect -3451 2613 -3258 2639
rect -3201 2798 -3008 2822
rect -3201 2639 -3176 2798
rect -3032 2639 -3008 2798
rect -3201 2613 -3008 2639
rect -2951 2798 -2758 2822
rect -2951 2639 -2926 2798
rect -2782 2639 -2758 2798
rect -2951 2613 -2758 2639
rect -2701 2798 -2508 2822
rect -2701 2639 -2676 2798
rect -2532 2639 -2508 2798
rect -2701 2613 -2508 2639
rect -2451 2798 -2258 2822
rect -2451 2639 -2426 2798
rect -2282 2639 -2258 2798
rect -2451 2613 -2258 2639
rect -2201 2798 -2008 2822
rect -2201 2639 -2176 2798
rect -2032 2639 -2008 2798
rect -2201 2613 -2008 2639
rect -1951 2798 -1758 2822
rect -1951 2639 -1926 2798
rect -1782 2639 -1758 2798
rect -1951 2613 -1758 2639
rect -1701 2798 -1508 2822
rect -1701 2639 -1676 2798
rect -1532 2639 -1508 2798
rect -1701 2613 -1508 2639
rect -1451 2798 -1258 2822
rect -1451 2639 -1426 2798
rect -1282 2639 -1258 2798
rect -1451 2613 -1258 2639
rect -1201 2798 -1008 2822
rect -1201 2639 -1176 2798
rect -1032 2639 -1008 2798
rect -1201 2613 -1008 2639
rect -951 2798 -758 2822
rect -951 2639 -926 2798
rect -782 2639 -758 2798
rect -951 2613 -758 2639
rect -701 2798 -508 2822
rect -701 2639 -676 2798
rect -532 2639 -508 2798
rect -701 2613 -508 2639
rect -451 2798 -258 2822
rect -451 2639 -426 2798
rect -282 2639 -258 2798
rect -451 2613 -258 2639
rect -201 2798 -8 2822
rect -201 2639 -176 2798
rect -32 2639 -8 2798
rect -201 2613 -8 2639
rect 49 2798 242 2822
rect 49 2639 74 2798
rect 218 2639 242 2798
rect 49 2613 242 2639
rect 299 2798 492 2822
rect 299 2639 324 2798
rect 468 2639 492 2798
rect 299 2613 492 2639
rect 549 2798 742 2822
rect 549 2639 574 2798
rect 718 2639 742 2798
rect 549 2613 742 2639
rect 799 2798 992 2822
rect 799 2639 824 2798
rect 968 2639 992 2798
rect 799 2613 992 2639
rect 1049 2798 1242 2822
rect 1049 2639 1074 2798
rect 1218 2639 1242 2798
rect 1049 2613 1242 2639
rect 1299 2798 1492 2822
rect 1299 2639 1324 2798
rect 1468 2639 1492 2798
rect 1299 2613 1492 2639
rect 1549 2798 1742 2822
rect 1549 2639 1574 2798
rect 1718 2639 1742 2798
rect 1549 2613 1742 2639
rect 1799 2798 1992 2822
rect 1799 2639 1824 2798
rect 1968 2639 1992 2798
rect 1799 2613 1992 2639
rect 2049 2798 2242 2822
rect 2049 2639 2074 2798
rect 2218 2639 2242 2798
rect 2049 2613 2242 2639
rect 2299 2798 2492 2822
rect 2299 2639 2324 2798
rect 2468 2639 2492 2798
rect 2299 2613 2492 2639
rect 2549 2798 2742 2822
rect 2549 2639 2574 2798
rect 2718 2639 2742 2798
rect 2549 2613 2742 2639
rect 2799 2798 2992 2822
rect 2799 2639 2824 2798
rect 2968 2639 2992 2798
rect 2799 2613 2992 2639
rect 3049 2798 3242 2822
rect 3049 2639 3074 2798
rect 3218 2639 3242 2798
rect 3049 2613 3242 2639
rect 3299 2798 3492 2822
rect 3299 2639 3324 2798
rect 3468 2639 3492 2798
rect 3299 2613 3492 2639
rect 3549 2798 3742 2822
rect 3549 2639 3574 2798
rect 3718 2639 3742 2798
rect 3549 2613 3742 2639
rect 3799 2798 3992 2822
rect 3799 2639 3824 2798
rect 3968 2639 3992 2798
rect 3799 2613 3992 2639
rect 4049 2798 4242 2822
rect 4049 2639 4074 2798
rect 4218 2639 4242 2798
rect 4049 2613 4242 2639
rect 4299 2798 4492 2822
rect 4299 2639 4324 2798
rect 4468 2639 4492 2798
rect 4299 2613 4492 2639
rect 4549 2798 4742 2822
rect 4549 2639 4574 2798
rect 4718 2639 4742 2798
rect 4549 2613 4742 2639
rect 4799 2798 4992 2822
rect 4799 2639 4824 2798
rect 4968 2639 4992 2798
rect 4799 2613 4992 2639
rect 5049 2798 5242 2822
rect 5049 2639 5074 2798
rect 5218 2639 5242 2798
rect 5049 2613 5242 2639
rect 5299 2798 5492 2822
rect 5299 2639 5324 2798
rect 5468 2639 5492 2798
rect 5299 2613 5492 2639
rect 5549 2798 5742 2822
rect 5549 2639 5574 2798
rect 5718 2639 5742 2798
rect 5549 2613 5742 2639
rect 5799 2798 5992 2822
rect 5799 2639 5824 2798
rect 5968 2639 5992 2798
rect 5799 2613 5992 2639
rect 6049 2798 6242 2822
rect 6049 2639 6074 2798
rect 6218 2639 6242 2798
rect 6049 2613 6242 2639
rect 6299 2798 6492 2822
rect 6299 2639 6324 2798
rect 6468 2639 6492 2798
rect 6299 2613 6492 2639
rect 6549 2798 6742 2822
rect 6549 2639 6574 2798
rect 6718 2639 6742 2798
rect 6549 2613 6742 2639
rect 6799 2798 6992 2822
rect 6799 2639 6824 2798
rect 6968 2639 6992 2798
rect 6799 2613 6992 2639
rect -3951 1693 -3758 1717
rect -3951 1534 -3926 1693
rect -3782 1534 -3758 1693
rect -3951 1508 -3758 1534
rect -3701 1693 -3508 1717
rect -3701 1534 -3676 1693
rect -3532 1534 -3508 1693
rect -3701 1508 -3508 1534
rect -3451 1693 -3258 1717
rect -3451 1534 -3426 1693
rect -3282 1534 -3258 1693
rect -3451 1508 -3258 1534
rect -3201 1693 -3008 1717
rect -3201 1534 -3176 1693
rect -3032 1534 -3008 1693
rect -3201 1508 -3008 1534
rect -2951 1693 -2758 1717
rect -2951 1534 -2926 1693
rect -2782 1534 -2758 1693
rect -2951 1508 -2758 1534
rect -2701 1693 -2508 1717
rect -2701 1534 -2676 1693
rect -2532 1534 -2508 1693
rect -2701 1508 -2508 1534
rect -2451 1693 -2258 1717
rect -2451 1534 -2426 1693
rect -2282 1534 -2258 1693
rect -2451 1508 -2258 1534
rect -2201 1693 -2008 1717
rect -2201 1534 -2176 1693
rect -2032 1534 -2008 1693
rect -2201 1508 -2008 1534
rect -1951 1693 -1758 1717
rect -1951 1534 -1926 1693
rect -1782 1534 -1758 1693
rect -1951 1508 -1758 1534
rect -1701 1693 -1508 1717
rect -1701 1534 -1676 1693
rect -1532 1534 -1508 1693
rect -1701 1508 -1508 1534
rect -1451 1693 -1258 1717
rect -1451 1534 -1426 1693
rect -1282 1534 -1258 1693
rect -1451 1508 -1258 1534
rect -1201 1693 -1008 1717
rect -1201 1534 -1176 1693
rect -1032 1534 -1008 1693
rect -1201 1508 -1008 1534
rect -951 1693 -758 1717
rect -951 1534 -926 1693
rect -782 1534 -758 1693
rect -951 1508 -758 1534
rect -701 1693 -508 1717
rect -701 1534 -676 1693
rect -532 1534 -508 1693
rect -701 1508 -508 1534
rect -451 1693 -258 1717
rect -451 1534 -426 1693
rect -282 1534 -258 1693
rect -451 1508 -258 1534
rect -201 1693 -8 1717
rect -201 1534 -176 1693
rect -32 1534 -8 1693
rect -201 1508 -8 1534
rect 49 1693 242 1717
rect 49 1534 74 1693
rect 218 1534 242 1693
rect 49 1508 242 1534
rect 299 1693 492 1717
rect 299 1534 324 1693
rect 468 1534 492 1693
rect 299 1508 492 1534
rect 549 1693 742 1717
rect 549 1534 574 1693
rect 718 1534 742 1693
rect 549 1508 742 1534
rect 799 1693 992 1717
rect 799 1534 824 1693
rect 968 1534 992 1693
rect 799 1508 992 1534
rect 1049 1693 1242 1717
rect 1049 1534 1074 1693
rect 1218 1534 1242 1693
rect 1049 1508 1242 1534
rect 1299 1693 1492 1717
rect 1299 1534 1324 1693
rect 1468 1534 1492 1693
rect 1299 1508 1492 1534
rect 1549 1693 1742 1717
rect 1549 1534 1574 1693
rect 1718 1534 1742 1693
rect 1549 1508 1742 1534
rect 1799 1693 1992 1717
rect 1799 1534 1824 1693
rect 1968 1534 1992 1693
rect 1799 1508 1992 1534
rect 2049 1693 2242 1717
rect 2049 1534 2074 1693
rect 2218 1534 2242 1693
rect 2049 1508 2242 1534
rect 2299 1693 2492 1717
rect 2299 1534 2324 1693
rect 2468 1534 2492 1693
rect 2299 1508 2492 1534
rect 2549 1693 2742 1717
rect 2549 1534 2574 1693
rect 2718 1534 2742 1693
rect 2549 1508 2742 1534
rect 2799 1693 2992 1717
rect 2799 1534 2824 1693
rect 2968 1534 2992 1693
rect 2799 1508 2992 1534
rect 3049 1693 3242 1717
rect 3049 1534 3074 1693
rect 3218 1534 3242 1693
rect 3049 1508 3242 1534
rect 3299 1693 3492 1717
rect 3299 1534 3324 1693
rect 3468 1534 3492 1693
rect 3299 1508 3492 1534
rect 3549 1693 3742 1717
rect 3549 1534 3574 1693
rect 3718 1534 3742 1693
rect 3549 1508 3742 1534
rect 3799 1693 3992 1717
rect 3799 1534 3824 1693
rect 3968 1534 3992 1693
rect 3799 1508 3992 1534
rect 4049 1693 4242 1717
rect 4049 1534 4074 1693
rect 4218 1534 4242 1693
rect 4049 1508 4242 1534
rect 4299 1693 4492 1717
rect 4299 1534 4324 1693
rect 4468 1534 4492 1693
rect 4299 1508 4492 1534
rect 4549 1693 4742 1717
rect 4549 1534 4574 1693
rect 4718 1534 4742 1693
rect 4549 1508 4742 1534
rect 4799 1693 4992 1717
rect 4799 1534 4824 1693
rect 4968 1534 4992 1693
rect 4799 1508 4992 1534
rect 5049 1693 5242 1717
rect 5049 1534 5074 1693
rect 5218 1534 5242 1693
rect 5049 1508 5242 1534
rect 5299 1693 5492 1717
rect 5299 1534 5324 1693
rect 5468 1534 5492 1693
rect 5299 1508 5492 1534
rect 5549 1693 5742 1717
rect 5549 1534 5574 1693
rect 5718 1534 5742 1693
rect 5549 1508 5742 1534
rect 5799 1693 5992 1717
rect 5799 1534 5824 1693
rect 5968 1534 5992 1693
rect 5799 1508 5992 1534
rect 6049 1693 6242 1717
rect 6049 1534 6074 1693
rect 6218 1534 6242 1693
rect 6049 1508 6242 1534
rect 6299 1693 6492 1717
rect 6299 1534 6324 1693
rect 6468 1534 6492 1693
rect 6299 1508 6492 1534
rect 6549 1693 6742 1717
rect 6549 1534 6574 1693
rect 6718 1534 6742 1693
rect 6549 1508 6742 1534
rect 6799 1693 6992 1717
rect 6799 1534 6824 1693
rect 6968 1534 6992 1693
rect 6799 1508 6992 1534
rect -3969 568 -3776 592
rect -3969 409 -3944 568
rect -3800 409 -3776 568
rect -3969 383 -3776 409
rect -3719 568 -3526 592
rect -3719 409 -3694 568
rect -3550 409 -3526 568
rect -3719 383 -3526 409
rect -3469 568 -3276 592
rect -3469 409 -3444 568
rect -3300 409 -3276 568
rect -3469 383 -3276 409
rect -3219 568 -3026 592
rect -3219 409 -3194 568
rect -3050 409 -3026 568
rect -3219 383 -3026 409
rect -2969 568 -2776 592
rect -2969 409 -2944 568
rect -2800 409 -2776 568
rect -2969 383 -2776 409
rect -2719 568 -2526 592
rect -2719 409 -2694 568
rect -2550 409 -2526 568
rect -2719 383 -2526 409
rect -2469 568 -2276 592
rect -2469 409 -2444 568
rect -2300 409 -2276 568
rect -2469 383 -2276 409
rect -2219 568 -2026 592
rect -2219 409 -2194 568
rect -2050 409 -2026 568
rect -2219 383 -2026 409
rect -1969 568 -1776 592
rect -1969 409 -1944 568
rect -1800 409 -1776 568
rect -1969 383 -1776 409
rect -1719 568 -1526 592
rect -1719 409 -1694 568
rect -1550 409 -1526 568
rect -1719 383 -1526 409
rect -1469 568 -1276 592
rect -1469 409 -1444 568
rect -1300 409 -1276 568
rect -1469 383 -1276 409
rect -1219 568 -1026 592
rect -1219 409 -1194 568
rect -1050 409 -1026 568
rect -1219 383 -1026 409
rect -969 568 -776 592
rect -969 409 -944 568
rect -800 409 -776 568
rect -969 383 -776 409
rect -719 568 -526 592
rect -719 409 -694 568
rect -550 409 -526 568
rect -719 383 -526 409
rect -469 568 -276 592
rect -469 409 -444 568
rect -300 409 -276 568
rect -469 383 -276 409
rect -219 568 -26 592
rect -219 409 -194 568
rect -50 409 -26 568
rect -219 383 -26 409
rect 31 568 224 592
rect 31 409 56 568
rect 200 409 224 568
rect 31 383 224 409
rect 281 568 474 592
rect 281 409 306 568
rect 450 409 474 568
rect 281 383 474 409
rect 531 568 724 592
rect 531 409 556 568
rect 700 409 724 568
rect 531 383 724 409
rect 781 568 974 592
rect 781 409 806 568
rect 950 409 974 568
rect 781 383 974 409
rect 1031 568 1224 592
rect 1031 409 1056 568
rect 1200 409 1224 568
rect 1031 383 1224 409
rect 1281 568 1474 592
rect 1281 409 1306 568
rect 1450 409 1474 568
rect 1281 383 1474 409
rect 1531 568 1724 592
rect 1531 409 1556 568
rect 1700 409 1724 568
rect 1531 383 1724 409
rect 1781 568 1974 592
rect 1781 409 1806 568
rect 1950 409 1974 568
rect 1781 383 1974 409
rect 2031 568 2224 592
rect 2031 409 2056 568
rect 2200 409 2224 568
rect 2031 383 2224 409
rect 2281 568 2474 592
rect 2281 409 2306 568
rect 2450 409 2474 568
rect 2281 383 2474 409
rect 2531 568 2724 592
rect 2531 409 2556 568
rect 2700 409 2724 568
rect 2531 383 2724 409
rect 2781 568 2974 592
rect 2781 409 2806 568
rect 2950 409 2974 568
rect 2781 383 2974 409
rect 3031 568 3224 592
rect 3031 409 3056 568
rect 3200 409 3224 568
rect 3031 383 3224 409
rect 3281 568 3474 592
rect 3281 409 3306 568
rect 3450 409 3474 568
rect 3281 383 3474 409
rect 3531 568 3724 592
rect 3531 409 3556 568
rect 3700 409 3724 568
rect 3531 383 3724 409
rect 3781 568 3974 592
rect 3781 409 3806 568
rect 3950 409 3974 568
rect 3781 383 3974 409
rect 4031 568 4224 592
rect 4031 409 4056 568
rect 4200 409 4224 568
rect 4031 383 4224 409
rect 4281 568 4474 592
rect 4281 409 4306 568
rect 4450 409 4474 568
rect 4281 383 4474 409
rect 4531 568 4724 592
rect 4531 409 4556 568
rect 4700 409 4724 568
rect 4531 383 4724 409
rect 4781 568 4974 592
rect 4781 409 4806 568
rect 4950 409 4974 568
rect 4781 383 4974 409
rect 5031 568 5224 592
rect 5031 409 5056 568
rect 5200 409 5224 568
rect 5031 383 5224 409
rect 5281 568 5474 592
rect 5281 409 5306 568
rect 5450 409 5474 568
rect 5281 383 5474 409
rect 5531 568 5724 592
rect 5531 409 5556 568
rect 5700 409 5724 568
rect 5531 383 5724 409
rect 5781 568 5974 592
rect 5781 409 5806 568
rect 5950 409 5974 568
rect 5781 383 5974 409
rect 6031 568 6224 592
rect 6031 409 6056 568
rect 6200 409 6224 568
rect 6031 383 6224 409
rect 6281 568 6474 592
rect 6281 409 6306 568
rect 6450 409 6474 568
rect 6281 383 6474 409
rect 6531 568 6724 592
rect 6531 409 6556 568
rect 6700 409 6724 568
rect 6531 383 6724 409
rect 6781 568 6974 592
rect 6781 409 6806 568
rect 6950 409 6974 568
rect 6781 383 6974 409
<< psubdiffcont >>
rect -3926 2639 -3782 2798
rect -3676 2639 -3532 2798
rect -3426 2639 -3282 2798
rect -3176 2639 -3032 2798
rect -2926 2639 -2782 2798
rect -2676 2639 -2532 2798
rect -2426 2639 -2282 2798
rect -2176 2639 -2032 2798
rect -1926 2639 -1782 2798
rect -1676 2639 -1532 2798
rect -1426 2639 -1282 2798
rect -1176 2639 -1032 2798
rect -926 2639 -782 2798
rect -676 2639 -532 2798
rect -426 2639 -282 2798
rect -176 2639 -32 2798
rect 74 2639 218 2798
rect 324 2639 468 2798
rect 574 2639 718 2798
rect 824 2639 968 2798
rect 1074 2639 1218 2798
rect 1324 2639 1468 2798
rect 1574 2639 1718 2798
rect 1824 2639 1968 2798
rect 2074 2639 2218 2798
rect 2324 2639 2468 2798
rect 2574 2639 2718 2798
rect 2824 2639 2968 2798
rect 3074 2639 3218 2798
rect 3324 2639 3468 2798
rect 3574 2639 3718 2798
rect 3824 2639 3968 2798
rect 4074 2639 4218 2798
rect 4324 2639 4468 2798
rect 4574 2639 4718 2798
rect 4824 2639 4968 2798
rect 5074 2639 5218 2798
rect 5324 2639 5468 2798
rect 5574 2639 5718 2798
rect 5824 2639 5968 2798
rect 6074 2639 6218 2798
rect 6324 2639 6468 2798
rect 6574 2639 6718 2798
rect 6824 2639 6968 2798
rect -3926 1534 -3782 1693
rect -3676 1534 -3532 1693
rect -3426 1534 -3282 1693
rect -3176 1534 -3032 1693
rect -2926 1534 -2782 1693
rect -2676 1534 -2532 1693
rect -2426 1534 -2282 1693
rect -2176 1534 -2032 1693
rect -1926 1534 -1782 1693
rect -1676 1534 -1532 1693
rect -1426 1534 -1282 1693
rect -1176 1534 -1032 1693
rect -926 1534 -782 1693
rect -676 1534 -532 1693
rect -426 1534 -282 1693
rect -176 1534 -32 1693
rect 74 1534 218 1693
rect 324 1534 468 1693
rect 574 1534 718 1693
rect 824 1534 968 1693
rect 1074 1534 1218 1693
rect 1324 1534 1468 1693
rect 1574 1534 1718 1693
rect 1824 1534 1968 1693
rect 2074 1534 2218 1693
rect 2324 1534 2468 1693
rect 2574 1534 2718 1693
rect 2824 1534 2968 1693
rect 3074 1534 3218 1693
rect 3324 1534 3468 1693
rect 3574 1534 3718 1693
rect 3824 1534 3968 1693
rect 4074 1534 4218 1693
rect 4324 1534 4468 1693
rect 4574 1534 4718 1693
rect 4824 1534 4968 1693
rect 5074 1534 5218 1693
rect 5324 1534 5468 1693
rect 5574 1534 5718 1693
rect 5824 1534 5968 1693
rect 6074 1534 6218 1693
rect 6324 1534 6468 1693
rect 6574 1534 6718 1693
rect 6824 1534 6968 1693
rect -3944 409 -3800 568
rect -3694 409 -3550 568
rect -3444 409 -3300 568
rect -3194 409 -3050 568
rect -2944 409 -2800 568
rect -2694 409 -2550 568
rect -2444 409 -2300 568
rect -2194 409 -2050 568
rect -1944 409 -1800 568
rect -1694 409 -1550 568
rect -1444 409 -1300 568
rect -1194 409 -1050 568
rect -944 409 -800 568
rect -694 409 -550 568
rect -444 409 -300 568
rect -194 409 -50 568
rect 56 409 200 568
rect 306 409 450 568
rect 556 409 700 568
rect 806 409 950 568
rect 1056 409 1200 568
rect 1306 409 1450 568
rect 1556 409 1700 568
rect 1806 409 1950 568
rect 2056 409 2200 568
rect 2306 409 2450 568
rect 2556 409 2700 568
rect 2806 409 2950 568
rect 3056 409 3200 568
rect 3306 409 3450 568
rect 3556 409 3700 568
rect 3806 409 3950 568
rect 4056 409 4200 568
rect 4306 409 4450 568
rect 4556 409 4700 568
rect 4806 409 4950 568
rect 5056 409 5200 568
rect 5306 409 5450 568
rect 5556 409 5700 568
rect 5806 409 5950 568
rect 6056 409 6200 568
rect 6306 409 6450 568
rect 6556 409 6700 568
rect 6806 409 6950 568
<< polysilicon >>
rect -4148 2545 7026 2565
rect -4148 2491 -4135 2545
rect -4077 2525 7026 2545
rect -4077 2502 -3638 2525
rect -4077 2491 -4062 2502
rect -4148 2477 -4062 2491
rect -3878 2464 -3638 2502
rect -2846 2464 -2606 2525
rect -2502 2464 -2262 2525
rect -1470 2464 -1230 2525
rect -1126 2464 -886 2525
rect -94 2464 146 2525
rect 250 2464 490 2525
rect 1282 2464 1522 2525
rect 1626 2464 1866 2525
rect 2658 2464 2898 2525
rect 3002 2464 3242 2525
rect 4034 2464 4274 2525
rect 4378 2464 4618 2525
rect 5410 2464 5650 2525
rect 5754 2464 5994 2525
rect 6786 2464 7026 2525
rect -4090 2194 -4010 2210
rect -4090 2141 -4076 2194
rect -4026 2187 -4010 2194
rect -3534 2187 -3294 2256
rect -3190 2187 -2950 2256
rect -2158 2187 -1918 2256
rect -1814 2187 -1574 2256
rect -782 2187 -542 2256
rect -438 2187 -198 2256
rect 594 2187 834 2256
rect 938 2187 1178 2256
rect 1970 2187 2210 2256
rect 2314 2187 2554 2256
rect 3346 2187 3586 2256
rect 3690 2187 3930 2256
rect 4722 2187 4962 2256
rect 5066 2187 5306 2256
rect 6098 2187 6338 2256
rect 6442 2187 6682 2256
rect -4026 2147 7026 2187
rect -4026 2141 -4010 2147
rect -4090 2125 -4010 2141
rect -3878 2097 -3638 2147
rect -2846 2097 -2606 2147
rect -2502 2097 -2262 2147
rect -1470 2097 -1230 2147
rect -1126 2097 -886 2147
rect -94 2097 146 2147
rect 250 2097 490 2147
rect 1282 2097 1522 2147
rect 1626 2097 1866 2147
rect 2658 2097 2898 2147
rect 3002 2097 3242 2147
rect 4034 2097 4274 2147
rect 4378 2097 4618 2147
rect 5410 2097 5650 2147
rect 5754 2097 5994 2147
rect 6786 2097 7026 2147
rect -4136 1828 -4060 1841
rect -4136 1776 -4123 1828
rect -4074 1822 -4060 1828
rect -3534 1822 -3294 1933
rect -3190 1822 -2950 1889
rect -2158 1822 -1918 1889
rect -1814 1822 -1574 1889
rect -782 1822 -542 1889
rect -438 1822 -198 1889
rect 594 1822 834 1889
rect 938 1822 1178 1889
rect 1970 1822 2210 1889
rect 2314 1822 2554 1889
rect 3346 1822 3586 1889
rect 3690 1822 3930 1889
rect 4722 1822 4962 1889
rect 5066 1822 5306 1889
rect 6098 1822 6338 1889
rect 6442 1822 6682 1889
rect -4074 1782 6682 1822
rect -4074 1776 -4060 1782
rect -4136 1763 -4060 1776
rect -4075 1455 7026 1460
rect -4149 1440 7026 1455
rect -4149 1386 -4135 1440
rect -4077 1420 7026 1440
rect -4077 1397 -3638 1420
rect -4077 1386 -4062 1397
rect -4149 1372 -4062 1386
rect -3878 1359 -3638 1397
rect -2846 1359 -2606 1420
rect -2502 1359 -2262 1420
rect -1470 1359 -1230 1420
rect -1126 1359 -886 1420
rect -94 1359 146 1420
rect 250 1359 490 1420
rect 1282 1359 1522 1420
rect 1626 1359 1866 1420
rect 2658 1359 2898 1420
rect 3002 1359 3242 1420
rect 4034 1359 4274 1420
rect 4378 1359 4618 1420
rect 5410 1359 5650 1420
rect 5754 1359 5994 1420
rect 6786 1359 7026 1420
rect -4104 1089 -4025 1106
rect -4104 1036 -4090 1089
rect -4038 1082 -4025 1089
rect -3534 1082 -3294 1151
rect -3190 1082 -2950 1151
rect -2158 1082 -1918 1151
rect -1814 1082 -1574 1151
rect -782 1082 -542 1151
rect -438 1082 -198 1151
rect 594 1082 834 1151
rect 938 1082 1178 1151
rect 1970 1082 2210 1151
rect 2314 1082 2554 1151
rect 3346 1082 3586 1151
rect 3690 1082 3930 1151
rect 4722 1082 4962 1151
rect 5066 1082 5306 1151
rect 6098 1082 6338 1151
rect 6442 1082 6682 1151
rect -4038 1042 7026 1082
rect -4038 1036 -4025 1042
rect -4104 1021 -4025 1036
rect -3878 992 -3638 1042
rect -2846 992 -2606 1042
rect -2502 992 -2262 1042
rect -1470 992 -1230 1042
rect -1126 992 -886 1042
rect -94 992 146 1042
rect 250 992 490 1042
rect 1282 992 1522 1042
rect 1626 992 1866 1042
rect 2658 992 2898 1042
rect 3002 992 3242 1042
rect 4034 992 4274 1042
rect 4378 992 4618 1042
rect 5410 992 5650 1042
rect 5754 992 5994 1042
rect 6786 992 7026 1042
rect -4136 723 -4060 736
rect -4136 671 -4123 723
rect -4074 717 -4060 723
rect -3534 717 -3294 828
rect -3190 717 -2950 784
rect -2158 717 -1918 784
rect -1814 717 -1574 784
rect -782 717 -542 784
rect -438 717 -198 784
rect 594 717 834 784
rect 938 717 1178 784
rect 1970 717 2210 784
rect 2314 717 2554 784
rect 3346 717 3586 784
rect 3690 717 3930 784
rect 4722 717 4962 784
rect 5066 717 5306 784
rect 6098 717 6338 784
rect 6442 717 6682 784
rect -4074 677 6682 717
rect -4074 671 -4060 677
rect -4136 658 -4060 671
<< polycontact >>
rect -4135 2491 -4077 2545
rect -4076 2141 -4026 2194
rect -4123 1776 -4074 1828
rect -4135 1386 -4077 1440
rect -4090 1036 -4038 1089
rect -4123 671 -4074 723
<< metal1 >>
rect -3991 2798 7115 2856
rect -3991 2639 -3926 2798
rect -3782 2639 -3676 2798
rect -3532 2639 -3426 2798
rect -3282 2639 -3176 2798
rect -3032 2639 -2926 2798
rect -2782 2639 -2676 2798
rect -2532 2639 -2426 2798
rect -2282 2639 -2176 2798
rect -2032 2639 -1926 2798
rect -1782 2639 -1676 2798
rect -1532 2639 -1426 2798
rect -1282 2639 -1176 2798
rect -1032 2639 -926 2798
rect -782 2639 -676 2798
rect -532 2639 -426 2798
rect -282 2639 -176 2798
rect -32 2639 74 2798
rect 218 2639 324 2798
rect 468 2639 574 2798
rect 718 2639 824 2798
rect 968 2639 1074 2798
rect 1218 2639 1324 2798
rect 1468 2639 1574 2798
rect 1718 2639 1824 2798
rect 1968 2639 2074 2798
rect 2218 2639 2324 2798
rect 2468 2639 2574 2798
rect 2718 2639 2824 2798
rect 2968 2639 3074 2798
rect 3218 2639 3324 2798
rect 3468 2639 3574 2798
rect 3718 2639 3824 2798
rect 3968 2639 4074 2798
rect 4218 2639 4324 2798
rect 4468 2639 4574 2798
rect 4718 2639 4824 2798
rect 4968 2639 5074 2798
rect 5218 2639 5324 2798
rect 5468 2639 5574 2798
rect 5718 2639 5824 2798
rect 5968 2639 6074 2798
rect 6218 2639 6324 2798
rect 6468 2639 6574 2798
rect 6718 2639 6824 2798
rect 6968 2795 7115 2798
rect 6968 2781 7113 2795
rect 6968 2779 7037 2781
rect 6985 2725 7037 2779
rect 7093 2725 7113 2781
rect 6968 2664 7113 2725
rect 6968 2661 7038 2664
rect -3991 2605 6930 2639
rect 6986 2610 7038 2661
rect 7092 2610 7113 2664
rect 6986 2605 7113 2610
rect -3991 2573 7113 2605
rect -4148 2546 -4062 2560
rect -4148 2489 -4137 2546
rect -4076 2489 -4062 2546
rect -4148 2477 -4062 2489
rect -3265 2418 -3219 2573
rect -1889 2418 -1843 2573
rect -513 2418 -467 2573
rect 863 2418 909 2573
rect 2239 2418 2285 2573
rect 3615 2418 3661 2573
rect 4991 2418 5037 2573
rect 6367 2418 6413 2573
rect -3622 2399 -3545 2408
rect -3622 2338 -3612 2399
rect -3556 2338 -3545 2399
rect -3622 2328 -3545 2338
rect -2941 2402 -2864 2411
rect -2941 2342 -2931 2402
rect -2875 2342 -2864 2402
rect -2941 2332 -2864 2342
rect -2259 2397 -2182 2406
rect -2259 2337 -2249 2397
rect -2193 2337 -2182 2397
rect -2259 2327 -2182 2337
rect -1568 2390 -1491 2399
rect -1568 2330 -1558 2390
rect -1502 2330 -1491 2390
rect -1568 2320 -1491 2330
rect -879 2389 -802 2398
rect -879 2329 -869 2389
rect -813 2329 -802 2389
rect -879 2319 -802 2329
rect -187 2389 -110 2398
rect -187 2329 -177 2389
rect -121 2329 -110 2389
rect -187 2319 -110 2329
rect 502 2389 579 2398
rect 502 2329 512 2389
rect 568 2329 579 2389
rect 502 2319 579 2329
rect 1192 2393 1269 2402
rect 1192 2333 1202 2393
rect 1258 2333 1269 2393
rect 1192 2323 1269 2333
rect 1878 2394 1955 2403
rect 1878 2334 1888 2394
rect 1944 2334 1955 2394
rect 1878 2324 1955 2334
rect 2565 2395 2642 2404
rect 2565 2335 2575 2395
rect 2631 2335 2642 2395
rect 2565 2325 2642 2335
rect 3254 2392 3331 2401
rect 3254 2332 3264 2392
rect 3320 2332 3331 2392
rect 3254 2322 3331 2332
rect 3949 2396 4026 2405
rect 3949 2336 3959 2396
rect 4015 2336 4026 2396
rect 3949 2326 4026 2336
rect 4629 2397 4706 2406
rect 4629 2337 4639 2397
rect 4695 2337 4706 2397
rect 4629 2327 4706 2337
rect 5315 2394 5392 2403
rect 5315 2334 5325 2394
rect 5381 2334 5392 2394
rect 5315 2324 5392 2334
rect 6004 2390 6081 2399
rect 6004 2330 6014 2390
rect 6070 2330 6081 2390
rect 6004 2320 6081 2330
rect 6691 2394 6768 2403
rect 6691 2334 6701 2394
rect 6757 2334 6768 2394
rect 6691 2324 6768 2334
rect -3953 2247 -3907 2308
rect -2577 2247 -2531 2302
rect -1201 2247 -1155 2303
rect 175 2247 221 2303
rect 1551 2247 1597 2303
rect 2927 2247 2973 2303
rect 4303 2247 4349 2302
rect 5679 2247 5725 2303
rect 7055 2247 7101 2303
rect -4339 2191 -4252 2210
rect -4090 2194 -4010 2210
rect -4090 2191 -4076 2194
rect -4339 2135 -4321 2191
rect -4265 2141 -4076 2191
rect -4026 2141 -4010 2194
rect -3953 2169 7410 2247
rect -4265 2135 -4010 2141
rect -4339 2124 -4252 2135
rect -4090 2125 -4010 2135
rect -3265 2051 -3219 2169
rect -1889 2051 -1843 2169
rect -513 2051 -467 2169
rect 863 2051 909 2169
rect 2239 2051 2285 2169
rect 3615 2051 3661 2169
rect 4991 2051 5037 2169
rect 6367 2051 6413 2169
rect -3625 2036 -3548 2045
rect -3625 1976 -3615 2036
rect -3559 1976 -3548 2036
rect -3625 1966 -3548 1976
rect -2943 2034 -2866 2043
rect -2943 1974 -2933 2034
rect -2877 1974 -2866 2034
rect -2943 1964 -2866 1974
rect -2254 2027 -2177 2036
rect -2254 1967 -2244 2027
rect -2188 1967 -2177 2027
rect -2254 1957 -2177 1967
rect -1568 2026 -1491 2035
rect -1568 1966 -1558 2026
rect -1502 1966 -1491 2026
rect -1568 1956 -1491 1966
rect -878 2022 -801 2031
rect -878 1962 -868 2022
rect -812 1962 -801 2022
rect -878 1952 -801 1962
rect -184 2025 -107 2034
rect -184 1965 -174 2025
rect -118 1965 -107 2025
rect -184 1955 -107 1965
rect 505 2025 582 2034
rect 505 1965 515 2025
rect 571 1965 582 2025
rect 505 1955 582 1965
rect 1194 2027 1271 2036
rect 1194 1967 1204 2027
rect 1260 1967 1271 2027
rect 1194 1957 1271 1967
rect 1877 2025 1954 2034
rect 1877 1965 1887 2025
rect 1943 1965 1954 2025
rect 1877 1955 1954 1965
rect 2567 2032 2644 2041
rect 2567 1972 2577 2032
rect 2633 1972 2644 2032
rect 2567 1962 2644 1972
rect 3256 2029 3333 2038
rect 3256 1969 3266 2029
rect 3322 1969 3333 2029
rect 3256 1959 3333 1969
rect 3942 2024 4019 2033
rect 3942 1964 3952 2024
rect 4008 1964 4019 2024
rect 3942 1954 4019 1964
rect 4629 2028 4706 2037
rect 4629 1968 4639 2028
rect 4695 1968 4706 2028
rect 4629 1958 4706 1968
rect 5321 2028 5398 2037
rect 5321 1968 5331 2028
rect 5387 1968 5398 2028
rect 5321 1958 5398 1968
rect 6010 2032 6087 2041
rect 6010 1972 6020 2032
rect 6076 1972 6087 2032
rect 6010 1962 6087 1972
rect 6690 2029 6767 2038
rect 6690 1969 6700 2029
rect 6756 1969 6767 2029
rect 6690 1959 6767 1969
rect -4136 1828 -4060 1841
rect -4136 1775 -4125 1828
rect -4072 1775 -4060 1828
rect -4136 1763 -4060 1775
rect -3953 1753 -3907 1935
rect -2577 1753 -2531 1935
rect -1201 1753 -1155 1935
rect 175 1753 221 1935
rect 1551 1753 1597 1935
rect 2927 1753 2973 1935
rect 4303 1753 4349 1935
rect 5679 1753 5725 1935
rect 7055 1753 7101 1935
rect -3991 1693 7113 1753
rect -3991 1534 -3926 1693
rect -3782 1534 -3676 1693
rect -3532 1534 -3426 1693
rect -3282 1534 -3176 1693
rect -3032 1534 -2926 1693
rect -2782 1534 -2676 1693
rect -2532 1534 -2426 1693
rect -2282 1534 -2176 1693
rect -2032 1534 -1926 1693
rect -1782 1534 -1676 1693
rect -1532 1534 -1426 1693
rect -1282 1534 -1176 1693
rect -1032 1534 -926 1693
rect -782 1534 -676 1693
rect -532 1534 -426 1693
rect -282 1534 -176 1693
rect -32 1534 74 1693
rect 218 1534 324 1693
rect 468 1534 574 1693
rect 718 1534 824 1693
rect 968 1534 1074 1693
rect 1218 1534 1324 1693
rect 1468 1534 1574 1693
rect 1718 1534 1824 1693
rect 1968 1534 2074 1693
rect 2218 1534 2324 1693
rect 2468 1534 2574 1693
rect 2718 1534 2824 1693
rect 2968 1534 3074 1693
rect 3218 1534 3324 1693
rect 3468 1534 3574 1693
rect 3718 1534 3824 1693
rect 3968 1534 4074 1693
rect 4218 1534 4324 1693
rect 4468 1534 4574 1693
rect 4718 1534 4824 1693
rect 4968 1534 5074 1693
rect 5218 1534 5324 1693
rect 5468 1534 5574 1693
rect 5718 1534 5824 1693
rect 5968 1534 6074 1693
rect 6218 1534 6324 1693
rect 6468 1534 6574 1693
rect 6718 1534 6824 1693
rect 6968 1676 7113 1693
rect 6968 1674 7037 1676
rect 6985 1620 7037 1674
rect 7093 1620 7113 1676
rect 6968 1559 7113 1620
rect 6968 1556 7038 1559
rect -3991 1500 6930 1534
rect 6986 1505 7038 1556
rect 7092 1505 7113 1559
rect 6986 1500 7113 1505
rect -3991 1468 7113 1500
rect -4149 1441 -4062 1455
rect -4149 1386 -4135 1441
rect -4077 1386 -4062 1441
rect -4149 1372 -4062 1386
rect -3265 1313 -3219 1468
rect -1889 1313 -1843 1468
rect -513 1313 -467 1468
rect 863 1313 909 1468
rect 2239 1313 2285 1468
rect 3615 1313 3661 1468
rect 4991 1313 5037 1468
rect 6367 1313 6413 1468
rect -3622 1294 -3545 1303
rect -3622 1233 -3612 1294
rect -3556 1233 -3545 1294
rect -3622 1223 -3545 1233
rect -2941 1297 -2864 1306
rect -2941 1237 -2931 1297
rect -2875 1237 -2864 1297
rect -2941 1227 -2864 1237
rect -2259 1292 -2182 1301
rect -2259 1232 -2249 1292
rect -2193 1232 -2182 1292
rect -2259 1222 -2182 1232
rect -1568 1285 -1491 1294
rect -1568 1225 -1558 1285
rect -1502 1225 -1491 1285
rect -1568 1215 -1491 1225
rect -879 1284 -802 1293
rect -879 1224 -869 1284
rect -813 1224 -802 1284
rect -879 1214 -802 1224
rect -187 1284 -110 1293
rect -187 1224 -177 1284
rect -121 1224 -110 1284
rect -187 1214 -110 1224
rect 502 1284 579 1293
rect 502 1224 512 1284
rect 568 1224 579 1284
rect 502 1214 579 1224
rect 1192 1288 1269 1297
rect 1192 1228 1202 1288
rect 1258 1228 1269 1288
rect 1192 1218 1269 1228
rect 1878 1289 1955 1298
rect 1878 1229 1888 1289
rect 1944 1229 1955 1289
rect 1878 1219 1955 1229
rect 2565 1290 2642 1299
rect 2565 1230 2575 1290
rect 2631 1230 2642 1290
rect 2565 1220 2642 1230
rect 3254 1287 3331 1296
rect 3254 1227 3264 1287
rect 3320 1227 3331 1287
rect 3254 1217 3331 1227
rect 3949 1291 4026 1300
rect 3949 1231 3959 1291
rect 4015 1231 4026 1291
rect 3949 1221 4026 1231
rect 4629 1292 4706 1301
rect 4629 1232 4639 1292
rect 4695 1232 4706 1292
rect 4629 1222 4706 1232
rect 5315 1289 5392 1298
rect 5315 1229 5325 1289
rect 5381 1229 5392 1289
rect 5315 1219 5392 1229
rect 6004 1285 6081 1294
rect 6004 1225 6014 1285
rect 6070 1225 6081 1285
rect 6004 1215 6081 1225
rect 6691 1289 6768 1298
rect 6691 1229 6701 1289
rect 6757 1229 6768 1289
rect 6691 1219 6768 1229
rect -3953 1142 -3907 1203
rect -2577 1142 -2531 1197
rect -1201 1142 -1155 1198
rect 175 1142 221 1198
rect 1551 1142 1597 1198
rect 2927 1142 2973 1198
rect 4303 1142 4349 1197
rect 5679 1142 5725 1198
rect 7055 1142 7101 1198
rect 7255 1142 7410 2169
rect -4333 1086 -4253 1096
rect -4333 1032 -4320 1086
rect -4266 1082 -4253 1086
rect -4104 1089 -4025 1106
rect -4104 1082 -4090 1089
rect -4266 1036 -4090 1082
rect -4038 1036 -4025 1089
rect -3953 1064 7410 1142
rect -4266 1032 -4253 1036
rect -4333 1009 -4253 1032
rect -4104 1021 -4025 1036
rect -3265 946 -3219 1064
rect -1889 946 -1843 1064
rect -513 946 -467 1064
rect 863 946 909 1064
rect 2239 946 2285 1064
rect 3615 946 3661 1064
rect 4991 946 5037 1064
rect 6367 946 6413 1064
rect -3625 931 -3548 940
rect -3625 871 -3615 931
rect -3559 871 -3548 931
rect -3625 861 -3548 871
rect -2943 929 -2866 938
rect -2943 869 -2933 929
rect -2877 869 -2866 929
rect -2943 859 -2866 869
rect -2254 922 -2177 931
rect -2254 862 -2244 922
rect -2188 862 -2177 922
rect -2254 852 -2177 862
rect -1568 921 -1491 930
rect -1568 861 -1558 921
rect -1502 861 -1491 921
rect -1568 851 -1491 861
rect -878 917 -801 926
rect -878 857 -868 917
rect -812 857 -801 917
rect -878 847 -801 857
rect -184 920 -107 929
rect -184 860 -174 920
rect -118 860 -107 920
rect -184 850 -107 860
rect 505 920 582 929
rect 505 860 515 920
rect 571 860 582 920
rect 505 850 582 860
rect 1194 922 1271 931
rect 1194 862 1204 922
rect 1260 862 1271 922
rect 1194 852 1271 862
rect 1877 920 1954 929
rect 1877 860 1887 920
rect 1943 860 1954 920
rect 1877 850 1954 860
rect 2567 927 2644 936
rect 2567 867 2577 927
rect 2633 867 2644 927
rect 2567 857 2644 867
rect 3256 924 3333 933
rect 3256 864 3266 924
rect 3322 864 3333 924
rect 3256 854 3333 864
rect 3942 919 4019 928
rect 3942 859 3952 919
rect 4008 859 4019 919
rect 3942 849 4019 859
rect 4629 923 4706 932
rect 4629 863 4639 923
rect 4695 863 4706 923
rect 4629 853 4706 863
rect 5321 923 5398 932
rect 5321 863 5331 923
rect 5387 863 5398 923
rect 5321 853 5398 863
rect 6010 927 6087 936
rect 6010 867 6020 927
rect 6076 867 6087 927
rect 6010 857 6087 867
rect 6690 924 6767 933
rect 6690 864 6700 924
rect 6756 864 6767 924
rect 6690 854 6767 864
rect -4136 723 -4060 737
rect -4136 671 -4124 723
rect -4072 671 -4060 723
rect -4136 658 -4060 671
rect -3953 648 -3907 830
rect -2577 648 -2531 830
rect -1201 648 -1155 830
rect 175 648 221 830
rect 1551 648 1597 830
rect 2927 648 2973 830
rect 4303 648 4349 830
rect 5679 648 5725 830
rect 6908 648 6992 649
rect 7055 648 7101 830
rect -3990 634 7116 648
rect -3990 632 7040 634
rect -3990 578 6934 632
rect 6988 578 7040 632
rect 7096 578 7116 634
rect -3990 568 7116 578
rect -3990 409 -3944 568
rect -3800 409 -3694 568
rect -3550 409 -3444 568
rect -3300 409 -3194 568
rect -3050 409 -2944 568
rect -2800 409 -2694 568
rect -2550 409 -2444 568
rect -2300 409 -2194 568
rect -2050 409 -1944 568
rect -1800 409 -1694 568
rect -1550 409 -1444 568
rect -1300 409 -1194 568
rect -1050 409 -944 568
rect -800 409 -694 568
rect -550 409 -444 568
rect -300 409 -194 568
rect -50 409 56 568
rect 200 409 306 568
rect 450 409 556 568
rect 700 409 806 568
rect 950 409 1056 568
rect 1200 409 1306 568
rect 1450 409 1556 568
rect 1700 409 1806 568
rect 1950 409 2056 568
rect 2200 409 2306 568
rect 2450 409 2556 568
rect 2700 409 2806 568
rect 2950 409 3056 568
rect 3200 409 3306 568
rect 3450 409 3556 568
rect 3700 409 3806 568
rect 3950 409 4056 568
rect 4200 409 4306 568
rect 4450 409 4556 568
rect 4700 409 4806 568
rect 4950 409 5056 568
rect 5200 409 5306 568
rect 5450 409 5556 568
rect 5700 409 5806 568
rect 5950 409 6056 568
rect 6200 409 6306 568
rect 6450 409 6556 568
rect 6700 409 6806 568
rect 6950 517 7116 568
rect 6950 514 7041 517
rect 6989 463 7041 514
rect 7095 463 7116 517
rect 6989 458 7116 463
rect 6950 409 7116 458
rect -3990 365 7116 409
<< via1 >>
rect 6931 2725 6968 2779
rect 6968 2725 6985 2779
rect 7037 2725 7093 2781
rect 6930 2639 6968 2661
rect 6968 2639 6986 2661
rect 6930 2605 6986 2639
rect 7038 2610 7092 2664
rect -4137 2545 -4076 2546
rect -4137 2491 -4135 2545
rect -4135 2491 -4077 2545
rect -4077 2491 -4076 2545
rect -4137 2489 -4076 2491
rect -3612 2338 -3556 2399
rect -2931 2342 -2875 2402
rect -2249 2337 -2193 2397
rect -1558 2330 -1502 2390
rect -869 2329 -813 2389
rect -177 2329 -121 2389
rect 512 2329 568 2389
rect 1202 2333 1258 2393
rect 1888 2334 1944 2394
rect 2575 2335 2631 2395
rect 3264 2332 3320 2392
rect 3959 2336 4015 2396
rect 4639 2337 4695 2397
rect 5325 2334 5381 2394
rect 6014 2330 6070 2390
rect 6701 2334 6757 2394
rect -4321 2135 -4265 2191
rect -3615 1976 -3559 2036
rect -2933 1974 -2877 2034
rect -2244 1967 -2188 2027
rect -1558 1966 -1502 2026
rect -868 1962 -812 2022
rect -174 1965 -118 2025
rect 515 1965 571 2025
rect 1204 1967 1260 2027
rect 1887 1965 1943 2025
rect 2577 1972 2633 2032
rect 3266 1969 3322 2029
rect 3952 1964 4008 2024
rect 4639 1968 4695 2028
rect 5331 1968 5387 2028
rect 6020 1972 6076 2032
rect 6700 1969 6756 2029
rect -4125 1776 -4123 1828
rect -4123 1776 -4074 1828
rect -4074 1776 -4072 1828
rect -4125 1775 -4072 1776
rect 6931 1620 6968 1674
rect 6968 1620 6985 1674
rect 7037 1620 7093 1676
rect 6930 1534 6968 1556
rect 6968 1534 6986 1556
rect 6930 1500 6986 1534
rect 7038 1505 7092 1559
rect -4135 1440 -4077 1441
rect -4135 1386 -4077 1440
rect -3612 1233 -3556 1294
rect -2931 1237 -2875 1297
rect -2249 1232 -2193 1292
rect -1558 1225 -1502 1285
rect -869 1224 -813 1284
rect -177 1224 -121 1284
rect 512 1224 568 1284
rect 1202 1228 1258 1288
rect 1888 1229 1944 1289
rect 2575 1230 2631 1290
rect 3264 1227 3320 1287
rect 3959 1231 4015 1291
rect 4639 1232 4695 1292
rect 5325 1229 5381 1289
rect 6014 1225 6070 1285
rect 6701 1229 6757 1289
rect -4320 1032 -4266 1086
rect -3615 871 -3559 931
rect -2933 869 -2877 929
rect -2244 862 -2188 922
rect -1558 861 -1502 921
rect -868 857 -812 917
rect -174 860 -118 920
rect 515 860 571 920
rect 1204 862 1260 922
rect 1887 860 1943 920
rect 2577 867 2633 927
rect 3266 864 3322 924
rect 3952 859 4008 919
rect 4639 863 4695 923
rect 5331 863 5387 923
rect 6020 867 6076 927
rect 6700 864 6756 924
rect -4124 671 -4123 723
rect -4123 671 -4074 723
rect -4074 671 -4072 723
rect 6934 578 6988 632
rect 7040 578 7096 634
rect 6933 458 6950 514
rect 6950 458 6989 514
rect 7041 463 7095 517
<< metal2 >>
rect 7030 2795 7086 2796
rect 6916 2781 7107 2795
rect 6916 2779 7037 2781
rect 6916 2725 6931 2779
rect 6985 2725 7037 2779
rect 7093 2725 7107 2781
rect 6916 2664 7107 2725
rect 6916 2661 7038 2664
rect 6916 2605 6930 2661
rect 6986 2610 7038 2661
rect 7092 2610 7107 2664
rect 6986 2605 7107 2610
rect 6916 2581 7107 2605
rect 6916 2573 7089 2581
rect -4148 2546 -4063 2560
rect -4148 2489 -4137 2546
rect -4076 2489 -4063 2546
rect -4148 2477 -4063 2489
rect -4339 2191 -4252 2210
rect -4339 2135 -4321 2191
rect -4265 2135 -4252 2191
rect -4339 2124 -4252 2135
rect -4321 1096 -4265 2124
rect -4133 1846 -4077 2477
rect -3622 2399 -3545 2408
rect -3622 2338 -3612 2399
rect -3556 2338 -3545 2399
rect -3622 2328 -3545 2338
rect -2941 2402 -2864 2411
rect -2941 2342 -2931 2402
rect -2875 2342 -2864 2402
rect -2941 2332 -2864 2342
rect -2259 2397 -2182 2406
rect -2259 2337 -2249 2397
rect -2193 2337 -2182 2397
rect -3619 2056 -3563 2328
rect -2933 2056 -2877 2332
rect -2259 2327 -2182 2337
rect -1568 2390 -1491 2399
rect -1568 2330 -1558 2390
rect -1502 2330 -1491 2390
rect -2246 2056 -2190 2327
rect -1568 2320 -1491 2330
rect -879 2389 -802 2398
rect -879 2329 -869 2389
rect -813 2329 -802 2389
rect -1556 2056 -1500 2320
rect -879 2319 -802 2329
rect -187 2389 -110 2398
rect -187 2329 -177 2389
rect -121 2329 -110 2389
rect -187 2319 -110 2329
rect 502 2389 579 2398
rect 502 2329 512 2389
rect 568 2329 579 2389
rect 502 2319 579 2329
rect 1192 2393 1269 2402
rect 1192 2333 1202 2393
rect 1258 2333 1269 2393
rect 1192 2323 1269 2333
rect 1878 2394 1955 2403
rect 1878 2334 1888 2394
rect 1944 2334 1955 2394
rect 1878 2324 1955 2334
rect 2565 2395 2642 2404
rect 2565 2335 2575 2395
rect 2631 2335 2642 2395
rect 2565 2325 2642 2335
rect 3254 2392 3331 2401
rect 3254 2332 3264 2392
rect 3320 2332 3331 2392
rect -867 2056 -811 2319
rect -174 2056 -118 2319
rect 514 2056 570 2319
rect 1201 2056 1257 2323
rect 1889 2056 1945 2324
rect 2582 2056 2638 2325
rect 3254 2322 3331 2332
rect 3949 2396 4026 2405
rect 3949 2336 3959 2396
rect 4015 2336 4026 2396
rect 3949 2326 4026 2336
rect 4629 2397 4706 2406
rect 4629 2337 4639 2397
rect 4695 2337 4706 2397
rect 4629 2327 4706 2337
rect 5315 2394 5392 2403
rect 5315 2334 5325 2394
rect 5381 2334 5392 2394
rect 3266 2056 3322 2322
rect 3955 2056 4011 2326
rect 4640 2056 4696 2327
rect 5315 2324 5392 2334
rect 6004 2390 6081 2399
rect 6004 2330 6014 2390
rect 6070 2330 6081 2390
rect 5331 2056 5387 2324
rect 6004 2320 6081 2330
rect 6691 2394 6768 2403
rect 6691 2334 6701 2394
rect 6757 2334 6768 2394
rect 6691 2324 6768 2334
rect 6018 2056 6074 2320
rect 6704 2056 6760 2324
rect -3619 2045 6777 2056
rect -3625 2036 6777 2045
rect -3625 1976 -3615 2036
rect -3559 2034 6777 2036
rect -3559 1976 -2933 2034
rect -3625 1974 -2933 1976
rect -2877 2032 6777 2034
rect -2877 2027 2577 2032
rect -2877 1974 -2244 2027
rect -3625 1967 -2244 1974
rect -2188 2026 1204 2027
rect -2188 1967 -1558 2026
rect -3625 1966 -3548 1967
rect -4139 1828 -4055 1846
rect -4139 1775 -4125 1828
rect -4072 1775 -4055 1828
rect -4139 1762 -4055 1775
rect -4133 1455 -4077 1762
rect -4149 1441 -4062 1455
rect -4149 1386 -4135 1441
rect -4077 1386 -4062 1441
rect -4149 1372 -4062 1386
rect -4333 1086 -4253 1096
rect -4333 1032 -4320 1086
rect -4266 1032 -4253 1086
rect -4333 1009 -4253 1032
rect -4133 737 -4077 1372
rect -3619 1303 -3563 1966
rect -2943 1964 -2866 1967
rect -2933 1306 -2877 1964
rect -2254 1957 -2177 1967
rect -1568 1966 -1558 1967
rect -1502 2025 1204 2026
rect -1502 2022 -174 2025
rect -1502 1967 -868 2022
rect -1502 1966 -1491 1967
rect -3622 1294 -3545 1303
rect -3622 1233 -3612 1294
rect -3556 1233 -3545 1294
rect -3622 1223 -3545 1233
rect -2941 1297 -2864 1306
rect -2246 1301 -2190 1957
rect -1568 1956 -1491 1966
rect -878 1962 -868 1967
rect -812 1967 -174 2022
rect -812 1962 -801 1967
rect -2941 1237 -2931 1297
rect -2875 1237 -2864 1297
rect -2941 1227 -2864 1237
rect -2259 1292 -2182 1301
rect -1556 1294 -1500 1956
rect -878 1952 -801 1962
rect -184 1965 -174 1967
rect -118 1967 515 2025
rect -118 1965 -107 1967
rect -184 1955 -107 1965
rect 505 1965 515 1967
rect 571 1967 1204 2025
rect 1260 2025 2577 2027
rect 1260 1967 1887 2025
rect 571 1965 582 1967
rect 505 1955 582 1965
rect 1194 1957 1271 1967
rect 1877 1965 1887 1967
rect 1943 1972 2577 2025
rect 2633 2029 6020 2032
rect 2633 1972 3266 2029
rect 1943 1969 3266 1972
rect 3322 2028 6020 2029
rect 3322 2024 4639 2028
rect 3322 1969 3952 2024
rect 1943 1967 3952 1969
rect 1943 1965 1954 1967
rect -2259 1232 -2249 1292
rect -2193 1232 -2182 1292
rect -3619 951 -3563 1223
rect -2933 951 -2877 1227
rect -2259 1222 -2182 1232
rect -1568 1285 -1491 1294
rect -867 1293 -811 1952
rect -174 1293 -118 1955
rect 514 1293 570 1955
rect 1201 1297 1257 1957
rect 1877 1955 1954 1965
rect 2567 1962 2644 1967
rect 1889 1298 1945 1955
rect 2582 1299 2638 1962
rect 3256 1959 3333 1967
rect 3942 1964 3952 1967
rect 4008 1968 4639 2024
rect 4695 1968 5331 2028
rect 5387 1972 6020 2028
rect 6076 2029 6777 2032
rect 6076 1972 6700 2029
rect 5387 1969 6700 1972
rect 6756 1969 6777 2029
rect 5387 1968 6777 1969
rect 4008 1967 6777 1968
rect 4008 1964 4019 1967
rect -1568 1225 -1558 1285
rect -1502 1225 -1491 1285
rect -2246 951 -2190 1222
rect -1568 1215 -1491 1225
rect -879 1284 -802 1293
rect -879 1224 -869 1284
rect -813 1224 -802 1284
rect -1556 951 -1500 1215
rect -879 1214 -802 1224
rect -187 1284 -110 1293
rect -187 1224 -177 1284
rect -121 1224 -110 1284
rect -187 1214 -110 1224
rect 502 1284 579 1293
rect 502 1224 512 1284
rect 568 1224 579 1284
rect 502 1214 579 1224
rect 1192 1288 1269 1297
rect 1192 1228 1202 1288
rect 1258 1228 1269 1288
rect 1192 1218 1269 1228
rect 1878 1289 1955 1298
rect 1878 1229 1888 1289
rect 1944 1229 1955 1289
rect 1878 1219 1955 1229
rect 2565 1290 2642 1299
rect 3266 1296 3322 1959
rect 3942 1954 4019 1964
rect 4629 1958 4706 1967
rect 5321 1958 5398 1967
rect 6010 1962 6087 1967
rect 3955 1300 4011 1954
rect 4640 1301 4696 1958
rect 2565 1230 2575 1290
rect 2631 1230 2642 1290
rect 2565 1220 2642 1230
rect 3254 1287 3331 1296
rect 3254 1227 3264 1287
rect 3320 1227 3331 1287
rect -867 951 -811 1214
rect -174 951 -118 1214
rect 514 951 570 1214
rect 1201 951 1257 1218
rect 1889 951 1945 1219
rect 2582 951 2638 1220
rect 3254 1217 3331 1227
rect 3949 1291 4026 1300
rect 3949 1231 3959 1291
rect 4015 1231 4026 1291
rect 3949 1221 4026 1231
rect 4629 1292 4706 1301
rect 5331 1298 5387 1958
rect 4629 1232 4639 1292
rect 4695 1232 4706 1292
rect 4629 1222 4706 1232
rect 5315 1289 5392 1298
rect 6018 1294 6074 1962
rect 6690 1959 6767 1967
rect 6704 1298 6760 1959
rect 6919 1690 7089 2573
rect 6916 1676 7107 1690
rect 6916 1674 7037 1676
rect 6916 1620 6931 1674
rect 6985 1620 7037 1674
rect 7093 1620 7107 1676
rect 6916 1559 7107 1620
rect 6916 1556 7038 1559
rect 6916 1500 6930 1556
rect 6986 1505 7038 1556
rect 7092 1505 7107 1559
rect 6986 1500 7107 1505
rect 6916 1476 7107 1500
rect 6916 1468 7089 1476
rect 5315 1229 5325 1289
rect 5381 1229 5392 1289
rect 3266 951 3322 1217
rect 3955 951 4011 1221
rect 4640 951 4696 1222
rect 5315 1219 5392 1229
rect 6004 1285 6081 1294
rect 6004 1225 6014 1285
rect 6070 1225 6081 1285
rect 5331 951 5387 1219
rect 6004 1215 6081 1225
rect 6691 1289 6768 1298
rect 6691 1229 6701 1289
rect 6757 1229 6768 1289
rect 6691 1219 6768 1229
rect 6018 951 6074 1215
rect 6704 951 6760 1219
rect -3619 940 6777 951
rect -3625 931 6777 940
rect -3625 871 -3615 931
rect -3559 929 6777 931
rect -3559 871 -2933 929
rect -3625 869 -2933 871
rect -2877 927 6777 929
rect -2877 922 2577 927
rect -2877 869 -2244 922
rect -3625 862 -2244 869
rect -2188 921 1204 922
rect -2188 862 -1558 921
rect -3625 861 -3548 862
rect -2943 859 -2866 862
rect -2254 852 -2177 862
rect -1568 861 -1558 862
rect -1502 920 1204 921
rect -1502 917 -174 920
rect -1502 862 -868 917
rect -1502 861 -1491 862
rect -1568 851 -1491 861
rect -878 857 -868 862
rect -812 862 -174 917
rect -812 857 -801 862
rect -878 847 -801 857
rect -184 860 -174 862
rect -118 862 515 920
rect -118 860 -107 862
rect -184 850 -107 860
rect 505 860 515 862
rect 571 862 1204 920
rect 1260 920 2577 922
rect 1260 862 1887 920
rect 571 860 582 862
rect 505 850 582 860
rect 1194 852 1271 862
rect 1877 860 1887 862
rect 1943 867 2577 920
rect 2633 924 6020 927
rect 2633 867 3266 924
rect 1943 864 3266 867
rect 3322 923 6020 924
rect 3322 919 4639 923
rect 3322 864 3952 919
rect 1943 862 3952 864
rect 1943 860 1954 862
rect 1877 850 1954 860
rect 2567 857 2644 862
rect 3256 854 3333 862
rect 3942 859 3952 862
rect 4008 863 4639 919
rect 4695 863 5331 923
rect 5387 867 6020 923
rect 6076 924 6777 927
rect 6076 867 6700 924
rect 5387 864 6700 867
rect 6756 864 6777 924
rect 5387 863 6777 864
rect 4008 862 6777 863
rect 4008 859 4019 862
rect 3942 849 4019 859
rect 4629 853 4706 862
rect 5321 853 5398 862
rect 6010 857 6087 862
rect 6690 854 6767 862
rect -4136 723 -4060 737
rect -4136 671 -4124 723
rect -4072 671 -4060 723
rect -4136 658 -4060 671
rect 6919 649 7089 1468
rect 6908 648 7089 649
rect 6908 634 7110 648
rect 6908 632 7040 634
rect 6908 578 6934 632
rect 6988 578 7040 632
rect 7096 578 7110 634
rect 6908 517 7110 578
rect 6908 514 7041 517
rect 6908 458 6933 514
rect 6989 463 7041 514
rect 7095 463 7110 517
rect 6989 458 7110 463
rect 6908 434 7110 458
rect 6908 431 6992 434
use nmos_3p3_9N32EK  nmos_3p3_9N32EK_0
timestamp 1693281404
transform 1 0 1574 0 1 2360
box -5564 -128 5564 128
use nmos_3p3_9N32EK  nmos_3p3_9N32EK_1
timestamp 1693281404
transform 1 0 1574 0 1 1993
box -5564 -128 5564 128
use nmos_3p3_9N32EK  nmos_3p3_9N32EK_2
timestamp 1693281404
transform 1 0 1574 0 1 888
box -5564 -128 5564 128
use nmos_3p3_9N32EK  nmos_3p3_9N32EK_3
timestamp 1693281404
transform 1 0 1574 0 1 1255
box -5564 -128 5564 128
<< labels >>
flabel via1 -4111 2524 -4111 2524 0 FreeSans 1600 0 0 0 IM_T
port 0 nsew
flabel via1 -4296 1055 -4296 1055 0 FreeSans 1600 0 0 0 IM
port 1 nsew
flabel psubdiffcont -2576 2763 -2576 2763 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 7347 1582 7347 1582 0 FreeSans 1600 0 0 0 OUT
port 3 nsew
flabel via1 -3600 2010 -3600 2010 0 FreeSans 1600 0 0 0 SD
port 4 nsew
<< end >>
