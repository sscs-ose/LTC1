* NGSPICE file created from CM_MSB_V2_flat_flat.ext - technology: gf180mcuC

.subckt CM_MSB_V2_flat_flat IM_T VSS OUT IM SD
X0 SD IM_T.t0 OUT.t27 VSS.t0 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X1 SD IM.t0 VSS.t77 VSS.t59 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X2 VSS IM.t1 SD.t52 VSS.t51 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X3 VSS IM.t2 SD.t60 VSS.t50 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X4 SD IM_T.t1 OUT.t26 VSS.t61 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X5 SD IM_T.t2 OUT.t25 VSS.t9 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X6 OUT IM_T.t3 SD.t48 VSS.t60 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X7 SD IM.t3 VSS.t1 VSS.t0 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X8 SD IM_T.t4 OUT.t24 VSS.t59 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X9 OUT IM_T.t5 SD.t46 VSS.t47 nfet_03v3 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
X10 VSS IM.t4 SD.t12 VSS.t31 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X11 SD IM.t5 VSS.t21 VSS.t20 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X12 SD IM.t6 VSS.t10 VSS.t9 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X13 VSS IM.t7 SD.t53 VSS.t60 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X14 SD IM_T.t6 OUT.t23 VSS.t34 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X15 OUT IM_T.t7 SD.t44 VSS.t31 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X16 SD IM_T.t8 OUT.t22 VSS.t20 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X17 SD IM.t8 VSS.t3 VSS.t2 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X18 OUT IM_T.t9 SD.t42 VSS.t11 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X19 SD IM.t9 VSS.t35 VSS.t34 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X20 VSS IM.t10 SD.t9 VSS.t22 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X21 SD IM_T.t10 OUT.t21 VSS.t2 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X22 VSS IM.t11 SD.t5 VSS.t11 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X23 OUT IM_T.t11 SD.t40 VSS.t58 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X24 OUT IM_T.t12 SD.t39 VSS.t22 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X25 VSS IM.t12 SD.t55 VSS.t58 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X26 SD IM_T.t13 OUT.t20 VSS.t57 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X27 SD IM.t13 VSS.t74 VSS.t56 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X28 VSS IM.t14 SD.t58 VSS.t55 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X29 SD IM_T.t14 OUT.t19 VSS.t41 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X30 SD IM.t15 VSS.t78 VSS.t57 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X31 SD IM_T.t15 OUT.t18 VSS.t36 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X32 OUT IM_T.t16 SD.t35 VSS.t25 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X33 SD IM.t16 VSS.t42 VSS.t41 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X34 SD IM_T.t17 OUT.t17 VSS.t56 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X35 OUT IM_T.t18 SD.t33 VSS.t55 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X36 SD IM.t17 VSS.t46 VSS.t45 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X37 VSS IM.t18 SD.t2 VSS.t4 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X38 SD IM.t19 VSS.t37 VSS.t36 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X39 VSS IM.t20 SD.t10 VSS.t25 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X40 VSS IM.t21 SD.t6 VSS.t14 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X41 SD IM_T.t19 OUT.t16 VSS.t54 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X42 SD IM_T.t20 OUT.t15 VSS.t45 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X43 OUT IM_T.t21 SD.t30 VSS.t4 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X44 OUT IM_T.t22 SD.t29 VSS.t53 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X45 SD IM.t22 VSS.t66 VSS.t52 nfet_03v3 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X46 OUT IM_T.t23 SD.t28 VSS.t17 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X47 SD IM.t23 VSS.t8 VSS.t7 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X48 VSS IM.t24 SD.t15 VSS.t38 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X49 OUT IM_T.t24 SD.t27 VSS.t14 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X50 SD IM.t25 VSS.t71 VSS.t54 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X51 VSS IM.t26 SD.t11 VSS.t28 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X52 SD IM_T.t25 OUT.t14 VSS.t43 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X53 SD IM_T.t26 OUT.t13 VSS.t52 nfet_03v3 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X54 VSS IM.t27 SD.t7 VSS.t17 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X55 SD IM_T.t27 OUT.t12 VSS.t7 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X56 OUT IM_T.t28 SD.t23 VSS.t38 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X57 VSS IM.t28 SD.t56 VSS.t53 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X58 OUT IM_T.t29 SD.t22 VSS.t51 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X59 OUT IM_T.t30 SD.t21 VSS.t50 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X60 SD IM.t29 VSS.t79 VSS.t61 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X61 OUT IM_T.t31 SD.t20 VSS.t28 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X62 SD IM.t30 VSS.t44 VSS.t43 nfet_03v3 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X63 VSS IM.t31 SD.t19 VSS.t47 nfet_03v3 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
R0 IM_T.n18 IM_T.t5 84.5899
R1 IM_T.n20 IM_T.n19 64.4419
R2 IM_T.n22 IM_T.n21 64.4419
R3 IM_T.n24 IM_T.n23 64.4419
R4 IM_T.n26 IM_T.n25 64.4419
R5 IM_T.n28 IM_T.n27 64.4419
R6 IM_T.n30 IM_T.n29 64.4419
R7 IM_T.n32 IM_T.n31 64.4419
R8 IM_T.n1 IM_T.n0 63.3497
R9 IM_T.n3 IM_T.n2 63.3497
R10 IM_T.n5 IM_T.n4 63.3497
R11 IM_T.n7 IM_T.n6 63.3497
R12 IM_T.n9 IM_T.n8 63.3497
R13 IM_T.n11 IM_T.n10 63.3497
R14 IM_T.n13 IM_T.n12 63.3497
R15 IM_T.n15 IM_T.n14 57.7181
R16 IM_T.n0 IM_T.t25 31.3373
R17 IM_T.n33 IM_T.n32 31.1676
R18 IM_T.n18 IM_T.t1 20.1485
R19 IM_T.n19 IM_T.t28 20.1485
R20 IM_T.n20 IM_T.t17 20.1485
R21 IM_T.n21 IM_T.t21 20.1485
R22 IM_T.n22 IM_T.t8 20.1485
R23 IM_T.n23 IM_T.t12 20.1485
R24 IM_T.n24 IM_T.t4 20.1485
R25 IM_T.n25 IM_T.t31 20.1485
R26 IM_T.n26 IM_T.t27 20.1485
R27 IM_T.n27 IM_T.t24 20.1485
R28 IM_T.n28 IM_T.t20 20.1485
R29 IM_T.n29 IM_T.t18 20.1485
R30 IM_T.n30 IM_T.t10 20.1485
R31 IM_T.n31 IM_T.t7 20.1485
R32 IM_T.n32 IM_T.t26 20.1485
R33 IM_T.n0 IM_T.t22 18.4695
R34 IM_T.n1 IM_T.t19 18.4695
R35 IM_T.n2 IM_T.t16 18.4695
R36 IM_T.n3 IM_T.t14 18.4695
R37 IM_T.n4 IM_T.t9 18.4695
R38 IM_T.n5 IM_T.t6 18.4695
R39 IM_T.n6 IM_T.t3 18.4695
R40 IM_T.n7 IM_T.t2 18.4695
R41 IM_T.n8 IM_T.t30 18.4695
R42 IM_T.n9 IM_T.t15 18.4695
R43 IM_T.n10 IM_T.t23 18.4695
R44 IM_T.n11 IM_T.t13 18.4695
R45 IM_T.n12 IM_T.t11 18.4695
R46 IM_T.n13 IM_T.t0 18.4695
R47 IM_T.n14 IM_T.t29 18.4695
R48 IM_T.n19 IM_T.n18 13.0902
R49 IM_T.n21 IM_T.n20 13.0902
R50 IM_T.n23 IM_T.n22 13.0902
R51 IM_T.n25 IM_T.n24 13.0902
R52 IM_T.n27 IM_T.n26 13.0902
R53 IM_T.n29 IM_T.n28 13.0902
R54 IM_T.n31 IM_T.n30 13.0902
R55 IM_T.n2 IM_T.n1 12.8683
R56 IM_T.n4 IM_T.n3 12.8683
R57 IM_T.n6 IM_T.n5 12.8683
R58 IM_T.n8 IM_T.n7 12.8683
R59 IM_T.n10 IM_T.n9 12.8683
R60 IM_T.n12 IM_T.n11 12.8683
R61 IM_T.n14 IM_T.n13 12.8683
R62 IM_T.n34 IM_T.n17 4.52219
R63 IM_T.n34 IM_T.n33 2.25726
R64 IM_T.n16 IM_T.n15 2.24422
R65 IM_T.n34 IM_T.n15 0.0145636
R66 IM_T.n17 IM_T.n16 0.00700602
R67 IM_T IM_T.n34 0.00154651
R68 OUT.n31 OUT.t13 5.37963
R69 OUT.n46 OUT.n0 4.86963
R70 OUT.n31 OUT.n30 3.61615
R71 OUT.n33 OUT.n26 3.61615
R72 OUT.n35 OUT.n22 3.61615
R73 OUT.n37 OUT.n18 3.61615
R74 OUT.n39 OUT.n14 3.61615
R75 OUT.n41 OUT.n10 3.61615
R76 OUT.n43 OUT.n6 3.61615
R77 OUT.n45 OUT.n2 3.61615
R78 OUT.n44 OUT.n4 3.50463
R79 OUT.n42 OUT.n8 3.50463
R80 OUT.n40 OUT.n12 3.50463
R81 OUT.n38 OUT.n16 3.50463
R82 OUT.n36 OUT.n20 3.50463
R83 OUT.n34 OUT.n24 3.50463
R84 OUT.n32 OUT.n28 3.50463
R85 OUT.n4 OUT.t26 1.3655
R86 OUT.n4 OUT.n3 1.3655
R87 OUT.n8 OUT.t17 1.3655
R88 OUT.n8 OUT.n7 1.3655
R89 OUT.n12 OUT.t22 1.3655
R90 OUT.n12 OUT.n11 1.3655
R91 OUT.n16 OUT.t24 1.3655
R92 OUT.n16 OUT.n15 1.3655
R93 OUT.n20 OUT.t12 1.3655
R94 OUT.n20 OUT.n19 1.3655
R95 OUT.n24 OUT.t15 1.3655
R96 OUT.n24 OUT.n23 1.3655
R97 OUT.n28 OUT.t21 1.3655
R98 OUT.n28 OUT.n27 1.3655
R99 OUT.n30 OUT.t27 1.3655
R100 OUT.n30 OUT.n29 1.3655
R101 OUT.n26 OUT.t20 1.3655
R102 OUT.n26 OUT.n25 1.3655
R103 OUT.n22 OUT.t18 1.3655
R104 OUT.n22 OUT.n21 1.3655
R105 OUT.n18 OUT.t25 1.3655
R106 OUT.n18 OUT.n17 1.3655
R107 OUT.n14 OUT.t23 1.3655
R108 OUT.n14 OUT.n13 1.3655
R109 OUT.n10 OUT.t19 1.3655
R110 OUT.n10 OUT.n9 1.3655
R111 OUT.n6 OUT.t16 1.3655
R112 OUT.n6 OUT.n5 1.3655
R113 OUT.n2 OUT.t14 1.3655
R114 OUT.n2 OUT.n1 1.3655
R115 OUT.n46 OUT.n45 0.5105
R116 OUT.n45 OUT.n44 0.5105
R117 OUT.n44 OUT.n43 0.5105
R118 OUT.n43 OUT.n42 0.5105
R119 OUT.n42 OUT.n41 0.5105
R120 OUT.n41 OUT.n40 0.5105
R121 OUT.n40 OUT.n39 0.5105
R122 OUT.n39 OUT.n38 0.5105
R123 OUT.n38 OUT.n37 0.5105
R124 OUT.n37 OUT.n36 0.5105
R125 OUT.n36 OUT.n35 0.5105
R126 OUT.n35 OUT.n34 0.5105
R127 OUT.n34 OUT.n33 0.5105
R128 OUT.n33 OUT.n32 0.5105
R129 OUT.n32 OUT.n31 0.5105
R130 OUT OUT.n46 0.33675
R131 SD.n81 SD.n79 6.36527
R132 SD.n85 SD.n84 4.5005
R133 SD.n67 SD.n12 3.63741
R134 SD.n41 SD.n40 3.28149
R135 SD.n52 SD.n26 3.28101
R136 SD.n64 SD.n17 3.27542
R137 SD.n78 SD.n1 3.26817
R138 SD.n109 SD.n91 3.258
R139 SD.n43 SD.n33 3.25644
R140 SD.n76 SD.n3 3.24511
R141 SD.n98 SD.n95 3.23798
R142 SD.n100 SD.n93 3.23061
R143 SD.n73 SD.n10 3.2111
R144 SD.n58 SD.n19 3.20644
R145 SD.n55 SD.n21 3.20496
R146 SD.n49 SD.n31 3.204
R147 SD.n111 SD.n89 3.19428
R148 SD.n116 SD.n87 3.16815
R149 SD.n114 SD.n113 2.58749
R150 SD.n75 SD.n5 2.5852
R151 SD.n41 SD.n38 2.57457
R152 SD.n98 SD.n97 2.56564
R153 SD.n48 SD.n47 2.24976
R154 SD.n62 SD.n61 2.24638
R155 SD.n104 SD.n103 2.24631
R156 SD.n71 SD.n70 2.24557
R157 SD.n120 SD.n119 2.24508
R158 SD.n84 SD.n83 1.85761
R159 SD.n54 SD.n24 1.49577
R160 SD.n108 SD.n107 1.49553
R161 SD.n74 SD.n8 1.49548
R162 SD.n42 SD.n36 1.49542
R163 SD.n65 SD.n15 1.49542
R164 SD.n51 SD.n29 1.49542
R165 SD.n113 SD.t58 1.47093
R166 SD.n26 SD.t10 1.47081
R167 SD.n1 SD.t27 1.4708
R168 SD.n17 SD.t39 1.46022
R169 SD.n5 SD.t21 1.4602
R170 SD.n91 SD.t55 1.46017
R171 SD.n33 SD.t56 1.46008
R172 SD.n69 SD.n68 1.45967
R173 SD.n46 SD.n45 1.45927
R174 SD.n3 SD.n2 1.45919
R175 SD.n60 SD.n59 1.45916
R176 SD.n119 SD.n118 1.4476
R177 SD.n107 SD.n106 1.44722
R178 SD.n15 SD.n14 1.44631
R179 SD.n36 SD.n35 1.4456
R180 SD.n29 SD.n28 1.44501
R181 SD.n8 SD.n7 1.44371
R182 SD.n24 SD.n23 1.44299
R183 SD.n102 SD.t12 1.42418
R184 SD.n40 SD.n39 1.41105
R185 SD.n118 SD.t28 1.3655
R186 SD.n118 SD.n117 1.3655
R187 SD.n106 SD.t40 1.3655
R188 SD.n106 SD.n105 1.3655
R189 SD.n97 SD.t22 1.3655
R190 SD.n97 SD.n96 1.3655
R191 SD.n95 SD.t52 1.3655
R192 SD.n95 SD.n94 1.3655
R193 SD.n93 SD.t44 1.3655
R194 SD.n93 SD.n92 1.3655
R195 SD.n89 SD.t33 1.3655
R196 SD.n89 SD.n88 1.3655
R197 SD.n87 SD.t7 1.3655
R198 SD.n87 SD.n86 1.3655
R199 SD.n7 SD.t11 1.3655
R200 SD.n7 SD.n6 1.3655
R201 SD.n14 SD.t9 1.3655
R202 SD.n14 SD.n13 1.3655
R203 SD.n23 SD.t2 1.3655
R204 SD.n23 SD.n22 1.3655
R205 SD.n28 SD.t35 1.3655
R206 SD.n28 SD.n27 1.3655
R207 SD.n35 SD.t29 1.3655
R208 SD.n35 SD.n34 1.3655
R209 SD.n38 SD.t19 1.3655
R210 SD.n38 SD.n37 1.3655
R211 SD.n31 SD.t23 1.3655
R212 SD.n31 SD.n30 1.3655
R213 SD.n21 SD.t30 1.3655
R214 SD.n21 SD.n20 1.3655
R215 SD.n19 SD.t5 1.3655
R216 SD.n19 SD.n18 1.3655
R217 SD.n12 SD.t53 1.3655
R218 SD.n12 SD.n11 1.3655
R219 SD.n10 SD.t20 1.3655
R220 SD.n10 SD.n9 1.3655
R221 SD.n83 SD.n82 1.34398
R222 SD.n40 SD.t46 1.28824
R223 SD.n102 SD.n101 1.2738
R224 SD.n60 SD.t42 1.23341
R225 SD.n3 SD.t60 1.23339
R226 SD.n46 SD.t15 1.23331
R227 SD.n69 SD.t48 1.23295
R228 SD.n33 SD.n32 1.23247
R229 SD.n91 SD.n90 1.23239
R230 SD.n5 SD.n4 1.23236
R231 SD.n17 SD.n16 1.23234
R232 SD.n1 SD.n0 1.21851
R233 SD.n26 SD.n25 1.21849
R234 SD.n113 SD.n112 1.21839
R235 SD.n70 SD.n69 1.09468
R236 SD.n47 SD.n46 1.09004
R237 SD.n61 SD.n60 1.08871
R238 SD.n103 SD.n102 1.08617
R239 SD.n80 SD.t6 0.81425
R240 SD.n77 SD.n76 0.605393
R241 SD.n99 SD.n98 0.603024
R242 SD.n66 SD.n65 0.590381
R243 SD.n48 SD.n44 0.57793
R244 SD.n111 SD.n110 0.571801
R245 SD.n42 SD.n41 0.571708
R246 SD.n57 SD.n56 0.570677
R247 SD.n75 SD.n74 0.57026
R248 SD.n115 SD.n114 0.56537
R249 SD.n54 SD.n53 0.560195
R250 SD.n108 SD.n104 0.558901
R251 SD.n51 SD.n50 0.553694
R252 SD.n81 SD.n80 0.55175
R253 SD.n121 SD.n120 0.551536
R254 SD.n72 SD.n71 0.54879
R255 SD.n63 SD.n62 0.545974
R256 SD.n73 SD.n72 0.0239783
R257 SD.n64 SD.n63 0.0232473
R258 SD.n83 SD.n81 0.0226604
R259 SD.n53 SD.n52 0.0202802
R260 SD.n110 SD.n109 0.0192912
R261 SD.n44 SD.n43 0.0192912
R262 SD.n56 SD.n55 0.0181289
R263 SD.n43 SD.n42 0.0164699
R264 SD.n104 SD.n100 0.0163101
R265 SD SD.n121 0.0153352
R266 SD.n109 SD.n108 0.0151457
R267 SD.n55 SD.n54 0.0149378
R268 SD.n52 SD.n51 0.0148219
R269 SD.n116 SD.n115 0.0148149
R270 SD.n50 SD.n49 0.0143462
R271 SD.n71 SD.n67 0.0138309
R272 SD.n76 SD.n75 0.0138281
R273 SD.n120 SD.n116 0.0138259
R274 SD.n114 SD.n111 0.0134986
R275 SD.n62 SD.n58 0.0119156
R276 SD.n65 SD.n64 0.0115197
R277 SD.n49 SD.n48 0.0113833
R278 SD.n74 SD.n73 0.011083
R279 SD SD.n85 0.00643407
R280 SD.n84 SD.n79 0.00579412
R281 SD.n67 SD.n66 0.00445604
R282 SD.n78 SD.n77 0.00445604
R283 SD.n58 SD.n57 0.00386449
R284 SD.n100 SD.n99 0.00247802
R285 SD.n85 SD.n78 0.00247802
R286 VSS.n159 VSS.t0 326.524
R287 VSS.n80 VSS.t38 317.817
R288 VSS.n105 VSS.t56 300.402
R289 VSS.n13 VSS.t43 291.695
R290 VSS.n172 VSS.t58 291.695
R291 VSS.n112 VSS.t11 274.281
R292 VSS.n145 VSS.t45 265.574
R293 VSS.n120 VSS.t34 248.159
R294 VSS.n136 VSS.t14 239.452
R295 VSS.n128 VSS.t28 222.036
R296 VSS.n127 VSS.t9 213.329
R297 VSS.n137 VSS.t7 195.915
R298 VSS.n119 VSS.t60 187.208
R299 VSS.n146 VSS.t17 169.792
R300 VSS.n63 VSS.t20 161.085
R301 VSS.n88 VSS.t47 143.671
R302 VSS.n173 VSS.t57 143.671
R303 VSS.n69 VSS.t4 134.964
R304 VSS.n95 VSS.t61 117.549
R305 VSS.n164 VSS.t31 117.549
R306 VSS.n76 VSS.t54 108.841
R307 VSS.n158 VSS.t51 108.841
R308 VSS.n102 VSS.t25 91.4272
R309 VSS.n157 VSS.t52 91.4272
R310 VSS.n83 VSS.t53 82.7199
R311 VSS.n167 VSS.t2 82.7199
R312 VSS.n108 VSS.t41 65.3053
R313 VSS.n149 VSS.t55 56.598
R314 VSS.n115 VSS.t22 39.1833
R315 VSS.n140 VSS.t36 30.4761
R316 VSS.n124 VSS.t59 13.0615
R317 VSS.n120 VSS.n119 8.7078
R318 VSS.n124 VSS.n123 8.7078
R319 VSS.n128 VSS.n127 8.7078
R320 VSS.n133 VSS.n132 8.7078
R321 VSS.n137 VSS.n136 8.7078
R322 VSS.n141 VSS.n140 8.7078
R323 VSS.n146 VSS.n145 8.7078
R324 VSS.n150 VSS.n149 8.7078
R325 VSS.n173 VSS.n172 8.7078
R326 VSS.n168 VSS.n167 8.7078
R327 VSS.n164 VSS.n163 8.7078
R328 VSS.n159 VSS.n158 8.7078
R329 VSS.n90 VSS.n87 6.30644
R330 VSS.n30 VSS.t66 5.13332
R331 VSS.n87 VSS.n12 5.10637
R332 VSS.n161 VSS.n157 4.46046
R333 VSS.n132 VSS.t50 4.35415
R334 VSS.n162 VSS.n156 3.78833
R335 VSS.n171 VSS.n154 3.78833
R336 VSS.n144 VSS.n1 3.78833
R337 VSS.n131 VSS.n3 3.78833
R338 VSS.n118 VSS.n5 3.78833
R339 VSS.n111 VSS.n7 3.78833
R340 VSS.n101 VSS.n9 3.78833
R341 VSS.n91 VSS.n11 3.78833
R342 VSS.n79 VSS.n16 3.74137
R343 VSS.n72 VSS.n18 3.74137
R344 VSS.n62 VSS.n20 3.74137
R345 VSS.n54 VSS.n22 3.74137
R346 VSS.n47 VSS.n24 3.74137
R347 VSS.n42 VSS.n26 3.74137
R348 VSS.n35 VSS.n28 3.74137
R349 VSS.n86 VSS.n14 2.6005
R350 VSS.n14 VSS.n13 2.6005
R351 VSS.n85 VSS.n84 2.6005
R352 VSS.n84 VSS.n83 2.6005
R353 VSS.n82 VSS.n81 2.6005
R354 VSS.n81 VSS.n80 2.6005
R355 VSS.n78 VSS.n77 2.6005
R356 VSS.n77 VSS.n76 2.6005
R357 VSS.n75 VSS.n74 2.6005
R358 VSS.n74 VSS.n73 2.6005
R359 VSS.n71 VSS.n70 2.6005
R360 VSS.n70 VSS.n69 2.6005
R361 VSS.n68 VSS.n67 2.6005
R362 VSS.n67 VSS.n66 2.6005
R363 VSS.n65 VSS.n64 2.6005
R364 VSS.n64 VSS.n63 2.6005
R365 VSS.n61 VSS.n60 2.6005
R366 VSS.n60 VSS.n59 2.6005
R367 VSS.n58 VSS.n57 2.6005
R368 VSS.n56 VSS.n55 2.6005
R369 VSS.n53 VSS.n52 2.6005
R370 VSS.n51 VSS.n50 2.6005
R371 VSS.n49 VSS.n48 2.6005
R372 VSS.n46 VSS.n45 2.6005
R373 VSS.n44 VSS.n43 2.6005
R374 VSS.n41 VSS.n40 2.6005
R375 VSS.n39 VSS.n38 2.6005
R376 VSS.n37 VSS.n36 2.6005
R377 VSS.n34 VSS.n33 2.6005
R378 VSS.n32 VSS.n31 2.6005
R379 VSS.n30 VSS.n29 2.6005
R380 VSS.n90 VSS.n89 2.6005
R381 VSS.n89 VSS.n88 2.6005
R382 VSS.n94 VSS.n93 2.6005
R383 VSS.n93 VSS.n92 2.6005
R384 VSS.n97 VSS.n96 2.6005
R385 VSS.n96 VSS.n95 2.6005
R386 VSS.n100 VSS.n99 2.6005
R387 VSS.n99 VSS.n98 2.6005
R388 VSS.n104 VSS.n103 2.6005
R389 VSS.n103 VSS.n102 2.6005
R390 VSS.n107 VSS.n106 2.6005
R391 VSS.n106 VSS.n105 2.6005
R392 VSS.n110 VSS.n109 2.6005
R393 VSS.n109 VSS.n108 2.6005
R394 VSS.n114 VSS.n113 2.6005
R395 VSS.n113 VSS.n112 2.6005
R396 VSS.n117 VSS.n116 2.6005
R397 VSS.n116 VSS.n115 2.6005
R398 VSS.n122 VSS.n121 2.6005
R399 VSS.n121 VSS.n120 2.6005
R400 VSS.n126 VSS.n125 2.6005
R401 VSS.n125 VSS.n124 2.6005
R402 VSS.n130 VSS.n129 2.6005
R403 VSS.n129 VSS.n128 2.6005
R404 VSS.n135 VSS.n134 2.6005
R405 VSS.n134 VSS.n133 2.6005
R406 VSS.n139 VSS.n138 2.6005
R407 VSS.n138 VSS.n137 2.6005
R408 VSS.n143 VSS.n142 2.6005
R409 VSS.n142 VSS.n141 2.6005
R410 VSS.n148 VSS.n147 2.6005
R411 VSS.n147 VSS.n146 2.6005
R412 VSS.n152 VSS.n151 2.6005
R413 VSS.n151 VSS.n150 2.6005
R414 VSS.n175 VSS.n174 2.6005
R415 VSS.n174 VSS.n173 2.6005
R416 VSS.n170 VSS.n169 2.6005
R417 VSS.n169 VSS.n168 2.6005
R418 VSS.n166 VSS.n165 2.6005
R419 VSS.n165 VSS.n164 2.6005
R420 VSS.n160 VSS.n159 2.6005
R421 VSS.n161 VSS.n160 1.76263
R422 VSS.n16 VSS.t79 1.3655
R423 VSS.n16 VSS.n15 1.3655
R424 VSS.n18 VSS.t74 1.3655
R425 VSS.n18 VSS.n17 1.3655
R426 VSS.n20 VSS.t21 1.3655
R427 VSS.n20 VSS.n19 1.3655
R428 VSS.n22 VSS.t77 1.3655
R429 VSS.n22 VSS.n21 1.3655
R430 VSS.n24 VSS.t8 1.3655
R431 VSS.n24 VSS.n23 1.3655
R432 VSS.n26 VSS.t46 1.3655
R433 VSS.n26 VSS.n25 1.3655
R434 VSS.n28 VSS.t3 1.3655
R435 VSS.n28 VSS.n27 1.3655
R436 VSS.n156 VSS.t1 1.3655
R437 VSS.n156 VSS.n155 1.3655
R438 VSS.n154 VSS.t78 1.3655
R439 VSS.n154 VSS.n153 1.3655
R440 VSS.n1 VSS.t37 1.3655
R441 VSS.n1 VSS.n0 1.3655
R442 VSS.n3 VSS.t10 1.3655
R443 VSS.n3 VSS.n2 1.3655
R444 VSS.n5 VSS.t35 1.3655
R445 VSS.n5 VSS.n4 1.3655
R446 VSS.n7 VSS.t42 1.3655
R447 VSS.n7 VSS.n6 1.3655
R448 VSS.n9 VSS.t71 1.3655
R449 VSS.n9 VSS.n8 1.3655
R450 VSS.n11 VSS.t44 1.3655
R451 VSS.n11 VSS.n10 1.3655
R452 VSS.n162 VSS.n161 0.454611
R453 VSS.n86 VSS.n85 0.144885
R454 VSS.n85 VSS.n82 0.144885
R455 VSS.n78 VSS.n75 0.144885
R456 VSS.n71 VSS.n68 0.144885
R457 VSS.n68 VSS.n65 0.144885
R458 VSS.n61 VSS.n58 0.144885
R459 VSS.n58 VSS.n56 0.144885
R460 VSS.n53 VSS.n51 0.144885
R461 VSS.n51 VSS.n49 0.144885
R462 VSS.n46 VSS.n44 0.144885
R463 VSS.n41 VSS.n39 0.144885
R464 VSS.n39 VSS.n37 0.144885
R465 VSS.n34 VSS.n32 0.144885
R466 VSS.n32 VSS.n30 0.144885
R467 VSS.n97 VSS.n94 0.144885
R468 VSS.n100 VSS.n97 0.144885
R469 VSS.n107 VSS.n104 0.144885
R470 VSS.n110 VSS.n107 0.144885
R471 VSS.n117 VSS.n114 0.144885
R472 VSS.n126 VSS.n122 0.144885
R473 VSS.n130 VSS.n126 0.144885
R474 VSS.n139 VSS.n135 0.144885
R475 VSS.n143 VSS.n139 0.144885
R476 VSS.n152 VSS.n148 0.144885
R477 VSS.n170 VSS.n166 0.144885
R478 VSS.n47 VSS.n46 0.141035
R479 VSS.n118 VSS.n117 0.13911
R480 VSS.n171 VSS.n170 0.127559
R481 VSS.n75 VSS.n72 0.125634
R482 VSS.n79 VSS.n78 0.123709
R483 VSS.n166 VSS.n162 0.121783
R484 VSS.n91 VSS.n90 0.116008
R485 VSS.n114 VSS.n111 0.110233
R486 VSS.n44 VSS.n42 0.108307
R487 VSS.n54 VSS.n53 0.100607
R488 VSS.n131 VSS.n130 0.0986818
R489 VSS.n148 VSS.n144 0.087131
R490 VSS.n65 VSS.n62 0.0852059
R491 VSS.n87 VSS.n86 0.0832807
R492 VSS.n35 VSS.n34 0.0775053
R493 VSS VSS.n175 0.0775053
R494 VSS.n101 VSS.n100 0.0755802
R495 VSS.n104 VSS.n101 0.0698048
R496 VSS.n37 VSS.n35 0.0678797
R497 VSS VSS.n152 0.0678797
R498 VSS.n62 VSS.n61 0.0601791
R499 VSS.n144 VSS.n143 0.058254
R500 VSS.n135 VSS.n131 0.0467032
R501 VSS.n56 VSS.n54 0.0447781
R502 VSS.n42 VSS.n41 0.0370775
R503 VSS.n111 VSS.n110 0.0351524
R504 VSS.n94 VSS.n91 0.029377
R505 VSS.n82 VSS.n79 0.0216765
R506 VSS.n72 VSS.n71 0.0197513
R507 VSS.n175 VSS.n171 0.0178262
R508 VSS.n122 VSS.n118 0.0062754
R509 VSS.n49 VSS.n47 0.00435027
R510 IM IM.n30 32.4348
R511 IM.n0 IM.t31 30.5343
R512 IM.n0 IM.t30 18.1775
R513 IM.n1 IM.t28 18.1775
R514 IM.n4 IM.t25 18.1775
R515 IM.n5 IM.t20 18.1775
R516 IM.n8 IM.t16 18.1775
R517 IM.n9 IM.t11 18.1775
R518 IM.n12 IM.t9 18.1775
R519 IM.n13 IM.t7 18.1775
R520 IM.n16 IM.t6 18.1775
R521 IM.n17 IM.t2 18.1775
R522 IM.n20 IM.t19 18.1775
R523 IM.n21 IM.t27 18.1775
R524 IM.n24 IM.t15 18.1775
R525 IM.n25 IM.t12 18.1775
R526 IM.n28 IM.t3 18.1775
R527 IM.n29 IM.t1 18.1775
R528 IM.n2 IM.t29 17.6665
R529 IM.n3 IM.t24 17.6665
R530 IM.n6 IM.t13 17.6665
R531 IM.n7 IM.t18 17.6665
R532 IM.n10 IM.t5 17.6665
R533 IM.n11 IM.t10 17.6665
R534 IM.n14 IM.t0 17.6665
R535 IM.n15 IM.t26 17.6665
R536 IM.n18 IM.t23 17.6665
R537 IM.n19 IM.t21 17.6665
R538 IM.n22 IM.t17 17.6665
R539 IM.n23 IM.t14 17.6665
R540 IM.n26 IM.t8 17.6665
R541 IM.n27 IM.t4 17.6665
R542 IM.n30 IM.t22 17.6665
R543 IM.n1 IM.n0 12.8683
R544 IM.n2 IM.n1 12.8683
R545 IM.n3 IM.n2 12.8683
R546 IM.n4 IM.n3 12.8683
R547 IM.n5 IM.n4 12.8683
R548 IM.n6 IM.n5 12.8683
R549 IM.n7 IM.n6 12.8683
R550 IM.n8 IM.n7 12.8683
R551 IM.n9 IM.n8 12.8683
R552 IM.n10 IM.n9 12.8683
R553 IM.n11 IM.n10 12.8683
R554 IM.n12 IM.n11 12.8683
R555 IM.n13 IM.n12 12.8683
R556 IM.n14 IM.n13 12.8683
R557 IM.n15 IM.n14 12.8683
R558 IM.n16 IM.n15 12.8683
R559 IM.n17 IM.n16 12.8683
R560 IM.n18 IM.n17 12.8683
R561 IM.n19 IM.n18 12.8683
R562 IM.n20 IM.n19 12.8683
R563 IM.n21 IM.n20 12.8683
R564 IM.n22 IM.n21 12.8683
R565 IM.n23 IM.n22 12.8683
R566 IM.n24 IM.n23 12.8683
R567 IM.n25 IM.n24 12.8683
R568 IM.n26 IM.n25 12.8683
R569 IM.n27 IM.n26 12.8683
R570 IM.n28 IM.n27 12.8683
R571 IM.n29 IM.n28 12.8683
R572 IM.n30 IM.n29 12.8683
C0 OUT IM 1.33f
C1 IM SD 0.916f
C2 IM IM_T 1.99f
C3 OUT SD 4.66f
C4 OUT IM_T 0.753f
C5 IM_T SD 1f
.ends

