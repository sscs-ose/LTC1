magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -2234 1019 2234
<< metal1 >>
rect -19 1228 19 1234
rect -19 1202 -13 1228
rect 13 1202 19 1228
rect -19 1174 19 1202
rect -19 1148 -13 1174
rect 13 1148 19 1174
rect -19 1120 19 1148
rect -19 1094 -13 1120
rect 13 1094 19 1120
rect -19 1066 19 1094
rect -19 1040 -13 1066
rect 13 1040 19 1066
rect -19 1012 19 1040
rect -19 986 -13 1012
rect 13 986 19 1012
rect -19 958 19 986
rect -19 932 -13 958
rect 13 932 19 958
rect -19 904 19 932
rect -19 878 -13 904
rect 13 878 19 904
rect -19 850 19 878
rect -19 824 -13 850
rect 13 824 19 850
rect -19 796 19 824
rect -19 770 -13 796
rect 13 770 19 796
rect -19 742 19 770
rect -19 716 -13 742
rect 13 716 19 742
rect -19 688 19 716
rect -19 662 -13 688
rect 13 662 19 688
rect -19 634 19 662
rect -19 608 -13 634
rect 13 608 19 634
rect -19 580 19 608
rect -19 554 -13 580
rect 13 554 19 580
rect -19 526 19 554
rect -19 500 -13 526
rect 13 500 19 526
rect -19 472 19 500
rect -19 446 -13 472
rect 13 446 19 472
rect -19 418 19 446
rect -19 392 -13 418
rect 13 392 19 418
rect -19 364 19 392
rect -19 338 -13 364
rect 13 338 19 364
rect -19 310 19 338
rect -19 284 -13 310
rect 13 284 19 310
rect -19 256 19 284
rect -19 230 -13 256
rect 13 230 19 256
rect -19 202 19 230
rect -19 176 -13 202
rect 13 176 19 202
rect -19 148 19 176
rect -19 122 -13 148
rect 13 122 19 148
rect -19 94 19 122
rect -19 68 -13 94
rect 13 68 19 94
rect -19 40 19 68
rect -19 14 -13 40
rect 13 14 19 40
rect -19 -14 19 14
rect -19 -40 -13 -14
rect 13 -40 19 -14
rect -19 -68 19 -40
rect -19 -94 -13 -68
rect 13 -94 19 -68
rect -19 -122 19 -94
rect -19 -148 -13 -122
rect 13 -148 19 -122
rect -19 -176 19 -148
rect -19 -202 -13 -176
rect 13 -202 19 -176
rect -19 -230 19 -202
rect -19 -256 -13 -230
rect 13 -256 19 -230
rect -19 -284 19 -256
rect -19 -310 -13 -284
rect 13 -310 19 -284
rect -19 -338 19 -310
rect -19 -364 -13 -338
rect 13 -364 19 -338
rect -19 -392 19 -364
rect -19 -418 -13 -392
rect 13 -418 19 -392
rect -19 -446 19 -418
rect -19 -472 -13 -446
rect 13 -472 19 -446
rect -19 -500 19 -472
rect -19 -526 -13 -500
rect 13 -526 19 -500
rect -19 -554 19 -526
rect -19 -580 -13 -554
rect 13 -580 19 -554
rect -19 -608 19 -580
rect -19 -634 -13 -608
rect 13 -634 19 -608
rect -19 -662 19 -634
rect -19 -688 -13 -662
rect 13 -688 19 -662
rect -19 -716 19 -688
rect -19 -742 -13 -716
rect 13 -742 19 -716
rect -19 -770 19 -742
rect -19 -796 -13 -770
rect 13 -796 19 -770
rect -19 -824 19 -796
rect -19 -850 -13 -824
rect 13 -850 19 -824
rect -19 -878 19 -850
rect -19 -904 -13 -878
rect 13 -904 19 -878
rect -19 -932 19 -904
rect -19 -958 -13 -932
rect 13 -958 19 -932
rect -19 -986 19 -958
rect -19 -1012 -13 -986
rect 13 -1012 19 -986
rect -19 -1040 19 -1012
rect -19 -1066 -13 -1040
rect 13 -1066 19 -1040
rect -19 -1094 19 -1066
rect -19 -1120 -13 -1094
rect 13 -1120 19 -1094
rect -19 -1148 19 -1120
rect -19 -1174 -13 -1148
rect 13 -1174 19 -1148
rect -19 -1202 19 -1174
rect -19 -1228 -13 -1202
rect 13 -1228 19 -1202
rect -19 -1234 19 -1228
<< via1 >>
rect -13 1202 13 1228
rect -13 1148 13 1174
rect -13 1094 13 1120
rect -13 1040 13 1066
rect -13 986 13 1012
rect -13 932 13 958
rect -13 878 13 904
rect -13 824 13 850
rect -13 770 13 796
rect -13 716 13 742
rect -13 662 13 688
rect -13 608 13 634
rect -13 554 13 580
rect -13 500 13 526
rect -13 446 13 472
rect -13 392 13 418
rect -13 338 13 364
rect -13 284 13 310
rect -13 230 13 256
rect -13 176 13 202
rect -13 122 13 148
rect -13 68 13 94
rect -13 14 13 40
rect -13 -40 13 -14
rect -13 -94 13 -68
rect -13 -148 13 -122
rect -13 -202 13 -176
rect -13 -256 13 -230
rect -13 -310 13 -284
rect -13 -364 13 -338
rect -13 -418 13 -392
rect -13 -472 13 -446
rect -13 -526 13 -500
rect -13 -580 13 -554
rect -13 -634 13 -608
rect -13 -688 13 -662
rect -13 -742 13 -716
rect -13 -796 13 -770
rect -13 -850 13 -824
rect -13 -904 13 -878
rect -13 -958 13 -932
rect -13 -1012 13 -986
rect -13 -1066 13 -1040
rect -13 -1120 13 -1094
rect -13 -1174 13 -1148
rect -13 -1228 13 -1202
<< metal2 >>
rect -19 1228 19 1234
rect -19 1202 -13 1228
rect 13 1202 19 1228
rect -19 1174 19 1202
rect -19 1148 -13 1174
rect 13 1148 19 1174
rect -19 1120 19 1148
rect -19 1094 -13 1120
rect 13 1094 19 1120
rect -19 1066 19 1094
rect -19 1040 -13 1066
rect 13 1040 19 1066
rect -19 1012 19 1040
rect -19 986 -13 1012
rect 13 986 19 1012
rect -19 958 19 986
rect -19 932 -13 958
rect 13 932 19 958
rect -19 904 19 932
rect -19 878 -13 904
rect 13 878 19 904
rect -19 850 19 878
rect -19 824 -13 850
rect 13 824 19 850
rect -19 796 19 824
rect -19 770 -13 796
rect 13 770 19 796
rect -19 742 19 770
rect -19 716 -13 742
rect 13 716 19 742
rect -19 688 19 716
rect -19 662 -13 688
rect 13 662 19 688
rect -19 634 19 662
rect -19 608 -13 634
rect 13 608 19 634
rect -19 580 19 608
rect -19 554 -13 580
rect 13 554 19 580
rect -19 526 19 554
rect -19 500 -13 526
rect 13 500 19 526
rect -19 472 19 500
rect -19 446 -13 472
rect 13 446 19 472
rect -19 418 19 446
rect -19 392 -13 418
rect 13 392 19 418
rect -19 364 19 392
rect -19 338 -13 364
rect 13 338 19 364
rect -19 310 19 338
rect -19 284 -13 310
rect 13 284 19 310
rect -19 256 19 284
rect -19 230 -13 256
rect 13 230 19 256
rect -19 202 19 230
rect -19 176 -13 202
rect 13 176 19 202
rect -19 148 19 176
rect -19 122 -13 148
rect 13 122 19 148
rect -19 94 19 122
rect -19 68 -13 94
rect 13 68 19 94
rect -19 40 19 68
rect -19 14 -13 40
rect 13 14 19 40
rect -19 -14 19 14
rect -19 -40 -13 -14
rect 13 -40 19 -14
rect -19 -68 19 -40
rect -19 -94 -13 -68
rect 13 -94 19 -68
rect -19 -122 19 -94
rect -19 -148 -13 -122
rect 13 -148 19 -122
rect -19 -176 19 -148
rect -19 -202 -13 -176
rect 13 -202 19 -176
rect -19 -230 19 -202
rect -19 -256 -13 -230
rect 13 -256 19 -230
rect -19 -284 19 -256
rect -19 -310 -13 -284
rect 13 -310 19 -284
rect -19 -338 19 -310
rect -19 -364 -13 -338
rect 13 -364 19 -338
rect -19 -392 19 -364
rect -19 -418 -13 -392
rect 13 -418 19 -392
rect -19 -446 19 -418
rect -19 -472 -13 -446
rect 13 -472 19 -446
rect -19 -500 19 -472
rect -19 -526 -13 -500
rect 13 -526 19 -500
rect -19 -554 19 -526
rect -19 -580 -13 -554
rect 13 -580 19 -554
rect -19 -608 19 -580
rect -19 -634 -13 -608
rect 13 -634 19 -608
rect -19 -662 19 -634
rect -19 -688 -13 -662
rect 13 -688 19 -662
rect -19 -716 19 -688
rect -19 -742 -13 -716
rect 13 -742 19 -716
rect -19 -770 19 -742
rect -19 -796 -13 -770
rect 13 -796 19 -770
rect -19 -824 19 -796
rect -19 -850 -13 -824
rect 13 -850 19 -824
rect -19 -878 19 -850
rect -19 -904 -13 -878
rect 13 -904 19 -878
rect -19 -932 19 -904
rect -19 -958 -13 -932
rect 13 -958 19 -932
rect -19 -986 19 -958
rect -19 -1012 -13 -986
rect 13 -1012 19 -986
rect -19 -1040 19 -1012
rect -19 -1066 -13 -1040
rect 13 -1066 19 -1040
rect -19 -1094 19 -1066
rect -19 -1120 -13 -1094
rect 13 -1120 19 -1094
rect -19 -1148 19 -1120
rect -19 -1174 -13 -1148
rect 13 -1174 19 -1148
rect -19 -1202 19 -1174
rect -19 -1228 -13 -1202
rect 13 -1228 19 -1202
rect -19 -1234 19 -1228
<< end >>
