* NGSPICE file created from NOR_Layout_flat.ext - technology: gf180mcuC

.subckt NOR_Layout_flat IN2 IN1 IN4 IN5 IN6 C1 B1 IN7 IN3 IN8 A1 OUT EN VSS VDD
X0 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t2 Transmission_Gate_Layout_3.VIN.t55 VSS.t112 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1 Transmission_Gate_Layout_15.CLKB EN.t0 VSS.t254 VSS.t253 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X2 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t6 Transmission_Gate_Layout_3.VIN.t109 VDD.t106 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t3 Transmission_Gate_Layout_5.VIN.t56 VSS.t117 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X4 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t2 Transmission_Gate_Layout_3.VIN.t8 VSS.t48 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X5 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t6 Transmission_Gate_Layout_2.VIN.t82 VDD.t73 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLK.t2 VSS.t64 VSS.t63 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X7 OUT Transmission_Gate_Layout_13.CLKB.t6 Transmission_Gate_Layout_13.VIN.t120 VDD.t47 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X8 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t6 Transmission_Gate_Layout_12.VIN.t140 VDD.t55 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X9 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t6 Transmission_Gate_Layout_11.VIN.t36 VDD.t3 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X10 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t2 Transmission_Gate_Layout_1.VIN.t15 VSS.t36 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X11 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t3 Transmission_Gate_Layout_3.VIN.t6 VSS.t55 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X12 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 Transmission_Gate_Layout_13.CLK.t3 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.t2 VDD.t48 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X13 Transmission_Gate_Layout_4.VIN EN.t1 IN7.t35 VSS.t241 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X14 IN2 Transmission_Gate_Layout_18.CLKB.t6 Transmission_Gate_Layout_7.VIN.t0 VDD.t171 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X15 VDD Transmission_Gate_Layout_11.CLK.t4 Transmission_Gate_Layout_8.CLKB.t2 VDD.t185 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X16 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t2 OUT.t72 VSS.t181 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X17 Transmission_Gate_Layout_11.VIN EN.t2 IN4.t47 VSS.t242 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X18 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t7 IN2.t22 VDD.t248 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X19 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t7 Transmission_Gate_Layout_11.VIN.t35 VDD.t144 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X20 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t2 Transmission_Gate_Layout_3.VIN.t68 VSS.t156 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X21 IN7 EN.t3 Transmission_Gate_Layout_4.VIN.t94 VSS.t240 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X22 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t4 Transmission_Gate_Layout_6.VIN.t45 VSS.t43 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X23 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t6 IN3.t23 VDD.t41 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X24 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t6 Transmission_Gate_Layout_9.VIN.t23 VDD.t59 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X25 Transmission_Gate_Layout_4.VIN EN.t4 IN7.t34 VSS.t252 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X26 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t6 Transmission_Gate_Layout_6.VIN.t18 VDD.t83 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X27 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t5 Transmission_Gate_Layout_8.VIN.t71 VSS.t113 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X28 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t7 Transmission_Gate_Layout_9.VOUT.t139 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X29 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT B1.t0 VDD.t150 VDD.t149 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X30 Transmission_Gate_Layout_10.VIN EN.t5 IN3.t47 VSS.t251 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X31 OUT Transmission_Gate_Layout_12.CLKB.t6 Transmission_Gate_Layout_12.VIN.t48 VDD.t92 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X32 Transmission_Gate_Layout_4.VIN EN.t6 IN7.t33 VSS.t237 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X33 IN1 Transmission_Gate_Layout_16.CLKB.t6 Transmission_Gate_Layout_6.VIN.t60 VDD.t241 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X34 Transmission_Gate_Layout_8.VIN EN.t7 IN6.t47 VSS.t238 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X35 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t7 IN3.t22 VDD.t40 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X36 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t7 OUT.t22 VDD.t54 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X37 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t6 IN4.t0 VDD.t154 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X38 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t5 Transmission_Gate_Layout_6.VIN.t44 VSS.t54 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X39 IN7 EN.t8 Transmission_Gate_Layout_4.VIN.t91 VSS.t239 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X40 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t6 Transmission_Gate_Layout_12.VIN.t49 VDD.t62 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X41 IN2 EN.t9 Transmission_Gate_Layout_7.VIN.t48 VSS.t232 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X42 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t7 Transmission_Gate_Layout_3.VIN.t39 VDD.t90 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X43 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t6 Transmission_Gate_Layout_5.VIN.t55 VSS.t117 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X44 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLK.t3 VSS.t57 VSS.t17 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X45 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t6 Transmission_Gate_Layout_5.VIN.t22 VDD.t117 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X46 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t6 Transmission_Gate_Layout_9.VOUT.t49 VDD.t53 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X47 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t6 Transmission_Gate_Layout_10.VIN.t46 VDD.t78 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X48 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t7 Transmission_Gate_Layout_9.VOUT.t50 VDD.t58 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X49 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t7 Transmission_Gate_Layout_1.VIN.t38 VDD.t65 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X50 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t7 Transmission_Gate_Layout_9.VOUT.t21 VSS.t122 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X51 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t7 Transmission_Gate_Layout_13.VIN.t97 VDD.t71 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X52 VSS EN.t10 Transmission_Gate_Layout_18.CLKB.t5 VSS.t233 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X53 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t7 IN4.t1 VDD.t155 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X54 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t8 Transmission_Gate_Layout_7.VIN.t23 VSS.t116 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X55 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t3 Transmission_Gate_Layout_12.VIN.t0 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X56 Transmission_Gate_Layout_10.VIN EN.t11 IN3.t46 VSS.t236 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X57 IN6 Transmission_Gate_Layout_21.CLKB.t6 Transmission_Gate_Layout_8.VIN.t8 VDD.t43 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X58 VDD Transmission_Gate_Layout_12.CLK.t3 Transmission_Gate_Layout_12.CLKB.t2 VDD.t214 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X59 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t6 IN7.t23 VDD.t31 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X60 OUT Transmission_Gate_Layout_12.CLK.t4 Transmission_Gate_Layout_12.VIN.t89 VSS.t182 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X61 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t9 Transmission_Gate_Layout_3.VIN.t54 VSS.t128 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X62 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t10 Transmission_Gate_Layout_11.VIN.t60 VSS.t116 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X63 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t6 Transmission_Gate_Layout_9.VOUT.t100 VSS.t53 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X64 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t11 Transmission_Gate_Layout_2.VIN.t111 VSS.t131 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X65 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t7 Transmission_Gate_Layout_9.VOUT.t73 VDD.t60 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X66 IN2 Transmission_Gate_Layout_18.CLKB.t8 Transmission_Gate_Layout_7.VIN.t26 VDD.t249 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X67 IN8 EN.t12 Transmission_Gate_Layout_5.VIN.t95 VSS.t230 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X68 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t7 Transmission_Gate_Layout_9.VIN.t46 VSS.t52 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X69 IN5 EN.t13 Transmission_Gate_Layout_9.VIN.t59 VSS.t231 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X70 Transmission_Gate_Layout_15.CLKB EN.t14 VDD.t290 VDD.t113 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X71 VSS Transmission_Gate_Layout_9.CLK.t8 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.t3 VSS.t49 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X72 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t9 Transmission_Gate_Layout_3.VIN.t7 VSS.t48 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X73 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t8 Transmission_Gate_Layout_3.VIN.t40 VDD.t85 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X74 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t12 Transmission_Gate_Layout_1.VIN.t109 VSS.t122 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X75 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t4 Transmission_Gate_Layout_1.VIN.t16 VSS.t19 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X76 IN7 EN.t15 Transmission_Gate_Layout_4.VIN.t90 VSS.t228 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X77 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLK.t4 VDD.t49 VDD.t14 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X78 VDD EN.t16 Transmission_Gate_Layout_21.CLKB.t2 VDD.t258 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X79 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t10 Transmission_Gate_Layout_9.VOUT.t99 VSS.t56 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X80 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t8 Transmission_Gate_Layout_11.VIN.t34 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X81 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t7 Transmission_Gate_Layout_2.VIN.t53 VDD.t74 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X82 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t7 OUT.t31 VDD.t91 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X83 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t6 Transmission_Gate_Layout_13.VIN.t39 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X84 IN7 Transmission_Gate_Layout_17.CLKB.t7 Transmission_Gate_Layout_4.VIN.t53 VDD.t29 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X85 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t4 Transmission_Gate_Layout_9.VOUT.t143 VSS.t161 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X86 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t11 Transmission_Gate_Layout_3.VIN.t2 VSS.t46 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X87 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t8 Transmission_Gate_Layout_8.VIN.t45 VDD.t52 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X88 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t8 Transmission_Gate_Layout_9.VOUT.t74 VDD.t61 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X89 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t9 Transmission_Gate_Layout_3.VIN.t41 VDD.t86 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X90 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t13 Transmission_Gate_Layout_2.VIN.t110 VSS.t112 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X91 Transmission_Gate_Layout_3.CLK Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.t2 VSS.t92 VSS.t91 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X92 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t14 Transmission_Gate_Layout_11.VIN.t57 VSS.t123 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X93 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t5 Transmission_Gate_Layout_12.VIN.t18 VSS.t16 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X94 OUT Transmission_Gate_Layout_12.CLKB.t8 Transmission_Gate_Layout_12.VIN.t33 VDD.t97 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X95 IN7 Transmission_Gate_Layout_17.CLKB.t8 Transmission_Gate_Layout_4.VIN.t54 VDD.t30 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X96 IN7 Transmission_Gate_Layout_17.CLKB.t9 Transmission_Gate_Layout_4.VIN.t55 VDD.t33 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X97 VDD Transmission_Gate_Layout_11.CLK.t15 Transmission_Gate_Layout_5.CLKB.t2 VDD.t182 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X98 VDD A1.t0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.t3 VDD.t107 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X99 IN5 EN.t17 Transmission_Gate_Layout_9.VIN.t58 VSS.t229 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X100 IN8 Transmission_Gate_Layout_20.CLKB.t6 Transmission_Gate_Layout_5.VIN.t24 VDD.t131 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X101 VSS Transmission_Gate_Layout_9.CLK.t12 Transmission_Gate_Layout_10.CLKB.t5 VSS.t13 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X102 VDD Transmission_Gate_Layout_1.CLK.t6 Transmission_Gate_Layout_2.CLKB.t4 VDD.t19 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X103 IN6 Transmission_Gate_Layout_21.CLKB.t7 Transmission_Gate_Layout_8.VIN.t9 VDD.t45 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X104 IN6 Transmission_Gate_Layout_21.CLKB.t8 Transmission_Gate_Layout_8.VIN.t10 VDD.t44 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X105 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t13 Transmission_Gate_Layout_10.VIN.t71 VSS.t43 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X106 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t14 Transmission_Gate_Layout_9.VOUT.t98 VSS.t70 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X107 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t5 Transmission_Gate_Layout_13.VIN.t0 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X108 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t8 Transmission_Gate_Layout_9.VOUT.t138 VDD.t57 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X109 Transmission_Gate_Layout_9.VIN EN.t18 IN5.t21 VSS.t224 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X110 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t8 IN3.t21 VDD.t41 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X111 Transmission_Gate_Layout_16.CLKB EN.t19 VSS.t226 VSS.t225 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X112 IN5 EN.t20 Transmission_Gate_Layout_9.VIN.t57 VSS.t227 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X113 OUT Transmission_Gate_Layout_12.CLKB.t9 Transmission_Gate_Layout_12.VIN.t34 VDD.t92 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X114 Transmission_Gate_Layout_6.VIN EN.t21 IN1.t47 VSS.t222 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X115 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_9.CLK.t15 VDD.t123 VDD.t122 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X116 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t6 Transmission_Gate_Layout_13.VIN.t1 VSS.t4 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X117 Transmission_Gate_Layout_9.VIN EN.t22 IN5.t19 VSS.t223 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X118 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t5 OUT.t71 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X119 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t16 Transmission_Gate_Layout_8.VIN.t69 VSS.t117 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X120 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t8 Transmission_Gate_Layout_10.VIN.t24 VDD.t72 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X121 Transmission_Gate_Layout_1.CLK Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.t2 VSS.t102 VSS.t101 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X122 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t9 Transmission_Gate_Layout_9.VIN.t20 VDD.t64 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X123 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t9 IN2.t20 VDD.t250 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X124 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.t2 VSS.t108 VSS.t85 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X125 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t7 IN8.t1 VDD.t132 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X126 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t17 Transmission_Gate_Layout_9.VOUT.t20 VSS.t133 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X127 IN6 EN.t23 Transmission_Gate_Layout_8.VIN.t95 VSS.t221 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X128 OUT Transmission_Gate_Layout_13.CLK.t6 Transmission_Gate_Layout_13.VIN.t43 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X129 IN3 Transmission_Gate_Layout_14.CLKB.t9 Transmission_Gate_Layout_10.VIN.t20 VDD.t42 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X130 IN4 Transmission_Gate_Layout_19.CLKB.t8 Transmission_Gate_Layout_11.VIN.t2 VDD.t156 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X131 Transmission_Gate_Layout_6.VIN EN.t24 IN1.t46 VSS.t219 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X132 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t10 OUT.t34 VDD.t98 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X133 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t8 Transmission_Gate_Layout_1.VIN.t39 VDD.t65 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X134 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t16 Transmission_Gate_Layout_6.VIN.t41 VSS.t54 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X135 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t7 Transmission_Gate_Layout_13.VIN.t31 VSS.t20 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X136 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t10 Transmission_Gate_Layout_6.VIN.t22 VDD.t88 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X137 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t7 Transmission_Gate_Layout_9.VOUT.t141 VSS.t163 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X138 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t18 Transmission_Gate_Layout_2.VIN.t109 VSS.t127 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X139 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t17 Transmission_Gate_Layout_2.VIN.t143 VSS.t48 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X140 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t8 Transmission_Gate_Layout_13.VIN.t96 VDD.t77 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X141 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t8 IN8.t2 VDD.t133 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X142 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t9 IN6.t11 VDD.t46 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X143 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t8 Transmission_Gate_Layout_9.VOUT.t142 VSS.t162 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X144 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t7 Transmission_Gate_Layout_13.VIN.t124 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X145 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t10 IN6.t12 VDD.t0 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X146 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t18 Transmission_Gate_Layout_6.VIN.t40 VSS.t47 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X147 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t6 IN5.t47 VDD.t297 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X148 Transmission_Gate_Layout_10.VIN EN.t25 IN3.t45 VSS.t220 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X149 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t11 Transmission_Gate_Layout_6.VIN.t23 VDD.t89 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X150 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t19 Transmission_Gate_Layout_2.VIN.t108 VSS.t131 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X151 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLK.t19 VDD.t121 VDD.t24 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X152 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t8 Transmission_Gate_Layout_13.VIN.t125 VDD.t162 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X153 IN8 EN.t26 Transmission_Gate_Layout_5.VIN.t94 VSS.t221 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X154 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t20 Transmission_Gate_Layout_2.VIN.t142 VSS.t48 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X155 IN8 Transmission_Gate_Layout_20.CLKB.t9 Transmission_Gate_Layout_5.VIN.t27 VDD.t134 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X156 OUT Transmission_Gate_Layout_13.CLK.t7 Transmission_Gate_Layout_13.VIN.t44 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X157 IN2 Transmission_Gate_Layout_18.CLKB.t10 Transmission_Gate_Layout_7.VIN.t28 VDD.t171 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X158 OUT Transmission_Gate_Layout_13.CLKB.t8 Transmission_Gate_Layout_13.VIN.t2 VDD.t12 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X159 IN1 EN.t27 Transmission_Gate_Layout_6.VIN.t83 VSS.t216 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X160 IN5 Transmission_Gate_Layout_15.CLKB.t7 Transmission_Gate_Layout_9.VIN.t87 VDD.t294 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X161 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t20 Transmission_Gate_Layout_3.VIN.t53 VSS.t127 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X162 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t8 Transmission_Gate_Layout_1.VIN.t18 VSS.t24 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X163 Transmission_Gate_Layout_6.VIN EN.t28 IN1.t44 VSS.t217 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X164 IN8 EN.t29 Transmission_Gate_Layout_5.VIN.t93 VSS.t218 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X165 VSS Transmission_Gate_Layout_12.CLK.t5 Transmission_Gate_Layout_12.CLKB.t5 VSS.t183 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X166 IN8 Transmission_Gate_Layout_20.CLKB.t10 Transmission_Gate_Layout_5.VIN.t28 VDD.t135 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X167 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t9 Transmission_Gate_Layout_11.VIN.t33 VDD.t5 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X168 IN1 EN.t30 Transmission_Gate_Layout_6.VIN.t82 VSS.t214 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X169 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLK.t21 VDD.t195 VDD.t180 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X170 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t9 Transmission_Gate_Layout_2.VIN.t23 VSS.t25 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X171 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t9 Transmission_Gate_Layout_13.VIN.t143 VSS.t165 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X172 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t9 Transmission_Gate_Layout_13.VIN.t126 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X173 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t22 Transmission_Gate_Layout_8.VIN.t67 VSS.t114 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X174 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t9 IN4.t3 VDD.t154 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X175 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t21 Transmission_Gate_Layout_2.VIN.t141 VSS.t46 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X176 Transmission_Gate_Layout_16.CLKB EN.t31 VDD.t287 VDD.t85 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X177 IN5 Transmission_Gate_Layout_15.CLKB.t8 Transmission_Gate_Layout_9.VIN.t86 VDD.t293 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X178 OUT Transmission_Gate_Layout_12.CLKB.t11 Transmission_Gate_Layout_12.VIN.t36 VDD.t94 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X179 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t10 Transmission_Gate_Layout_3.VIN.t92 VDD.t144 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X180 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t11 IN8.t5 VDD.t136 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X181 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t23 Transmission_Gate_Layout_7.VIN.t20 VSS.t126 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X182 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t9 Transmission_Gate_Layout_10.VIN.t25 VDD.t73 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X183 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t22 Transmission_Gate_Layout_1.VIN.t84 VSS.t56 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X184 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t9 Transmission_Gate_Layout_9.VOUT.t52 VDD.t55 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X185 IN5 EN.t32 Transmission_Gate_Layout_9.VIN.t56 VSS.t215 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X186 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t24 Transmission_Gate_Layout_11.VIN.t54 VSS.t130 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X187 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t11 Transmission_Gate_Layout_3.VIN.t93 VDD.t3 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X188 VDD Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.t3 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.t1 VDD.t163 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X189 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t25 Transmission_Gate_Layout_1.VIN.t108 VSS.t133 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X190 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t23 Transmission_Gate_Layout_4.VIN.t51 VSS.t89 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X191 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t10 Transmission_Gate_Layout_9.VOUT.t53 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X192 Transmission_Gate_Layout_5.VIN EN.t33 IN8.t44 VSS.t265 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X193 IN1 Transmission_Gate_Layout_16.CLKB.t7 Transmission_Gate_Layout_6.VIN.t61 VDD.t242 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X194 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t9 OUT.t20 VDD.t13 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X195 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t9 Transmission_Gate_Layout_9.VOUT.t137 VDD.t57 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X196 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t12 IN8.t6 VDD.t137 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X197 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t24 Transmission_Gate_Layout_6.VIN.t39 VSS.t43 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X198 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t9 Transmission_Gate_Layout_2.VIN.t81 VDD.t78 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X199 OUT Transmission_Gate_Layout_12.CLK.t6 Transmission_Gate_Layout_12.VIN.t90 VSS.t186 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X200 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t10 Transmission_Gate_Layout_12.VIN.t139 VDD.t58 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X201 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t10 Transmission_Gate_Layout_3.VIN.t80 VSS.t170 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X202 Transmission_Gate_Layout_15.CLKB EN.t34 VDD.t286 VDD.t113 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X203 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t25 Transmission_Gate_Layout_6.VIN.t38 VSS.t90 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X204 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT Transmission_Gate_Layout_13.CLK.t8 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.t0 VDD.t50 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X205 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t10 Transmission_Gate_Layout_9.VOUT.t76 VDD.t62 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X206 IN3 Transmission_Gate_Layout_14.CLKB.t10 Transmission_Gate_Layout_10.VIN.t19 VDD.t43 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X207 IN5 Transmission_Gate_Layout_15.CLKB.t9 Transmission_Gate_Layout_9.VIN.t85 VDD.t296 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X208 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_11.CLK.t26 VSS.t149 VSS.t118 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X209 OUT Transmission_Gate_Layout_12.CLK.t7 Transmission_Gate_Layout_12.VIN.t91 VSS.t187 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X210 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t27 Transmission_Gate_Layout_9.VOUT.t19 VSS.t133 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X211 VSS Transmission_Gate_Layout_3.CLK.t11 Transmission_Gate_Layout_0.CLKB.t4 VSS.t166 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X212 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t11 Transmission_Gate_Layout_12.VIN.t138 VDD.t53 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X213 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_11.CLK.t28 VDD.t194 VDD.t178 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X214 OUT Transmission_Gate_Layout_13.CLK.t9 Transmission_Gate_Layout_13.VIN.t45 VSS.t8 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X215 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t26 Transmission_Gate_Layout_3.VIN.t11 VSS.t62 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X216 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t27 Transmission_Gate_Layout_10.VIN.t67 VSS.t54 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X217 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t10 Transmission_Gate_Layout_2.VIN.t32 VDD.t71 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X218 VSS Transmission_Gate_Layout_1.CLK.t10 Transmission_Gate_Layout_2.CLKB.t5 VSS.t21 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X219 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t11 Transmission_Gate_Layout_1.VIN.t19 VSS.t27 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X220 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t28 Transmission_Gate_Layout_2.VIN.t140 VSS.t62 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X221 IN7 Transmission_Gate_Layout_17.CLKB.t10 Transmission_Gate_Layout_4.VIN.t0 VDD.t29 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X222 IN8 Transmission_Gate_Layout_20.CLKB.t13 Transmission_Gate_Layout_5.VIN.t31 VDD.t138 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X223 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 Transmission_Gate_Layout_3.CLK.t12 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.t0 VDD.t48 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X224 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t8 IN1.t21 VDD.t246 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X225 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t7 Transmission_Gate_Layout_5.VIN.t23 VDD.t120 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X226 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t29 Transmission_Gate_Layout_3.VIN.t10 VSS.t46 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X227 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t12 Transmission_Gate_Layout_2.VIN.t24 VSS.t32 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X228 Transmission_Gate_Layout_9.VIN EN.t35 IN5.t17 VSS.t299 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X229 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_11.CLK.t29 VSS.t148 VSS.t118 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X230 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t11 Transmission_Gate_Layout_8.VIN.t42 VDD.t10 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X231 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t13 Transmission_Gate_Layout_12.VIN.t85 VSS.t171 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X232 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t30 Transmission_Gate_Layout_3.VIN.t52 VSS.t131 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X233 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t30 Transmission_Gate_Layout_10.VIN.t65 VSS.t47 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X234 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t12 Transmission_Gate_Layout_13.VIN.t129 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X235 VDD EN.t36 Transmission_Gate_Layout_14.CLKB.t2 VDD.t258 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X236 IN3 EN.t37 Transmission_Gate_Layout_10.VIN.t92 VSS.t276 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X237 OUT Transmission_Gate_Layout_12.CLKB.t12 Transmission_Gate_Layout_12.VIN.t37 VDD.t95 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X238 IN7 Transmission_Gate_Layout_17.CLKB.t11 Transmission_Gate_Layout_4.VIN.t1 VDD.t30 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X239 IN8 EN.t38 Transmission_Gate_Layout_5.VIN.t92 VSS.t218 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X240 IN6 EN.t39 Transmission_Gate_Layout_8.VIN.t94 VSS.t221 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X241 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t10 Transmission_Gate_Layout_13.VIN.t94 VDD.t74 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X242 VSS Transmission_Gate_Layout_9.CLK.t31 Transmission_Gate_Layout_6.CLKB.t5 VSS.t13 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X243 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t11 Transmission_Gate_Layout_9.VOUT.t77 VDD.t63 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X244 Transmission_Gate_Layout_9.VIN EN.t40 IN5.t16 VSS.t296 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X245 IN3 EN.t41 Transmission_Gate_Layout_10.VIN.t91 VSS.t280 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X246 VDD Transmission_Gate_Layout_9.CLK.t32 Transmission_Gate_Layout_6.CLKB.t2 VDD.t227 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X247 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t11 Transmission_Gate_Layout_2.VIN.t33 VDD.t75 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X248 Transmission_Gate_Layout_19.CLKB EN.t42 VSS.t320 VSS.t292 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X249 Transmission_Gate_Layout_5.VIN EN.t43 IN8.t42 VSS.t238 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X250 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t31 Transmission_Gate_Layout_11.VIN.t53 VSS.t123 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X251 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t8 OUT.t76 VSS.t188 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X252 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t13 Transmission_Gate_Layout_3.VIN.t95 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X253 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t32 Transmission_Gate_Layout_7.VIN.t18 VSS.t130 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X254 IN6 EN.t44 Transmission_Gate_Layout_8.VIN.t93 VSS.t218 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X255 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t13 Transmission_Gate_Layout_13.VIN.t34 VSS.t26 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X256 Transmission_Gate_Layout_7.VIN EN.t45 IN2.t46 VSS.t273 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X257 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t10 IN5.t43 VDD.t295 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X258 Transmission_Gate_Layout_5.VIN EN.t46 IN8.t41 VSS.t289 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X259 VSS EN.t47 Transmission_Gate_Layout_20.CLKB.t5 VSS.t283 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X260 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t33 Transmission_Gate_Layout_1.VIN.t36 VSS.t82 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X261 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t14 Transmission_Gate_Layout_12.VIN.t21 VSS.t31 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X262 VSS EN.t48 Transmission_Gate_Layout_14.CLKB.t5 VSS.t268 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X263 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t10 OUT.t19 VDD.t56 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X264 IN2 EN.t49 Transmission_Gate_Layout_7.VIN.t94 VSS.t271 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X265 IN4 EN.t50 Transmission_Gate_Layout_11.VIN.t84 VSS.t264 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X266 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t6 Transmission_Gate_Layout_4.VIN.t56 VDD.t32 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X267 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t34 Transmission_Gate_Layout_9.VOUT.t97 VSS.t70 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X268 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t9 Transmission_Gate_Layout_12.VIN.t52 VDD.t61 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X269 Transmission_Gate_Layout_17.CLKB EN.t51 VSS.t315 VSS.t294 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X270 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t33 Transmission_Gate_Layout_5.VIN.t54 VSS.t113 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X271 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t10 Transmission_Gate_Layout_2.VIN.t59 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X272 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t15 Transmission_Gate_Layout_13.VIN.t35 VSS.t33 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X273 OUT Transmission_Gate_Layout_12.CLK.t9 Transmission_Gate_Layout_12.VIN.t93 VSS.t189 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X274 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t35 Transmission_Gate_Layout_1.VIN.t24 VSS.t70 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X275 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t14 Transmission_Gate_Layout_13.VIN.t112 VSS.t164 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X276 OUT Transmission_Gate_Layout_12.CLKB.t13 Transmission_Gate_Layout_12.VIN.t38 VDD.t94 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X277 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t14 Transmission_Gate_Layout_3.VIN.t96 VDD.t144 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X278 IN3 Transmission_Gate_Layout_14.CLKB.t11 Transmission_Gate_Layout_10.VIN.t18 VDD.t44 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X279 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t11 IN5.t42 VDD.t182 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X280 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t8 Transmission_Gate_Layout_1.VIN.t63 VDD.t113 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X281 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t34 Transmission_Gate_Layout_1.VIN.t106 VSS.t125 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X282 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t14 OUT.t38 VDD.t96 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X283 Transmission_Gate_Layout_19.CLKB EN.t52 VDD.t283 VDD.t131 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X284 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t12 Transmission_Gate_Layout_9.VIN.t17 VDD.t66 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X285 VDD EN.t53 Transmission_Gate_Layout_20.CLKB.t2 VDD.t161 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X286 IN6 EN.t54 Transmission_Gate_Layout_8.VIN.t92 VSS.t218 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X287 OUT Transmission_Gate_Layout_13.CLK.t10 Transmission_Gate_Layout_13.VIN.t46 VSS.t9 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X288 IN3 Transmission_Gate_Layout_14.CLKB.t12 Transmission_Gate_Layout_10.VIN.t17 VDD.t45 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X289 IN1 EN.t55 Transmission_Gate_Layout_6.VIN.t81 VSS.t288 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X290 Transmission_Gate_Layout_8.VIN EN.t56 IN6.t42 VSS.t265 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X291 VSS Transmission_Gate_Layout_11.CLK.t35 Transmission_Gate_Layout_8.CLKB.t5 VSS.t120 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X292 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t12 Transmission_Gate_Layout_10.VIN.t28 VDD.t76 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X293 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t15 OUT.t39 VDD.t93 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X294 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t7 Transmission_Gate_Layout_7.VIN.t65 VDD.t100 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X295 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t36 Transmission_Gate_Layout_4.VIN.t48 VSS.t81 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X296 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t11 IN6.t13 VDD.t41 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X297 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t7 Transmission_Gate_Layout_1.VIN.t113 VDD.t29 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X298 IN6 EN.t57 Transmission_Gate_Layout_8.VIN.t91 VSS.t279 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X299 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t15 Transmission_Gate_Layout_9.VOUT.t47 VSS.t173 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X300 IN2 EN.t58 Transmission_Gate_Layout_7.VIN.t93 VSS.t263 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X301 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t12 Transmission_Gate_Layout_8.VIN.t41 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X302 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t11 Transmission_Gate_Layout_2.VIN.t80 VDD.t78 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X303 Transmission_Gate_Layout_6.VIN EN.t59 IN1.t41 VSS.t262 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X304 Transmission_Gate_Layout_17.CLKB EN.t60 VDD.t280 VDD.t122 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X305 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t12 Transmission_Gate_Layout_12.VIN.t137 VDD.t58 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X306 IN1 EN.t61 Transmission_Gate_Layout_6.VIN.t80 VSS.t286 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X307 IN3 EN.t62 Transmission_Gate_Layout_10.VIN.t90 VSS.t258 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X308 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t12 IN6.t14 VDD.t40 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X309 IN3 Transmission_Gate_Layout_14.CLKB.t13 Transmission_Gate_Layout_10.VIN.t16 VDD.t43 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X310 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLK.t36 VSS.t145 VSS.t118 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X311 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t37 Transmission_Gate_Layout_9.VIN.t42 VSS.t81 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X312 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t10 Transmission_Gate_Layout_1.VIN.t41 VDD.t64 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X313 Transmission_Gate_Layout_11.VIN EN.t63 IN4.t45 VSS.t282 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X314 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t8 Transmission_Gate_Layout_1.VIN.t114 VDD.t30 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X315 VSS Transmission_Gate_Layout_13.CLK.t11 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.t0 VSS.t65 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X316 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t10 OUT.t78 VSS.t190 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X317 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLK.t38 VSS.t80 VSS.t78 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X318 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t16 Transmission_Gate_Layout_3.VIN.t82 VSS.t169 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X319 Transmission_Gate_Layout_11.VIN EN.t64 IN4.t44 VSS.t259 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X320 IN5 Transmission_Gate_Layout_15.CLKB.t12 Transmission_Gate_Layout_9.VIN.t84 VDD.t294 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X321 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t13 Transmission_Gate_Layout_9.VIN.t16 VDD.t65 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X322 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t14 IN3.t20 VDD.t0 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X323 IN1 Transmission_Gate_Layout_16.CLKB.t9 Transmission_Gate_Layout_6.VIN.t63 VDD.t243 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X324 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t9 Transmission_Gate_Layout_1.VIN.t115 VDD.t34 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X325 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t37 Transmission_Gate_Layout_3.VIN.t51 VSS.t131 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X326 IN4 EN.t65 Transmission_Gate_Layout_11.VIN.t83 VSS.t260 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X327 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t8 Transmission_Gate_Layout_3.VIN.t113 VDD.t105 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X328 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t9 Transmission_Gate_Layout_1.VIN.t64 VDD.t115 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X329 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t39 Transmission_Gate_Layout_4.VIN.t47 VSS.t52 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X330 Transmission_Gate_Layout_8.VIN EN.t66 IN6.t40 VSS.t289 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X331 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t12 OUT.t66 VSS.t10 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X332 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t15 IN3.t19 VDD.t46 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X333 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t9 Transmission_Gate_Layout_3.VIN.t126 VDD.t106 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X334 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t10 Transmission_Gate_Layout_4.VIN.t60 VDD.t31 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X335 Transmission_Gate_Layout_16.CLKB EN.t67 VDD.t279 VDD.t85 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X336 IN5 Transmission_Gate_Layout_15.CLKB.t13 Transmission_Gate_Layout_9.VIN.t83 VDD.t293 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X337 IN8 EN.t68 Transmission_Gate_Layout_5.VIN.t91 VSS.t279 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X338 VDD EN.t69 Transmission_Gate_Layout_14.CLKB.t1 VDD.t258 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X339 IN2 Transmission_Gate_Layout_18.CLKB.t11 Transmission_Gate_Layout_7.VIN.t29 VDD.t178 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X340 IN1 Transmission_Gate_Layout_16.CLKB.t10 Transmission_Gate_Layout_6.VIN.t64 VDD.t240 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X341 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t16 Transmission_Gate_Layout_2.VIN.t27 VSS.t35 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X342 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t10 Transmission_Gate_Layout_7.VIN.t67 VDD.t104 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X343 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLK.t40 VSS.t79 VSS.t78 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X344 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLK.t17 VDD.t39 VDD.t24 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X345 Transmission_Gate_Layout_7.VIN EN.t70 IN2.t43 VSS.t255 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X346 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t10 Transmission_Gate_Layout_1.VIN.t65 VDD.t116 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X347 VDD Transmission_Gate_Layout_11.CLK.t38 Transmission_Gate_Layout_8.CLKB.t1 VDD.t185 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X348 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t12 Transmission_Gate_Layout_13.VIN.t92 VDD.t74 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X349 OUT Transmission_Gate_Layout_12.CLKB.t16 Transmission_Gate_Layout_12.VIN.t41 VDD.t95 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X350 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t10 IN4.t4 VDD.t157 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X351 Transmission_Gate_Layout_5.VIN EN.t71 IN8.t39 VSS.t265 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X352 VSS Transmission_Gate_Layout_9.CLK.t41 Transmission_Gate_Layout_10.CLKB.t4 VSS.t13 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X353 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t17 Transmission_Gate_Layout_12.VIN.t87 VSS.t172 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X354 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t15 Transmission_Gate_Layout_3.VIN.t97 VDD.t5 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X355 Transmission_Gate_Layout_10.VIN EN.t72 IN3.t44 VSS.t257 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X356 VDD C1.t0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.t3 VDD.t200 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X357 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t14 Transmission_Gate_Layout_9.VIN.t15 VDD.t59 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X358 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t12 Transmission_Gate_Layout_6.VIN.t0 VDD.t83 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X359 Transmission_Gate_Layout_5.VIN EN.t73 IN8.t38 VSS.t275 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X360 Transmission_Gate_Layout_15.CLKB EN.t74 VSS.t314 VSS.t253 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X361 VSS Transmission_Gate_Layout_3.CLK.t18 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.t2 VSS.t97 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X362 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t39 Transmission_Gate_Layout_7.VIN.t16 VSS.t123 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X363 IN4 EN.t75 Transmission_Gate_Layout_11.VIN.t82 VSS.t281 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X364 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t11 Transmission_Gate_Layout_7.VIN.t79 VDD.t103 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X365 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t11 Transmission_Gate_Layout_2.VIN.t60 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X366 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t11 Transmission_Gate_Layout_5.VIN.t5 VDD.t117 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X367 Transmission_Gate_Layout_11.VIN EN.t76 IN4.t41 VSS.t242 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X368 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t11 IN1.t18 VDD.t227 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X369 IN7 EN.t77 Transmission_Gate_Layout_4.VIN.t89 VSS.t240 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X370 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t19 Transmission_Gate_Layout_3.VIN.t83 VSS.t156 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X371 IN3 Transmission_Gate_Layout_14.CLKB.t16 Transmission_Gate_Layout_10.VIN.t13 VDD.t44 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X372 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t13 Transmission_Gate_Layout_12.VIN.t136 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X373 IN4 EN.t78 Transmission_Gate_Layout_11.VIN.t81 VSS.t277 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X374 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t42 Transmission_Gate_Layout_1.VIN.t87 VSS.t70 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X375 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t40 Transmission_Gate_Layout_7.VIN.t15 VSS.t123 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X376 Transmission_Gate_Layout_4.VIN EN.t79 IN7.t32 VSS.t252 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X377 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t11 Transmission_Gate_Layout_1.VIN.t117 VDD.t33 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X378 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.t2 VSS.t100 VSS.t99 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X379 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t20 Transmission_Gate_Layout_3.VIN.t69 VSS.t157 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X380 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t17 OUT.t41 VDD.t96 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X381 VDD Transmission_Gate_Layout_9.CLK.t43 Transmission_Gate_Layout_10.CLKB.t2 VDD.t19 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X382 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t41 Transmission_Gate_Layout_3.VIN.t50 VSS.t112 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X383 Transmission_Gate_Layout_8.VIN EN.t80 IN6.t39 VSS.t289 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X384 IN7 EN.t81 Transmission_Gate_Layout_4.VIN.t87 VSS.t239 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X385 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t12 Transmission_Gate_Layout_3.VIN.t111 VDD.t102 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X386 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t12 Transmission_Gate_Layout_5.VIN.t6 VDD.t118 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X387 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t15 Transmission_Gate_Layout_9.VOUT.t110 VDD.t60 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X388 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLK.t21 VSS.t159 VSS.t158 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X389 IN2 EN.t82 Transmission_Gate_Layout_7.VIN.t90 VSS.t232 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X390 IN4 Transmission_Gate_Layout_19.CLKB.t11 Transmission_Gate_Layout_11.VIN.t5 VDD.t158 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X391 IN4 Transmission_Gate_Layout_19.CLKB.t12 Transmission_Gate_Layout_11.VIN.t6 VDD.t159 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X392 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t12 IN1.t17 VDD.t246 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X393 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t12 Transmission_Gate_Layout_4.VIN.t62 VDD.t35 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X394 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t13 Transmission_Gate_Layout_8.VIN.t40 VDD.t57 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X395 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t13 OUT.t65 VSS.t12 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X396 Transmission_Gate_Layout_7.VIN EN.t83 IN2.t41 VSS.t278 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X397 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t13 Transmission_Gate_Layout_6.VIN.t1 VDD.t84 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X398 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t42 Transmission_Gate_Layout_1.VIN.t105 VSS.t133 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X399 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT Transmission_Gate_Layout_11.CLK.t43 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.t1 VDD.t27 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X400 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t13 Transmission_Gate_Layout_1.VIN.t68 VDD.t119 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X401 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t18 Transmission_Gate_Layout_12.VIN.t22 VSS.t34 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X402 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t14 Transmission_Gate_Layout_3.VIN.t15 VDD.t85 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X403 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t19 Transmission_Gate_Layout_2.VIN.t28 VSS.t38 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X404 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t22 Transmission_Gate_Layout_12.VIN.t73 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X405 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t23 Transmission_Gate_Layout_12.VIN.t74 VSS.t160 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X406 IN4 Transmission_Gate_Layout_19.CLKB.t13 Transmission_Gate_Layout_11.VIN.t7 VDD.t160 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X407 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t13 Transmission_Gate_Layout_4.VIN.t63 VDD.t36 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X408 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t12 IN2.t17 VDD.t248 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X409 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t44 Transmission_Gate_Layout_3.VIN.t49 VSS.t127 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X410 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t13 Transmission_Gate_Layout_3.VIN.t110 VDD.t101 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X411 IN6 Transmission_Gate_Layout_21.CLKB.t13 Transmission_Gate_Layout_8.VIN.t15 VDD.t42 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X412 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t14 Transmission_Gate_Layout_9.VOUT.t132 VDD.t10 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X413 IN3 EN.t84 Transmission_Gate_Layout_10.VIN.t88 VSS.t256 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X414 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t17 IN3.t18 VDD.t0 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X415 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t45 Transmission_Gate_Layout_2.VIN.t107 VSS.t131 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X416 VSS Transmission_Gate_Layout_11.CLK.t46 Transmission_Gate_Layout_5.CLKB.t5 VSS.t120 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X417 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t11 OUT.t79 VSS.t191 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X418 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t44 Transmission_Gate_Layout_9.VIN.t41 VSS.t52 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X419 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t14 Transmission_Gate_Layout_8.VIN.t39 VDD.t52 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X420 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t13 IN2.t16 VDD.t251 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X421 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t15 Transmission_Gate_Layout_3.VIN.t16 VDD.t86 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X422 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t14 Transmission_Gate_Layout_7.VIN.t64 VDD.t99 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X423 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t13 Transmission_Gate_Layout_2.VIN.t35 VDD.t77 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X424 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t14 OUT.t64 VSS.t11 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X425 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t11 Transmission_Gate_Layout_12.VIN.t54 VDD.t63 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X426 IN7 EN.t85 Transmission_Gate_Layout_4.VIN.t86 VSS.t228 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X427 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t12 Transmission_Gate_Layout_2.VIN.t61 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X428 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t20 Transmission_Gate_Layout_12.VIN.t23 VSS.t39 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X429 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t11 OUT.t18 VDD.t17 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X430 Transmission_Gate_Layout_4.VIN EN.t86 IN7.t31 VSS.t274 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X431 IN6 EN.t87 Transmission_Gate_Layout_8.VIN.t90 VSS.t230 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X432 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.t3 VDD.t140 VDD.t139 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X433 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t13 Transmission_Gate_Layout_2.VIN.t62 VDD.t162 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X434 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t14 IN4.t8 VDD.t155 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X435 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t21 Transmission_Gate_Layout_1.VIN.t23 VSS.t36 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X436 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t16 Transmission_Gate_Layout_3.VIN.t98 VDD.t5 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X437 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t22 Transmission_Gate_Layout_13.VIN.t38 VSS.t40 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X438 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t24 Transmission_Gate_Layout_9.VOUT.t36 VSS.t161 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X439 IN2 EN.t88 Transmission_Gate_Layout_7.VIN.t89 VSS.t272 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X440 Transmission_Gate_Layout_3.CLK Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.t3 VDD.t125 VDD.t124 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X441 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t47 Transmission_Gate_Layout_5.VIN.t53 VSS.t114 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X442 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT Transmission_Gate_Layout_3.CLK.t25 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.t0 VDD.t50 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X443 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t12 IN7.t2 VDD.t31 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X444 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t16 Transmission_Gate_Layout_3.VIN.t17 VDD.t87 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X445 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t45 Transmission_Gate_Layout_2.VIN.t139 VSS.t55 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X446 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t13 Transmission_Gate_Layout_13.VIN.t91 VDD.t75 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X447 Transmission_Gate_Layout_11.VIN EN.t89 IN4.t39 VSS.t267 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X448 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 Transmission_Gate_Layout_11.CLK.t48 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.t2 VDD.t28 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X449 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t14 Transmission_Gate_Layout_5.VIN.t8 VDD.t114 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X450 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1 Transmission_Gate_Layout_12.CLK.t12 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.t1 VDD.t217 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X451 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t17 Transmission_Gate_Layout_13.VIN.t134 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X452 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t49 Transmission_Gate_Layout_11.VIN.t51 VSS.t123 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X453 Transmission_Gate_Layout_10.VIN EN.t90 IN3.t43 VSS.t251 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X454 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t23 Transmission_Gate_Layout_12.VIN.t1 VSS.t16 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X455 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t46 Transmission_Gate_Layout_6.VIN.t35 VSS.t47 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X456 IN2 Transmission_Gate_Layout_18.CLKB.t14 Transmission_Gate_Layout_7.VIN.t32 VDD.t249 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X457 VSS Transmission_Gate_Layout_9.CLK.t47 Transmission_Gate_Layout_6.CLKB.t4 VSS.t13 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X458 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t14 Transmission_Gate_Layout_10.VIN.t30 VDD.t72 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X459 IN5 EN.t91 Transmission_Gate_Layout_9.VIN.t55 VSS.t229 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X460 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t13 IN7.t3 VDD.t32 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X461 OUT Transmission_Gate_Layout_13.CLKB.t12 Transmission_Gate_Layout_13.VIN.t40 VDD.t47 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X462 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 A1.t1 VDD.t111 VDD.t110 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X463 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLK.t24 VSS.t18 VSS.t17 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X464 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t48 Transmission_Gate_Layout_9.VOUT.t96 VSS.t70 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X465 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t14 Transmission_Gate_Layout_11.VIN.t28 VDD.t144 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X466 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t15 Transmission_Gate_Layout_12.VIN.t135 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X467 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLK.t15 VSS.t68 VSS.t63 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X468 OUT Transmission_Gate_Layout_13.CLKB.t13 Transmission_Gate_Layout_13.VIN.t41 VDD.t16 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X469 IN2 Transmission_Gate_Layout_18.CLKB.t15 Transmission_Gate_Layout_7.VIN.t33 VDD.t252 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X470 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t17 Transmission_Gate_Layout_6.VIN.t5 VDD.t88 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X471 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t49 Transmission_Gate_Layout_9.VIN.t39 VSS.t71 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X472 Transmission_Gate_Layout_16.CLKB EN.t92 VSS.t313 VSS.t225 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X473 IN5 EN.t93 Transmission_Gate_Layout_9.VIN.t54 VSS.t227 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X474 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT B1.t1 VSS.t106 VSS.t105 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X475 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t50 Transmission_Gate_Layout_9.VIN.t38 VSS.t89 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X476 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t15 Transmission_Gate_Layout_11.VIN.t27 VDD.t3 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X477 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t12 Transmission_Gate_Layout_1.VIN.t43 VDD.t66 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X478 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t16 Transmission_Gate_Layout_9.VOUT.t130 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X479 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t15 IN4.t9 VDD.t161 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X480 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t51 Transmission_Gate_Layout_4.VIN.t45 VSS.t71 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X481 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t13 OUT.t80 VSS.t181 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X482 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t26 Transmission_Gate_Layout_13.VIN.t101 VSS.t4 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X483 Transmission_Gate_Layout_7.VIN EN.t94 IN2.t39 VSS.t266 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X484 IN7 EN.t95 Transmission_Gate_Layout_4.VIN.t84 VSS.t261 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X485 Transmission_Gate_Layout_9.VIN EN.t96 IN5.t13 VSS.t223 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X486 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t18 IN3.t17 VDD.t40 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X487 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t52 Transmission_Gate_Layout_10.VIN.t63 VSS.t54 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X488 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t14 Transmission_Gate_Layout_2.VIN.t79 VDD.t76 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X489 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t18 Transmission_Gate_Layout_6.VIN.t6 VDD.t89 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X490 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t53 Transmission_Gate_Layout_4.VIN.t44 VSS.t52 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X491 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t50 Transmission_Gate_Layout_9.VOUT.t18 VSS.t133 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X492 VSS EN.t97 Transmission_Gate_Layout_21.CLKB.t5 VSS.t283 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X493 OUT Transmission_Gate_Layout_13.CLK.t16 Transmission_Gate_Layout_13.VIN.t50 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X494 IN2 Transmission_Gate_Layout_18.CLKB.t16 Transmission_Gate_Layout_7.VIN.t34 VDD.t178 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X495 IN8 Transmission_Gate_Layout_20.CLKB.t14 Transmission_Gate_Layout_5.VIN.t32 VDD.t134 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X496 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t15 Transmission_Gate_Layout_10.VIN.t31 VDD.t78 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X497 IN7 Transmission_Gate_Layout_17.CLKB.t14 Transmission_Gate_Layout_4.VIN.t4 VDD.t33 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X498 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t15 Transmission_Gate_Layout_9.VOUT.t58 VDD.t58 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X499 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t54 Transmission_Gate_Layout_1.VIN.t129 VSS.t53 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X500 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT Transmission_Gate_Layout_9.CLK.t55 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.t3 VDD.t298 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X501 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t56 Transmission_Gate_Layout_3.VIN.t132 VSS.t62 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X502 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t51 Transmission_Gate_Layout_2.VIN.t106 VSS.t127 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X503 IN6 Transmission_Gate_Layout_21.CLKB.t14 Transmission_Gate_Layout_8.VIN.t16 VDD.t43 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X504 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT A1.t2 VSS.t84 VSS.t83 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X505 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t19 Transmission_Gate_Layout_3.VIN.t20 VDD.t90 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X506 VDD Transmission_Gate_Layout_12.CLK.t14 Transmission_Gate_Layout_12.CLKB.t1 VDD.t214 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X507 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t52 Transmission_Gate_Layout_5.VIN.t52 VSS.t124 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X508 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t16 Transmission_Gate_Layout_9.VOUT.t59 VDD.t53 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X509 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t27 Transmission_Gate_Layout_9.VOUT.t37 VSS.t162 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X510 IN8 Transmission_Gate_Layout_20.CLKB.t15 Transmission_Gate_Layout_5.VIN.t61 VDD.t135 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X511 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t17 Transmission_Gate_Layout_9.VOUT.t129 VDD.t10 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X512 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t17 IN2.t12 VDD.t253 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X513 IN7 Transmission_Gate_Layout_17.CLKB.t15 Transmission_Gate_Layout_4.VIN.t5 VDD.t34 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X514 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLK.t53 VDD.t191 VDD.t180 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X515 Transmission_Gate_Layout_10.VIN EN.t98 IN3.t42 VSS.t220 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X516 Transmission_Gate_Layout_10.VIN EN.t99 IN3.t41 VSS.t236 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X517 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t54 Transmission_Gate_Layout_5.VIN.t51 VSS.t114 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X518 OUT Transmission_Gate_Layout_12.CLK.t15 Transmission_Gate_Layout_12.VIN.t97 VSS.t182 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X519 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t13 Transmission_Gate_Layout_12.VIN.t56 VDD.t63 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X520 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t57 Transmission_Gate_Layout_3.VIN.t133 VSS.t48 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X521 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t58 Transmission_Gate_Layout_9.VOUT.t95 VSS.t82 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X522 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t16 Transmission_Gate_Layout_10.VIN.t32 VDD.t73 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X523 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t13 IN1.t16 VDD.t227 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X524 VDD EN.t100 Transmission_Gate_Layout_21.CLKB.t1 VDD.t258 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X525 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t17 Transmission_Gate_Layout_9.VOUT.t60 VDD.t55 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X526 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t55 Transmission_Gate_Layout_9.VOUT.t17 VSS.t125 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X527 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t17 Transmission_Gate_Layout_2.VIN.t39 VDD.t74 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X528 VSS Transmission_Gate_Layout_12.CLK.t16 Transmission_Gate_Layout_12.CLKB.t4 VSS.t183 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X529 Transmission_Gate_Layout_6.VIN EN.t101 IN1.t39 VSS.t217 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X530 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_9.CLK.t59 VSS.t243 VSS.t78 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X531 VSS Transmission_Gate_Layout_11.CLK.t56 Transmission_Gate_Layout_8.CLKB.t4 VSS.t120 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X532 VDD Transmission_Gate_Layout_3.CLK.t28 Transmission_Gate_Layout_0.CLKB.t0 VDD.t185 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X533 OUT Transmission_Gate_Layout_13.CLKB.t14 Transmission_Gate_Layout_13.VIN.t69 VDD.t18 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X534 IN1 EN.t102 Transmission_Gate_Layout_6.VIN.t79 VSS.t214 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X535 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t25 Transmission_Gate_Layout_1.VIN.t1 VSS.t19 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X536 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t57 Transmission_Gate_Layout_8.VIN.t63 VSS.t114 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X537 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t60 Transmission_Gate_Layout_9.VIN.t36 VSS.t71 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X538 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t58 Transmission_Gate_Layout_11.VIN.t49 VSS.t130 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X539 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t14 Transmission_Gate_Layout_1.VIN.t47 VDD.t59 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X540 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t16 IN8.t14 VDD.t137 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X541 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t59 Transmission_Gate_Layout_9.VOUT.t16 VSS.t115 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X542 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t16 Transmission_Gate_Layout_11.VIN.t26 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X543 IN4 Transmission_Gate_Layout_19.CLKB.t16 Transmission_Gate_Layout_11.VIN.t10 VDD.t158 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X544 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t18 Transmission_Gate_Layout_13.VIN.t135 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X545 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t14 IN5.t39 VDD.t297 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X546 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 Transmission_Gate_Layout_9.CLK.t61 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.t2 VDD.t299 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X547 Transmission_Gate_Layout_4.VIN EN.t103 IN7.t30 VSS.t241 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X548 IN5 EN.t104 Transmission_Gate_Layout_9.VIN.t53 VSS.t215 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X549 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t16 Transmission_Gate_Layout_9.VOUT.t111 VDD.t62 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X550 OUT Transmission_Gate_Layout_12.CLKB.t18 Transmission_Gate_Layout_12.VIN.t43 VDD.t97 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X551 IN8 EN.t105 Transmission_Gate_Layout_5.VIN.t90 VSS.t221 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X552 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t17 OUT.t62 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X553 OUT Transmission_Gate_Layout_13.CLKB.t15 Transmission_Gate_Layout_13.VIN.t70 VDD.t47 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X554 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t17 Transmission_Gate_Layout_9.VOUT.t112 VDD.t61 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X555 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_11.CLK.t60 VDD.t190 VDD.t178 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X556 VDD Transmission_Gate_Layout_1.CLK.t26 Transmission_Gate_Layout_2.CLKB.t0 VDD.t19 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X557 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t18 IN2.t11 VDD.t248 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X558 VSS Transmission_Gate_Layout_11.CLK.t61 Transmission_Gate_Layout_5.CLKB.t4 VSS.t120 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X559 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t18 Transmission_Gate_Layout_2.VIN.t40 VDD.t71 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X560 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.t4 VDD.t167 VDD.t166 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X561 IN6 Transmission_Gate_Layout_21.CLKB.t15 Transmission_Gate_Layout_8.VIN.t17 VDD.t44 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X562 Transmission_Gate_Layout_4.VIN EN.t106 IN7.t29 VSS.t237 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X563 VDD Transmission_Gate_Layout_11.CLK.t62 Transmission_Gate_Layout_5.CLKB.t1 VDD.t182 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X564 IN8 EN.t107 Transmission_Gate_Layout_5.VIN.t89 VSS.t279 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X565 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t27 Transmission_Gate_Layout_13.VIN.t15 VSS.t20 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X566 IN8 Transmission_Gate_Layout_20.CLKB.t17 Transmission_Gate_Layout_5.VIN.t63 VDD.t131 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X567 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t18 Transmission_Gate_Layout_9.VOUT.t128 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X568 IN6 Transmission_Gate_Layout_21.CLKB.t16 Transmission_Gate_Layout_8.VIN.t18 VDD.t45 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X569 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.t2 VSS.t98 VSS.t97 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X570 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t63 Transmission_Gate_Layout_3.VIN.t48 VSS.t128 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X571 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t62 Transmission_Gate_Layout_9.VOUT.t94 VSS.t53 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X572 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t29 Transmission_Gate_Layout_13.VIN.t102 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X573 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t19 IN3.t16 VDD.t40 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X574 OUT Transmission_Gate_Layout_12.CLK.t17 Transmission_Gate_Layout_12.VIN.t98 VSS.t187 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X575 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t15 Transmission_Gate_Layout_12.VIN.t58 VDD.t60 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X576 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t16 IN7.t6 VDD.t35 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X577 VSS EN.t108 Transmission_Gate_Layout_18.CLKB.t4 VSS.t233 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X578 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t18 IN8.t16 VDD.t132 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X579 IN3 Transmission_Gate_Layout_14.CLKB.t20 Transmission_Gate_Layout_10.VIN.t9 VDD.t42 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X580 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_9.CLK.t63 VSS.t244 VSS.t78 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X581 VSS Transmission_Gate_Layout_1.CLK.t28 Transmission_Gate_Layout_2.CLKB.t1 VSS.t21 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X582 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_9.CLK.t64 VDD.t300 VDD.t122 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X583 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t64 Transmission_Gate_Layout_2.VIN.t105 VSS.t128 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X584 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t65 Transmission_Gate_Layout_8.VIN.t61 VSS.t124 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X585 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t19 OUT.t43 VDD.t98 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X586 VDD Transmission_Gate_Layout_9.CLK.t65 Transmission_Gate_Layout_6.CLKB.t1 VDD.t227 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X587 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t66 Transmission_Gate_Layout_2.VIN.t138 VSS.t62 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X588 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t67 Transmission_Gate_Layout_9.VIN.t34 VSS.t81 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X589 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t17 IN4.t11 VDD.t155 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X590 OUT Transmission_Gate_Layout_13.CLK.t18 Transmission_Gate_Layout_13.VIN.t52 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X591 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t17 IN7.t7 VDD.t36 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X592 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t68 Transmission_Gate_Layout_10.VIN.t61 VSS.t90 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X593 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t18 Transmission_Gate_Layout_9.VIN.t11 VDD.t64 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X594 VDD Transmission_Gate_Layout_12.CLK.t18 Transmission_Gate_Layout_12.CLKB.t0 VDD.t214 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X595 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t15 Transmission_Gate_Layout_13.VIN.t89 VDD.t77 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X596 Transmission_Gate_Layout_9.VIN EN.t109 IN5.t11 VSS.t299 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X597 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t18 IN7.t8 VDD.t31 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X598 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t19 IN8.t17 VDD.t133 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X599 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t29 Transmission_Gate_Layout_1.VIN.t2 VSS.t24 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X600 IN1 Transmission_Gate_Layout_16.CLKB.t14 Transmission_Gate_Layout_6.VIN.t68 VDD.t242 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X601 IN5 EN.t110 Transmission_Gate_Layout_9.VIN.t52 VSS.t231 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X602 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t17 IN6.t19 VDD.t0 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X603 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t69 Transmission_Gate_Layout_9.VIN.t33 VSS.t89 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X604 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t30 Transmission_Gate_Layout_9.VOUT.t38 VSS.t163 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X605 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t66 Transmission_Gate_Layout_8.VIN.t60 VSS.t124 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X606 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t30 Transmission_Gate_Layout_2.VIN.t7 VSS.t25 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X607 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t19 Transmission_Gate_Layout_9.VOUT.t127 VDD.t52 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X608 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t19 Transmission_Gate_Layout_13.VIN.t136 VDD.t162 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X609 IN2 Transmission_Gate_Layout_18.CLKB.t19 Transmission_Gate_Layout_7.VIN.t37 VDD.t249 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X610 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t18 IN6.t20 VDD.t46 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X611 Transmission_Gate_Layout_9.VIN EN.t111 IN5.t9 VSS.t296 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X612 VDD EN.t112 Transmission_Gate_Layout_18.CLKB.t2 VDD.t99 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X613 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1 C1.t1 VDD.t204 VDD.t203 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X614 IN3 EN.t113 Transmission_Gate_Layout_10.VIN.t84 VSS.t280 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X615 VSS Transmission_Gate_Layout_11.CLK.t67 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.t3 VSS.t49 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X616 IN5 Transmission_Gate_Layout_15.CLKB.t15 Transmission_Gate_Layout_9.VIN.t82 VDD.t296 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X617 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t19 OUT.t83 VSS.t188 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X618 Transmission_Gate_Layout_19.CLKB EN.t114 VSS.t307 VSS.t292 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X619 OUT Transmission_Gate_Layout_13.CLKB.t16 Transmission_Gate_Layout_13.VIN.t60 VDD.t12 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X620 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t68 Transmission_Gate_Layout_11.VIN.t47 VSS.t126 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X621 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLK.t70 VDD.t303 VDD.t24 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X622 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t31 Transmission_Gate_Layout_13.VIN.t17 VSS.t26 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X623 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t17 Transmission_Gate_Layout_11.VIN.t25 VDD.t5 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X624 IN2 EN.t115 Transmission_Gate_Layout_7.VIN.t87 VSS.t271 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X625 IN5 Transmission_Gate_Layout_15.CLKB.t16 Transmission_Gate_Layout_9.VIN.t81 VDD.t292 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X626 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t19 IN6.t21 VDD.t41 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X627 Transmission_Gate_Layout_17.CLKB EN.t116 VSS.t308 VSS.t294 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X628 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t31 Transmission_Gate_Layout_13.VIN.t103 VSS.t164 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X629 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t32 Transmission_Gate_Layout_13.VIN.t104 VSS.t165 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X630 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t71 Transmission_Gate_Layout_2.VIN.t137 VSS.t55 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X631 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t72 Transmission_Gate_Layout_10.VIN.t59 VSS.t47 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X632 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t16 Transmission_Gate_Layout_2.VIN.t78 VDD.t72 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X633 OUT Transmission_Gate_Layout_12.CLKB.t20 Transmission_Gate_Layout_12.VIN.t45 VDD.t97 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X634 IN7 Transmission_Gate_Layout_17.CLKB.t19 Transmission_Gate_Layout_4.VIN.t9 VDD.t33 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X635 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t20 Transmission_Gate_Layout_3.VIN.t102 VDD.t3 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X636 OUT Transmission_Gate_Layout_13.CLK.t19 Transmission_Gate_Layout_13.VIN.t53 VSS.t9 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X637 Transmission_Gate_Layout_9.VIN EN.t117 IN5.t8 VSS.t224 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X638 Transmission_Gate_Layout_5.VIN EN.t118 IN8.t35 VSS.t289 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X639 VDD Transmission_Gate_Layout_1.CLK.t32 Transmission_Gate_Layout_2.CLKB.t2 VDD.t19 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X640 IN1 EN.t119 Transmission_Gate_Layout_6.VIN.t78 VSS.t288 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X641 VSS Transmission_Gate_Layout_11.CLK.t69 Transmission_Gate_Layout_8.CLKB.t3 VSS.t120 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X642 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t18 Transmission_Gate_Layout_9.VOUT.t61 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X643 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t19 Transmission_Gate_Layout_9.VIN.t10 VDD.t65 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X644 VSS Transmission_Gate_Layout_3.CLK.t33 Transmission_Gate_Layout_0.CLKB.t1 VSS.t166 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X645 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t20 IN8.t18 VDD.t136 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X646 OUT Transmission_Gate_Layout_13.CLK.t20 Transmission_Gate_Layout_13.VIN.t54 VSS.t8 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X647 Transmission_Gate_Layout_6.VIN EN.t120 IN1.t36 VSS.t222 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X648 Transmission_Gate_Layout_9.CLK Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.t2 VDD.t127 VDD.t126 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X649 IN6 EN.t121 Transmission_Gate_Layout_8.VIN.t89 VSS.t279 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X650 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t17 OUT.t12 VDD.t13 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X651 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t15 Transmission_Gate_Layout_3.VIN.t118 VDD.t105 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X652 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.t3 VDD.t175 VDD.t139 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X653 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t33 Transmission_Gate_Layout_1.VIN.t3 VSS.t27 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X654 Transmission_Gate_Layout_6.VIN EN.t122 IN1.t35 VSS.t262 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X655 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t17 IN5.t36 VDD.t295 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X656 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t14 Transmission_Gate_Layout_4.VIN.t64 VDD.t31 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X657 IN1 EN.t123 Transmission_Gate_Layout_6.VIN.t77 VSS.t286 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X658 Transmission_Gate_Layout_6.VIN EN.t124 IN1.t33 VSS.t219 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X659 Transmission_Gate_Layout_11.VIN EN.t125 IN4.t38 VSS.t282 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X660 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT A1.t3 VSS.t86 VSS.t85 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X661 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLK.t73 VSS.t245 VSS.t78 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X662 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t34 Transmission_Gate_Layout_3.VIN.t74 VSS.t169 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X663 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t20 Transmission_Gate_Layout_12.VIN.t134 VDD.t53 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X664 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t18 IN5.t35 VDD.t182 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X665 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t19 IN5.t34 VDD.t291 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X666 OUT Transmission_Gate_Layout_12.CLK.t20 Transmission_Gate_Layout_12.VIN.t100 VSS.t186 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X667 IN3 Transmission_Gate_Layout_14.CLKB.t21 Transmission_Gate_Layout_10.VIN.t8 VDD.t42 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X668 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t35 Transmission_Gate_Layout_3.VIN.t75 VSS.t170 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X669 IN4 EN.t126 Transmission_Gate_Layout_11.VIN.t80 VSS.t260 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X670 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t21 OUT.t45 VDD.t98 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X671 Transmission_Gate_Layout_19.CLKB EN.t127 VDD.t272 VDD.t131 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X672 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t15 IN1.t14 VDD.t244 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X673 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t21 OUT.t58 VSS.t10 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X674 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t15 Transmission_Gate_Layout_5.VIN.t9 VDD.t120 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X675 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t17 Transmission_Gate_Layout_13.VIN.t87 VDD.t77 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X676 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t19 Transmission_Gate_Layout_8.VIN.t34 VDD.t10 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X677 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t16 Transmission_Gate_Layout_7.VIN.t71 VDD.t103 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X678 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLK.t70 VSS.t134 VSS.t118 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X679 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t18 Transmission_Gate_Layout_2.VIN.t3 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X680 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLK.t36 VDD.t211 VDD.t180 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X681 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t20 IN5.t33 VDD.t297 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X682 VSS Transmission_Gate_Layout_1.CLK.t34 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.t3 VSS.t28 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X683 Transmission_Gate_Layout_7.VIN EN.t128 IN2.t37 VSS.t255 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X684 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t16 IN1.t13 VDD.t245 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X685 IN8 EN.t129 Transmission_Gate_Layout_5.VIN.t88 VSS.t230 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X686 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t35 Transmission_Gate_Layout_12.VIN.t5 VSS.t31 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X687 Transmission_Gate_Layout_17.CLKB EN.t130 VDD.t271 VDD.t122 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X688 IN8 Transmission_Gate_Layout_20.CLKB.t21 Transmission_Gate_Layout_5.VIN.t67 VDD.t138 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X689 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t36 Transmission_Gate_Layout_2.VIN.t9 VSS.t32 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X690 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t21 Transmission_Gate_Layout_13.VIN.t138 VDD.t162 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X691 IN1 EN.t131 Transmission_Gate_Layout_6.VIN.t76 VSS.t216 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X692 Transmission_Gate_Layout_12.CLK Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.t2 VDD.t231 VDD.t230 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X693 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t37 Transmission_Gate_Layout_12.VIN.t78 VSS.t171 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X694 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t38 Transmission_Gate_Layout_12.VIN.t79 VSS.t172 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X695 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t74 Transmission_Gate_Layout_10.VIN.t58 VSS.t43 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X696 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t20 Transmission_Gate_Layout_9.VOUT.t115 VDD.t63 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X697 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t18 Transmission_Gate_Layout_2.VIN.t77 VDD.t73 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X698 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t71 Transmission_Gate_Layout_9.VOUT.t15 VSS.t122 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X699 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t21 Transmission_Gate_Layout_12.VIN.t133 VDD.t55 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X700 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t15 Transmission_Gate_Layout_1.VIN.t121 VDD.t33 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X701 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t72 Transmission_Gate_Layout_1.VIN.t101 VSS.t115 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X702 IN3 EN.t132 Transmission_Gate_Layout_10.VIN.t83 VSS.t276 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X703 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t22 Transmission_Gate_Layout_3.VIN.t104 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X704 OUT Transmission_Gate_Layout_13.CLKB.t18 Transmission_Gate_Layout_13.VIN.t64 VDD.t12 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X705 IN1 Transmission_Gate_Layout_16.CLKB.t17 Transmission_Gate_Layout_6.VIN.t71 VDD.t243 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X706 IN4 EN.t133 Transmission_Gate_Layout_11.VIN.t79 VSS.t281 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X707 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t73 Transmission_Gate_Layout_1.VIN.t100 VSS.t133 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X708 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t19 OUT.t10 VDD.t56 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X709 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t75 Transmission_Gate_Layout_4.VIN.t42 VSS.t89 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X710 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t20 Transmission_Gate_Layout_8.VIN.t33 VDD.t57 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X711 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t19 Transmission_Gate_Layout_2.VIN.t41 VDD.t75 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X712 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t16 Transmission_Gate_Layout_12.VIN.t59 VDD.t61 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X713 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t76 Transmission_Gate_Layout_6.VIN.t32 VSS.t43 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X714 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t19 Transmission_Gate_Layout_2.VIN.t4 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X715 Transmission_Gate_Layout_11.VIN EN.t134 IN4.t35 VSS.t242 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X716 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t16 Transmission_Gate_Layout_1.VIN.t71 VDD.t119 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X717 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t74 Transmission_Gate_Layout_5.VIN.t50 VSS.t117 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X718 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t39 Transmission_Gate_Layout_9.VOUT.t41 VSS.t173 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X719 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t20 OUT.t9 VDD.t54 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X720 IN1 Transmission_Gate_Layout_16.CLKB.t18 Transmission_Gate_Layout_6.VIN.t48 VDD.t240 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X721 IN1 Transmission_Gate_Layout_16.CLKB.t19 Transmission_Gate_Layout_6.VIN.t49 VDD.t241 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X722 IN4 EN.t135 Transmission_Gate_Layout_11.VIN.t78 VSS.t277 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X723 Transmission_Gate_Layout_4.VIN EN.t136 IN7.t28 VSS.t252 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X724 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t77 Transmission_Gate_Layout_9.VOUT.t93 VSS.t56 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X725 VSS EN.t137 Transmission_Gate_Layout_14.CLKB.t4 VSS.t268 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X726 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t17 Transmission_Gate_Layout_12.VIN.t60 VDD.t62 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X727 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t18 IN4.t12 VDD.t157 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X728 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t17 Transmission_Gate_Layout_1.VIN.t72 VDD.t113 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X729 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t78 Transmission_Gate_Layout_4.VIN.t41 VSS.t71 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X730 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t79 Transmission_Gate_Layout_3.VIN.t135 VSS.t55 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X731 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t16 Transmission_Gate_Layout_4.VIN.t66 VDD.t32 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X732 OUT Transmission_Gate_Layout_12.CLK.t21 Transmission_Gate_Layout_12.VIN.t101 VSS.t189 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X733 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t37 Transmission_Gate_Layout_13.VIN.t19 VSS.t33 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X734 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t40 Transmission_Gate_Layout_3.VIN.t76 VSS.t157 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X735 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t23 Transmission_Gate_Layout_3.VIN.t105 VDD.t3 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X736 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t17 Transmission_Gate_Layout_3.VIN.t129 VDD.t101 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X737 Transmission_Gate_Layout_8.VIN EN.t138 IN6.t36 VSS.t289 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X738 IN3 Transmission_Gate_Layout_14.CLKB.t22 Transmission_Gate_Layout_10.VIN.t7 VDD.t45 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X739 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t80 Transmission_Gate_Layout_2.VIN.t136 VSS.t62 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X740 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t19 Transmission_Gate_Layout_13.VIN.t85 VDD.t71 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X741 IN2 EN.t139 Transmission_Gate_Layout_7.VIN.t84 VSS.t232 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X742 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t81 Transmission_Gate_Layout_3.VIN.t136 VSS.t62 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X743 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t22 OUT.t46 VDD.t93 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X744 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t18 Transmission_Gate_Layout_7.VIN.t63 VDD.t100 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X745 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t22 OUT.t57 VSS.t12 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X746 Transmission_Gate_Layout_7.VIN EN.t140 IN2.t35 VSS.t278 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X747 IN1 Transmission_Gate_Layout_16.CLKB.t20 Transmission_Gate_Layout_6.VIN.t50 VDD.t242 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X748 VSS EN.t141 Transmission_Gate_Layout_20.CLKB.t4 VSS.t283 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X749 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t21 OUT.t8 VDD.t13 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X750 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t17 Transmission_Gate_Layout_1.VIN.t123 VDD.t29 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X751 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t21 Transmission_Gate_Layout_8.VIN.t32 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X752 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t21 Transmission_Gate_Layout_9.VIN.t8 VDD.t66 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X753 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t38 Transmission_Gate_Layout_12.VIN.t6 VSS.t34 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X754 VDD EN.t142 Transmission_Gate_Layout_20.CLKB.t1 VDD.t161 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X755 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT B1.t2 VSS.t107 VSS.t28 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X756 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_11.CLK.t75 VSS.t132 VSS.t118 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X757 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t82 Transmission_Gate_Layout_6.VIN.t29 VSS.t54 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X758 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t20 IN6.t22 VDD.t40 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X759 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t20 Transmission_Gate_Layout_2.VIN.t5 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X760 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t76 Transmission_Gate_Layout_3.VIN.t47 VSS.t131 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X761 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t20 Transmission_Gate_Layout_10.VIN.t36 VDD.t76 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X762 VDD B1.t3 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.t1 VDD.t107 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X763 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t18 Transmission_Gate_Layout_1.VIN.t51 VDD.t64 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X764 IN5 Transmission_Gate_Layout_15.CLKB.t21 Transmission_Gate_Layout_9.VIN.t80 VDD.t296 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X765 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t18 Transmission_Gate_Layout_1.VIN.t124 VDD.t30 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X766 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t39 Transmission_Gate_Layout_2.VIN.t11 VSS.t35 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X767 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t22 Transmission_Gate_Layout_12.VIN.t132 VDD.t53 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X768 IN3 EN.t143 Transmission_Gate_Layout_10.VIN.t82 VSS.t256 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X769 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t77 Transmission_Gate_Layout_7.VIN.t10 VSS.t116 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X770 IN3 EN.t144 Transmission_Gate_Layout_10.VIN.t81 VSS.t258 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X771 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLK.t23 VDD.t51 VDD.t14 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X772 Transmission_Gate_Layout_11.CLK Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.t2 VSS.t88 VSS.t87 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X773 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t22 OUT.t86 VSS.t191 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X774 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t18 Transmission_Gate_Layout_5.VIN.t12 VDD.t114 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X775 Transmission_Gate_Layout_5.VIN EN.t145 IN8.t33 VSS.t238 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X776 Transmission_Gate_Layout_8.VIN EN.t146 IN6.t35 VSS.t275 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X777 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t23 OUT.t87 VSS.t190 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X778 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t78 Transmission_Gate_Layout_7.VIN.t9 VSS.t130 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X779 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t23 OUT.t24 VDD.t91 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X780 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t23 IN3.t15 VDD.t46 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X781 IN7 EN.t147 Transmission_Gate_Layout_4.VIN.t80 VSS.t228 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X782 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t19 Transmission_Gate_Layout_3.VIN.t112 VDD.t106 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X783 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t83 Transmission_Gate_Layout_1.VIN.t132 VSS.t82 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X784 IN4 Transmission_Gate_Layout_19.CLKB.t19 Transmission_Gate_Layout_11.VIN.t61 VDD.t159 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X785 Transmission_Gate_Layout_4.VIN EN.t148 IN7.t27 VSS.t274 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X786 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t19 Transmission_Gate_Layout_1.VIN.t125 VDD.t34 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X787 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t79 Transmission_Gate_Layout_1.VIN.t98 VSS.t125 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X788 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t84 Transmission_Gate_Layout_1.VIN.t133 VSS.t82 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X789 IN8 EN.t149 Transmission_Gate_Layout_5.VIN.t87 VSS.t230 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X790 IN6 EN.t150 Transmission_Gate_Layout_8.VIN.t88 VSS.t230 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X791 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLK.t40 VDD.t25 VDD.t24 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X792 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t19 Transmission_Gate_Layout_1.VIN.t74 VDD.t115 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X793 Transmission_Gate_Layout_8.VIN EN.t151 IN6.t33 VSS.t238 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X794 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t41 Transmission_Gate_Layout_1.VIN.t6 VSS.t36 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X795 IN2 EN.t152 Transmission_Gate_Layout_7.VIN.t83 VSS.t272 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X796 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t80 Transmission_Gate_Layout_1.VIN.t97 VSS.t122 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X797 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t21 Transmission_Gate_Layout_11.VIN.t21 VDD.t144 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X798 IN4 Transmission_Gate_Layout_19.CLKB.t20 Transmission_Gate_Layout_11.VIN.t62 VDD.t160 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X799 Transmission_Gate_Layout_7.VIN EN.t153 IN2.t33 VSS.t273 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X800 Transmission_Gate_Layout_11.VIN EN.t154 IN4.t33 VSS.t267 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X801 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t81 Transmission_Gate_Layout_7.VIN.t8 VSS.t130 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X802 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t82 Transmission_Gate_Layout_1.VIN.t96 VSS.t115 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X803 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t20 Transmission_Gate_Layout_7.VIN.t61 VDD.t104 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X804 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t20 Transmission_Gate_Layout_6.VIN.t8 VDD.t83 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X805 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t83 Transmission_Gate_Layout_1.VIN.t95 VSS.t125 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X806 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t24 Transmission_Gate_Layout_3.VIN.t106 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X807 IN4 EN.t155 Transmission_Gate_Layout_11.VIN.t77 VSS.t264 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X808 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t20 Transmission_Gate_Layout_1.VIN.t75 VDD.t116 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X809 VDD Transmission_Gate_Layout_11.CLK.t84 Transmission_Gate_Layout_8.CLKB.t0 VDD.t185 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X810 Transmission_Gate_Layout_10.VIN EN.t156 IN3.t40 VSS.t251 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X811 Transmission_Gate_Layout_10.VIN EN.t157 IN3.t39 VSS.t257 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X812 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t22 IN5.t31 VDD.t295 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X813 Transmission_Gate_Layout_8.VIN EN.t158 IN6.t32 VSS.t265 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X814 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t22 Transmission_Gate_Layout_9.VIN.t7 VDD.t59 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X815 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t24 IN3.t14 VDD.t41 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X816 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t22 OUT.t7 VDD.t56 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X817 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t20 IN2.t9 VDD.t251 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X818 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLK.t41 VSS.t174 VSS.t158 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X819 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLK.t42 VSS.t37 VSS.t17 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X820 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t21 Transmission_Gate_Layout_5.VIN.t15 VDD.t117 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X821 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t21 Transmission_Gate_Layout_10.VIN.t37 VDD.t78 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X822 OUT Transmission_Gate_Layout_12.CLKB.t24 Transmission_Gate_Layout_12.VIN.t26 VDD.t92 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X823 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t19 Transmission_Gate_Layout_12.VIN.t62 VDD.t61 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X824 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t22 Transmission_Gate_Layout_9.VOUT.t65 VDD.t58 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X825 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t23 IN5.t30 VDD.t182 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X826 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t85 Transmission_Gate_Layout_9.VIN.t31 VSS.t71 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X827 IN6 Transmission_Gate_Layout_21.CLKB.t21 Transmission_Gate_Layout_8.VIN.t23 VDD.t43 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X828 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t43 Transmission_Gate_Layout_2.VIN.t12 VSS.t38 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X829 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t21 IN2.t8 VDD.t250 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X830 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t21 Transmission_Gate_Layout_3.VIN.t22 VDD.t90 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X831 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t42 Transmission_Gate_Layout_12.VIN.t81 VSS.t160 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X832 Transmission_Gate_Layout_7.VIN EN.t159 IN2.t32 VSS.t266 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X833 IN7 EN.t160 Transmission_Gate_Layout_4.VIN.t78 VSS.t261 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X834 Transmission_Gate_Layout_9.VIN EN.t161 IN5.t7 VSS.t223 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X835 Transmission_Gate_Layout_19.CLKB EN.t162 VDD.t268 VDD.t131 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X836 VDD Transmission_Gate_Layout_9.CLK.t86 Transmission_Gate_Layout_10.CLKB.t1 VDD.t19 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X837 IN3 Transmission_Gate_Layout_14.CLKB.t25 Transmission_Gate_Layout_10.VIN.t4 VDD.t45 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X838 IN4 Transmission_Gate_Layout_19.CLKB.t21 Transmission_Gate_Layout_11.VIN.t63 VDD.t156 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X839 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t87 Transmission_Gate_Layout_9.VIN.t30 VSS.t52 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X840 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t43 Transmission_Gate_Layout_3.VIN.t77 VSS.t156 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X841 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t20 Transmission_Gate_Layout_1.VIN.t53 VDD.t65 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X842 IN2 EN.t163 Transmission_Gate_Layout_7.VIN.t80 VSS.t263 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X843 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t25 OUT.t26 VDD.t93 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X844 VSS EN.t164 Transmission_Gate_Layout_21.CLKB.t4 VSS.t283 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X845 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT A1.t4 VDD.t177 VDD.t176 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X846 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t85 Transmission_Gate_Layout_3.VIN.t46 VSS.t128 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X847 Transmission_Gate_Layout_17.CLKB EN.t165 VDD.t267 VDD.t122 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X848 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t22 Transmission_Gate_Layout_3.VIN.t23 VDD.t85 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X849 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t86 Transmission_Gate_Layout_5.VIN.t49 VSS.t124 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X850 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t20 IN7.t10 VDD.t32 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X851 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t21 Transmission_Gate_Layout_3.VIN.t119 VDD.t102 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X852 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t22 Transmission_Gate_Layout_5.VIN.t16 VDD.t118 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X853 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t88 Transmission_Gate_Layout_4.VIN.t38 VSS.t81 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X854 VDD EN.t166 Transmission_Gate_Layout_21.CLKB.t0 VDD.t258 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X855 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t23 Transmission_Gate_Layout_9.VOUT.t2 VDD.t60 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X856 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t24 OUT.t56 VSS.t11 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X857 Transmission_Gate_Layout_11.VIN EN.t167 IN4.t31 VSS.t259 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X858 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t20 Transmission_Gate_Layout_4.VIN.t70 VDD.t35 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X859 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t89 Transmission_Gate_Layout_6.VIN.t28 VSS.t90 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X860 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t22 Transmission_Gate_Layout_2.VIN.t44 VDD.t74 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X861 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t44 Transmission_Gate_Layout_12.VIN.t8 VSS.t39 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X862 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t21 Transmission_Gate_Layout_1.VIN.t54 VDD.t64 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X863 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t23 Transmission_Gate_Layout_6.VIN.t11 VDD.t84 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X864 IN6 Transmission_Gate_Layout_21.CLKB.t22 Transmission_Gate_Layout_8.VIN.t0 VDD.t42 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X865 IN2 Transmission_Gate_Layout_18.CLKB.t22 Transmission_Gate_Layout_7.VIN.t40 VDD.t252 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X866 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t44 Transmission_Gate_Layout_12.VIN.t82 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X867 Transmission_Gate_Layout_5.VIN EN.t168 IN8.t31 VSS.t265 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X868 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t22 IN4.t16 VDD.t161 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X869 IN2 Transmission_Gate_Layout_18.CLKB.t23 Transmission_Gate_Layout_7.VIN.t41 VDD.t171 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X870 IN1 Transmission_Gate_Layout_16.CLKB.t21 Transmission_Gate_Layout_6.VIN.t51 VDD.t243 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X871 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t90 Transmission_Gate_Layout_4.VIN.t37 VSS.t89 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X872 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t45 Transmission_Gate_Layout_13.VIN.t22 VSS.t40 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X873 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t21 Transmission_Gate_Layout_4.VIN.t16 VDD.t36 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X874 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t24 Transmission_Gate_Layout_3.VIN.t25 VDD.t86 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X875 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t23 Transmission_Gate_Layout_2.VIN.t45 VDD.t77 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X876 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t26 IN3.t13 VDD.t46 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X877 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t91 Transmission_Gate_Layout_9.VOUT.t92 VSS.t82 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X878 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t87 Transmission_Gate_Layout_2.VIN.t104 VSS.t128 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X879 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t25 Transmission_Gate_Layout_13.VIN.t142 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X880 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t88 Transmission_Gate_Layout_9.VOUT.t14 VSS.t125 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X881 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t23 OUT.t6 VDD.t17 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X882 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t23 IN4.t17 VDD.t154 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X883 IN1 Transmission_Gate_Layout_16.CLKB.t22 Transmission_Gate_Layout_6.VIN.t52 VDD.t240 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X884 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLK.t46 VDD.t26 VDD.t24 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X885 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t89 Transmission_Gate_Layout_7.VIN.t6 VSS.t126 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X886 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t90 Transmission_Gate_Layout_8.VIN.t57 VSS.t113 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X887 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t22 Transmission_Gate_Layout_2.VIN.t113 VDD.t162 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X888 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t23 Transmission_Gate_Layout_8.VIN.t30 VDD.t52 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X889 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t24 IN4.t18 VDD.t157 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X890 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t22 Transmission_Gate_Layout_7.VIN.t55 VDD.t99 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X891 IN1 EN.t169 Transmission_Gate_Layout_6.VIN.t75 VSS.t214 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X892 IN6 Transmission_Gate_Layout_21.CLKB.t23 Transmission_Gate_Layout_8.VIN.t1 VDD.t44 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X893 Transmission_Gate_Layout_15.CLKB EN.t170 VSS.t300 VSS.t253 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X894 VDD Transmission_Gate_Layout_11.CLK.t91 Transmission_Gate_Layout_5.CLKB.t0 VDD.t182 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X895 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t92 Transmission_Gate_Layout_11.VIN.t45 VSS.t130 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X896 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t93 Transmission_Gate_Layout_9.VOUT.t13 VSS.t115 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X897 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t20 Transmission_Gate_Layout_13.VIN.t84 VDD.t75 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X898 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t94 Transmission_Gate_Layout_3.VIN.t45 VSS.t127 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X899 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLK.t25 VSS.t69 VSS.t63 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X900 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t24 IN2.t5 VDD.t253 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X901 IN7 Transmission_Gate_Layout_17.CLKB.t21 Transmission_Gate_Layout_4.VIN.t11 VDD.t34 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X902 IN8 Transmission_Gate_Layout_20.CLKB.t22 Transmission_Gate_Layout_5.VIN.t68 VDD.t131 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X903 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t45 Transmission_Gate_Layout_9.VOUT.t44 VSS.t161 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X904 Transmission_Gate_Layout_4.VIN EN.t171 IN7.t26 VSS.t241 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X905 IN5 EN.t172 Transmission_Gate_Layout_9.VIN.t51 VSS.t215 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X906 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t92 Transmission_Gate_Layout_3.VIN.t139 VSS.t55 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X907 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t24 OUT.t88 VSS.t181 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X908 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK.t95 Transmission_Gate_Layout_3.VIN.t44 VSS.t112 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X909 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t96 Transmission_Gate_Layout_8.VIN.t55 VSS.t114 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X910 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t26 OUT.t55 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X911 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t23 Transmission_Gate_Layout_9.VOUT.t123 VDD.t57 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X912 IN7 EN.t173 Transmission_Gate_Layout_4.VIN.t76 VSS.t240 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X913 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t25 Transmission_Gate_Layout_3.VIN.t26 VDD.t87 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X914 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t47 Transmission_Gate_Layout_12.VIN.t9 VSS.t16 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X915 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_9.CLK.t93 VDD.t306 VDD.t122 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X916 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t97 Transmission_Gate_Layout_7.VIN.t3 VSS.t126 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X917 Transmission_Gate_Layout_4.VIN EN.t174 IN7.t25 VSS.t237 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X918 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t94 Transmission_Gate_Layout_1.VIN.t136 VSS.t56 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X919 OUT Transmission_Gate_Layout_13.CLKB.t24 Transmission_Gate_Layout_13.VIN.t12 VDD.t16 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X920 Transmission_Gate_Layout_15.CLKB EN.t175 VDD.t264 VDD.t113 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X921 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t26 Transmission_Gate_Layout_6.VIN.t14 VDD.t88 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X922 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t24 Transmission_Gate_Layout_10.VIN.t40 VDD.t72 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X923 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t48 Transmission_Gate_Layout_13.VIN.t23 VSS.t20 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X924 IN7 EN.t176 Transmission_Gate_Layout_4.VIN.t74 VSS.t239 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X925 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t23 Transmission_Gate_Layout_11.VIN.t19 VDD.t3 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X926 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t22 Transmission_Gate_Layout_1.VIN.t55 VDD.t66 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X927 Transmission_Gate_Layout_1.CLK Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.t3 VDD.t146 VDD.t145 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X928 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT C1.t2 VSS.t151 VSS.t150 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X929 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t24 IN6.t2 VDD.t0 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X930 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t98 Transmission_Gate_Layout_9.VOUT.t12 VSS.t122 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X931 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t21 Transmission_Gate_Layout_2.VIN.t76 VDD.t76 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X932 VSS EN.t177 Transmission_Gate_Layout_18.CLKB.t3 VSS.t233 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X933 IN4 Transmission_Gate_Layout_19.CLKB.t25 Transmission_Gate_Layout_11.VIN.t67 VDD.t159 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X934 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t27 Transmission_Gate_Layout_6.VIN.t15 VDD.t89 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X935 IN7 Transmission_Gate_Layout_17.CLKB.t22 Transmission_Gate_Layout_4.VIN.t12 VDD.t29 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X936 VSS Transmission_Gate_Layout_11.CLK.t99 Transmission_Gate_Layout_5.CLKB.t3 VSS.t120 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X937 Transmission_Gate_Layout_10.VIN EN.t178 IN3.t38 VSS.t236 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X938 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t46 Transmission_Gate_Layout_13.VIN.t109 VSS.t4 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X939 IN8 Transmission_Gate_Layout_20.CLKB.t23 Transmission_Gate_Layout_5.VIN.t69 VDD.t134 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X940 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t100 Transmission_Gate_Layout_2.VIN.t103 VSS.t128 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X941 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t101 Transmission_Gate_Layout_8.VIN.t53 VSS.t124 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X942 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t95 Transmission_Gate_Layout_6.VIN.t26 VSS.t90 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X943 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t102 Transmission_Gate_Layout_2.VIN.t102 VSS.t127 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X944 OUT Transmission_Gate_Layout_12.CLK.t25 Transmission_Gate_Layout_12.VIN.t105 VSS.t182 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X945 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t26 Transmission_Gate_Layout_13.VIN.t71 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X946 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t96 Transmission_Gate_Layout_9.VIN.t28 VSS.t81 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X947 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t103 Transmission_Gate_Layout_11.VIN.t42 VSS.t116 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X948 OUT Transmission_Gate_Layout_13.CLK.t27 Transmission_Gate_Layout_13.VIN.t5 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X949 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t97 Transmission_Gate_Layout_10.VIN.t56 VSS.t90 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X950 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t98 Transmission_Gate_Layout_9.VOUT.t91 VSS.t53 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X951 OUT Transmission_Gate_Layout_13.CLK.t28 Transmission_Gate_Layout_13.VIN.t6 VSS.t7 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X952 IN4 Transmission_Gate_Layout_19.CLKB.t26 Transmission_Gate_Layout_11.VIN.t68 VDD.t160 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X953 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t49 Transmission_Gate_Layout_1.VIN.t9 VSS.t24 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X954 Transmission_Gate_Layout_9.VIN EN.t179 IN5.t5 VSS.t299 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X955 IN7 Transmission_Gate_Layout_17.CLKB.t23 Transmission_Gate_Layout_4.VIN.t13 VDD.t30 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X956 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t24 Transmission_Gate_Layout_9.VOUT.t67 VDD.t53 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X957 IN5 EN.t180 Transmission_Gate_Layout_9.VIN.t50 VSS.t231 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X958 IN8 Transmission_Gate_Layout_20.CLKB.t24 Transmission_Gate_Layout_5.VIN.t70 VDD.t135 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X959 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t24 Transmission_Gate_Layout_11.VIN.t18 VDD.t5 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X960 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLK.t99 Transmission_Gate_Layout_9.VIN.t26 VSS.t89 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X961 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t50 Transmission_Gate_Layout_1.VIN.t10 VSS.t19 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X962 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t51 Transmission_Gate_Layout_2.VIN.t15 VSS.t25 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X963 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK.t100 Transmission_Gate_Layout_3.VIN.t141 VSS.t46 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X964 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t101 Transmission_Gate_Layout_9.VOUT.t90 VSS.t56 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X965 VDD Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.t4 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.t3 VDD.t141 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X966 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t47 Transmission_Gate_Layout_9.VOUT.t45 VSS.t162 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X967 Transmission_Gate_Layout_9.VIN EN.t181 IN5.t3 VSS.t296 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X968 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t25 IN2.t4 VDD.t251 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X969 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t24 IN7.t14 VDD.t35 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X970 Transmission_Gate_Layout_10.VIN EN.t182 IN3.t37 VSS.t220 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X971 Transmission_Gate_Layout_19.CLKB EN.t183 VSS.t293 VSS.t292 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X972 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLK.t104 VDD.t181 VDD.t180 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X973 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t25 OUT.t4 VDD.t17 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X974 IN8 EN.t184 Transmission_Gate_Layout_5.VIN.t86 VSS.t218 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X975 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t105 Transmission_Gate_Layout_11.VIN.t41 VSS.t126 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X976 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t106 Transmission_Gate_Layout_2.VIN.t101 VSS.t112 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X977 OUT Transmission_Gate_Layout_12.CLKB.t26 Transmission_Gate_Layout_12.VIN.t28 VDD.t94 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X978 VDD Transmission_Gate_Layout_3.CLK.t48 Transmission_Gate_Layout_0.CLKB.t2 VDD.t185 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X979 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t25 IN8.t23 VDD.t136 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X980 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t107 Transmission_Gate_Layout_11.VIN.t39 VSS.t126 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X981 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t25 Transmission_Gate_Layout_9.VOUT.t68 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X982 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t27 Transmission_Gate_Layout_3.VIN.t35 VDD.t144 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X983 OUT Transmission_Gate_Layout_13.CLKB.t26 Transmission_Gate_Layout_13.VIN.t14 VDD.t18 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X984 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t25 IN7.t15 VDD.t36 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X985 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t25 Transmission_Gate_Layout_10.VIN.t41 VDD.t73 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X986 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB.t26 Transmission_Gate_Layout_9.VOUT.t69 VDD.t55 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X987 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t22 Transmission_Gate_Layout_13.VIN.t82 VDD.t75 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X988 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t23 Transmission_Gate_Layout_1.VIN.t56 VDD.t59 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X989 Transmission_Gate_Layout_17.CLKB EN.t185 VSS.t295 VSS.t294 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X990 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t26 IN8.t9 VDD.t137 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X991 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLKB.t25 Transmission_Gate_Layout_11.VIN.t17 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X992 VSS Transmission_Gate_Layout_12.CLK.t26 Transmission_Gate_Layout_12.CLKB.t3 VSS.t183 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X993 IN5 EN.t186 Transmission_Gate_Layout_9.VIN.t49 VSS.t229 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X994 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t102 Transmission_Gate_Layout_4.VIN.t35 VSS.t71 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X995 Transmission_Gate_Layout_5.VIN EN.t187 IN8.t29 VSS.t289 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X996 VSS EN.t188 Transmission_Gate_Layout_20.CLKB.t3 VSS.t283 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X997 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t103 Transmission_Gate_Layout_2.VIN.t135 VSS.t55 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X998 VDD EN.t189 Transmission_Gate_Layout_18.CLKB.t1 VDD.t99 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X999 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t108 Transmission_Gate_Layout_5.VIN.t48 VSS.t113 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1000 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t104 Transmission_Gate_Layout_10.VIN.t54 VSS.t43 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1001 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t49 Transmission_Gate_Layout_13.VIN.t110 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1002 Transmission_Gate_Layout_9.VIN EN.t190 IN5.t1 VSS.t224 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1003 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t26 IN7.t16 VDD.t32 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1004 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t105 Transmission_Gate_Layout_1.VIN.t138 VSS.t70 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1005 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t106 Transmission_Gate_Layout_10.VIN.t53 VSS.t90 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1006 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t24 Transmission_Gate_Layout_9.VOUT.t3 VDD.t61 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1007 IN1 EN.t191 Transmission_Gate_Layout_6.VIN.t74 VSS.t288 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1008 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_11.CLK.t109 VDD.t179 VDD.t178 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1009 VSS Transmission_Gate_Layout_3.CLK.t50 Transmission_Gate_Layout_0.CLKB.t3 VSS.t166 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1010 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t23 Transmission_Gate_Layout_2.VIN.t75 VDD.t78 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1011 Transmission_Gate_Layout_16.CLKB EN.t192 VSS.t287 VSS.t225 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1012 IN5 EN.t193 Transmission_Gate_Layout_9.VIN.t48 VSS.t227 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1013 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t110 Transmission_Gate_Layout_9.VOUT.t11 VSS.t125 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1014 OUT Transmission_Gate_Layout_13.CLK.t29 Transmission_Gate_Layout_13.VIN.t7 VSS.t8 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1015 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t24 Transmission_Gate_Layout_12.VIN.t131 VDD.t58 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1016 Transmission_Gate_Layout_6.VIN EN.t194 IN1.t29 VSS.t222 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1017 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT Transmission_Gate_Layout_12.CLK.t27 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.t1 VDD.t222 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1018 OUT Transmission_Gate_Layout_13.CLKB.t27 Transmission_Gate_Layout_13.VIN.t66 VDD.t16 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1019 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t107 Transmission_Gate_Layout_1.VIN.t139 VSS.t53 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1020 IN6 EN.t195 Transmission_Gate_Layout_8.VIN.t87 VSS.t230 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1021 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t25 Transmission_Gate_Layout_9.VOUT.t4 VDD.t62 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1022 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLK.t52 Transmission_Gate_Layout_1.VIN.t11 VSS.t27 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1023 IN3 Transmission_Gate_Layout_14.CLKB.t27 Transmission_Gate_Layout_10.VIN.t2 VDD.t43 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1024 IN2 Transmission_Gate_Layout_18.CLKB.t26 Transmission_Gate_Layout_7.VIN.t44 VDD.t252 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1025 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t111 Transmission_Gate_Layout_8.VIN.t51 VSS.t117 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1026 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t24 Transmission_Gate_Layout_1.VIN.t57 VDD.t66 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1027 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_19.CLKB.t27 IN4.t21 VDD.t161 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1028 VSS Transmission_Gate_Layout_12.CLK.t28 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.t2 VSS.t65 nfet_03v3 ad=0.22p pd=1.88u as=0.13p ps=1.02u w=0.5u l=0.28u
X1029 IN1 EN.t196 Transmission_Gate_Layout_6.VIN.t73 VSS.t286 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1030 IN5 Transmission_Gate_Layout_15.CLKB.t24 Transmission_Gate_Layout_9.VIN.t79 VDD.t292 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1031 IN6 Transmission_Gate_Layout_21.CLKB.t25 Transmission_Gate_Layout_8.VIN.t3 VDD.t45 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1032 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t27 Transmission_Gate_Layout_8.VIN.t26 VDD.t10 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1033 IN5 Transmission_Gate_Layout_15.CLKB.t25 Transmission_Gate_Layout_9.VIN.t78 VDD.t294 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1034 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t112 Transmission_Gate_Layout_5.VIN.t47 VSS.t124 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1035 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t26 Transmission_Gate_Layout_2.VIN.t48 VDD.t71 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1036 Transmission_Gate_Layout_6.VIN EN.t197 IN1.t27 VSS.t219 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1037 Transmission_Gate_Layout_11.VIN EN.t198 IN4.t30 VSS.t282 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1038 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t108 Transmission_Gate_Layout_4.VIN.t32 VSS.t81 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1039 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t24 Transmission_Gate_Layout_2.VIN.t74 VDD.t76 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1040 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t25 Transmission_Gate_Layout_12.VIN.t68 VDD.t60 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1041 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t51 Transmission_Gate_Layout_9.VOUT.t79 VSS.t163 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1042 IN8 Transmission_Gate_Layout_20.CLKB.t27 Transmission_Gate_Layout_5.VIN.t58 VDD.t138 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1043 Transmission_Gate_Layout_13.CLK Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.t2 VDD.t239 VDD.t238 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1044 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB.t26 Transmission_Gate_Layout_9.VOUT.t5 VDD.t63 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1045 Transmission_Gate_Layout_16.CLKB EN.t199 VDD.t261 VDD.t85 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1046 IN5 Transmission_Gate_Layout_15.CLKB.t26 Transmission_Gate_Layout_9.VIN.t77 VDD.t293 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1047 VDD Transmission_Gate_Layout_9.CLK.t109 Transmission_Gate_Layout_6.CLKB.t0 VDD.t227 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1048 VSS EN.t200 Transmission_Gate_Layout_21.CLKB.t3 VSS.t283 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1049 OUT Transmission_Gate_Layout_12.CLK.t29 Transmission_Gate_Layout_12.VIN.t106 VSS.t187 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1050 VDD EN.t201 Transmission_Gate_Layout_14.CLKB.t0 VDD.t258 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1051 Transmission_Gate_Layout_5.VIN EN.t202 IN8.t28 VSS.t275 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1052 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t110 Transmission_Gate_Layout_2.VIN.t134 VSS.t46 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1053 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t27 Transmission_Gate_Layout_9.VIN.t2 VDD.t64 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1054 OUT Transmission_Gate_Layout_12.CLKB.t27 Transmission_Gate_Layout_12.VIN.t29 VDD.t95 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1055 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t28 IN8.t11 VDD.t132 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1056 VSS Transmission_Gate_Layout_1.CLK.t53 Transmission_Gate_Layout_2.CLKB.t3 VSS.t21 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1057 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t25 Transmission_Gate_Layout_13.VIN.t79 VDD.t74 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1058 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT C1.t3 VDD.t205 VDD.t149 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1059 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t111 Transmission_Gate_Layout_2.VIN.t133 VSS.t48 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1060 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t27 IN2.t2 VDD.t253 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1061 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_9.CLK.t112 VSS.t246 VSS.t78 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1062 IN7 Transmission_Gate_Layout_17.CLKB.t27 Transmission_Gate_Layout_4.VIN.t26 VDD.t34 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1063 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t54 Transmission_Gate_Layout_12.VIN.t13 VSS.t31 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1064 IN1 EN.t203 Transmission_Gate_Layout_6.VIN.t72 VSS.t216 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1065 Transmission_Gate_Layout_5.VIN EN.t204 IN8.t27 VSS.t238 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1066 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t26 Transmission_Gate_Layout_2.VIN.t117 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1067 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t25 Transmission_Gate_Layout_9.VOUT.t121 VDD.t52 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1068 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_20.CLKB.t29 IN8.t12 VDD.t133 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1069 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t26 IN6.t4 VDD.t46 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1070 Transmission_Gate_Layout_6.VIN EN.t205 IN1.t25 VSS.t217 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1071 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT Transmission_Gate_Layout_1.CLK.t55 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.t3 VDD.t27 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1072 IN8 EN.t206 Transmission_Gate_Layout_5.VIN.t85 VSS.t279 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1073 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t52 Transmission_Gate_Layout_13.VIN.t115 VSS.t165 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1074 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t27 IN5.t26 VDD.t291 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1075 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t22 Transmission_Gate_Layout_4.VIN.t17 VDD.t32 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1076 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLK.t113 Transmission_Gate_Layout_2.VIN.t132 VSS.t46 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1077 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLK.t114 VDD.t309 VDD.t24 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1078 IN8 EN.t207 Transmission_Gate_Layout_5.VIN.t84 VSS.t221 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1079 IN3 EN.t208 Transmission_Gate_Layout_10.VIN.t76 VSS.t280 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1080 VDD Transmission_Gate_Layout_3.CLK.t53 Transmission_Gate_Layout_0.CLKB.t5 VDD.t185 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1081 IN4 EN.t209 Transmission_Gate_Layout_11.VIN.t76 VSS.t281 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1082 IN6 EN.t210 Transmission_Gate_Layout_8.VIN.t86 VSS.t279 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1083 OUT Transmission_Gate_Layout_13.CLKB.t28 Transmission_Gate_Layout_13.VIN.t67 VDD.t18 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1084 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t23 IN1.t6 VDD.t244 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1085 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t30 OUT.t91 VSS.t188 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1086 IN3 Transmission_Gate_Layout_14.CLKB.t28 Transmission_Gate_Layout_10.VIN.t1 VDD.t44 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1087 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT C1.t4 VSS.t152 VSS.t99 nfet_03v3 ad=0.13p pd=1.02u as=0.22p ps=1.88u w=0.5u l=0.28u
X1088 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_1.CLKB.t26 Transmission_Gate_Layout_1.VIN.t59 VDD.t59 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1089 Transmission_Gate_Layout_5.VIN EN.t211 IN8.t24 VSS.t275 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1090 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t28 OUT.t29 VDD.t96 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1091 VDD EN.t212 Transmission_Gate_Layout_20.CLKB.t0 VDD.t161 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1092 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t28 Transmission_Gate_Layout_8.VIN.t25 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1093 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t56 Transmission_Gate_Layout_13.VIN.t25 VSS.t26 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1094 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_3.CLK.t54 Transmission_Gate_Layout_9.VOUT.t80 VSS.t173 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1095 IN4 EN.t213 Transmission_Gate_Layout_11.VIN.t75 VSS.t277 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1096 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t27 IN6.t5 VDD.t40 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1097 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t24 IN1.t5 VDD.t245 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1098 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t25 IN1.t4 VDD.t246 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1099 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t26 Transmission_Gate_Layout_2.VIN.t73 VDD.t72 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1100 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB.t28 IN6.t6 VDD.t41 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1101 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK.t55 Transmission_Gate_Layout_13.VIN.t116 VSS.t164 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1102 Transmission_Gate_Layout_9.CLK Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.t3 VSS.t94 VSS.t93 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X1103 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t113 Transmission_Gate_Layout_7.VIN.t2 VSS.t123 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1104 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t56 Transmission_Gate_Layout_3.VIN.t86 VSS.t170 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1105 OUT Transmission_Gate_Layout_12.CLK.t31 Transmission_Gate_Layout_12.VIN.t108 VSS.t186 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1106 Transmission_Gate_Layout_7.VIN EN.t214 IN2.t30 VSS.t278 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1107 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 Transmission_Gate_Layout_1.CLK.t57 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.t2 VDD.t28 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X1108 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t23 Transmission_Gate_Layout_3.VIN.t130 VDD.t105 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1109 OUT Transmission_Gate_Layout_13.CLK.t30 Transmission_Gate_Layout_13.VIN.t8 VSS.t9 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1110 Transmission_Gate_Layout_13.CLK Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.t3 VSS.t210 VSS.t209 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X1111 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t23 Transmission_Gate_Layout_4.VIN.t18 VDD.t31 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1112 Transmission_Gate_Layout_8.VIN EN.t215 IN6.t29 VSS.t275 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1113 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t28 Transmission_Gate_Layout_9.VIN.t1 VDD.t65 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1114 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB.t29 IN3.t12 VDD.t0 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1115 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t24 Transmission_Gate_Layout_1.VIN.t28 VDD.t34 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1116 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t115 Transmission_Gate_Layout_10.VIN.t49 VSS.t54 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1117 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t27 Transmission_Gate_Layout_12.VIN.t70 VDD.t60 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1118 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t28 IN7.t18 VDD.t35 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1119 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t58 Transmission_Gate_Layout_2.VIN.t17 VSS.t35 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1120 IN1 Transmission_Gate_Layout_16.CLKB.t26 Transmission_Gate_Layout_6.VIN.t56 VDD.t241 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1121 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t23 Transmission_Gate_Layout_1.VIN.t78 VDD.t115 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1122 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 B1.t4 VDD.t153 VDD.t110 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1123 Transmission_Gate_Layout_11.CLK Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.t3 VDD.t235 VDD.t234 pfet_03v3 ad=0.44p pd=2.88u as=0.44p ps=2.88u w=1u l=0.28u
X1124 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t59 Transmission_Gate_Layout_2.VIN.t18 VSS.t32 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1125 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t57 Transmission_Gate_Layout_12.VIN.t114 VSS.t171 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1126 Transmission_Gate_Layout_8.VIN EN.t216 IN6.t28 VSS.t275 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1127 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLK.t116 Transmission_Gate_Layout_10.VIN.t48 VSS.t47 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1128 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_17.CLKB.t29 IN7.t19 VDD.t36 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1129 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t24 Transmission_Gate_Layout_7.VIN.t60 VDD.t104 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1130 IN3 EN.t217 Transmission_Gate_Layout_10.VIN.t75 VSS.t276 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1131 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t58 Transmission_Gate_Layout_3.VIN.t87 VSS.t169 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1132 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t24 Transmission_Gate_Layout_1.VIN.t79 VDD.t116 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1133 IN6 EN.t218 Transmission_Gate_Layout_8.VIN.t85 VSS.t221 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1134 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_11.CLK.t114 Transmission_Gate_Layout_11.VIN.t38 VSS.t116 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1135 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLKB.t28 Transmission_Gate_Layout_3.VIN.t36 VDD.t5 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1136 Transmission_Gate_Layout_4.VIN EN.t219 IN7.t24 VSS.t274 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1137 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLK.t59 VDD.t225 VDD.t180 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1138 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t25 Transmission_Gate_Layout_7.VIN.t54 VDD.t103 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1139 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t115 Transmission_Gate_Layout_5.VIN.t46 VSS.t113 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1140 Transmission_Gate_Layout_8.VIN EN.t220 IN6.t26 VSS.t238 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1141 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t31 OUT.t50 VSS.t10 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1142 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t26 Transmission_Gate_Layout_9.VOUT.t120 VDD.t52 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1143 VDD EN.t221 Transmission_Gate_Layout_18.CLKB.t0 VDD.t99 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1144 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t25 Transmission_Gate_Layout_5.VIN.t19 VDD.t120 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1145 IN6 EN.t222 Transmission_Gate_Layout_8.VIN.t84 VSS.t218 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1146 IN2 EN.t223 Transmission_Gate_Layout_7.VIN.t76 VSS.t272 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1147 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t27 Transmission_Gate_Layout_2.VIN.t72 VDD.t73 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1148 Transmission_Gate_Layout_7.VIN EN.t224 IN2.t28 VSS.t273 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1149 Transmission_Gate_Layout_11.VIN EN.t225 IN4.t27 VSS.t267 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1150 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t27 Transmission_Gate_Layout_2.VIN.t118 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1151 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t27 Transmission_Gate_Layout_12.VIN.t130 VDD.t55 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1152 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t25 Transmission_Gate_Layout_1.VIN.t29 VDD.t33 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1153 VSS EN.t226 Transmission_Gate_Layout_14.CLKB.t3 VSS.t268 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1154 IN2 EN.t227 Transmission_Gate_Layout_7.VIN.t75 VSS.t271 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1155 IN4 EN.t228 Transmission_Gate_Layout_11.VIN.t74 VSS.t264 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1156 VDD Transmission_Gate_Layout_9.CLK.t117 Transmission_Gate_Layout_10.CLKB.t0 VDD.t19 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1157 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t60 Transmission_Gate_Layout_12.VIN.t115 VSS.t172 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1158 OUT Transmission_Gate_Layout_12.CLK.t32 Transmission_Gate_Layout_12.VIN.t109 VSS.t189 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1159 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_11.CLK.t116 Transmission_Gate_Layout_9.VOUT.t10 VSS.t115 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1160 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t60 Transmission_Gate_Layout_13.VIN.t28 VSS.t33 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1161 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB.t28 Transmission_Gate_Layout_12.VIN.t129 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1162 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLK.t61 VSS.t198 VSS.t158 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1163 IN5 Transmission_Gate_Layout_15.CLKB.t28 Transmission_Gate_Layout_9.VIN.t76 VDD.t292 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1164 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t27 Transmission_Gate_Layout_2.VIN.t49 VDD.t75 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1165 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t26 Transmission_Gate_Layout_1.VIN.t81 VDD.t119 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1166 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_9.CLK.t118 Transmission_Gate_Layout_6.VIN.t24 VSS.t47 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1167 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLKB.t29 OUT.t0 VDD.t54 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1168 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t26 Transmission_Gate_Layout_3.VIN.t116 VDD.t102 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1169 VSS Transmission_Gate_Layout_9.CLK.t119 Transmission_Gate_Layout_6.CLKB.t3 VSS.t13 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1170 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t27 Transmission_Gate_Layout_5.VIN.t21 VDD.t118 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1171 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_1.CLK.t61 Transmission_Gate_Layout_2.VIN.t20 VSS.t38 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1172 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t28 Transmission_Gate_Layout_12.VIN.t71 VDD.t62 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1173 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t26 Transmission_Gate_Layout_4.VIN.t21 VDD.t35 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1174 Transmission_Gate_Layout_8.VIN EN.t229 IN6.t24 VSS.t265 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1175 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB.t29 Transmission_Gate_Layout_8.VIN.t24 VDD.t57 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1176 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_3.CLK.t62 Transmission_Gate_Layout_12.VIN.t116 VSS.t160 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1177 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_2.CLKB.t28 Transmission_Gate_Layout_2.VIN.t71 VDD.t72 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1178 Transmission_Gate_Layout_7.VIN EN.t230 IN2.t26 VSS.t266 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1179 VDD Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.t4 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.t2 VDD.t141 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X1180 IN7 EN.t231 Transmission_Gate_Layout_4.VIN.t72 VSS.t261 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1181 IN2 Transmission_Gate_Layout_18.CLKB.t28 Transmission_Gate_Layout_7.VIN.t46 VDD.t178 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1182 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_6.CLKB.t28 Transmission_Gate_Layout_6.VIN.t16 VDD.t84 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1183 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB.t27 Transmission_Gate_Layout_3.VIN.t128 VDD.t101 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1184 IN6 Transmission_Gate_Layout_21.CLKB.t29 Transmission_Gate_Layout_8.VIN.t7 VDD.t42 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1185 Transmission_Gate_Layout_6.VIN EN.t232 IN1.t24 VSS.t262 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1186 IN2 EN.t233 Transmission_Gate_Layout_7.VIN.t73 VSS.t263 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1187 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB.t29 Transmission_Gate_Layout_13.VIN.t75 VDD.t71 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1188 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t117 Transmission_Gate_Layout_1.VIN.t90 VSS.t122 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1189 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.CLKB.t28 Transmission_Gate_Layout_1.VIN.t45 VDD.t113 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1190 IN3 EN.t234 Transmission_Gate_Layout_10.VIN.t74 VSS.t258 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1191 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_4.CLKB.t27 Transmission_Gate_Layout_4.VIN.t22 VDD.t36 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1192 Transmission_Gate_Layout_12.CLK Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.t3 VSS.t200 VSS.t199 nfet_03v3 ad=0.176p pd=1.68u as=0.176p ps=1.68u w=0.4u l=0.28u
X1193 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_3.CLK.t63 Transmission_Gate_Layout_3.VIN.t88 VSS.t157 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1194 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLK.t118 VSS.t119 VSS.t118 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1195 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.CLKB.t29 Transmission_Gate_Layout_9.VIN.t0 VDD.t66 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1196 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB.t28 Transmission_Gate_Layout_2.VIN.t50 VDD.t77 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1197 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t33 OUT.t94 VSS.t190 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1198 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t119 Transmission_Gate_Layout_8.VIN.t49 VSS.t117 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X1199 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_0.CLKB.t29 Transmission_Gate_Layout_9.VOUT.t117 VDD.t10 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1200 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLK.t120 Transmission_Gate_Layout_7.VIN.t1 VSS.t116 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1201 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t32 OUT.t49 VSS.t11 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1202 Transmission_Gate_Layout_11.VIN EN.t235 IN4.t25 VSS.t259 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1203 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLK.t120 Transmission_Gate_Layout_4.VIN.t31 VSS.t52 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1204 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.CLK.t33 OUT.t48 VSS.t12 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1205 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t28 Transmission_Gate_Layout_7.VIN.t62 VDD.t100 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1206 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t121 Transmission_Gate_Layout_1.VIN.t142 VSS.t53 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1207 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB.t29 Transmission_Gate_Layout_10.VIN.t45 VDD.t76 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1208 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t62 Transmission_Gate_Layout_12.VIN.t14 VSS.t39 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1209 IN4 EN.t236 Transmission_Gate_Layout_11.VIN.t73 VSS.t260 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1210 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t28 Transmission_Gate_Layout_1.VIN.t32 VDD.t29 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1211 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t28 Transmission_Gate_Layout_2.VIN.t119 VDD.t162 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1212 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK.t63 Transmission_Gate_Layout_12.VIN.t15 VSS.t34 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1213 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_7.CLKB.t29 Transmission_Gate_Layout_7.VIN.t57 VDD.t99 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1214 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_15.CLKB.t29 IN5.t24 VDD.t291 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1215 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK.t122 Transmission_Gate_Layout_9.VOUT.t89 VSS.t82 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1216 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB.t29 Transmission_Gate_Layout_12.VIN.t72 VDD.t63 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X1217 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB.t29 IN2.t0 VDD.t250 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1218 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t27 IN1.t2 VDD.t227 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X1219 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB.t29 Transmission_Gate_Layout_2.VIN.t54 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1220 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_1.CLK.t64 Transmission_Gate_Layout_13.VIN.t30 VSS.t40 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1221 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLK.t34 VDD.t15 VDD.t14 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1222 IN4 Transmission_Gate_Layout_19.CLKB.t28 Transmission_Gate_Layout_11.VIN.t70 VDD.t156 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1223 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t28 IN1.t1 VDD.t244 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1224 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.CLKB.t29 Transmission_Gate_Layout_5.VIN.t1 VDD.t114 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1225 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK.t123 Transmission_Gate_Layout_1.VIN.t143 VSS.t56 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1226 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_11.CLK.t121 Transmission_Gate_Layout_1.VIN.t89 VSS.t115 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1227 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB.t29 Transmission_Gate_Layout_1.VIN.t33 VDD.t30 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1228 Transmission_Gate_Layout_7.VIN EN.t237 IN2.t24 VSS.t255 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1229 IN3 EN.t238 Transmission_Gate_Layout_10.VIN.t73 VSS.t256 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1230 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLKB.t29 OUT.t30 VDD.t91 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1231 VSS Transmission_Gate_Layout_9.CLK.t124 Transmission_Gate_Layout_10.CLKB.t3 VSS.t13 nfet_03v3 ad=0.55p pd=3.38u as=0.55p ps=3.38u w=1.25u l=0.28u
X1232 Transmission_Gate_Layout_10.VIN EN.t239 IN3.t36 VSS.t257 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1233 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.CLK.t34 OUT.t95 VSS.t191 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X1234 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLK.t64 VDD.t226 VDD.t180 pfet_03v3 ad=1.1p pd=5.88u as=1.1p ps=5.88u w=2.5u l=0.28u
X1235 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB.t29 Transmission_Gate_Layout_3.VIN.t30 VDD.t87 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1236 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_11.CLK.t122 Transmission_Gate_Layout_5.VIN.t45 VSS.t114 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1237 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_11.CLK.t123 Transmission_Gate_Layout_8.VIN.t48 VSS.t113 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1238 IN4 Transmission_Gate_Layout_19.CLKB.t29 Transmission_Gate_Layout_11.VIN.t71 VDD.t158 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1239 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_16.CLKB.t29 IN1.t0 VDD.t245 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1240 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK.t124 Transmission_Gate_Layout_2.VIN.t100 VSS.t112 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1241 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB.t29 Transmission_Gate_Layout_13.VIN.t74 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
R0 Transmission_Gate_Layout_11.CLK.t28 Transmission_Gate_Layout_11.CLK.t60 82.9076
R1 Transmission_Gate_Layout_11.CLK.t109 Transmission_Gate_Layout_11.CLK.t28 82.9076
R2 Transmission_Gate_Layout_11.CLK.t62 Transmission_Gate_Layout_11.CLK.t91 82.9076
R3 Transmission_Gate_Layout_11.CLK.t15 Transmission_Gate_Layout_11.CLK.t62 82.9076
R4 Transmission_Gate_Layout_11.CLK.t38 Transmission_Gate_Layout_11.CLK.t84 82.9076
R5 Transmission_Gate_Layout_11.CLK.t4 Transmission_Gate_Layout_11.CLK.t38 82.9076
R6 Transmission_Gate_Layout_11.CLK.t53 Transmission_Gate_Layout_11.CLK.t104 82.9076
R7 Transmission_Gate_Layout_11.CLK.t21 Transmission_Gate_Layout_11.CLK.t53 82.9076
R8 Transmission_Gate_Layout_11.CLK.t29 Transmission_Gate_Layout_11.CLK.n10 56.4451
R9 Transmission_Gate_Layout_11.CLK.t46 Transmission_Gate_Layout_11.CLK.n67 56.4451
R10 Transmission_Gate_Layout_11.CLK.t69 Transmission_Gate_Layout_11.CLK.n38 56.4451
R11 Transmission_Gate_Layout_11.CLK.t36 Transmission_Gate_Layout_11.CLK.n96 56.4451
R12 Transmission_Gate_Layout_11.CLK.n29 Transmission_Gate_Layout_11.CLK.t109 49.7969
R13 Transmission_Gate_Layout_11.CLK.n86 Transmission_Gate_Layout_11.CLK.t15 49.7969
R14 Transmission_Gate_Layout_11.CLK.n57 Transmission_Gate_Layout_11.CLK.t4 49.7969
R15 Transmission_Gate_Layout_11.CLK.n115 Transmission_Gate_Layout_11.CLK.t21 49.7969
R16 Transmission_Gate_Layout_11.CLK.n4 Transmission_Gate_Layout_11.CLK.t97 39.7594
R17 Transmission_Gate_Layout_11.CLK.n61 Transmission_Gate_Layout_11.CLK.t80 39.7594
R18 Transmission_Gate_Layout_11.CLK.n32 Transmission_Gate_Layout_11.CLK.t7 39.7594
R19 Transmission_Gate_Layout_11.CLK.n90 Transmission_Gate_Layout_11.CLK.t105 39.7594
R20 Transmission_Gate_Layout_11.CLK.n12 Transmission_Gate_Layout_11.CLK.n11 35.0405
R21 Transmission_Gate_Layout_11.CLK.n28 Transmission_Gate_Layout_11.CLK.n27 35.0405
R22 Transmission_Gate_Layout_11.CLK.n69 Transmission_Gate_Layout_11.CLK.n68 35.0405
R23 Transmission_Gate_Layout_11.CLK.n85 Transmission_Gate_Layout_11.CLK.n84 35.0405
R24 Transmission_Gate_Layout_11.CLK.n40 Transmission_Gate_Layout_11.CLK.n39 35.0405
R25 Transmission_Gate_Layout_11.CLK.n56 Transmission_Gate_Layout_11.CLK.n55 35.0405
R26 Transmission_Gate_Layout_11.CLK.n98 Transmission_Gate_Layout_11.CLK.n97 35.0405
R27 Transmission_Gate_Layout_11.CLK.n114 Transmission_Gate_Layout_11.CLK.n113 35.0405
R28 Transmission_Gate_Layout_11.CLK.n29 Transmission_Gate_Layout_11.CLK.t26 31.1559
R29 Transmission_Gate_Layout_11.CLK.n86 Transmission_Gate_Layout_11.CLK.t61 31.1559
R30 Transmission_Gate_Layout_11.CLK.n57 Transmission_Gate_Layout_11.CLK.t56 31.1559
R31 Transmission_Gate_Layout_11.CLK.n115 Transmission_Gate_Layout_11.CLK.t70 31.1559
R32 Transmission_Gate_Layout_11.CLK.n122 Transmission_Gate_Layout_11.CLK.n121 24.3453
R33 Transmission_Gate_Layout_11.CLK.n120 Transmission_Gate_Layout_11.CLK.t67 22.0309
R34 Transmission_Gate_Layout_11.CLK.t23 Transmission_Gate_Layout_11.CLK.n19 21.9005
R35 Transmission_Gate_Layout_11.CLK.n18 Transmission_Gate_Layout_11.CLK.t95 21.9005
R36 Transmission_Gate_Layout_11.CLK.n17 Transmission_Gate_Layout_11.CLK.t40 21.9005
R37 Transmission_Gate_Layout_11.CLK.n16 Transmission_Gate_Layout_11.CLK.t20 21.9005
R38 Transmission_Gate_Layout_11.CLK.n15 Transmission_Gate_Layout_11.CLK.t78 21.9005
R39 Transmission_Gate_Layout_11.CLK.n14 Transmission_Gate_Layout_11.CLK.t63 21.9005
R40 Transmission_Gate_Layout_11.CLK.n13 Transmission_Gate_Layout_11.CLK.t8 21.9005
R41 Transmission_Gate_Layout_11.CLK.n11 Transmission_Gate_Layout_11.CLK.t75 21.9005
R42 Transmission_Gate_Layout_11.CLK.n12 Transmission_Gate_Layout_11.CLK.t76 21.9005
R43 Transmission_Gate_Layout_11.CLK.n68 Transmission_Gate_Layout_11.CLK.t99 21.9005
R44 Transmission_Gate_Layout_11.CLK.n69 Transmission_Gate_Layout_11.CLK.t3 21.9005
R45 Transmission_Gate_Layout_11.CLK.n70 Transmission_Gate_Layout_11.CLK.t73 21.9005
R46 Transmission_Gate_Layout_11.CLK.n71 Transmission_Gate_Layout_11.CLK.t54 21.9005
R47 Transmission_Gate_Layout_11.CLK.n72 Transmission_Gate_Layout_11.CLK.t121 21.9005
R48 Transmission_Gate_Layout_11.CLK.n73 Transmission_Gate_Layout_11.CLK.t112 21.9005
R49 Transmission_Gate_Layout_11.CLK.n74 Transmission_Gate_Layout_11.CLK.t83 21.9005
R50 Transmission_Gate_Layout_11.CLK.n75 Transmission_Gate_Layout_11.CLK.t33 21.9005
R51 Transmission_Gate_Layout_11.CLK.t12 Transmission_Gate_Layout_11.CLK.n76 21.9005
R52 Transmission_Gate_Layout_11.CLK.n39 Transmission_Gate_Layout_11.CLK.t35 21.9005
R53 Transmission_Gate_Layout_11.CLK.n40 Transmission_Gate_Layout_11.CLK.t111 21.9005
R54 Transmission_Gate_Layout_11.CLK.n41 Transmission_Gate_Layout_11.CLK.t17 21.9005
R55 Transmission_Gate_Layout_11.CLK.n42 Transmission_Gate_Layout_11.CLK.t22 21.9005
R56 Transmission_Gate_Layout_11.CLK.n43 Transmission_Gate_Layout_11.CLK.t59 21.9005
R57 Transmission_Gate_Layout_11.CLK.n44 Transmission_Gate_Layout_11.CLK.t65 21.9005
R58 Transmission_Gate_Layout_11.CLK.n45 Transmission_Gate_Layout_11.CLK.t55 21.9005
R59 Transmission_Gate_Layout_11.CLK.n46 Transmission_Gate_Layout_11.CLK.t90 21.9005
R60 Transmission_Gate_Layout_11.CLK.t98 Transmission_Gate_Layout_11.CLK.n47 21.9005
R61 Transmission_Gate_Layout_11.CLK.t68 Transmission_Gate_Layout_11.CLK.n105 21.9005
R62 Transmission_Gate_Layout_11.CLK.n104 Transmission_Gate_Layout_11.CLK.t106 21.9005
R63 Transmission_Gate_Layout_11.CLK.n103 Transmission_Gate_Layout_11.CLK.t14 21.9005
R64 Transmission_Gate_Layout_11.CLK.n102 Transmission_Gate_Layout_11.CLK.t18 21.9005
R65 Transmission_Gate_Layout_11.CLK.n101 Transmission_Gate_Layout_11.CLK.t58 21.9005
R66 Transmission_Gate_Layout_11.CLK.n100 Transmission_Gate_Layout_11.CLK.t64 21.9005
R67 Transmission_Gate_Layout_11.CLK.n99 Transmission_Gate_Layout_11.CLK.t103 21.9005
R68 Transmission_Gate_Layout_11.CLK.n97 Transmission_Gate_Layout_11.CLK.t118 21.9005
R69 Transmission_Gate_Layout_11.CLK.n98 Transmission_Gate_Layout_11.CLK.t11 21.9005
R70 Transmission_Gate_Layout_11.CLK.n20 Transmission_Gate_Layout_11.CLK.t23 21.5094
R71 Transmission_Gate_Layout_11.CLK.n21 Transmission_Gate_Layout_11.CLK.t95 21.5094
R72 Transmission_Gate_Layout_11.CLK.n22 Transmission_Gate_Layout_11.CLK.t40 21.5094
R73 Transmission_Gate_Layout_11.CLK.n23 Transmission_Gate_Layout_11.CLK.t20 21.5094
R74 Transmission_Gate_Layout_11.CLK.n24 Transmission_Gate_Layout_11.CLK.t78 21.5094
R75 Transmission_Gate_Layout_11.CLK.n25 Transmission_Gate_Layout_11.CLK.t63 21.5094
R76 Transmission_Gate_Layout_11.CLK.n26 Transmission_Gate_Layout_11.CLK.t8 21.5094
R77 Transmission_Gate_Layout_11.CLK.n28 Transmission_Gate_Layout_11.CLK.t75 21.5094
R78 Transmission_Gate_Layout_11.CLK.n27 Transmission_Gate_Layout_11.CLK.t76 21.5094
R79 Transmission_Gate_Layout_11.CLK.n85 Transmission_Gate_Layout_11.CLK.t99 21.5094
R80 Transmission_Gate_Layout_11.CLK.n84 Transmission_Gate_Layout_11.CLK.t3 21.5094
R81 Transmission_Gate_Layout_11.CLK.n83 Transmission_Gate_Layout_11.CLK.t73 21.5094
R82 Transmission_Gate_Layout_11.CLK.n82 Transmission_Gate_Layout_11.CLK.t54 21.5094
R83 Transmission_Gate_Layout_11.CLK.n81 Transmission_Gate_Layout_11.CLK.t121 21.5094
R84 Transmission_Gate_Layout_11.CLK.n80 Transmission_Gate_Layout_11.CLK.t112 21.5094
R85 Transmission_Gate_Layout_11.CLK.n79 Transmission_Gate_Layout_11.CLK.t83 21.5094
R86 Transmission_Gate_Layout_11.CLK.n78 Transmission_Gate_Layout_11.CLK.t33 21.5094
R87 Transmission_Gate_Layout_11.CLK.n77 Transmission_Gate_Layout_11.CLK.t12 21.5094
R88 Transmission_Gate_Layout_11.CLK.n56 Transmission_Gate_Layout_11.CLK.t35 21.5094
R89 Transmission_Gate_Layout_11.CLK.n55 Transmission_Gate_Layout_11.CLK.t111 21.5094
R90 Transmission_Gate_Layout_11.CLK.n54 Transmission_Gate_Layout_11.CLK.t17 21.5094
R91 Transmission_Gate_Layout_11.CLK.n53 Transmission_Gate_Layout_11.CLK.t22 21.5094
R92 Transmission_Gate_Layout_11.CLK.n52 Transmission_Gate_Layout_11.CLK.t59 21.5094
R93 Transmission_Gate_Layout_11.CLK.n51 Transmission_Gate_Layout_11.CLK.t65 21.5094
R94 Transmission_Gate_Layout_11.CLK.n50 Transmission_Gate_Layout_11.CLK.t55 21.5094
R95 Transmission_Gate_Layout_11.CLK.n49 Transmission_Gate_Layout_11.CLK.t90 21.5094
R96 Transmission_Gate_Layout_11.CLK.n48 Transmission_Gate_Layout_11.CLK.t98 21.5094
R97 Transmission_Gate_Layout_11.CLK.n106 Transmission_Gate_Layout_11.CLK.t68 21.5094
R98 Transmission_Gate_Layout_11.CLK.n107 Transmission_Gate_Layout_11.CLK.t106 21.5094
R99 Transmission_Gate_Layout_11.CLK.n108 Transmission_Gate_Layout_11.CLK.t14 21.5094
R100 Transmission_Gate_Layout_11.CLK.n109 Transmission_Gate_Layout_11.CLK.t18 21.5094
R101 Transmission_Gate_Layout_11.CLK.n110 Transmission_Gate_Layout_11.CLK.t58 21.5094
R102 Transmission_Gate_Layout_11.CLK.n111 Transmission_Gate_Layout_11.CLK.t64 21.5094
R103 Transmission_Gate_Layout_11.CLK.n112 Transmission_Gate_Layout_11.CLK.t103 21.5094
R104 Transmission_Gate_Layout_11.CLK.n114 Transmission_Gate_Layout_11.CLK.t118 21.5094
R105 Transmission_Gate_Layout_11.CLK.n113 Transmission_Gate_Layout_11.CLK.t11 21.5094
R106 Transmission_Gate_Layout_11.CLK.n120 Transmission_Gate_Layout_11.CLK.t43 21.3791
R107 Transmission_Gate_Layout_11.CLK.n121 Transmission_Gate_Layout_11.CLK.t48 21.3791
R108 Transmission_Gate_Layout_11.CLK.n20 Transmission_Gate_Layout_11.CLK.t89 20.988
R109 Transmission_Gate_Layout_11.CLK.n21 Transmission_Gate_Layout_11.CLK.t2 20.988
R110 Transmission_Gate_Layout_11.CLK.n22 Transmission_Gate_Layout_11.CLK.t39 20.988
R111 Transmission_Gate_Layout_11.CLK.n23 Transmission_Gate_Layout_11.CLK.t44 20.988
R112 Transmission_Gate_Layout_11.CLK.n24 Transmission_Gate_Layout_11.CLK.t81 20.988
R113 Transmission_Gate_Layout_11.CLK.n25 Transmission_Gate_Layout_11.CLK.t85 20.988
R114 Transmission_Gate_Layout_11.CLK.n26 Transmission_Gate_Layout_11.CLK.t120 20.988
R115 Transmission_Gate_Layout_11.CLK.n27 Transmission_Gate_Layout_11.CLK.t37 20.988
R116 Transmission_Gate_Layout_11.CLK.t26 Transmission_Gate_Layout_11.CLK.n28 20.988
R117 Transmission_Gate_Layout_11.CLK.n84 Transmission_Gate_Layout_11.CLK.t6 20.988
R118 Transmission_Gate_Layout_11.CLK.n83 Transmission_Gate_Layout_11.CLK.t42 20.988
R119 Transmission_Gate_Layout_11.CLK.n82 Transmission_Gate_Layout_11.CLK.t47 20.988
R120 Transmission_Gate_Layout_11.CLK.n81 Transmission_Gate_Layout_11.CLK.t82 20.988
R121 Transmission_Gate_Layout_11.CLK.n80 Transmission_Gate_Layout_11.CLK.t86 20.988
R122 Transmission_Gate_Layout_11.CLK.n79 Transmission_Gate_Layout_11.CLK.t79 20.988
R123 Transmission_Gate_Layout_11.CLK.n78 Transmission_Gate_Layout_11.CLK.t115 20.988
R124 Transmission_Gate_Layout_11.CLK.n77 Transmission_Gate_Layout_11.CLK.t117 20.988
R125 Transmission_Gate_Layout_11.CLK.t61 Transmission_Gate_Layout_11.CLK.n85 20.988
R126 Transmission_Gate_Layout_11.CLK.n55 Transmission_Gate_Layout_11.CLK.t119 20.988
R127 Transmission_Gate_Layout_11.CLK.n54 Transmission_Gate_Layout_11.CLK.t27 20.988
R128 Transmission_Gate_Layout_11.CLK.n53 Transmission_Gate_Layout_11.CLK.t96 20.988
R129 Transmission_Gate_Layout_11.CLK.n52 Transmission_Gate_Layout_11.CLK.t116 20.988
R130 Transmission_Gate_Layout_11.CLK.n51 Transmission_Gate_Layout_11.CLK.t66 20.988
R131 Transmission_Gate_Layout_11.CLK.n50 Transmission_Gate_Layout_11.CLK.t110 20.988
R132 Transmission_Gate_Layout_11.CLK.n49 Transmission_Gate_Layout_11.CLK.t5 20.988
R133 Transmission_Gate_Layout_11.CLK.n48 Transmission_Gate_Layout_11.CLK.t71 20.988
R134 Transmission_Gate_Layout_11.CLK.t56 Transmission_Gate_Layout_11.CLK.n56 20.988
R135 Transmission_Gate_Layout_11.CLK.n106 Transmission_Gate_Layout_11.CLK.t107 20.988
R136 Transmission_Gate_Layout_11.CLK.n107 Transmission_Gate_Layout_11.CLK.t124 20.988
R137 Transmission_Gate_Layout_11.CLK.n108 Transmission_Gate_Layout_11.CLK.t31 20.988
R138 Transmission_Gate_Layout_11.CLK.n109 Transmission_Gate_Layout_11.CLK.t102 20.988
R139 Transmission_Gate_Layout_11.CLK.n110 Transmission_Gate_Layout_11.CLK.t24 20.988
R140 Transmission_Gate_Layout_11.CLK.n111 Transmission_Gate_Layout_11.CLK.t87 20.988
R141 Transmission_Gate_Layout_11.CLK.n112 Transmission_Gate_Layout_11.CLK.t114 20.988
R142 Transmission_Gate_Layout_11.CLK.n113 Transmission_Gate_Layout_11.CLK.t19 20.988
R143 Transmission_Gate_Layout_11.CLK.t70 Transmission_Gate_Layout_11.CLK.n114 20.988
R144 Transmission_Gate_Layout_11.CLK.n121 Transmission_Gate_Layout_11.CLK.n120 20.8576
R145 Transmission_Gate_Layout_11.CLK.n5 Transmission_Gate_Layout_11.CLK.n4 20.8576
R146 Transmission_Gate_Layout_11.CLK.n6 Transmission_Gate_Layout_11.CLK.n5 20.8576
R147 Transmission_Gate_Layout_11.CLK.n7 Transmission_Gate_Layout_11.CLK.n6 20.8576
R148 Transmission_Gate_Layout_11.CLK.n8 Transmission_Gate_Layout_11.CLK.n7 20.8576
R149 Transmission_Gate_Layout_11.CLK.n9 Transmission_Gate_Layout_11.CLK.n8 20.8576
R150 Transmission_Gate_Layout_11.CLK.n10 Transmission_Gate_Layout_11.CLK.n9 20.8576
R151 Transmission_Gate_Layout_11.CLK.n67 Transmission_Gate_Layout_11.CLK.n66 20.8576
R152 Transmission_Gate_Layout_11.CLK.n66 Transmission_Gate_Layout_11.CLK.n65 20.8576
R153 Transmission_Gate_Layout_11.CLK.n65 Transmission_Gate_Layout_11.CLK.n64 20.8576
R154 Transmission_Gate_Layout_11.CLK.n64 Transmission_Gate_Layout_11.CLK.n63 20.8576
R155 Transmission_Gate_Layout_11.CLK.n63 Transmission_Gate_Layout_11.CLK.n62 20.8576
R156 Transmission_Gate_Layout_11.CLK.n62 Transmission_Gate_Layout_11.CLK.n61 20.8576
R157 Transmission_Gate_Layout_11.CLK.n38 Transmission_Gate_Layout_11.CLK.n37 20.8576
R158 Transmission_Gate_Layout_11.CLK.n37 Transmission_Gate_Layout_11.CLK.n36 20.8576
R159 Transmission_Gate_Layout_11.CLK.n36 Transmission_Gate_Layout_11.CLK.n35 20.8576
R160 Transmission_Gate_Layout_11.CLK.n35 Transmission_Gate_Layout_11.CLK.n34 20.8576
R161 Transmission_Gate_Layout_11.CLK.n34 Transmission_Gate_Layout_11.CLK.n33 20.8576
R162 Transmission_Gate_Layout_11.CLK.n33 Transmission_Gate_Layout_11.CLK.n32 20.8576
R163 Transmission_Gate_Layout_11.CLK.n91 Transmission_Gate_Layout_11.CLK.n90 20.8576
R164 Transmission_Gate_Layout_11.CLK.n92 Transmission_Gate_Layout_11.CLK.n91 20.8576
R165 Transmission_Gate_Layout_11.CLK.n93 Transmission_Gate_Layout_11.CLK.n92 20.8576
R166 Transmission_Gate_Layout_11.CLK.n94 Transmission_Gate_Layout_11.CLK.n93 20.8576
R167 Transmission_Gate_Layout_11.CLK.n95 Transmission_Gate_Layout_11.CLK.n94 20.8576
R168 Transmission_Gate_Layout_11.CLK.n96 Transmission_Gate_Layout_11.CLK.n95 20.8576
R169 Transmission_Gate_Layout_11.CLK.n19 Transmission_Gate_Layout_11.CLK.t97 20.5969
R170 Transmission_Gate_Layout_11.CLK.n18 Transmission_Gate_Layout_11.CLK.t41 20.5969
R171 Transmission_Gate_Layout_11.CLK.n17 Transmission_Gate_Layout_11.CLK.t113 20.5969
R172 Transmission_Gate_Layout_11.CLK.n16 Transmission_Gate_Layout_11.CLK.t94 20.5969
R173 Transmission_Gate_Layout_11.CLK.n15 Transmission_Gate_Layout_11.CLK.t32 20.5969
R174 Transmission_Gate_Layout_11.CLK.n14 Transmission_Gate_Layout_11.CLK.t9 20.5969
R175 Transmission_Gate_Layout_11.CLK.n13 Transmission_Gate_Layout_11.CLK.t77 20.5969
R176 Transmission_Gate_Layout_11.CLK.n12 Transmission_Gate_Layout_11.CLK.t30 20.5969
R177 Transmission_Gate_Layout_11.CLK.n11 Transmission_Gate_Layout_11.CLK.t29 20.5969
R178 Transmission_Gate_Layout_11.CLK.n68 Transmission_Gate_Layout_11.CLK.t46 20.5969
R179 Transmission_Gate_Layout_11.CLK.n69 Transmission_Gate_Layout_11.CLK.t74 20.5969
R180 Transmission_Gate_Layout_11.CLK.n70 Transmission_Gate_Layout_11.CLK.t25 20.5969
R181 Transmission_Gate_Layout_11.CLK.n71 Transmission_Gate_Layout_11.CLK.t122 20.5969
R182 Transmission_Gate_Layout_11.CLK.n72 Transmission_Gate_Layout_11.CLK.t72 20.5969
R183 Transmission_Gate_Layout_11.CLK.n73 Transmission_Gate_Layout_11.CLK.t52 20.5969
R184 Transmission_Gate_Layout_11.CLK.n74 Transmission_Gate_Layout_11.CLK.t34 20.5969
R185 Transmission_Gate_Layout_11.CLK.n76 Transmission_Gate_Layout_11.CLK.t80 20.5969
R186 Transmission_Gate_Layout_11.CLK.n75 Transmission_Gate_Layout_11.CLK.t108 20.5969
R187 Transmission_Gate_Layout_11.CLK.n47 Transmission_Gate_Layout_11.CLK.t7 20.5969
R188 Transmission_Gate_Layout_11.CLK.n45 Transmission_Gate_Layout_11.CLK.t88 20.5969
R189 Transmission_Gate_Layout_11.CLK.n44 Transmission_Gate_Layout_11.CLK.t101 20.5969
R190 Transmission_Gate_Layout_11.CLK.n43 Transmission_Gate_Layout_11.CLK.t93 20.5969
R191 Transmission_Gate_Layout_11.CLK.n42 Transmission_Gate_Layout_11.CLK.t57 20.5969
R192 Transmission_Gate_Layout_11.CLK.n41 Transmission_Gate_Layout_11.CLK.t50 20.5969
R193 Transmission_Gate_Layout_11.CLK.n40 Transmission_Gate_Layout_11.CLK.t16 20.5969
R194 Transmission_Gate_Layout_11.CLK.n39 Transmission_Gate_Layout_11.CLK.t69 20.5969
R195 Transmission_Gate_Layout_11.CLK.n46 Transmission_Gate_Layout_11.CLK.t123 20.5969
R196 Transmission_Gate_Layout_11.CLK.n98 Transmission_Gate_Layout_11.CLK.t45 20.5969
R197 Transmission_Gate_Layout_11.CLK.n99 Transmission_Gate_Layout_11.CLK.t10 20.5969
R198 Transmission_Gate_Layout_11.CLK.n100 Transmission_Gate_Layout_11.CLK.t100 20.5969
R199 Transmission_Gate_Layout_11.CLK.n101 Transmission_Gate_Layout_11.CLK.t92 20.5969
R200 Transmission_Gate_Layout_11.CLK.n102 Transmission_Gate_Layout_11.CLK.t51 20.5969
R201 Transmission_Gate_Layout_11.CLK.n103 Transmission_Gate_Layout_11.CLK.t49 20.5969
R202 Transmission_Gate_Layout_11.CLK.n104 Transmission_Gate_Layout_11.CLK.t13 20.5969
R203 Transmission_Gate_Layout_11.CLK.n105 Transmission_Gate_Layout_11.CLK.t105 20.5969
R204 Transmission_Gate_Layout_11.CLK.n97 Transmission_Gate_Layout_11.CLK.t36 20.5969
R205 Transmission_Gate_Layout_11.CLK.n19 Transmission_Gate_Layout_11.CLK.n18 19.4672
R206 Transmission_Gate_Layout_11.CLK.n18 Transmission_Gate_Layout_11.CLK.n17 19.4672
R207 Transmission_Gate_Layout_11.CLK.n17 Transmission_Gate_Layout_11.CLK.n16 19.4672
R208 Transmission_Gate_Layout_11.CLK.n16 Transmission_Gate_Layout_11.CLK.n15 19.4672
R209 Transmission_Gate_Layout_11.CLK.n15 Transmission_Gate_Layout_11.CLK.n14 19.4672
R210 Transmission_Gate_Layout_11.CLK.n14 Transmission_Gate_Layout_11.CLK.n13 19.4672
R211 Transmission_Gate_Layout_11.CLK.n13 Transmission_Gate_Layout_11.CLK.n12 19.4672
R212 Transmission_Gate_Layout_11.CLK.n21 Transmission_Gate_Layout_11.CLK.n20 19.4672
R213 Transmission_Gate_Layout_11.CLK.n22 Transmission_Gate_Layout_11.CLK.n21 19.4672
R214 Transmission_Gate_Layout_11.CLK.n23 Transmission_Gate_Layout_11.CLK.n22 19.4672
R215 Transmission_Gate_Layout_11.CLK.n24 Transmission_Gate_Layout_11.CLK.n23 19.4672
R216 Transmission_Gate_Layout_11.CLK.n25 Transmission_Gate_Layout_11.CLK.n24 19.4672
R217 Transmission_Gate_Layout_11.CLK.n26 Transmission_Gate_Layout_11.CLK.n25 19.4672
R218 Transmission_Gate_Layout_11.CLK.n27 Transmission_Gate_Layout_11.CLK.n26 19.4672
R219 Transmission_Gate_Layout_11.CLK.n70 Transmission_Gate_Layout_11.CLK.n69 19.4672
R220 Transmission_Gate_Layout_11.CLK.n71 Transmission_Gate_Layout_11.CLK.n70 19.4672
R221 Transmission_Gate_Layout_11.CLK.n72 Transmission_Gate_Layout_11.CLK.n71 19.4672
R222 Transmission_Gate_Layout_11.CLK.n73 Transmission_Gate_Layout_11.CLK.n72 19.4672
R223 Transmission_Gate_Layout_11.CLK.n74 Transmission_Gate_Layout_11.CLK.n73 19.4672
R224 Transmission_Gate_Layout_11.CLK.n75 Transmission_Gate_Layout_11.CLK.n74 19.4672
R225 Transmission_Gate_Layout_11.CLK.n76 Transmission_Gate_Layout_11.CLK.n75 19.4672
R226 Transmission_Gate_Layout_11.CLK.n84 Transmission_Gate_Layout_11.CLK.n83 19.4672
R227 Transmission_Gate_Layout_11.CLK.n83 Transmission_Gate_Layout_11.CLK.n82 19.4672
R228 Transmission_Gate_Layout_11.CLK.n82 Transmission_Gate_Layout_11.CLK.n81 19.4672
R229 Transmission_Gate_Layout_11.CLK.n81 Transmission_Gate_Layout_11.CLK.n80 19.4672
R230 Transmission_Gate_Layout_11.CLK.n80 Transmission_Gate_Layout_11.CLK.n79 19.4672
R231 Transmission_Gate_Layout_11.CLK.n79 Transmission_Gate_Layout_11.CLK.n78 19.4672
R232 Transmission_Gate_Layout_11.CLK.n78 Transmission_Gate_Layout_11.CLK.n77 19.4672
R233 Transmission_Gate_Layout_11.CLK.n41 Transmission_Gate_Layout_11.CLK.n40 19.4672
R234 Transmission_Gate_Layout_11.CLK.n42 Transmission_Gate_Layout_11.CLK.n41 19.4672
R235 Transmission_Gate_Layout_11.CLK.n43 Transmission_Gate_Layout_11.CLK.n42 19.4672
R236 Transmission_Gate_Layout_11.CLK.n44 Transmission_Gate_Layout_11.CLK.n43 19.4672
R237 Transmission_Gate_Layout_11.CLK.n45 Transmission_Gate_Layout_11.CLK.n44 19.4672
R238 Transmission_Gate_Layout_11.CLK.n46 Transmission_Gate_Layout_11.CLK.n45 19.4672
R239 Transmission_Gate_Layout_11.CLK.n47 Transmission_Gate_Layout_11.CLK.n46 19.4672
R240 Transmission_Gate_Layout_11.CLK.n55 Transmission_Gate_Layout_11.CLK.n54 19.4672
R241 Transmission_Gate_Layout_11.CLK.n54 Transmission_Gate_Layout_11.CLK.n53 19.4672
R242 Transmission_Gate_Layout_11.CLK.n53 Transmission_Gate_Layout_11.CLK.n52 19.4672
R243 Transmission_Gate_Layout_11.CLK.n52 Transmission_Gate_Layout_11.CLK.n51 19.4672
R244 Transmission_Gate_Layout_11.CLK.n51 Transmission_Gate_Layout_11.CLK.n50 19.4672
R245 Transmission_Gate_Layout_11.CLK.n50 Transmission_Gate_Layout_11.CLK.n49 19.4672
R246 Transmission_Gate_Layout_11.CLK.n49 Transmission_Gate_Layout_11.CLK.n48 19.4672
R247 Transmission_Gate_Layout_11.CLK.n105 Transmission_Gate_Layout_11.CLK.n104 19.4672
R248 Transmission_Gate_Layout_11.CLK.n104 Transmission_Gate_Layout_11.CLK.n103 19.4672
R249 Transmission_Gate_Layout_11.CLK.n103 Transmission_Gate_Layout_11.CLK.n102 19.4672
R250 Transmission_Gate_Layout_11.CLK.n102 Transmission_Gate_Layout_11.CLK.n101 19.4672
R251 Transmission_Gate_Layout_11.CLK.n101 Transmission_Gate_Layout_11.CLK.n100 19.4672
R252 Transmission_Gate_Layout_11.CLK.n100 Transmission_Gate_Layout_11.CLK.n99 19.4672
R253 Transmission_Gate_Layout_11.CLK.n99 Transmission_Gate_Layout_11.CLK.n98 19.4672
R254 Transmission_Gate_Layout_11.CLK.n107 Transmission_Gate_Layout_11.CLK.n106 19.4672
R255 Transmission_Gate_Layout_11.CLK.n108 Transmission_Gate_Layout_11.CLK.n107 19.4672
R256 Transmission_Gate_Layout_11.CLK.n109 Transmission_Gate_Layout_11.CLK.n108 19.4672
R257 Transmission_Gate_Layout_11.CLK.n110 Transmission_Gate_Layout_11.CLK.n109 19.4672
R258 Transmission_Gate_Layout_11.CLK.n111 Transmission_Gate_Layout_11.CLK.n110 19.4672
R259 Transmission_Gate_Layout_11.CLK.n112 Transmission_Gate_Layout_11.CLK.n111 19.4672
R260 Transmission_Gate_Layout_11.CLK.n113 Transmission_Gate_Layout_11.CLK.n112 19.4672
R261 Transmission_Gate_Layout_11.CLK.n4 Transmission_Gate_Layout_11.CLK.t41 18.9023
R262 Transmission_Gate_Layout_11.CLK.n5 Transmission_Gate_Layout_11.CLK.t113 18.9023
R263 Transmission_Gate_Layout_11.CLK.n6 Transmission_Gate_Layout_11.CLK.t94 18.9023
R264 Transmission_Gate_Layout_11.CLK.n7 Transmission_Gate_Layout_11.CLK.t32 18.9023
R265 Transmission_Gate_Layout_11.CLK.n8 Transmission_Gate_Layout_11.CLK.t9 18.9023
R266 Transmission_Gate_Layout_11.CLK.n9 Transmission_Gate_Layout_11.CLK.t77 18.9023
R267 Transmission_Gate_Layout_11.CLK.n10 Transmission_Gate_Layout_11.CLK.t30 18.9023
R268 Transmission_Gate_Layout_11.CLK.n67 Transmission_Gate_Layout_11.CLK.t74 18.9023
R269 Transmission_Gate_Layout_11.CLK.n66 Transmission_Gate_Layout_11.CLK.t25 18.9023
R270 Transmission_Gate_Layout_11.CLK.n65 Transmission_Gate_Layout_11.CLK.t122 18.9023
R271 Transmission_Gate_Layout_11.CLK.n64 Transmission_Gate_Layout_11.CLK.t72 18.9023
R272 Transmission_Gate_Layout_11.CLK.n63 Transmission_Gate_Layout_11.CLK.t52 18.9023
R273 Transmission_Gate_Layout_11.CLK.n62 Transmission_Gate_Layout_11.CLK.t34 18.9023
R274 Transmission_Gate_Layout_11.CLK.n61 Transmission_Gate_Layout_11.CLK.t108 18.9023
R275 Transmission_Gate_Layout_11.CLK.n33 Transmission_Gate_Layout_11.CLK.t88 18.9023
R276 Transmission_Gate_Layout_11.CLK.n34 Transmission_Gate_Layout_11.CLK.t101 18.9023
R277 Transmission_Gate_Layout_11.CLK.n35 Transmission_Gate_Layout_11.CLK.t93 18.9023
R278 Transmission_Gate_Layout_11.CLK.n36 Transmission_Gate_Layout_11.CLK.t57 18.9023
R279 Transmission_Gate_Layout_11.CLK.n37 Transmission_Gate_Layout_11.CLK.t50 18.9023
R280 Transmission_Gate_Layout_11.CLK.n38 Transmission_Gate_Layout_11.CLK.t16 18.9023
R281 Transmission_Gate_Layout_11.CLK.n32 Transmission_Gate_Layout_11.CLK.t123 18.9023
R282 Transmission_Gate_Layout_11.CLK.n96 Transmission_Gate_Layout_11.CLK.t45 18.9023
R283 Transmission_Gate_Layout_11.CLK.n95 Transmission_Gate_Layout_11.CLK.t10 18.9023
R284 Transmission_Gate_Layout_11.CLK.n94 Transmission_Gate_Layout_11.CLK.t100 18.9023
R285 Transmission_Gate_Layout_11.CLK.n93 Transmission_Gate_Layout_11.CLK.t92 18.9023
R286 Transmission_Gate_Layout_11.CLK.n92 Transmission_Gate_Layout_11.CLK.t51 18.9023
R287 Transmission_Gate_Layout_11.CLK.n91 Transmission_Gate_Layout_11.CLK.t49 18.9023
R288 Transmission_Gate_Layout_11.CLK.n90 Transmission_Gate_Layout_11.CLK.t13 18.9023
R289 Transmission_Gate_Layout_11.CLK.n116 Transmission_Gate_Layout_11.CLK.n115 16.4443
R290 Transmission_Gate_Layout_11.CLK.n58 Transmission_Gate_Layout_11.CLK.n57 16.4436
R291 Transmission_Gate_Layout_11.CLK.n30 Transmission_Gate_Layout_11.CLK.n29 16.4376
R292 Transmission_Gate_Layout_11.CLK.n87 Transmission_Gate_Layout_11.CLK.n86 16.4376
R293 Transmission_Gate_Layout_11.CLK.n0 Transmission_Gate_Layout_11.CLK.n2 11.313
R294 Transmission_Gate_Layout_11.CLK.n123 Transmission_Gate_Layout_11.CLK.n122 7.84627
R295 Transmission_Gate_Layout_11.CLK.n126 Transmission_Gate_Layout_11.CLK.n124 7.70137
R296 Transmission_Gate_Layout_11.CLK.n123 Transmission_Gate_Layout_11.CLK 7.5343
R297 Transmission_Gate_Layout_11.CLK.n59 Transmission_Gate_Layout_11.CLK.n58 5.33122
R298 Transmission_Gate_Layout_11.CLK.n117 Transmission_Gate_Layout_11.CLK.n116 5.33034
R299 Transmission_Gate_Layout_11.CLK.n126 Transmission_Gate_Layout_11.CLK.n125 4.70224
R300 Transmission_Gate_Layout_11.CLK.n1 Transmission_Gate_Layout_11.CLK.n0 0.903854
R301 Transmission_Gate_Layout_11.CLK.n3 Transmission_Gate_Layout_11.CLK.n2 0.902576
R302 Transmission_Gate_Layout_11.CLK.n59 Transmission_Gate_Layout_11.CLK.n2 4.5005
R303 Transmission_Gate_Layout_11.CLK.n0 Transmission_Gate_Layout_11.CLK.n117 4.5005
R304 Transmission_Gate_Layout_11.CLK.n119 Transmission_Gate_Layout_11.CLK.n118 4.5005
R305 Transmission_Gate_Layout_11.CLK.n87 Transmission_Gate_Layout_11.CLK.n60 2.25186
R306 Transmission_Gate_Layout_11.CLK.n31 Transmission_Gate_Layout_11.CLK.n30 2.25154
R307 Transmission_Gate_Layout_11.CLK.n89 Transmission_Gate_Layout_11.CLK.n88 2.24309
R308 Transmission_Gate_Layout_11.CLK.n127 Transmission_Gate_Layout_11.CLK.n123 1.2535
R309 Transmission_Gate_Layout_11.CLK.n3 Transmission_Gate_Layout_11.CLK.n89 0.00392645
R310 Transmission_Gate_Layout_11.CLK.n127 Transmission_Gate_Layout_11.CLK 0.493543
R311 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_11.CLK.n127 0.248978
R312 Transmission_Gate_Layout_11.CLK.n122 Transmission_Gate_Layout_11.CLK 0.147067
R313 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_11.CLK.n126 0.115935
R314 Transmission_Gate_Layout_11.CLK.n116 Transmission_Gate_Layout_11.CLK 0.0895398
R315 Transmission_Gate_Layout_11.CLK.n58 Transmission_Gate_Layout_11.CLK 0.0883538
R316 Transmission_Gate_Layout_11.CLK.n88 Transmission_Gate_Layout_11.CLK 0.0770183
R317 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_11.CLK.n119 0.0593683
R318 Transmission_Gate_Layout_11.CLK.n119 Transmission_Gate_Layout_11.CLK.n30 0.0335882
R319 Transmission_Gate_Layout_11.CLK.n117 Transmission_Gate_Layout_11.CLK.n31 0.0180708
R320 Transmission_Gate_Layout_11.CLK.n60 Transmission_Gate_Layout_11.CLK.n59 0.0180687
R321 Transmission_Gate_Layout_11.CLK.n88 Transmission_Gate_Layout_11.CLK.n87 0.0168265
R322 Transmission_Gate_Layout_11.CLK.n89 Transmission_Gate_Layout_11.CLK.n60 0.0158083
R323 Transmission_Gate_Layout_11.CLK.n118 Transmission_Gate_Layout_11.CLK.n31 0.0158062
R324 Transmission_Gate_Layout_11.CLK.n3 Transmission_Gate_Layout_11.CLK.n87 2.25612
R325 Transmission_Gate_Layout_11.CLK.n118 Transmission_Gate_Layout_11.CLK.n1 0.00304887
R326 Transmission_Gate_Layout_11.CLK.n1 Transmission_Gate_Layout_11.CLK.n30 1.50352
R327 Transmission_Gate_Layout_3.VIN.n212 Transmission_Gate_Layout_3.VIN 16.6454
R328 Transmission_Gate_Layout_3.VIN.n46 Transmission_Gate_Layout_3.VIN.t7 5.21612
R329 Transmission_Gate_Layout_3.VIN.n113 Transmission_Gate_Layout_3.VIN.n111 5.21612
R330 Transmission_Gate_Layout_3.VIN.n127 Transmission_Gate_Layout_3.VIN.t51 4.4609
R331 Transmission_Gate_Layout_3.VIN.n126 Transmission_Gate_Layout_3.VIN.t47 4.4609
R332 Transmission_Gate_Layout_3.VIN.n125 Transmission_Gate_Layout_3.VIN.t52 4.4609
R333 Transmission_Gate_Layout_3.VIN.n51 Transmission_Gate_Layout_3.VIN.n35 4.4609
R334 Transmission_Gate_Layout_3.VIN.n50 Transmission_Gate_Layout_3.VIN.n36 4.4609
R335 Transmission_Gate_Layout_3.VIN.n49 Transmission_Gate_Layout_3.VIN.n37 4.4609
R336 Transmission_Gate_Layout_3.VIN.n47 Transmission_Gate_Layout_3.VIN.t8 4.4609
R337 Transmission_Gate_Layout_3.VIN.n46 Transmission_Gate_Layout_3.VIN.t133 4.4609
R338 Transmission_Gate_Layout_3.VIN.n115 Transmission_Gate_Layout_3.VIN.n114 4.4609
R339 Transmission_Gate_Layout_3.VIN.n113 Transmission_Gate_Layout_3.VIN.n112 4.4609
R340 Transmission_Gate_Layout_3.VIN.n156 Transmission_Gate_Layout_3.VIN.n155 3.90572
R341 Transmission_Gate_Layout_3.VIN.n194 Transmission_Gate_Layout_3.VIN.n191 3.90572
R342 Transmission_Gate_Layout_3.VIN.n202 Transmission_Gate_Layout_3.VIN.n199 3.90572
R343 Transmission_Gate_Layout_3.VIN.n25 Transmission_Gate_Layout_3.VIN.n24 3.90572
R344 Transmission_Gate_Layout_3.VIN.n33 Transmission_Gate_Layout_3.VIN.n32 3.90572
R345 Transmission_Gate_Layout_3.VIN.n42 Transmission_Gate_Layout_3.VIN.n39 3.90572
R346 Transmission_Gate_Layout_3.VIN.n101 Transmission_Gate_Layout_3.VIN.n100 3.90572
R347 Transmission_Gate_Layout_3.VIN.n109 Transmission_Gate_Layout_3.VIN.n108 3.90572
R348 Transmission_Gate_Layout_3.VIN.n120 Transmission_Gate_Layout_3.VIN.n117 3.90572
R349 Transmission_Gate_Layout_3.VIN.n91 Transmission_Gate_Layout_3.VIN.n88 3.84485
R350 Transmission_Gate_Layout_3.VIN.n83 Transmission_Gate_Layout_3.VIN.n80 3.84485
R351 Transmission_Gate_Layout_3.VIN.n77 Transmission_Gate_Layout_3.VIN.n76 3.84485
R352 Transmission_Gate_Layout_3.VIN.n146 Transmission_Gate_Layout_3.VIN.n143 3.84485
R353 Transmission_Gate_Layout_3.VIN.n172 Transmission_Gate_Layout_3.VIN.n171 3.84485
R354 Transmission_Gate_Layout_3.VIN.n164 Transmission_Gate_Layout_3.VIN.n163 3.84485
R355 Transmission_Gate_Layout_3.VIN.n7 Transmission_Gate_Layout_3.VIN.n4 3.84485
R356 Transmission_Gate_Layout_3.VIN.n15 Transmission_Gate_Layout_3.VIN.n12 3.84485
R357 Transmission_Gate_Layout_3.VIN.n65 Transmission_Gate_Layout_3.VIN.n64 3.84485
R358 Transmission_Gate_Layout_3.VIN.n134 Transmission_Gate_Layout_3.VIN.t118 3.3285
R359 Transmission_Gate_Layout_3.VIN.n133 Transmission_Gate_Layout_3.VIN.t113 3.3285
R360 Transmission_Gate_Layout_3.VIN.n132 Transmission_Gate_Layout_3.VIN.t130 3.3285
R361 Transmission_Gate_Layout_3.VIN.n137 Transmission_Gate_Layout_3.VIN.n136 3.3285
R362 Transmission_Gate_Layout_3.VIN.n139 Transmission_Gate_Layout_3.VIN.n138 3.3285
R363 Transmission_Gate_Layout_3.VIN.n141 Transmission_Gate_Layout_3.VIN.n140 3.3285
R364 Transmission_Gate_Layout_3.VIN.n70 Transmission_Gate_Layout_3.VIN.t23 3.3285
R365 Transmission_Gate_Layout_3.VIN.n69 Transmission_Gate_Layout_3.VIN.t40 3.3285
R366 Transmission_Gate_Layout_3.VIN.n68 Transmission_Gate_Layout_3.VIN.t15 3.3285
R367 Transmission_Gate_Layout_3.VIN.n58 Transmission_Gate_Layout_3.VIN.n0 3.3285
R368 Transmission_Gate_Layout_3.VIN.n57 Transmission_Gate_Layout_3.VIN.n1 3.3285
R369 Transmission_Gate_Layout_3.VIN.n56 Transmission_Gate_Layout_3.VIN.n2 3.3285
R370 Transmission_Gate_Layout_3.VIN.n156 Transmission_Gate_Layout_3.VIN.n153 3.1505
R371 Transmission_Gate_Layout_3.VIN.n157 Transmission_Gate_Layout_3.VIN.n151 3.1505
R372 Transmission_Gate_Layout_3.VIN.n194 Transmission_Gate_Layout_3.VIN.n193 3.1505
R373 Transmission_Gate_Layout_3.VIN.n197 Transmission_Gate_Layout_3.VIN.n196 3.1505
R374 Transmission_Gate_Layout_3.VIN.n202 Transmission_Gate_Layout_3.VIN.n201 3.1505
R375 Transmission_Gate_Layout_3.VIN.n205 Transmission_Gate_Layout_3.VIN.n204 3.1505
R376 Transmission_Gate_Layout_3.VIN.n207 Transmission_Gate_Layout_3.VIN.n189 3.1505
R377 Transmission_Gate_Layout_3.VIN.n208 Transmission_Gate_Layout_3.VIN.n187 3.1505
R378 Transmission_Gate_Layout_3.VIN.n209 Transmission_Gate_Layout_3.VIN.n185 3.1505
R379 Transmission_Gate_Layout_3.VIN.n25 Transmission_Gate_Layout_3.VIN.n22 3.1505
R380 Transmission_Gate_Layout_3.VIN.n26 Transmission_Gate_Layout_3.VIN.n20 3.1505
R381 Transmission_Gate_Layout_3.VIN.n33 Transmission_Gate_Layout_3.VIN.n30 3.1505
R382 Transmission_Gate_Layout_3.VIN.n34 Transmission_Gate_Layout_3.VIN.n28 3.1505
R383 Transmission_Gate_Layout_3.VIN.n42 Transmission_Gate_Layout_3.VIN.n41 3.1505
R384 Transmission_Gate_Layout_3.VIN.n45 Transmission_Gate_Layout_3.VIN.n44 3.1505
R385 Transmission_Gate_Layout_3.VIN.n101 Transmission_Gate_Layout_3.VIN.n98 3.1505
R386 Transmission_Gate_Layout_3.VIN.n102 Transmission_Gate_Layout_3.VIN.n96 3.1505
R387 Transmission_Gate_Layout_3.VIN.n109 Transmission_Gate_Layout_3.VIN.n106 3.1505
R388 Transmission_Gate_Layout_3.VIN.n110 Transmission_Gate_Layout_3.VIN.n104 3.1505
R389 Transmission_Gate_Layout_3.VIN.n120 Transmission_Gate_Layout_3.VIN.n119 3.1505
R390 Transmission_Gate_Layout_3.VIN.n123 Transmission_Gate_Layout_3.VIN.n122 3.1505
R391 Transmission_Gate_Layout_3.VIN.n67 Transmission_Gate_Layout_3.VIN.n58 2.72398
R392 Transmission_Gate_Layout_3.VIN.n135 Transmission_Gate_Layout_3.VIN.n134 2.72398
R393 Transmission_Gate_Layout_3.VIN.n91 Transmission_Gate_Layout_3.VIN.n90 2.6005
R394 Transmission_Gate_Layout_3.VIN.n94 Transmission_Gate_Layout_3.VIN.n93 2.6005
R395 Transmission_Gate_Layout_3.VIN.n83 Transmission_Gate_Layout_3.VIN.n82 2.6005
R396 Transmission_Gate_Layout_3.VIN.n86 Transmission_Gate_Layout_3.VIN.n85 2.6005
R397 Transmission_Gate_Layout_3.VIN.n77 Transmission_Gate_Layout_3.VIN.n74 2.6005
R398 Transmission_Gate_Layout_3.VIN.n78 Transmission_Gate_Layout_3.VIN.n72 2.6005
R399 Transmission_Gate_Layout_3.VIN.n146 Transmission_Gate_Layout_3.VIN.n145 2.6005
R400 Transmission_Gate_Layout_3.VIN.n149 Transmission_Gate_Layout_3.VIN.n148 2.6005
R401 Transmission_Gate_Layout_3.VIN.n172 Transmission_Gate_Layout_3.VIN.n169 2.6005
R402 Transmission_Gate_Layout_3.VIN.n173 Transmission_Gate_Layout_3.VIN.n167 2.6005
R403 Transmission_Gate_Layout_3.VIN.n164 Transmission_Gate_Layout_3.VIN.n161 2.6005
R404 Transmission_Gate_Layout_3.VIN.n165 Transmission_Gate_Layout_3.VIN.n159 2.6005
R405 Transmission_Gate_Layout_3.VIN.n177 Transmission_Gate_Layout_3.VIN.n176 2.6005
R406 Transmission_Gate_Layout_3.VIN.n180 Transmission_Gate_Layout_3.VIN.n179 2.6005
R407 Transmission_Gate_Layout_3.VIN.n183 Transmission_Gate_Layout_3.VIN.n182 2.6005
R408 Transmission_Gate_Layout_3.VIN.n7 Transmission_Gate_Layout_3.VIN.n6 2.6005
R409 Transmission_Gate_Layout_3.VIN.n10 Transmission_Gate_Layout_3.VIN.n9 2.6005
R410 Transmission_Gate_Layout_3.VIN.n15 Transmission_Gate_Layout_3.VIN.n14 2.6005
R411 Transmission_Gate_Layout_3.VIN.n18 Transmission_Gate_Layout_3.VIN.n17 2.6005
R412 Transmission_Gate_Layout_3.VIN.n65 Transmission_Gate_Layout_3.VIN.n62 2.6005
R413 Transmission_Gate_Layout_3.VIN.n66 Transmission_Gate_Layout_3.VIN.n60 2.6005
R414 Transmission_Gate_Layout_3.VIN.n49 Transmission_Gate_Layout_3.VIN.n48 2.47941
R415 Transmission_Gate_Layout_3.VIN.n125 Transmission_Gate_Layout_3.VIN.n124 2.47941
R416 Transmission_Gate_Layout_3.VIN.n122 Transmission_Gate_Layout_3.VIN.t50 1.3109
R417 Transmission_Gate_Layout_3.VIN.n122 Transmission_Gate_Layout_3.VIN.n121 1.3109
R418 Transmission_Gate_Layout_3.VIN.n119 Transmission_Gate_Layout_3.VIN.t44 1.3109
R419 Transmission_Gate_Layout_3.VIN.n119 Transmission_Gate_Layout_3.VIN.n118 1.3109
R420 Transmission_Gate_Layout_3.VIN.n96 Transmission_Gate_Layout_3.VIN.t49 1.3109
R421 Transmission_Gate_Layout_3.VIN.n96 Transmission_Gate_Layout_3.VIN.n95 1.3109
R422 Transmission_Gate_Layout_3.VIN.n98 Transmission_Gate_Layout_3.VIN.t53 1.3109
R423 Transmission_Gate_Layout_3.VIN.n98 Transmission_Gate_Layout_3.VIN.n97 1.3109
R424 Transmission_Gate_Layout_3.VIN.n100 Transmission_Gate_Layout_3.VIN.t45 1.3109
R425 Transmission_Gate_Layout_3.VIN.n100 Transmission_Gate_Layout_3.VIN.n99 1.3109
R426 Transmission_Gate_Layout_3.VIN.n151 Transmission_Gate_Layout_3.VIN.t80 1.3109
R427 Transmission_Gate_Layout_3.VIN.n151 Transmission_Gate_Layout_3.VIN.n150 1.3109
R428 Transmission_Gate_Layout_3.VIN.n153 Transmission_Gate_Layout_3.VIN.t86 1.3109
R429 Transmission_Gate_Layout_3.VIN.n153 Transmission_Gate_Layout_3.VIN.n152 1.3109
R430 Transmission_Gate_Layout_3.VIN.n155 Transmission_Gate_Layout_3.VIN.t75 1.3109
R431 Transmission_Gate_Layout_3.VIN.n155 Transmission_Gate_Layout_3.VIN.n154 1.3109
R432 Transmission_Gate_Layout_3.VIN.n185 Transmission_Gate_Layout_3.VIN.t76 1.3109
R433 Transmission_Gate_Layout_3.VIN.n185 Transmission_Gate_Layout_3.VIN.n184 1.3109
R434 Transmission_Gate_Layout_3.VIN.n187 Transmission_Gate_Layout_3.VIN.t69 1.3109
R435 Transmission_Gate_Layout_3.VIN.n187 Transmission_Gate_Layout_3.VIN.n186 1.3109
R436 Transmission_Gate_Layout_3.VIN.n189 Transmission_Gate_Layout_3.VIN.t88 1.3109
R437 Transmission_Gate_Layout_3.VIN.n189 Transmission_Gate_Layout_3.VIN.n188 1.3109
R438 Transmission_Gate_Layout_3.VIN.n196 Transmission_Gate_Layout_3.VIN.t87 1.3109
R439 Transmission_Gate_Layout_3.VIN.n196 Transmission_Gate_Layout_3.VIN.n195 1.3109
R440 Transmission_Gate_Layout_3.VIN.n193 Transmission_Gate_Layout_3.VIN.t82 1.3109
R441 Transmission_Gate_Layout_3.VIN.n193 Transmission_Gate_Layout_3.VIN.n192 1.3109
R442 Transmission_Gate_Layout_3.VIN.n191 Transmission_Gate_Layout_3.VIN.t74 1.3109
R443 Transmission_Gate_Layout_3.VIN.n191 Transmission_Gate_Layout_3.VIN.n190 1.3109
R444 Transmission_Gate_Layout_3.VIN.n204 Transmission_Gate_Layout_3.VIN.t77 1.3109
R445 Transmission_Gate_Layout_3.VIN.n204 Transmission_Gate_Layout_3.VIN.n203 1.3109
R446 Transmission_Gate_Layout_3.VIN.n201 Transmission_Gate_Layout_3.VIN.t68 1.3109
R447 Transmission_Gate_Layout_3.VIN.n201 Transmission_Gate_Layout_3.VIN.n200 1.3109
R448 Transmission_Gate_Layout_3.VIN.n199 Transmission_Gate_Layout_3.VIN.t83 1.3109
R449 Transmission_Gate_Layout_3.VIN.n199 Transmission_Gate_Layout_3.VIN.n198 1.3109
R450 Transmission_Gate_Layout_3.VIN.n20 Transmission_Gate_Layout_3.VIN.t132 1.3109
R451 Transmission_Gate_Layout_3.VIN.n20 Transmission_Gate_Layout_3.VIN.n19 1.3109
R452 Transmission_Gate_Layout_3.VIN.n22 Transmission_Gate_Layout_3.VIN.t136 1.3109
R453 Transmission_Gate_Layout_3.VIN.n22 Transmission_Gate_Layout_3.VIN.n21 1.3109
R454 Transmission_Gate_Layout_3.VIN.n24 Transmission_Gate_Layout_3.VIN.t11 1.3109
R455 Transmission_Gate_Layout_3.VIN.n24 Transmission_Gate_Layout_3.VIN.n23 1.3109
R456 Transmission_Gate_Layout_3.VIN.n28 Transmission_Gate_Layout_3.VIN.t2 1.3109
R457 Transmission_Gate_Layout_3.VIN.n28 Transmission_Gate_Layout_3.VIN.n27 1.3109
R458 Transmission_Gate_Layout_3.VIN.n30 Transmission_Gate_Layout_3.VIN.t10 1.3109
R459 Transmission_Gate_Layout_3.VIN.n30 Transmission_Gate_Layout_3.VIN.n29 1.3109
R460 Transmission_Gate_Layout_3.VIN.n32 Transmission_Gate_Layout_3.VIN.t141 1.3109
R461 Transmission_Gate_Layout_3.VIN.n32 Transmission_Gate_Layout_3.VIN.n31 1.3109
R462 Transmission_Gate_Layout_3.VIN.n44 Transmission_Gate_Layout_3.VIN.t135 1.3109
R463 Transmission_Gate_Layout_3.VIN.n44 Transmission_Gate_Layout_3.VIN.n43 1.3109
R464 Transmission_Gate_Layout_3.VIN.n41 Transmission_Gate_Layout_3.VIN.t6 1.3109
R465 Transmission_Gate_Layout_3.VIN.n41 Transmission_Gate_Layout_3.VIN.n40 1.3109
R466 Transmission_Gate_Layout_3.VIN.n39 Transmission_Gate_Layout_3.VIN.t139 1.3109
R467 Transmission_Gate_Layout_3.VIN.n39 Transmission_Gate_Layout_3.VIN.n38 1.3109
R468 Transmission_Gate_Layout_3.VIN.n104 Transmission_Gate_Layout_3.VIN.t46 1.3109
R469 Transmission_Gate_Layout_3.VIN.n104 Transmission_Gate_Layout_3.VIN.n103 1.3109
R470 Transmission_Gate_Layout_3.VIN.n106 Transmission_Gate_Layout_3.VIN.t48 1.3109
R471 Transmission_Gate_Layout_3.VIN.n106 Transmission_Gate_Layout_3.VIN.n105 1.3109
R472 Transmission_Gate_Layout_3.VIN.n108 Transmission_Gate_Layout_3.VIN.t54 1.3109
R473 Transmission_Gate_Layout_3.VIN.n108 Transmission_Gate_Layout_3.VIN.n107 1.3109
R474 Transmission_Gate_Layout_3.VIN.n117 Transmission_Gate_Layout_3.VIN.t55 1.3109
R475 Transmission_Gate_Layout_3.VIN.n117 Transmission_Gate_Layout_3.VIN.n116 1.3109
R476 Transmission_Gate_Layout_3.VIN.n94 Transmission_Gate_Layout_3.VIN.n91 1.24485
R477 Transmission_Gate_Layout_3.VIN.n86 Transmission_Gate_Layout_3.VIN.n83 1.24485
R478 Transmission_Gate_Layout_3.VIN.n78 Transmission_Gate_Layout_3.VIN.n77 1.24485
R479 Transmission_Gate_Layout_3.VIN.n149 Transmission_Gate_Layout_3.VIN.n146 1.24485
R480 Transmission_Gate_Layout_3.VIN.n173 Transmission_Gate_Layout_3.VIN.n172 1.24485
R481 Transmission_Gate_Layout_3.VIN.n165 Transmission_Gate_Layout_3.VIN.n164 1.24485
R482 Transmission_Gate_Layout_3.VIN.n180 Transmission_Gate_Layout_3.VIN.n177 1.24485
R483 Transmission_Gate_Layout_3.VIN.n183 Transmission_Gate_Layout_3.VIN.n180 1.24485
R484 Transmission_Gate_Layout_3.VIN.n10 Transmission_Gate_Layout_3.VIN.n7 1.24485
R485 Transmission_Gate_Layout_3.VIN.n18 Transmission_Gate_Layout_3.VIN.n15 1.24485
R486 Transmission_Gate_Layout_3.VIN.n58 Transmission_Gate_Layout_3.VIN.n57 1.24485
R487 Transmission_Gate_Layout_3.VIN.n57 Transmission_Gate_Layout_3.VIN.n56 1.24485
R488 Transmission_Gate_Layout_3.VIN.n66 Transmission_Gate_Layout_3.VIN.n65 1.24485
R489 Transmission_Gate_Layout_3.VIN.n69 Transmission_Gate_Layout_3.VIN.n68 1.24485
R490 Transmission_Gate_Layout_3.VIN.n70 Transmission_Gate_Layout_3.VIN.n69 1.24485
R491 Transmission_Gate_Layout_3.VIN.n139 Transmission_Gate_Layout_3.VIN.n137 1.24485
R492 Transmission_Gate_Layout_3.VIN.n141 Transmission_Gate_Layout_3.VIN.n139 1.24485
R493 Transmission_Gate_Layout_3.VIN.n134 Transmission_Gate_Layout_3.VIN.n133 1.24485
R494 Transmission_Gate_Layout_3.VIN.n133 Transmission_Gate_Layout_3.VIN.n132 1.24485
R495 Transmission_Gate_Layout_3.VIN.n174 Transmission_Gate_Layout_3.VIN.n173 1.2018
R496 Transmission_Gate_Layout_3.VIN.n177 Transmission_Gate_Layout_3.VIN.n174 1.2018
R497 Transmission_Gate_Layout_3.VIN.n56 Transmission_Gate_Layout_3.VIN.n55 1.2018
R498 Transmission_Gate_Layout_3.VIN.n68 Transmission_Gate_Layout_3.VIN.n67 1.2018
R499 Transmission_Gate_Layout_3.VIN.n137 Transmission_Gate_Layout_3.VIN.n135 1.2018
R500 Transmission_Gate_Layout_3.VIN.n132 Transmission_Gate_Layout_3.VIN.n131 1.2018
R501 Transmission_Gate_Layout_3.VIN.n206 Transmission_Gate_Layout_3.VIN.n205 0.957239
R502 Transmission_Gate_Layout_3.VIN.n207 Transmission_Gate_Layout_3.VIN.n206 0.957239
R503 Transmission_Gate_Layout_3.VIN.n48 Transmission_Gate_Layout_3.VIN.n47 0.957239
R504 Transmission_Gate_Layout_3.VIN.n52 Transmission_Gate_Layout_3.VIN.n51 0.957239
R505 Transmission_Gate_Layout_3.VIN.n128 Transmission_Gate_Layout_3.VIN.n127 0.957239
R506 Transmission_Gate_Layout_3.VIN.n124 Transmission_Gate_Layout_3.VIN.n115 0.957239
R507 Transmission_Gate_Layout_3.VIN.n211 Transmission_Gate_Layout_3.VIN.n149 0.806587
R508 Transmission_Gate_Layout_3.VIN.n210 Transmission_Gate_Layout_3.VIN.n183 0.806587
R509 Transmission_Gate_Layout_3.VIN.n157 Transmission_Gate_Layout_3.VIN.n156 0.755717
R510 Transmission_Gate_Layout_3.VIN.n197 Transmission_Gate_Layout_3.VIN.n194 0.755717
R511 Transmission_Gate_Layout_3.VIN.n205 Transmission_Gate_Layout_3.VIN.n202 0.755717
R512 Transmission_Gate_Layout_3.VIN.n209 Transmission_Gate_Layout_3.VIN.n208 0.755717
R513 Transmission_Gate_Layout_3.VIN.n208 Transmission_Gate_Layout_3.VIN.n207 0.755717
R514 Transmission_Gate_Layout_3.VIN.n26 Transmission_Gate_Layout_3.VIN.n25 0.755717
R515 Transmission_Gate_Layout_3.VIN.n34 Transmission_Gate_Layout_3.VIN.n33 0.755717
R516 Transmission_Gate_Layout_3.VIN.n45 Transmission_Gate_Layout_3.VIN.n42 0.755717
R517 Transmission_Gate_Layout_3.VIN.n47 Transmission_Gate_Layout_3.VIN.n46 0.755717
R518 Transmission_Gate_Layout_3.VIN.n51 Transmission_Gate_Layout_3.VIN.n50 0.755717
R519 Transmission_Gate_Layout_3.VIN.n50 Transmission_Gate_Layout_3.VIN.n49 0.755717
R520 Transmission_Gate_Layout_3.VIN.n102 Transmission_Gate_Layout_3.VIN.n101 0.755717
R521 Transmission_Gate_Layout_3.VIN.n110 Transmission_Gate_Layout_3.VIN.n109 0.755717
R522 Transmission_Gate_Layout_3.VIN.n127 Transmission_Gate_Layout_3.VIN.n126 0.755717
R523 Transmission_Gate_Layout_3.VIN.n126 Transmission_Gate_Layout_3.VIN.n125 0.755717
R524 Transmission_Gate_Layout_3.VIN.n115 Transmission_Gate_Layout_3.VIN.n113 0.755717
R525 Transmission_Gate_Layout_3.VIN.n123 Transmission_Gate_Layout_3.VIN.n120 0.755717
R526 Transmission_Gate_Layout_3.VIN.n93 Transmission_Gate_Layout_3.VIN.t128 0.7285
R527 Transmission_Gate_Layout_3.VIN.n93 Transmission_Gate_Layout_3.VIN.n92 0.7285
R528 Transmission_Gate_Layout_3.VIN.n90 Transmission_Gate_Layout_3.VIN.t110 0.7285
R529 Transmission_Gate_Layout_3.VIN.n90 Transmission_Gate_Layout_3.VIN.n89 0.7285
R530 Transmission_Gate_Layout_3.VIN.n88 Transmission_Gate_Layout_3.VIN.t129 0.7285
R531 Transmission_Gate_Layout_3.VIN.n88 Transmission_Gate_Layout_3.VIN.n87 0.7285
R532 Transmission_Gate_Layout_3.VIN.n85 Transmission_Gate_Layout_3.VIN.t111 0.7285
R533 Transmission_Gate_Layout_3.VIN.n85 Transmission_Gate_Layout_3.VIN.n84 0.7285
R534 Transmission_Gate_Layout_3.VIN.n82 Transmission_Gate_Layout_3.VIN.t119 0.7285
R535 Transmission_Gate_Layout_3.VIN.n82 Transmission_Gate_Layout_3.VIN.n81 0.7285
R536 Transmission_Gate_Layout_3.VIN.n80 Transmission_Gate_Layout_3.VIN.t116 0.7285
R537 Transmission_Gate_Layout_3.VIN.n80 Transmission_Gate_Layout_3.VIN.n79 0.7285
R538 Transmission_Gate_Layout_3.VIN.n72 Transmission_Gate_Layout_3.VIN.t126 0.7285
R539 Transmission_Gate_Layout_3.VIN.n72 Transmission_Gate_Layout_3.VIN.n71 0.7285
R540 Transmission_Gate_Layout_3.VIN.n74 Transmission_Gate_Layout_3.VIN.t109 0.7285
R541 Transmission_Gate_Layout_3.VIN.n74 Transmission_Gate_Layout_3.VIN.n73 0.7285
R542 Transmission_Gate_Layout_3.VIN.n76 Transmission_Gate_Layout_3.VIN.t112 0.7285
R543 Transmission_Gate_Layout_3.VIN.n76 Transmission_Gate_Layout_3.VIN.n75 0.7285
R544 Transmission_Gate_Layout_3.VIN.n148 Transmission_Gate_Layout_3.VIN.t35 0.7285
R545 Transmission_Gate_Layout_3.VIN.n148 Transmission_Gate_Layout_3.VIN.n147 0.7285
R546 Transmission_Gate_Layout_3.VIN.n145 Transmission_Gate_Layout_3.VIN.t96 0.7285
R547 Transmission_Gate_Layout_3.VIN.n145 Transmission_Gate_Layout_3.VIN.n144 0.7285
R548 Transmission_Gate_Layout_3.VIN.n143 Transmission_Gate_Layout_3.VIN.t92 0.7285
R549 Transmission_Gate_Layout_3.VIN.n143 Transmission_Gate_Layout_3.VIN.n142 0.7285
R550 Transmission_Gate_Layout_3.VIN.n182 Transmission_Gate_Layout_3.VIN.t95 0.7285
R551 Transmission_Gate_Layout_3.VIN.n182 Transmission_Gate_Layout_3.VIN.n181 0.7285
R552 Transmission_Gate_Layout_3.VIN.n179 Transmission_Gate_Layout_3.VIN.t106 0.7285
R553 Transmission_Gate_Layout_3.VIN.n179 Transmission_Gate_Layout_3.VIN.n178 0.7285
R554 Transmission_Gate_Layout_3.VIN.n176 Transmission_Gate_Layout_3.VIN.t104 0.7285
R555 Transmission_Gate_Layout_3.VIN.n176 Transmission_Gate_Layout_3.VIN.n175 0.7285
R556 Transmission_Gate_Layout_3.VIN.n167 Transmission_Gate_Layout_3.VIN.t97 0.7285
R557 Transmission_Gate_Layout_3.VIN.n167 Transmission_Gate_Layout_3.VIN.n166 0.7285
R558 Transmission_Gate_Layout_3.VIN.n169 Transmission_Gate_Layout_3.VIN.t98 0.7285
R559 Transmission_Gate_Layout_3.VIN.n169 Transmission_Gate_Layout_3.VIN.n168 0.7285
R560 Transmission_Gate_Layout_3.VIN.n171 Transmission_Gate_Layout_3.VIN.t36 0.7285
R561 Transmission_Gate_Layout_3.VIN.n171 Transmission_Gate_Layout_3.VIN.n170 0.7285
R562 Transmission_Gate_Layout_3.VIN.n159 Transmission_Gate_Layout_3.VIN.t102 0.7285
R563 Transmission_Gate_Layout_3.VIN.n159 Transmission_Gate_Layout_3.VIN.n158 0.7285
R564 Transmission_Gate_Layout_3.VIN.n161 Transmission_Gate_Layout_3.VIN.t105 0.7285
R565 Transmission_Gate_Layout_3.VIN.n161 Transmission_Gate_Layout_3.VIN.n160 0.7285
R566 Transmission_Gate_Layout_3.VIN.n163 Transmission_Gate_Layout_3.VIN.t93 0.7285
R567 Transmission_Gate_Layout_3.VIN.n163 Transmission_Gate_Layout_3.VIN.n162 0.7285
R568 Transmission_Gate_Layout_3.VIN.n60 Transmission_Gate_Layout_3.VIN.t30 0.7285
R569 Transmission_Gate_Layout_3.VIN.n60 Transmission_Gate_Layout_3.VIN.n59 0.7285
R570 Transmission_Gate_Layout_3.VIN.n62 Transmission_Gate_Layout_3.VIN.t26 0.7285
R571 Transmission_Gate_Layout_3.VIN.n62 Transmission_Gate_Layout_3.VIN.n61 0.7285
R572 Transmission_Gate_Layout_3.VIN.n64 Transmission_Gate_Layout_3.VIN.t17 0.7285
R573 Transmission_Gate_Layout_3.VIN.n64 Transmission_Gate_Layout_3.VIN.n63 0.7285
R574 Transmission_Gate_Layout_3.VIN.n9 Transmission_Gate_Layout_3.VIN.t25 0.7285
R575 Transmission_Gate_Layout_3.VIN.n9 Transmission_Gate_Layout_3.VIN.n8 0.7285
R576 Transmission_Gate_Layout_3.VIN.n6 Transmission_Gate_Layout_3.VIN.t41 0.7285
R577 Transmission_Gate_Layout_3.VIN.n6 Transmission_Gate_Layout_3.VIN.n5 0.7285
R578 Transmission_Gate_Layout_3.VIN.n4 Transmission_Gate_Layout_3.VIN.t16 0.7285
R579 Transmission_Gate_Layout_3.VIN.n4 Transmission_Gate_Layout_3.VIN.n3 0.7285
R580 Transmission_Gate_Layout_3.VIN.n17 Transmission_Gate_Layout_3.VIN.t39 0.7285
R581 Transmission_Gate_Layout_3.VIN.n17 Transmission_Gate_Layout_3.VIN.n16 0.7285
R582 Transmission_Gate_Layout_3.VIN.n14 Transmission_Gate_Layout_3.VIN.t20 0.7285
R583 Transmission_Gate_Layout_3.VIN.n14 Transmission_Gate_Layout_3.VIN.n13 0.7285
R584 Transmission_Gate_Layout_3.VIN.n12 Transmission_Gate_Layout_3.VIN.t22 0.7285
R585 Transmission_Gate_Layout_3.VIN.n12 Transmission_Gate_Layout_3.VIN.n11 0.7285
R586 Transmission_Gate_Layout_3.VIN.n211 Transmission_Gate_Layout_3.VIN.n210 0.626587
R587 Transmission_Gate_Layout_3.VIN.n53 Transmission_Gate_Layout_3.VIN.n52 0.626587
R588 Transmission_Gate_Layout_3.VIN.n55 Transmission_Gate_Layout_3.VIN.n54 0.626587
R589 Transmission_Gate_Layout_3.VIN.n131 Transmission_Gate_Layout_3.VIN.n130 0.626587
R590 Transmission_Gate_Layout_3.VIN.n129 Transmission_Gate_Layout_3.VIN.n128 0.626587
R591 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.VIN.n70 0.607022
R592 Transmission_Gate_Layout_3.VIN.n130 Transmission_Gate_Layout_3.VIN.n94 0.575717
R593 Transmission_Gate_Layout_3.VIN.n131 Transmission_Gate_Layout_3.VIN.n86 0.575717
R594 Transmission_Gate_Layout_3.VIN.n135 Transmission_Gate_Layout_3.VIN.n78 0.575717
R595 Transmission_Gate_Layout_3.VIN.n174 Transmission_Gate_Layout_3.VIN.n165 0.575717
R596 Transmission_Gate_Layout_3.VIN.n55 Transmission_Gate_Layout_3.VIN.n10 0.575717
R597 Transmission_Gate_Layout_3.VIN.n54 Transmission_Gate_Layout_3.VIN.n18 0.575717
R598 Transmission_Gate_Layout_3.VIN.n67 Transmission_Gate_Layout_3.VIN.n66 0.575717
R599 Transmission_Gate_Layout_3.VIN.n212 Transmission_Gate_Layout_3.VIN.n141 0.459
R600 Transmission_Gate_Layout_3.VIN.n211 Transmission_Gate_Layout_3.VIN.n157 0.428978
R601 Transmission_Gate_Layout_3.VIN.n210 Transmission_Gate_Layout_3.VIN.n209 0.428978
R602 Transmission_Gate_Layout_3.VIN.n206 Transmission_Gate_Layout_3.VIN.n197 0.331152
R603 Transmission_Gate_Layout_3.VIN.n53 Transmission_Gate_Layout_3.VIN.n26 0.331152
R604 Transmission_Gate_Layout_3.VIN.n52 Transmission_Gate_Layout_3.VIN.n34 0.331152
R605 Transmission_Gate_Layout_3.VIN.n48 Transmission_Gate_Layout_3.VIN.n45 0.331152
R606 Transmission_Gate_Layout_3.VIN.n129 Transmission_Gate_Layout_3.VIN.n102 0.331152
R607 Transmission_Gate_Layout_3.VIN.n128 Transmission_Gate_Layout_3.VIN.n110 0.331152
R608 Transmission_Gate_Layout_3.VIN.n124 Transmission_Gate_Layout_3.VIN.n123 0.331152
R609 Transmission_Gate_Layout_3.VIN.n54 Transmission_Gate_Layout_3.VIN.n53 0.239196
R610 Transmission_Gate_Layout_3.VIN.n130 Transmission_Gate_Layout_3.VIN.n129 0.239196
R611 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.VIN.n211 0.192239
R612 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.VIN.n212 0.108109
R613 Transmission_Gate_Layout_7.VIN.n97 Transmission_Gate_Layout_7.VIN.n96 5.32175
R614 Transmission_Gate_Layout_7.VIN.n57 Transmission_Gate_Layout_7.VIN.t87 5.21612
R615 Transmission_Gate_Layout_7.VIN.n61 Transmission_Gate_Layout_7.VIN.n60 4.4609
R616 Transmission_Gate_Layout_7.VIN.n63 Transmission_Gate_Layout_7.VIN.n62 4.4609
R617 Transmission_Gate_Layout_7.VIN.n65 Transmission_Gate_Layout_7.VIN.n64 4.4609
R618 Transmission_Gate_Layout_7.VIN.n58 Transmission_Gate_Layout_7.VIN.t75 4.4609
R619 Transmission_Gate_Layout_7.VIN.n57 Transmission_Gate_Layout_7.VIN.t94 4.4609
R620 Transmission_Gate_Layout_7.VIN.n117 Transmission_Gate_Layout_7.VIN.n114 3.90572
R621 Transmission_Gate_Layout_7.VIN.n125 Transmission_Gate_Layout_7.VIN.n122 3.90572
R622 Transmission_Gate_Layout_7.VIN.n37 Transmission_Gate_Layout_7.VIN.n34 3.90572
R623 Transmission_Gate_Layout_7.VIN.n55 Transmission_Gate_Layout_7.VIN.n54 3.90572
R624 Transmission_Gate_Layout_7.VIN.n45 Transmission_Gate_Layout_7.VIN.n42 3.90572
R625 Transmission_Gate_Layout_7.VIN.n138 Transmission_Gate_Layout_7.VIN.n137 3.90572
R626 Transmission_Gate_Layout_7.VIN.n4 Transmission_Gate_Layout_7.VIN.n1 3.84485
R627 Transmission_Gate_Layout_7.VIN.n88 Transmission_Gate_Layout_7.VIN.n85 3.84485
R628 Transmission_Gate_Layout_7.VIN.n74 Transmission_Gate_Layout_7.VIN.n73 3.84485
R629 Transmission_Gate_Layout_7.VIN.n31 Transmission_Gate_Layout_7.VIN.n30 3.84485
R630 Transmission_Gate_Layout_7.VIN.n22 Transmission_Gate_Layout_7.VIN.n21 3.84485
R631 Transmission_Gate_Layout_7.VIN.n14 Transmission_Gate_Layout_7.VIN.n13 3.84485
R632 Transmission_Gate_Layout_7.VIN.n94 Transmission_Gate_Layout_7.VIN.t34 3.3285
R633 Transmission_Gate_Layout_7.VIN.n93 Transmission_Gate_Layout_7.VIN.t46 3.3285
R634 Transmission_Gate_Layout_7.VIN.n92 Transmission_Gate_Layout_7.VIN.t29 3.3285
R635 Transmission_Gate_Layout_7.VIN.n79 Transmission_Gate_Layout_7.VIN.n78 3.3285
R636 Transmission_Gate_Layout_7.VIN.n81 Transmission_Gate_Layout_7.VIN.n80 3.3285
R637 Transmission_Gate_Layout_7.VIN.n83 Transmission_Gate_Layout_7.VIN.n82 3.3285
R638 Transmission_Gate_Layout_7.VIN.n117 Transmission_Gate_Layout_7.VIN.n116 3.1505
R639 Transmission_Gate_Layout_7.VIN.n120 Transmission_Gate_Layout_7.VIN.n119 3.1505
R640 Transmission_Gate_Layout_7.VIN.n125 Transmission_Gate_Layout_7.VIN.n124 3.1505
R641 Transmission_Gate_Layout_7.VIN.n128 Transmission_Gate_Layout_7.VIN.n127 3.1505
R642 Transmission_Gate_Layout_7.VIN.n37 Transmission_Gate_Layout_7.VIN.n36 3.1505
R643 Transmission_Gate_Layout_7.VIN.n40 Transmission_Gate_Layout_7.VIN.n39 3.1505
R644 Transmission_Gate_Layout_7.VIN.n55 Transmission_Gate_Layout_7.VIN.n52 3.1505
R645 Transmission_Gate_Layout_7.VIN.n56 Transmission_Gate_Layout_7.VIN.n50 3.1505
R646 Transmission_Gate_Layout_7.VIN.n45 Transmission_Gate_Layout_7.VIN.n44 3.1505
R647 Transmission_Gate_Layout_7.VIN.n48 Transmission_Gate_Layout_7.VIN.n47 3.1505
R648 Transmission_Gate_Layout_7.VIN.n130 Transmission_Gate_Layout_7.VIN.n112 3.1505
R649 Transmission_Gate_Layout_7.VIN.n131 Transmission_Gate_Layout_7.VIN.n110 3.1505
R650 Transmission_Gate_Layout_7.VIN.n132 Transmission_Gate_Layout_7.VIN.n108 3.1505
R651 Transmission_Gate_Layout_7.VIN.n138 Transmission_Gate_Layout_7.VIN.n135 3.1505
R652 Transmission_Gate_Layout_7.VIN.n141 Transmission_Gate_Layout_7.VIN.n140 3.1505
R653 Transmission_Gate_Layout_7.VIN.n4 Transmission_Gate_Layout_7.VIN.n3 2.6005
R654 Transmission_Gate_Layout_7.VIN.n7 Transmission_Gate_Layout_7.VIN.n6 2.6005
R655 Transmission_Gate_Layout_7.VIN.n88 Transmission_Gate_Layout_7.VIN.n87 2.6005
R656 Transmission_Gate_Layout_7.VIN.n91 Transmission_Gate_Layout_7.VIN.n90 2.6005
R657 Transmission_Gate_Layout_7.VIN.n74 Transmission_Gate_Layout_7.VIN.n71 2.6005
R658 Transmission_Gate_Layout_7.VIN.n75 Transmission_Gate_Layout_7.VIN.n69 2.6005
R659 Transmission_Gate_Layout_7.VIN.n31 Transmission_Gate_Layout_7.VIN.n28 2.6005
R660 Transmission_Gate_Layout_7.VIN.n32 Transmission_Gate_Layout_7.VIN.n26 2.6005
R661 Transmission_Gate_Layout_7.VIN.n22 Transmission_Gate_Layout_7.VIN.n19 2.6005
R662 Transmission_Gate_Layout_7.VIN.n23 Transmission_Gate_Layout_7.VIN.n17 2.6005
R663 Transmission_Gate_Layout_7.VIN.n14 Transmission_Gate_Layout_7.VIN.n11 2.6005
R664 Transmission_Gate_Layout_7.VIN.n15 Transmission_Gate_Layout_7.VIN.n9 2.6005
R665 Transmission_Gate_Layout_7.VIN.n106 Transmission_Gate_Layout_7.VIN.n105 2.6005
R666 Transmission_Gate_Layout_7.VIN.n103 Transmission_Gate_Layout_7.VIN.n102 2.6005
R667 Transmission_Gate_Layout_7.VIN.n100 Transmission_Gate_Layout_7.VIN.n99 2.6005
R668 Transmission_Gate_Layout_7.VIN.n61 Transmission_Gate_Layout_7.VIN.n59 2.47941
R669 Transmission_Gate_Layout_7.VIN.n96 Transmission_Gate_Layout_7.VIN.n95 1.90239
R670 Transmission_Gate_Layout_7.VIN.n135 Transmission_Gate_Layout_7.VIN.t20 1.3109
R671 Transmission_Gate_Layout_7.VIN.n135 Transmission_Gate_Layout_7.VIN.n134 1.3109
R672 Transmission_Gate_Layout_7.VIN.n137 Transmission_Gate_Layout_7.VIN.t3 1.3109
R673 Transmission_Gate_Layout_7.VIN.n137 Transmission_Gate_Layout_7.VIN.n136 1.3109
R674 Transmission_Gate_Layout_7.VIN.n108 Transmission_Gate_Layout_7.VIN.t16 1.3109
R675 Transmission_Gate_Layout_7.VIN.n108 Transmission_Gate_Layout_7.VIN.n107 1.3109
R676 Transmission_Gate_Layout_7.VIN.n110 Transmission_Gate_Layout_7.VIN.t15 1.3109
R677 Transmission_Gate_Layout_7.VIN.n110 Transmission_Gate_Layout_7.VIN.n109 1.3109
R678 Transmission_Gate_Layout_7.VIN.n112 Transmission_Gate_Layout_7.VIN.t2 1.3109
R679 Transmission_Gate_Layout_7.VIN.n112 Transmission_Gate_Layout_7.VIN.n111 1.3109
R680 Transmission_Gate_Layout_7.VIN.n119 Transmission_Gate_Layout_7.VIN.t18 1.3109
R681 Transmission_Gate_Layout_7.VIN.n119 Transmission_Gate_Layout_7.VIN.n118 1.3109
R682 Transmission_Gate_Layout_7.VIN.n116 Transmission_Gate_Layout_7.VIN.t9 1.3109
R683 Transmission_Gate_Layout_7.VIN.n116 Transmission_Gate_Layout_7.VIN.n115 1.3109
R684 Transmission_Gate_Layout_7.VIN.n114 Transmission_Gate_Layout_7.VIN.t8 1.3109
R685 Transmission_Gate_Layout_7.VIN.n114 Transmission_Gate_Layout_7.VIN.n113 1.3109
R686 Transmission_Gate_Layout_7.VIN.n127 Transmission_Gate_Layout_7.VIN.t10 1.3109
R687 Transmission_Gate_Layout_7.VIN.n127 Transmission_Gate_Layout_7.VIN.n126 1.3109
R688 Transmission_Gate_Layout_7.VIN.n124 Transmission_Gate_Layout_7.VIN.t23 1.3109
R689 Transmission_Gate_Layout_7.VIN.n124 Transmission_Gate_Layout_7.VIN.n123 1.3109
R690 Transmission_Gate_Layout_7.VIN.n122 Transmission_Gate_Layout_7.VIN.t1 1.3109
R691 Transmission_Gate_Layout_7.VIN.n122 Transmission_Gate_Layout_7.VIN.n121 1.3109
R692 Transmission_Gate_Layout_7.VIN.n39 Transmission_Gate_Layout_7.VIN.t84 1.3109
R693 Transmission_Gate_Layout_7.VIN.n39 Transmission_Gate_Layout_7.VIN.n38 1.3109
R694 Transmission_Gate_Layout_7.VIN.n36 Transmission_Gate_Layout_7.VIN.t90 1.3109
R695 Transmission_Gate_Layout_7.VIN.n36 Transmission_Gate_Layout_7.VIN.n35 1.3109
R696 Transmission_Gate_Layout_7.VIN.n34 Transmission_Gate_Layout_7.VIN.t48 1.3109
R697 Transmission_Gate_Layout_7.VIN.n34 Transmission_Gate_Layout_7.VIN.n33 1.3109
R698 Transmission_Gate_Layout_7.VIN.n50 Transmission_Gate_Layout_7.VIN.t89 1.3109
R699 Transmission_Gate_Layout_7.VIN.n50 Transmission_Gate_Layout_7.VIN.n49 1.3109
R700 Transmission_Gate_Layout_7.VIN.n52 Transmission_Gate_Layout_7.VIN.t83 1.3109
R701 Transmission_Gate_Layout_7.VIN.n52 Transmission_Gate_Layout_7.VIN.n51 1.3109
R702 Transmission_Gate_Layout_7.VIN.n54 Transmission_Gate_Layout_7.VIN.t76 1.3109
R703 Transmission_Gate_Layout_7.VIN.n54 Transmission_Gate_Layout_7.VIN.n53 1.3109
R704 Transmission_Gate_Layout_7.VIN.n47 Transmission_Gate_Layout_7.VIN.t93 1.3109
R705 Transmission_Gate_Layout_7.VIN.n47 Transmission_Gate_Layout_7.VIN.n46 1.3109
R706 Transmission_Gate_Layout_7.VIN.n44 Transmission_Gate_Layout_7.VIN.t73 1.3109
R707 Transmission_Gate_Layout_7.VIN.n44 Transmission_Gate_Layout_7.VIN.n43 1.3109
R708 Transmission_Gate_Layout_7.VIN.n42 Transmission_Gate_Layout_7.VIN.t80 1.3109
R709 Transmission_Gate_Layout_7.VIN.n42 Transmission_Gate_Layout_7.VIN.n41 1.3109
R710 Transmission_Gate_Layout_7.VIN.n140 Transmission_Gate_Layout_7.VIN.t6 1.3109
R711 Transmission_Gate_Layout_7.VIN.n140 Transmission_Gate_Layout_7.VIN.n139 1.3109
R712 Transmission_Gate_Layout_7.VIN.n7 Transmission_Gate_Layout_7.VIN.n4 1.24485
R713 Transmission_Gate_Layout_7.VIN.n91 Transmission_Gate_Layout_7.VIN.n88 1.24485
R714 Transmission_Gate_Layout_7.VIN.n93 Transmission_Gate_Layout_7.VIN.n92 1.24485
R715 Transmission_Gate_Layout_7.VIN.n94 Transmission_Gate_Layout_7.VIN.n93 1.24485
R716 Transmission_Gate_Layout_7.VIN.n75 Transmission_Gate_Layout_7.VIN.n74 1.24485
R717 Transmission_Gate_Layout_7.VIN.n32 Transmission_Gate_Layout_7.VIN.n31 1.24485
R718 Transmission_Gate_Layout_7.VIN.n81 Transmission_Gate_Layout_7.VIN.n79 1.24485
R719 Transmission_Gate_Layout_7.VIN.n83 Transmission_Gate_Layout_7.VIN.n81 1.24485
R720 Transmission_Gate_Layout_7.VIN.n23 Transmission_Gate_Layout_7.VIN.n22 1.24485
R721 Transmission_Gate_Layout_7.VIN.n15 Transmission_Gate_Layout_7.VIN.n14 1.24485
R722 Transmission_Gate_Layout_7.VIN.n103 Transmission_Gate_Layout_7.VIN.n100 1.24485
R723 Transmission_Gate_Layout_7.VIN.n106 Transmission_Gate_Layout_7.VIN.n103 1.24485
R724 Transmission_Gate_Layout_7.VIN.n95 Transmission_Gate_Layout_7.VIN.n94 1.2018
R725 Transmission_Gate_Layout_7.VIN.n79 Transmission_Gate_Layout_7.VIN.n77 1.2018
R726 Transmission_Gate_Layout_7.VIN.n24 Transmission_Gate_Layout_7.VIN.n23 1.2018
R727 Transmission_Gate_Layout_7.VIN.n129 Transmission_Gate_Layout_7.VIN.n128 0.957239
R728 Transmission_Gate_Layout_7.VIN.n130 Transmission_Gate_Layout_7.VIN.n129 0.957239
R729 Transmission_Gate_Layout_7.VIN.n59 Transmission_Gate_Layout_7.VIN.n58 0.957239
R730 Transmission_Gate_Layout_7.VIN.n66 Transmission_Gate_Layout_7.VIN.n65 0.957239
R731 Transmission_Gate_Layout_7.VIN.n142 Transmission_Gate_Layout_7.VIN.n7 0.806587
R732 Transmission_Gate_Layout_7.VIN.n133 Transmission_Gate_Layout_7.VIN.n106 0.806587
R733 Transmission_Gate_Layout_7.VIN.n120 Transmission_Gate_Layout_7.VIN.n117 0.755717
R734 Transmission_Gate_Layout_7.VIN.n128 Transmission_Gate_Layout_7.VIN.n125 0.755717
R735 Transmission_Gate_Layout_7.VIN.n40 Transmission_Gate_Layout_7.VIN.n37 0.755717
R736 Transmission_Gate_Layout_7.VIN.n56 Transmission_Gate_Layout_7.VIN.n55 0.755717
R737 Transmission_Gate_Layout_7.VIN.n58 Transmission_Gate_Layout_7.VIN.n57 0.755717
R738 Transmission_Gate_Layout_7.VIN.n63 Transmission_Gate_Layout_7.VIN.n61 0.755717
R739 Transmission_Gate_Layout_7.VIN.n65 Transmission_Gate_Layout_7.VIN.n63 0.755717
R740 Transmission_Gate_Layout_7.VIN.n48 Transmission_Gate_Layout_7.VIN.n45 0.755717
R741 Transmission_Gate_Layout_7.VIN.n132 Transmission_Gate_Layout_7.VIN.n131 0.755717
R742 Transmission_Gate_Layout_7.VIN.n131 Transmission_Gate_Layout_7.VIN.n130 0.755717
R743 Transmission_Gate_Layout_7.VIN.n141 Transmission_Gate_Layout_7.VIN.n138 0.755717
R744 Transmission_Gate_Layout_7.VIN.n96 Transmission_Gate_Layout_7.VIN.n83 0.742022
R745 Transmission_Gate_Layout_7.VIN.n6 Transmission_Gate_Layout_7.VIN.t64 0.7285
R746 Transmission_Gate_Layout_7.VIN.n6 Transmission_Gate_Layout_7.VIN.n5 0.7285
R747 Transmission_Gate_Layout_7.VIN.n3 Transmission_Gate_Layout_7.VIN.t55 0.7285
R748 Transmission_Gate_Layout_7.VIN.n3 Transmission_Gate_Layout_7.VIN.n2 0.7285
R749 Transmission_Gate_Layout_7.VIN.n1 Transmission_Gate_Layout_7.VIN.t57 0.7285
R750 Transmission_Gate_Layout_7.VIN.n1 Transmission_Gate_Layout_7.VIN.n0 0.7285
R751 Transmission_Gate_Layout_7.VIN.n99 Transmission_Gate_Layout_7.VIN.t71 0.7285
R752 Transmission_Gate_Layout_7.VIN.n99 Transmission_Gate_Layout_7.VIN.n98 0.7285
R753 Transmission_Gate_Layout_7.VIN.n102 Transmission_Gate_Layout_7.VIN.t79 0.7285
R754 Transmission_Gate_Layout_7.VIN.n102 Transmission_Gate_Layout_7.VIN.n101 0.7285
R755 Transmission_Gate_Layout_7.VIN.n105 Transmission_Gate_Layout_7.VIN.t54 0.7285
R756 Transmission_Gate_Layout_7.VIN.n105 Transmission_Gate_Layout_7.VIN.n104 0.7285
R757 Transmission_Gate_Layout_7.VIN.n90 Transmission_Gate_Layout_7.VIN.t44 0.7285
R758 Transmission_Gate_Layout_7.VIN.n90 Transmission_Gate_Layout_7.VIN.n89 0.7285
R759 Transmission_Gate_Layout_7.VIN.n87 Transmission_Gate_Layout_7.VIN.t33 0.7285
R760 Transmission_Gate_Layout_7.VIN.n87 Transmission_Gate_Layout_7.VIN.n86 0.7285
R761 Transmission_Gate_Layout_7.VIN.n85 Transmission_Gate_Layout_7.VIN.t40 0.7285
R762 Transmission_Gate_Layout_7.VIN.n85 Transmission_Gate_Layout_7.VIN.n84 0.7285
R763 Transmission_Gate_Layout_7.VIN.n69 Transmission_Gate_Layout_7.VIN.t32 0.7285
R764 Transmission_Gate_Layout_7.VIN.n69 Transmission_Gate_Layout_7.VIN.n68 0.7285
R765 Transmission_Gate_Layout_7.VIN.n71 Transmission_Gate_Layout_7.VIN.t26 0.7285
R766 Transmission_Gate_Layout_7.VIN.n71 Transmission_Gate_Layout_7.VIN.n70 0.7285
R767 Transmission_Gate_Layout_7.VIN.n73 Transmission_Gate_Layout_7.VIN.t37 0.7285
R768 Transmission_Gate_Layout_7.VIN.n73 Transmission_Gate_Layout_7.VIN.n72 0.7285
R769 Transmission_Gate_Layout_7.VIN.n26 Transmission_Gate_Layout_7.VIN.t0 0.7285
R770 Transmission_Gate_Layout_7.VIN.n26 Transmission_Gate_Layout_7.VIN.n25 0.7285
R771 Transmission_Gate_Layout_7.VIN.n28 Transmission_Gate_Layout_7.VIN.t41 0.7285
R772 Transmission_Gate_Layout_7.VIN.n28 Transmission_Gate_Layout_7.VIN.n27 0.7285
R773 Transmission_Gate_Layout_7.VIN.n30 Transmission_Gate_Layout_7.VIN.t28 0.7285
R774 Transmission_Gate_Layout_7.VIN.n30 Transmission_Gate_Layout_7.VIN.n29 0.7285
R775 Transmission_Gate_Layout_7.VIN.n17 Transmission_Gate_Layout_7.VIN.t65 0.7285
R776 Transmission_Gate_Layout_7.VIN.n17 Transmission_Gate_Layout_7.VIN.n16 0.7285
R777 Transmission_Gate_Layout_7.VIN.n19 Transmission_Gate_Layout_7.VIN.t62 0.7285
R778 Transmission_Gate_Layout_7.VIN.n19 Transmission_Gate_Layout_7.VIN.n18 0.7285
R779 Transmission_Gate_Layout_7.VIN.n21 Transmission_Gate_Layout_7.VIN.t63 0.7285
R780 Transmission_Gate_Layout_7.VIN.n21 Transmission_Gate_Layout_7.VIN.n20 0.7285
R781 Transmission_Gate_Layout_7.VIN.n9 Transmission_Gate_Layout_7.VIN.t60 0.7285
R782 Transmission_Gate_Layout_7.VIN.n9 Transmission_Gate_Layout_7.VIN.n8 0.7285
R783 Transmission_Gate_Layout_7.VIN.n11 Transmission_Gate_Layout_7.VIN.t61 0.7285
R784 Transmission_Gate_Layout_7.VIN.n11 Transmission_Gate_Layout_7.VIN.n10 0.7285
R785 Transmission_Gate_Layout_7.VIN.n13 Transmission_Gate_Layout_7.VIN.t67 0.7285
R786 Transmission_Gate_Layout_7.VIN.n13 Transmission_Gate_Layout_7.VIN.n12 0.7285
R787 Transmission_Gate_Layout_7.VIN.n67 Transmission_Gate_Layout_7.VIN.n66 0.626587
R788 Transmission_Gate_Layout_7.VIN.n77 Transmission_Gate_Layout_7.VIN.n76 0.626587
R789 Transmission_Gate_Layout_7.VIN.n142 Transmission_Gate_Layout_7.VIN.n133 0.626587
R790 Transmission_Gate_Layout_7.VIN.n92 Transmission_Gate_Layout_7.VIN 0.607022
R791 Transmission_Gate_Layout_7.VIN.n95 Transmission_Gate_Layout_7.VIN.n91 0.575717
R792 Transmission_Gate_Layout_7.VIN.n76 Transmission_Gate_Layout_7.VIN.n75 0.575717
R793 Transmission_Gate_Layout_7.VIN.n77 Transmission_Gate_Layout_7.VIN.n32 0.575717
R794 Transmission_Gate_Layout_7.VIN.n24 Transmission_Gate_Layout_7.VIN.n15 0.575717
R795 Transmission_Gate_Layout_7.VIN.n97 Transmission_Gate_Layout_7.VIN.n24 0.570002
R796 Transmission_Gate_Layout_7.VIN.n100 Transmission_Gate_Layout_7.VIN.n97 0.562022
R797 Transmission_Gate_Layout_7.VIN.n133 Transmission_Gate_Layout_7.VIN.n132 0.428978
R798 Transmission_Gate_Layout_7.VIN.n142 Transmission_Gate_Layout_7.VIN.n141 0.428978
R799 Transmission_Gate_Layout_7.VIN.n129 Transmission_Gate_Layout_7.VIN.n120 0.331152
R800 Transmission_Gate_Layout_7.VIN.n67 Transmission_Gate_Layout_7.VIN.n40 0.331152
R801 Transmission_Gate_Layout_7.VIN.n59 Transmission_Gate_Layout_7.VIN.n56 0.331152
R802 Transmission_Gate_Layout_7.VIN.n66 Transmission_Gate_Layout_7.VIN.n48 0.331152
R803 Transmission_Gate_Layout_7.VIN.n76 Transmission_Gate_Layout_7.VIN.n67 0.239196
R804 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.VIN.n142 0.192239
R805 VSS.n166 VSS.n165 3274.56
R806 VSS.n361 VSS.t87 1488.24
R807 VSS.n361 VSS.t93 1488.24
R808 VSS.n341 VSS.t91 1488.24
R809 VSS.n341 VSS.t101 1488.24
R810 VSS.n341 VSS.t199 1488.24
R811 VSS.n341 VSS.t209 1488.24
R812 VSS.n615 VSS.n614 832.628
R813 VSS.n1155 VSS.n1154 519.736
R814 VSS.n341 VSS.n328 476.067
R815 VSS.n506 VSS.t28 372.284
R816 VSS.n506 VSS.t97 372.284
R817 VSS.n83 VSS.n82 286.959
R818 VSS.n328 VSS.n327 213.668
R819 VSS.n399 VSS.t49 161.036
R820 VSS.n397 VSS.t85 161.036
R821 VSS.n178 VSS.t65 161.036
R822 VSS.n176 VSS.t99 161.036
R823 VSS.n388 VSS.n387 97.5981
R824 VSS.n167 VSS.n166 97.5981
R825 VSS.n883 VSS.t220 95.3395
R826 VSS.n808 VSS.t163 95.3395
R827 VSS.n747 VSS.t34 95.3395
R828 VSS.n702 VSS.t25 95.3395
R829 VSS.n640 VSS.t3 95.3395
R830 VSS.n592 VSS.t187 95.3395
R831 VSS.n283 VSS.t11 95.3395
R832 VSS.n843 VSS.t280 82.6276
R833 VSS.n790 VSS.t171 82.6276
R834 VSS.n765 VSS.t36 82.6276
R835 VSS.n684 VSS.t20 82.6276
R836 VSS.n659 VSS.t157 82.6276
R837 VSS.n247 VSS.t188 82.6276
R838 VSS.n301 VSS.t7 82.6276
R839 VSS.n1389 VSS.t277 73.8269
R840 VSS.n1334 VSS.t227 73.8269
R841 VSS.n1281 VSS.t228 73.8269
R842 VSS.n1228 VSS.t216 73.8269
R843 VSS.n1183 VSS.t255 73.8269
R844 VSS.n10 VSS.t259 63.9833
R845 VSS.n1352 VSS.t299 63.9833
R846 VSS.n1299 VSS.t241 63.9833
R847 VSS.n1246 VSS.t219 63.9833
R848 VSS.n1165 VSS.t272 63.9833
R849 VSS.n840 VSS.t236 57.2039
R850 VSS.n787 VSS.t162 57.2039
R851 VSS.n768 VSS.t39 57.2039
R852 VSS.n681 VSS.t38 57.2039
R853 VSS.n662 VSS.t4 57.2039
R854 VSS.n250 VSS.t186 57.2039
R855 VSS.n304 VSS.t12 57.2039
R856 VSS.n1004 VSS.t70 53.874
R857 VSS.n1114 VSS.t128 53.874
R858 VSS.n104 VSS.t238 49.4761
R859 VSS.n944 VSS.t114 49.4761
R860 VSS.n1054 VSS.t54 49.4761
R861 VSS.n880 VSS.t276 44.492
R862 VSS.n811 VSS.t172 44.492
R863 VSS.n744 VSS.t27 44.492
R864 VSS.n705 VSS.t33 44.492
R865 VSS.n637 VSS.t156 44.492
R866 VSS.n595 VSS.t181 44.492
R867 VSS.n280 VSS.t6 44.492
R868 VSS.n7 VSS.t264 44.2963
R869 VSS.n1355 VSS.t215 44.2963
R870 VSS.n1302 VSS.t239 44.2963
R871 VSS.n1249 VSS.t286 44.2963
R872 VSS.n1162 VSS.t273 44.2963
R873 VSS.n907 VSS.t221 42.8794
R874 VSS.n962 VSS.t125 42.8794
R875 VSS.n989 VSS.t81 42.8794
R876 VSS.n1072 VSS.t55 42.8794
R877 VSS.n1099 VSS.t123 42.8794
R878 VSS.n114 VSS.t256 36.0174
R879 VSS.n803 VSS.t0 36.0174
R880 VSS.n753 VSS.t19 36.0174
R881 VSS.n697 VSS.t40 36.0174
R882 VSS.n647 VSS.t169 36.0174
R883 VSS.n587 VSS.t190 36.0174
R884 VSS.n289 VSS.t9 36.0174
R885 VSS.n1386 VSS.t282 34.4528
R886 VSS.n1331 VSS.t223 34.4528
R887 VSS.n1278 VSS.t274 34.4528
R888 VSS.n1225 VSS.t217 34.4528
R889 VSS.n1186 VSS.t263 34.4528
R890 VSS.n910 VSS.t265 29.6859
R891 VSS.n965 VSS.t113 29.6859
R892 VSS.n986 VSS.t56 29.6859
R893 VSS.n1075 VSS.t43 29.6859
R894 VSS.n1096 VSS.t112 29.6859
R895 VSS.n23 VSS.t242 27.8905
R896 VSS.n1340 VSS.t224 27.8905
R897 VSS.n1287 VSS.t252 27.8905
R898 VSS.n1234 VSS.t222 27.8905
R899 VSS.n1178 VSS.t232 27.8905
R900 VSS.t97 VSS.t105 23.5357
R901 VSS.n849 VSS.t257 23.3056
R902 VSS.n796 VSS.t173 23.3056
R903 VSS.n759 VSS.t31 23.3056
R904 VSS.n690 VSS.t32 23.3056
R905 VSS.n653 VSS.t165 23.3056
R906 VSS.n295 VSS.t5 23.3056
R907 VSS.n101 VSS.t230 23.0891
R908 VSS.n941 VSS.t133 23.0891
R909 VSS.n1010 VSS.t71 23.0891
R910 VSS.n1051 VSS.t46 23.0891
R911 VSS.n1138 VSS.t116 23.0891
R912 VSS.n895 VSS.t218 18.6913
R913 VSS.n950 VSS.t115 18.6913
R914 VSS.n1002 VSS.t52 18.6913
R915 VSS.n1060 VSS.t62 18.6913
R916 VSS.n1112 VSS.t130 18.6913
R917 VSS.n16 VSS.t260 18.0469
R918 VSS.n1346 VSS.t231 18.0469
R919 VSS.n1293 VSS.t240 18.0469
R920 VSS.n1240 VSS.t288 18.0469
R921 VSS.n1171 VSS.t278 18.0469
R922 VSS.n874 VSS.t251 14.831
R923 VSS.n817 VSS.t161 14.831
R924 VSS.n738 VSS.t16 14.831
R925 VSS.n711 VSS.t35 14.831
R926 VSS.n631 VSS.t164 14.831
R927 VSS.n601 VSS.t189 14.831
R928 VSS.n274 VSS.t10 14.831
R929 VSS.n901 VSS.t275 12.0945
R930 VSS.n956 VSS.t124 12.0945
R931 VSS.n995 VSS.t53 12.0945
R932 VSS.n1066 VSS.t90 12.0945
R933 VSS.n1105 VSS.t127 12.0945
R934 VSS.n1380 VSS.t281 11.4846
R935 VSS.n1325 VSS.t229 11.4846
R936 VSS.n1272 VSS.t261 11.4846
R937 VSS.n1219 VSS.t214 11.4846
R938 VSS.n1192 VSS.t266 11.4846
R939 VSS.n235 VSS.t182 10.5937
R940 VSS.n483 VSS.t202 9.32958
R941 VSS.n483 VSS.t96 9.32958
R942 VSS.n536 VSS.t204 9.32958
R943 VSS.n536 VSS.t207 9.32958
R944 VSS.n511 VSS.t212 9.32958
R945 VSS.n511 VSS.t73 9.32958
R946 VSS.n460 VSS.t154 9.32958
R947 VSS.n460 VSS.t211 9.32958
R948 VSS.n430 VSS.t206 9.32958
R949 VSS.n430 VSS.t213 9.32958
R950 VSS.n407 VSS.t2 9.32958
R951 VSS.n407 VSS.t111 9.32958
R952 VSS.n570 VSS.t104 9.32958
R953 VSS.n570 VSS.t201 9.32958
R954 VSS.n216 VSS.t75 9.32958
R955 VSS.n216 VSS.t208 9.32958
R956 VSS.n186 VSS.t110 9.32958
R957 VSS.n186 VSS.t155 9.32958
R958 VSS.n1341 VSS.n1339 9.13939
R959 VSS.n1288 VSS.n1286 9.13939
R960 VSS.n1235 VSS.n1233 9.13939
R961 VSS.n1179 VSS.n47 9.13939
R962 VSS.n951 VSS.n949 9.13939
R963 VSS.n1005 VSS.n1003 9.13939
R964 VSS.n1061 VSS.n1059 9.13939
R965 VSS.n1115 VSS.n1113 9.13939
R966 VSS.n896 VSS.n894 9.13939
R967 VSS.n290 VSS.n288 9.13939
R968 VSS.n590 VSS.n588 9.13939
R969 VSS.n648 VSS.n646 9.13939
R970 VSS.n700 VSS.n698 9.13939
R971 VSS.n754 VSS.n752 9.13939
R972 VSS.n806 VSS.n804 9.13939
R973 VSS.n169 VSS.n163 9.13939
R974 VSS.n169 VSS.n168 9.13939
R975 VSS.n179 VSS.n177 9.13939
R976 VSS.n196 VSS.n194 9.13939
R977 VSS.n194 VSS.n192 9.13939
R978 VSS.n227 VSS.n225 9.13939
R979 VSS.n225 VSS.n223 9.13939
R980 VSS.n575 VSS.n153 9.13939
R981 VSS.n390 VSS.n385 9.13939
R982 VSS.n390 VSS.n389 9.13939
R983 VSS.n400 VSS.n398 9.13939
R984 VSS.n417 VSS.n415 9.13939
R985 VSS.n415 VSS.n413 9.13939
R986 VSS.n468 VSS.n466 9.13939
R987 VSS.n441 VSS.n439 9.13939
R988 VSS.n439 VSS.n437 9.13939
R989 VSS.n521 VSS.n519 9.13939
R990 VSS.n519 VSS.n517 9.13939
R991 VSS.n478 VSS.n476 9.13939
R992 VSS.n547 VSS.n545 9.13939
R993 VSS.n545 VSS.n543 9.13939
R994 VSS.n115 VSS.n113 9.13939
R995 VSS.n95 VSS.t289 7.69671
R996 VSS.n935 VSS.t117 7.69671
R997 VSS.n1016 VSS.t82 7.69671
R998 VSS.n1045 VSS.t47 7.69671
R999 VSS.n1132 VSS.t131 7.69671
R1000 VSS.n343 VSS.t92 7.49789
R1001 VSS.n343 VSS.t102 7.49789
R1002 VSS.n500 VSS.t106 7.49789
R1003 VSS.n360 VSS.t88 7.49789
R1004 VSS.n360 VSS.t94 7.49789
R1005 VSS.n386 VSS.t84 7.49789
R1006 VSS.n339 VSS.t200 7.49789
R1007 VSS.n339 VSS.t210 7.49789
R1008 VSS.n164 VSS.t151 7.49789
R1009 VSS.n467 VSS.t153 7.12769
R1010 VSS.n438 VSS.t205 7.12769
R1011 VSS.n414 VSS.t1 7.12769
R1012 VSS.n475 VSS.t95 7.12769
R1013 VSS.n544 VSS.t203 7.12769
R1014 VSS.n518 VSS.t72 7.12769
R1015 VSS.n152 VSS.t103 7.12769
R1016 VSS.n224 VSS.t74 7.12769
R1017 VSS.n193 VSS.t109 7.12769
R1018 VSS.n509 VSS.n492 6.65737
R1019 VSS.n509 VSS.n493 6.65737
R1020 VSS.n503 VSS.t107 6.65737
R1021 VSS.n503 VSS.t98 6.65737
R1022 VSS.n403 VSS.n380 6.65737
R1023 VSS.n403 VSS.n381 6.65737
R1024 VSS.n392 VSS.t108 6.65737
R1025 VSS.n392 VSS.t86 6.65737
R1026 VSS.n182 VSS.n158 6.65737
R1027 VSS.n182 VSS.n159 6.65737
R1028 VSS.n171 VSS.t100 6.65737
R1029 VSS.n171 VSS.t152 6.65737
R1030 VSS.n561 VSS.n321 6.46636
R1031 VSS.n582 VSS.n581 6.45126
R1032 VSS.n891 VSS.n110 5.87352
R1033 VSS.n889 VSS.n888 5.8598
R1034 VSS.n1149 VSS.n1148 5.8598
R1035 VSS.n1152 VSS.n1151 5.8497
R1036 VSS.n859 VSS.n857 5.21612
R1037 VSS.n120 VSS.n118 5.21612
R1038 VSS.n125 VSS.t37 5.21612
R1039 VSS.n131 VSS.n129 5.21612
R1040 VSS.n137 VSS.t198 5.21612
R1041 VSS.n141 VSS.n139 5.21612
R1042 VSS.n260 VSS.t64 5.21612
R1043 VSS.n74 VSS.n72 5.21612
R1044 VSS.n80 VSS.n79 5.21612
R1045 VSS.n64 VSS.n62 5.21612
R1046 VSS.n70 VSS.n69 5.21612
R1047 VSS.n58 VSS.t244 5.21612
R1048 VSS.n60 VSS.t79 5.21612
R1049 VSS.n50 VSS.n48 5.21612
R1050 VSS.n56 VSS.n55 5.21612
R1051 VSS.n1116 VSS.t149 5.21612
R1052 VSS.n1118 VSS.t134 5.21612
R1053 VSS.n44 VSS.n43 5.21612
R1054 VSS.n37 VSS.t313 5.21612
R1055 VSS.n33 VSS.t295 5.21612
R1056 VSS.n29 VSS.t314 5.21612
R1057 VSS.n27 VSS.t293 5.21612
R1058 VSS.n240 VSS.n239 5.2005
R1059 VSS.n239 VSS.n238 5.2005
R1060 VSS.n243 VSS.n242 5.2005
R1061 VSS.n242 VSS.n241 5.2005
R1062 VSS.n355 VSS.n354 4.5005
R1063 VSS.n373 VSS.n359 4.5005
R1064 VSS.n469 VSS 4.5005
R1065 VSS.n151 VSS.n149 4.5005
R1066 VSS.n237 VSS.n236 4.5005
R1067 VSS.n236 VSS.n235 4.5005
R1068 VSS.n861 VSS.n860 4.4609
R1069 VSS.n859 VSS.n858 4.4609
R1070 VSS.n122 VSS.n121 4.4609
R1071 VSS.n120 VSS.n119 4.4609
R1072 VSS.n126 VSS.t57 4.4609
R1073 VSS.n125 VSS.t18 4.4609
R1074 VSS.n133 VSS.n132 4.4609
R1075 VSS.n131 VSS.n130 4.4609
R1076 VSS.n138 VSS.t159 4.4609
R1077 VSS.n137 VSS.t174 4.4609
R1078 VSS.n143 VSS.n142 4.4609
R1079 VSS.n141 VSS.n140 4.4609
R1080 VSS.n261 VSS.t68 4.4609
R1081 VSS.n260 VSS.t69 4.4609
R1082 VSS.n81 VSS.n77 4.4609
R1083 VSS.n80 VSS.n78 4.4609
R1084 VSS.n76 VSS.n75 4.4609
R1085 VSS.n74 VSS.n73 4.4609
R1086 VSS.n71 VSS.n67 4.4609
R1087 VSS.n70 VSS.n68 4.4609
R1088 VSS.n66 VSS.n65 4.4609
R1089 VSS.n64 VSS.n63 4.4609
R1090 VSS.n61 VSS.t245 4.4609
R1091 VSS.n60 VSS.t80 4.4609
R1092 VSS.n59 VSS.t243 4.4609
R1093 VSS.n58 VSS.t246 4.4609
R1094 VSS.n57 VSS.n53 4.4609
R1095 VSS.n56 VSS.n54 4.4609
R1096 VSS.n52 VSS.n51 4.4609
R1097 VSS.n50 VSS.n49 4.4609
R1098 VSS.n1119 VSS.t145 4.4609
R1099 VSS.n1118 VSS.t119 4.4609
R1100 VSS.n1117 VSS.t148 4.4609
R1101 VSS.n1116 VSS.t132 4.4609
R1102 VSS.n45 VSS.n41 4.4609
R1103 VSS.n44 VSS.n42 4.4609
R1104 VSS.n38 VSS.t287 4.4609
R1105 VSS.n37 VSS.t226 4.4609
R1106 VSS.n34 VSS.t315 4.4609
R1107 VSS.n33 VSS.t308 4.4609
R1108 VSS.n30 VSS.t300 4.4609
R1109 VSS.n29 VSS.t254 4.4609
R1110 VSS.n28 VSS.t320 4.4609
R1111 VSS.n27 VSS.t307 4.4609
R1112 VSS.n363 VSS.n362 4.45263
R1113 VSS.n340 VSS.n338 4.45095
R1114 VSS.n3 VSS.n2 4.29799
R1115 VSS.n1158 VSS.n1155 4.29732
R1116 VSS.n500 VSS.n496 4.27004
R1117 VSS.n505 VSS.n504 4.25879
R1118 VSS.n508 VSS.n507 4.25811
R1119 VSS.n864 VSS.n863 2.61255
R1120 VSS.n264 VSS.n263 2.61255
R1121 VSS.n85 VSS.n84 2.61255
R1122 VSS.n1122 VSS.n1121 2.61255
R1123 VSS.n389 VSS.n386 2.61175
R1124 VSS.n168 VSS.n164 2.61175
R1125 VSS.n551 VSS.n550 2.6005
R1126 VSS.n550 VSS.n549 2.6005
R1127 VSS.n548 VSS.n547 2.6005
R1128 VSS.n547 VSS.n546 2.6005
R1129 VSS.n545 VSS 2.6005
R1130 VSS.n545 VSS.n544 2.6005
R1131 VSS.n543 VSS.n541 2.6005
R1132 VSS.n543 VSS.n542 2.6005
R1133 VSS.n540 VSS.n539 2.6005
R1134 VSS.n539 VSS.n538 2.6005
R1135 VSS.n479 VSS.n478 2.6005
R1136 VSS.n478 VSS.n477 2.6005
R1137 VSS.n482 VSS.n481 2.6005
R1138 VSS.n481 VSS.n480 2.6005
R1139 VSS.n486 VSS.n485 2.6005
R1140 VSS.n485 VSS.n484 2.6005
R1141 VSS.n347 VSS.n346 2.6005
R1142 VSS.n346 VSS.n345 2.6005
R1143 VSS.n350 VSS.n349 2.6005
R1144 VSS.n349 VSS.n348 2.6005
R1145 VSS.n353 VSS.n352 2.6005
R1146 VSS.n352 VSS.n351 2.6005
R1147 VSS VSS.n501 2.6005
R1148 VSS.n506 VSS.n497 2.6005
R1149 VSS.n495 VSS.n494 2.6005
R1150 VSS.n499 VSS.n498 2.6005
R1151 VSS.n510 VSS.n491 2.6005
R1152 VSS.n491 VSS.n490 2.6005
R1153 VSS.n525 VSS.n524 2.6005
R1154 VSS.n524 VSS.n523 2.6005
R1155 VSS.n522 VSS.n521 2.6005
R1156 VSS.n521 VSS.n520 2.6005
R1157 VSS.n519 VSS 2.6005
R1158 VSS.n519 VSS.n518 2.6005
R1159 VSS.n517 VSS.n515 2.6005
R1160 VSS.n517 VSS.n516 2.6005
R1161 VSS.n514 VSS.n513 2.6005
R1162 VSS.n513 VSS.n512 2.6005
R1163 VSS.n528 VSS.n527 2.6005
R1164 VSS.n527 VSS.n526 2.6005
R1165 VSS.n466 VSS.n464 2.6005
R1166 VSS.n466 VSS.n465 2.6005
R1167 VSS.n422 VSS.n379 2.6005
R1168 VSS.n379 VSS.n378 2.6005
R1169 VSS.n421 VSS.n420 2.6005
R1170 VSS.n420 VSS.n419 2.6005
R1171 VSS.n418 VSS.n417 2.6005
R1172 VSS.n417 VSS.n416 2.6005
R1173 VSS.n415 VSS 2.6005
R1174 VSS.n415 VSS.n414 2.6005
R1175 VSS.n413 VSS.n411 2.6005
R1176 VSS.n413 VSS.n412 2.6005
R1177 VSS.n410 VSS.n409 2.6005
R1178 VSS.n409 VSS.n408 2.6005
R1179 VSS.n406 VSS.n405 2.6005
R1180 VSS.n405 VSS.n404 2.6005
R1181 VSS.n402 VSS.n383 2.6005
R1182 VSS.n383 VSS.n382 2.6005
R1183 VSS.n401 VSS.n400 2.6005
R1184 VSS.n400 VSS.n399 2.6005
R1185 VSS.n398 VSS.n396 2.6005
R1186 VSS.n398 VSS.n397 2.6005
R1187 VSS.n395 VSS.n394 2.6005
R1188 VSS.n394 VSS.n393 2.6005
R1189 VSS.n391 VSS.n385 2.6005
R1190 VSS.n385 VSS.n384 2.6005
R1191 VSS VSS.n390 2.6005
R1192 VSS.n390 VSS.t83 2.6005
R1193 VSS.n389 VSS.n388 2.6005
R1194 VSS.n442 VSS.n441 2.6005
R1195 VSS.n441 VSS.n440 2.6005
R1196 VSS.n439 VSS 2.6005
R1197 VSS.n439 VSS.n438 2.6005
R1198 VSS.n437 VSS.n435 2.6005
R1199 VSS.n437 VSS.n436 2.6005
R1200 VSS.n434 VSS.n433 2.6005
R1201 VSS.n433 VSS.n432 2.6005
R1202 VSS.n445 VSS.n444 2.6005
R1203 VSS.n444 VSS.n443 2.6005
R1204 VSS.n369 VSS.n368 2.6005
R1205 VSS.n368 VSS.n367 2.6005
R1206 VSS.n372 VSS.n371 2.6005
R1207 VSS.n371 VSS.n370 2.6005
R1208 VSS.n463 VSS.n462 2.6005
R1209 VSS.n462 VSS.n461 2.6005
R1210 VSS.n459 VSS.n458 2.6005
R1211 VSS.n458 VSS.n457 2.6005
R1212 VSS.n366 VSS.n365 2.6005
R1213 VSS.n365 VSS.n364 2.6005
R1214 VSS.n231 VSS.n230 2.6005
R1215 VSS.n230 VSS.n229 2.6005
R1216 VSS.n228 VSS.n227 2.6005
R1217 VSS.n227 VSS.n226 2.6005
R1218 VSS.n225 VSS 2.6005
R1219 VSS.n225 VSS.n224 2.6005
R1220 VSS.n223 VSS.n221 2.6005
R1221 VSS.n223 VSS.n222 2.6005
R1222 VSS.n220 VSS.n219 2.6005
R1223 VSS.n219 VSS.n218 2.6005
R1224 VSS.n201 VSS.n157 2.6005
R1225 VSS.n157 VSS.n156 2.6005
R1226 VSS.n200 VSS.n199 2.6005
R1227 VSS.n199 VSS.n198 2.6005
R1228 VSS.n197 VSS.n196 2.6005
R1229 VSS.n196 VSS.n195 2.6005
R1230 VSS.n194 VSS 2.6005
R1231 VSS.n194 VSS.n193 2.6005
R1232 VSS.n192 VSS.n190 2.6005
R1233 VSS.n192 VSS.n191 2.6005
R1234 VSS.n189 VSS.n188 2.6005
R1235 VSS.n188 VSS.n187 2.6005
R1236 VSS.n185 VSS.n184 2.6005
R1237 VSS.n184 VSS.n183 2.6005
R1238 VSS.n573 VSS.n572 2.6005
R1239 VSS.n572 VSS.n571 2.6005
R1240 VSS.n569 VSS.n568 2.6005
R1241 VSS.n568 VSS.n567 2.6005
R1242 VSS.n337 VSS.n336 2.6005
R1243 VSS.n336 VSS.n335 2.6005
R1244 VSS.n334 VSS.n333 2.6005
R1245 VSS.n333 VSS.n332 2.6005
R1246 VSS.n331 VSS.n330 2.6005
R1247 VSS.n330 VSS.n329 2.6005
R1248 VSS.n576 VSS.n575 2.6005
R1249 VSS.n575 VSS.n574 2.6005
R1250 VSS.n181 VSS.n161 2.6005
R1251 VSS.n161 VSS.n160 2.6005
R1252 VSS.n180 VSS.n179 2.6005
R1253 VSS.n179 VSS.n178 2.6005
R1254 VSS.n177 VSS.n175 2.6005
R1255 VSS.n177 VSS.n176 2.6005
R1256 VSS.n174 VSS.n173 2.6005
R1257 VSS.n173 VSS.n172 2.6005
R1258 VSS.n170 VSS.n163 2.6005
R1259 VSS.n163 VSS.n162 2.6005
R1260 VSS VSS.n169 2.6005
R1261 VSS.n169 VSS.t150 2.6005
R1262 VSS.n168 VSS.n167 2.6005
R1263 VSS.n855 VSS.n115 2.6005
R1264 VSS.n115 VSS.n114 2.6005
R1265 VSS.n830 VSS.n117 2.6005
R1266 VSS.n117 VSS.n116 2.6005
R1267 VSS.n828 VSS.n827 2.6005
R1268 VSS.n827 VSS.n826 2.6005
R1269 VSS.n825 VSS.n824 2.6005
R1270 VSS.n824 VSS.n823 2.6005
R1271 VSS.n822 VSS.n821 2.6005
R1272 VSS.n821 VSS.n820 2.6005
R1273 VSS.n819 VSS.n818 2.6005
R1274 VSS.n818 VSS.n817 2.6005
R1275 VSS.n816 VSS.n815 2.6005
R1276 VSS.n815 VSS.n814 2.6005
R1277 VSS.n813 VSS.n812 2.6005
R1278 VSS.n812 VSS.n811 2.6005
R1279 VSS.n810 VSS.n809 2.6005
R1280 VSS.n809 VSS.n808 2.6005
R1281 VSS.n807 VSS.n806 2.6005
R1282 VSS.n806 VSS.n805 2.6005
R1283 VSS.n804 VSS.n802 2.6005
R1284 VSS.n804 VSS.n803 2.6005
R1285 VSS.n801 VSS.n800 2.6005
R1286 VSS.n800 VSS.n799 2.6005
R1287 VSS.n798 VSS.n797 2.6005
R1288 VSS.n797 VSS.n796 2.6005
R1289 VSS.n795 VSS.n794 2.6005
R1290 VSS.n794 VSS.n793 2.6005
R1291 VSS.n792 VSS.n791 2.6005
R1292 VSS.n791 VSS.n790 2.6005
R1293 VSS.n789 VSS.n788 2.6005
R1294 VSS.n788 VSS.n787 2.6005
R1295 VSS.n786 VSS.n785 2.6005
R1296 VSS.n785 VSS.n784 2.6005
R1297 VSS.n783 VSS.n782 2.6005
R1298 VSS.n782 VSS.n781 2.6005
R1299 VSS.n780 VSS.n779 2.6005
R1300 VSS.n779 VSS.n778 2.6005
R1301 VSS.n777 VSS.n124 2.6005
R1302 VSS.n124 VSS.n123 2.6005
R1303 VSS.n776 VSS.n775 2.6005
R1304 VSS.n775 VSS.n774 2.6005
R1305 VSS.n773 VSS.n772 2.6005
R1306 VSS.n772 VSS.n771 2.6005
R1307 VSS.n770 VSS.n769 2.6005
R1308 VSS.n769 VSS.n768 2.6005
R1309 VSS.n767 VSS.n766 2.6005
R1310 VSS.n766 VSS.n765 2.6005
R1311 VSS.n764 VSS.n763 2.6005
R1312 VSS.n763 VSS.n762 2.6005
R1313 VSS.n761 VSS.n760 2.6005
R1314 VSS.n760 VSS.n759 2.6005
R1315 VSS.n758 VSS.n757 2.6005
R1316 VSS.n757 VSS.n756 2.6005
R1317 VSS.n755 VSS.n754 2.6005
R1318 VSS.n754 VSS.n753 2.6005
R1319 VSS.n752 VSS.n750 2.6005
R1320 VSS.n752 VSS.n751 2.6005
R1321 VSS.n749 VSS.n748 2.6005
R1322 VSS.n748 VSS.n747 2.6005
R1323 VSS.n746 VSS.n745 2.6005
R1324 VSS.n745 VSS.n744 2.6005
R1325 VSS.n743 VSS.n742 2.6005
R1326 VSS.n742 VSS.n741 2.6005
R1327 VSS.n740 VSS.n739 2.6005
R1328 VSS.n739 VSS.n738 2.6005
R1329 VSS.n737 VSS.n736 2.6005
R1330 VSS.n736 VSS.n735 2.6005
R1331 VSS.n734 VSS.n733 2.6005
R1332 VSS.n733 VSS.n732 2.6005
R1333 VSS.n731 VSS.n730 2.6005
R1334 VSS.n730 VSS.n729 2.6005
R1335 VSS.n727 VSS.n726 2.6005
R1336 VSS.n726 VSS.n725 2.6005
R1337 VSS.n724 VSS.n128 2.6005
R1338 VSS.n128 VSS.n127 2.6005
R1339 VSS.n722 VSS.n721 2.6005
R1340 VSS.n721 VSS.n720 2.6005
R1341 VSS.n719 VSS.n718 2.6005
R1342 VSS.n718 VSS.n717 2.6005
R1343 VSS.n716 VSS.n715 2.6005
R1344 VSS.n715 VSS.n714 2.6005
R1345 VSS.n713 VSS.n712 2.6005
R1346 VSS.n712 VSS.n711 2.6005
R1347 VSS.n710 VSS.n709 2.6005
R1348 VSS.n709 VSS.n708 2.6005
R1349 VSS.n707 VSS.n706 2.6005
R1350 VSS.n706 VSS.n705 2.6005
R1351 VSS.n704 VSS.n703 2.6005
R1352 VSS.n703 VSS.n702 2.6005
R1353 VSS.n701 VSS.n700 2.6005
R1354 VSS.n700 VSS.n699 2.6005
R1355 VSS.n698 VSS.n696 2.6005
R1356 VSS.n698 VSS.n697 2.6005
R1357 VSS.n695 VSS.n694 2.6005
R1358 VSS.n694 VSS.n693 2.6005
R1359 VSS.n692 VSS.n691 2.6005
R1360 VSS.n691 VSS.n690 2.6005
R1361 VSS.n689 VSS.n688 2.6005
R1362 VSS.n688 VSS.n687 2.6005
R1363 VSS.n686 VSS.n685 2.6005
R1364 VSS.n685 VSS.n684 2.6005
R1365 VSS.n683 VSS.n682 2.6005
R1366 VSS.n682 VSS.n681 2.6005
R1367 VSS.n680 VSS.n679 2.6005
R1368 VSS.n679 VSS.n678 2.6005
R1369 VSS.n677 VSS.n676 2.6005
R1370 VSS.n676 VSS.n675 2.6005
R1371 VSS.n674 VSS.n673 2.6005
R1372 VSS.n673 VSS.n672 2.6005
R1373 VSS.n671 VSS.n135 2.6005
R1374 VSS.n135 VSS.n134 2.6005
R1375 VSS.n854 VSS.n853 2.6005
R1376 VSS.n853 VSS.n852 2.6005
R1377 VSS.n851 VSS.n850 2.6005
R1378 VSS.n850 VSS.n849 2.6005
R1379 VSS.n848 VSS.n847 2.6005
R1380 VSS.n847 VSS.n846 2.6005
R1381 VSS.n845 VSS.n844 2.6005
R1382 VSS.n844 VSS.n843 2.6005
R1383 VSS.n842 VSS.n841 2.6005
R1384 VSS.n841 VSS.n840 2.6005
R1385 VSS.n839 VSS.n838 2.6005
R1386 VSS.n838 VSS.n837 2.6005
R1387 VSS.n836 VSS.n835 2.6005
R1388 VSS.n835 VSS.n834 2.6005
R1389 VSS.n833 VSS.n832 2.6005
R1390 VSS.n832 VSS.n831 2.6005
R1391 VSS.n863 VSS.n862 2.6005
R1392 VSS.n867 VSS.n866 2.6005
R1393 VSS.n866 VSS.n865 2.6005
R1394 VSS.n870 VSS.n869 2.6005
R1395 VSS.n869 VSS.n868 2.6005
R1396 VSS.n873 VSS.n872 2.6005
R1397 VSS.n872 VSS.n871 2.6005
R1398 VSS.n876 VSS.n875 2.6005
R1399 VSS.n875 VSS.n874 2.6005
R1400 VSS.n879 VSS.n878 2.6005
R1401 VSS.n878 VSS.n877 2.6005
R1402 VSS.n882 VSS.n881 2.6005
R1403 VSS.n881 VSS.n880 2.6005
R1404 VSS.n885 VSS.n884 2.6005
R1405 VSS.n884 VSS.n883 2.6005
R1406 VSS.n585 VSS.n145 2.6005
R1407 VSS.n145 VSS.n144 2.6005
R1408 VSS.n612 VSS.n611 2.6005
R1409 VSS.n611 VSS.n610 2.6005
R1410 VSS.n609 VSS.n608 2.6005
R1411 VSS.n608 VSS.n607 2.6005
R1412 VSS.n606 VSS.n605 2.6005
R1413 VSS.n605 VSS.n604 2.6005
R1414 VSS.n603 VSS.n602 2.6005
R1415 VSS.n602 VSS.n601 2.6005
R1416 VSS.n600 VSS.n599 2.6005
R1417 VSS.n599 VSS.n598 2.6005
R1418 VSS.n597 VSS.n596 2.6005
R1419 VSS.n596 VSS.n595 2.6005
R1420 VSS.n594 VSS.n593 2.6005
R1421 VSS.n593 VSS.n592 2.6005
R1422 VSS.n591 VSS.n590 2.6005
R1423 VSS.n590 VSS.n589 2.6005
R1424 VSS.n588 VSS.n586 2.6005
R1425 VSS.n588 VSS.n587 2.6005
R1426 VSS.n313 VSS.n259 2.6005
R1427 VSS.n259 VSS.n258 2.6005
R1428 VSS.n312 VSS.n311 2.6005
R1429 VSS.n311 VSS.n310 2.6005
R1430 VSS.n309 VSS.n308 2.6005
R1431 VSS.n308 VSS.n307 2.6005
R1432 VSS.n306 VSS.n305 2.6005
R1433 VSS.n305 VSS.n304 2.6005
R1434 VSS.n303 VSS.n302 2.6005
R1435 VSS.n302 VSS.n301 2.6005
R1436 VSS.n300 VSS.n299 2.6005
R1437 VSS.n299 VSS.n298 2.6005
R1438 VSS.n297 VSS.n296 2.6005
R1439 VSS.n296 VSS.n295 2.6005
R1440 VSS.n294 VSS.n293 2.6005
R1441 VSS.n293 VSS.n292 2.6005
R1442 VSS.n291 VSS.n290 2.6005
R1443 VSS.n290 VSS.n289 2.6005
R1444 VSS.n288 VSS.n286 2.6005
R1445 VSS.n288 VSS.n287 2.6005
R1446 VSS.n285 VSS.n284 2.6005
R1447 VSS.n284 VSS.n283 2.6005
R1448 VSS.n282 VSS.n281 2.6005
R1449 VSS.n281 VSS.n280 2.6005
R1450 VSS.n279 VSS.n278 2.6005
R1451 VSS.n278 VSS.n277 2.6005
R1452 VSS.n276 VSS.n275 2.6005
R1453 VSS.n275 VSS.n274 2.6005
R1454 VSS.n273 VSS.n272 2.6005
R1455 VSS.n272 VSS.n271 2.6005
R1456 VSS.n270 VSS.n269 2.6005
R1457 VSS.n269 VSS.n268 2.6005
R1458 VSS.n267 VSS.n266 2.6005
R1459 VSS.n266 VSS.n265 2.6005
R1460 VSS.n263 VSS.n262 2.6005
R1461 VSS.n246 VSS.n245 2.6005
R1462 VSS.n245 VSS.n244 2.6005
R1463 VSS.n249 VSS.n248 2.6005
R1464 VSS.n248 VSS.n247 2.6005
R1465 VSS.n252 VSS.n251 2.6005
R1466 VSS.n251 VSS.n250 2.6005
R1467 VSS.n255 VSS.n254 2.6005
R1468 VSS.n254 VSS.n253 2.6005
R1469 VSS.n316 VSS.n315 2.6005
R1470 VSS.n315 VSS.n314 2.6005
R1471 VSS.n617 VSS.n616 2.6005
R1472 VSS.n616 VSS.n615 2.6005
R1473 VSS.n639 VSS.n638 2.6005
R1474 VSS.n638 VSS.n637 2.6005
R1475 VSS.n636 VSS.n635 2.6005
R1476 VSS.n635 VSS.n634 2.6005
R1477 VSS.n633 VSS.n632 2.6005
R1478 VSS.n632 VSS.n631 2.6005
R1479 VSS.n630 VSS.n629 2.6005
R1480 VSS.n629 VSS.n628 2.6005
R1481 VSS.n627 VSS.n626 2.6005
R1482 VSS.n626 VSS.n625 2.6005
R1483 VSS.n624 VSS.n623 2.6005
R1484 VSS.n623 VSS.n622 2.6005
R1485 VSS.n620 VSS.n619 2.6005
R1486 VSS.n619 VSS.n618 2.6005
R1487 VSS.n670 VSS.n669 2.6005
R1488 VSS.n669 VSS.n668 2.6005
R1489 VSS.n667 VSS.n666 2.6005
R1490 VSS.n666 VSS.n665 2.6005
R1491 VSS.n664 VSS.n663 2.6005
R1492 VSS.n663 VSS.n662 2.6005
R1493 VSS.n661 VSS.n660 2.6005
R1494 VSS.n660 VSS.n659 2.6005
R1495 VSS.n658 VSS.n657 2.6005
R1496 VSS.n657 VSS.n656 2.6005
R1497 VSS.n655 VSS.n654 2.6005
R1498 VSS.n654 VSS.n653 2.6005
R1499 VSS.n652 VSS.n651 2.6005
R1500 VSS.n651 VSS.n650 2.6005
R1501 VSS.n649 VSS.n648 2.6005
R1502 VSS.n648 VSS.n647 2.6005
R1503 VSS.n642 VSS.n641 2.6005
R1504 VSS.n641 VSS.n640 2.6005
R1505 VSS.n1113 VSS.n1111 2.6005
R1506 VSS.n1113 VSS.n1112 2.6005
R1507 VSS.n1092 VSS.n1091 2.6005
R1508 VSS.n1091 VSS.n1090 2.6005
R1509 VSS.n1095 VSS.n1094 2.6005
R1510 VSS.n1094 VSS.n1093 2.6005
R1511 VSS.n1098 VSS.n1097 2.6005
R1512 VSS.n1097 VSS.n1096 2.6005
R1513 VSS.n1101 VSS.n1100 2.6005
R1514 VSS.n1100 VSS.n1099 2.6005
R1515 VSS.n1104 VSS.n1103 2.6005
R1516 VSS.n1103 VSS.n1102 2.6005
R1517 VSS.n1107 VSS.n1106 2.6005
R1518 VSS.n1106 VSS.n1105 2.6005
R1519 VSS.n1110 VSS.n1109 2.6005
R1520 VSS.n1109 VSS.n1108 2.6005
R1521 VSS.n1143 VSS.n1142 2.6005
R1522 VSS.n1142 VSS.n1141 2.6005
R1523 VSS.n1140 VSS.n1139 2.6005
R1524 VSS.n1139 VSS.n1138 2.6005
R1525 VSS.n1137 VSS.n1136 2.6005
R1526 VSS.n1136 VSS.n1135 2.6005
R1527 VSS.n1134 VSS.n1133 2.6005
R1528 VSS.n1133 VSS.n1132 2.6005
R1529 VSS.n1131 VSS.n1130 2.6005
R1530 VSS.n1130 VSS.n1129 2.6005
R1531 VSS.n1128 VSS.n1127 2.6005
R1532 VSS.n1127 VSS.n1126 2.6005
R1533 VSS.n1125 VSS.n1124 2.6005
R1534 VSS.n1124 VSS.n1123 2.6005
R1535 VSS.n1121 VSS.n1120 2.6005
R1536 VSS.n1089 VSS.n1088 2.6005
R1537 VSS.n1088 VSS.n1087 2.6005
R1538 VSS.n1086 VSS.n1085 2.6005
R1539 VSS.n1085 VSS.n1084 2.6005
R1540 VSS.n1038 VSS.n1037 2.6005
R1541 VSS.n1037 VSS.n1036 2.6005
R1542 VSS.n1041 VSS.n1040 2.6005
R1543 VSS.n1040 VSS.n1039 2.6005
R1544 VSS.n1044 VSS.n1043 2.6005
R1545 VSS.n1043 VSS.n1042 2.6005
R1546 VSS.n1047 VSS.n1046 2.6005
R1547 VSS.n1046 VSS.n1045 2.6005
R1548 VSS.n1050 VSS.n1049 2.6005
R1549 VSS.n1049 VSS.n1048 2.6005
R1550 VSS.n1053 VSS.n1052 2.6005
R1551 VSS.n1052 VSS.n1051 2.6005
R1552 VSS.n1056 VSS.n1055 2.6005
R1553 VSS.n1055 VSS.n1054 2.6005
R1554 VSS.n1059 VSS.n1057 2.6005
R1555 VSS.n1059 VSS.n1058 2.6005
R1556 VSS.n1062 VSS.n1061 2.6005
R1557 VSS.n1061 VSS.n1060 2.6005
R1558 VSS.n1065 VSS.n1064 2.6005
R1559 VSS.n1064 VSS.n1063 2.6005
R1560 VSS.n1068 VSS.n1067 2.6005
R1561 VSS.n1067 VSS.n1066 2.6005
R1562 VSS.n1071 VSS.n1070 2.6005
R1563 VSS.n1070 VSS.n1069 2.6005
R1564 VSS.n1074 VSS.n1073 2.6005
R1565 VSS.n1073 VSS.n1072 2.6005
R1566 VSS.n1077 VSS.n1076 2.6005
R1567 VSS.n1076 VSS.n1075 2.6005
R1568 VSS.n1080 VSS.n1079 2.6005
R1569 VSS.n1079 VSS.n1078 2.6005
R1570 VSS.n1083 VSS.n1082 2.6005
R1571 VSS.n1082 VSS.n1081 2.6005
R1572 VSS.n1034 VSS.n1033 2.6005
R1573 VSS.n1033 VSS.n1032 2.6005
R1574 VSS.n1031 VSS.n1030 2.6005
R1575 VSS.n1030 VSS.n1029 2.6005
R1576 VSS.n982 VSS.n981 2.6005
R1577 VSS.n981 VSS.n980 2.6005
R1578 VSS.n985 VSS.n984 2.6005
R1579 VSS.n984 VSS.n983 2.6005
R1580 VSS.n988 VSS.n987 2.6005
R1581 VSS.n987 VSS.n986 2.6005
R1582 VSS.n991 VSS.n990 2.6005
R1583 VSS.n990 VSS.n989 2.6005
R1584 VSS.n994 VSS.n993 2.6005
R1585 VSS.n993 VSS.n992 2.6005
R1586 VSS.n997 VSS.n996 2.6005
R1587 VSS.n996 VSS.n995 2.6005
R1588 VSS.n1000 VSS.n999 2.6005
R1589 VSS.n999 VSS.n998 2.6005
R1590 VSS.n1003 VSS.n1001 2.6005
R1591 VSS.n1003 VSS.n1002 2.6005
R1592 VSS.n1006 VSS.n1005 2.6005
R1593 VSS.n1005 VSS.n1004 2.6005
R1594 VSS.n1009 VSS.n1008 2.6005
R1595 VSS.n1008 VSS.n1007 2.6005
R1596 VSS.n1012 VSS.n1011 2.6005
R1597 VSS.n1011 VSS.n1010 2.6005
R1598 VSS.n1015 VSS.n1014 2.6005
R1599 VSS.n1014 VSS.n1013 2.6005
R1600 VSS.n1018 VSS.n1017 2.6005
R1601 VSS.n1017 VSS.n1016 2.6005
R1602 VSS.n1021 VSS.n1020 2.6005
R1603 VSS.n1020 VSS.n1019 2.6005
R1604 VSS.n1024 VSS.n1023 2.6005
R1605 VSS.n1023 VSS.n1022 2.6005
R1606 VSS.n1027 VSS.n1026 2.6005
R1607 VSS.n1026 VSS.n1025 2.6005
R1608 VSS.n979 VSS.n978 2.6005
R1609 VSS.n978 VSS.n977 2.6005
R1610 VSS.n976 VSS.n975 2.6005
R1611 VSS.n975 VSS.n974 2.6005
R1612 VSS.n928 VSS.n927 2.6005
R1613 VSS.n927 VSS.n926 2.6005
R1614 VSS.n931 VSS.n930 2.6005
R1615 VSS.n930 VSS.n929 2.6005
R1616 VSS.n934 VSS.n933 2.6005
R1617 VSS.n933 VSS.n932 2.6005
R1618 VSS.n937 VSS.n936 2.6005
R1619 VSS.n936 VSS.n935 2.6005
R1620 VSS.n940 VSS.n939 2.6005
R1621 VSS.n939 VSS.n938 2.6005
R1622 VSS.n943 VSS.n942 2.6005
R1623 VSS.n942 VSS.n941 2.6005
R1624 VSS.n946 VSS.n945 2.6005
R1625 VSS.n945 VSS.n944 2.6005
R1626 VSS.n949 VSS.n947 2.6005
R1627 VSS.n949 VSS.n948 2.6005
R1628 VSS.n952 VSS.n951 2.6005
R1629 VSS.n951 VSS.n950 2.6005
R1630 VSS.n955 VSS.n954 2.6005
R1631 VSS.n954 VSS.n953 2.6005
R1632 VSS.n958 VSS.n957 2.6005
R1633 VSS.n957 VSS.n956 2.6005
R1634 VSS.n961 VSS.n960 2.6005
R1635 VSS.n960 VSS.n959 2.6005
R1636 VSS.n964 VSS.n963 2.6005
R1637 VSS.n963 VSS.n962 2.6005
R1638 VSS.n967 VSS.n966 2.6005
R1639 VSS.n966 VSS.n965 2.6005
R1640 VSS.n970 VSS.n969 2.6005
R1641 VSS.n969 VSS.n968 2.6005
R1642 VSS.n973 VSS.n972 2.6005
R1643 VSS.n972 VSS.n971 2.6005
R1644 VSS.n924 VSS.n923 2.6005
R1645 VSS.n923 VSS.n922 2.6005
R1646 VSS.n900 VSS.n899 2.6005
R1647 VSS.n899 VSS.n898 2.6005
R1648 VSS.n903 VSS.n902 2.6005
R1649 VSS.n902 VSS.n901 2.6005
R1650 VSS.n906 VSS.n905 2.6005
R1651 VSS.n905 VSS.n904 2.6005
R1652 VSS.n909 VSS.n908 2.6005
R1653 VSS.n908 VSS.n907 2.6005
R1654 VSS.n912 VSS.n911 2.6005
R1655 VSS.n911 VSS.n910 2.6005
R1656 VSS.n915 VSS.n914 2.6005
R1657 VSS.n914 VSS.n913 2.6005
R1658 VSS.n918 VSS.n917 2.6005
R1659 VSS.n917 VSS.n916 2.6005
R1660 VSS.n921 VSS.n920 2.6005
R1661 VSS.n920 VSS.n919 2.6005
R1662 VSS.n84 VSS.n83 2.6005
R1663 VSS.n88 VSS.n87 2.6005
R1664 VSS.n87 VSS.n86 2.6005
R1665 VSS.n91 VSS.n90 2.6005
R1666 VSS.n90 VSS.n89 2.6005
R1667 VSS.n94 VSS.n93 2.6005
R1668 VSS.n93 VSS.n92 2.6005
R1669 VSS.n97 VSS.n96 2.6005
R1670 VSS.n96 VSS.n95 2.6005
R1671 VSS.n100 VSS.n99 2.6005
R1672 VSS.n99 VSS.n98 2.6005
R1673 VSS.n103 VSS.n102 2.6005
R1674 VSS.n102 VSS.n101 2.6005
R1675 VSS.n106 VSS.n105 2.6005
R1676 VSS.n105 VSS.n104 2.6005
R1677 VSS.n897 VSS.n896 2.6005
R1678 VSS.n896 VSS.n895 2.6005
R1679 VSS.n1182 VSS.n47 2.6005
R1680 VSS.n47 VSS.n46 2.6005
R1681 VSS.n1185 VSS.n1184 2.6005
R1682 VSS.n1184 VSS.n1183 2.6005
R1683 VSS.n1188 VSS.n1187 2.6005
R1684 VSS.n1187 VSS.n1186 2.6005
R1685 VSS.n1191 VSS.n1190 2.6005
R1686 VSS.n1190 VSS.n1189 2.6005
R1687 VSS.n1194 VSS.n1193 2.6005
R1688 VSS.n1193 VSS.n1192 2.6005
R1689 VSS.n1197 VSS.n1196 2.6005
R1690 VSS.n1196 VSS.n1195 2.6005
R1691 VSS.n1200 VSS.n1199 2.6005
R1692 VSS.n1199 VSS.n1198 2.6005
R1693 VSS.n1203 VSS.n1202 2.6005
R1694 VSS.n1202 VSS.n1201 2.6005
R1695 VSS.n1207 VSS.n1206 2.6005
R1696 VSS.n1206 VSS.n1205 2.6005
R1697 VSS.n1208 VSS.n40 2.6005
R1698 VSS.n40 VSS.n39 2.6005
R1699 VSS.n1257 VSS.n1256 2.6005
R1700 VSS.n1256 VSS.n1255 2.6005
R1701 VSS.n1254 VSS.n1253 2.6005
R1702 VSS.n1253 VSS.n1252 2.6005
R1703 VSS.n1251 VSS.n1250 2.6005
R1704 VSS.n1250 VSS.n1249 2.6005
R1705 VSS.n1248 VSS.n1247 2.6005
R1706 VSS.n1247 VSS.n1246 2.6005
R1707 VSS.n1245 VSS.n1244 2.6005
R1708 VSS.n1244 VSS.n1243 2.6005
R1709 VSS.n1242 VSS.n1241 2.6005
R1710 VSS.n1241 VSS.n1240 2.6005
R1711 VSS.n1239 VSS.n1238 2.6005
R1712 VSS.n1238 VSS.n1237 2.6005
R1713 VSS.n1236 VSS.n1235 2.6005
R1714 VSS.n1235 VSS.n1234 2.6005
R1715 VSS.n1233 VSS.n1231 2.6005
R1716 VSS.n1233 VSS.n1232 2.6005
R1717 VSS.n1230 VSS.n1229 2.6005
R1718 VSS.n1229 VSS.n1228 2.6005
R1719 VSS.n1227 VSS.n1226 2.6005
R1720 VSS.n1226 VSS.n1225 2.6005
R1721 VSS.n1224 VSS.n1223 2.6005
R1722 VSS.n1223 VSS.n1222 2.6005
R1723 VSS.n1221 VSS.n1220 2.6005
R1724 VSS.n1220 VSS.n1219 2.6005
R1725 VSS.n1218 VSS.n1217 2.6005
R1726 VSS.n1217 VSS.n1216 2.6005
R1727 VSS.n1215 VSS.n1214 2.6005
R1728 VSS.n1214 VSS.n1213 2.6005
R1729 VSS.n1212 VSS.n1211 2.6005
R1730 VSS.n1211 VSS.n1210 2.6005
R1731 VSS.n1260 VSS.n1259 2.6005
R1732 VSS.n1259 VSS.n1258 2.6005
R1733 VSS.n1261 VSS.n36 2.6005
R1734 VSS.n36 VSS.n35 2.6005
R1735 VSS.n1310 VSS.n1309 2.6005
R1736 VSS.n1309 VSS.n1308 2.6005
R1737 VSS.n1307 VSS.n1306 2.6005
R1738 VSS.n1306 VSS.n1305 2.6005
R1739 VSS.n1304 VSS.n1303 2.6005
R1740 VSS.n1303 VSS.n1302 2.6005
R1741 VSS.n1301 VSS.n1300 2.6005
R1742 VSS.n1300 VSS.n1299 2.6005
R1743 VSS.n1298 VSS.n1297 2.6005
R1744 VSS.n1297 VSS.n1296 2.6005
R1745 VSS.n1295 VSS.n1294 2.6005
R1746 VSS.n1294 VSS.n1293 2.6005
R1747 VSS.n1292 VSS.n1291 2.6005
R1748 VSS.n1291 VSS.n1290 2.6005
R1749 VSS.n1289 VSS.n1288 2.6005
R1750 VSS.n1288 VSS.n1287 2.6005
R1751 VSS.n1286 VSS.n1284 2.6005
R1752 VSS.n1286 VSS.n1285 2.6005
R1753 VSS.n1283 VSS.n1282 2.6005
R1754 VSS.n1282 VSS.n1281 2.6005
R1755 VSS.n1280 VSS.n1279 2.6005
R1756 VSS.n1279 VSS.n1278 2.6005
R1757 VSS.n1277 VSS.n1276 2.6005
R1758 VSS.n1276 VSS.n1275 2.6005
R1759 VSS.n1274 VSS.n1273 2.6005
R1760 VSS.n1273 VSS.n1272 2.6005
R1761 VSS.n1271 VSS.n1270 2.6005
R1762 VSS.n1270 VSS.n1269 2.6005
R1763 VSS.n1268 VSS.n1267 2.6005
R1764 VSS.n1267 VSS.n1266 2.6005
R1765 VSS.n1265 VSS.n1264 2.6005
R1766 VSS.n1264 VSS.n1263 2.6005
R1767 VSS.n1313 VSS.n1312 2.6005
R1768 VSS.n1312 VSS.n1311 2.6005
R1769 VSS.n1314 VSS.n32 2.6005
R1770 VSS.n32 VSS.n31 2.6005
R1771 VSS.n1363 VSS.n1362 2.6005
R1772 VSS.n1362 VSS.n1361 2.6005
R1773 VSS.n1360 VSS.n1359 2.6005
R1774 VSS.n1359 VSS.n1358 2.6005
R1775 VSS.n1357 VSS.n1356 2.6005
R1776 VSS.n1356 VSS.n1355 2.6005
R1777 VSS.n1354 VSS.n1353 2.6005
R1778 VSS.n1353 VSS.n1352 2.6005
R1779 VSS.n1351 VSS.n1350 2.6005
R1780 VSS.n1350 VSS.n1349 2.6005
R1781 VSS.n1348 VSS.n1347 2.6005
R1782 VSS.n1347 VSS.n1346 2.6005
R1783 VSS.n1345 VSS.n1344 2.6005
R1784 VSS.n1344 VSS.n1343 2.6005
R1785 VSS.n1342 VSS.n1341 2.6005
R1786 VSS.n1341 VSS.n1340 2.6005
R1787 VSS.n1339 VSS.n1337 2.6005
R1788 VSS.n1339 VSS.n1338 2.6005
R1789 VSS.n1336 VSS.n1335 2.6005
R1790 VSS.n1335 VSS.n1334 2.6005
R1791 VSS.n1333 VSS.n1332 2.6005
R1792 VSS.n1332 VSS.n1331 2.6005
R1793 VSS.n1330 VSS.n1329 2.6005
R1794 VSS.n1329 VSS.n1328 2.6005
R1795 VSS.n1327 VSS.n1326 2.6005
R1796 VSS.n1326 VSS.n1325 2.6005
R1797 VSS.n1324 VSS.n1323 2.6005
R1798 VSS.n1323 VSS.n1322 2.6005
R1799 VSS.n1321 VSS.n1320 2.6005
R1800 VSS.n1320 VSS.n1319 2.6005
R1801 VSS.n1318 VSS.n1317 2.6005
R1802 VSS.n1317 VSS.n1316 2.6005
R1803 VSS.n1366 VSS.n1365 2.6005
R1804 VSS.n1365 VSS.n1364 2.6005
R1805 VSS.n1391 VSS.n1390 2.6005
R1806 VSS.n1390 VSS.n1389 2.6005
R1807 VSS.n1388 VSS.n1387 2.6005
R1808 VSS.n1387 VSS.n1386 2.6005
R1809 VSS.n1385 VSS.n1384 2.6005
R1810 VSS.n1384 VSS.n1383 2.6005
R1811 VSS.n1382 VSS.n1381 2.6005
R1812 VSS.n1381 VSS.n1380 2.6005
R1813 VSS.n1379 VSS.n1378 2.6005
R1814 VSS.n1378 VSS.n1377 2.6005
R1815 VSS.n1376 VSS.n1375 2.6005
R1816 VSS.n1375 VSS.n1374 2.6005
R1817 VSS.n1373 VSS.n1372 2.6005
R1818 VSS.n1372 VSS.n1371 2.6005
R1819 VSS.n1369 VSS.n1368 2.6005
R1820 VSS.n1368 VSS.n1367 2.6005
R1821 VSS.n1 VSS.n0 2.6005
R1822 VSS.n6 VSS.n5 2.6005
R1823 VSS.n5 VSS.n4 2.6005
R1824 VSS.n9 VSS.n8 2.6005
R1825 VSS.n8 VSS.n7 2.6005
R1826 VSS.n12 VSS.n11 2.6005
R1827 VSS.n11 VSS.n10 2.6005
R1828 VSS.n15 VSS.n14 2.6005
R1829 VSS.n14 VSS.n13 2.6005
R1830 VSS.n18 VSS.n17 2.6005
R1831 VSS.n17 VSS.n16 2.6005
R1832 VSS.n21 VSS.n20 2.6005
R1833 VSS.n20 VSS.n19 2.6005
R1834 VSS.n1394 VSS.n1393 2.6005
R1835 VSS.n1393 VSS.n1392 2.6005
R1836 VSS.n1176 VSS.n1175 2.6005
R1837 VSS.n1175 VSS.n1174 2.6005
R1838 VSS.n1173 VSS.n1172 2.6005
R1839 VSS.n1172 VSS.n1171 2.6005
R1840 VSS.n1170 VSS.n1169 2.6005
R1841 VSS.n1169 VSS.n1168 2.6005
R1842 VSS.n1167 VSS.n1166 2.6005
R1843 VSS.n1166 VSS.n1165 2.6005
R1844 VSS.n1164 VSS.n1163 2.6005
R1845 VSS.n1163 VSS.n1162 2.6005
R1846 VSS.n1161 VSS.n1160 2.6005
R1847 VSS.n1160 VSS.n1159 2.6005
R1848 VSS.n1157 VSS.n1156 2.6005
R1849 VSS.n530 VSS.n489 2.41287
R1850 VSS.n489 VSS.n488 2.41287
R1851 VSS.n476 VSS 2.41287
R1852 VSS.n476 VSS.n475 2.41287
R1853 VSS.n555 VSS.n554 2.41287
R1854 VSS.n554 VSS.n553 2.41287
R1855 VSS.n455 VSS.n448 2.41287
R1856 VSS.n448 VSS.n447 2.41287
R1857 VSS.n429 VSS.n377 2.41287
R1858 VSS.n377 VSS.n376 2.41287
R1859 VSS VSS.n468 2.41287
R1860 VSS.n468 VSS.n467 2.41287
R1861 VSS VSS.n153 2.41287
R1862 VSS.n153 VSS.n152 2.41287
R1863 VSS.n233 VSS.n155 2.41287
R1864 VSS.n155 VSS.n154 2.41287
R1865 VSS.n205 VSS.n204 2.41287
R1866 VSS.n204 VSS.n203 2.41287
R1867 VSS.n318 VSS.n257 2.41287
R1868 VSS.n257 VSS.n256 2.41287
R1869 VSS.n113 VSS.n111 2.41287
R1870 VSS.n113 VSS.n112 2.41287
R1871 VSS.n894 VSS.n892 2.41287
R1872 VSS.n894 VSS.n893 2.41287
R1873 VSS.n1145 VSS.n1115 2.41287
R1874 VSS.n646 VSS.n644 2.41287
R1875 VSS.n646 VSS.n645 2.41287
R1876 VSS.n1115 VSS.n1114 2.41287
R1877 VSS.n25 VSS.n24 2.41287
R1878 VSS.n24 VSS.n23 2.41287
R1879 VSS.n1180 VSS.n1179 2.41287
R1880 VSS.n1179 VSS.n1178 2.41287
R1881 VSS.n888 VSS.n111 2.2512
R1882 VSS.n583 VSS.n582 2.24619
R1883 VSS.n887 VSS.n886 2.24619
R1884 VSS.n887 VSS.n856 2.24599
R1885 VSS.n109 VSS.n26 2.24599
R1886 VSS.n474 VSS.n473 2.24559
R1887 VSS VSS.n342 2.2449
R1888 VSS.n340 VSS 2.24431
R1889 VSS.n357 VSS.n356 2.24421
R1890 VSS.n362 VSS 2.24347
R1891 VSS.n865 VSS.t268 2.11914
R1892 VSS.n834 VSS.t258 2.11914
R1893 VSS.n826 VSS.t166 2.11914
R1894 VSS.n781 VSS.t160 2.11914
R1895 VSS.n774 VSS.t24 2.11914
R1896 VSS.n729 VSS.t17 2.11914
R1897 VSS.n720 VSS.t21 2.11914
R1898 VSS.n675 VSS.t26 2.11914
R1899 VSS.n668 VSS.t170 2.11914
R1900 VSS.n622 VSS.t158 2.11914
R1901 VSS.n610 VSS.t183 2.11914
R1902 VSS.n256 VSS.t191 2.11914
R1903 VSS.n310 VSS.t8 2.11914
R1904 VSS.n265 VSS.t63 2.11914
R1905 VSS.n501 VSS.n496 1.65822
R1906 VSS.n505 VSS.n499 1.65822
R1907 VSS.n3 VSS.n1 1.64953
R1908 VSS.n1158 VSS.n1157 1.64943
R1909 VSS.n0 VSS.t267 1.64109
R1910 VSS.n1371 VSS.t292 1.64109
R1911 VSS.n1361 VSS.t296 1.64109
R1912 VSS.n1316 VSS.t253 1.64109
R1913 VSS.n1308 VSS.t237 1.64109
R1914 VSS.n1263 VSS.t294 1.64109
R1915 VSS.n1255 VSS.t262 1.64109
R1916 VSS.n1210 VSS.t225 1.64109
R1917 VSS.n1201 VSS.t233 1.64109
R1918 VSS.n1156 VSS.t271 1.64109
R1919 VSS.n535 VSS.n534 1.5005
R1920 VSS.n557 VSS.n556 1.5005
R1921 VSS.n565 VSS.n564 1.5005
R1922 VSS.n215 VSS.n214 1.5005
R1923 VSS.n320 VSS.n319 1.49906
R1924 VSS.n892 VSS.n891 1.49673
R1925 VSS.n1150 VSS.n1146 1.49673
R1926 VSS.n558 VSS.n557 1.49619
R1927 VSS.n564 VSS.n561 1.49619
R1928 VSS.n579 VSS.n578 1.49619
R1929 VSS.n473 VSS.n472 1.35924
R1930 VSS.n452 VSS.n451 1.34792
R1931 VSS.n559 VSS.n558 1.34613
R1932 VSS.n579 VSS.n148 1.34613
R1933 VSS.n209 VSS.n208 1.33121
R1934 VSS.n429 VSS.n428 1.1255
R1935 VSS.n455 VSS.n454 1.1255
R1936 VSS VSS.n474 1.1255
R1937 VSS.n578 VSS 1.1255
R1938 VSS.n454 VSS.n452 1.12386
R1939 VSS.n1177 VSS.n1153 1.12363
R1940 VSS.n428 VSS.n426 1.12348
R1941 VSS.n472 VSS.n471 1.12329
R1942 VSS.n211 VSS.n210 1.12283
R1943 VSS.n86 VSS.t283 1.09996
R1944 VSS.n916 VSS.t279 1.09996
R1945 VSS.n926 VSS.t120 1.09996
R1946 VSS.n971 VSS.t122 1.09996
R1947 VSS.n980 VSS.t89 1.09996
R1948 VSS.n1025 VSS.t78 1.09996
R1949 VSS.n1036 VSS.t13 1.09996
R1950 VSS.n1081 VSS.t48 1.09996
R1951 VSS.n1090 VSS.t126 1.09996
R1952 VSS.n1123 VSS.t118 1.09996
R1953 VSS.n861 VSS.n859 0.755717
R1954 VSS.n122 VSS.n120 0.755717
R1955 VSS.n126 VSS.n125 0.755717
R1956 VSS.n133 VSS.n131 0.755717
R1957 VSS.n138 VSS.n137 0.755717
R1958 VSS.n143 VSS.n141 0.755717
R1959 VSS.n261 VSS.n260 0.755717
R1960 VSS.n76 VSS.n74 0.755717
R1961 VSS.n81 VSS.n80 0.755717
R1962 VSS.n66 VSS.n64 0.755717
R1963 VSS.n71 VSS.n70 0.755717
R1964 VSS.n59 VSS.n58 0.755717
R1965 VSS.n61 VSS.n60 0.755717
R1966 VSS.n52 VSS.n50 0.755717
R1967 VSS.n57 VSS.n56 0.755717
R1968 VSS.n1117 VSS.n1116 0.755717
R1969 VSS.n1119 VSS.n1118 0.755717
R1970 VSS.n45 VSS.n44 0.755717
R1971 VSS.n38 VSS.n37 0.755717
R1972 VSS.n34 VSS.n33 0.755717
R1973 VSS.n30 VSS.n29 0.755717
R1974 VSS.n28 VSS.n27 0.755717
R1975 VSS.n864 VSS.n861 0.691152
R1976 VSS.n829 VSS.n122 0.691152
R1977 VSS.n728 VSS.n126 0.691152
R1978 VSS.n723 VSS.n133 0.691152
R1979 VSS.n621 VSS.n138 0.691152
R1980 VSS.n613 VSS.n143 0.691152
R1981 VSS.n264 VSS.n261 0.691152
R1982 VSS.n85 VSS.n76 0.691152
R1983 VSS.n85 VSS.n81 0.691152
R1984 VSS.n925 VSS.n66 0.691152
R1985 VSS.n925 VSS.n71 0.691152
R1986 VSS.n1028 VSS.n59 0.691152
R1987 VSS.n1028 VSS.n61 0.691152
R1988 VSS.n1035 VSS.n52 0.691152
R1989 VSS.n1035 VSS.n57 0.691152
R1990 VSS.n1122 VSS.n1117 0.691152
R1991 VSS.n1122 VSS.n1119 0.691152
R1992 VSS.n1204 VSS.n45 0.691152
R1993 VSS.n1209 VSS.n38 0.691152
R1994 VSS.n1262 VSS.n34 0.691152
R1995 VSS.n1315 VSS.n30 0.691152
R1996 VSS.n1370 VSS.n28 0.691152
R1997 VSS.n620 VSS.n617 0.632911
R1998 VSS.n6 VSS.n3 0.559375
R1999 VSS.n1161 VSS.n1158 0.559135
R2000 VSS.n506 VSS.n496 0.472687
R2001 VSS.n506 VSS.n505 0.472687
R2002 VSS.n507 VSS.n506 0.472445
R2003 VSS.n503 VSS.n502 0.3155
R2004 VSS.n392 VSS.n391 0.3155
R2005 VSS.n171 VSS.n170 0.3155
R2006 VSS.n510 VSS.n509 0.306661
R2007 VSS.n406 VSS.n403 0.306661
R2008 VSS.n185 VSS.n182 0.306661
R2009 VSS.n342 VSS.n341 0.252261
R2010 VSS.n362 VSS.n361 0.252237
R2011 VSS.n341 VSS.n340 0.252153
R2012 VSS.n347 VSS.n344 0.186929
R2013 VSS.n366 VSS.n363 0.186929
R2014 VSS.n338 VSS.n337 0.186929
R2015 VSS.n833 VSS.n830 0.172464
R2016 VSS.n780 VSS.n777 0.172464
R2017 VSS.n727 VSS.n724 0.172464
R2018 VSS.n674 VSS.n671 0.172464
R2019 VSS.n316 VSS.n313 0.172464
R2020 VSS.n924 VSS.n921 0.172464
R2021 VSS.n979 VSS.n976 0.172464
R2022 VSS.n1034 VSS.n1031 0.172464
R2023 VSS.n1089 VSS.n1086 0.172464
R2024 VSS.n1369 VSS.n1366 0.172464
R2025 VSS.n1314 VSS.n1313 0.172464
R2026 VSS.n1208 VSS.n1207 0.172464
R2027 VSS.n529 VSS.n528 0.159607
R2028 VSS.n459 VSS.n456 0.159607
R2029 VSS.n202 VSS.n201 0.159607
R2030 VSS.n487 VSS.n486 0.158804
R2031 VSS.n423 VSS.n422 0.158804
R2032 VSS.n569 VSS.n566 0.158804
R2033 VSS.n1261 VSS 0.096125
R2034 VSS VSS.n1260 0.0768393
R2035 VSS.n350 VSS.n347 0.0760357
R2036 VSS.n353 VSS.n350 0.0760357
R2037 VSS.n482 VSS.n479 0.0760357
R2038 VSS.n551 VSS.n548 0.0760357
R2039 VSS.n548 VSS 0.0760357
R2040 VSS.n541 VSS 0.0760357
R2041 VSS.n541 VSS.n540 0.0760357
R2042 VSS.n528 VSS.n525 0.0760357
R2043 VSS.n525 VSS.n522 0.0760357
R2044 VSS.n522 VSS 0.0760357
R2045 VSS.n515 VSS 0.0760357
R2046 VSS.n515 VSS.n514 0.0760357
R2047 VSS.n508 VSS.n495 0.0760357
R2048 VSS.n502 VSS 0.0760357
R2049 VSS.n369 VSS.n366 0.0760357
R2050 VSS.n372 VSS.n369 0.0760357
R2051 VSS.n464 VSS.n463 0.0760357
R2052 VSS.n445 VSS.n442 0.0760357
R2053 VSS.n442 VSS 0.0760357
R2054 VSS.n435 VSS 0.0760357
R2055 VSS.n435 VSS.n434 0.0760357
R2056 VSS.n422 VSS.n421 0.0760357
R2057 VSS.n421 VSS.n418 0.0760357
R2058 VSS.n418 VSS 0.0760357
R2059 VSS.n411 VSS 0.0760357
R2060 VSS.n411 VSS.n410 0.0760357
R2061 VSS.n402 VSS.n401 0.0760357
R2062 VSS.n396 VSS.n395 0.0760357
R2063 VSS.n391 VSS 0.0760357
R2064 VSS.n337 VSS.n334 0.0760357
R2065 VSS.n334 VSS.n331 0.0760357
R2066 VSS.n576 VSS.n573 0.0760357
R2067 VSS.n231 VSS.n228 0.0760357
R2068 VSS.n228 VSS 0.0760357
R2069 VSS.n221 VSS 0.0760357
R2070 VSS.n221 VSS.n220 0.0760357
R2071 VSS.n201 VSS.n200 0.0760357
R2072 VSS.n200 VSS.n197 0.0760357
R2073 VSS.n197 VSS 0.0760357
R2074 VSS.n190 VSS 0.0760357
R2075 VSS.n190 VSS.n189 0.0760357
R2076 VSS.n181 VSS.n180 0.0760357
R2077 VSS.n175 VSS.n174 0.0760357
R2078 VSS.n170 VSS 0.0760357
R2079 VSS.n870 VSS.n867 0.0760357
R2080 VSS.n873 VSS.n870 0.0760357
R2081 VSS.n876 VSS.n873 0.0760357
R2082 VSS.n879 VSS.n876 0.0760357
R2083 VSS.n882 VSS.n879 0.0760357
R2084 VSS.n885 VSS.n882 0.0760357
R2085 VSS.n855 VSS.n854 0.0760357
R2086 VSS.n854 VSS.n851 0.0760357
R2087 VSS.n851 VSS.n848 0.0760357
R2088 VSS.n848 VSS.n845 0.0760357
R2089 VSS.n845 VSS.n842 0.0760357
R2090 VSS.n842 VSS.n839 0.0760357
R2091 VSS.n839 VSS.n836 0.0760357
R2092 VSS.n836 VSS.n833 0.0760357
R2093 VSS.n828 VSS.n825 0.0760357
R2094 VSS.n825 VSS.n822 0.0760357
R2095 VSS.n822 VSS.n819 0.0760357
R2096 VSS.n819 VSS.n816 0.0760357
R2097 VSS.n816 VSS.n813 0.0760357
R2098 VSS.n813 VSS.n810 0.0760357
R2099 VSS.n810 VSS.n807 0.0760357
R2100 VSS.n802 VSS.n801 0.0760357
R2101 VSS.n801 VSS.n798 0.0760357
R2102 VSS.n798 VSS.n795 0.0760357
R2103 VSS.n795 VSS.n792 0.0760357
R2104 VSS.n792 VSS.n789 0.0760357
R2105 VSS.n789 VSS.n786 0.0760357
R2106 VSS.n786 VSS.n783 0.0760357
R2107 VSS.n783 VSS.n780 0.0760357
R2108 VSS.n777 VSS.n776 0.0760357
R2109 VSS.n776 VSS.n773 0.0760357
R2110 VSS.n773 VSS.n770 0.0760357
R2111 VSS.n770 VSS.n767 0.0760357
R2112 VSS.n767 VSS.n764 0.0760357
R2113 VSS.n764 VSS.n761 0.0760357
R2114 VSS.n761 VSS.n758 0.0760357
R2115 VSS.n758 VSS.n755 0.0760357
R2116 VSS.n750 VSS.n749 0.0760357
R2117 VSS.n749 VSS.n746 0.0760357
R2118 VSS.n746 VSS.n743 0.0760357
R2119 VSS.n743 VSS.n740 0.0760357
R2120 VSS.n740 VSS.n737 0.0760357
R2121 VSS.n737 VSS.n734 0.0760357
R2122 VSS.n734 VSS.n731 0.0760357
R2123 VSS.n722 VSS.n719 0.0760357
R2124 VSS.n719 VSS.n716 0.0760357
R2125 VSS.n716 VSS.n713 0.0760357
R2126 VSS.n713 VSS.n710 0.0760357
R2127 VSS.n710 VSS.n707 0.0760357
R2128 VSS.n707 VSS.n704 0.0760357
R2129 VSS.n704 VSS.n701 0.0760357
R2130 VSS.n696 VSS.n695 0.0760357
R2131 VSS.n695 VSS.n692 0.0760357
R2132 VSS.n692 VSS.n689 0.0760357
R2133 VSS.n689 VSS.n686 0.0760357
R2134 VSS.n686 VSS.n683 0.0760357
R2135 VSS.n683 VSS.n680 0.0760357
R2136 VSS.n680 VSS.n677 0.0760357
R2137 VSS.n677 VSS.n674 0.0760357
R2138 VSS.n671 VSS.n670 0.0760357
R2139 VSS.n670 VSS.n667 0.0760357
R2140 VSS.n667 VSS.n664 0.0760357
R2141 VSS.n664 VSS.n661 0.0760357
R2142 VSS.n661 VSS.n658 0.0760357
R2143 VSS.n658 VSS.n655 0.0760357
R2144 VSS.n655 VSS.n652 0.0760357
R2145 VSS.n652 VSS.n649 0.0760357
R2146 VSS.n642 VSS.n639 0.0760357
R2147 VSS.n639 VSS.n636 0.0760357
R2148 VSS.n636 VSS.n633 0.0760357
R2149 VSS.n633 VSS.n630 0.0760357
R2150 VSS.n630 VSS.n627 0.0760357
R2151 VSS.n627 VSS.n624 0.0760357
R2152 VSS.n612 VSS.n609 0.0760357
R2153 VSS.n609 VSS.n606 0.0760357
R2154 VSS.n606 VSS.n603 0.0760357
R2155 VSS.n603 VSS.n600 0.0760357
R2156 VSS.n600 VSS.n597 0.0760357
R2157 VSS.n597 VSS.n594 0.0760357
R2158 VSS.n594 VSS.n591 0.0760357
R2159 VSS.n586 VSS.n585 0.0760357
R2160 VSS.n249 VSS.n246 0.0760357
R2161 VSS.n252 VSS.n249 0.0760357
R2162 VSS.n255 VSS.n252 0.0760357
R2163 VSS.n313 VSS.n312 0.0760357
R2164 VSS.n312 VSS.n309 0.0760357
R2165 VSS.n309 VSS.n306 0.0760357
R2166 VSS.n306 VSS.n303 0.0760357
R2167 VSS.n303 VSS.n300 0.0760357
R2168 VSS.n300 VSS.n297 0.0760357
R2169 VSS.n297 VSS.n294 0.0760357
R2170 VSS.n294 VSS.n291 0.0760357
R2171 VSS.n286 VSS.n285 0.0760357
R2172 VSS.n285 VSS.n282 0.0760357
R2173 VSS.n282 VSS.n279 0.0760357
R2174 VSS.n279 VSS.n276 0.0760357
R2175 VSS.n276 VSS.n273 0.0760357
R2176 VSS.n273 VSS.n270 0.0760357
R2177 VSS.n270 VSS.n267 0.0760357
R2178 VSS.n91 VSS.n88 0.0760357
R2179 VSS.n94 VSS.n91 0.0760357
R2180 VSS.n97 VSS.n94 0.0760357
R2181 VSS.n100 VSS.n97 0.0760357
R2182 VSS.n103 VSS.n100 0.0760357
R2183 VSS.n106 VSS.n103 0.0760357
R2184 VSS.n900 VSS.n897 0.0760357
R2185 VSS.n903 VSS.n900 0.0760357
R2186 VSS.n906 VSS.n903 0.0760357
R2187 VSS.n909 VSS.n906 0.0760357
R2188 VSS.n912 VSS.n909 0.0760357
R2189 VSS.n915 VSS.n912 0.0760357
R2190 VSS.n918 VSS.n915 0.0760357
R2191 VSS.n921 VSS.n918 0.0760357
R2192 VSS.n931 VSS.n928 0.0760357
R2193 VSS.n934 VSS.n931 0.0760357
R2194 VSS.n937 VSS.n934 0.0760357
R2195 VSS.n940 VSS.n937 0.0760357
R2196 VSS.n943 VSS.n940 0.0760357
R2197 VSS.n946 VSS.n943 0.0760357
R2198 VSS.n947 VSS.n946 0.0760357
R2199 VSS.n955 VSS.n952 0.0760357
R2200 VSS.n958 VSS.n955 0.0760357
R2201 VSS.n961 VSS.n958 0.0760357
R2202 VSS.n964 VSS.n961 0.0760357
R2203 VSS.n967 VSS.n964 0.0760357
R2204 VSS.n970 VSS.n967 0.0760357
R2205 VSS.n973 VSS.n970 0.0760357
R2206 VSS.n976 VSS.n973 0.0760357
R2207 VSS.n982 VSS.n979 0.0760357
R2208 VSS.n985 VSS.n982 0.0760357
R2209 VSS.n988 VSS.n985 0.0760357
R2210 VSS.n991 VSS.n988 0.0760357
R2211 VSS.n994 VSS.n991 0.0760357
R2212 VSS.n997 VSS.n994 0.0760357
R2213 VSS.n1000 VSS.n997 0.0760357
R2214 VSS.n1001 VSS.n1000 0.0760357
R2215 VSS.n1009 VSS.n1006 0.0760357
R2216 VSS.n1012 VSS.n1009 0.0760357
R2217 VSS.n1015 VSS.n1012 0.0760357
R2218 VSS.n1018 VSS.n1015 0.0760357
R2219 VSS.n1021 VSS.n1018 0.0760357
R2220 VSS.n1024 VSS.n1021 0.0760357
R2221 VSS.n1027 VSS.n1024 0.0760357
R2222 VSS.n1041 VSS.n1038 0.0760357
R2223 VSS.n1044 VSS.n1041 0.0760357
R2224 VSS.n1047 VSS.n1044 0.0760357
R2225 VSS.n1050 VSS.n1047 0.0760357
R2226 VSS.n1053 VSS.n1050 0.0760357
R2227 VSS.n1056 VSS.n1053 0.0760357
R2228 VSS.n1057 VSS.n1056 0.0760357
R2229 VSS.n1065 VSS.n1062 0.0760357
R2230 VSS.n1068 VSS.n1065 0.0760357
R2231 VSS.n1071 VSS.n1068 0.0760357
R2232 VSS.n1074 VSS.n1071 0.0760357
R2233 VSS.n1077 VSS.n1074 0.0760357
R2234 VSS.n1080 VSS.n1077 0.0760357
R2235 VSS.n1083 VSS.n1080 0.0760357
R2236 VSS.n1086 VSS.n1083 0.0760357
R2237 VSS.n1092 VSS.n1089 0.0760357
R2238 VSS.n1095 VSS.n1092 0.0760357
R2239 VSS.n1098 VSS.n1095 0.0760357
R2240 VSS.n1101 VSS.n1098 0.0760357
R2241 VSS.n1104 VSS.n1101 0.0760357
R2242 VSS.n1107 VSS.n1104 0.0760357
R2243 VSS.n1110 VSS.n1107 0.0760357
R2244 VSS.n1111 VSS.n1110 0.0760357
R2245 VSS.n1143 VSS.n1140 0.0760357
R2246 VSS.n1140 VSS.n1137 0.0760357
R2247 VSS.n1137 VSS.n1134 0.0760357
R2248 VSS.n1134 VSS.n1131 0.0760357
R2249 VSS.n1131 VSS.n1128 0.0760357
R2250 VSS.n1128 VSS.n1125 0.0760357
R2251 VSS.n9 VSS.n6 0.0760357
R2252 VSS.n12 VSS.n9 0.0760357
R2253 VSS.n15 VSS.n12 0.0760357
R2254 VSS.n18 VSS.n15 0.0760357
R2255 VSS.n21 VSS.n18 0.0760357
R2256 VSS.n1394 VSS.n1391 0.0760357
R2257 VSS.n1391 VSS.n1388 0.0760357
R2258 VSS.n1388 VSS.n1385 0.0760357
R2259 VSS.n1385 VSS.n1382 0.0760357
R2260 VSS.n1382 VSS.n1379 0.0760357
R2261 VSS.n1379 VSS.n1376 0.0760357
R2262 VSS.n1376 VSS.n1373 0.0760357
R2263 VSS.n1366 VSS.n1363 0.0760357
R2264 VSS.n1363 VSS.n1360 0.0760357
R2265 VSS.n1360 VSS.n1357 0.0760357
R2266 VSS.n1357 VSS.n1354 0.0760357
R2267 VSS.n1354 VSS.n1351 0.0760357
R2268 VSS.n1351 VSS.n1348 0.0760357
R2269 VSS.n1348 VSS.n1345 0.0760357
R2270 VSS.n1345 VSS.n1342 0.0760357
R2271 VSS.n1337 VSS.n1336 0.0760357
R2272 VSS.n1336 VSS.n1333 0.0760357
R2273 VSS.n1333 VSS.n1330 0.0760357
R2274 VSS.n1330 VSS.n1327 0.0760357
R2275 VSS.n1327 VSS.n1324 0.0760357
R2276 VSS.n1324 VSS.n1321 0.0760357
R2277 VSS.n1321 VSS.n1318 0.0760357
R2278 VSS.n1313 VSS.n1310 0.0760357
R2279 VSS.n1310 VSS.n1307 0.0760357
R2280 VSS.n1307 VSS.n1304 0.0760357
R2281 VSS.n1304 VSS.n1301 0.0760357
R2282 VSS.n1301 VSS.n1298 0.0760357
R2283 VSS.n1298 VSS.n1295 0.0760357
R2284 VSS.n1295 VSS.n1292 0.0760357
R2285 VSS.n1292 VSS.n1289 0.0760357
R2286 VSS.n1284 VSS.n1283 0.0760357
R2287 VSS.n1283 VSS.n1280 0.0760357
R2288 VSS.n1280 VSS.n1277 0.0760357
R2289 VSS.n1277 VSS.n1274 0.0760357
R2290 VSS.n1274 VSS.n1271 0.0760357
R2291 VSS.n1271 VSS.n1268 0.0760357
R2292 VSS.n1268 VSS.n1265 0.0760357
R2293 VSS.n1260 VSS.n1257 0.0760357
R2294 VSS.n1257 VSS.n1254 0.0760357
R2295 VSS.n1254 VSS.n1251 0.0760357
R2296 VSS.n1251 VSS.n1248 0.0760357
R2297 VSS.n1248 VSS.n1245 0.0760357
R2298 VSS.n1245 VSS.n1242 0.0760357
R2299 VSS.n1242 VSS.n1239 0.0760357
R2300 VSS.n1239 VSS.n1236 0.0760357
R2301 VSS.n1231 VSS.n1230 0.0760357
R2302 VSS.n1230 VSS.n1227 0.0760357
R2303 VSS.n1227 VSS.n1224 0.0760357
R2304 VSS.n1224 VSS.n1221 0.0760357
R2305 VSS.n1221 VSS.n1218 0.0760357
R2306 VSS.n1218 VSS.n1215 0.0760357
R2307 VSS.n1215 VSS.n1212 0.0760357
R2308 VSS.n1203 VSS.n1200 0.0760357
R2309 VSS.n1200 VSS.n1197 0.0760357
R2310 VSS.n1197 VSS.n1194 0.0760357
R2311 VSS.n1194 VSS.n1191 0.0760357
R2312 VSS.n1191 VSS.n1188 0.0760357
R2313 VSS.n1188 VSS.n1185 0.0760357
R2314 VSS.n1185 VSS.n1182 0.0760357
R2315 VSS.n1176 VSS.n1173 0.0760357
R2316 VSS.n1173 VSS.n1170 0.0760357
R2317 VSS.n1170 VSS.n1167 0.0760357
R2318 VSS.n1167 VSS.n1164 0.0760357
R2319 VSS.n1164 VSS.n1161 0.0760357
R2320 VSS.n1177 VSS.n1176 0.0728317
R2321 VSS.n483 VSS.n482 0.0728214
R2322 VSS.n514 VSS.n511 0.0728214
R2323 VSS.n463 VSS.n460 0.0728214
R2324 VSS.n410 VSS.n407 0.0728214
R2325 VSS.n573 VSS.n570 0.0728214
R2326 VSS.n189 VSS.n186 0.0728214
R2327 VSS.n319 VSS.n255 0.070727
R2328 VSS.n246 VSS.n243 0.0704107
R2329 VSS.n886 VSS.n885 0.0668722
R2330 VSS.n22 VSS.n21 0.0668722
R2331 VSS.n643 VSS.n642 0.0664687
R2332 VSS.n343 VSS 0.0647857
R2333 VSS VSS.n500 0.0647857
R2334 VSS VSS.n360 0.0647857
R2335 VSS VSS.n386 0.0647857
R2336 VSS VSS.n339 0.0647857
R2337 VSS VSS.n164 0.0647857
R2338 VSS.n867 VSS.n864 0.0639821
R2339 VSS.n829 VSS.n828 0.0639821
R2340 VSS.n731 VSS.n728 0.0639821
R2341 VSS.n723 VSS.n722 0.0639821
R2342 VSS.n624 VSS.n621 0.0639821
R2343 VSS.n613 VSS.n612 0.0639821
R2344 VSS.n267 VSS.n264 0.0639821
R2345 VSS.n88 VSS.n85 0.0639821
R2346 VSS.n928 VSS.n925 0.0639821
R2347 VSS.n1028 VSS.n1027 0.0639821
R2348 VSS.n1038 VSS.n1035 0.0639821
R2349 VSS.n1125 VSS.n1122 0.0639821
R2350 VSS.n1373 VSS.n1370 0.0639821
R2351 VSS.n1318 VSS.n1315 0.0639821
R2352 VSS.n1265 VSS.n1262 0.0639821
R2353 VSS.n1212 VSS.n1209 0.0639821
R2354 VSS.n1204 VSS.n1203 0.0639821
R2355 VSS.n354 VSS.n353 0.05675
R2356 VSS.n552 VSS.n551 0.05675
R2357 VSS.n373 VSS.n372 0.05675
R2358 VSS.n434 VSS.n431 0.05675
R2359 VSS.n331 VSS.n151 0.05675
R2360 VSS.n232 VSS.n231 0.05675
R2361 VSS.n107 VSS.n106 0.05675
R2362 VSS.n479 VSS.n326 0.0559464
R2363 VSS.n540 VSS.n537 0.0559464
R2364 VSS.n464 VSS.n375 0.0559464
R2365 VSS.n446 VSS.n445 0.0559464
R2366 VSS.n577 VSS.n576 0.0559464
R2367 VSS.n220 VSS.n217 0.0559464
R2368 VSS.n317 VSS.n316 0.0559464
R2369 VSS.n1144 VSS.n1143 0.0559464
R2370 VSS VSS.n495 0.0422857
R2371 VSS.n401 VSS 0.0422857
R2372 VSS.n180 VSS 0.0422857
R2373 VSS.n807 VSS 0.0422857
R2374 VSS.n750 VSS 0.0422857
R2375 VSS.n701 VSS 0.0422857
R2376 VSS.n591 VSS 0.0422857
R2377 VSS.n585 VSS.n584 0.0422857
R2378 VSS.n286 VSS 0.0422857
R2379 VSS.n947 VSS 0.0422857
R2380 VSS.n1006 VSS 0.0422857
R2381 VSS.n1057 VSS 0.0422857
R2382 VSS VSS.n1394 0.0422857
R2383 VSS.n1337 VSS 0.0422857
R2384 VSS.n1284 VSS 0.0422857
R2385 VSS.n1231 VSS 0.0422857
R2386 VSS.n1182 VSS 0.0422857
R2387 VSS.n1146 VSS 0.0363205
R2388 VSS.n498 VSS 0.03425
R2389 VSS.n396 VSS 0.03425
R2390 VSS.n175 VSS 0.03425
R2391 VSS VSS.n855 0.03425
R2392 VSS.n802 VSS 0.03425
R2393 VSS.n755 VSS 0.03425
R2394 VSS.n696 VSS 0.03425
R2395 VSS.n649 VSS 0.03425
R2396 VSS.n586 VSS 0.03425
R2397 VSS.n291 VSS 0.03425
R2398 VSS.n897 VSS 0.03425
R2399 VSS.n952 VSS 0.03425
R2400 VSS.n1001 VSS 0.03425
R2401 VSS.n1062 VSS 0.03425
R2402 VSS.n1111 VSS 0.03425
R2403 VSS.n1342 VSS 0.03425
R2404 VSS.n1289 VSS 0.03425
R2405 VSS.n1236 VSS 0.03425
R2406 VSS.n136 VSS 0.0331222
R2407 VSS.n856 VSS 0.0327187
R2408 VSS.n428 VSS.n427 0.0301053
R2409 VSS.n454 VSS.n453 0.0301053
R2410 VSS.n578 VSS.n150 0.0301053
R2411 VSS.n474 VSS.n355 0.0289211
R2412 VSS.n428 VSS.n424 0.0289211
R2413 VSS.n213 VSS.n212 0.0289211
R2414 VSS.n534 VSS.n531 0.0289211
R2415 VSS.n533 VSS.n532 0.0289211
R2416 VSS.n557 VSS.n323 0.0289211
R2417 VSS.n325 VSS.n324 0.0289211
R2418 VSS.n564 VSS.n234 0.0289211
R2419 VSS.n563 VSS.n562 0.0289211
R2420 VSS.n454 VSS.n449 0.0289211
R2421 VSS.n469 VSS.n359 0.0289211
R2422 VSS.n471 VSS.n470 0.0289211
R2423 VSS.n578 VSS.n149 0.0289211
R2424 VSS VSS.n26 0.024683
R2425 VSS.n208 VSS.n207 0.0221964
R2426 VSS.n210 VSS.n209 0.0221964
R2427 VSS.n451 VSS.n322 0.0221964
R2428 VSS.n560 VSS.n559 0.0221964
R2429 VSS.n357 VSS.n148 0.0221964
R2430 VSS.n581 VSS.n580 0.0221964
R2431 VSS.n108 VSS 0.0221964
R2432 VSS VSS.n326 0.0205893
R2433 VSS.n455 VSS.n446 0.0205893
R2434 VSS.n429 VSS.n423 0.0205893
R2435 VSS VSS.n577 0.0205893
R2436 VSS.n318 VSS.n317 0.0205893
R2437 VSS.n890 VSS.n889 0.0205893
R2438 VSS.n892 VSS.n108 0.0205893
R2439 VSS.n1145 VSS.n1144 0.0205893
R2440 VSS.n1153 VSS.n1152 0.0205893
R2441 VSS.n1150 VSS.n1149 0.0205893
R2442 VSS VSS.n354 0.0197857
R2443 VSS.n556 VSS.n487 0.0197857
R2444 VSS.n555 VSS.n552 0.0197857
R2445 VSS.n530 VSS.n529 0.0197857
R2446 VSS VSS.n373 0.0197857
R2447 VSS.n375 VSS.n374 0.0197857
R2448 VSS.n456 VSS.n455 0.0197857
R2449 VSS VSS.n151 0.0197857
R2450 VSS.n566 VSS.n565 0.0197857
R2451 VSS.n233 VSS.n232 0.0197857
R2452 VSS.n205 VSS.n202 0.0197857
R2453 VSS.n892 VSS.n107 0.0197857
R2454 VSS.n1151 VSS.n1150 0.0197857
R2455 VSS.n1181 VSS.n1180 0.0197857
R2456 VSS.n537 VSS.n536 0.017375
R2457 VSS.n217 VSS.n216 0.017375
R2458 VSS.n431 VSS.n430 0.0165714
R2459 VSS.n509 VSS.n508 0.0157679
R2460 VSS.n504 VSS.n503 0.0157679
R2461 VSS.n403 VSS.n402 0.0157679
R2462 VSS.n395 VSS.n392 0.0157679
R2463 VSS.n182 VSS.n181 0.0157679
R2464 VSS.n174 VSS.n171 0.0157679
R2465 VSS VSS.n1181 0.0149643
R2466 VSS.n240 VSS.n237 0.0133571
R2467 VSS.n830 VSS.n829 0.0125536
R2468 VSS.n728 VSS.n727 0.0125536
R2469 VSS.n724 VSS.n723 0.0125536
R2470 VSS.n621 VSS.n620 0.0125536
R2471 VSS.n617 VSS.n613 0.0125536
R2472 VSS.n925 VSS.n924 0.0125536
R2473 VSS.n1031 VSS.n1028 0.0125536
R2474 VSS.n1035 VSS.n1034 0.0125536
R2475 VSS.n1370 VSS.n1369 0.0125536
R2476 VSS.n1315 VSS.n1314 0.0125536
R2477 VSS.n1262 VSS.n1261 0.0125536
R2478 VSS.n1209 VSS.n1208 0.0125536
R2479 VSS.n1207 VSS.n1204 0.0125536
R2480 VSS.n473 VSS.n357 0.0118221
R2481 VSS.n344 VSS.n343 0.01175
R2482 VSS.n363 VSS.n360 0.01175
R2483 VSS.n339 VSS.n338 0.01175
R2484 VSS.n110 VSS.n109 0.0110437
R2485 VSS.n644 VSS.n643 0.0110223
R2486 VSS.n26 VSS.n25 0.0110223
R2487 VSS.n888 VSS.n887 0.0106437
R2488 VSS.n1148 VSS.n1147 0.0106437
R2489 VSS.n582 VSS.n147 0.0106222
R2490 VSS.n321 VSS.n320 0.0106222
R2491 VSS.n644 VSS.n136 0.0106222
R2492 VSS.n25 VSS.n22 0.0106222
R2493 VSS.n583 VSS.n146 0.00903929
R2494 VSS.n237 VSS.n146 0.00900356
R2495 VSS.n207 VSS.n206 0.00820897
R2496 VSS.n561 VSS.n560 0.00820897
R2497 VSS.n558 VSS.n322 0.00820897
R2498 VSS.n580 VSS.n579 0.00820897
R2499 VSS.n214 VSS.n211 0.00807964
R2500 VSS.n319 VSS.n318 0.00775238
R2501 VSS.n891 VSS.n890 0.00741026
R2502 VSS.n1146 VSS.n1145 0.00741026
R2503 VSS.n426 VSS.n425 0.00703287
R2504 VSS.n1180 VSS.n1177 0.0066335
R2505 VSS.n452 VSS.n450 0.00641377
R2506 VSS.n472 VSS.n358 0.00641106
R2507 VSS.n243 VSS.n240 0.006125
R2508 VSS.n584 VSS.n583 0.00532143
R2509 VSS.n486 VSS.n483 0.00371429
R2510 VSS.n511 VSS.n510 0.00371429
R2511 VSS.n460 VSS.n459 0.00371429
R2512 VSS.n430 VSS.n429 0.00371429
R2513 VSS.n407 VSS.n406 0.00371429
R2514 VSS.n570 VSS.n569 0.00371429
R2515 VSS.n186 VSS.n185 0.00371429
R2516 VSS.n536 VSS.n535 0.00291071
R2517 VSS.n216 VSS.n215 0.00291071
R2518 VSS.n214 VSS.n213 0.00168421
R2519 VSS.n534 VSS.n533 0.00168421
R2520 VSS.n557 VSS.n325 0.00168421
R2521 VSS.n564 VSS.n563 0.00168421
R2522 VSS.n471 VSS.n469 0.00168421
R2523 VSS.n556 VSS.n555 0.00130357
R2524 VSS.n535 VSS.n530 0.00130357
R2525 VSS VSS.n374 0.00130357
R2526 VSS.n565 VSS.n233 0.00130357
R2527 VSS.n215 VSS.n205 0.00130357
R2528 EN.t142 EN.t212 82.9076
R2529 EN.t53 EN.t142 82.9076
R2530 EN.t166 EN.t16 82.9076
R2531 EN.t100 EN.t166 82.9076
R2532 EN.t69 EN.t36 82.9076
R2533 EN.t201 EN.t69 82.9076
R2534 EN.t52 EN.t162 82.9076
R2535 EN.t127 EN.t52 82.9076
R2536 EN.t175 EN.t34 82.9076
R2537 EN.t14 EN.t175 82.9076
R2538 EN.t60 EN.t165 82.9076
R2539 EN.t130 EN.t60 82.9076
R2540 EN.t199 EN.t67 82.9076
R2541 EN.t31 EN.t199 82.9076
R2542 EN.t112 EN.t221 82.9076
R2543 EN.t189 EN.t112 82.9076
R2544 EN.t108 EN.n225 56.4451
R2545 EN.n112 EN.t53 49.7969
R2546 EN.n82 EN.t100 49.7969
R2547 EN.n53 EN.t201 49.7969
R2548 EN.n143 EN.t127 49.7969
R2549 EN.n177 EN.t14 49.7969
R2550 EN.n211 EN.t130 49.7969
R2551 EN.n25 EN.t31 49.7969
R2552 EN.n244 EN.t189 49.7969
R2553 EN.n219 EN.t227 39.7594
R2554 EN.n111 EN.n110 35.0405
R2555 EN.n59 EN.n58 35.0405
R2556 EN.n81 EN.n80 35.0405
R2557 EN.n52 EN.n51 35.0405
R2558 EN.n120 EN.n119 35.0405
R2559 EN.n142 EN.n141 35.0405
R2560 EN.n154 EN.n153 35.0405
R2561 EN.n176 EN.n175 35.0405
R2562 EN.n210 EN.n209 35.0405
R2563 EN.n2 EN.n1 35.0405
R2564 EN.n24 EN.n23 35.0405
R2565 EN.n227 EN.n226 35.0405
R2566 EN.n243 EN.n242 35.0405
R2567 EN.n112 EN.t141 31.1559
R2568 EN.n82 EN.t200 31.1559
R2569 EN.n53 EN.t48 31.1559
R2570 EN.n143 EN.t183 31.1559
R2571 EN.n177 EN.t74 31.1559
R2572 EN.n211 EN.t185 31.1559
R2573 EN.n25 EN.t92 31.1559
R2574 EN.n244 EN.t10 31.1559
R2575 EN.t47 EN.n87 21.9005
R2576 EN.t46 EN.n95 21.9005
R2577 EN.t73 EN.n97 21.9005
R2578 EN.t207 EN.n101 21.9005
R2579 EN.t68 EN.n102 21.9005
R2580 EN.t97 EN.n59 21.9005
R2581 EN.t87 EN.n63 21.9005
R2582 EN.t222 EN.n65 21.9005
R2583 EN.t146 EN.n67 21.9005
R2584 EN.t218 EN.n72 21.9005
R2585 EN.t226 EN.n28 21.9005
R2586 EN.t90 EN.n30 21.9005
R2587 EN.t217 EN.n34 21.9005
R2588 EN.t84 EN.n36 21.9005
R2589 EN.t239 EN.n38 21.9005
R2590 EN.t41 EN.n40 21.9005
R2591 EN.t178 EN.n43 21.9005
R2592 EN.t235 EN.n133 21.9005
R2593 EN.t135 EN.n128 21.9005
R2594 EN.t125 EN.n122 21.9005
R2595 EN.t114 EN.n120 21.9005
R2596 EN.t104 EN.n167 21.9005
R2597 EN.t190 EN.n164 21.9005
R2598 EN.t96 EN.n158 21.9005
R2599 EN.t0 EN.n154 21.9005
R2600 EN.t171 EN.n201 21.9005
R2601 EN.t3 EN.n196 21.9005
R2602 EN.t85 EN.n194 21.9005
R2603 EN.t148 EN.n190 21.9005
R2604 EN.t116 EN.n186 21.9005
R2605 EN.t160 EN.n188 21.9005
R2606 EN.t59 EN.n15 21.9005
R2607 EN.t197 EN.n14 21.9005
R2608 EN.t194 EN.n10 21.9005
R2609 EN.t203 EN.n6 21.9005
R2610 EN.t28 EN.n4 21.9005
R2611 EN.t19 EN.n2 21.9005
R2612 EN.n226 EN.t177 21.9005
R2613 EN.n227 EN.t159 21.9005
R2614 EN.n228 EN.t233 21.9005
R2615 EN.n229 EN.t70 21.9005
R2616 EN.n230 EN.t82 21.9005
R2617 EN.n231 EN.t140 21.9005
R2618 EN.n232 EN.t152 21.9005
R2619 EN.n233 EN.t224 21.9005
R2620 EN.t49 EN.n234 21.9005
R2621 EN.n111 EN.t47 21.5094
R2622 EN.n110 EN.t46 21.5094
R2623 EN.n109 EN.t12 21.5094
R2624 EN.n108 EN.t145 21.5094
R2625 EN.n107 EN.t38 21.5094
R2626 EN.n106 EN.t73 21.5094
R2627 EN.n105 EN.t207 21.5094
R2628 EN.n104 EN.t168 21.5094
R2629 EN.n103 EN.t68 21.5094
R2630 EN.n81 EN.t97 21.5094
R2631 EN.n80 EN.t80 21.5094
R2632 EN.n79 EN.t87 21.5094
R2633 EN.n78 EN.t151 21.5094
R2634 EN.n77 EN.t222 21.5094
R2635 EN.n76 EN.t146 21.5094
R2636 EN.n75 EN.t218 21.5094
R2637 EN.n74 EN.t229 21.5094
R2638 EN.n73 EN.t57 21.5094
R2639 EN.n52 EN.t226 21.5094
R2640 EN.n51 EN.t90 21.5094
R2641 EN.n50 EN.t217 21.5094
R2642 EN.n49 EN.t25 21.5094
R2643 EN.n48 EN.t84 21.5094
R2644 EN.n47 EN.t239 21.5094
R2645 EN.n46 EN.t41 21.5094
R2646 EN.n45 EN.t178 21.5094
R2647 EN.n44 EN.t234 21.5094
R2648 EN.n134 EN.t154 21.5094
R2649 EN.n135 EN.t228 21.5094
R2650 EN.n136 EN.t235 21.5094
R2651 EN.n137 EN.t65 21.5094
R2652 EN.n138 EN.t76 21.5094
R2653 EN.n139 EN.t135 21.5094
R2654 EN.n140 EN.t125 21.5094
R2655 EN.n142 EN.t114 21.5094
R2656 EN.n141 EN.t133 21.5094
R2657 EN.n168 EN.t111 21.5094
R2658 EN.n169 EN.t104 21.5094
R2659 EN.n170 EN.t109 21.5094
R2660 EN.n171 EN.t180 21.5094
R2661 EN.n172 EN.t190 21.5094
R2662 EN.n173 EN.t20 21.5094
R2663 EN.n174 EN.t96 21.5094
R2664 EN.n176 EN.t0 21.5094
R2665 EN.n175 EN.t17 21.5094
R2666 EN.n202 EN.t174 21.5094
R2667 EN.n203 EN.t8 21.5094
R2668 EN.n204 EN.t171 21.5094
R2669 EN.n205 EN.t3 21.5094
R2670 EN.n206 EN.t79 21.5094
R2671 EN.n207 EN.t85 21.5094
R2672 EN.n208 EN.t148 21.5094
R2673 EN.n210 EN.t116 21.5094
R2674 EN.n209 EN.t160 21.5094
R2675 EN.n16 EN.t59 21.5094
R2676 EN.n17 EN.t123 21.5094
R2677 EN.n18 EN.t197 21.5094
R2678 EN.n19 EN.t119 21.5094
R2679 EN.n20 EN.t194 21.5094
R2680 EN.n21 EN.t203 21.5094
R2681 EN.n22 EN.t28 21.5094
R2682 EN.n24 EN.t19 21.5094
R2683 EN.n23 EN.t102 21.5094
R2684 EN.n243 EN.t177 21.5094
R2685 EN.n242 EN.t159 21.5094
R2686 EN.n241 EN.t233 21.5094
R2687 EN.n240 EN.t70 21.5094
R2688 EN.n239 EN.t82 21.5094
R2689 EN.n238 EN.t140 21.5094
R2690 EN.n237 EN.t152 21.5094
R2691 EN.n236 EN.t224 21.5094
R2692 EN.n235 EN.t49 21.5094
R2693 EN.n110 EN.t118 20.988
R2694 EN.n109 EN.t129 20.988
R2695 EN.n108 EN.t204 20.988
R2696 EN.n107 EN.t29 20.988
R2697 EN.n106 EN.t202 20.988
R2698 EN.n105 EN.t26 20.988
R2699 EN.n104 EN.t33 20.988
R2700 EN.n103 EN.t107 20.988
R2701 EN.t141 EN.n111 20.988
R2702 EN.n80 EN.t66 20.988
R2703 EN.n79 EN.t195 20.988
R2704 EN.n78 EN.t7 20.988
R2705 EN.n77 EN.t54 20.988
R2706 EN.n76 EN.t215 20.988
R2707 EN.n75 EN.t23 20.988
R2708 EN.n74 EN.t158 20.988
R2709 EN.n73 EN.t210 20.988
R2710 EN.t200 EN.n81 20.988
R2711 EN.n51 EN.t156 20.988
R2712 EN.n50 EN.t37 20.988
R2713 EN.n49 EN.t98 20.988
R2714 EN.n48 EN.t143 20.988
R2715 EN.n47 EN.t72 20.988
R2716 EN.n46 EN.t113 20.988
R2717 EN.n45 EN.t11 20.988
R2718 EN.n44 EN.t62 20.988
R2719 EN.t48 EN.n52 20.988
R2720 EN.n134 EN.t225 20.988
R2721 EN.n135 EN.t50 20.988
R2722 EN.n136 EN.t64 20.988
R2723 EN.n137 EN.t126 20.988
R2724 EN.n138 EN.t134 20.988
R2725 EN.n139 EN.t213 20.988
R2726 EN.n140 EN.t198 20.988
R2727 EN.n141 EN.t209 20.988
R2728 EN.t183 EN.n142 20.988
R2729 EN.n168 EN.t181 20.988
R2730 EN.n169 EN.t172 20.988
R2731 EN.n170 EN.t179 20.988
R2732 EN.n171 EN.t13 20.988
R2733 EN.n172 EN.t18 20.988
R2734 EN.n173 EN.t93 20.988
R2735 EN.n174 EN.t161 20.988
R2736 EN.n175 EN.t91 20.988
R2737 EN.t74 EN.n176 20.988
R2738 EN.n202 EN.t6 20.988
R2739 EN.n203 EN.t81 20.988
R2740 EN.n204 EN.t1 20.988
R2741 EN.n205 EN.t77 20.988
R2742 EN.n206 EN.t136 20.988
R2743 EN.n207 EN.t147 20.988
R2744 EN.n208 EN.t219 20.988
R2745 EN.n209 EN.t231 20.988
R2746 EN.t185 EN.n210 20.988
R2747 EN.n16 EN.t122 20.988
R2748 EN.n17 EN.t196 20.988
R2749 EN.n18 EN.t24 20.988
R2750 EN.n19 EN.t191 20.988
R2751 EN.n20 EN.t21 20.988
R2752 EN.n21 EN.t27 20.988
R2753 EN.n22 EN.t101 20.988
R2754 EN.n23 EN.t169 20.988
R2755 EN.t92 EN.n24 20.988
R2756 EN.n242 EN.t230 20.988
R2757 EN.n241 EN.t58 20.988
R2758 EN.n240 EN.t128 20.988
R2759 EN.n239 EN.t139 20.988
R2760 EN.n238 EN.t214 20.988
R2761 EN.n237 EN.t223 20.988
R2762 EN.n236 EN.t45 20.988
R2763 EN.n235 EN.t115 20.988
R2764 EN.t10 EN.n243 20.988
R2765 EN.n225 EN.n224 20.8576
R2766 EN.n224 EN.n223 20.8576
R2767 EN.n223 EN.n222 20.8576
R2768 EN.n222 EN.n221 20.8576
R2769 EN.n221 EN.n220 20.8576
R2770 EN.n220 EN.n219 20.8576
R2771 EN.n87 EN.t188 20.5969
R2772 EN.n95 EN.t187 20.5969
R2773 EN.n94 EN.t149 20.5969
R2774 EN.n93 EN.t43 20.5969
R2775 EN.n92 EN.t184 20.5969
R2776 EN.n97 EN.t211 20.5969
R2777 EN.n101 EN.t105 20.5969
R2778 EN.n102 EN.t206 20.5969
R2779 EN.n100 EN.t71 20.5969
R2780 EN.n70 EN.t121 20.5969
R2781 EN.n72 EN.t39 20.5969
R2782 EN.n67 EN.t216 20.5969
R2783 EN.n65 EN.t44 20.5969
R2784 EN.n62 EN.t220 20.5969
R2785 EN.n63 EN.t150 20.5969
R2786 EN.n58 EN.t138 20.5969
R2787 EN.n59 EN.t164 20.5969
R2788 EN.n71 EN.t56 20.5969
R2789 EN.n28 EN.t137 20.5969
R2790 EN.n30 EN.t5 20.5969
R2791 EN.n34 EN.t132 20.5969
R2792 EN.n33 EN.t182 20.5969
R2793 EN.n36 EN.t238 20.5969
R2794 EN.n38 EN.t157 20.5969
R2795 EN.n40 EN.t208 20.5969
R2796 EN.n42 EN.t144 20.5969
R2797 EN.n43 EN.t99 20.5969
R2798 EN.n119 EN.t75 20.5969
R2799 EN.n122 EN.t63 20.5969
R2800 EN.n128 EN.t78 20.5969
R2801 EN.n127 EN.t2 20.5969
R2802 EN.n126 EN.t236 20.5969
R2803 EN.n133 EN.t167 20.5969
R2804 EN.n132 EN.t155 20.5969
R2805 EN.n131 EN.t89 20.5969
R2806 EN.n120 EN.t42 20.5969
R2807 EN.n153 EN.t186 20.5969
R2808 EN.n158 EN.t22 20.5969
R2809 EN.n157 EN.t193 20.5969
R2810 EN.n164 EN.t117 20.5969
R2811 EN.n163 EN.t110 20.5969
R2812 EN.n162 EN.t35 20.5969
R2813 EN.n167 EN.t32 20.5969
R2814 EN.n166 EN.t40 20.5969
R2815 EN.n154 EN.t170 20.5969
R2816 EN.n188 EN.t95 20.5969
R2817 EN.n190 EN.t86 20.5969
R2818 EN.n194 EN.t15 20.5969
R2819 EN.n193 EN.t4 20.5969
R2820 EN.n196 EN.t173 20.5969
R2821 EN.n201 EN.t103 20.5969
R2822 EN.n200 EN.t176 20.5969
R2823 EN.n199 EN.t106 20.5969
R2824 EN.n186 EN.t51 20.5969
R2825 EN.n1 EN.t30 20.5969
R2826 EN.n4 EN.t205 20.5969
R2827 EN.n6 EN.t131 20.5969
R2828 EN.n10 EN.t120 20.5969
R2829 EN.n9 EN.t55 20.5969
R2830 EN.n14 EN.t124 20.5969
R2831 EN.n13 EN.t61 20.5969
R2832 EN.n15 EN.t232 20.5969
R2833 EN.n2 EN.t192 20.5969
R2834 EN.n234 EN.t227 20.5969
R2835 EN.n232 EN.t88 20.5969
R2836 EN.n231 EN.t83 20.5969
R2837 EN.n230 EN.t9 20.5969
R2838 EN.n229 EN.t237 20.5969
R2839 EN.n228 EN.t163 20.5969
R2840 EN.n227 EN.t94 20.5969
R2841 EN.n226 EN.t108 20.5969
R2842 EN.n233 EN.t153 20.5969
R2843 EN.n95 EN.n94 19.4672
R2844 EN.n94 EN.n93 19.4672
R2845 EN.n93 EN.n92 19.4672
R2846 EN.n101 EN.n100 19.4672
R2847 EN.n110 EN.n109 19.4672
R2848 EN.n109 EN.n108 19.4672
R2849 EN.n108 EN.n107 19.4672
R2850 EN.n107 EN.n106 19.4672
R2851 EN.n106 EN.n105 19.4672
R2852 EN.n105 EN.n104 19.4672
R2853 EN.n104 EN.n103 19.4672
R2854 EN.n63 EN.n62 19.4672
R2855 EN.n72 EN.n71 19.4672
R2856 EN.n71 EN.n70 19.4672
R2857 EN.n80 EN.n79 19.4672
R2858 EN.n79 EN.n78 19.4672
R2859 EN.n78 EN.n77 19.4672
R2860 EN.n77 EN.n76 19.4672
R2861 EN.n76 EN.n75 19.4672
R2862 EN.n75 EN.n74 19.4672
R2863 EN.n74 EN.n73 19.4672
R2864 EN.n34 EN.n33 19.4672
R2865 EN.n43 EN.n42 19.4672
R2866 EN.n51 EN.n50 19.4672
R2867 EN.n50 EN.n49 19.4672
R2868 EN.n49 EN.n48 19.4672
R2869 EN.n48 EN.n47 19.4672
R2870 EN.n47 EN.n46 19.4672
R2871 EN.n46 EN.n45 19.4672
R2872 EN.n45 EN.n44 19.4672
R2873 EN.n132 EN.n131 19.4672
R2874 EN.n133 EN.n132 19.4672
R2875 EN.n127 EN.n126 19.4672
R2876 EN.n128 EN.n127 19.4672
R2877 EN.n135 EN.n134 19.4672
R2878 EN.n136 EN.n135 19.4672
R2879 EN.n137 EN.n136 19.4672
R2880 EN.n138 EN.n137 19.4672
R2881 EN.n139 EN.n138 19.4672
R2882 EN.n140 EN.n139 19.4672
R2883 EN.n141 EN.n140 19.4672
R2884 EN.n167 EN.n166 19.4672
R2885 EN.n163 EN.n162 19.4672
R2886 EN.n164 EN.n163 19.4672
R2887 EN.n158 EN.n157 19.4672
R2888 EN.n169 EN.n168 19.4672
R2889 EN.n170 EN.n169 19.4672
R2890 EN.n171 EN.n170 19.4672
R2891 EN.n172 EN.n171 19.4672
R2892 EN.n173 EN.n172 19.4672
R2893 EN.n174 EN.n173 19.4672
R2894 EN.n175 EN.n174 19.4672
R2895 EN.n200 EN.n199 19.4672
R2896 EN.n201 EN.n200 19.4672
R2897 EN.n194 EN.n193 19.4672
R2898 EN.n203 EN.n202 19.4672
R2899 EN.n204 EN.n203 19.4672
R2900 EN.n205 EN.n204 19.4672
R2901 EN.n206 EN.n205 19.4672
R2902 EN.n207 EN.n206 19.4672
R2903 EN.n208 EN.n207 19.4672
R2904 EN.n209 EN.n208 19.4672
R2905 EN.n14 EN.n13 19.4672
R2906 EN.n10 EN.n9 19.4672
R2907 EN.n17 EN.n16 19.4672
R2908 EN.n18 EN.n17 19.4672
R2909 EN.n19 EN.n18 19.4672
R2910 EN.n20 EN.n19 19.4672
R2911 EN.n21 EN.n20 19.4672
R2912 EN.n22 EN.n21 19.4672
R2913 EN.n23 EN.n22 19.4672
R2914 EN.n228 EN.n227 19.4672
R2915 EN.n229 EN.n228 19.4672
R2916 EN.n230 EN.n229 19.4672
R2917 EN.n231 EN.n230 19.4672
R2918 EN.n232 EN.n231 19.4672
R2919 EN.n233 EN.n232 19.4672
R2920 EN.n234 EN.n233 19.4672
R2921 EN.n242 EN.n241 19.4672
R2922 EN.n241 EN.n240 19.4672
R2923 EN.n240 EN.n239 19.4672
R2924 EN.n239 EN.n238 19.4672
R2925 EN.n238 EN.n237 19.4672
R2926 EN.n237 EN.n236 19.4672
R2927 EN.n236 EN.n235 19.4672
R2928 EN.t187 EN.n88 18.9023
R2929 EN.t149 EN.n89 18.9023
R2930 EN.t43 EN.n90 18.9023
R2931 EN.t184 EN.n91 18.9023
R2932 EN.t211 EN.n96 18.9023
R2933 EN.t105 EN.n98 18.9023
R2934 EN.t71 EN.n99 18.9023
R2935 EN.t39 EN.n68 18.9023
R2936 EN.t216 EN.n66 18.9023
R2937 EN.t44 EN.n64 18.9023
R2938 EN.t220 EN.n61 18.9023
R2939 EN.t150 EN.n60 18.9023
R2940 EN.t138 EN.n57 18.9023
R2941 EN.t56 EN.n69 18.9023
R2942 EN.t5 EN.n29 18.9023
R2943 EN.t132 EN.n31 18.9023
R2944 EN.t182 EN.n32 18.9023
R2945 EN.t238 EN.n35 18.9023
R2946 EN.t157 EN.n37 18.9023
R2947 EN.t208 EN.n39 18.9023
R2948 EN.t99 EN.n41 18.9023
R2949 EN.t75 EN.n118 18.9023
R2950 EN.t63 EN.n121 18.9023
R2951 EN.t78 EN.n123 18.9023
R2952 EN.t2 EN.n124 18.9023
R2953 EN.t236 EN.n125 18.9023
R2954 EN.t167 EN.n129 18.9023
R2955 EN.t155 EN.n130 18.9023
R2956 EN.t186 EN.n152 18.9023
R2957 EN.t22 EN.n155 18.9023
R2958 EN.t193 EN.n156 18.9023
R2959 EN.t117 EN.n159 18.9023
R2960 EN.t110 EN.n160 18.9023
R2961 EN.t35 EN.n161 18.9023
R2962 EN.t32 EN.n165 18.9023
R2963 EN.t95 EN.n187 18.9023
R2964 EN.t86 EN.n189 18.9023
R2965 EN.t15 EN.n191 18.9023
R2966 EN.t4 EN.n192 18.9023
R2967 EN.t173 EN.n195 18.9023
R2968 EN.t103 EN.n197 18.9023
R2969 EN.t176 EN.n198 18.9023
R2970 EN.t30 EN.n0 18.9023
R2971 EN.t205 EN.n3 18.9023
R2972 EN.t131 EN.n5 18.9023
R2973 EN.t120 EN.n7 18.9023
R2974 EN.t55 EN.n8 18.9023
R2975 EN.t124 EN.n11 18.9023
R2976 EN.t61 EN.n12 18.9023
R2977 EN.n220 EN.t88 18.9023
R2978 EN.n221 EN.t83 18.9023
R2979 EN.n222 EN.t9 18.9023
R2980 EN.n223 EN.t237 18.9023
R2981 EN.n224 EN.t163 18.9023
R2982 EN.n225 EN.t94 18.9023
R2983 EN.n219 EN.t153 18.9023
R2984 EN EN.n244 17.6496
R2985 EN.n218 EN.n25 16.4431
R2986 EN.n54 EN.n53 16.443
R2987 EN.n113 EN.n112 16.4376
R2988 EN.n83 EN.n82 16.4376
R2989 EN.n144 EN.n143 16.4376
R2990 EN.n178 EN.n177 16.4376
R2991 EN.n212 EN.n211 16.4376
R2992 EN.n115 EN.n114 9.32902
R2993 EN.n55 EN.n54 7.81778
R2994 EN.n85 EN.n84 4.59449
R2995 EN.n218 EN.n217 4.33887
R2996 EN.n115 EN 3.32688
R2997 EN.n184 EN.n183 2.81655
R2998 EN.n150 EN.n149 2.81655
R2999 EN.n116 EN.n115 2.55924
R3000 EN.n84 EN.n83 2.25216
R3001 EN.n114 EN.n113 2.25216
R3002 EN.n56 EN.n27 2.24309
R3003 EN.n86 EN.n26 2.24309
R3004 EN.n216 EN.n215 1.1255
R3005 EN.n182 EN.n181 1.1255
R3006 EN.n148 EN.n147 1.1255
R3007 EN.n145 EN.n144 0.897624
R3008 EN.n179 EN.n178 0.897624
R3009 EN.n213 EN.n212 0.897624
R3010 EN.n54 EN 0.0811151
R3011 EN EN.n218 0.0800508
R3012 EN.n26 EN 0.0770183
R3013 EN.n27 EN 0.0770183
R3014 EN.n117 EN 0.0550252
R3015 EN.n151 EN 0.0550252
R3016 EN.n185 EN 0.0550252
R3017 EN.n216 EN.n184 0.0324737
R3018 EN.n217 EN.n216 0.0324737
R3019 EN.n182 EN.n150 0.0324737
R3020 EN.n183 EN.n182 0.0324737
R3021 EN.n148 EN.n116 0.0324737
R3022 EN.n149 EN.n148 0.0324737
R3023 EN.n144 EN.n117 0.0301053
R3024 EN.n147 EN.n146 0.0301053
R3025 EN.n178 EN.n151 0.0301053
R3026 EN.n181 EN.n180 0.0301053
R3027 EN.n212 EN.n185 0.0301053
R3028 EN.n215 EN.n214 0.0301053
R3029 EN.n56 EN.n55 0.0157541
R3030 EN.n86 EN.n85 0.0157541
R3031 EN.n114 EN.n86 0.0152178
R3032 EN.n84 EN.n56 0.0152178
R3033 EN.n215 EN.n213 0.00662734
R3034 EN.n181 EN.n179 0.00662734
R3035 EN.n147 EN.n145 0.00662734
R3036 Transmission_Gate_Layout_15.CLKB.n27 Transmission_Gate_Layout_15.CLKB.t15 54.5477
R3037 Transmission_Gate_Layout_15.CLKB.n27 Transmission_Gate_Layout_15.CLKB.t17 38.3255
R3038 Transmission_Gate_Layout_15.CLKB.n28 Transmission_Gate_Layout_15.CLKB.t24 38.3255
R3039 Transmission_Gate_Layout_15.CLKB.n29 Transmission_Gate_Layout_15.CLKB.t27 38.3255
R3040 Transmission_Gate_Layout_15.CLKB.n30 Transmission_Gate_Layout_15.CLKB.t8 38.3255
R3041 Transmission_Gate_Layout_15.CLKB.n31 Transmission_Gate_Layout_15.CLKB.t14 38.3255
R3042 Transmission_Gate_Layout_15.CLKB.n32 Transmission_Gate_Layout_15.CLKB.t7 38.3255
R3043 Transmission_Gate_Layout_15.CLKB.t11 Transmission_Gate_Layout_15.CLKB.n24 37.9344
R3044 Transmission_Gate_Layout_15.CLKB.t9 Transmission_Gate_Layout_15.CLKB.n23 37.9344
R3045 Transmission_Gate_Layout_15.CLKB.t10 Transmission_Gate_Layout_15.CLKB.n20 37.9344
R3046 Transmission_Gate_Layout_15.CLKB.t16 Transmission_Gate_Layout_15.CLKB.n17 37.9344
R3047 Transmission_Gate_Layout_15.CLKB.t19 Transmission_Gate_Layout_15.CLKB.n14 37.9344
R3048 Transmission_Gate_Layout_15.CLKB.t26 Transmission_Gate_Layout_15.CLKB.n11 37.9344
R3049 Transmission_Gate_Layout_15.CLKB.t6 Transmission_Gate_Layout_15.CLKB.n8 37.9344
R3050 Transmission_Gate_Layout_15.CLKB.t25 Transmission_Gate_Layout_15.CLKB.n5 37.9344
R3051 Transmission_Gate_Layout_15.CLKB.n25 Transmission_Gate_Layout_15.CLKB.t11 37.5434
R3052 Transmission_Gate_Layout_15.CLKB.n26 Transmission_Gate_Layout_15.CLKB.t9 37.5434
R3053 Transmission_Gate_Layout_15.CLKB.n21 Transmission_Gate_Layout_15.CLKB.t10 37.5434
R3054 Transmission_Gate_Layout_15.CLKB.n18 Transmission_Gate_Layout_15.CLKB.t16 37.5434
R3055 Transmission_Gate_Layout_15.CLKB.n15 Transmission_Gate_Layout_15.CLKB.t19 37.5434
R3056 Transmission_Gate_Layout_15.CLKB.n12 Transmission_Gate_Layout_15.CLKB.t26 37.5434
R3057 Transmission_Gate_Layout_15.CLKB.n9 Transmission_Gate_Layout_15.CLKB.t6 37.5434
R3058 Transmission_Gate_Layout_15.CLKB.n6 Transmission_Gate_Layout_15.CLKB.t25 37.5434
R3059 Transmission_Gate_Layout_15.CLKB.n25 Transmission_Gate_Layout_15.CLKB.t18 37.413
R3060 Transmission_Gate_Layout_15.CLKB.t17 Transmission_Gate_Layout_15.CLKB.n21 37.413
R3061 Transmission_Gate_Layout_15.CLKB.t24 Transmission_Gate_Layout_15.CLKB.n18 37.413
R3062 Transmission_Gate_Layout_15.CLKB.t27 Transmission_Gate_Layout_15.CLKB.n15 37.413
R3063 Transmission_Gate_Layout_15.CLKB.t8 Transmission_Gate_Layout_15.CLKB.n12 37.413
R3064 Transmission_Gate_Layout_15.CLKB.t14 Transmission_Gate_Layout_15.CLKB.n9 37.413
R3065 Transmission_Gate_Layout_15.CLKB.t7 Transmission_Gate_Layout_15.CLKB.n6 37.413
R3066 Transmission_Gate_Layout_15.CLKB.t15 Transmission_Gate_Layout_15.CLKB.n26 37.413
R3067 Transmission_Gate_Layout_15.CLKB.n24 Transmission_Gate_Layout_15.CLKB.t23 37.0219
R3068 Transmission_Gate_Layout_15.CLKB.n23 Transmission_Gate_Layout_15.CLKB.t21 37.0219
R3069 Transmission_Gate_Layout_15.CLKB.n20 Transmission_Gate_Layout_15.CLKB.t22 37.0219
R3070 Transmission_Gate_Layout_15.CLKB.n17 Transmission_Gate_Layout_15.CLKB.t28 37.0219
R3071 Transmission_Gate_Layout_15.CLKB.n14 Transmission_Gate_Layout_15.CLKB.t29 37.0219
R3072 Transmission_Gate_Layout_15.CLKB.n11 Transmission_Gate_Layout_15.CLKB.t13 37.0219
R3073 Transmission_Gate_Layout_15.CLKB.n5 Transmission_Gate_Layout_15.CLKB.t12 37.0219
R3074 Transmission_Gate_Layout_15.CLKB.n8 Transmission_Gate_Layout_15.CLKB.t20 37.0219
R3075 Transmission_Gate_Layout_15.CLKB.t21 Transmission_Gate_Layout_15.CLKB.n22 35.1969
R3076 Transmission_Gate_Layout_15.CLKB.t22 Transmission_Gate_Layout_15.CLKB.n19 35.1969
R3077 Transmission_Gate_Layout_15.CLKB.t28 Transmission_Gate_Layout_15.CLKB.n16 35.1969
R3078 Transmission_Gate_Layout_15.CLKB.t29 Transmission_Gate_Layout_15.CLKB.n13 35.1969
R3079 Transmission_Gate_Layout_15.CLKB.t13 Transmission_Gate_Layout_15.CLKB.n10 35.1969
R3080 Transmission_Gate_Layout_15.CLKB.t20 Transmission_Gate_Layout_15.CLKB.n7 35.1969
R3081 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_15.CLKB.n32 26.6826
R3082 Transmission_Gate_Layout_15.CLKB.n26 Transmission_Gate_Layout_15.CLKB.n25 19.148
R3083 Transmission_Gate_Layout_15.CLKB.n28 Transmission_Gate_Layout_15.CLKB.n27 16.2227
R3084 Transmission_Gate_Layout_15.CLKB.n29 Transmission_Gate_Layout_15.CLKB.n28 16.2227
R3085 Transmission_Gate_Layout_15.CLKB.n30 Transmission_Gate_Layout_15.CLKB.n29 16.2227
R3086 Transmission_Gate_Layout_15.CLKB.n31 Transmission_Gate_Layout_15.CLKB.n30 16.2227
R3087 Transmission_Gate_Layout_15.CLKB.n32 Transmission_Gate_Layout_15.CLKB.n31 16.2227
R3088 Transmission_Gate_Layout_15.CLKB.n2 Transmission_Gate_Layout_15.CLKB.n0 5.21612
R3089 Transmission_Gate_Layout_15.CLKB.n36 Transmission_Gate_Layout_15.CLKB.n35 4.57285
R3090 Transmission_Gate_Layout_15.CLKB.n4 Transmission_Gate_Layout_15.CLKB.n3 4.4609
R3091 Transmission_Gate_Layout_15.CLKB.n2 Transmission_Gate_Layout_15.CLKB.n1 4.4609
R3092 Transmission_Gate_Layout_15.CLKB.n37 Transmission_Gate_Layout_15.CLKB.n33 3.3285
R3093 Transmission_Gate_Layout_15.CLKB.n36 Transmission_Gate_Layout_15.CLKB.n34 3.3285
R3094 Transmission_Gate_Layout_15.CLKB.n37 Transmission_Gate_Layout_15.CLKB.n36 1.24485
R3095 Transmission_Gate_Layout_15.CLKB.n4 Transmission_Gate_Layout_15.CLKB.n2 0.755717
R3096 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_15.CLKB.n37 0.750969
R3097 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_15.CLKB.n4 0.510317
R3098 Transmission_Gate_Layout_7.CLKB.n27 Transmission_Gate_Layout_7.CLKB.t19 54.5477
R3099 Transmission_Gate_Layout_7.CLKB.n27 Transmission_Gate_Layout_7.CLKB.t25 38.3255
R3100 Transmission_Gate_Layout_7.CLKB.n28 Transmission_Gate_Layout_7.CLKB.t27 38.3255
R3101 Transmission_Gate_Layout_7.CLKB.n29 Transmission_Gate_Layout_7.CLKB.t10 38.3255
R3102 Transmission_Gate_Layout_7.CLKB.n30 Transmission_Gate_Layout_7.CLKB.t12 38.3255
R3103 Transmission_Gate_Layout_7.CLKB.n32 Transmission_Gate_Layout_7.CLKB.t23 38.3255
R3104 Transmission_Gate_Layout_7.CLKB.n31 Transmission_Gate_Layout_7.CLKB.t18 38.3255
R3105 Transmission_Gate_Layout_7.CLKB.t22 Transmission_Gate_Layout_7.CLKB.n24 37.9344
R3106 Transmission_Gate_Layout_7.CLKB.t6 Transmission_Gate_Layout_7.CLKB.n23 37.9344
R3107 Transmission_Gate_Layout_7.CLKB.t11 Transmission_Gate_Layout_7.CLKB.n20 37.9344
R3108 Transmission_Gate_Layout_7.CLKB.t13 Transmission_Gate_Layout_7.CLKB.n17 37.9344
R3109 Transmission_Gate_Layout_7.CLKB.t20 Transmission_Gate_Layout_7.CLKB.n14 37.9344
R3110 Transmission_Gate_Layout_7.CLKB.t21 Transmission_Gate_Layout_7.CLKB.n11 37.9344
R3111 Transmission_Gate_Layout_7.CLKB.t28 Transmission_Gate_Layout_7.CLKB.n8 37.9344
R3112 Transmission_Gate_Layout_7.CLKB.t8 Transmission_Gate_Layout_7.CLKB.n5 37.9344
R3113 Transmission_Gate_Layout_7.CLKB.n25 Transmission_Gate_Layout_7.CLKB.t22 37.5434
R3114 Transmission_Gate_Layout_7.CLKB.n26 Transmission_Gate_Layout_7.CLKB.t6 37.5434
R3115 Transmission_Gate_Layout_7.CLKB.n21 Transmission_Gate_Layout_7.CLKB.t11 37.5434
R3116 Transmission_Gate_Layout_7.CLKB.n18 Transmission_Gate_Layout_7.CLKB.t13 37.5434
R3117 Transmission_Gate_Layout_7.CLKB.n15 Transmission_Gate_Layout_7.CLKB.t20 37.5434
R3118 Transmission_Gate_Layout_7.CLKB.n12 Transmission_Gate_Layout_7.CLKB.t21 37.5434
R3119 Transmission_Gate_Layout_7.CLKB.n9 Transmission_Gate_Layout_7.CLKB.t28 37.5434
R3120 Transmission_Gate_Layout_7.CLKB.n6 Transmission_Gate_Layout_7.CLKB.t8 37.5434
R3121 Transmission_Gate_Layout_7.CLKB.n25 Transmission_Gate_Layout_7.CLKB.t14 37.413
R3122 Transmission_Gate_Layout_7.CLKB.t19 Transmission_Gate_Layout_7.CLKB.n26 37.413
R3123 Transmission_Gate_Layout_7.CLKB.t25 Transmission_Gate_Layout_7.CLKB.n21 37.413
R3124 Transmission_Gate_Layout_7.CLKB.t27 Transmission_Gate_Layout_7.CLKB.n18 37.413
R3125 Transmission_Gate_Layout_7.CLKB.t10 Transmission_Gate_Layout_7.CLKB.n15 37.413
R3126 Transmission_Gate_Layout_7.CLKB.t12 Transmission_Gate_Layout_7.CLKB.n12 37.413
R3127 Transmission_Gate_Layout_7.CLKB.t23 Transmission_Gate_Layout_7.CLKB.n6 37.413
R3128 Transmission_Gate_Layout_7.CLKB.t18 Transmission_Gate_Layout_7.CLKB.n9 37.413
R3129 Transmission_Gate_Layout_7.CLKB.n5 Transmission_Gate_Layout_7.CLKB.t15 37.0219
R3130 Transmission_Gate_Layout_7.CLKB.n11 Transmission_Gate_Layout_7.CLKB.t26 37.0219
R3131 Transmission_Gate_Layout_7.CLKB.n14 Transmission_Gate_Layout_7.CLKB.t24 37.0219
R3132 Transmission_Gate_Layout_7.CLKB.n17 Transmission_Gate_Layout_7.CLKB.t17 37.0219
R3133 Transmission_Gate_Layout_7.CLKB.n20 Transmission_Gate_Layout_7.CLKB.t16 37.0219
R3134 Transmission_Gate_Layout_7.CLKB.n23 Transmission_Gate_Layout_7.CLKB.t9 37.0219
R3135 Transmission_Gate_Layout_7.CLKB.n24 Transmission_Gate_Layout_7.CLKB.t29 37.0219
R3136 Transmission_Gate_Layout_7.CLKB.n8 Transmission_Gate_Layout_7.CLKB.t7 37.0219
R3137 Transmission_Gate_Layout_7.CLKB.t26 Transmission_Gate_Layout_7.CLKB.n10 35.1969
R3138 Transmission_Gate_Layout_7.CLKB.t24 Transmission_Gate_Layout_7.CLKB.n13 35.1969
R3139 Transmission_Gate_Layout_7.CLKB.t17 Transmission_Gate_Layout_7.CLKB.n16 35.1969
R3140 Transmission_Gate_Layout_7.CLKB.t16 Transmission_Gate_Layout_7.CLKB.n19 35.1969
R3141 Transmission_Gate_Layout_7.CLKB.t9 Transmission_Gate_Layout_7.CLKB.n22 35.1969
R3142 Transmission_Gate_Layout_7.CLKB.t7 Transmission_Gate_Layout_7.CLKB.n7 35.1969
R3143 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_7.CLKB.n32 26.6826
R3144 Transmission_Gate_Layout_7.CLKB.n26 Transmission_Gate_Layout_7.CLKB.n25 19.148
R3145 Transmission_Gate_Layout_7.CLKB.n28 Transmission_Gate_Layout_7.CLKB.n27 16.2227
R3146 Transmission_Gate_Layout_7.CLKB.n29 Transmission_Gate_Layout_7.CLKB.n28 16.2227
R3147 Transmission_Gate_Layout_7.CLKB.n30 Transmission_Gate_Layout_7.CLKB.n29 16.2227
R3148 Transmission_Gate_Layout_7.CLKB.n31 Transmission_Gate_Layout_7.CLKB.n30 16.2227
R3149 Transmission_Gate_Layout_7.CLKB.n32 Transmission_Gate_Layout_7.CLKB.n31 16.2227
R3150 Transmission_Gate_Layout_7.CLKB.n35 Transmission_Gate_Layout_7.CLKB.n34 5.21612
R3151 Transmission_Gate_Layout_7.CLKB.n2 Transmission_Gate_Layout_7.CLKB.n0 4.57285
R3152 Transmission_Gate_Layout_7.CLKB.n35 Transmission_Gate_Layout_7.CLKB.n33 4.4609
R3153 Transmission_Gate_Layout_7.CLKB.n37 Transmission_Gate_Layout_7.CLKB.n36 4.4609
R3154 Transmission_Gate_Layout_7.CLKB.n2 Transmission_Gate_Layout_7.CLKB.n1 3.3285
R3155 Transmission_Gate_Layout_7.CLKB.n4 Transmission_Gate_Layout_7.CLKB.n3 3.3285
R3156 Transmission_Gate_Layout_7.CLKB.n4 Transmission_Gate_Layout_7.CLKB.n2 1.24485
R3157 Transmission_Gate_Layout_7.CLKB.n37 Transmission_Gate_Layout_7.CLKB.n35 0.755717
R3158 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_7.CLKB.n4 0.750969
R3159 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_7.CLKB.n37 0.510317
R3160 VDD.n580 VDD.n579 111.675
R3161 VDD.n579 VDD.t176 105.912
R3162 VDD.n67 VDD.t238 100.427
R3163 VDD.n86 VDD.t147 91.8808
R3164 VDD.n110 VDD.t69 91.8808
R3165 VDD.n895 VDD.t168 91.8808
R3166 VDD.n767 VDD.t129 81.4337
R3167 VDD.n767 VDD.t207 81.4337
R3168 VDD.n660 VDD.t1 81.4337
R3169 VDD.n660 VDD.t67 81.4337
R3170 VDD.n798 VDD.t200 74.01
R3171 VDD.n846 VDD.t217 71.0665
R3172 VDD.n558 VDD.t299 71.0665
R3173 VDD.n576 VDD.t163 71.0665
R3174 VDD.n552 VDD.n191 59.7182
R3175 VDD.n698 VDD.t149 49.2667
R3176 VDD.n773 VDD.t48 44.0257
R3177 VDD.n791 VDD.t141 44.0257
R3178 VDD.n684 VDD.t107 43.0365
R3179 VDD.n666 VDD.t28 40.2304
R3180 VDD.n806 VDD.t203 23.6892
R3181 VDD.n565 VDD.t298 23.6892
R3182 VDD.n569 VDD.t166 23.6892
R3183 VDD.n191 VDD.t81 21.716
R3184 VDD.n993 VDD.t214 20.4814
R3185 VDD.n952 VDD.t93 20.4814
R3186 VDD.n937 VDD.t18 20.4814
R3187 VDD.n835 VDD.t14 20.4814
R3188 VDD.n984 VDD.t95 17.8099
R3189 VDD.n967 VDD.t92 16.029
R3190 VDD.n880 VDD.t17 16.029
R3191 VDD.n780 VDD.t50 14.6756
R3192 VDD.n784 VDD.t139 14.6756
R3193 VDD.n301 VDD.t155 14.6391
R3194 VDD.n356 VDD.t291 14.6391
R3195 VDD.n468 VDD.t244 14.6391
R3196 VDD.n523 VDD.t104 14.6391
R3197 VDD.n673 VDD.t27 13.4105
R3198 VDD.n677 VDD.t110 13.4105
R3199 VDD.n970 VDD.t96 13.3576
R3200 VDD.n883 VDD.t12 13.3576
R3201 VDD.n981 VDD.t91 11.5766
R3202 VDD.n864 VDD.t16 11.5766
R3203 VDD.n152 VDD.t13 10.6862
R3204 VDD.n14 VDD.t258 10.522
R3205 VDD.n1233 VDD.t44 10.522
R3206 VDD.n1217 VDD.t185 10.522
R3207 VDD.n1176 VDD.t55 10.522
R3208 VDD.n1161 VDD.t66 10.522
R3209 VDD.n1120 VDD.t24 10.522
R3210 VDD.n1103 VDD.t19 10.522
R3211 VDD.n1062 VDD.t77 10.522
R3212 VDD.n1047 VDD.t144 10.522
R3213 VDD.n1006 VDD.t180 10.522
R3214 VDD.n282 VDD.t161 10.522
R3215 VDD.n320 VDD.t131 10.522
R3216 VDD.n337 VDD.t182 10.522
R3217 VDD.n375 VDD.t113 10.522
R3218 VDD.n391 VDD.t36 10.522
R3219 VDD.n432 VDD.t122 10.522
R3220 VDD.n449 VDD.t227 10.522
R3221 VDD.n487 VDD.t85 10.522
R3222 VDD.n504 VDD.t99 10.522
R3223 VDD.n542 VDD.t178 10.522
R3224 VDD.n1057 VDD.n1055 10.5005
R3225 VDD.n23 VDD.t46 9.14963
R3226 VDD.n1208 VDD.t10 9.14963
R3227 VDD.n1129 VDD.t63 9.14963
R3228 VDD.n1094 VDD.t72 9.14963
R3229 VDD.n1015 VDD.t162 9.14963
R3230 VDD.n423 VDD.t34 9.14963
R3231 VDD.n955 VDD.t94 8.90522
R3232 VDD.n68 VDD.n66 8.25278
R3233 VDD.n1248 VDD.t0 8.23472
R3234 VDD.n1191 VDD.t52 8.23472
R3235 VDD.n1146 VDD.t60 8.23472
R3236 VDD.n1077 VDD.t78 8.23472
R3237 VDD.n1032 VDD.t8 8.23472
R3238 VDD.n297 VDD.t158 8.23472
R3239 VDD.n305 VDD.t132 8.23472
R3240 VDD.n352 VDD.t292 8.23472
R3241 VDD.n360 VDD.t118 8.23472
R3242 VDD.n406 VDD.t29 8.23472
R3243 VDD.n464 VDD.t243 8.23472
R3244 VDD.n472 VDD.t84 8.23472
R3245 VDD.n519 VDD.t101 8.23472
R3246 VDD.n527 VDD.t251 8.23472
R3247 VDD.n1203 VDD.n1201 8.2255
R3248 VDD.n1201 VDD.n1199 8.2255
R3249 VDD.n1141 VDD.n1139 8.2255
R3250 VDD.n1139 VDD.n1137 8.2255
R3251 VDD.n1089 VDD.n1087 8.2255
R3252 VDD.n1087 VDD.n1085 8.2255
R3253 VDD.n1027 VDD.n1025 8.2255
R3254 VDD.n1025 VDD.n1023 8.2255
R3255 VDD.n979 VDD.n977 8.2255
R3256 VDD.n977 VDD.n975 8.2255
R3257 VDD.n87 VDD.n85 8.2255
R3258 VDD.n89 VDD.n87 8.2255
R3259 VDD.n111 VDD.n109 8.2255
R3260 VDD.n113 VDD.n111 8.2255
R3261 VDD.n898 VDD.n896 8.2255
R3262 VDD.n809 VDD.n807 8.2255
R3263 VDD.n699 VDD.n697 8.2255
R3264 VDD.n783 VDD.n781 8.2255
R3265 VDD.n785 VDD.n783 8.2255
R3266 VDD.n676 VDD.n674 8.2255
R3267 VDD.n678 VDD.n676 8.2255
R3268 VDD.n298 VDD.n272 8.2255
R3269 VDD.n302 VDD.n272 8.2255
R3270 VDD.n304 VDD.n302 8.2255
R3271 VDD.n306 VDD.n304 8.2255
R3272 VDD.n353 VDD.n263 8.2255
R3273 VDD.n357 VDD.n263 8.2255
R3274 VDD.n359 VDD.n357 8.2255
R3275 VDD.n361 VDD.n359 8.2255
R3276 VDD.n416 VDD.n414 8.2255
R3277 VDD.n418 VDD.n416 8.2255
R3278 VDD.n465 VDD.n250 8.2255
R3279 VDD.n469 VDD.n250 8.2255
R3280 VDD.n471 VDD.n469 8.2255
R3281 VDD.n473 VDD.n471 8.2255
R3282 VDD.n520 VDD.n241 8.2255
R3283 VDD.n524 VDD.n241 8.2255
R3284 VDD.n526 VDD.n524 8.2255
R3285 VDD.n528 VDD.n526 8.2255
R3286 VDD.n568 VDD.n566 8.2255
R3287 VDD.n570 VDD.n568 8.2255
R3288 VDD.t129 VDD.t145 7.96286
R3289 VDD.t207 VDD.t230 7.96286
R3290 VDD.t1 VDD.t126 7.96286
R3291 VDD.t67 VDD.t124 7.96286
R3292 VDD.t81 VDD.t234 7.96286
R3293 VDD.n872 VDD.n870 7.613
R3294 VDD.n811 VDD.n809 7.3505
R3295 VDD.t154 VDD.t136 7.3198
R3296 VDD.t134 VDD.t159 7.3198
R3297 VDD.t295 VDD.t117 7.3198
R3298 VDD.t115 VDD.t294 7.3198
R3299 VDD.t245 VDD.t89 7.3198
R3300 VDD.t87 VDD.t242 7.3198
R3301 VDD.t103 VDD.t253 7.3198
R3302 VDD.t252 VDD.t105 7.3198
R3303 VDD.n744 VDD.t233 7.06752
R3304 VDD.n744 VDD.t232 7.06752
R3305 VDD.n726 VDD.t130 7.06752
R3306 VDD.n726 VDD.t237 7.06752
R3307 VDD.n709 VDD.t247 7.06752
R3308 VDD.n709 VDD.t208 7.06752
R3309 VDD.n637 VDD.t206 7.06752
R3310 VDD.n637 VDD.t128 7.06752
R3311 VDD.n619 VDD.t236 7.06752
R3312 VDD.n619 VDD.t170 7.06752
R3313 VDD.n602 VDD.t2 7.06752
R3314 VDD.n602 VDD.t68 7.06752
R3315 VDD.n178 VDD.t172 7.06752
R3316 VDD.n186 VDD.t82 7.06752
R3317 VDD.n181 VDD.t112 7.06752
R3318 VDD.n94 VDD.t148 7.06752
R3319 VDD.n118 VDD.t70 7.06752
R3320 VDD.n169 VDD.t169 7.06752
R3321 VDD.n1251 VDD.t45 6.86235
R3322 VDD.n1194 VDD.t9 6.86235
R3323 VDD.n1143 VDD.t65 6.86235
R3324 VDD.n1080 VDD.t71 6.86235
R3325 VDD.n1029 VDD.t3 6.86235
R3326 VDD.n303 VDD.t135 6.86235
R3327 VDD.n358 VDD.t116 6.86235
R3328 VDD.n409 VDD.t31 6.86235
R3329 VDD.n470 VDD.t90 6.86235
R3330 VDD.n525 VDD.t249 6.86235
R3331 VDD.n810 VDD.t222 6.76869
R3332 VDD.n812 VDD.n811 6.3005
R3333 VDD.n811 VDD.n810 6.3005
R3334 VDD.n165 VDD.n164 6.3005
R3335 VDD.n164 VDD.n163 6.3005
R3336 VDD.n134 VDD.n133 6.3005
R3337 VDD.n133 VDD.n132 6.3005
R3338 VDD.n128 VDD.n127 6.3005
R3339 VDD.n127 VDD.n126 6.3005
R3340 VDD.n137 VDD.n136 6.3005
R3341 VDD.n815 VDD.n814 6.3005
R3342 VDD.n854 VDD.n853 6.3005
R3343 VDD.n853 VDD.n852 6.3005
R3344 VDD.n851 VDD.n850 6.3005
R3345 VDD.n850 VDD.n849 6.3005
R3346 VDD.n147 VDD.n146 6.3005
R3347 VDD.n125 VDD.n124 6.3005
R3348 VDD.n124 VDD.n123 6.3005
R3349 VDD.n154 VDD.n153 6.3005
R3350 VDD.n153 VDD.n152 6.3005
R3351 VDD.n910 VDD.n909 6.3005
R3352 VDD.n874 VDD 6.3005
R3353 VDD.n874 VDD.n873 6.3005
R3354 VDD.n157 VDD.n156 6.3005
R3355 VDD.n872 VDD.n871 6.3005
R3356 VDD.n917 VDD.n916 6.3005
R3357 VDD.n916 VDD.n915 6.3005
R3358 VDD.n929 VDD.n928 6.3005
R3359 VDD.n936 VDD.n935 6.3005
R3360 VDD.n935 VDD.n934 6.3005
R3361 VDD.n26 VDD.t43 5.94744
R3362 VDD.n1205 VDD.t53 5.94744
R3363 VDD.n1132 VDD.t59 5.94744
R3364 VDD.n1091 VDD.t74 5.94744
R3365 VDD.n1018 VDD.t5 5.94744
R3366 VDD.n294 VDD.t138 5.94744
R3367 VDD.n308 VDD.t157 5.94744
R3368 VDD.n349 VDD.t119 5.94744
R3369 VDD.n363 VDD.t297 5.94744
R3370 VDD.n420 VDD.t32 5.94744
R3371 VDD.n461 VDD.t86 5.94744
R3372 VDD.n475 VDD.t246 5.94744
R3373 VDD.n516 VDD.t171 5.94744
R3374 VDD.n530 VDD.t100 5.94744
R3375 VDD.n760 VDD.n759 4.9354
R3376 VDD.n742 VDD.n741 4.9354
R3377 VDD.n724 VDD.n723 4.9354
R3378 VDD.n653 VDD.n652 4.9354
R3379 VDD.n635 VDD.n634 4.9354
R3380 VDD.n617 VDD.n616 4.9354
R3381 VDD.n554 VDD.n553 4.9354
R3382 VDD.n190 VDD.n189 4.9354
R3383 VDD.n185 VDD.n184 4.9354
R3384 VDD.n180 VDD.n179 4.9354
R3385 VDD.n590 VDD.n582 4.9354
R3386 VDD.n206 VDD.n205 4.93487
R3387 VDD.n219 VDD.n218 4.93487
R3388 VDD.n232 VDD.n231 4.93487
R3389 VDD.n551 VDD.n550 4.93487
R3390 VDD.n769 VDD.n768 4.93474
R3391 VDD.n729 VDD.n725 4.93474
R3392 VDD.n747 VDD.n743 4.93474
R3393 VDD.n762 VDD.n761 4.93474
R3394 VDD.n662 VDD.n661 4.93474
R3395 VDD.n622 VDD.n618 4.93474
R3396 VDD.n640 VDD.n636 4.93474
R3397 VDD.n655 VDD.n654 4.93474
R3398 VDD.n763 VDD.t146 4.7942
R3399 VDD.n763 VDD.t231 4.7942
R3400 VDD.n694 VDD.t150 4.7942
R3401 VDD.n694 VDD.t205 4.7942
R3402 VDD.n656 VDD.t127 4.7942
R3403 VDD.n656 VDD.t125 4.7942
R3404 VDD.n583 VDD.t177 4.7942
R3405 VDD.n233 VDD.t235 4.7942
R3406 VDD.n70 VDD.t239 4.7942
R3407 VDD.n1236 VDD.t41 4.57507
R3408 VDD.n1179 VDD.t11 4.57507
R3409 VDD.n1158 VDD.t62 4.57507
R3410 VDD.n1065 VDD.t73 4.57507
R3411 VDD.n1044 VDD.t7 4.57507
R3412 VDD.n285 VDD.t156 4.57507
R3413 VDD.n317 VDD.t137 4.57507
R3414 VDD.n340 VDD.t296 4.57507
R3415 VDD.n372 VDD.t120 4.57507
R3416 VDD.n394 VDD.t30 4.57507
R3417 VDD.n452 VDD.t240 4.57507
R3418 VDD.n484 VDD.t83 4.57507
R3419 VDD.n507 VDD.t106 4.57507
R3420 VDD.n539 VDD.t250 4.57507
R3421 VDD.n269 VDD.t272 4.57285
R3422 VDD.n260 VDD.t290 4.57285
R3423 VDD.n256 VDD.t271 4.57285
R3424 VDD.n258 VDD.t123 4.57285
R3425 VDD.n247 VDD.t287 4.57285
R3426 VDD.n244 VDD.n242 4.57285
R3427 VDD.n238 VDD.t179 4.57285
R3428 VDD.n254 VDD.n253 4.57285
R3429 VDD.n267 VDD.n266 4.57285
R3430 VDD.n276 VDD.n275 4.57285
R3431 VDD.n2 VDD.n0 4.57285
R3432 VDD.n8 VDD.n7 4.57285
R3433 VDD.n34 VDD.n32 4.57285
R3434 VDD.n40 VDD.n39 4.57285
R3435 VDD.n42 VDD.t309 4.57285
R3436 VDD.n44 VDD.t39 4.57285
R3437 VDD.n48 VDD.n46 4.57285
R3438 VDD.n54 VDD.n53 4.57285
R3439 VDD.n56 VDD.t195 4.57285
R3440 VDD.n58 VDD.t211 4.57285
R3441 VDD.n828 VDD.t51 4.57285
R3442 VDD.n63 VDD.n62 4.57285
R3443 VDD.n857 VDD.n856 4.5005
R3444 VDD.n856 VDD.n855 4.5005
R3445 VDD.n150 VDD.n149 4.5005
R3446 VDD.n149 VDD.n148 4.5005
R3447 VDD.n122 VDD.n121 4.5005
R3448 VDD.n121 VDD.n120 4.5005
R3449 VDD.n140 VDD.n139 4.5005
R3450 VDD.n139 VDD.n138 4.5005
R3451 VDD.n818 VDD.n817 4.5005
R3452 VDD.n817 VDD.n816 4.5005
R3453 VDD.n160 VDD.n159 4.5005
R3454 VDD.n159 VDD.n158 4.5005
R3455 VDD.n877 VDD.n876 4.5005
R3456 VDD.n876 VDD.n875 4.5005
R3457 VDD.n913 VDD.n912 4.5005
R3458 VDD.n912 VDD.n911 4.5005
R3459 VDD.n932 VDD.n931 4.5005
R3460 VDD.n931 VDD.n930 4.5005
R3461 VDD.n930 VDD.t56 4.45286
R3462 VDD.n961 VDD.t98 3.56239
R3463 VDD.n918 VDD.t47 3.56239
R3464 VDD.n797 VDD.n796 3.42899
R3465 VDD.n270 VDD.t268 3.3285
R3466 VDD.n269 VDD.t283 3.3285
R3467 VDD.n261 VDD.t286 3.3285
R3468 VDD.n260 VDD.t264 3.3285
R3469 VDD.n259 VDD.t306 3.3285
R3470 VDD.n258 VDD.t300 3.3285
R3471 VDD.n257 VDD.t267 3.3285
R3472 VDD.n256 VDD.t280 3.3285
R3473 VDD.n248 VDD.t279 3.3285
R3474 VDD.n247 VDD.t261 3.3285
R3475 VDD.n244 VDD.n243 3.3285
R3476 VDD.n246 VDD.n245 3.3285
R3477 VDD.n239 VDD.t190 3.3285
R3478 VDD.n238 VDD.t194 3.3285
R3479 VDD.n255 VDD.n251 3.3285
R3480 VDD.n254 VDD.n252 3.3285
R3481 VDD.n268 VDD.n264 3.3285
R3482 VDD.n267 VDD.n265 3.3285
R3483 VDD.n277 VDD.n273 3.3285
R3484 VDD.n276 VDD.n274 3.3285
R3485 VDD.n9 VDD.n5 3.3285
R3486 VDD.n8 VDD.n6 3.3285
R3487 VDD.n4 VDD.n3 3.3285
R3488 VDD.n2 VDD.n1 3.3285
R3489 VDD.n41 VDD.n37 3.3285
R3490 VDD.n40 VDD.n38 3.3285
R3491 VDD.n36 VDD.n35 3.3285
R3492 VDD.n34 VDD.n33 3.3285
R3493 VDD.n45 VDD.t25 3.3285
R3494 VDD.n44 VDD.t26 3.3285
R3495 VDD.n43 VDD.t303 3.3285
R3496 VDD.n42 VDD.t121 3.3285
R3497 VDD.n55 VDD.n51 3.3285
R3498 VDD.n54 VDD.n52 3.3285
R3499 VDD.n50 VDD.n49 3.3285
R3500 VDD.n48 VDD.n47 3.3285
R3501 VDD.n59 VDD.t225 3.3285
R3502 VDD.n58 VDD.t226 3.3285
R3503 VDD.n57 VDD.t181 3.3285
R3504 VDD.n56 VDD.t191 3.3285
R3505 VDD.n829 VDD.t15 3.3285
R3506 VDD.n828 VDD.t49 3.3285
R3507 VDD.n64 VDD.n60 3.3285
R3508 VDD.n63 VDD.n61 3.3285
R3509 VDD.n765 VDD.n764 3.1505
R3510 VDD.n758 VDD.n757 3.1505
R3511 VDD.n755 VDD.n754 3.1505
R3512 VDD.n753 VDD.n752 3.1505
R3513 VDD VDD.n751 3.1505
R3514 VDD.n750 VDD.n749 3.1505
R3515 VDD.n746 VDD.n745 3.1505
R3516 VDD.n740 VDD.n739 3.1505
R3517 VDD.n737 VDD.n736 3.1505
R3518 VDD.n735 VDD.n734 3.1505
R3519 VDD VDD.n733 3.1505
R3520 VDD.n732 VDD.n731 3.1505
R3521 VDD.n728 VDD.n727 3.1505
R3522 VDD.n722 VDD.n721 3.1505
R3523 VDD.n719 VDD.n718 3.1505
R3524 VDD.n717 VDD.n716 3.1505
R3525 VDD VDD.n715 3.1505
R3526 VDD.n713 VDD.n712 3.1505
R3527 VDD.n711 VDD.n710 3.1505
R3528 VDD.n772 VDD.n771 3.1505
R3529 VDD.n771 VDD.n770 3.1505
R3530 VDD.n775 VDD.n774 3.1505
R3531 VDD.n774 VDD.n773 3.1505
R3532 VDD.n778 VDD.n777 3.1505
R3533 VDD.n777 VDD.n776 3.1505
R3534 VDD.n781 VDD.n779 3.1505
R3535 VDD.n781 VDD.n780 3.1505
R3536 VDD.n783 VDD 3.1505
R3537 VDD.n783 VDD.n782 3.1505
R3538 VDD.n786 VDD.n785 3.1505
R3539 VDD.n785 VDD.n784 3.1505
R3540 VDD.n790 VDD.n789 3.1505
R3541 VDD.n789 VDD.n788 3.1505
R3542 VDD.n793 VDD.n792 3.1505
R3543 VDD.n792 VDD.n791 3.1505
R3544 VDD.n700 VDD.n699 3.1505
R3545 VDD.n699 VDD.n698 3.1505
R3546 VDD.n697 VDD.n695 3.1505
R3547 VDD.n703 VDD.n702 3.1505
R3548 VDD.n702 VDD.n701 3.1505
R3549 VDD.n658 VDD.n657 3.1505
R3550 VDD.n651 VDD.n650 3.1505
R3551 VDD.n648 VDD.n647 3.1505
R3552 VDD.n646 VDD.n645 3.1505
R3553 VDD VDD.n644 3.1505
R3554 VDD.n643 VDD.n642 3.1505
R3555 VDD.n639 VDD.n638 3.1505
R3556 VDD.n633 VDD.n632 3.1505
R3557 VDD.n630 VDD.n629 3.1505
R3558 VDD.n628 VDD.n627 3.1505
R3559 VDD VDD.n626 3.1505
R3560 VDD.n625 VDD.n624 3.1505
R3561 VDD.n621 VDD.n620 3.1505
R3562 VDD.n615 VDD.n614 3.1505
R3563 VDD.n612 VDD.n611 3.1505
R3564 VDD.n610 VDD.n609 3.1505
R3565 VDD VDD.n608 3.1505
R3566 VDD.n606 VDD.n605 3.1505
R3567 VDD.n604 VDD.n603 3.1505
R3568 VDD.n665 VDD.n664 3.1505
R3569 VDD.n664 VDD.n663 3.1505
R3570 VDD.n668 VDD.n667 3.1505
R3571 VDD.n667 VDD.n666 3.1505
R3572 VDD.n671 VDD.n670 3.1505
R3573 VDD.n670 VDD.n669 3.1505
R3574 VDD.n674 VDD.n672 3.1505
R3575 VDD.n674 VDD.n673 3.1505
R3576 VDD.n676 VDD 3.1505
R3577 VDD.n676 VDD.n675 3.1505
R3578 VDD.n679 VDD.n678 3.1505
R3579 VDD.n678 VDD.n677 3.1505
R3580 VDD.n683 VDD.n682 3.1505
R3581 VDD.n682 VDD.n681 3.1505
R3582 VDD.n686 VDD.n685 3.1505
R3583 VDD.n578 VDD.n577 3.1505
R3584 VDD.n577 VDD.n576 3.1505
R3585 VDD.n204 VDD.n203 3.1505
R3586 VDD.n193 VDD.n192 3.1505
R3587 VDD.n201 VDD.n200 3.1505
R3588 VDD VDD.n199 3.1505
R3589 VDD.n197 VDD.n196 3.1505
R3590 VDD.n195 VDD.n194 3.1505
R3591 VDD.n217 VDD.n216 3.1505
R3592 VDD.n209 VDD.n208 3.1505
R3593 VDD.n214 VDD.n213 3.1505
R3594 VDD VDD.n212 3.1505
R3595 VDD.n211 VDD.n210 3.1505
R3596 VDD.n188 VDD.n187 3.1505
R3597 VDD.n230 VDD.n229 3.1505
R3598 VDD.n222 VDD.n221 3.1505
R3599 VDD.n227 VDD.n226 3.1505
R3600 VDD VDD.n225 3.1505
R3601 VDD.n224 VDD.n223 3.1505
R3602 VDD.n183 VDD.n182 3.1505
R3603 VDD.n237 VDD.n236 3.1505
R3604 VDD.n235 VDD.n234 3.1505
R3605 VDD.n281 VDD.n280 3.1505
R3606 VDD.n284 VDD.n283 3.1505
R3607 VDD.n283 VDD.n282 3.1505
R3608 VDD.n287 VDD.n286 3.1505
R3609 VDD.n286 VDD.n285 3.1505
R3610 VDD.n290 VDD.n289 3.1505
R3611 VDD.n289 VDD.n288 3.1505
R3612 VDD.n293 VDD.n292 3.1505
R3613 VDD.n292 VDD.n291 3.1505
R3614 VDD.n296 VDD.n295 3.1505
R3615 VDD.n295 VDD.n294 3.1505
R3616 VDD.n299 VDD.n298 3.1505
R3617 VDD.n298 VDD.n297 3.1505
R3618 VDD VDD.n272 3.1505
R3619 VDD.n272 VDD.n271 3.1505
R3620 VDD.n302 VDD.n300 3.1505
R3621 VDD.n302 VDD.n301 3.1505
R3622 VDD.n304 VDD 3.1505
R3623 VDD.n304 VDD.n303 3.1505
R3624 VDD.n307 VDD.n306 3.1505
R3625 VDD.n306 VDD.n305 3.1505
R3626 VDD.n310 VDD.n309 3.1505
R3627 VDD.n309 VDD.n308 3.1505
R3628 VDD.n313 VDD.n312 3.1505
R3629 VDD.n312 VDD.n311 3.1505
R3630 VDD.n316 VDD.n315 3.1505
R3631 VDD.n315 VDD.n314 3.1505
R3632 VDD.n319 VDD.n318 3.1505
R3633 VDD.n318 VDD.n317 3.1505
R3634 VDD.n322 VDD.n321 3.1505
R3635 VDD.n321 VDD.n320 3.1505
R3636 VDD.n325 VDD.n324 3.1505
R3637 VDD.n324 VDD.n323 3.1505
R3638 VDD.n329 VDD.n328 3.1505
R3639 VDD.n328 VDD.n327 3.1505
R3640 VDD.n332 VDD.n331 3.1505
R3641 VDD.n331 VDD.n330 3.1505
R3642 VDD.n336 VDD.n335 3.1505
R3643 VDD.n335 VDD.n334 3.1505
R3644 VDD.n339 VDD.n338 3.1505
R3645 VDD.n338 VDD.n337 3.1505
R3646 VDD.n342 VDD.n341 3.1505
R3647 VDD.n341 VDD.n340 3.1505
R3648 VDD.n345 VDD.n344 3.1505
R3649 VDD.n344 VDD.n343 3.1505
R3650 VDD.n348 VDD.n347 3.1505
R3651 VDD.n347 VDD.n346 3.1505
R3652 VDD.n351 VDD.n350 3.1505
R3653 VDD.n350 VDD.n349 3.1505
R3654 VDD.n354 VDD.n353 3.1505
R3655 VDD.n353 VDD.n352 3.1505
R3656 VDD VDD.n263 3.1505
R3657 VDD.n263 VDD.n262 3.1505
R3658 VDD.n357 VDD.n355 3.1505
R3659 VDD.n357 VDD.n356 3.1505
R3660 VDD.n359 VDD 3.1505
R3661 VDD.n359 VDD.n358 3.1505
R3662 VDD.n362 VDD.n361 3.1505
R3663 VDD.n361 VDD.n360 3.1505
R3664 VDD.n365 VDD.n364 3.1505
R3665 VDD.n364 VDD.n363 3.1505
R3666 VDD.n368 VDD.n367 3.1505
R3667 VDD.n367 VDD.n366 3.1505
R3668 VDD.n371 VDD.n370 3.1505
R3669 VDD.n370 VDD.n369 3.1505
R3670 VDD.n374 VDD.n373 3.1505
R3671 VDD.n373 VDD.n372 3.1505
R3672 VDD.n377 VDD.n376 3.1505
R3673 VDD.n376 VDD.n375 3.1505
R3674 VDD.n380 VDD.n379 3.1505
R3675 VDD.n379 VDD.n378 3.1505
R3676 VDD.n384 VDD.n383 3.1505
R3677 VDD.n383 VDD.n382 3.1505
R3678 VDD.n387 VDD.n386 3.1505
R3679 VDD.n386 VDD.n385 3.1505
R3680 VDD.n390 VDD.n389 3.1505
R3681 VDD.n389 VDD.n388 3.1505
R3682 VDD.n393 VDD.n392 3.1505
R3683 VDD.n392 VDD.n391 3.1505
R3684 VDD.n396 VDD.n395 3.1505
R3685 VDD.n395 VDD.n394 3.1505
R3686 VDD.n399 VDD.n398 3.1505
R3687 VDD.n398 VDD.n397 3.1505
R3688 VDD.n402 VDD.n401 3.1505
R3689 VDD.n401 VDD.n400 3.1505
R3690 VDD.n405 VDD.n404 3.1505
R3691 VDD.n404 VDD.n403 3.1505
R3692 VDD.n408 VDD.n407 3.1505
R3693 VDD.n407 VDD.n406 3.1505
R3694 VDD.n411 VDD.n410 3.1505
R3695 VDD.n410 VDD.n409 3.1505
R3696 VDD.n414 VDD.n412 3.1505
R3697 VDD.n414 VDD.n413 3.1505
R3698 VDD.n416 VDD 3.1505
R3699 VDD.n416 VDD.n415 3.1505
R3700 VDD.n419 VDD.n418 3.1505
R3701 VDD.n418 VDD.n417 3.1505
R3702 VDD.n422 VDD.n421 3.1505
R3703 VDD.n421 VDD.n420 3.1505
R3704 VDD.n425 VDD.n424 3.1505
R3705 VDD.n424 VDD.n423 3.1505
R3706 VDD.n428 VDD.n427 3.1505
R3707 VDD.n427 VDD.n426 3.1505
R3708 VDD.n431 VDD.n430 3.1505
R3709 VDD.n430 VDD.n429 3.1505
R3710 VDD.n434 VDD.n433 3.1505
R3711 VDD.n433 VDD.n432 3.1505
R3712 VDD.n437 VDD.n436 3.1505
R3713 VDD.n436 VDD.n435 3.1505
R3714 VDD.n441 VDD.n440 3.1505
R3715 VDD.n440 VDD.n439 3.1505
R3716 VDD.n444 VDD.n443 3.1505
R3717 VDD.n443 VDD.n442 3.1505
R3718 VDD.n448 VDD.n447 3.1505
R3719 VDD.n447 VDD.n446 3.1505
R3720 VDD.n451 VDD.n450 3.1505
R3721 VDD.n450 VDD.n449 3.1505
R3722 VDD.n454 VDD.n453 3.1505
R3723 VDD.n453 VDD.n452 3.1505
R3724 VDD.n457 VDD.n456 3.1505
R3725 VDD.n456 VDD.n455 3.1505
R3726 VDD.n460 VDD.n459 3.1505
R3727 VDD.n459 VDD.n458 3.1505
R3728 VDD.n463 VDD.n462 3.1505
R3729 VDD.n462 VDD.n461 3.1505
R3730 VDD.n466 VDD.n465 3.1505
R3731 VDD.n465 VDD.n464 3.1505
R3732 VDD VDD.n250 3.1505
R3733 VDD.n250 VDD.n249 3.1505
R3734 VDD.n469 VDD.n467 3.1505
R3735 VDD.n469 VDD.n468 3.1505
R3736 VDD.n471 VDD 3.1505
R3737 VDD.n471 VDD.n470 3.1505
R3738 VDD.n474 VDD.n473 3.1505
R3739 VDD.n473 VDD.n472 3.1505
R3740 VDD.n477 VDD.n476 3.1505
R3741 VDD.n476 VDD.n475 3.1505
R3742 VDD.n480 VDD.n479 3.1505
R3743 VDD.n479 VDD.n478 3.1505
R3744 VDD.n483 VDD.n482 3.1505
R3745 VDD.n482 VDD.n481 3.1505
R3746 VDD.n486 VDD.n485 3.1505
R3747 VDD.n485 VDD.n484 3.1505
R3748 VDD.n489 VDD.n488 3.1505
R3749 VDD.n488 VDD.n487 3.1505
R3750 VDD.n492 VDD.n491 3.1505
R3751 VDD.n491 VDD.n490 3.1505
R3752 VDD.n496 VDD.n495 3.1505
R3753 VDD.n495 VDD.n494 3.1505
R3754 VDD.n499 VDD.n498 3.1505
R3755 VDD.n498 VDD.n497 3.1505
R3756 VDD.n503 VDD.n502 3.1505
R3757 VDD.n502 VDD.n501 3.1505
R3758 VDD.n506 VDD.n505 3.1505
R3759 VDD.n505 VDD.n504 3.1505
R3760 VDD.n509 VDD.n508 3.1505
R3761 VDD.n508 VDD.n507 3.1505
R3762 VDD.n512 VDD.n511 3.1505
R3763 VDD.n511 VDD.n510 3.1505
R3764 VDD.n515 VDD.n514 3.1505
R3765 VDD.n514 VDD.n513 3.1505
R3766 VDD.n518 VDD.n517 3.1505
R3767 VDD.n517 VDD.n516 3.1505
R3768 VDD.n521 VDD.n520 3.1505
R3769 VDD.n520 VDD.n519 3.1505
R3770 VDD VDD.n241 3.1505
R3771 VDD.n241 VDD.n240 3.1505
R3772 VDD.n524 VDD.n522 3.1505
R3773 VDD.n524 VDD.n523 3.1505
R3774 VDD.n526 VDD 3.1505
R3775 VDD.n526 VDD.n525 3.1505
R3776 VDD.n529 VDD.n528 3.1505
R3777 VDD.n528 VDD.n527 3.1505
R3778 VDD.n532 VDD.n531 3.1505
R3779 VDD.n531 VDD.n530 3.1505
R3780 VDD.n535 VDD.n534 3.1505
R3781 VDD.n534 VDD.n533 3.1505
R3782 VDD.n538 VDD.n537 3.1505
R3783 VDD.n537 VDD.n536 3.1505
R3784 VDD.n541 VDD.n540 3.1505
R3785 VDD.n540 VDD.n539 3.1505
R3786 VDD.n544 VDD.n543 3.1505
R3787 VDD.n543 VDD.n542 3.1505
R3788 VDD.n547 VDD.n546 3.1505
R3789 VDD.n557 VDD.n556 3.1505
R3790 VDD.n556 VDD.n555 3.1505
R3791 VDD.n560 VDD.n559 3.1505
R3792 VDD.n559 VDD.n558 3.1505
R3793 VDD.n563 VDD.n562 3.1505
R3794 VDD.n562 VDD.n561 3.1505
R3795 VDD.n566 VDD.n564 3.1505
R3796 VDD.n566 VDD.n565 3.1505
R3797 VDD.n568 VDD 3.1505
R3798 VDD.n568 VDD.n567 3.1505
R3799 VDD.n571 VDD.n570 3.1505
R3800 VDD.n570 VDD.n569 3.1505
R3801 VDD.n575 VDD.n574 3.1505
R3802 VDD.n574 VDD.n573 3.1505
R3803 VDD.n589 VDD.n588 3.1505
R3804 VDD.n587 VDD.n586 3.1505
R3805 VDD.n69 VDD.n68 3.1505
R3806 VDD.n68 VDD.n67 3.1505
R3807 VDD.n73 VDD.n72 3.1505
R3808 VDD.n72 VDD.n71 3.1505
R3809 VDD.n76 VDD.n75 3.1505
R3810 VDD.n75 VDD.n74 3.1505
R3811 VDD.n79 VDD.n78 3.1505
R3812 VDD.n78 VDD.n77 3.1505
R3813 VDD.n82 VDD.n81 3.1505
R3814 VDD.n81 VDD.n80 3.1505
R3815 VDD.n85 VDD.n83 3.1505
R3816 VDD.n85 VDD.n84 3.1505
R3817 VDD.n87 VDD 3.1505
R3818 VDD.n87 VDD.n86 3.1505
R3819 VDD.n90 VDD.n89 3.1505
R3820 VDD.n89 VDD.n88 3.1505
R3821 VDD.n93 VDD.n92 3.1505
R3822 VDD.n92 VDD.n91 3.1505
R3823 VDD.n97 VDD.n96 3.1505
R3824 VDD.n96 VDD.n95 3.1505
R3825 VDD.n100 VDD.n99 3.1505
R3826 VDD.n99 VDD.n98 3.1505
R3827 VDD.n103 VDD.n102 3.1505
R3828 VDD.n102 VDD.n101 3.1505
R3829 VDD.n106 VDD.n105 3.1505
R3830 VDD.n105 VDD.n104 3.1505
R3831 VDD.n109 VDD.n107 3.1505
R3832 VDD.n109 VDD.n108 3.1505
R3833 VDD.n111 VDD 3.1505
R3834 VDD.n111 VDD.n110 3.1505
R3835 VDD.n114 VDD.n113 3.1505
R3836 VDD.n113 VDD.n112 3.1505
R3837 VDD.n117 VDD.n116 3.1505
R3838 VDD.n116 VDD.n115 3.1505
R3839 VDD.n848 VDD.n847 3.1505
R3840 VDD.n847 VDD.n846 3.1505
R3841 VDD.n845 VDD.n844 3.1505
R3842 VDD.n844 VDD.n843 3.1505
R3843 VDD.n809 VDD 3.1505
R3844 VDD.n809 VDD.n808 3.1505
R3845 VDD.n807 VDD.n805 3.1505
R3846 VDD.n807 VDD.n806 3.1505
R3847 VDD.n803 VDD.n802 3.1505
R3848 VDD.n802 VDD.n801 3.1505
R3849 VDD.n800 VDD.n799 3.1505
R3850 VDD.n899 VDD.n898 3.1505
R3851 VDD.n898 VDD.n897 3.1505
R3852 VDD.n896 VDD 3.1505
R3853 VDD.n896 VDD.n895 3.1505
R3854 VDD.n168 VDD.n167 3.1505
R3855 VDD.n167 VDD.n166 3.1505
R3856 VDD.n172 VDD.n171 3.1505
R3857 VDD.n171 VDD.n170 3.1505
R3858 VDD.n131 VDD.n130 3.1505
R3859 VDD.n130 VDD.n129 3.1505
R3860 VDD.n902 VDD.n901 3.1505
R3861 VDD.n901 VDD.n900 3.1505
R3862 VDD.n13 VDD.n12 3.1505
R3863 VDD.n16 VDD.n15 3.1505
R3864 VDD.n15 VDD.n14 3.1505
R3865 VDD.n19 VDD.n18 3.1505
R3866 VDD.n18 VDD.n17 3.1505
R3867 VDD.n22 VDD.n21 3.1505
R3868 VDD.n21 VDD.n20 3.1505
R3869 VDD.n25 VDD.n24 3.1505
R3870 VDD.n24 VDD.n23 3.1505
R3871 VDD.n28 VDD.n27 3.1505
R3872 VDD.n27 VDD.n26 3.1505
R3873 VDD.n31 VDD.n30 3.1505
R3874 VDD.n30 VDD.n29 3.1505
R3875 VDD VDD.n1258 3.1505
R3876 VDD.n1258 VDD.n1257 3.1505
R3877 VDD.n1256 VDD.n1255 3.1505
R3878 VDD.n1255 VDD.n1254 3.1505
R3879 VDD.n1253 VDD.n1252 3.1505
R3880 VDD.n1252 VDD.n1251 3.1505
R3881 VDD.n1250 VDD.n1249 3.1505
R3882 VDD.n1249 VDD.n1248 3.1505
R3883 VDD.n1247 VDD.n1246 3.1505
R3884 VDD.n1246 VDD.n1245 3.1505
R3885 VDD.n1244 VDD.n1243 3.1505
R3886 VDD.n1243 VDD.n1242 3.1505
R3887 VDD.n1241 VDD.n1240 3.1505
R3888 VDD.n1240 VDD.n1239 3.1505
R3889 VDD.n1238 VDD.n1237 3.1505
R3890 VDD.n1237 VDD.n1236 3.1505
R3891 VDD.n1235 VDD.n1234 3.1505
R3892 VDD.n1234 VDD.n1233 3.1505
R3893 VDD.n1232 VDD.n1231 3.1505
R3894 VDD.n1231 VDD.n1230 3.1505
R3895 VDD.n1229 VDD.n1228 3.1505
R3896 VDD.n1228 VDD.n1227 3.1505
R3897 VDD.n1226 VDD.n1225 3.1505
R3898 VDD.n1225 VDD.n1224 3.1505
R3899 VDD.n1222 VDD.n1221 3.1505
R3900 VDD.n1221 VDD.n1220 3.1505
R3901 VDD.n1219 VDD.n1218 3.1505
R3902 VDD.n1218 VDD.n1217 3.1505
R3903 VDD.n1216 VDD.n1215 3.1505
R3904 VDD.n1215 VDD.n1214 3.1505
R3905 VDD.n1213 VDD.n1212 3.1505
R3906 VDD.n1212 VDD.n1211 3.1505
R3907 VDD.n1210 VDD.n1209 3.1505
R3908 VDD.n1209 VDD.n1208 3.1505
R3909 VDD.n1207 VDD.n1206 3.1505
R3910 VDD.n1206 VDD.n1205 3.1505
R3911 VDD.n1204 VDD.n1203 3.1505
R3912 VDD.n1203 VDD.n1202 3.1505
R3913 VDD.n1201 VDD 3.1505
R3914 VDD.n1201 VDD.n1200 3.1505
R3915 VDD.n1199 VDD.n1197 3.1505
R3916 VDD.n1199 VDD.n1198 3.1505
R3917 VDD.n1196 VDD.n1195 3.1505
R3918 VDD.n1195 VDD.n1194 3.1505
R3919 VDD.n1193 VDD.n1192 3.1505
R3920 VDD.n1192 VDD.n1191 3.1505
R3921 VDD.n1190 VDD.n1189 3.1505
R3922 VDD.n1189 VDD.n1188 3.1505
R3923 VDD.n1187 VDD.n1186 3.1505
R3924 VDD.n1186 VDD.n1185 3.1505
R3925 VDD.n1184 VDD.n1183 3.1505
R3926 VDD.n1183 VDD.n1182 3.1505
R3927 VDD.n1181 VDD.n1180 3.1505
R3928 VDD.n1180 VDD.n1179 3.1505
R3929 VDD.n1178 VDD.n1177 3.1505
R3930 VDD.n1177 VDD.n1176 3.1505
R3931 VDD.n1175 VDD.n1174 3.1505
R3932 VDD.n1174 VDD.n1173 3.1505
R3933 VDD.n1172 VDD.n1171 3.1505
R3934 VDD.n1171 VDD.n1170 3.1505
R3935 VDD.n1169 VDD.n1168 3.1505
R3936 VDD.n1168 VDD.n1167 3.1505
R3937 VDD.n1166 VDD.n1165 3.1505
R3938 VDD.n1165 VDD.n1164 3.1505
R3939 VDD.n1163 VDD.n1162 3.1505
R3940 VDD.n1162 VDD.n1161 3.1505
R3941 VDD.n1160 VDD.n1159 3.1505
R3942 VDD.n1159 VDD.n1158 3.1505
R3943 VDD.n1157 VDD.n1156 3.1505
R3944 VDD.n1156 VDD.n1155 3.1505
R3945 VDD.n1154 VDD.n1153 3.1505
R3946 VDD.n1153 VDD.n1152 3.1505
R3947 VDD.n1151 VDD.n1150 3.1505
R3948 VDD.n1150 VDD.n1149 3.1505
R3949 VDD.n1148 VDD.n1147 3.1505
R3950 VDD.n1147 VDD.n1146 3.1505
R3951 VDD.n1145 VDD.n1144 3.1505
R3952 VDD.n1144 VDD.n1143 3.1505
R3953 VDD.n1142 VDD.n1141 3.1505
R3954 VDD.n1141 VDD.n1140 3.1505
R3955 VDD.n1139 VDD 3.1505
R3956 VDD.n1139 VDD.n1138 3.1505
R3957 VDD.n1137 VDD.n1135 3.1505
R3958 VDD.n1137 VDD.n1136 3.1505
R3959 VDD.n1134 VDD.n1133 3.1505
R3960 VDD.n1133 VDD.n1132 3.1505
R3961 VDD.n1131 VDD.n1130 3.1505
R3962 VDD.n1130 VDD.n1129 3.1505
R3963 VDD.n1128 VDD.n1127 3.1505
R3964 VDD.n1127 VDD.n1126 3.1505
R3965 VDD.n1125 VDD.n1124 3.1505
R3966 VDD.n1124 VDD.n1123 3.1505
R3967 VDD.n1122 VDD.n1121 3.1505
R3968 VDD.n1121 VDD.n1120 3.1505
R3969 VDD.n1119 VDD.n1118 3.1505
R3970 VDD.n1118 VDD.n1117 3.1505
R3971 VDD.n1115 VDD.n1114 3.1505
R3972 VDD.n1114 VDD.n1113 3.1505
R3973 VDD.n1112 VDD.n1111 3.1505
R3974 VDD.n1111 VDD.n1110 3.1505
R3975 VDD.n1108 VDD.n1107 3.1505
R3976 VDD.n1107 VDD.n1106 3.1505
R3977 VDD.n1105 VDD.n1104 3.1505
R3978 VDD.n1104 VDD.n1103 3.1505
R3979 VDD.n1102 VDD.n1101 3.1505
R3980 VDD.n1101 VDD.n1100 3.1505
R3981 VDD.n1099 VDD.n1098 3.1505
R3982 VDD.n1098 VDD.n1097 3.1505
R3983 VDD.n1096 VDD.n1095 3.1505
R3984 VDD.n1095 VDD.n1094 3.1505
R3985 VDD.n1093 VDD.n1092 3.1505
R3986 VDD.n1092 VDD.n1091 3.1505
R3987 VDD.n1090 VDD.n1089 3.1505
R3988 VDD.n1089 VDD.n1088 3.1505
R3989 VDD.n1087 VDD 3.1505
R3990 VDD.n1087 VDD.n1086 3.1505
R3991 VDD.n1085 VDD.n1083 3.1505
R3992 VDD.n1085 VDD.n1084 3.1505
R3993 VDD.n1082 VDD.n1081 3.1505
R3994 VDD.n1081 VDD.n1080 3.1505
R3995 VDD.n1079 VDD.n1078 3.1505
R3996 VDD.n1078 VDD.n1077 3.1505
R3997 VDD.n1076 VDD.n1075 3.1505
R3998 VDD.n1075 VDD.n1074 3.1505
R3999 VDD.n1073 VDD.n1072 3.1505
R4000 VDD.n1072 VDD.n1071 3.1505
R4001 VDD.n1070 VDD.n1069 3.1505
R4002 VDD.n1069 VDD.n1068 3.1505
R4003 VDD.n1067 VDD.n1066 3.1505
R4004 VDD.n1066 VDD.n1065 3.1505
R4005 VDD.n1064 VDD.n1063 3.1505
R4006 VDD.n1063 VDD.n1062 3.1505
R4007 VDD.n1061 VDD.n1060 3.1505
R4008 VDD.n1060 VDD.n1059 3.1505
R4009 VDD.n1058 VDD.n1057 3.1505
R4010 VDD.n1057 VDD.n1056 3.1505
R4011 VDD.n1055 VDD.n1053 3.1505
R4012 VDD.n1055 VDD.n1054 3.1505
R4013 VDD.n1052 VDD.n1051 3.1505
R4014 VDD.n1051 VDD.n1050 3.1505
R4015 VDD.n1049 VDD.n1048 3.1505
R4016 VDD.n1048 VDD.n1047 3.1505
R4017 VDD.n1046 VDD.n1045 3.1505
R4018 VDD.n1045 VDD.n1044 3.1505
R4019 VDD.n1043 VDD.n1042 3.1505
R4020 VDD.n1042 VDD.n1041 3.1505
R4021 VDD.n1040 VDD.n1039 3.1505
R4022 VDD.n1039 VDD.n1038 3.1505
R4023 VDD.n1037 VDD.n1036 3.1505
R4024 VDD.n1036 VDD.n1035 3.1505
R4025 VDD.n1034 VDD.n1033 3.1505
R4026 VDD.n1033 VDD.n1032 3.1505
R4027 VDD.n1031 VDD.n1030 3.1505
R4028 VDD.n1030 VDD.n1029 3.1505
R4029 VDD.n1028 VDD.n1027 3.1505
R4030 VDD.n1027 VDD.n1026 3.1505
R4031 VDD.n1025 VDD 3.1505
R4032 VDD.n1025 VDD.n1024 3.1505
R4033 VDD.n1023 VDD.n1021 3.1505
R4034 VDD.n1023 VDD.n1022 3.1505
R4035 VDD.n1020 VDD.n1019 3.1505
R4036 VDD.n1019 VDD.n1018 3.1505
R4037 VDD.n1017 VDD.n1016 3.1505
R4038 VDD.n1016 VDD.n1015 3.1505
R4039 VDD.n1014 VDD.n1013 3.1505
R4040 VDD.n1013 VDD.n1012 3.1505
R4041 VDD.n1011 VDD.n1010 3.1505
R4042 VDD.n1010 VDD.n1009 3.1505
R4043 VDD.n1008 VDD.n1007 3.1505
R4044 VDD.n1007 VDD.n1006 3.1505
R4045 VDD.n1005 VDD.n1004 3.1505
R4046 VDD.n882 VDD.n881 3.1505
R4047 VDD.n881 VDD.n880 3.1505
R4048 VDD.n885 VDD.n884 3.1505
R4049 VDD.n884 VDD.n883 3.1505
R4050 VDD.n888 VDD.n887 3.1505
R4051 VDD.n887 VDD.n886 3.1505
R4052 VDD.n823 VDD.n822 3.1505
R4053 VDD.n822 VDD.n821 3.1505
R4054 VDD.n826 VDD.n825 3.1505
R4055 VDD.n825 VDD.n824 3.1505
R4056 VDD.n866 VDD.n865 3.1505
R4057 VDD.n865 VDD.n864 3.1505
R4058 VDD.n870 VDD.n869 3.1505
R4059 VDD.n920 VDD.n919 3.1505
R4060 VDD.n919 VDD.n918 3.1505
R4061 VDD.n923 VDD.n922 3.1505
R4062 VDD.n922 VDD.n921 3.1505
R4063 VDD.n833 VDD.n832 3.1505
R4064 VDD.n998 VDD.n997 3.1505
R4065 VDD.n995 VDD.n994 3.1505
R4066 VDD.n994 VDD.n993 3.1505
R4067 VDD.n992 VDD.n991 3.1505
R4068 VDD.n991 VDD.n990 3.1505
R4069 VDD.n989 VDD.n988 3.1505
R4070 VDD.n988 VDD.n987 3.1505
R4071 VDD.n986 VDD.n985 3.1505
R4072 VDD.n985 VDD.n984 3.1505
R4073 VDD.n983 VDD.n982 3.1505
R4074 VDD.n982 VDD.n981 3.1505
R4075 VDD.n980 VDD.n979 3.1505
R4076 VDD.n979 VDD.n978 3.1505
R4077 VDD.n977 VDD 3.1505
R4078 VDD.n977 VDD.n976 3.1505
R4079 VDD.n975 VDD.n973 3.1505
R4080 VDD.n975 VDD.n974 3.1505
R4081 VDD.n972 VDD.n971 3.1505
R4082 VDD.n971 VDD.n970 3.1505
R4083 VDD.n969 VDD.n968 3.1505
R4084 VDD.n968 VDD.n967 3.1505
R4085 VDD.n966 VDD.n965 3.1505
R4086 VDD.n965 VDD.n964 3.1505
R4087 VDD.n963 VDD.n962 3.1505
R4088 VDD.n962 VDD.n961 3.1505
R4089 VDD.n960 VDD.n959 3.1505
R4090 VDD.n959 VDD.n958 3.1505
R4091 VDD.n957 VDD.n956 3.1505
R4092 VDD.n956 VDD.n955 3.1505
R4093 VDD.n954 VDD.n953 3.1505
R4094 VDD.n953 VDD.n952 3.1505
R4095 VDD.n951 VDD.n950 3.1505
R4096 VDD.n950 VDD.n949 3.1505
R4097 VDD.n948 VDD.n947 3.1505
R4098 VDD.n947 VDD.n946 3.1505
R4099 VDD.n945 VDD.n944 3.1505
R4100 VDD.n944 VDD.n943 3.1505
R4101 VDD.n942 VDD.n941 3.1505
R4102 VDD.n941 VDD.n940 3.1505
R4103 VDD.n939 VDD.n938 3.1505
R4104 VDD.n938 VDD.n937 3.1505
R4105 VDD.n787 VDD.n706 3.06224
R4106 VDD.n787 VDD.n708 3.06224
R4107 VDD.n680 VDD.n599 3.06224
R4108 VDD.n680 VDD.n601 3.06224
R4109 VDD.n572 VDD.n177 3.06224
R4110 VDD.n804 VDD.n175 3.06224
R4111 VDD.n690 VDD.n689 2.6738
R4112 VDD.n596 VDD.n595 2.67318
R4113 VDD.n592 VDD.n581 2.6255
R4114 VDD.n581 VDD.n580 2.6255
R4115 VDD.n693 VDD.n692 2.6255
R4116 VDD.n692 VDD.n691 2.6255
R4117 VDD.n837 VDD.n836 2.6255
R4118 VDD.n836 VDD.n835 2.6255
R4119 VDD.n66 VDD 2.4698
R4120 VDD.n925 VDD.n143 2.2512
R4121 VDD.n891 VDD.n890 2.2512
R4122 VDD.n862 VDD.n861 2.2512
R4123 VDD.n889 VDD.n878 2.2498
R4124 VDD.n842 VDD.n841 2.24899
R4125 VDD.n927 VDD.n926 2.24859
R4126 VDD.n908 VDD.n907 2.24679
R4127 VDD.n795 VDD.n794 2.24619
R4128 VDD.n795 VDD.n704 2.24599
R4129 VDD.n689 VDD.n688 2.24362
R4130 VDD.n1242 VDD.t42 1.83033
R4131 VDD.n1185 VDD.t58 1.83033
R4132 VDD.n1152 VDD.t64 1.83033
R4133 VDD.n1071 VDD.t75 1.83033
R4134 VDD.n1038 VDD.t4 1.83033
R4135 VDD.n291 VDD.t154 1.83033
R4136 VDD.n311 VDD.t134 1.83033
R4137 VDD.n346 VDD.t295 1.83033
R4138 VDD.n366 VDD.t115 1.83033
R4139 VDD.n400 VDD.t35 1.83033
R4140 VDD.n458 VDD.t245 1.83033
R4141 VDD.n478 VDD.t87 1.83033
R4142 VDD.n513 VDD.t103 1.83033
R4143 VDD.n533 VDD.t252 1.83033
R4144 VDD.n708 VDD.t140 1.8205
R4145 VDD.n708 VDD.n707 1.8205
R4146 VDD.n706 VDD.t175 1.8205
R4147 VDD.n706 VDD.n705 1.8205
R4148 VDD.n601 VDD.t153 1.8205
R4149 VDD.n601 VDD.n600 1.8205
R4150 VDD.n599 VDD.t111 1.8205
R4151 VDD.n599 VDD.n598 1.8205
R4152 VDD.n177 VDD.t167 1.8205
R4153 VDD.n177 VDD.n176 1.8205
R4154 VDD.n175 VDD.t204 1.8205
R4155 VDD.n175 VDD.n174 1.8205
R4156 VDD.n206 VDD.n204 1.7854
R4157 VDD.n202 VDD.n193 1.7854
R4158 VDD.n199 VDD.n198 1.7854
R4159 VDD.n219 VDD.n217 1.7854
R4160 VDD.n215 VDD.n209 1.7854
R4161 VDD.n212 VDD.n207 1.7854
R4162 VDD.n232 VDD.n230 1.7854
R4163 VDD.n228 VDD.n222 1.7854
R4164 VDD.n225 VDD.n220 1.7854
R4165 VDD.n551 VDD.n237 1.7854
R4166 VDD.n760 VDD.n758 1.78487
R4167 VDD.n742 VDD.n740 1.78487
R4168 VDD.n724 VDD.n722 1.78487
R4169 VDD.n653 VDD.n651 1.78487
R4170 VDD.n635 VDD.n633 1.78487
R4171 VDD.n617 VDD.n615 1.78487
R4172 VDD.n190 VDD.n188 1.78487
R4173 VDD.n185 VDD.n183 1.78487
R4174 VDD.n234 VDD.n180 1.78487
R4175 VDD.n198 VDD.n197 1.78487
R4176 VDD.n202 VDD.n201 1.78487
R4177 VDD.n210 VDD.n207 1.78487
R4178 VDD.n215 VDD.n214 1.78487
R4179 VDD.n223 VDD.n220 1.78487
R4180 VDD.n228 VDD.n227 1.78487
R4181 VDD.n720 VDD.n717 1.78473
R4182 VDD.n714 VDD.n713 1.78473
R4183 VDD.n738 VDD.n735 1.78473
R4184 VDD.n731 VDD.n730 1.78473
R4185 VDD.n756 VDD.n753 1.78473
R4186 VDD.n749 VDD.n748 1.78473
R4187 VDD.n764 VDD.n762 1.78473
R4188 VDD.n756 VDD.n755 1.78473
R4189 VDD.n751 VDD.n748 1.78473
R4190 VDD.n747 VDD.n746 1.78473
R4191 VDD.n738 VDD.n737 1.78473
R4192 VDD.n733 VDD.n730 1.78473
R4193 VDD.n729 VDD.n728 1.78473
R4194 VDD.n720 VDD.n719 1.78473
R4195 VDD.n715 VDD.n714 1.78473
R4196 VDD.n613 VDD.n610 1.78473
R4197 VDD.n607 VDD.n606 1.78473
R4198 VDD.n631 VDD.n628 1.78473
R4199 VDD.n624 VDD.n623 1.78473
R4200 VDD.n649 VDD.n646 1.78473
R4201 VDD.n642 VDD.n641 1.78473
R4202 VDD.n657 VDD.n655 1.78473
R4203 VDD.n649 VDD.n648 1.78473
R4204 VDD.n644 VDD.n641 1.78473
R4205 VDD.n640 VDD.n639 1.78473
R4206 VDD.n631 VDD.n630 1.78473
R4207 VDD.n626 VDD.n623 1.78473
R4208 VDD.n622 VDD.n621 1.78473
R4209 VDD.n613 VDD.n612 1.78473
R4210 VDD.n608 VDD.n607 1.78473
R4211 VDD.n586 VDD.n585 1.78473
R4212 VDD.n143 VDD.n142 1.75132
R4213 VDD.n906 VDD.n905 1.75132
R4214 VDD.n892 VDD.n891 1.75132
R4215 VDD.n861 VDD.n859 1.75132
R4216 VDD.n840 VDD.n839 1.74291
R4217 VDD.n912 VDD.n910 1.663
R4218 VDD.n766 VDD 1.6259
R4219 VDD.n659 VDD 1.6259
R4220 VDD.n767 VDD.n766 1.58417
R4221 VDD.n660 VDD.n659 1.58417
R4222 VDD.n142 VDD.n141 1.49913
R4223 VDD.n905 VDD.n904 1.49913
R4224 VDD.n893 VDD.n892 1.49913
R4225 VDD.n859 VDD.n858 1.49913
R4226 VDD.n876 VDD.n874 1.4005
R4227 VDD.n139 VDD.n137 1.313
R4228 VDD.n270 VDD.n269 1.24485
R4229 VDD.n261 VDD.n260 1.24485
R4230 VDD.n257 VDD.n256 1.24485
R4231 VDD.n259 VDD.n258 1.24485
R4232 VDD.n248 VDD.n247 1.24485
R4233 VDD.n246 VDD.n244 1.24485
R4234 VDD.n239 VDD.n238 1.24485
R4235 VDD.n255 VDD.n254 1.24485
R4236 VDD.n268 VDD.n267 1.24485
R4237 VDD.n277 VDD.n276 1.24485
R4238 VDD.n4 VDD.n2 1.24485
R4239 VDD.n9 VDD.n8 1.24485
R4240 VDD.n36 VDD.n34 1.24485
R4241 VDD.n41 VDD.n40 1.24485
R4242 VDD.n43 VDD.n42 1.24485
R4243 VDD.n45 VDD.n44 1.24485
R4244 VDD.n50 VDD.n48 1.24485
R4245 VDD.n55 VDD.n54 1.24485
R4246 VDD.n57 VDD.n56 1.24485
R4247 VDD.n59 VDD.n58 1.24485
R4248 VDD.n829 VDD.n828 1.24485
R4249 VDD.n64 VDD.n63 1.24485
R4250 VDD.n149 VDD.n147 1.2255
R4251 VDD.n817 VDD.n815 1.138
R4252 VDD.n594 VDD.n593 1.12416
R4253 VDD.n839 VDD.n837 1.12383
R4254 VDD.n326 VDD.n270 0.935717
R4255 VDD.n381 VDD.n261 0.935717
R4256 VDD.n438 VDD.n257 0.935717
R4257 VDD.n438 VDD.n259 0.935717
R4258 VDD.n493 VDD.n248 0.935717
R4259 VDD.n500 VDD.n246 0.935717
R4260 VDD.n548 VDD.n239 0.935717
R4261 VDD.n445 VDD.n255 0.935717
R4262 VDD.n333 VDD.n268 0.935717
R4263 VDD.n278 VDD.n277 0.935717
R4264 VDD.n10 VDD.n4 0.935717
R4265 VDD.n10 VDD.n9 0.935717
R4266 VDD.n1223 VDD.n36 0.935717
R4267 VDD.n1223 VDD.n41 0.935717
R4268 VDD.n1116 VDD.n43 0.935717
R4269 VDD.n1116 VDD.n45 0.935717
R4270 VDD.n1109 VDD.n50 0.935717
R4271 VDD.n1109 VDD.n55 0.935717
R4272 VDD.n1002 VDD.n57 0.935717
R4273 VDD.n1002 VDD.n59 0.935717
R4274 VDD.n830 VDD.n829 0.935717
R4275 VDD.n999 VDD.n64 0.935717
R4276 VDD.n976 VDD.t97 0.890972
R4277 VDD.n873 VDD.t54 0.890972
R4278 VDD.n931 VDD.n929 0.8755
R4279 VDD.n550 VDD.n549 0.794429
R4280 VDD.n546 VDD.n545 0.720389
R4281 VDD.n12 VDD.n11 0.720389
R4282 VDD.n280 VDD.n279 0.720179
R4283 VDD.n1004 VDD.n1003 0.720179
R4284 VDD.n767 VDD.n760 0.684371
R4285 VDD.n767 VDD.n742 0.684371
R4286 VDD.n767 VDD.n724 0.684371
R4287 VDD.n660 VDD.n653 0.684371
R4288 VDD.n660 VDD.n635 0.684371
R4289 VDD.n660 VDD.n617 0.684371
R4290 VDD.n553 VDD.n552 0.684371
R4291 VDD.n552 VDD.n190 0.684371
R4292 VDD.n552 VDD.n185 0.684371
R4293 VDD.n552 VDD.n180 0.684371
R4294 VDD.n584 VDD.n582 0.684371
R4295 VDD.n552 VDD.n202 0.684371
R4296 VDD.n552 VDD.n206 0.684371
R4297 VDD.n552 VDD.n215 0.684371
R4298 VDD.n552 VDD.n207 0.684371
R4299 VDD.n552 VDD.n219 0.684371
R4300 VDD.n552 VDD.n228 0.684371
R4301 VDD.n552 VDD.n220 0.684371
R4302 VDD.n552 VDD.n232 0.684371
R4303 VDD.n552 VDD.n551 0.684371
R4304 VDD.n767 VDD.n762 0.684132
R4305 VDD.n767 VDD.n756 0.684132
R4306 VDD.n767 VDD.n748 0.684132
R4307 VDD.n767 VDD.n747 0.684132
R4308 VDD.n767 VDD.n738 0.684132
R4309 VDD.n767 VDD.n730 0.684132
R4310 VDD.n767 VDD.n729 0.684132
R4311 VDD.n767 VDD.n720 0.684132
R4312 VDD.n768 VDD.n767 0.684132
R4313 VDD.n660 VDD.n655 0.684132
R4314 VDD.n660 VDD.n649 0.684132
R4315 VDD.n660 VDD.n641 0.684132
R4316 VDD.n660 VDD.n640 0.684132
R4317 VDD.n660 VDD.n631 0.684132
R4318 VDD.n660 VDD.n623 0.684132
R4319 VDD.n660 VDD.n622 0.684132
R4320 VDD.n660 VDD.n613 0.684132
R4321 VDD.n661 VDD.n660 0.684132
R4322 VDD.n585 VDD.n584 0.684132
R4323 VDD.n874 VDD.n872 0.613
R4324 VDD.n159 VDD.n157 0.613
R4325 VDD.n1001 VDD.n1000 0.557375
R4326 VDD.n997 VDD.n996 0.460561
R4327 VDD.n832 VDD.n831 0.460561
R4328 VDD.n1257 VDD.t40 0.457957
R4329 VDD.n1200 VDD.t57 0.457957
R4330 VDD.n1138 VDD.t61 0.457957
R4331 VDD.n1086 VDD.t76 0.457957
R4332 VDD.n1024 VDD.t6 0.457957
R4333 VDD.n271 VDD.t133 0.457957
R4334 VDD.n303 VDD.t160 0.457957
R4335 VDD.n262 VDD.t114 0.457957
R4336 VDD.n358 VDD.t293 0.457957
R4337 VDD.n415 VDD.t33 0.457957
R4338 VDD.n249 VDD.t88 0.457957
R4339 VDD.n470 VDD.t241 0.457957
R4340 VDD.n240 VDD.t248 0.457957
R4341 VDD.n525 VDD.t102 0.457957
R4342 VDD.n685 VDD.n684 0.250031
R4343 VDD.n697 VDD.n696 0.230164
R4344 VDD.n799 VDD.n798 0.150959
R4345 VDD.n772 VDD.n769 0.103357
R4346 VDD.n665 VDD.n662 0.103357
R4347 VDD.n557 VDD.n554 0.103357
R4348 VDD.n76 VDD.n73 0.103357
R4349 VDD.n100 VDD.n97 0.103357
R4350 VDD.n332 VDD.n329 0.0969286
R4351 VDD.n387 VDD.n384 0.0969286
R4352 VDD.n444 VDD.n441 0.0969286
R4353 VDD.n499 VDD.n496 0.0969286
R4354 VDD.n134 VDD.n131 0.0969286
R4355 VDD.n1229 VDD.n1226 0.0969286
R4356 VDD.n1172 VDD.n1169 0.0969286
R4357 VDD.n1115 VDD.n1112 0.0969286
R4358 VDD.n948 VDD.n945 0.0969286
R4359 VDD.n704 VDD.n703 0.0945937
R4360 VDD.n591 VDD.n590 0.0840714
R4361 VDD.n752 VDD 0.0760357
R4362 VDD VDD.n750 0.0760357
R4363 VDD.n734 VDD 0.0760357
R4364 VDD VDD.n732 0.0760357
R4365 VDD.n716 VDD 0.0760357
R4366 VDD VDD.n712 0.0760357
R4367 VDD.n712 VDD.n711 0.0760357
R4368 VDD.n775 VDD.n772 0.0760357
R4369 VDD.n778 VDD.n775 0.0760357
R4370 VDD.n779 VDD.n778 0.0760357
R4371 VDD.n779 VDD 0.0760357
R4372 VDD.n786 VDD 0.0760357
R4373 VDD.n793 VDD.n790 0.0760357
R4374 VDD.n703 VDD.n700 0.0760357
R4375 VDD.n645 VDD 0.0760357
R4376 VDD VDD.n643 0.0760357
R4377 VDD.n627 VDD 0.0760357
R4378 VDD VDD.n625 0.0760357
R4379 VDD.n609 VDD 0.0760357
R4380 VDD VDD.n605 0.0760357
R4381 VDD.n605 VDD.n604 0.0760357
R4382 VDD.n668 VDD.n665 0.0760357
R4383 VDD.n671 VDD.n668 0.0760357
R4384 VDD.n672 VDD.n671 0.0760357
R4385 VDD.n672 VDD 0.0760357
R4386 VDD.n679 VDD 0.0760357
R4387 VDD.n686 VDD.n683 0.0760357
R4388 VDD.n284 VDD.n281 0.0760357
R4389 VDD.n287 VDD.n284 0.0760357
R4390 VDD.n290 VDD.n287 0.0760357
R4391 VDD.n293 VDD.n290 0.0760357
R4392 VDD.n296 VDD.n293 0.0760357
R4393 VDD.n299 VDD.n296 0.0760357
R4394 VDD VDD.n299 0.0760357
R4395 VDD.n300 VDD 0.0760357
R4396 VDD.n300 VDD 0.0760357
R4397 VDD.n307 VDD 0.0760357
R4398 VDD.n310 VDD.n307 0.0760357
R4399 VDD.n313 VDD.n310 0.0760357
R4400 VDD.n316 VDD.n313 0.0760357
R4401 VDD.n319 VDD.n316 0.0760357
R4402 VDD.n322 VDD.n319 0.0760357
R4403 VDD.n325 VDD.n322 0.0760357
R4404 VDD.n339 VDD.n336 0.0760357
R4405 VDD.n342 VDD.n339 0.0760357
R4406 VDD.n345 VDD.n342 0.0760357
R4407 VDD.n348 VDD.n345 0.0760357
R4408 VDD.n351 VDD.n348 0.0760357
R4409 VDD.n354 VDD.n351 0.0760357
R4410 VDD VDD.n354 0.0760357
R4411 VDD.n355 VDD 0.0760357
R4412 VDD.n355 VDD 0.0760357
R4413 VDD.n362 VDD 0.0760357
R4414 VDD.n365 VDD.n362 0.0760357
R4415 VDD.n368 VDD.n365 0.0760357
R4416 VDD.n371 VDD.n368 0.0760357
R4417 VDD.n374 VDD.n371 0.0760357
R4418 VDD.n377 VDD.n374 0.0760357
R4419 VDD.n380 VDD.n377 0.0760357
R4420 VDD.n390 VDD.n387 0.0760357
R4421 VDD.n393 VDD.n390 0.0760357
R4422 VDD.n396 VDD.n393 0.0760357
R4423 VDD.n399 VDD.n396 0.0760357
R4424 VDD.n402 VDD.n399 0.0760357
R4425 VDD.n405 VDD.n402 0.0760357
R4426 VDD.n408 VDD.n405 0.0760357
R4427 VDD.n411 VDD.n408 0.0760357
R4428 VDD.n412 VDD.n411 0.0760357
R4429 VDD.n412 VDD 0.0760357
R4430 VDD.n419 VDD 0.0760357
R4431 VDD.n422 VDD.n419 0.0760357
R4432 VDD.n425 VDD.n422 0.0760357
R4433 VDD.n428 VDD.n425 0.0760357
R4434 VDD.n431 VDD.n428 0.0760357
R4435 VDD.n434 VDD.n431 0.0760357
R4436 VDD.n437 VDD.n434 0.0760357
R4437 VDD.n451 VDD.n448 0.0760357
R4438 VDD.n454 VDD.n451 0.0760357
R4439 VDD.n457 VDD.n454 0.0760357
R4440 VDD.n460 VDD.n457 0.0760357
R4441 VDD.n463 VDD.n460 0.0760357
R4442 VDD.n466 VDD.n463 0.0760357
R4443 VDD VDD.n466 0.0760357
R4444 VDD.n467 VDD 0.0760357
R4445 VDD.n467 VDD 0.0760357
R4446 VDD.n474 VDD 0.0760357
R4447 VDD.n477 VDD.n474 0.0760357
R4448 VDD.n480 VDD.n477 0.0760357
R4449 VDD.n483 VDD.n480 0.0760357
R4450 VDD.n486 VDD.n483 0.0760357
R4451 VDD.n489 VDD.n486 0.0760357
R4452 VDD.n492 VDD.n489 0.0760357
R4453 VDD.n506 VDD.n503 0.0760357
R4454 VDD.n509 VDD.n506 0.0760357
R4455 VDD.n512 VDD.n509 0.0760357
R4456 VDD.n515 VDD.n512 0.0760357
R4457 VDD.n518 VDD.n515 0.0760357
R4458 VDD.n521 VDD.n518 0.0760357
R4459 VDD VDD.n521 0.0760357
R4460 VDD.n522 VDD 0.0760357
R4461 VDD.n522 VDD 0.0760357
R4462 VDD.n529 VDD 0.0760357
R4463 VDD.n532 VDD.n529 0.0760357
R4464 VDD.n535 VDD.n532 0.0760357
R4465 VDD.n538 VDD.n535 0.0760357
R4466 VDD.n541 VDD.n538 0.0760357
R4467 VDD.n544 VDD.n541 0.0760357
R4468 VDD.n547 VDD.n544 0.0760357
R4469 VDD.n226 VDD 0.0760357
R4470 VDD VDD.n224 0.0760357
R4471 VDD.n213 VDD 0.0760357
R4472 VDD VDD.n211 0.0760357
R4473 VDD.n200 VDD 0.0760357
R4474 VDD VDD.n196 0.0760357
R4475 VDD.n196 VDD.n195 0.0760357
R4476 VDD.n560 VDD.n557 0.0760357
R4477 VDD.n563 VDD.n560 0.0760357
R4478 VDD.n564 VDD.n563 0.0760357
R4479 VDD.n564 VDD 0.0760357
R4480 VDD.n571 VDD 0.0760357
R4481 VDD.n578 VDD.n575 0.0760357
R4482 VDD.n590 VDD.n589 0.0760357
R4483 VDD.n79 VDD.n76 0.0760357
R4484 VDD.n82 VDD.n79 0.0760357
R4485 VDD.n83 VDD.n82 0.0760357
R4486 VDD.n83 VDD 0.0760357
R4487 VDD.n90 VDD 0.0760357
R4488 VDD.n93 VDD.n90 0.0760357
R4489 VDD.n103 VDD.n100 0.0760357
R4490 VDD.n106 VDD.n103 0.0760357
R4491 VDD.n107 VDD.n106 0.0760357
R4492 VDD.n107 VDD 0.0760357
R4493 VDD.n114 VDD 0.0760357
R4494 VDD.n117 VDD.n114 0.0760357
R4495 VDD.n902 VDD.n899 0.0760357
R4496 VDD.n899 VDD 0.0760357
R4497 VDD.n848 VDD.n845 0.0760357
R4498 VDD.n805 VDD 0.0760357
R4499 VDD.n803 VDD.n800 0.0760357
R4500 VDD.n16 VDD.n13 0.0760357
R4501 VDD.n19 VDD.n16 0.0760357
R4502 VDD.n22 VDD.n19 0.0760357
R4503 VDD.n25 VDD.n22 0.0760357
R4504 VDD.n28 VDD.n25 0.0760357
R4505 VDD.n31 VDD.n28 0.0760357
R4506 VDD VDD.n31 0.0760357
R4507 VDD VDD.n1256 0.0760357
R4508 VDD.n1256 VDD.n1253 0.0760357
R4509 VDD.n1253 VDD.n1250 0.0760357
R4510 VDD.n1250 VDD.n1247 0.0760357
R4511 VDD.n1247 VDD.n1244 0.0760357
R4512 VDD.n1244 VDD.n1241 0.0760357
R4513 VDD.n1241 VDD.n1238 0.0760357
R4514 VDD.n1238 VDD.n1235 0.0760357
R4515 VDD.n1235 VDD.n1232 0.0760357
R4516 VDD.n1232 VDD.n1229 0.0760357
R4517 VDD.n1222 VDD.n1219 0.0760357
R4518 VDD.n1219 VDD.n1216 0.0760357
R4519 VDD.n1216 VDD.n1213 0.0760357
R4520 VDD.n1213 VDD.n1210 0.0760357
R4521 VDD.n1210 VDD.n1207 0.0760357
R4522 VDD.n1207 VDD.n1204 0.0760357
R4523 VDD.n1204 VDD 0.0760357
R4524 VDD.n1197 VDD 0.0760357
R4525 VDD.n1197 VDD.n1196 0.0760357
R4526 VDD.n1196 VDD.n1193 0.0760357
R4527 VDD.n1193 VDD.n1190 0.0760357
R4528 VDD.n1190 VDD.n1187 0.0760357
R4529 VDD.n1187 VDD.n1184 0.0760357
R4530 VDD.n1184 VDD.n1181 0.0760357
R4531 VDD.n1181 VDD.n1178 0.0760357
R4532 VDD.n1178 VDD.n1175 0.0760357
R4533 VDD.n1175 VDD.n1172 0.0760357
R4534 VDD.n1169 VDD.n1166 0.0760357
R4535 VDD.n1166 VDD.n1163 0.0760357
R4536 VDD.n1163 VDD.n1160 0.0760357
R4537 VDD.n1160 VDD.n1157 0.0760357
R4538 VDD.n1157 VDD.n1154 0.0760357
R4539 VDD.n1154 VDD.n1151 0.0760357
R4540 VDD.n1151 VDD.n1148 0.0760357
R4541 VDD.n1148 VDD.n1145 0.0760357
R4542 VDD.n1145 VDD.n1142 0.0760357
R4543 VDD.n1142 VDD 0.0760357
R4544 VDD.n1135 VDD 0.0760357
R4545 VDD.n1135 VDD.n1134 0.0760357
R4546 VDD.n1134 VDD.n1131 0.0760357
R4547 VDD.n1131 VDD.n1128 0.0760357
R4548 VDD.n1128 VDD.n1125 0.0760357
R4549 VDD.n1125 VDD.n1122 0.0760357
R4550 VDD.n1122 VDD.n1119 0.0760357
R4551 VDD.n1108 VDD.n1105 0.0760357
R4552 VDD.n1105 VDD.n1102 0.0760357
R4553 VDD.n1102 VDD.n1099 0.0760357
R4554 VDD.n1099 VDD.n1096 0.0760357
R4555 VDD.n1096 VDD.n1093 0.0760357
R4556 VDD.n1093 VDD.n1090 0.0760357
R4557 VDD.n1090 VDD 0.0760357
R4558 VDD.n1083 VDD 0.0760357
R4559 VDD.n1083 VDD.n1082 0.0760357
R4560 VDD.n1082 VDD.n1079 0.0760357
R4561 VDD.n1079 VDD.n1076 0.0760357
R4562 VDD.n1076 VDD.n1073 0.0760357
R4563 VDD.n1073 VDD.n1070 0.0760357
R4564 VDD.n1070 VDD.n1067 0.0760357
R4565 VDD.n1067 VDD.n1064 0.0760357
R4566 VDD.n1064 VDD.n1061 0.0760357
R4567 VDD.n1061 VDD.n1058 0.0760357
R4568 VDD.n1053 VDD.n1052 0.0760357
R4569 VDD.n1052 VDD.n1049 0.0760357
R4570 VDD.n1049 VDD.n1046 0.0760357
R4571 VDD.n1046 VDD.n1043 0.0760357
R4572 VDD.n1043 VDD.n1040 0.0760357
R4573 VDD.n1040 VDD.n1037 0.0760357
R4574 VDD.n1037 VDD.n1034 0.0760357
R4575 VDD.n1034 VDD.n1031 0.0760357
R4576 VDD.n1031 VDD.n1028 0.0760357
R4577 VDD.n1028 VDD 0.0760357
R4578 VDD.n1021 VDD 0.0760357
R4579 VDD.n1021 VDD.n1020 0.0760357
R4580 VDD.n1020 VDD.n1017 0.0760357
R4581 VDD.n1017 VDD.n1014 0.0760357
R4582 VDD.n1014 VDD.n1011 0.0760357
R4583 VDD.n1011 VDD.n1008 0.0760357
R4584 VDD.n1008 VDD.n1005 0.0760357
R4585 VDD.n998 VDD.n995 0.0760357
R4586 VDD.n995 VDD.n992 0.0760357
R4587 VDD.n992 VDD.n989 0.0760357
R4588 VDD.n989 VDD.n986 0.0760357
R4589 VDD.n986 VDD.n983 0.0760357
R4590 VDD.n983 VDD.n980 0.0760357
R4591 VDD.n980 VDD 0.0760357
R4592 VDD.n973 VDD 0.0760357
R4593 VDD.n973 VDD.n972 0.0760357
R4594 VDD.n972 VDD.n969 0.0760357
R4595 VDD.n969 VDD.n966 0.0760357
R4596 VDD.n966 VDD.n963 0.0760357
R4597 VDD.n963 VDD.n960 0.0760357
R4598 VDD.n960 VDD.n957 0.0760357
R4599 VDD.n957 VDD.n954 0.0760357
R4600 VDD.n954 VDD.n951 0.0760357
R4601 VDD.n951 VDD.n948 0.0760357
R4602 VDD.n945 VDD.n942 0.0760357
R4603 VDD.n942 VDD.n939 0.0760357
R4604 VDD.n923 VDD.n920 0.0760357
R4605 VDD.n885 VDD.n882 0.0760357
R4606 VDD.n888 VDD.n885 0.0760357
R4607 VDD.n867 VDD.n866 0.0760357
R4608 VDD.n826 VDD.n823 0.0760357
R4609 VDD.n851 VDD.n848 0.0752321
R4610 VDD.n131 VDD.n128 0.0744286
R4611 VDD.n800 VDD.n797 0.073274
R4612 VDD.n920 VDD.n917 0.0728214
R4613 VDD.n593 VDD.n578 0.0716604
R4614 VDD.n868 VDD.n867 0.0704107
R4615 VDD.n168 VDD.n165 0.0688036
R4616 VDD.n812 VDD 0.068
R4617 VDD.n794 VDD.n793 0.0668722
R4618 VDD.n687 VDD.n686 0.0668722
R4619 VDD.n939 VDD.n936 0.0655893
R4620 VDD.n173 VDD.n172 0.0647857
R4621 VDD.n827 VDD.n826 0.05675
R4622 VDD.n866 VDD.n863 0.0560366
R4623 VDD.n834 VDD.n833 0.0559464
R4624 VDD.n787 VDD.n786 0.0535357
R4625 VDD.n680 VDD.n679 0.0535357
R4626 VDD.n572 VDD.n571 0.0535357
R4627 VDD.n805 VDD.n804 0.0535357
R4628 VDD.n1058 VDD 0.051125
R4629 VDD.n329 VDD.n326 0.0503214
R4630 VDD.n333 VDD.n332 0.0503214
R4631 VDD.n384 VDD.n381 0.0503214
R4632 VDD.n441 VDD.n438 0.0503214
R4633 VDD.n445 VDD.n444 0.0503214
R4634 VDD.n496 VDD.n493 0.0503214
R4635 VDD.n500 VDD.n499 0.0503214
R4636 VDD.n549 VDD.n548 0.0503214
R4637 VDD.n1226 VDD.n1223 0.0503214
R4638 VDD.n1116 VDD.n1115 0.0503214
R4639 VDD.n1112 VDD.n1109 0.0503214
R4640 VDD.n1002 VDD.n1001 0.0503214
R4641 VDD.n1000 VDD.n999 0.0503214
R4642 VDD.n73 VDD.n70 0.0495179
R4643 VDD.n845 VDD.n842 0.0492107
R4644 VDD.n924 VDD.n923 0.0471071
R4645 VDD.n1053 VDD 0.0463036
R4646 VDD.n889 VDD.n888 0.0451951
R4647 VDD VDD.n894 0.0438929
R4648 VDD.n769 VDD.n709 0.039875
R4649 VDD.n662 VDD.n602 0.039875
R4650 VDD.n554 VDD.n178 0.039875
R4651 VDD.n97 VDD.n94 0.039875
R4652 VDD.n172 VDD.n169 0.039875
R4653 VDD.n882 VDD.n879 0.039875
R4654 VDD VDD.n765 0.0382679
R4655 VDD.n700 VDD 0.0382679
R4656 VDD.n695 VDD 0.0382679
R4657 VDD VDD.n658 0.0382679
R4658 VDD.n236 VDD 0.0382679
R4659 VDD VDD.n235 0.0382679
R4660 VDD.n589 VDD 0.0382679
R4661 VDD VDD.n587 0.0382679
R4662 VDD.n69 VDD 0.0382679
R4663 VDD.n903 VDD.n902 0.0382679
R4664 VDD.n745 VDD.n744 0.0366607
R4665 VDD.n727 VDD.n726 0.0366607
R4666 VDD.n711 VDD.n709 0.0366607
R4667 VDD.n638 VDD.n637 0.0366607
R4668 VDD.n620 VDD.n619 0.0366607
R4669 VDD.n604 VDD.n602 0.0366607
R4670 VDD.n182 VDD.n181 0.0366607
R4671 VDD.n187 VDD.n186 0.0366607
R4672 VDD.n195 VDD.n178 0.0366607
R4673 VDD.n94 VDD.n93 0.0366607
R4674 VDD.n118 VDD.n117 0.0366607
R4675 VDD.n169 VDD.n168 0.0366607
R4676 VDD.n595 VDD.n594 0.0301053
R4677 VDD.n796 VDD.n795 0.0301053
R4678 VDD.n795 VDD.n690 0.0289211
R4679 VDD.n765 VDD.n763 0.0270179
R4680 VDD.n695 VDD.n694 0.0270179
R4681 VDD.n658 VDD.n656 0.0270179
R4682 VDD.n235 VDD.n233 0.0270179
R4683 VDD.n587 VDD.n583 0.0270179
R4684 VDD.n70 VDD.n69 0.0270179
R4685 VDD.n281 VDD.n278 0.0262143
R4686 VDD.n326 VDD.n325 0.0262143
R4687 VDD.n336 VDD.n333 0.0262143
R4688 VDD.n381 VDD.n380 0.0262143
R4689 VDD.n438 VDD.n437 0.0262143
R4690 VDD.n448 VDD.n445 0.0262143
R4691 VDD.n493 VDD.n492 0.0262143
R4692 VDD.n503 VDD.n500 0.0262143
R4693 VDD.n548 VDD.n547 0.0262143
R4694 VDD.n13 VDD.n10 0.0262143
R4695 VDD.n1223 VDD.n1222 0.0262143
R4696 VDD.n1119 VDD.n1116 0.0262143
R4697 VDD.n1109 VDD.n1108 0.0262143
R4698 VDD.n1005 VDD.n1002 0.0262143
R4699 VDD.n999 VDD.n998 0.0262143
R4700 VDD.n833 VDD.n830 0.0262143
R4701 VDD.n790 VDD.n787 0.023
R4702 VDD.n683 VDD.n680 0.023
R4703 VDD.n575 VDD.n572 0.023
R4704 VDD.n804 VDD.n803 0.023
R4705 VDD.n592 VDD.n591 0.0205893
R4706 VDD.n858 VDD.n857 0.0205893
R4707 VDD.n841 VDD.n840 0.0205893
R4708 VDD.n837 VDD.n834 0.0205893
R4709 VDD.n837 VDD.n827 0.0197857
R4710 VDD.n857 VDD.n854 0.0181786
R4711 VDD.n125 VDD.n122 0.017375
R4712 VDD.n890 VDD.n877 0.0165714
R4713 VDD.n914 VDD.n913 0.0157679
R4714 VDD.n689 VDD.n597 0.0157541
R4715 VDD.n597 VDD.n596 0.0151974
R4716 VDD.n141 VDD.n140 0.0149643
R4717 VDD.n893 VDD.n150 0.0141607
R4718 VDD.n877 VDD 0.0133571
R4719 VDD.n155 VDD.n154 0.0133571
R4720 VDD.n140 VDD.n135 0.0125536
R4721 VDD.n162 VDD.n150 0.01175
R4722 VDD.n925 VDD.n924 0.01175
R4723 VDD.n704 VDD.n693 0.0110223
R4724 VDD.n818 VDD.n813 0.0109464
R4725 VDD.n936 VDD.n933 0.0109464
R4726 VDD.n907 VDD.n906 0.0106437
R4727 VDD.n861 VDD.n860 0.0106437
R4728 VDD.n688 VDD.n687 0.0106222
R4729 VDD.n913 VDD.n908 0.00942171
R4730 VDD.n908 VDD.n144 0.00942171
R4731 VDD.n862 VDD.n160 0.00933929
R4732 VDD.n813 VDD.n812 0.00853571
R4733 VDD.n933 VDD.n932 0.00853571
R4734 VDD.n894 VDD.n893 0.00773214
R4735 VDD.n165 VDD.n162 0.00773214
R4736 VDD.n142 VDD.n65 0.00768806
R4737 VDD.n905 VDD.n145 0.00768806
R4738 VDD.n892 VDD.n151 0.00768806
R4739 VDD.n859 VDD.n161 0.00768806
R4740 VDD.n820 VDD.n819 0.00743315
R4741 VDD.n819 VDD.n818 0.00740569
R4742 VDD.n863 VDD.n862 0.00701873
R4743 VDD.n119 VDD.n118 0.00692857
R4744 VDD.n141 VDD.n119 0.00692857
R4745 VDD.n135 VDD.n134 0.00692857
R4746 VDD.n839 VDD.n838 0.00618576
R4747 VDD VDD.n868 0.006125
R4748 VDD.n160 VDD.n155 0.006125
R4749 VDD.n932 VDD.n927 0.00581627
R4750 VDD.n927 VDD.n925 0.00581627
R4751 VDD.n593 VDD.n592 0.00581354
R4752 VDD.n842 VDD.n820 0.00501427
R4753 VDD.n879 VDD.n144 0.00451786
R4754 VDD.n917 VDD.n914 0.00371429
R4755 VDD.n890 VDD.n889 0.00340942
R4756 VDD.n128 VDD.n125 0.00210714
R4757 VDD.n904 VDD.n903 0.00210714
R4758 VDD.n858 VDD.n173 0.00130357
R4759 VDD.n854 VDD.n851 0.00130357
R4760 Transmission_Gate_Layout_5.VIN.n105 Transmission_Gate_Layout_5.VIN.n104 8.08758
R4761 Transmission_Gate_Layout_5.VIN.n79 Transmission_Gate_Layout_5.VIN.t89 5.21612
R4762 Transmission_Gate_Layout_5.VIN.n84 Transmission_Gate_Layout_5.VIN.n68 4.4609
R4763 Transmission_Gate_Layout_5.VIN.n83 Transmission_Gate_Layout_5.VIN.n69 4.4609
R4764 Transmission_Gate_Layout_5.VIN.n82 Transmission_Gate_Layout_5.VIN.n70 4.4609
R4765 Transmission_Gate_Layout_5.VIN.n80 Transmission_Gate_Layout_5.VIN.t85 4.4609
R4766 Transmission_Gate_Layout_5.VIN.n79 Transmission_Gate_Layout_5.VIN.t91 4.4609
R4767 Transmission_Gate_Layout_5.VIN.n125 Transmission_Gate_Layout_5.VIN.n122 3.90572
R4768 Transmission_Gate_Layout_5.VIN.n58 Transmission_Gate_Layout_5.VIN.n57 3.90572
R4769 Transmission_Gate_Layout_5.VIN.n66 Transmission_Gate_Layout_5.VIN.n65 3.90572
R4770 Transmission_Gate_Layout_5.VIN.n75 Transmission_Gate_Layout_5.VIN.n72 3.90572
R4771 Transmission_Gate_Layout_5.VIN.n14 Transmission_Gate_Layout_5.VIN.n13 3.90572
R4772 Transmission_Gate_Layout_5.VIN.n133 Transmission_Gate_Layout_5.VIN.n130 3.90572
R4773 Transmission_Gate_Layout_5.VIN.n40 Transmission_Gate_Layout_5.VIN.n37 3.84485
R4774 Transmission_Gate_Layout_5.VIN.n48 Transmission_Gate_Layout_5.VIN.n45 3.84485
R4775 Transmission_Gate_Layout_5.VIN.n98 Transmission_Gate_Layout_5.VIN.n97 3.84485
R4776 Transmission_Gate_Layout_5.VIN.n22 Transmission_Gate_Layout_5.VIN.n21 3.84485
R4777 Transmission_Gate_Layout_5.VIN.n30 Transmission_Gate_Layout_5.VIN.n29 3.84485
R4778 Transmission_Gate_Layout_5.VIN.n4 Transmission_Gate_Layout_5.VIN.n1 3.84485
R4779 Transmission_Gate_Layout_5.VIN.n91 Transmission_Gate_Layout_5.VIN.n33 3.3285
R4780 Transmission_Gate_Layout_5.VIN.n90 Transmission_Gate_Layout_5.VIN.n34 3.3285
R4781 Transmission_Gate_Layout_5.VIN.n89 Transmission_Gate_Layout_5.VIN.n35 3.3285
R4782 Transmission_Gate_Layout_5.VIN.n103 Transmission_Gate_Layout_5.VIN.t68 3.3285
R4783 Transmission_Gate_Layout_5.VIN.n102 Transmission_Gate_Layout_5.VIN.t63 3.3285
R4784 Transmission_Gate_Layout_5.VIN.n101 Transmission_Gate_Layout_5.VIN.t24 3.3285
R4785 Transmission_Gate_Layout_5.VIN.n125 Transmission_Gate_Layout_5.VIN.n124 3.1505
R4786 Transmission_Gate_Layout_5.VIN.n128 Transmission_Gate_Layout_5.VIN.n127 3.1505
R4787 Transmission_Gate_Layout_5.VIN.n58 Transmission_Gate_Layout_5.VIN.n55 3.1505
R4788 Transmission_Gate_Layout_5.VIN.n59 Transmission_Gate_Layout_5.VIN.n53 3.1505
R4789 Transmission_Gate_Layout_5.VIN.n66 Transmission_Gate_Layout_5.VIN.n63 3.1505
R4790 Transmission_Gate_Layout_5.VIN.n67 Transmission_Gate_Layout_5.VIN.n61 3.1505
R4791 Transmission_Gate_Layout_5.VIN.n75 Transmission_Gate_Layout_5.VIN.n74 3.1505
R4792 Transmission_Gate_Layout_5.VIN.n78 Transmission_Gate_Layout_5.VIN.n77 3.1505
R4793 Transmission_Gate_Layout_5.VIN.n14 Transmission_Gate_Layout_5.VIN.n11 3.1505
R4794 Transmission_Gate_Layout_5.VIN.n15 Transmission_Gate_Layout_5.VIN.n9 3.1505
R4795 Transmission_Gate_Layout_5.VIN.n138 Transmission_Gate_Layout_5.VIN.n120 3.1505
R4796 Transmission_Gate_Layout_5.VIN.n139 Transmission_Gate_Layout_5.VIN.n118 3.1505
R4797 Transmission_Gate_Layout_5.VIN.n140 Transmission_Gate_Layout_5.VIN.n116 3.1505
R4798 Transmission_Gate_Layout_5.VIN.n136 Transmission_Gate_Layout_5.VIN.n135 3.1505
R4799 Transmission_Gate_Layout_5.VIN.n133 Transmission_Gate_Layout_5.VIN.n132 3.1505
R4800 Transmission_Gate_Layout_5.VIN.n100 Transmission_Gate_Layout_5.VIN.n91 2.72398
R4801 Transmission_Gate_Layout_5.VIN.n40 Transmission_Gate_Layout_5.VIN.n39 2.6005
R4802 Transmission_Gate_Layout_5.VIN.n43 Transmission_Gate_Layout_5.VIN.n42 2.6005
R4803 Transmission_Gate_Layout_5.VIN.n48 Transmission_Gate_Layout_5.VIN.n47 2.6005
R4804 Transmission_Gate_Layout_5.VIN.n51 Transmission_Gate_Layout_5.VIN.n50 2.6005
R4805 Transmission_Gate_Layout_5.VIN.n98 Transmission_Gate_Layout_5.VIN.n95 2.6005
R4806 Transmission_Gate_Layout_5.VIN.n99 Transmission_Gate_Layout_5.VIN.n93 2.6005
R4807 Transmission_Gate_Layout_5.VIN.n22 Transmission_Gate_Layout_5.VIN.n19 2.6005
R4808 Transmission_Gate_Layout_5.VIN.n23 Transmission_Gate_Layout_5.VIN.n17 2.6005
R4809 Transmission_Gate_Layout_5.VIN.n30 Transmission_Gate_Layout_5.VIN.n27 2.6005
R4810 Transmission_Gate_Layout_5.VIN.n31 Transmission_Gate_Layout_5.VIN.n25 2.6005
R4811 Transmission_Gate_Layout_5.VIN.n108 Transmission_Gate_Layout_5.VIN.n107 2.6005
R4812 Transmission_Gate_Layout_5.VIN.n111 Transmission_Gate_Layout_5.VIN.n110 2.6005
R4813 Transmission_Gate_Layout_5.VIN.n114 Transmission_Gate_Layout_5.VIN.n113 2.6005
R4814 Transmission_Gate_Layout_5.VIN.n7 Transmission_Gate_Layout_5.VIN.n6 2.6005
R4815 Transmission_Gate_Layout_5.VIN.n4 Transmission_Gate_Layout_5.VIN.n3 2.6005
R4816 Transmission_Gate_Layout_5.VIN.n82 Transmission_Gate_Layout_5.VIN.n81 2.47941
R4817 Transmission_Gate_Layout_5.VIN.n135 Transmission_Gate_Layout_5.VIN.t50 1.3109
R4818 Transmission_Gate_Layout_5.VIN.n135 Transmission_Gate_Layout_5.VIN.n134 1.3109
R4819 Transmission_Gate_Layout_5.VIN.n130 Transmission_Gate_Layout_5.VIN.t55 1.3109
R4820 Transmission_Gate_Layout_5.VIN.n130 Transmission_Gate_Layout_5.VIN.n129 1.3109
R4821 Transmission_Gate_Layout_5.VIN.n127 Transmission_Gate_Layout_5.VIN.t45 1.3109
R4822 Transmission_Gate_Layout_5.VIN.n127 Transmission_Gate_Layout_5.VIN.n126 1.3109
R4823 Transmission_Gate_Layout_5.VIN.n124 Transmission_Gate_Layout_5.VIN.t51 1.3109
R4824 Transmission_Gate_Layout_5.VIN.n124 Transmission_Gate_Layout_5.VIN.n123 1.3109
R4825 Transmission_Gate_Layout_5.VIN.n122 Transmission_Gate_Layout_5.VIN.t53 1.3109
R4826 Transmission_Gate_Layout_5.VIN.n122 Transmission_Gate_Layout_5.VIN.n121 1.3109
R4827 Transmission_Gate_Layout_5.VIN.n116 Transmission_Gate_Layout_5.VIN.t49 1.3109
R4828 Transmission_Gate_Layout_5.VIN.n116 Transmission_Gate_Layout_5.VIN.n115 1.3109
R4829 Transmission_Gate_Layout_5.VIN.n118 Transmission_Gate_Layout_5.VIN.t47 1.3109
R4830 Transmission_Gate_Layout_5.VIN.n118 Transmission_Gate_Layout_5.VIN.n117 1.3109
R4831 Transmission_Gate_Layout_5.VIN.n120 Transmission_Gate_Layout_5.VIN.t52 1.3109
R4832 Transmission_Gate_Layout_5.VIN.n120 Transmission_Gate_Layout_5.VIN.n119 1.3109
R4833 Transmission_Gate_Layout_5.VIN.n53 Transmission_Gate_Layout_5.VIN.t93 1.3109
R4834 Transmission_Gate_Layout_5.VIN.n53 Transmission_Gate_Layout_5.VIN.n52 1.3109
R4835 Transmission_Gate_Layout_5.VIN.n55 Transmission_Gate_Layout_5.VIN.t92 1.3109
R4836 Transmission_Gate_Layout_5.VIN.n55 Transmission_Gate_Layout_5.VIN.n54 1.3109
R4837 Transmission_Gate_Layout_5.VIN.n57 Transmission_Gate_Layout_5.VIN.t86 1.3109
R4838 Transmission_Gate_Layout_5.VIN.n57 Transmission_Gate_Layout_5.VIN.n56 1.3109
R4839 Transmission_Gate_Layout_5.VIN.n61 Transmission_Gate_Layout_5.VIN.t88 1.3109
R4840 Transmission_Gate_Layout_5.VIN.n61 Transmission_Gate_Layout_5.VIN.n60 1.3109
R4841 Transmission_Gate_Layout_5.VIN.n63 Transmission_Gate_Layout_5.VIN.t95 1.3109
R4842 Transmission_Gate_Layout_5.VIN.n63 Transmission_Gate_Layout_5.VIN.n62 1.3109
R4843 Transmission_Gate_Layout_5.VIN.n65 Transmission_Gate_Layout_5.VIN.t87 1.3109
R4844 Transmission_Gate_Layout_5.VIN.n65 Transmission_Gate_Layout_5.VIN.n64 1.3109
R4845 Transmission_Gate_Layout_5.VIN.n77 Transmission_Gate_Layout_5.VIN.t90 1.3109
R4846 Transmission_Gate_Layout_5.VIN.n77 Transmission_Gate_Layout_5.VIN.n76 1.3109
R4847 Transmission_Gate_Layout_5.VIN.n74 Transmission_Gate_Layout_5.VIN.t84 1.3109
R4848 Transmission_Gate_Layout_5.VIN.n74 Transmission_Gate_Layout_5.VIN.n73 1.3109
R4849 Transmission_Gate_Layout_5.VIN.n72 Transmission_Gate_Layout_5.VIN.t94 1.3109
R4850 Transmission_Gate_Layout_5.VIN.n72 Transmission_Gate_Layout_5.VIN.n71 1.3109
R4851 Transmission_Gate_Layout_5.VIN.n9 Transmission_Gate_Layout_5.VIN.t46 1.3109
R4852 Transmission_Gate_Layout_5.VIN.n9 Transmission_Gate_Layout_5.VIN.n8 1.3109
R4853 Transmission_Gate_Layout_5.VIN.n11 Transmission_Gate_Layout_5.VIN.t54 1.3109
R4854 Transmission_Gate_Layout_5.VIN.n11 Transmission_Gate_Layout_5.VIN.n10 1.3109
R4855 Transmission_Gate_Layout_5.VIN.n13 Transmission_Gate_Layout_5.VIN.t48 1.3109
R4856 Transmission_Gate_Layout_5.VIN.n13 Transmission_Gate_Layout_5.VIN.n12 1.3109
R4857 Transmission_Gate_Layout_5.VIN.n132 Transmission_Gate_Layout_5.VIN.t56 1.3109
R4858 Transmission_Gate_Layout_5.VIN.n132 Transmission_Gate_Layout_5.VIN.n131 1.3109
R4859 Transmission_Gate_Layout_5.VIN.n43 Transmission_Gate_Layout_5.VIN.n40 1.24485
R4860 Transmission_Gate_Layout_5.VIN.n51 Transmission_Gate_Layout_5.VIN.n48 1.24485
R4861 Transmission_Gate_Layout_5.VIN.n91 Transmission_Gate_Layout_5.VIN.n90 1.24485
R4862 Transmission_Gate_Layout_5.VIN.n90 Transmission_Gate_Layout_5.VIN.n89 1.24485
R4863 Transmission_Gate_Layout_5.VIN.n99 Transmission_Gate_Layout_5.VIN.n98 1.24485
R4864 Transmission_Gate_Layout_5.VIN.n103 Transmission_Gate_Layout_5.VIN.n102 1.24485
R4865 Transmission_Gate_Layout_5.VIN.n102 Transmission_Gate_Layout_5.VIN.n101 1.24485
R4866 Transmission_Gate_Layout_5.VIN.n23 Transmission_Gate_Layout_5.VIN.n22 1.24485
R4867 Transmission_Gate_Layout_5.VIN.n31 Transmission_Gate_Layout_5.VIN.n30 1.24485
R4868 Transmission_Gate_Layout_5.VIN.n111 Transmission_Gate_Layout_5.VIN.n108 1.24485
R4869 Transmission_Gate_Layout_5.VIN.n114 Transmission_Gate_Layout_5.VIN.n111 1.24485
R4870 Transmission_Gate_Layout_5.VIN.n7 Transmission_Gate_Layout_5.VIN.n4 1.24485
R4871 Transmission_Gate_Layout_5.VIN.n89 Transmission_Gate_Layout_5.VIN.n88 1.2018
R4872 Transmission_Gate_Layout_5.VIN.n32 Transmission_Gate_Layout_5.VIN.n31 1.2018
R4873 Transmission_Gate_Layout_5.VIN.n81 Transmission_Gate_Layout_5.VIN.n80 0.957239
R4874 Transmission_Gate_Layout_5.VIN.n85 Transmission_Gate_Layout_5.VIN.n84 0.957239
R4875 Transmission_Gate_Layout_5.VIN.n138 Transmission_Gate_Layout_5.VIN.n137 0.957239
R4876 Transmission_Gate_Layout_5.VIN.n137 Transmission_Gate_Layout_5.VIN.n136 0.957239
R4877 Transmission_Gate_Layout_5.VIN.n141 Transmission_Gate_Layout_5.VIN.n114 0.806587
R4878 Transmission_Gate_Layout_5.VIN.n142 Transmission_Gate_Layout_5.VIN.n7 0.806587
R4879 Transmission_Gate_Layout_5.VIN.n128 Transmission_Gate_Layout_5.VIN.n125 0.755717
R4880 Transmission_Gate_Layout_5.VIN.n59 Transmission_Gate_Layout_5.VIN.n58 0.755717
R4881 Transmission_Gate_Layout_5.VIN.n67 Transmission_Gate_Layout_5.VIN.n66 0.755717
R4882 Transmission_Gate_Layout_5.VIN.n78 Transmission_Gate_Layout_5.VIN.n75 0.755717
R4883 Transmission_Gate_Layout_5.VIN.n80 Transmission_Gate_Layout_5.VIN.n79 0.755717
R4884 Transmission_Gate_Layout_5.VIN.n84 Transmission_Gate_Layout_5.VIN.n83 0.755717
R4885 Transmission_Gate_Layout_5.VIN.n83 Transmission_Gate_Layout_5.VIN.n82 0.755717
R4886 Transmission_Gate_Layout_5.VIN.n15 Transmission_Gate_Layout_5.VIN.n14 0.755717
R4887 Transmission_Gate_Layout_5.VIN.n140 Transmission_Gate_Layout_5.VIN.n139 0.755717
R4888 Transmission_Gate_Layout_5.VIN.n139 Transmission_Gate_Layout_5.VIN.n138 0.755717
R4889 Transmission_Gate_Layout_5.VIN.n136 Transmission_Gate_Layout_5.VIN.n133 0.755717
R4890 Transmission_Gate_Layout_5.VIN.n113 Transmission_Gate_Layout_5.VIN.t6 0.7285
R4891 Transmission_Gate_Layout_5.VIN.n113 Transmission_Gate_Layout_5.VIN.n112 0.7285
R4892 Transmission_Gate_Layout_5.VIN.n110 Transmission_Gate_Layout_5.VIN.t16 0.7285
R4893 Transmission_Gate_Layout_5.VIN.n110 Transmission_Gate_Layout_5.VIN.n109 0.7285
R4894 Transmission_Gate_Layout_5.VIN.n107 Transmission_Gate_Layout_5.VIN.t21 0.7285
R4895 Transmission_Gate_Layout_5.VIN.n107 Transmission_Gate_Layout_5.VIN.n106 0.7285
R4896 Transmission_Gate_Layout_5.VIN.n93 Transmission_Gate_Layout_5.VIN.t32 0.7285
R4897 Transmission_Gate_Layout_5.VIN.n93 Transmission_Gate_Layout_5.VIN.n92 0.7285
R4898 Transmission_Gate_Layout_5.VIN.n95 Transmission_Gate_Layout_5.VIN.t27 0.7285
R4899 Transmission_Gate_Layout_5.VIN.n95 Transmission_Gate_Layout_5.VIN.n94 0.7285
R4900 Transmission_Gate_Layout_5.VIN.n97 Transmission_Gate_Layout_5.VIN.t69 0.7285
R4901 Transmission_Gate_Layout_5.VIN.n97 Transmission_Gate_Layout_5.VIN.n96 0.7285
R4902 Transmission_Gate_Layout_5.VIN.n42 Transmission_Gate_Layout_5.VIN.t31 0.7285
R4903 Transmission_Gate_Layout_5.VIN.n42 Transmission_Gate_Layout_5.VIN.n41 0.7285
R4904 Transmission_Gate_Layout_5.VIN.n39 Transmission_Gate_Layout_5.VIN.t67 0.7285
R4905 Transmission_Gate_Layout_5.VIN.n39 Transmission_Gate_Layout_5.VIN.n38 0.7285
R4906 Transmission_Gate_Layout_5.VIN.n37 Transmission_Gate_Layout_5.VIN.t58 0.7285
R4907 Transmission_Gate_Layout_5.VIN.n37 Transmission_Gate_Layout_5.VIN.n36 0.7285
R4908 Transmission_Gate_Layout_5.VIN.n50 Transmission_Gate_Layout_5.VIN.t70 0.7285
R4909 Transmission_Gate_Layout_5.VIN.n50 Transmission_Gate_Layout_5.VIN.n49 0.7285
R4910 Transmission_Gate_Layout_5.VIN.n47 Transmission_Gate_Layout_5.VIN.t28 0.7285
R4911 Transmission_Gate_Layout_5.VIN.n47 Transmission_Gate_Layout_5.VIN.n46 0.7285
R4912 Transmission_Gate_Layout_5.VIN.n45 Transmission_Gate_Layout_5.VIN.t61 0.7285
R4913 Transmission_Gate_Layout_5.VIN.n45 Transmission_Gate_Layout_5.VIN.n44 0.7285
R4914 Transmission_Gate_Layout_5.VIN.n17 Transmission_Gate_Layout_5.VIN.t12 0.7285
R4915 Transmission_Gate_Layout_5.VIN.n17 Transmission_Gate_Layout_5.VIN.n16 0.7285
R4916 Transmission_Gate_Layout_5.VIN.n19 Transmission_Gate_Layout_5.VIN.t8 0.7285
R4917 Transmission_Gate_Layout_5.VIN.n19 Transmission_Gate_Layout_5.VIN.n18 0.7285
R4918 Transmission_Gate_Layout_5.VIN.n21 Transmission_Gate_Layout_5.VIN.t1 0.7285
R4919 Transmission_Gate_Layout_5.VIN.n21 Transmission_Gate_Layout_5.VIN.n20 0.7285
R4920 Transmission_Gate_Layout_5.VIN.n25 Transmission_Gate_Layout_5.VIN.t5 0.7285
R4921 Transmission_Gate_Layout_5.VIN.n25 Transmission_Gate_Layout_5.VIN.n24 0.7285
R4922 Transmission_Gate_Layout_5.VIN.n27 Transmission_Gate_Layout_5.VIN.t22 0.7285
R4923 Transmission_Gate_Layout_5.VIN.n27 Transmission_Gate_Layout_5.VIN.n26 0.7285
R4924 Transmission_Gate_Layout_5.VIN.n29 Transmission_Gate_Layout_5.VIN.t15 0.7285
R4925 Transmission_Gate_Layout_5.VIN.n29 Transmission_Gate_Layout_5.VIN.n28 0.7285
R4926 Transmission_Gate_Layout_5.VIN.n1 Transmission_Gate_Layout_5.VIN.t23 0.7285
R4927 Transmission_Gate_Layout_5.VIN.n1 Transmission_Gate_Layout_5.VIN.n0 0.7285
R4928 Transmission_Gate_Layout_5.VIN.n3 Transmission_Gate_Layout_5.VIN.t19 0.7285
R4929 Transmission_Gate_Layout_5.VIN.n3 Transmission_Gate_Layout_5.VIN.n2 0.7285
R4930 Transmission_Gate_Layout_5.VIN.n6 Transmission_Gate_Layout_5.VIN.t9 0.7285
R4931 Transmission_Gate_Layout_5.VIN.n6 Transmission_Gate_Layout_5.VIN.n5 0.7285
R4932 Transmission_Gate_Layout_5.VIN.n86 Transmission_Gate_Layout_5.VIN.n85 0.626587
R4933 Transmission_Gate_Layout_5.VIN.n88 Transmission_Gate_Layout_5.VIN.n87 0.626587
R4934 Transmission_Gate_Layout_5.VIN.n142 Transmission_Gate_Layout_5.VIN.n141 0.626587
R4935 Transmission_Gate_Layout_5.VIN.n101 Transmission_Gate_Layout_5.VIN 0.607022
R4936 Transmission_Gate_Layout_5.VIN.n104 Transmission_Gate_Layout_5.VIN.n100 0.579785
R4937 Transmission_Gate_Layout_5.VIN.n88 Transmission_Gate_Layout_5.VIN.n43 0.575717
R4938 Transmission_Gate_Layout_5.VIN.n87 Transmission_Gate_Layout_5.VIN.n51 0.575717
R4939 Transmission_Gate_Layout_5.VIN.n100 Transmission_Gate_Layout_5.VIN.n99 0.575717
R4940 Transmission_Gate_Layout_5.VIN.n32 Transmission_Gate_Layout_5.VIN.n23 0.575717
R4941 Transmission_Gate_Layout_5.VIN.n105 Transmission_Gate_Layout_5.VIN.n32 0.570002
R4942 Transmission_Gate_Layout_5.VIN.n104 Transmission_Gate_Layout_5.VIN.n103 0.562022
R4943 Transmission_Gate_Layout_5.VIN.n108 Transmission_Gate_Layout_5.VIN.n105 0.562022
R4944 Transmission_Gate_Layout_5.VIN.n142 Transmission_Gate_Layout_5.VIN.n15 0.428978
R4945 Transmission_Gate_Layout_5.VIN.n141 Transmission_Gate_Layout_5.VIN.n140 0.428978
R4946 Transmission_Gate_Layout_5.VIN.n137 Transmission_Gate_Layout_5.VIN.n128 0.331152
R4947 Transmission_Gate_Layout_5.VIN.n86 Transmission_Gate_Layout_5.VIN.n59 0.331152
R4948 Transmission_Gate_Layout_5.VIN.n85 Transmission_Gate_Layout_5.VIN.n67 0.331152
R4949 Transmission_Gate_Layout_5.VIN.n81 Transmission_Gate_Layout_5.VIN.n78 0.331152
R4950 Transmission_Gate_Layout_5.VIN.n87 Transmission_Gate_Layout_5.VIN.n86 0.239196
R4951 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_5.VIN.n142 0.192239
R4952 Transmission_Gate_Layout_1.VIN.n186 Transmission_Gate_Layout_1.VIN 14.3992
R4953 Transmission_Gate_Layout_1.VIN.n113 Transmission_Gate_Layout_1.VIN.n111 5.21612
R4954 Transmission_Gate_Layout_1.VIN.n53 Transmission_Gate_Layout_1.VIN.t90 5.21612
R4955 Transmission_Gate_Layout_1.VIN.n59 Transmission_Gate_Layout_1.VIN.n43 4.4609
R4956 Transmission_Gate_Layout_1.VIN.n56 Transmission_Gate_Layout_1.VIN.n44 4.4609
R4957 Transmission_Gate_Layout_1.VIN.n190 Transmission_Gate_Layout_1.VIN.t132 4.4609
R4958 Transmission_Gate_Layout_1.VIN.n189 Transmission_Gate_Layout_1.VIN.t133 4.4609
R4959 Transmission_Gate_Layout_1.VIN.n188 Transmission_Gate_Layout_1.VIN.t36 4.4609
R4960 Transmission_Gate_Layout_1.VIN.n115 Transmission_Gate_Layout_1.VIN.n114 4.4609
R4961 Transmission_Gate_Layout_1.VIN.n113 Transmission_Gate_Layout_1.VIN.n112 4.4609
R4962 Transmission_Gate_Layout_1.VIN.n54 Transmission_Gate_Layout_1.VIN.t97 4.4609
R4963 Transmission_Gate_Layout_1.VIN.n53 Transmission_Gate_Layout_1.VIN.t109 4.4609
R4964 Transmission_Gate_Layout_1.VIN.n58 Transmission_Gate_Layout_1.VIN.n57 4.4609
R4965 Transmission_Gate_Layout_1.VIN.n93 Transmission_Gate_Layout_1.VIN.n92 3.90572
R4966 Transmission_Gate_Layout_1.VIN.n107 Transmission_Gate_Layout_1.VIN.n104 3.90572
R4967 Transmission_Gate_Layout_1.VIN.n130 Transmission_Gate_Layout_1.VIN.n129 3.90572
R4968 Transmission_Gate_Layout_1.VIN.n168 Transmission_Gate_Layout_1.VIN.n165 3.90572
R4969 Transmission_Gate_Layout_1.VIN.n176 Transmission_Gate_Layout_1.VIN.n173 3.90572
R4970 Transmission_Gate_Layout_1.VIN.n101 Transmission_Gate_Layout_1.VIN.n100 3.90572
R4971 Transmission_Gate_Layout_1.VIN.n33 Transmission_Gate_Layout_1.VIN.n32 3.90572
R4972 Transmission_Gate_Layout_1.VIN.n41 Transmission_Gate_Layout_1.VIN.n40 3.90572
R4973 Transmission_Gate_Layout_1.VIN.n49 Transmission_Gate_Layout_1.VIN.n46 3.90572
R4974 Transmission_Gate_Layout_1.VIN.n23 Transmission_Gate_Layout_1.VIN.n20 3.84485
R4975 Transmission_Gate_Layout_1.VIN.n6 Transmission_Gate_Layout_1.VIN.n5 3.84485
R4976 Transmission_Gate_Layout_1.VIN.n120 Transmission_Gate_Layout_1.VIN.n117 3.84485
R4977 Transmission_Gate_Layout_1.VIN.n146 Transmission_Gate_Layout_1.VIN.n145 3.84485
R4978 Transmission_Gate_Layout_1.VIN.n138 Transmission_Gate_Layout_1.VIN.n137 3.84485
R4979 Transmission_Gate_Layout_1.VIN.n83 Transmission_Gate_Layout_1.VIN.n80 3.84485
R4980 Transmission_Gate_Layout_1.VIN.n75 Transmission_Gate_Layout_1.VIN.n72 3.84485
R4981 Transmission_Gate_Layout_1.VIN.n204 Transmission_Gate_Layout_1.VIN.n203 3.84485
R4982 Transmission_Gate_Layout_1.VIN.n15 Transmission_Gate_Layout_1.VIN.n12 3.84485
R4983 Transmission_Gate_Layout_1.VIN.n66 Transmission_Gate_Layout_1.VIN.n8 3.3285
R4984 Transmission_Gate_Layout_1.VIN.n65 Transmission_Gate_Layout_1.VIN.n9 3.3285
R4985 Transmission_Gate_Layout_1.VIN.n64 Transmission_Gate_Layout_1.VIN.n10 3.3285
R4986 Transmission_Gate_Layout_1.VIN.n70 Transmission_Gate_Layout_1.VIN.t72 3.3285
R4987 Transmission_Gate_Layout_1.VIN.n69 Transmission_Gate_Layout_1.VIN.t45 3.3285
R4988 Transmission_Gate_Layout_1.VIN.n68 Transmission_Gate_Layout_1.VIN.t63 3.3285
R4989 Transmission_Gate_Layout_1.VIN.n208 Transmission_Gate_Layout_1.VIN.n207 3.3285
R4990 Transmission_Gate_Layout_1.VIN.n210 Transmission_Gate_Layout_1.VIN.n209 3.3285
R4991 Transmission_Gate_Layout_1.VIN.n212 Transmission_Gate_Layout_1.VIN.n211 3.3285
R4992 Transmission_Gate_Layout_1.VIN.n197 Transmission_Gate_Layout_1.VIN.t28 3.3285
R4993 Transmission_Gate_Layout_1.VIN.n196 Transmission_Gate_Layout_1.VIN.t125 3.3285
R4994 Transmission_Gate_Layout_1.VIN.n195 Transmission_Gate_Layout_1.VIN.t115 3.3285
R4995 Transmission_Gate_Layout_1.VIN.n93 Transmission_Gate_Layout_1.VIN.n90 3.1505
R4996 Transmission_Gate_Layout_1.VIN.n94 Transmission_Gate_Layout_1.VIN.n88 3.1505
R4997 Transmission_Gate_Layout_1.VIN.n107 Transmission_Gate_Layout_1.VIN.n106 3.1505
R4998 Transmission_Gate_Layout_1.VIN.n110 Transmission_Gate_Layout_1.VIN.n109 3.1505
R4999 Transmission_Gate_Layout_1.VIN.n130 Transmission_Gate_Layout_1.VIN.n127 3.1505
R5000 Transmission_Gate_Layout_1.VIN.n131 Transmission_Gate_Layout_1.VIN.n125 3.1505
R5001 Transmission_Gate_Layout_1.VIN.n168 Transmission_Gate_Layout_1.VIN.n167 3.1505
R5002 Transmission_Gate_Layout_1.VIN.n171 Transmission_Gate_Layout_1.VIN.n170 3.1505
R5003 Transmission_Gate_Layout_1.VIN.n176 Transmission_Gate_Layout_1.VIN.n175 3.1505
R5004 Transmission_Gate_Layout_1.VIN.n179 Transmission_Gate_Layout_1.VIN.n178 3.1505
R5005 Transmission_Gate_Layout_1.VIN.n181 Transmission_Gate_Layout_1.VIN.n163 3.1505
R5006 Transmission_Gate_Layout_1.VIN.n182 Transmission_Gate_Layout_1.VIN.n161 3.1505
R5007 Transmission_Gate_Layout_1.VIN.n183 Transmission_Gate_Layout_1.VIN.n159 3.1505
R5008 Transmission_Gate_Layout_1.VIN.n101 Transmission_Gate_Layout_1.VIN.n98 3.1505
R5009 Transmission_Gate_Layout_1.VIN.n102 Transmission_Gate_Layout_1.VIN.n96 3.1505
R5010 Transmission_Gate_Layout_1.VIN.n33 Transmission_Gate_Layout_1.VIN.n30 3.1505
R5011 Transmission_Gate_Layout_1.VIN.n34 Transmission_Gate_Layout_1.VIN.n28 3.1505
R5012 Transmission_Gate_Layout_1.VIN.n41 Transmission_Gate_Layout_1.VIN.n38 3.1505
R5013 Transmission_Gate_Layout_1.VIN.n42 Transmission_Gate_Layout_1.VIN.n36 3.1505
R5014 Transmission_Gate_Layout_1.VIN.n49 Transmission_Gate_Layout_1.VIN.n48 3.1505
R5015 Transmission_Gate_Layout_1.VIN.n52 Transmission_Gate_Layout_1.VIN.n51 3.1505
R5016 Transmission_Gate_Layout_1.VIN.n206 Transmission_Gate_Layout_1.VIN.n197 2.72398
R5017 Transmission_Gate_Layout_1.VIN.n67 Transmission_Gate_Layout_1.VIN.n66 2.72398
R5018 Transmission_Gate_Layout_1.VIN.n23 Transmission_Gate_Layout_1.VIN.n22 2.6005
R5019 Transmission_Gate_Layout_1.VIN.n26 Transmission_Gate_Layout_1.VIN.n25 2.6005
R5020 Transmission_Gate_Layout_1.VIN.n6 Transmission_Gate_Layout_1.VIN.n3 2.6005
R5021 Transmission_Gate_Layout_1.VIN.n7 Transmission_Gate_Layout_1.VIN.n1 2.6005
R5022 Transmission_Gate_Layout_1.VIN.n120 Transmission_Gate_Layout_1.VIN.n119 2.6005
R5023 Transmission_Gate_Layout_1.VIN.n123 Transmission_Gate_Layout_1.VIN.n122 2.6005
R5024 Transmission_Gate_Layout_1.VIN.n146 Transmission_Gate_Layout_1.VIN.n143 2.6005
R5025 Transmission_Gate_Layout_1.VIN.n147 Transmission_Gate_Layout_1.VIN.n141 2.6005
R5026 Transmission_Gate_Layout_1.VIN.n138 Transmission_Gate_Layout_1.VIN.n135 2.6005
R5027 Transmission_Gate_Layout_1.VIN.n139 Transmission_Gate_Layout_1.VIN.n133 2.6005
R5028 Transmission_Gate_Layout_1.VIN.n151 Transmission_Gate_Layout_1.VIN.n150 2.6005
R5029 Transmission_Gate_Layout_1.VIN.n154 Transmission_Gate_Layout_1.VIN.n153 2.6005
R5030 Transmission_Gate_Layout_1.VIN.n157 Transmission_Gate_Layout_1.VIN.n156 2.6005
R5031 Transmission_Gate_Layout_1.VIN.n83 Transmission_Gate_Layout_1.VIN.n82 2.6005
R5032 Transmission_Gate_Layout_1.VIN.n86 Transmission_Gate_Layout_1.VIN.n85 2.6005
R5033 Transmission_Gate_Layout_1.VIN.n75 Transmission_Gate_Layout_1.VIN.n74 2.6005
R5034 Transmission_Gate_Layout_1.VIN.n78 Transmission_Gate_Layout_1.VIN.n77 2.6005
R5035 Transmission_Gate_Layout_1.VIN.n204 Transmission_Gate_Layout_1.VIN.n201 2.6005
R5036 Transmission_Gate_Layout_1.VIN.n205 Transmission_Gate_Layout_1.VIN.n199 2.6005
R5037 Transmission_Gate_Layout_1.VIN.n15 Transmission_Gate_Layout_1.VIN.n14 2.6005
R5038 Transmission_Gate_Layout_1.VIN.n18 Transmission_Gate_Layout_1.VIN.n17 2.6005
R5039 Transmission_Gate_Layout_1.VIN.n188 Transmission_Gate_Layout_1.VIN.n187 2.47941
R5040 Transmission_Gate_Layout_1.VIN.n56 Transmission_Gate_Layout_1.VIN.n55 2.47941
R5041 Transmission_Gate_Layout_1.VIN.n28 Transmission_Gate_Layout_1.VIN.t96 1.3109
R5042 Transmission_Gate_Layout_1.VIN.n28 Transmission_Gate_Layout_1.VIN.n27 1.3109
R5043 Transmission_Gate_Layout_1.VIN.n30 Transmission_Gate_Layout_1.VIN.t89 1.3109
R5044 Transmission_Gate_Layout_1.VIN.n30 Transmission_Gate_Layout_1.VIN.n29 1.3109
R5045 Transmission_Gate_Layout_1.VIN.n32 Transmission_Gate_Layout_1.VIN.t101 1.3109
R5046 Transmission_Gate_Layout_1.VIN.n32 Transmission_Gate_Layout_1.VIN.n31 1.3109
R5047 Transmission_Gate_Layout_1.VIN.n88 Transmission_Gate_Layout_1.VIN.t142 1.3109
R5048 Transmission_Gate_Layout_1.VIN.n88 Transmission_Gate_Layout_1.VIN.n87 1.3109
R5049 Transmission_Gate_Layout_1.VIN.n90 Transmission_Gate_Layout_1.VIN.t139 1.3109
R5050 Transmission_Gate_Layout_1.VIN.n90 Transmission_Gate_Layout_1.VIN.n89 1.3109
R5051 Transmission_Gate_Layout_1.VIN.n92 Transmission_Gate_Layout_1.VIN.t129 1.3109
R5052 Transmission_Gate_Layout_1.VIN.n92 Transmission_Gate_Layout_1.VIN.n91 1.3109
R5053 Transmission_Gate_Layout_1.VIN.n109 Transmission_Gate_Layout_1.VIN.t136 1.3109
R5054 Transmission_Gate_Layout_1.VIN.n109 Transmission_Gate_Layout_1.VIN.n108 1.3109
R5055 Transmission_Gate_Layout_1.VIN.n106 Transmission_Gate_Layout_1.VIN.t84 1.3109
R5056 Transmission_Gate_Layout_1.VIN.n106 Transmission_Gate_Layout_1.VIN.n105 1.3109
R5057 Transmission_Gate_Layout_1.VIN.n104 Transmission_Gate_Layout_1.VIN.t143 1.3109
R5058 Transmission_Gate_Layout_1.VIN.n104 Transmission_Gate_Layout_1.VIN.n103 1.3109
R5059 Transmission_Gate_Layout_1.VIN.n125 Transmission_Gate_Layout_1.VIN.t9 1.3109
R5060 Transmission_Gate_Layout_1.VIN.n125 Transmission_Gate_Layout_1.VIN.n124 1.3109
R5061 Transmission_Gate_Layout_1.VIN.n127 Transmission_Gate_Layout_1.VIN.t2 1.3109
R5062 Transmission_Gate_Layout_1.VIN.n127 Transmission_Gate_Layout_1.VIN.n126 1.3109
R5063 Transmission_Gate_Layout_1.VIN.n129 Transmission_Gate_Layout_1.VIN.t18 1.3109
R5064 Transmission_Gate_Layout_1.VIN.n129 Transmission_Gate_Layout_1.VIN.n128 1.3109
R5065 Transmission_Gate_Layout_1.VIN.n159 Transmission_Gate_Layout_1.VIN.t6 1.3109
R5066 Transmission_Gate_Layout_1.VIN.n159 Transmission_Gate_Layout_1.VIN.n158 1.3109
R5067 Transmission_Gate_Layout_1.VIN.n161 Transmission_Gate_Layout_1.VIN.t23 1.3109
R5068 Transmission_Gate_Layout_1.VIN.n161 Transmission_Gate_Layout_1.VIN.n160 1.3109
R5069 Transmission_Gate_Layout_1.VIN.n163 Transmission_Gate_Layout_1.VIN.t15 1.3109
R5070 Transmission_Gate_Layout_1.VIN.n163 Transmission_Gate_Layout_1.VIN.n162 1.3109
R5071 Transmission_Gate_Layout_1.VIN.n170 Transmission_Gate_Layout_1.VIN.t1 1.3109
R5072 Transmission_Gate_Layout_1.VIN.n170 Transmission_Gate_Layout_1.VIN.n169 1.3109
R5073 Transmission_Gate_Layout_1.VIN.n167 Transmission_Gate_Layout_1.VIN.t10 1.3109
R5074 Transmission_Gate_Layout_1.VIN.n167 Transmission_Gate_Layout_1.VIN.n166 1.3109
R5075 Transmission_Gate_Layout_1.VIN.n165 Transmission_Gate_Layout_1.VIN.t16 1.3109
R5076 Transmission_Gate_Layout_1.VIN.n165 Transmission_Gate_Layout_1.VIN.n164 1.3109
R5077 Transmission_Gate_Layout_1.VIN.n178 Transmission_Gate_Layout_1.VIN.t19 1.3109
R5078 Transmission_Gate_Layout_1.VIN.n178 Transmission_Gate_Layout_1.VIN.n177 1.3109
R5079 Transmission_Gate_Layout_1.VIN.n175 Transmission_Gate_Layout_1.VIN.t3 1.3109
R5080 Transmission_Gate_Layout_1.VIN.n175 Transmission_Gate_Layout_1.VIN.n174 1.3109
R5081 Transmission_Gate_Layout_1.VIN.n173 Transmission_Gate_Layout_1.VIN.t11 1.3109
R5082 Transmission_Gate_Layout_1.VIN.n173 Transmission_Gate_Layout_1.VIN.n172 1.3109
R5083 Transmission_Gate_Layout_1.VIN.n96 Transmission_Gate_Layout_1.VIN.t87 1.3109
R5084 Transmission_Gate_Layout_1.VIN.n96 Transmission_Gate_Layout_1.VIN.n95 1.3109
R5085 Transmission_Gate_Layout_1.VIN.n98 Transmission_Gate_Layout_1.VIN.t24 1.3109
R5086 Transmission_Gate_Layout_1.VIN.n98 Transmission_Gate_Layout_1.VIN.n97 1.3109
R5087 Transmission_Gate_Layout_1.VIN.n100 Transmission_Gate_Layout_1.VIN.t138 1.3109
R5088 Transmission_Gate_Layout_1.VIN.n100 Transmission_Gate_Layout_1.VIN.n99 1.3109
R5089 Transmission_Gate_Layout_1.VIN.n36 Transmission_Gate_Layout_1.VIN.t105 1.3109
R5090 Transmission_Gate_Layout_1.VIN.n36 Transmission_Gate_Layout_1.VIN.n35 1.3109
R5091 Transmission_Gate_Layout_1.VIN.n38 Transmission_Gate_Layout_1.VIN.t100 1.3109
R5092 Transmission_Gate_Layout_1.VIN.n38 Transmission_Gate_Layout_1.VIN.n37 1.3109
R5093 Transmission_Gate_Layout_1.VIN.n40 Transmission_Gate_Layout_1.VIN.t108 1.3109
R5094 Transmission_Gate_Layout_1.VIN.n40 Transmission_Gate_Layout_1.VIN.n39 1.3109
R5095 Transmission_Gate_Layout_1.VIN.n51 Transmission_Gate_Layout_1.VIN.t106 1.3109
R5096 Transmission_Gate_Layout_1.VIN.n51 Transmission_Gate_Layout_1.VIN.n50 1.3109
R5097 Transmission_Gate_Layout_1.VIN.n48 Transmission_Gate_Layout_1.VIN.t95 1.3109
R5098 Transmission_Gate_Layout_1.VIN.n48 Transmission_Gate_Layout_1.VIN.n47 1.3109
R5099 Transmission_Gate_Layout_1.VIN.n46 Transmission_Gate_Layout_1.VIN.t98 1.3109
R5100 Transmission_Gate_Layout_1.VIN.n46 Transmission_Gate_Layout_1.VIN.n45 1.3109
R5101 Transmission_Gate_Layout_1.VIN.n26 Transmission_Gate_Layout_1.VIN.n23 1.24485
R5102 Transmission_Gate_Layout_1.VIN.n7 Transmission_Gate_Layout_1.VIN.n6 1.24485
R5103 Transmission_Gate_Layout_1.VIN.n123 Transmission_Gate_Layout_1.VIN.n120 1.24485
R5104 Transmission_Gate_Layout_1.VIN.n147 Transmission_Gate_Layout_1.VIN.n146 1.24485
R5105 Transmission_Gate_Layout_1.VIN.n139 Transmission_Gate_Layout_1.VIN.n138 1.24485
R5106 Transmission_Gate_Layout_1.VIN.n154 Transmission_Gate_Layout_1.VIN.n151 1.24485
R5107 Transmission_Gate_Layout_1.VIN.n157 Transmission_Gate_Layout_1.VIN.n154 1.24485
R5108 Transmission_Gate_Layout_1.VIN.n86 Transmission_Gate_Layout_1.VIN.n83 1.24485
R5109 Transmission_Gate_Layout_1.VIN.n78 Transmission_Gate_Layout_1.VIN.n75 1.24485
R5110 Transmission_Gate_Layout_1.VIN.n197 Transmission_Gate_Layout_1.VIN.n196 1.24485
R5111 Transmission_Gate_Layout_1.VIN.n196 Transmission_Gate_Layout_1.VIN.n195 1.24485
R5112 Transmission_Gate_Layout_1.VIN.n205 Transmission_Gate_Layout_1.VIN.n204 1.24485
R5113 Transmission_Gate_Layout_1.VIN.n210 Transmission_Gate_Layout_1.VIN.n208 1.24485
R5114 Transmission_Gate_Layout_1.VIN.n212 Transmission_Gate_Layout_1.VIN.n210 1.24485
R5115 Transmission_Gate_Layout_1.VIN.n69 Transmission_Gate_Layout_1.VIN.n68 1.24485
R5116 Transmission_Gate_Layout_1.VIN.n70 Transmission_Gate_Layout_1.VIN.n69 1.24485
R5117 Transmission_Gate_Layout_1.VIN.n66 Transmission_Gate_Layout_1.VIN.n65 1.24485
R5118 Transmission_Gate_Layout_1.VIN.n65 Transmission_Gate_Layout_1.VIN.n64 1.24485
R5119 Transmission_Gate_Layout_1.VIN.n18 Transmission_Gate_Layout_1.VIN.n15 1.24485
R5120 Transmission_Gate_Layout_1.VIN.n148 Transmission_Gate_Layout_1.VIN.n147 1.2018
R5121 Transmission_Gate_Layout_1.VIN.n151 Transmission_Gate_Layout_1.VIN.n148 1.2018
R5122 Transmission_Gate_Layout_1.VIN.n195 Transmission_Gate_Layout_1.VIN.n194 1.2018
R5123 Transmission_Gate_Layout_1.VIN.n208 Transmission_Gate_Layout_1.VIN.n206 1.2018
R5124 Transmission_Gate_Layout_1.VIN.n68 Transmission_Gate_Layout_1.VIN.n67 1.2018
R5125 Transmission_Gate_Layout_1.VIN.n64 Transmission_Gate_Layout_1.VIN.n63 1.2018
R5126 Transmission_Gate_Layout_1.VIN.n180 Transmission_Gate_Layout_1.VIN.n179 0.957239
R5127 Transmission_Gate_Layout_1.VIN.n181 Transmission_Gate_Layout_1.VIN.n180 0.957239
R5128 Transmission_Gate_Layout_1.VIN.n191 Transmission_Gate_Layout_1.VIN.n190 0.957239
R5129 Transmission_Gate_Layout_1.VIN.n60 Transmission_Gate_Layout_1.VIN.n59 0.957239
R5130 Transmission_Gate_Layout_1.VIN.n55 Transmission_Gate_Layout_1.VIN.n54 0.957239
R5131 Transmission_Gate_Layout_1.VIN.n185 Transmission_Gate_Layout_1.VIN.n123 0.806587
R5132 Transmission_Gate_Layout_1.VIN.n184 Transmission_Gate_Layout_1.VIN.n157 0.806587
R5133 Transmission_Gate_Layout_1.VIN.n94 Transmission_Gate_Layout_1.VIN.n93 0.755717
R5134 Transmission_Gate_Layout_1.VIN.n110 Transmission_Gate_Layout_1.VIN.n107 0.755717
R5135 Transmission_Gate_Layout_1.VIN.n115 Transmission_Gate_Layout_1.VIN.n113 0.755717
R5136 Transmission_Gate_Layout_1.VIN.n131 Transmission_Gate_Layout_1.VIN.n130 0.755717
R5137 Transmission_Gate_Layout_1.VIN.n171 Transmission_Gate_Layout_1.VIN.n168 0.755717
R5138 Transmission_Gate_Layout_1.VIN.n179 Transmission_Gate_Layout_1.VIN.n176 0.755717
R5139 Transmission_Gate_Layout_1.VIN.n183 Transmission_Gate_Layout_1.VIN.n182 0.755717
R5140 Transmission_Gate_Layout_1.VIN.n182 Transmission_Gate_Layout_1.VIN.n181 0.755717
R5141 Transmission_Gate_Layout_1.VIN.n190 Transmission_Gate_Layout_1.VIN.n189 0.755717
R5142 Transmission_Gate_Layout_1.VIN.n189 Transmission_Gate_Layout_1.VIN.n188 0.755717
R5143 Transmission_Gate_Layout_1.VIN.n102 Transmission_Gate_Layout_1.VIN.n101 0.755717
R5144 Transmission_Gate_Layout_1.VIN.n34 Transmission_Gate_Layout_1.VIN.n33 0.755717
R5145 Transmission_Gate_Layout_1.VIN.n42 Transmission_Gate_Layout_1.VIN.n41 0.755717
R5146 Transmission_Gate_Layout_1.VIN.n52 Transmission_Gate_Layout_1.VIN.n49 0.755717
R5147 Transmission_Gate_Layout_1.VIN.n54 Transmission_Gate_Layout_1.VIN.n53 0.755717
R5148 Transmission_Gate_Layout_1.VIN.n59 Transmission_Gate_Layout_1.VIN.n58 0.755717
R5149 Transmission_Gate_Layout_1.VIN.n58 Transmission_Gate_Layout_1.VIN.n56 0.755717
R5150 Transmission_Gate_Layout_1.VIN.n25 Transmission_Gate_Layout_1.VIN.t65 0.7285
R5151 Transmission_Gate_Layout_1.VIN.n25 Transmission_Gate_Layout_1.VIN.n24 0.7285
R5152 Transmission_Gate_Layout_1.VIN.n22 Transmission_Gate_Layout_1.VIN.t75 0.7285
R5153 Transmission_Gate_Layout_1.VIN.n22 Transmission_Gate_Layout_1.VIN.n21 0.7285
R5154 Transmission_Gate_Layout_1.VIN.n20 Transmission_Gate_Layout_1.VIN.t79 0.7285
R5155 Transmission_Gate_Layout_1.VIN.n20 Transmission_Gate_Layout_1.VIN.n19 0.7285
R5156 Transmission_Gate_Layout_1.VIN.n1 Transmission_Gate_Layout_1.VIN.t78 0.7285
R5157 Transmission_Gate_Layout_1.VIN.n1 Transmission_Gate_Layout_1.VIN.n0 0.7285
R5158 Transmission_Gate_Layout_1.VIN.n3 Transmission_Gate_Layout_1.VIN.t74 0.7285
R5159 Transmission_Gate_Layout_1.VIN.n3 Transmission_Gate_Layout_1.VIN.n2 0.7285
R5160 Transmission_Gate_Layout_1.VIN.n5 Transmission_Gate_Layout_1.VIN.t64 0.7285
R5161 Transmission_Gate_Layout_1.VIN.n5 Transmission_Gate_Layout_1.VIN.n4 0.7285
R5162 Transmission_Gate_Layout_1.VIN.n199 Transmission_Gate_Layout_1.VIN.t114 0.7285
R5163 Transmission_Gate_Layout_1.VIN.n199 Transmission_Gate_Layout_1.VIN.n198 0.7285
R5164 Transmission_Gate_Layout_1.VIN.n201 Transmission_Gate_Layout_1.VIN.t33 0.7285
R5165 Transmission_Gate_Layout_1.VIN.n201 Transmission_Gate_Layout_1.VIN.n200 0.7285
R5166 Transmission_Gate_Layout_1.VIN.n203 Transmission_Gate_Layout_1.VIN.t124 0.7285
R5167 Transmission_Gate_Layout_1.VIN.n203 Transmission_Gate_Layout_1.VIN.n202 0.7285
R5168 Transmission_Gate_Layout_1.VIN.n122 Transmission_Gate_Layout_1.VIN.t43 0.7285
R5169 Transmission_Gate_Layout_1.VIN.n122 Transmission_Gate_Layout_1.VIN.n121 0.7285
R5170 Transmission_Gate_Layout_1.VIN.n119 Transmission_Gate_Layout_1.VIN.t57 0.7285
R5171 Transmission_Gate_Layout_1.VIN.n119 Transmission_Gate_Layout_1.VIN.n118 0.7285
R5172 Transmission_Gate_Layout_1.VIN.n117 Transmission_Gate_Layout_1.VIN.t55 0.7285
R5173 Transmission_Gate_Layout_1.VIN.n117 Transmission_Gate_Layout_1.VIN.n116 0.7285
R5174 Transmission_Gate_Layout_1.VIN.n156 Transmission_Gate_Layout_1.VIN.t41 0.7285
R5175 Transmission_Gate_Layout_1.VIN.n156 Transmission_Gate_Layout_1.VIN.n155 0.7285
R5176 Transmission_Gate_Layout_1.VIN.n153 Transmission_Gate_Layout_1.VIN.t54 0.7285
R5177 Transmission_Gate_Layout_1.VIN.n153 Transmission_Gate_Layout_1.VIN.n152 0.7285
R5178 Transmission_Gate_Layout_1.VIN.n150 Transmission_Gate_Layout_1.VIN.t51 0.7285
R5179 Transmission_Gate_Layout_1.VIN.n150 Transmission_Gate_Layout_1.VIN.n149 0.7285
R5180 Transmission_Gate_Layout_1.VIN.n141 Transmission_Gate_Layout_1.VIN.t56 0.7285
R5181 Transmission_Gate_Layout_1.VIN.n141 Transmission_Gate_Layout_1.VIN.n140 0.7285
R5182 Transmission_Gate_Layout_1.VIN.n143 Transmission_Gate_Layout_1.VIN.t59 0.7285
R5183 Transmission_Gate_Layout_1.VIN.n143 Transmission_Gate_Layout_1.VIN.n142 0.7285
R5184 Transmission_Gate_Layout_1.VIN.n145 Transmission_Gate_Layout_1.VIN.t47 0.7285
R5185 Transmission_Gate_Layout_1.VIN.n145 Transmission_Gate_Layout_1.VIN.n144 0.7285
R5186 Transmission_Gate_Layout_1.VIN.n133 Transmission_Gate_Layout_1.VIN.t38 0.7285
R5187 Transmission_Gate_Layout_1.VIN.n133 Transmission_Gate_Layout_1.VIN.n132 0.7285
R5188 Transmission_Gate_Layout_1.VIN.n135 Transmission_Gate_Layout_1.VIN.t39 0.7285
R5189 Transmission_Gate_Layout_1.VIN.n135 Transmission_Gate_Layout_1.VIN.n134 0.7285
R5190 Transmission_Gate_Layout_1.VIN.n137 Transmission_Gate_Layout_1.VIN.t53 0.7285
R5191 Transmission_Gate_Layout_1.VIN.n137 Transmission_Gate_Layout_1.VIN.n136 0.7285
R5192 Transmission_Gate_Layout_1.VIN.n85 Transmission_Gate_Layout_1.VIN.t123 0.7285
R5193 Transmission_Gate_Layout_1.VIN.n85 Transmission_Gate_Layout_1.VIN.n84 0.7285
R5194 Transmission_Gate_Layout_1.VIN.n82 Transmission_Gate_Layout_1.VIN.t32 0.7285
R5195 Transmission_Gate_Layout_1.VIN.n82 Transmission_Gate_Layout_1.VIN.n81 0.7285
R5196 Transmission_Gate_Layout_1.VIN.n80 Transmission_Gate_Layout_1.VIN.t113 0.7285
R5197 Transmission_Gate_Layout_1.VIN.n80 Transmission_Gate_Layout_1.VIN.n79 0.7285
R5198 Transmission_Gate_Layout_1.VIN.n77 Transmission_Gate_Layout_1.VIN.t29 0.7285
R5199 Transmission_Gate_Layout_1.VIN.n77 Transmission_Gate_Layout_1.VIN.n76 0.7285
R5200 Transmission_Gate_Layout_1.VIN.n74 Transmission_Gate_Layout_1.VIN.t117 0.7285
R5201 Transmission_Gate_Layout_1.VIN.n74 Transmission_Gate_Layout_1.VIN.n73 0.7285
R5202 Transmission_Gate_Layout_1.VIN.n72 Transmission_Gate_Layout_1.VIN.t121 0.7285
R5203 Transmission_Gate_Layout_1.VIN.n72 Transmission_Gate_Layout_1.VIN.n71 0.7285
R5204 Transmission_Gate_Layout_1.VIN.n17 Transmission_Gate_Layout_1.VIN.t81 0.7285
R5205 Transmission_Gate_Layout_1.VIN.n17 Transmission_Gate_Layout_1.VIN.n16 0.7285
R5206 Transmission_Gate_Layout_1.VIN.n14 Transmission_Gate_Layout_1.VIN.t68 0.7285
R5207 Transmission_Gate_Layout_1.VIN.n14 Transmission_Gate_Layout_1.VIN.n13 0.7285
R5208 Transmission_Gate_Layout_1.VIN.n12 Transmission_Gate_Layout_1.VIN.t71 0.7285
R5209 Transmission_Gate_Layout_1.VIN.n12 Transmission_Gate_Layout_1.VIN.n11 0.7285
R5210 Transmission_Gate_Layout_1.VIN.n185 Transmission_Gate_Layout_1.VIN.n184 0.626587
R5211 Transmission_Gate_Layout_1.VIN.n192 Transmission_Gate_Layout_1.VIN.n191 0.626587
R5212 Transmission_Gate_Layout_1.VIN.n194 Transmission_Gate_Layout_1.VIN.n193 0.626587
R5213 Transmission_Gate_Layout_1.VIN.n63 Transmission_Gate_Layout_1.VIN.n62 0.626587
R5214 Transmission_Gate_Layout_1.VIN.n61 Transmission_Gate_Layout_1.VIN.n60 0.626587
R5215 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.VIN.n212 0.607022
R5216 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.VIN.n70 0.607022
R5217 Transmission_Gate_Layout_1.VIN.n187 Transmission_Gate_Layout_1.VIN.n186 0.597239
R5218 Transmission_Gate_Layout_1.VIN.n62 Transmission_Gate_Layout_1.VIN.n26 0.575717
R5219 Transmission_Gate_Layout_1.VIN.n67 Transmission_Gate_Layout_1.VIN.n7 0.575717
R5220 Transmission_Gate_Layout_1.VIN.n148 Transmission_Gate_Layout_1.VIN.n139 0.575717
R5221 Transmission_Gate_Layout_1.VIN.n193 Transmission_Gate_Layout_1.VIN.n86 0.575717
R5222 Transmission_Gate_Layout_1.VIN.n194 Transmission_Gate_Layout_1.VIN.n78 0.575717
R5223 Transmission_Gate_Layout_1.VIN.n206 Transmission_Gate_Layout_1.VIN.n205 0.575717
R5224 Transmission_Gate_Layout_1.VIN.n63 Transmission_Gate_Layout_1.VIN.n18 0.575717
R5225 Transmission_Gate_Layout_1.VIN.n185 Transmission_Gate_Layout_1.VIN.n131 0.428978
R5226 Transmission_Gate_Layout_1.VIN.n184 Transmission_Gate_Layout_1.VIN.n183 0.428978
R5227 Transmission_Gate_Layout_1.VIN.n192 Transmission_Gate_Layout_1.VIN.n94 0.331152
R5228 Transmission_Gate_Layout_1.VIN.n187 Transmission_Gate_Layout_1.VIN.n110 0.331152
R5229 Transmission_Gate_Layout_1.VIN.n180 Transmission_Gate_Layout_1.VIN.n171 0.331152
R5230 Transmission_Gate_Layout_1.VIN.n191 Transmission_Gate_Layout_1.VIN.n102 0.331152
R5231 Transmission_Gate_Layout_1.VIN.n61 Transmission_Gate_Layout_1.VIN.n34 0.331152
R5232 Transmission_Gate_Layout_1.VIN.n60 Transmission_Gate_Layout_1.VIN.n42 0.331152
R5233 Transmission_Gate_Layout_1.VIN.n55 Transmission_Gate_Layout_1.VIN.n52 0.331152
R5234 Transmission_Gate_Layout_1.VIN.n186 Transmission_Gate_Layout_1.VIN.n115 0.301804
R5235 Transmission_Gate_Layout_1.VIN.n193 Transmission_Gate_Layout_1.VIN.n192 0.239196
R5236 Transmission_Gate_Layout_1.VIN.n62 Transmission_Gate_Layout_1.VIN.n61 0.239196
R5237 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.VIN.n185 0.192239
R5238 Transmission_Gate_Layout_9.CLK.t117 Transmission_Gate_Layout_9.CLK.t43 82.9076
R5239 Transmission_Gate_Layout_9.CLK.t86 Transmission_Gate_Layout_9.CLK.t117 82.9076
R5240 Transmission_Gate_Layout_9.CLK.t19 Transmission_Gate_Layout_9.CLK.t70 82.9076
R5241 Transmission_Gate_Layout_9.CLK.t114 Transmission_Gate_Layout_9.CLK.t19 82.9076
R5242 Transmission_Gate_Layout_9.CLK.t32 Transmission_Gate_Layout_9.CLK.t65 82.9076
R5243 Transmission_Gate_Layout_9.CLK.t109 Transmission_Gate_Layout_9.CLK.t32 82.9076
R5244 Transmission_Gate_Layout_9.CLK.t64 Transmission_Gate_Layout_9.CLK.t93 82.9076
R5245 Transmission_Gate_Layout_9.CLK.t15 Transmission_Gate_Layout_9.CLK.t64 82.9076
R5246 Transmission_Gate_Layout_9.CLK.t73 Transmission_Gate_Layout_9.CLK.n86 56.4451
R5247 Transmission_Gate_Layout_9.CLK.t59 Transmission_Gate_Layout_9.CLK.n60 56.4451
R5248 Transmission_Gate_Layout_9.CLK.n26 Transmission_Gate_Layout_9.CLK.t86 49.7969
R5249 Transmission_Gate_Layout_9.CLK.n105 Transmission_Gate_Layout_9.CLK.t114 49.7969
R5250 Transmission_Gate_Layout_9.CLK.n53 Transmission_Gate_Layout_9.CLK.t109 49.7969
R5251 Transmission_Gate_Layout_9.CLK.n79 Transmission_Gate_Layout_9.CLK.t15 49.7969
R5252 Transmission_Gate_Layout_9.CLK.n80 Transmission_Gate_Layout_9.CLK.t99 39.7594
R5253 Transmission_Gate_Layout_9.CLK.n54 Transmission_Gate_Layout_9.CLK.t23 39.7594
R5254 Transmission_Gate_Layout_9.CLK.n25 Transmission_Gate_Layout_9.CLK.n24 35.0405
R5255 Transmission_Gate_Layout_9.CLK.n88 Transmission_Gate_Layout_9.CLK.n87 35.0405
R5256 Transmission_Gate_Layout_9.CLK.n104 Transmission_Gate_Layout_9.CLK.n103 35.0405
R5257 Transmission_Gate_Layout_9.CLK.n52 Transmission_Gate_Layout_9.CLK.n51 35.0405
R5258 Transmission_Gate_Layout_9.CLK.n62 Transmission_Gate_Layout_9.CLK.n61 35.0405
R5259 Transmission_Gate_Layout_9.CLK.n78 Transmission_Gate_Layout_9.CLK.n77 35.0405
R5260 Transmission_Gate_Layout_9.CLK.n26 Transmission_Gate_Layout_9.CLK.t12 31.1559
R5261 Transmission_Gate_Layout_9.CLK.n105 Transmission_Gate_Layout_9.CLK.t40 31.1559
R5262 Transmission_Gate_Layout_9.CLK.n53 Transmission_Gate_Layout_9.CLK.t31 31.1559
R5263 Transmission_Gate_Layout_9.CLK.n79 Transmission_Gate_Layout_9.CLK.t63 31.1559
R5264 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.CLK.n107 24.3453
R5265 Transmission_Gate_Layout_9.CLK.n106 Transmission_Gate_Layout_9.CLK.t8 22.0309
R5266 Transmission_Gate_Layout_9.CLK.t124 Transmission_Gate_Layout_9.CLK.n1 21.9005
R5267 Transmission_Gate_Layout_9.CLK.t116 Transmission_Gate_Layout_9.CLK.n3 21.9005
R5268 Transmission_Gate_Layout_9.CLK.t113 Transmission_Gate_Layout_9.CLK.n11 21.9005
R5269 Transmission_Gate_Layout_9.CLK.t71 Transmission_Gate_Layout_9.CLK.n13 21.9005
R5270 Transmission_Gate_Layout_9.CLK.t104 Transmission_Gate_Layout_9.CLK.n16 21.9005
R5271 Transmission_Gate_Layout_9.CLK.t69 Transmission_Gate_Layout_9.CLK.n95 21.9005
R5272 Transmission_Gate_Layout_9.CLK.n94 Transmission_Gate_Layout_9.CLK.t101 21.9005
R5273 Transmission_Gate_Layout_9.CLK.n93 Transmission_Gate_Layout_9.CLK.t67 21.9005
R5274 Transmission_Gate_Layout_9.CLK.n92 Transmission_Gate_Layout_9.CLK.t98 21.9005
R5275 Transmission_Gate_Layout_9.CLK.n91 Transmission_Gate_Layout_9.CLK.t7 21.9005
R5276 Transmission_Gate_Layout_9.CLK.n90 Transmission_Gate_Layout_9.CLK.t14 21.9005
R5277 Transmission_Gate_Layout_9.CLK.n89 Transmission_Gate_Layout_9.CLK.t49 21.9005
R5278 Transmission_Gate_Layout_9.CLK.n87 Transmission_Gate_Layout_9.CLK.t38 21.9005
R5279 Transmission_Gate_Layout_9.CLK.n88 Transmission_Gate_Layout_9.CLK.t58 21.9005
R5280 Transmission_Gate_Layout_9.CLK.t47 Transmission_Gate_Layout_9.CLK.n28 21.9005
R5281 Transmission_Gate_Layout_9.CLK.t46 Transmission_Gate_Layout_9.CLK.n36 21.9005
R5282 Transmission_Gate_Layout_9.CLK.t25 Transmission_Gate_Layout_9.CLK.n38 21.9005
R5283 Transmission_Gate_Layout_9.CLK.t3 Transmission_Gate_Layout_9.CLK.n40 21.9005
R5284 Transmission_Gate_Layout_9.CLK.t76 Transmission_Gate_Layout_9.CLK.n43 21.9005
R5285 Transmission_Gate_Layout_9.CLK.t75 Transmission_Gate_Layout_9.CLK.n69 21.9005
R5286 Transmission_Gate_Layout_9.CLK.n68 Transmission_Gate_Layout_9.CLK.t22 21.9005
R5287 Transmission_Gate_Layout_9.CLK.n67 Transmission_Gate_Layout_9.CLK.t36 21.9005
R5288 Transmission_Gate_Layout_9.CLK.n66 Transmission_Gate_Layout_9.CLK.t107 21.9005
R5289 Transmission_Gate_Layout_9.CLK.n65 Transmission_Gate_Layout_9.CLK.t53 21.9005
R5290 Transmission_Gate_Layout_9.CLK.n64 Transmission_Gate_Layout_9.CLK.t35 21.9005
R5291 Transmission_Gate_Layout_9.CLK.n63 Transmission_Gate_Layout_9.CLK.t102 21.9005
R5292 Transmission_Gate_Layout_9.CLK.n61 Transmission_Gate_Layout_9.CLK.t112 21.9005
R5293 Transmission_Gate_Layout_9.CLK.n62 Transmission_Gate_Layout_9.CLK.t84 21.9005
R5294 Transmission_Gate_Layout_9.CLK.n25 Transmission_Gate_Layout_9.CLK.t124 21.5094
R5295 Transmission_Gate_Layout_9.CLK.n24 Transmission_Gate_Layout_9.CLK.t116 21.5094
R5296 Transmission_Gate_Layout_9.CLK.n23 Transmission_Gate_Layout_9.CLK.t113 21.5094
R5297 Transmission_Gate_Layout_9.CLK.n22 Transmission_Gate_Layout_9.CLK.t115 21.5094
R5298 Transmission_Gate_Layout_9.CLK.n21 Transmission_Gate_Layout_9.CLK.t28 21.5094
R5299 Transmission_Gate_Layout_9.CLK.n20 Transmission_Gate_Layout_9.CLK.t68 21.5094
R5300 Transmission_Gate_Layout_9.CLK.n19 Transmission_Gate_Layout_9.CLK.t71 21.5094
R5301 Transmission_Gate_Layout_9.CLK.n18 Transmission_Gate_Layout_9.CLK.t104 21.5094
R5302 Transmission_Gate_Layout_9.CLK.n17 Transmission_Gate_Layout_9.CLK.t111 21.5094
R5303 Transmission_Gate_Layout_9.CLK.n96 Transmission_Gate_Layout_9.CLK.t69 21.5094
R5304 Transmission_Gate_Layout_9.CLK.n97 Transmission_Gate_Layout_9.CLK.t101 21.5094
R5305 Transmission_Gate_Layout_9.CLK.n98 Transmission_Gate_Layout_9.CLK.t67 21.5094
R5306 Transmission_Gate_Layout_9.CLK.n99 Transmission_Gate_Layout_9.CLK.t98 21.5094
R5307 Transmission_Gate_Layout_9.CLK.n100 Transmission_Gate_Layout_9.CLK.t7 21.5094
R5308 Transmission_Gate_Layout_9.CLK.n101 Transmission_Gate_Layout_9.CLK.t14 21.5094
R5309 Transmission_Gate_Layout_9.CLK.n102 Transmission_Gate_Layout_9.CLK.t49 21.5094
R5310 Transmission_Gate_Layout_9.CLK.n104 Transmission_Gate_Layout_9.CLK.t38 21.5094
R5311 Transmission_Gate_Layout_9.CLK.n103 Transmission_Gate_Layout_9.CLK.t58 21.5094
R5312 Transmission_Gate_Layout_9.CLK.n52 Transmission_Gate_Layout_9.CLK.t47 21.5094
R5313 Transmission_Gate_Layout_9.CLK.n51 Transmission_Gate_Layout_9.CLK.t46 21.5094
R5314 Transmission_Gate_Layout_9.CLK.n50 Transmission_Gate_Layout_9.CLK.t29 21.5094
R5315 Transmission_Gate_Layout_9.CLK.n49 Transmission_Gate_Layout_9.CLK.t5 21.5094
R5316 Transmission_Gate_Layout_9.CLK.n48 Transmission_Gate_Layout_9.CLK.t81 21.5094
R5317 Transmission_Gate_Layout_9.CLK.n47 Transmission_Gate_Layout_9.CLK.t25 21.5094
R5318 Transmission_Gate_Layout_9.CLK.n46 Transmission_Gate_Layout_9.CLK.t3 21.5094
R5319 Transmission_Gate_Layout_9.CLK.n45 Transmission_Gate_Layout_9.CLK.t76 21.5094
R5320 Transmission_Gate_Layout_9.CLK.n44 Transmission_Gate_Layout_9.CLK.t57 21.5094
R5321 Transmission_Gate_Layout_9.CLK.n70 Transmission_Gate_Layout_9.CLK.t75 21.5094
R5322 Transmission_Gate_Layout_9.CLK.n71 Transmission_Gate_Layout_9.CLK.t22 21.5094
R5323 Transmission_Gate_Layout_9.CLK.n72 Transmission_Gate_Layout_9.CLK.t36 21.5094
R5324 Transmission_Gate_Layout_9.CLK.n73 Transmission_Gate_Layout_9.CLK.t107 21.5094
R5325 Transmission_Gate_Layout_9.CLK.n74 Transmission_Gate_Layout_9.CLK.t53 21.5094
R5326 Transmission_Gate_Layout_9.CLK.n75 Transmission_Gate_Layout_9.CLK.t35 21.5094
R5327 Transmission_Gate_Layout_9.CLK.n76 Transmission_Gate_Layout_9.CLK.t102 21.5094
R5328 Transmission_Gate_Layout_9.CLK.n78 Transmission_Gate_Layout_9.CLK.t112 21.5094
R5329 Transmission_Gate_Layout_9.CLK.n77 Transmission_Gate_Layout_9.CLK.t84 21.5094
R5330 Transmission_Gate_Layout_9.CLK.n107 Transmission_Gate_Layout_9.CLK.t61 21.3791
R5331 Transmission_Gate_Layout_9.CLK.n106 Transmission_Gate_Layout_9.CLK.t55 21.3791
R5332 Transmission_Gate_Layout_9.CLK.n24 Transmission_Gate_Layout_9.CLK.t72 20.988
R5333 Transmission_Gate_Layout_9.CLK.n23 Transmission_Gate_Layout_9.CLK.t110 20.988
R5334 Transmission_Gate_Layout_9.CLK.n22 Transmission_Gate_Layout_9.CLK.t52 20.988
R5335 Transmission_Gate_Layout_9.CLK.n21 Transmission_Gate_Layout_9.CLK.t80 20.988
R5336 Transmission_Gate_Layout_9.CLK.n20 Transmission_Gate_Layout_9.CLK.t106 20.988
R5337 Transmission_Gate_Layout_9.CLK.n19 Transmission_Gate_Layout_9.CLK.t45 20.988
R5338 Transmission_Gate_Layout_9.CLK.n18 Transmission_Gate_Layout_9.CLK.t74 20.988
R5339 Transmission_Gate_Layout_9.CLK.n17 Transmission_Gate_Layout_9.CLK.t17 20.988
R5340 Transmission_Gate_Layout_9.CLK.t12 Transmission_Gate_Layout_9.CLK.n25 20.988
R5341 Transmission_Gate_Layout_9.CLK.n96 Transmission_Gate_Layout_9.CLK.t50 20.988
R5342 Transmission_Gate_Layout_9.CLK.n97 Transmission_Gate_Layout_9.CLK.t77 20.988
R5343 Transmission_Gate_Layout_9.CLK.n98 Transmission_Gate_Layout_9.CLK.t37 20.988
R5344 Transmission_Gate_Layout_9.CLK.n99 Transmission_Gate_Layout_9.CLK.t62 20.988
R5345 Transmission_Gate_Layout_9.CLK.n100 Transmission_Gate_Layout_9.CLK.t87 20.988
R5346 Transmission_Gate_Layout_9.CLK.n101 Transmission_Gate_Layout_9.CLK.t34 20.988
R5347 Transmission_Gate_Layout_9.CLK.n102 Transmission_Gate_Layout_9.CLK.t60 20.988
R5348 Transmission_Gate_Layout_9.CLK.n103 Transmission_Gate_Layout_9.CLK.t122 20.988
R5349 Transmission_Gate_Layout_9.CLK.t40 Transmission_Gate_Layout_9.CLK.n104 20.988
R5350 Transmission_Gate_Layout_9.CLK.n51 Transmission_Gate_Layout_9.CLK.t18 20.988
R5351 Transmission_Gate_Layout_9.CLK.n50 Transmission_Gate_Layout_9.CLK.t11 20.988
R5352 Transmission_Gate_Layout_9.CLK.n49 Transmission_Gate_Layout_9.CLK.t16 20.988
R5353 Transmission_Gate_Layout_9.CLK.n48 Transmission_Gate_Layout_9.CLK.t56 20.988
R5354 Transmission_Gate_Layout_9.CLK.n47 Transmission_Gate_Layout_9.CLK.t89 20.988
R5355 Transmission_Gate_Layout_9.CLK.n46 Transmission_Gate_Layout_9.CLK.t92 20.988
R5356 Transmission_Gate_Layout_9.CLK.n45 Transmission_Gate_Layout_9.CLK.t4 20.988
R5357 Transmission_Gate_Layout_9.CLK.n44 Transmission_Gate_Layout_9.CLK.t9 20.988
R5358 Transmission_Gate_Layout_9.CLK.t31 Transmission_Gate_Layout_9.CLK.n52 20.988
R5359 Transmission_Gate_Layout_9.CLK.n70 Transmission_Gate_Layout_9.CLK.t90 20.988
R5360 Transmission_Gate_Layout_9.CLK.n71 Transmission_Gate_Layout_9.CLK.t123 20.988
R5361 Transmission_Gate_Layout_9.CLK.n72 Transmission_Gate_Layout_9.CLK.t88 20.988
R5362 Transmission_Gate_Layout_9.CLK.n73 Transmission_Gate_Layout_9.CLK.t121 20.988
R5363 Transmission_Gate_Layout_9.CLK.n74 Transmission_Gate_Layout_9.CLK.t39 20.988
R5364 Transmission_Gate_Layout_9.CLK.n75 Transmission_Gate_Layout_9.CLK.t42 20.988
R5365 Transmission_Gate_Layout_9.CLK.n76 Transmission_Gate_Layout_9.CLK.t78 20.988
R5366 Transmission_Gate_Layout_9.CLK.n77 Transmission_Gate_Layout_9.CLK.t83 20.988
R5367 Transmission_Gate_Layout_9.CLK.t63 Transmission_Gate_Layout_9.CLK.n78 20.988
R5368 Transmission_Gate_Layout_9.CLK.n81 Transmission_Gate_Layout_9.CLK.n80 20.8576
R5369 Transmission_Gate_Layout_9.CLK.n82 Transmission_Gate_Layout_9.CLK.n81 20.8576
R5370 Transmission_Gate_Layout_9.CLK.n83 Transmission_Gate_Layout_9.CLK.n82 20.8576
R5371 Transmission_Gate_Layout_9.CLK.n84 Transmission_Gate_Layout_9.CLK.n83 20.8576
R5372 Transmission_Gate_Layout_9.CLK.n85 Transmission_Gate_Layout_9.CLK.n84 20.8576
R5373 Transmission_Gate_Layout_9.CLK.n86 Transmission_Gate_Layout_9.CLK.n85 20.8576
R5374 Transmission_Gate_Layout_9.CLK.n55 Transmission_Gate_Layout_9.CLK.n54 20.8576
R5375 Transmission_Gate_Layout_9.CLK.n56 Transmission_Gate_Layout_9.CLK.n55 20.8576
R5376 Transmission_Gate_Layout_9.CLK.n57 Transmission_Gate_Layout_9.CLK.n56 20.8576
R5377 Transmission_Gate_Layout_9.CLK.n58 Transmission_Gate_Layout_9.CLK.n57 20.8576
R5378 Transmission_Gate_Layout_9.CLK.n59 Transmission_Gate_Layout_9.CLK.n58 20.8576
R5379 Transmission_Gate_Layout_9.CLK.n60 Transmission_Gate_Layout_9.CLK.n59 20.8576
R5380 Transmission_Gate_Layout_9.CLK.n107 Transmission_Gate_Layout_9.CLK.n106 20.8576
R5381 Transmission_Gate_Layout_9.CLK.n15 Transmission_Gate_Layout_9.CLK.t20 20.5969
R5382 Transmission_Gate_Layout_9.CLK.n13 Transmission_Gate_Layout_9.CLK.t103 20.5969
R5383 Transmission_Gate_Layout_9.CLK.n8 Transmission_Gate_Layout_9.CLK.t97 20.5969
R5384 Transmission_Gate_Layout_9.CLK.n9 Transmission_Gate_Layout_9.CLK.t66 20.5969
R5385 Transmission_Gate_Layout_9.CLK.n10 Transmission_Gate_Layout_9.CLK.t27 20.5969
R5386 Transmission_Gate_Layout_9.CLK.n11 Transmission_Gate_Layout_9.CLK.t21 20.5969
R5387 Transmission_Gate_Layout_9.CLK.n3 Transmission_Gate_Layout_9.CLK.t30 20.5969
R5388 Transmission_Gate_Layout_9.CLK.n1 Transmission_Gate_Layout_9.CLK.t41 20.5969
R5389 Transmission_Gate_Layout_9.CLK.n16 Transmission_Gate_Layout_9.CLK.t13 20.5969
R5390 Transmission_Gate_Layout_9.CLK.n88 Transmission_Gate_Layout_9.CLK.t91 20.5969
R5391 Transmission_Gate_Layout_9.CLK.n89 Transmission_Gate_Layout_9.CLK.t85 20.5969
R5392 Transmission_Gate_Layout_9.CLK.n90 Transmission_Gate_Layout_9.CLK.t48 20.5969
R5393 Transmission_Gate_Layout_9.CLK.n91 Transmission_Gate_Layout_9.CLK.t44 20.5969
R5394 Transmission_Gate_Layout_9.CLK.n92 Transmission_Gate_Layout_9.CLK.t6 20.5969
R5395 Transmission_Gate_Layout_9.CLK.n93 Transmission_Gate_Layout_9.CLK.t96 20.5969
R5396 Transmission_Gate_Layout_9.CLK.n94 Transmission_Gate_Layout_9.CLK.t10 20.5969
R5397 Transmission_Gate_Layout_9.CLK.n95 Transmission_Gate_Layout_9.CLK.t99 20.5969
R5398 Transmission_Gate_Layout_9.CLK.n87 Transmission_Gate_Layout_9.CLK.t73 20.5969
R5399 Transmission_Gate_Layout_9.CLK.n28 Transmission_Gate_Layout_9.CLK.t119 20.5969
R5400 Transmission_Gate_Layout_9.CLK.n36 Transmission_Gate_Layout_9.CLK.t118 20.5969
R5401 Transmission_Gate_Layout_9.CLK.n35 Transmission_Gate_Layout_9.CLK.t100 20.5969
R5402 Transmission_Gate_Layout_9.CLK.n34 Transmission_Gate_Layout_9.CLK.t82 20.5969
R5403 Transmission_Gate_Layout_9.CLK.n33 Transmission_Gate_Layout_9.CLK.t26 20.5969
R5404 Transmission_Gate_Layout_9.CLK.n38 Transmission_Gate_Layout_9.CLK.t95 20.5969
R5405 Transmission_Gate_Layout_9.CLK.n40 Transmission_Gate_Layout_9.CLK.t79 20.5969
R5406 Transmission_Gate_Layout_9.CLK.n42 Transmission_Gate_Layout_9.CLK.t2 20.5969
R5407 Transmission_Gate_Layout_9.CLK.n43 Transmission_Gate_Layout_9.CLK.t24 20.5969
R5408 Transmission_Gate_Layout_9.CLK.n69 Transmission_Gate_Layout_9.CLK.t23 20.5969
R5409 Transmission_Gate_Layout_9.CLK.n68 Transmission_Gate_Layout_9.CLK.t94 20.5969
R5410 Transmission_Gate_Layout_9.CLK.n67 Transmission_Gate_Layout_9.CLK.t108 20.5969
R5411 Transmission_Gate_Layout_9.CLK.n66 Transmission_Gate_Layout_9.CLK.t54 20.5969
R5412 Transmission_Gate_Layout_9.CLK.n65 Transmission_Gate_Layout_9.CLK.t120 20.5969
R5413 Transmission_Gate_Layout_9.CLK.n64 Transmission_Gate_Layout_9.CLK.t105 20.5969
R5414 Transmission_Gate_Layout_9.CLK.n63 Transmission_Gate_Layout_9.CLK.t51 20.5969
R5415 Transmission_Gate_Layout_9.CLK.n62 Transmission_Gate_Layout_9.CLK.t33 20.5969
R5416 Transmission_Gate_Layout_9.CLK.n61 Transmission_Gate_Layout_9.CLK.t59 20.5969
R5417 Transmission_Gate_Layout_9.CLK.n11 Transmission_Gate_Layout_9.CLK.n10 19.4672
R5418 Transmission_Gate_Layout_9.CLK.n10 Transmission_Gate_Layout_9.CLK.n9 19.4672
R5419 Transmission_Gate_Layout_9.CLK.n9 Transmission_Gate_Layout_9.CLK.n8 19.4672
R5420 Transmission_Gate_Layout_9.CLK.n16 Transmission_Gate_Layout_9.CLK.n15 19.4672
R5421 Transmission_Gate_Layout_9.CLK.n24 Transmission_Gate_Layout_9.CLK.n23 19.4672
R5422 Transmission_Gate_Layout_9.CLK.n23 Transmission_Gate_Layout_9.CLK.n22 19.4672
R5423 Transmission_Gate_Layout_9.CLK.n22 Transmission_Gate_Layout_9.CLK.n21 19.4672
R5424 Transmission_Gate_Layout_9.CLK.n21 Transmission_Gate_Layout_9.CLK.n20 19.4672
R5425 Transmission_Gate_Layout_9.CLK.n20 Transmission_Gate_Layout_9.CLK.n19 19.4672
R5426 Transmission_Gate_Layout_9.CLK.n19 Transmission_Gate_Layout_9.CLK.n18 19.4672
R5427 Transmission_Gate_Layout_9.CLK.n18 Transmission_Gate_Layout_9.CLK.n17 19.4672
R5428 Transmission_Gate_Layout_9.CLK.n95 Transmission_Gate_Layout_9.CLK.n94 19.4672
R5429 Transmission_Gate_Layout_9.CLK.n94 Transmission_Gate_Layout_9.CLK.n93 19.4672
R5430 Transmission_Gate_Layout_9.CLK.n93 Transmission_Gate_Layout_9.CLK.n92 19.4672
R5431 Transmission_Gate_Layout_9.CLK.n92 Transmission_Gate_Layout_9.CLK.n91 19.4672
R5432 Transmission_Gate_Layout_9.CLK.n91 Transmission_Gate_Layout_9.CLK.n90 19.4672
R5433 Transmission_Gate_Layout_9.CLK.n90 Transmission_Gate_Layout_9.CLK.n89 19.4672
R5434 Transmission_Gate_Layout_9.CLK.n89 Transmission_Gate_Layout_9.CLK.n88 19.4672
R5435 Transmission_Gate_Layout_9.CLK.n97 Transmission_Gate_Layout_9.CLK.n96 19.4672
R5436 Transmission_Gate_Layout_9.CLK.n98 Transmission_Gate_Layout_9.CLK.n97 19.4672
R5437 Transmission_Gate_Layout_9.CLK.n99 Transmission_Gate_Layout_9.CLK.n98 19.4672
R5438 Transmission_Gate_Layout_9.CLK.n100 Transmission_Gate_Layout_9.CLK.n99 19.4672
R5439 Transmission_Gate_Layout_9.CLK.n101 Transmission_Gate_Layout_9.CLK.n100 19.4672
R5440 Transmission_Gate_Layout_9.CLK.n102 Transmission_Gate_Layout_9.CLK.n101 19.4672
R5441 Transmission_Gate_Layout_9.CLK.n103 Transmission_Gate_Layout_9.CLK.n102 19.4672
R5442 Transmission_Gate_Layout_9.CLK.n36 Transmission_Gate_Layout_9.CLK.n35 19.4672
R5443 Transmission_Gate_Layout_9.CLK.n35 Transmission_Gate_Layout_9.CLK.n34 19.4672
R5444 Transmission_Gate_Layout_9.CLK.n34 Transmission_Gate_Layout_9.CLK.n33 19.4672
R5445 Transmission_Gate_Layout_9.CLK.n43 Transmission_Gate_Layout_9.CLK.n42 19.4672
R5446 Transmission_Gate_Layout_9.CLK.n51 Transmission_Gate_Layout_9.CLK.n50 19.4672
R5447 Transmission_Gate_Layout_9.CLK.n50 Transmission_Gate_Layout_9.CLK.n49 19.4672
R5448 Transmission_Gate_Layout_9.CLK.n49 Transmission_Gate_Layout_9.CLK.n48 19.4672
R5449 Transmission_Gate_Layout_9.CLK.n48 Transmission_Gate_Layout_9.CLK.n47 19.4672
R5450 Transmission_Gate_Layout_9.CLK.n47 Transmission_Gate_Layout_9.CLK.n46 19.4672
R5451 Transmission_Gate_Layout_9.CLK.n46 Transmission_Gate_Layout_9.CLK.n45 19.4672
R5452 Transmission_Gate_Layout_9.CLK.n45 Transmission_Gate_Layout_9.CLK.n44 19.4672
R5453 Transmission_Gate_Layout_9.CLK.n69 Transmission_Gate_Layout_9.CLK.n68 19.4672
R5454 Transmission_Gate_Layout_9.CLK.n68 Transmission_Gate_Layout_9.CLK.n67 19.4672
R5455 Transmission_Gate_Layout_9.CLK.n67 Transmission_Gate_Layout_9.CLK.n66 19.4672
R5456 Transmission_Gate_Layout_9.CLK.n66 Transmission_Gate_Layout_9.CLK.n65 19.4672
R5457 Transmission_Gate_Layout_9.CLK.n65 Transmission_Gate_Layout_9.CLK.n64 19.4672
R5458 Transmission_Gate_Layout_9.CLK.n64 Transmission_Gate_Layout_9.CLK.n63 19.4672
R5459 Transmission_Gate_Layout_9.CLK.n63 Transmission_Gate_Layout_9.CLK.n62 19.4672
R5460 Transmission_Gate_Layout_9.CLK.n71 Transmission_Gate_Layout_9.CLK.n70 19.4672
R5461 Transmission_Gate_Layout_9.CLK.n72 Transmission_Gate_Layout_9.CLK.n71 19.4672
R5462 Transmission_Gate_Layout_9.CLK.n73 Transmission_Gate_Layout_9.CLK.n72 19.4672
R5463 Transmission_Gate_Layout_9.CLK.n74 Transmission_Gate_Layout_9.CLK.n73 19.4672
R5464 Transmission_Gate_Layout_9.CLK.n75 Transmission_Gate_Layout_9.CLK.n74 19.4672
R5465 Transmission_Gate_Layout_9.CLK.n76 Transmission_Gate_Layout_9.CLK.n75 19.4672
R5466 Transmission_Gate_Layout_9.CLK.n77 Transmission_Gate_Layout_9.CLK.n76 19.4672
R5467 Transmission_Gate_Layout_9.CLK.t103 Transmission_Gate_Layout_9.CLK.n12 18.9023
R5468 Transmission_Gate_Layout_9.CLK.t97 Transmission_Gate_Layout_9.CLK.n7 18.9023
R5469 Transmission_Gate_Layout_9.CLK.t66 Transmission_Gate_Layout_9.CLK.n6 18.9023
R5470 Transmission_Gate_Layout_9.CLK.t27 Transmission_Gate_Layout_9.CLK.n5 18.9023
R5471 Transmission_Gate_Layout_9.CLK.t21 Transmission_Gate_Layout_9.CLK.n4 18.9023
R5472 Transmission_Gate_Layout_9.CLK.t30 Transmission_Gate_Layout_9.CLK.n2 18.9023
R5473 Transmission_Gate_Layout_9.CLK.t13 Transmission_Gate_Layout_9.CLK.n14 18.9023
R5474 Transmission_Gate_Layout_9.CLK.n86 Transmission_Gate_Layout_9.CLK.t91 18.9023
R5475 Transmission_Gate_Layout_9.CLK.n85 Transmission_Gate_Layout_9.CLK.t85 18.9023
R5476 Transmission_Gate_Layout_9.CLK.n84 Transmission_Gate_Layout_9.CLK.t48 18.9023
R5477 Transmission_Gate_Layout_9.CLK.n83 Transmission_Gate_Layout_9.CLK.t44 18.9023
R5478 Transmission_Gate_Layout_9.CLK.n82 Transmission_Gate_Layout_9.CLK.t6 18.9023
R5479 Transmission_Gate_Layout_9.CLK.n81 Transmission_Gate_Layout_9.CLK.t96 18.9023
R5480 Transmission_Gate_Layout_9.CLK.n80 Transmission_Gate_Layout_9.CLK.t10 18.9023
R5481 Transmission_Gate_Layout_9.CLK.t118 Transmission_Gate_Layout_9.CLK.n29 18.9023
R5482 Transmission_Gate_Layout_9.CLK.t100 Transmission_Gate_Layout_9.CLK.n30 18.9023
R5483 Transmission_Gate_Layout_9.CLK.t82 Transmission_Gate_Layout_9.CLK.n31 18.9023
R5484 Transmission_Gate_Layout_9.CLK.t26 Transmission_Gate_Layout_9.CLK.n32 18.9023
R5485 Transmission_Gate_Layout_9.CLK.t95 Transmission_Gate_Layout_9.CLK.n37 18.9023
R5486 Transmission_Gate_Layout_9.CLK.t79 Transmission_Gate_Layout_9.CLK.n39 18.9023
R5487 Transmission_Gate_Layout_9.CLK.t24 Transmission_Gate_Layout_9.CLK.n41 18.9023
R5488 Transmission_Gate_Layout_9.CLK.n54 Transmission_Gate_Layout_9.CLK.t94 18.9023
R5489 Transmission_Gate_Layout_9.CLK.n55 Transmission_Gate_Layout_9.CLK.t108 18.9023
R5490 Transmission_Gate_Layout_9.CLK.n56 Transmission_Gate_Layout_9.CLK.t54 18.9023
R5491 Transmission_Gate_Layout_9.CLK.n57 Transmission_Gate_Layout_9.CLK.t120 18.9023
R5492 Transmission_Gate_Layout_9.CLK.n58 Transmission_Gate_Layout_9.CLK.t105 18.9023
R5493 Transmission_Gate_Layout_9.CLK.n59 Transmission_Gate_Layout_9.CLK.t51 18.9023
R5494 Transmission_Gate_Layout_9.CLK.n60 Transmission_Gate_Layout_9.CLK.t33 18.9023
R5495 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.CLK.n0 18.6041
R5496 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.CLK.n105 17.6496
R5497 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.CLK.n79 17.6496
R5498 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.CLK.n53 16.4436
R5499 Transmission_Gate_Layout_9.CLK.n27 Transmission_Gate_Layout_9.CLK.n26 16.4376
R5500 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.CLK.n108 7.70137
R5501 Transmission_Gate_Layout_9.CLK.n0 Transmission_Gate_Layout_9.CLK 5.54464
R5502 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.CLK.n109 4.70224
R5503 Transmission_Gate_Layout_9.CLK.n0 Transmission_Gate_Layout_9.CLK 2.44482
R5504 Transmission_Gate_Layout_9.CLK.n0 Transmission_Gate_Layout_9.CLK.n27 2.24392
R5505 Transmission_Gate_Layout_6.VIN.n97 Transmission_Gate_Layout_6.VIN.n96 5.32175
R5506 Transmission_Gate_Layout_6.VIN.n60 Transmission_Gate_Layout_6.VIN.n59 5.21612
R5507 Transmission_Gate_Layout_6.VIN.n63 Transmission_Gate_Layout_6.VIN.t82 4.4609
R5508 Transmission_Gate_Layout_6.VIN.n64 Transmission_Gate_Layout_6.VIN.t79 4.4609
R5509 Transmission_Gate_Layout_6.VIN.n65 Transmission_Gate_Layout_6.VIN.t75 4.4609
R5510 Transmission_Gate_Layout_6.VIN.n61 Transmission_Gate_Layout_6.VIN.n57 4.4609
R5511 Transmission_Gate_Layout_6.VIN.n60 Transmission_Gate_Layout_6.VIN.n58 4.4609
R5512 Transmission_Gate_Layout_6.VIN.n125 Transmission_Gate_Layout_6.VIN.n122 3.90572
R5513 Transmission_Gate_Layout_6.VIN.n117 Transmission_Gate_Layout_6.VIN.n114 3.90572
R5514 Transmission_Gate_Layout_6.VIN.n37 Transmission_Gate_Layout_6.VIN.n34 3.90572
R5515 Transmission_Gate_Layout_6.VIN.n45 Transmission_Gate_Layout_6.VIN.n42 3.90572
R5516 Transmission_Gate_Layout_6.VIN.n55 Transmission_Gate_Layout_6.VIN.n54 3.90572
R5517 Transmission_Gate_Layout_6.VIN.n140 Transmission_Gate_Layout_6.VIN.n139 3.90572
R5518 Transmission_Gate_Layout_6.VIN.n4 Transmission_Gate_Layout_6.VIN.n1 3.84485
R5519 Transmission_Gate_Layout_6.VIN.n85 Transmission_Gate_Layout_6.VIN.n82 3.84485
R5520 Transmission_Gate_Layout_6.VIN.n74 Transmission_Gate_Layout_6.VIN.n73 3.84485
R5521 Transmission_Gate_Layout_6.VIN.n31 Transmission_Gate_Layout_6.VIN.n30 3.84485
R5522 Transmission_Gate_Layout_6.VIN.n14 Transmission_Gate_Layout_6.VIN.n13 3.84485
R5523 Transmission_Gate_Layout_6.VIN.n22 Transmission_Gate_Layout_6.VIN.n21 3.84485
R5524 Transmission_Gate_Layout_6.VIN.n94 Transmission_Gate_Layout_6.VIN.n93 3.3285
R5525 Transmission_Gate_Layout_6.VIN.n92 Transmission_Gate_Layout_6.VIN.n91 3.3285
R5526 Transmission_Gate_Layout_6.VIN.n90 Transmission_Gate_Layout_6.VIN.n89 3.3285
R5527 Transmission_Gate_Layout_6.VIN.n78 Transmission_Gate_Layout_6.VIN.t68 3.3285
R5528 Transmission_Gate_Layout_6.VIN.n79 Transmission_Gate_Layout_6.VIN.t61 3.3285
R5529 Transmission_Gate_Layout_6.VIN.n80 Transmission_Gate_Layout_6.VIN.t50 3.3285
R5530 Transmission_Gate_Layout_6.VIN.n125 Transmission_Gate_Layout_6.VIN.n124 3.1505
R5531 Transmission_Gate_Layout_6.VIN.n128 Transmission_Gate_Layout_6.VIN.n127 3.1505
R5532 Transmission_Gate_Layout_6.VIN.n117 Transmission_Gate_Layout_6.VIN.n116 3.1505
R5533 Transmission_Gate_Layout_6.VIN.n120 Transmission_Gate_Layout_6.VIN.n119 3.1505
R5534 Transmission_Gate_Layout_6.VIN.n37 Transmission_Gate_Layout_6.VIN.n36 3.1505
R5535 Transmission_Gate_Layout_6.VIN.n40 Transmission_Gate_Layout_6.VIN.n39 3.1505
R5536 Transmission_Gate_Layout_6.VIN.n45 Transmission_Gate_Layout_6.VIN.n44 3.1505
R5537 Transmission_Gate_Layout_6.VIN.n48 Transmission_Gate_Layout_6.VIN.n47 3.1505
R5538 Transmission_Gate_Layout_6.VIN.n55 Transmission_Gate_Layout_6.VIN.n52 3.1505
R5539 Transmission_Gate_Layout_6.VIN.n56 Transmission_Gate_Layout_6.VIN.n50 3.1505
R5540 Transmission_Gate_Layout_6.VIN.n130 Transmission_Gate_Layout_6.VIN.n112 3.1505
R5541 Transmission_Gate_Layout_6.VIN.n131 Transmission_Gate_Layout_6.VIN.n110 3.1505
R5542 Transmission_Gate_Layout_6.VIN.n132 Transmission_Gate_Layout_6.VIN.n108 3.1505
R5543 Transmission_Gate_Layout_6.VIN.n140 Transmission_Gate_Layout_6.VIN.n137 3.1505
R5544 Transmission_Gate_Layout_6.VIN.n141 Transmission_Gate_Layout_6.VIN.n135 3.1505
R5545 Transmission_Gate_Layout_6.VIN.n4 Transmission_Gate_Layout_6.VIN.n3 2.6005
R5546 Transmission_Gate_Layout_6.VIN.n7 Transmission_Gate_Layout_6.VIN.n6 2.6005
R5547 Transmission_Gate_Layout_6.VIN.n85 Transmission_Gate_Layout_6.VIN.n84 2.6005
R5548 Transmission_Gate_Layout_6.VIN.n88 Transmission_Gate_Layout_6.VIN.n87 2.6005
R5549 Transmission_Gate_Layout_6.VIN.n74 Transmission_Gate_Layout_6.VIN.n71 2.6005
R5550 Transmission_Gate_Layout_6.VIN.n75 Transmission_Gate_Layout_6.VIN.n69 2.6005
R5551 Transmission_Gate_Layout_6.VIN.n31 Transmission_Gate_Layout_6.VIN.n28 2.6005
R5552 Transmission_Gate_Layout_6.VIN.n32 Transmission_Gate_Layout_6.VIN.n26 2.6005
R5553 Transmission_Gate_Layout_6.VIN.n14 Transmission_Gate_Layout_6.VIN.n11 2.6005
R5554 Transmission_Gate_Layout_6.VIN.n15 Transmission_Gate_Layout_6.VIN.n9 2.6005
R5555 Transmission_Gate_Layout_6.VIN.n22 Transmission_Gate_Layout_6.VIN.n19 2.6005
R5556 Transmission_Gate_Layout_6.VIN.n23 Transmission_Gate_Layout_6.VIN.n17 2.6005
R5557 Transmission_Gate_Layout_6.VIN.n106 Transmission_Gate_Layout_6.VIN.n105 2.6005
R5558 Transmission_Gate_Layout_6.VIN.n103 Transmission_Gate_Layout_6.VIN.n102 2.6005
R5559 Transmission_Gate_Layout_6.VIN.n100 Transmission_Gate_Layout_6.VIN.n99 2.6005
R5560 Transmission_Gate_Layout_6.VIN.n63 Transmission_Gate_Layout_6.VIN.n62 2.47941
R5561 Transmission_Gate_Layout_6.VIN.n96 Transmission_Gate_Layout_6.VIN.n95 1.90239
R5562 Transmission_Gate_Layout_6.VIN.n135 Transmission_Gate_Layout_6.VIN.t45 1.3109
R5563 Transmission_Gate_Layout_6.VIN.n135 Transmission_Gate_Layout_6.VIN.n134 1.3109
R5564 Transmission_Gate_Layout_6.VIN.n137 Transmission_Gate_Layout_6.VIN.t32 1.3109
R5565 Transmission_Gate_Layout_6.VIN.n137 Transmission_Gate_Layout_6.VIN.n136 1.3109
R5566 Transmission_Gate_Layout_6.VIN.n108 Transmission_Gate_Layout_6.VIN.t28 1.3109
R5567 Transmission_Gate_Layout_6.VIN.n108 Transmission_Gate_Layout_6.VIN.n107 1.3109
R5568 Transmission_Gate_Layout_6.VIN.n110 Transmission_Gate_Layout_6.VIN.t38 1.3109
R5569 Transmission_Gate_Layout_6.VIN.n110 Transmission_Gate_Layout_6.VIN.n109 1.3109
R5570 Transmission_Gate_Layout_6.VIN.n112 Transmission_Gate_Layout_6.VIN.t26 1.3109
R5571 Transmission_Gate_Layout_6.VIN.n112 Transmission_Gate_Layout_6.VIN.n111 1.3109
R5572 Transmission_Gate_Layout_6.VIN.n127 Transmission_Gate_Layout_6.VIN.t24 1.3109
R5573 Transmission_Gate_Layout_6.VIN.n127 Transmission_Gate_Layout_6.VIN.n126 1.3109
R5574 Transmission_Gate_Layout_6.VIN.n124 Transmission_Gate_Layout_6.VIN.t35 1.3109
R5575 Transmission_Gate_Layout_6.VIN.n124 Transmission_Gate_Layout_6.VIN.n123 1.3109
R5576 Transmission_Gate_Layout_6.VIN.n122 Transmission_Gate_Layout_6.VIN.t40 1.3109
R5577 Transmission_Gate_Layout_6.VIN.n122 Transmission_Gate_Layout_6.VIN.n121 1.3109
R5578 Transmission_Gate_Layout_6.VIN.n119 Transmission_Gate_Layout_6.VIN.t29 1.3109
R5579 Transmission_Gate_Layout_6.VIN.n119 Transmission_Gate_Layout_6.VIN.n118 1.3109
R5580 Transmission_Gate_Layout_6.VIN.n116 Transmission_Gate_Layout_6.VIN.t44 1.3109
R5581 Transmission_Gate_Layout_6.VIN.n116 Transmission_Gate_Layout_6.VIN.n115 1.3109
R5582 Transmission_Gate_Layout_6.VIN.n114 Transmission_Gate_Layout_6.VIN.t41 1.3109
R5583 Transmission_Gate_Layout_6.VIN.n114 Transmission_Gate_Layout_6.VIN.n113 1.3109
R5584 Transmission_Gate_Layout_6.VIN.n39 Transmission_Gate_Layout_6.VIN.t74 1.3109
R5585 Transmission_Gate_Layout_6.VIN.n39 Transmission_Gate_Layout_6.VIN.n38 1.3109
R5586 Transmission_Gate_Layout_6.VIN.n36 Transmission_Gate_Layout_6.VIN.t78 1.3109
R5587 Transmission_Gate_Layout_6.VIN.n36 Transmission_Gate_Layout_6.VIN.n35 1.3109
R5588 Transmission_Gate_Layout_6.VIN.n34 Transmission_Gate_Layout_6.VIN.t81 1.3109
R5589 Transmission_Gate_Layout_6.VIN.n34 Transmission_Gate_Layout_6.VIN.n33 1.3109
R5590 Transmission_Gate_Layout_6.VIN.n47 Transmission_Gate_Layout_6.VIN.t83 1.3109
R5591 Transmission_Gate_Layout_6.VIN.n47 Transmission_Gate_Layout_6.VIN.n46 1.3109
R5592 Transmission_Gate_Layout_6.VIN.n44 Transmission_Gate_Layout_6.VIN.t72 1.3109
R5593 Transmission_Gate_Layout_6.VIN.n44 Transmission_Gate_Layout_6.VIN.n43 1.3109
R5594 Transmission_Gate_Layout_6.VIN.n42 Transmission_Gate_Layout_6.VIN.t76 1.3109
R5595 Transmission_Gate_Layout_6.VIN.n42 Transmission_Gate_Layout_6.VIN.n41 1.3109
R5596 Transmission_Gate_Layout_6.VIN.n50 Transmission_Gate_Layout_6.VIN.t80 1.3109
R5597 Transmission_Gate_Layout_6.VIN.n50 Transmission_Gate_Layout_6.VIN.n49 1.3109
R5598 Transmission_Gate_Layout_6.VIN.n52 Transmission_Gate_Layout_6.VIN.t77 1.3109
R5599 Transmission_Gate_Layout_6.VIN.n52 Transmission_Gate_Layout_6.VIN.n51 1.3109
R5600 Transmission_Gate_Layout_6.VIN.n54 Transmission_Gate_Layout_6.VIN.t73 1.3109
R5601 Transmission_Gate_Layout_6.VIN.n54 Transmission_Gate_Layout_6.VIN.n53 1.3109
R5602 Transmission_Gate_Layout_6.VIN.n139 Transmission_Gate_Layout_6.VIN.t39 1.3109
R5603 Transmission_Gate_Layout_6.VIN.n139 Transmission_Gate_Layout_6.VIN.n138 1.3109
R5604 Transmission_Gate_Layout_6.VIN.n7 Transmission_Gate_Layout_6.VIN.n4 1.24485
R5605 Transmission_Gate_Layout_6.VIN.n88 Transmission_Gate_Layout_6.VIN.n85 1.24485
R5606 Transmission_Gate_Layout_6.VIN.n92 Transmission_Gate_Layout_6.VIN.n90 1.24485
R5607 Transmission_Gate_Layout_6.VIN.n94 Transmission_Gate_Layout_6.VIN.n92 1.24485
R5608 Transmission_Gate_Layout_6.VIN.n75 Transmission_Gate_Layout_6.VIN.n74 1.24485
R5609 Transmission_Gate_Layout_6.VIN.n32 Transmission_Gate_Layout_6.VIN.n31 1.24485
R5610 Transmission_Gate_Layout_6.VIN.n79 Transmission_Gate_Layout_6.VIN.n78 1.24485
R5611 Transmission_Gate_Layout_6.VIN.n80 Transmission_Gate_Layout_6.VIN.n79 1.24485
R5612 Transmission_Gate_Layout_6.VIN.n15 Transmission_Gate_Layout_6.VIN.n14 1.24485
R5613 Transmission_Gate_Layout_6.VIN.n23 Transmission_Gate_Layout_6.VIN.n22 1.24485
R5614 Transmission_Gate_Layout_6.VIN.n103 Transmission_Gate_Layout_6.VIN.n100 1.24485
R5615 Transmission_Gate_Layout_6.VIN.n106 Transmission_Gate_Layout_6.VIN.n103 1.24485
R5616 Transmission_Gate_Layout_6.VIN.n95 Transmission_Gate_Layout_6.VIN.n94 1.2018
R5617 Transmission_Gate_Layout_6.VIN.n78 Transmission_Gate_Layout_6.VIN.n77 1.2018
R5618 Transmission_Gate_Layout_6.VIN.n24 Transmission_Gate_Layout_6.VIN.n23 1.2018
R5619 Transmission_Gate_Layout_6.VIN.n129 Transmission_Gate_Layout_6.VIN.n128 0.957239
R5620 Transmission_Gate_Layout_6.VIN.n130 Transmission_Gate_Layout_6.VIN.n129 0.957239
R5621 Transmission_Gate_Layout_6.VIN.n62 Transmission_Gate_Layout_6.VIN.n61 0.957239
R5622 Transmission_Gate_Layout_6.VIN.n66 Transmission_Gate_Layout_6.VIN.n65 0.957239
R5623 Transmission_Gate_Layout_6.VIN.n142 Transmission_Gate_Layout_6.VIN.n7 0.806587
R5624 Transmission_Gate_Layout_6.VIN.n133 Transmission_Gate_Layout_6.VIN.n106 0.806587
R5625 Transmission_Gate_Layout_6.VIN.n128 Transmission_Gate_Layout_6.VIN.n125 0.755717
R5626 Transmission_Gate_Layout_6.VIN.n120 Transmission_Gate_Layout_6.VIN.n117 0.755717
R5627 Transmission_Gate_Layout_6.VIN.n40 Transmission_Gate_Layout_6.VIN.n37 0.755717
R5628 Transmission_Gate_Layout_6.VIN.n48 Transmission_Gate_Layout_6.VIN.n45 0.755717
R5629 Transmission_Gate_Layout_6.VIN.n56 Transmission_Gate_Layout_6.VIN.n55 0.755717
R5630 Transmission_Gate_Layout_6.VIN.n61 Transmission_Gate_Layout_6.VIN.n60 0.755717
R5631 Transmission_Gate_Layout_6.VIN.n64 Transmission_Gate_Layout_6.VIN.n63 0.755717
R5632 Transmission_Gate_Layout_6.VIN.n65 Transmission_Gate_Layout_6.VIN.n64 0.755717
R5633 Transmission_Gate_Layout_6.VIN.n132 Transmission_Gate_Layout_6.VIN.n131 0.755717
R5634 Transmission_Gate_Layout_6.VIN.n131 Transmission_Gate_Layout_6.VIN.n130 0.755717
R5635 Transmission_Gate_Layout_6.VIN.n141 Transmission_Gate_Layout_6.VIN.n140 0.755717
R5636 Transmission_Gate_Layout_6.VIN.n96 Transmission_Gate_Layout_6.VIN.n80 0.742022
R5637 Transmission_Gate_Layout_6.VIN.n6 Transmission_Gate_Layout_6.VIN.t8 0.7285
R5638 Transmission_Gate_Layout_6.VIN.n6 Transmission_Gate_Layout_6.VIN.n5 0.7285
R5639 Transmission_Gate_Layout_6.VIN.n3 Transmission_Gate_Layout_6.VIN.t18 0.7285
R5640 Transmission_Gate_Layout_6.VIN.n3 Transmission_Gate_Layout_6.VIN.n2 0.7285
R5641 Transmission_Gate_Layout_6.VIN.n1 Transmission_Gate_Layout_6.VIN.t0 0.7285
R5642 Transmission_Gate_Layout_6.VIN.n1 Transmission_Gate_Layout_6.VIN.n0 0.7285
R5643 Transmission_Gate_Layout_6.VIN.n99 Transmission_Gate_Layout_6.VIN.t16 0.7285
R5644 Transmission_Gate_Layout_6.VIN.n99 Transmission_Gate_Layout_6.VIN.n98 0.7285
R5645 Transmission_Gate_Layout_6.VIN.n102 Transmission_Gate_Layout_6.VIN.t11 0.7285
R5646 Transmission_Gate_Layout_6.VIN.n102 Transmission_Gate_Layout_6.VIN.n101 0.7285
R5647 Transmission_Gate_Layout_6.VIN.n105 Transmission_Gate_Layout_6.VIN.t1 0.7285
R5648 Transmission_Gate_Layout_6.VIN.n105 Transmission_Gate_Layout_6.VIN.n104 0.7285
R5649 Transmission_Gate_Layout_6.VIN.n87 Transmission_Gate_Layout_6.VIN.t52 0.7285
R5650 Transmission_Gate_Layout_6.VIN.n87 Transmission_Gate_Layout_6.VIN.n86 0.7285
R5651 Transmission_Gate_Layout_6.VIN.n84 Transmission_Gate_Layout_6.VIN.t64 0.7285
R5652 Transmission_Gate_Layout_6.VIN.n84 Transmission_Gate_Layout_6.VIN.n83 0.7285
R5653 Transmission_Gate_Layout_6.VIN.n82 Transmission_Gate_Layout_6.VIN.t48 0.7285
R5654 Transmission_Gate_Layout_6.VIN.n82 Transmission_Gate_Layout_6.VIN.n81 0.7285
R5655 Transmission_Gate_Layout_6.VIN.n69 Transmission_Gate_Layout_6.VIN.t71 0.7285
R5656 Transmission_Gate_Layout_6.VIN.n69 Transmission_Gate_Layout_6.VIN.n68 0.7285
R5657 Transmission_Gate_Layout_6.VIN.n71 Transmission_Gate_Layout_6.VIN.t63 0.7285
R5658 Transmission_Gate_Layout_6.VIN.n71 Transmission_Gate_Layout_6.VIN.n70 0.7285
R5659 Transmission_Gate_Layout_6.VIN.n73 Transmission_Gate_Layout_6.VIN.t51 0.7285
R5660 Transmission_Gate_Layout_6.VIN.n73 Transmission_Gate_Layout_6.VIN.n72 0.7285
R5661 Transmission_Gate_Layout_6.VIN.n26 Transmission_Gate_Layout_6.VIN.t56 0.7285
R5662 Transmission_Gate_Layout_6.VIN.n26 Transmission_Gate_Layout_6.VIN.n25 0.7285
R5663 Transmission_Gate_Layout_6.VIN.n28 Transmission_Gate_Layout_6.VIN.t49 0.7285
R5664 Transmission_Gate_Layout_6.VIN.n28 Transmission_Gate_Layout_6.VIN.n27 0.7285
R5665 Transmission_Gate_Layout_6.VIN.n30 Transmission_Gate_Layout_6.VIN.t60 0.7285
R5666 Transmission_Gate_Layout_6.VIN.n30 Transmission_Gate_Layout_6.VIN.n29 0.7285
R5667 Transmission_Gate_Layout_6.VIN.n9 Transmission_Gate_Layout_6.VIN.t5 0.7285
R5668 Transmission_Gate_Layout_6.VIN.n9 Transmission_Gate_Layout_6.VIN.n8 0.7285
R5669 Transmission_Gate_Layout_6.VIN.n11 Transmission_Gate_Layout_6.VIN.t22 0.7285
R5670 Transmission_Gate_Layout_6.VIN.n11 Transmission_Gate_Layout_6.VIN.n10 0.7285
R5671 Transmission_Gate_Layout_6.VIN.n13 Transmission_Gate_Layout_6.VIN.t14 0.7285
R5672 Transmission_Gate_Layout_6.VIN.n13 Transmission_Gate_Layout_6.VIN.n12 0.7285
R5673 Transmission_Gate_Layout_6.VIN.n17 Transmission_Gate_Layout_6.VIN.t6 0.7285
R5674 Transmission_Gate_Layout_6.VIN.n17 Transmission_Gate_Layout_6.VIN.n16 0.7285
R5675 Transmission_Gate_Layout_6.VIN.n19 Transmission_Gate_Layout_6.VIN.t23 0.7285
R5676 Transmission_Gate_Layout_6.VIN.n19 Transmission_Gate_Layout_6.VIN.n18 0.7285
R5677 Transmission_Gate_Layout_6.VIN.n21 Transmission_Gate_Layout_6.VIN.t15 0.7285
R5678 Transmission_Gate_Layout_6.VIN.n21 Transmission_Gate_Layout_6.VIN.n20 0.7285
R5679 Transmission_Gate_Layout_6.VIN.n67 Transmission_Gate_Layout_6.VIN.n66 0.626587
R5680 Transmission_Gate_Layout_6.VIN.n77 Transmission_Gate_Layout_6.VIN.n76 0.626587
R5681 Transmission_Gate_Layout_6.VIN.n142 Transmission_Gate_Layout_6.VIN.n133 0.626587
R5682 Transmission_Gate_Layout_6.VIN.n90 Transmission_Gate_Layout_6.VIN 0.607022
R5683 Transmission_Gate_Layout_6.VIN.n95 Transmission_Gate_Layout_6.VIN.n88 0.575717
R5684 Transmission_Gate_Layout_6.VIN.n76 Transmission_Gate_Layout_6.VIN.n75 0.575717
R5685 Transmission_Gate_Layout_6.VIN.n77 Transmission_Gate_Layout_6.VIN.n32 0.575717
R5686 Transmission_Gate_Layout_6.VIN.n24 Transmission_Gate_Layout_6.VIN.n15 0.575717
R5687 Transmission_Gate_Layout_6.VIN.n97 Transmission_Gate_Layout_6.VIN.n24 0.570002
R5688 Transmission_Gate_Layout_6.VIN.n100 Transmission_Gate_Layout_6.VIN.n97 0.562022
R5689 Transmission_Gate_Layout_6.VIN.n133 Transmission_Gate_Layout_6.VIN.n132 0.428978
R5690 Transmission_Gate_Layout_6.VIN.n142 Transmission_Gate_Layout_6.VIN.n141 0.428978
R5691 Transmission_Gate_Layout_6.VIN.n129 Transmission_Gate_Layout_6.VIN.n120 0.331152
R5692 Transmission_Gate_Layout_6.VIN.n67 Transmission_Gate_Layout_6.VIN.n40 0.331152
R5693 Transmission_Gate_Layout_6.VIN.n66 Transmission_Gate_Layout_6.VIN.n48 0.331152
R5694 Transmission_Gate_Layout_6.VIN.n62 Transmission_Gate_Layout_6.VIN.n56 0.331152
R5695 Transmission_Gate_Layout_6.VIN.n76 Transmission_Gate_Layout_6.VIN.n67 0.239196
R5696 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.VIN.n142 0.192239
R5697 Transmission_Gate_Layout_2.CLKB.n24 Transmission_Gate_Layout_2.CLKB.t18 54.5477
R5698 Transmission_Gate_Layout_2.CLKB.n29 Transmission_Gate_Layout_2.CLKB.t16 38.3255
R5699 Transmission_Gate_Layout_2.CLKB.n28 Transmission_Gate_Layout_2.CLKB.t25 38.3255
R5700 Transmission_Gate_Layout_2.CLKB.n27 Transmission_Gate_Layout_2.CLKB.t14 38.3255
R5701 Transmission_Gate_Layout_2.CLKB.n26 Transmission_Gate_Layout_2.CLKB.t19 38.3255
R5702 Transmission_Gate_Layout_2.CLKB.n25 Transmission_Gate_Layout_2.CLKB.t23 38.3255
R5703 Transmission_Gate_Layout_2.CLKB.n24 Transmission_Gate_Layout_2.CLKB.t13 38.3255
R5704 Transmission_Gate_Layout_2.CLKB.t28 Transmission_Gate_Layout_2.CLKB.n2 37.9344
R5705 Transmission_Gate_Layout_2.CLKB.t12 Transmission_Gate_Layout_2.CLKB.n5 37.9344
R5706 Transmission_Gate_Layout_2.CLKB.t24 Transmission_Gate_Layout_2.CLKB.n8 37.9344
R5707 Transmission_Gate_Layout_2.CLKB.t7 Transmission_Gate_Layout_2.CLKB.n11 37.9344
R5708 Transmission_Gate_Layout_2.CLKB.t11 Transmission_Gate_Layout_2.CLKB.n14 37.9344
R5709 Transmission_Gate_Layout_2.CLKB.t22 Transmission_Gate_Layout_2.CLKB.n17 37.9344
R5710 Transmission_Gate_Layout_2.CLKB.t6 Transmission_Gate_Layout_2.CLKB.n20 37.9344
R5711 Transmission_Gate_Layout_2.CLKB.t17 Transmission_Gate_Layout_2.CLKB.n21 37.9344
R5712 Transmission_Gate_Layout_2.CLKB.n3 Transmission_Gate_Layout_2.CLKB.t28 37.5434
R5713 Transmission_Gate_Layout_2.CLKB.n6 Transmission_Gate_Layout_2.CLKB.t12 37.5434
R5714 Transmission_Gate_Layout_2.CLKB.n9 Transmission_Gate_Layout_2.CLKB.t24 37.5434
R5715 Transmission_Gate_Layout_2.CLKB.n12 Transmission_Gate_Layout_2.CLKB.t7 37.5434
R5716 Transmission_Gate_Layout_2.CLKB.n15 Transmission_Gate_Layout_2.CLKB.t11 37.5434
R5717 Transmission_Gate_Layout_2.CLKB.n18 Transmission_Gate_Layout_2.CLKB.t22 37.5434
R5718 Transmission_Gate_Layout_2.CLKB.n23 Transmission_Gate_Layout_2.CLKB.t6 37.5434
R5719 Transmission_Gate_Layout_2.CLKB.n22 Transmission_Gate_Layout_2.CLKB.t17 37.5434
R5720 Transmission_Gate_Layout_2.CLKB.t16 Transmission_Gate_Layout_2.CLKB.n3 37.413
R5721 Transmission_Gate_Layout_2.CLKB.t25 Transmission_Gate_Layout_2.CLKB.n6 37.413
R5722 Transmission_Gate_Layout_2.CLKB.t14 Transmission_Gate_Layout_2.CLKB.n9 37.413
R5723 Transmission_Gate_Layout_2.CLKB.t19 Transmission_Gate_Layout_2.CLKB.n12 37.413
R5724 Transmission_Gate_Layout_2.CLKB.t23 Transmission_Gate_Layout_2.CLKB.n15 37.413
R5725 Transmission_Gate_Layout_2.CLKB.t13 Transmission_Gate_Layout_2.CLKB.n18 37.413
R5726 Transmission_Gate_Layout_2.CLKB.n22 Transmission_Gate_Layout_2.CLKB.t8 37.413
R5727 Transmission_Gate_Layout_2.CLKB.t18 Transmission_Gate_Layout_2.CLKB.n23 37.413
R5728 Transmission_Gate_Layout_2.CLKB.n21 Transmission_Gate_Layout_2.CLKB.t15 37.0219
R5729 Transmission_Gate_Layout_2.CLKB.n17 Transmission_Gate_Layout_2.CLKB.t20 37.0219
R5730 Transmission_Gate_Layout_2.CLKB.n14 Transmission_Gate_Layout_2.CLKB.t9 37.0219
R5731 Transmission_Gate_Layout_2.CLKB.n11 Transmission_Gate_Layout_2.CLKB.t29 37.0219
R5732 Transmission_Gate_Layout_2.CLKB.n8 Transmission_Gate_Layout_2.CLKB.t21 37.0219
R5733 Transmission_Gate_Layout_2.CLKB.n5 Transmission_Gate_Layout_2.CLKB.t10 37.0219
R5734 Transmission_Gate_Layout_2.CLKB.n2 Transmission_Gate_Layout_2.CLKB.t26 37.0219
R5735 Transmission_Gate_Layout_2.CLKB.n20 Transmission_Gate_Layout_2.CLKB.t27 37.0219
R5736 Transmission_Gate_Layout_2.CLKB.t20 Transmission_Gate_Layout_2.CLKB.n16 35.1969
R5737 Transmission_Gate_Layout_2.CLKB.t9 Transmission_Gate_Layout_2.CLKB.n13 35.1969
R5738 Transmission_Gate_Layout_2.CLKB.t29 Transmission_Gate_Layout_2.CLKB.n10 35.1969
R5739 Transmission_Gate_Layout_2.CLKB.t21 Transmission_Gate_Layout_2.CLKB.n7 35.1969
R5740 Transmission_Gate_Layout_2.CLKB.t10 Transmission_Gate_Layout_2.CLKB.n4 35.1969
R5741 Transmission_Gate_Layout_2.CLKB.t27 Transmission_Gate_Layout_2.CLKB.n19 35.1969
R5742 Transmission_Gate_Layout_2.CLKB Transmission_Gate_Layout_2.CLKB.n29 26.6826
R5743 Transmission_Gate_Layout_2.CLKB.n23 Transmission_Gate_Layout_2.CLKB.n22 19.148
R5744 Transmission_Gate_Layout_2.CLKB.n29 Transmission_Gate_Layout_2.CLKB.n28 16.2227
R5745 Transmission_Gate_Layout_2.CLKB.n28 Transmission_Gate_Layout_2.CLKB.n27 16.2227
R5746 Transmission_Gate_Layout_2.CLKB.n27 Transmission_Gate_Layout_2.CLKB.n26 16.2227
R5747 Transmission_Gate_Layout_2.CLKB.n26 Transmission_Gate_Layout_2.CLKB.n25 16.2227
R5748 Transmission_Gate_Layout_2.CLKB.n25 Transmission_Gate_Layout_2.CLKB.n24 16.2227
R5749 Transmission_Gate_Layout_2.CLKB.n30 Transmission_Gate_Layout_2.CLKB.t3 5.21612
R5750 Transmission_Gate_Layout_2.CLKB.n0 Transmission_Gate_Layout_2.CLKB.t0 4.57285
R5751 Transmission_Gate_Layout_2.CLKB.n31 Transmission_Gate_Layout_2.CLKB.t1 4.4609
R5752 Transmission_Gate_Layout_2.CLKB.n30 Transmission_Gate_Layout_2.CLKB.t5 4.4609
R5753 Transmission_Gate_Layout_2.CLKB.n0 Transmission_Gate_Layout_2.CLKB.t2 3.3285
R5754 Transmission_Gate_Layout_2.CLKB.n1 Transmission_Gate_Layout_2.CLKB.t4 3.3285
R5755 Transmission_Gate_Layout_2.CLKB.n1 Transmission_Gate_Layout_2.CLKB.n0 1.24485
R5756 Transmission_Gate_Layout_2.CLKB.n31 Transmission_Gate_Layout_2.CLKB.n30 0.755717
R5757 Transmission_Gate_Layout_2.CLKB Transmission_Gate_Layout_2.CLKB.n1 0.750969
R5758 Transmission_Gate_Layout_2.CLKB Transmission_Gate_Layout_2.CLKB.n31 0.510317
R5759 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.VIN.n212 8.51067
R5760 Transmission_Gate_Layout_2.VIN.n116 Transmission_Gate_Layout_2.VIN.n115 5.21612
R5761 Transmission_Gate_Layout_2.VIN.n184 Transmission_Gate_Layout_2.VIN.t143 5.21612
R5762 Transmission_Gate_Layout_2.VIN.n119 Transmission_Gate_Layout_2.VIN.t107 4.4609
R5763 Transmission_Gate_Layout_2.VIN.n120 Transmission_Gate_Layout_2.VIN.t111 4.4609
R5764 Transmission_Gate_Layout_2.VIN.n121 Transmission_Gate_Layout_2.VIN.t108 4.4609
R5765 Transmission_Gate_Layout_2.VIN.n117 Transmission_Gate_Layout_2.VIN.n113 4.4609
R5766 Transmission_Gate_Layout_2.VIN.n116 Transmission_Gate_Layout_2.VIN.n114 4.4609
R5767 Transmission_Gate_Layout_2.VIN.n192 Transmission_Gate_Layout_2.VIN.n191 4.4609
R5768 Transmission_Gate_Layout_2.VIN.n190 Transmission_Gate_Layout_2.VIN.n189 4.4609
R5769 Transmission_Gate_Layout_2.VIN.n188 Transmission_Gate_Layout_2.VIN.n187 4.4609
R5770 Transmission_Gate_Layout_2.VIN.n185 Transmission_Gate_Layout_2.VIN.t142 4.4609
R5771 Transmission_Gate_Layout_2.VIN.n184 Transmission_Gate_Layout_2.VIN.t133 4.4609
R5772 Transmission_Gate_Layout_2.VIN.n6 Transmission_Gate_Layout_2.VIN.n5 3.90572
R5773 Transmission_Gate_Layout_2.VIN.n93 Transmission_Gate_Layout_2.VIN.n90 3.90572
R5774 Transmission_Gate_Layout_2.VIN.n101 Transmission_Gate_Layout_2.VIN.n98 3.90572
R5775 Transmission_Gate_Layout_2.VIN.n111 Transmission_Gate_Layout_2.VIN.n110 3.90572
R5776 Transmission_Gate_Layout_2.VIN.n164 Transmission_Gate_Layout_2.VIN.n161 3.90572
R5777 Transmission_Gate_Layout_2.VIN.n182 Transmission_Gate_Layout_2.VIN.n181 3.90572
R5778 Transmission_Gate_Layout_2.VIN.n172 Transmission_Gate_Layout_2.VIN.n169 3.90572
R5779 Transmission_Gate_Layout_2.VIN.n52 Transmission_Gate_Layout_2.VIN.n49 3.90572
R5780 Transmission_Gate_Layout_2.VIN.n44 Transmission_Gate_Layout_2.VIN.n41 3.90572
R5781 Transmission_Gate_Layout_2.VIN.n130 Transmission_Gate_Layout_2.VIN.n129 3.84485
R5782 Transmission_Gate_Layout_2.VIN.n87 Transmission_Gate_Layout_2.VIN.n86 3.84485
R5783 Transmission_Gate_Layout_2.VIN.n77 Transmission_Gate_Layout_2.VIN.n74 3.84485
R5784 Transmission_Gate_Layout_2.VIN.n201 Transmission_Gate_Layout_2.VIN.n200 3.84485
R5785 Transmission_Gate_Layout_2.VIN.n158 Transmission_Gate_Layout_2.VIN.n157 3.84485
R5786 Transmission_Gate_Layout_2.VIN.n148 Transmission_Gate_Layout_2.VIN.n145 3.84485
R5787 Transmission_Gate_Layout_2.VIN.n14 Transmission_Gate_Layout_2.VIN.n13 3.84485
R5788 Transmission_Gate_Layout_2.VIN.n22 Transmission_Gate_Layout_2.VIN.n21 3.84485
R5789 Transmission_Gate_Layout_2.VIN.n65 Transmission_Gate_Layout_2.VIN.n62 3.84485
R5790 Transmission_Gate_Layout_2.VIN.n141 Transmission_Gate_Layout_2.VIN.t45 3.3285
R5791 Transmission_Gate_Layout_2.VIN.n142 Transmission_Gate_Layout_2.VIN.t50 3.3285
R5792 Transmission_Gate_Layout_2.VIN.n143 Transmission_Gate_Layout_2.VIN.t35 3.3285
R5793 Transmission_Gate_Layout_2.VIN.n138 Transmission_Gate_Layout_2.VIN.n72 3.3285
R5794 Transmission_Gate_Layout_2.VIN.n139 Transmission_Gate_Layout_2.VIN.n71 3.3285
R5795 Transmission_Gate_Layout_2.VIN.n140 Transmission_Gate_Layout_2.VIN.n70 3.3285
R5796 Transmission_Gate_Layout_2.VIN.n134 Transmission_Gate_Layout_2.VIN.t113 3.3285
R5797 Transmission_Gate_Layout_2.VIN.n135 Transmission_Gate_Layout_2.VIN.t119 3.3285
R5798 Transmission_Gate_Layout_2.VIN.n136 Transmission_Gate_Layout_2.VIN.t62 3.3285
R5799 Transmission_Gate_Layout_2.VIN.n210 Transmission_Gate_Layout_2.VIN.n209 3.3285
R5800 Transmission_Gate_Layout_2.VIN.n208 Transmission_Gate_Layout_2.VIN.n207 3.3285
R5801 Transmission_Gate_Layout_2.VIN.n206 Transmission_Gate_Layout_2.VIN.n205 3.3285
R5802 Transmission_Gate_Layout_2.VIN.n6 Transmission_Gate_Layout_2.VIN.n3 3.1505
R5803 Transmission_Gate_Layout_2.VIN.n7 Transmission_Gate_Layout_2.VIN.n1 3.1505
R5804 Transmission_Gate_Layout_2.VIN.n93 Transmission_Gate_Layout_2.VIN.n92 3.1505
R5805 Transmission_Gate_Layout_2.VIN.n96 Transmission_Gate_Layout_2.VIN.n95 3.1505
R5806 Transmission_Gate_Layout_2.VIN.n101 Transmission_Gate_Layout_2.VIN.n100 3.1505
R5807 Transmission_Gate_Layout_2.VIN.n104 Transmission_Gate_Layout_2.VIN.n103 3.1505
R5808 Transmission_Gate_Layout_2.VIN.n111 Transmission_Gate_Layout_2.VIN.n108 3.1505
R5809 Transmission_Gate_Layout_2.VIN.n112 Transmission_Gate_Layout_2.VIN.n106 3.1505
R5810 Transmission_Gate_Layout_2.VIN.n164 Transmission_Gate_Layout_2.VIN.n163 3.1505
R5811 Transmission_Gate_Layout_2.VIN.n167 Transmission_Gate_Layout_2.VIN.n166 3.1505
R5812 Transmission_Gate_Layout_2.VIN.n182 Transmission_Gate_Layout_2.VIN.n179 3.1505
R5813 Transmission_Gate_Layout_2.VIN.n183 Transmission_Gate_Layout_2.VIN.n177 3.1505
R5814 Transmission_Gate_Layout_2.VIN.n172 Transmission_Gate_Layout_2.VIN.n171 3.1505
R5815 Transmission_Gate_Layout_2.VIN.n175 Transmission_Gate_Layout_2.VIN.n174 3.1505
R5816 Transmission_Gate_Layout_2.VIN.n52 Transmission_Gate_Layout_2.VIN.n51 3.1505
R5817 Transmission_Gate_Layout_2.VIN.n55 Transmission_Gate_Layout_2.VIN.n54 3.1505
R5818 Transmission_Gate_Layout_2.VIN.n44 Transmission_Gate_Layout_2.VIN.n43 3.1505
R5819 Transmission_Gate_Layout_2.VIN.n47 Transmission_Gate_Layout_2.VIN.n46 3.1505
R5820 Transmission_Gate_Layout_2.VIN.n57 Transmission_Gate_Layout_2.VIN.n39 3.1505
R5821 Transmission_Gate_Layout_2.VIN.n58 Transmission_Gate_Layout_2.VIN.n37 3.1505
R5822 Transmission_Gate_Layout_2.VIN.n59 Transmission_Gate_Layout_2.VIN.n35 3.1505
R5823 Transmission_Gate_Layout_2.VIN.n137 Transmission_Gate_Layout_2.VIN.n136 2.72398
R5824 Transmission_Gate_Layout_2.VIN.n211 Transmission_Gate_Layout_2.VIN.n210 2.72398
R5825 Transmission_Gate_Layout_2.VIN.n130 Transmission_Gate_Layout_2.VIN.n127 2.6005
R5826 Transmission_Gate_Layout_2.VIN.n131 Transmission_Gate_Layout_2.VIN.n125 2.6005
R5827 Transmission_Gate_Layout_2.VIN.n87 Transmission_Gate_Layout_2.VIN.n84 2.6005
R5828 Transmission_Gate_Layout_2.VIN.n88 Transmission_Gate_Layout_2.VIN.n82 2.6005
R5829 Transmission_Gate_Layout_2.VIN.n77 Transmission_Gate_Layout_2.VIN.n76 2.6005
R5830 Transmission_Gate_Layout_2.VIN.n80 Transmission_Gate_Layout_2.VIN.n79 2.6005
R5831 Transmission_Gate_Layout_2.VIN.n201 Transmission_Gate_Layout_2.VIN.n198 2.6005
R5832 Transmission_Gate_Layout_2.VIN.n202 Transmission_Gate_Layout_2.VIN.n196 2.6005
R5833 Transmission_Gate_Layout_2.VIN.n158 Transmission_Gate_Layout_2.VIN.n155 2.6005
R5834 Transmission_Gate_Layout_2.VIN.n159 Transmission_Gate_Layout_2.VIN.n153 2.6005
R5835 Transmission_Gate_Layout_2.VIN.n148 Transmission_Gate_Layout_2.VIN.n147 2.6005
R5836 Transmission_Gate_Layout_2.VIN.n151 Transmission_Gate_Layout_2.VIN.n150 2.6005
R5837 Transmission_Gate_Layout_2.VIN.n14 Transmission_Gate_Layout_2.VIN.n11 2.6005
R5838 Transmission_Gate_Layout_2.VIN.n15 Transmission_Gate_Layout_2.VIN.n9 2.6005
R5839 Transmission_Gate_Layout_2.VIN.n22 Transmission_Gate_Layout_2.VIN.n19 2.6005
R5840 Transmission_Gate_Layout_2.VIN.n23 Transmission_Gate_Layout_2.VIN.n17 2.6005
R5841 Transmission_Gate_Layout_2.VIN.n27 Transmission_Gate_Layout_2.VIN.n26 2.6005
R5842 Transmission_Gate_Layout_2.VIN.n30 Transmission_Gate_Layout_2.VIN.n29 2.6005
R5843 Transmission_Gate_Layout_2.VIN.n33 Transmission_Gate_Layout_2.VIN.n32 2.6005
R5844 Transmission_Gate_Layout_2.VIN.n68 Transmission_Gate_Layout_2.VIN.n67 2.6005
R5845 Transmission_Gate_Layout_2.VIN.n65 Transmission_Gate_Layout_2.VIN.n64 2.6005
R5846 Transmission_Gate_Layout_2.VIN.n119 Transmission_Gate_Layout_2.VIN.n118 2.47941
R5847 Transmission_Gate_Layout_2.VIN.n188 Transmission_Gate_Layout_2.VIN.n186 2.47941
R5848 Transmission_Gate_Layout_2.VIN.n1 Transmission_Gate_Layout_2.VIN.t20 1.3109
R5849 Transmission_Gate_Layout_2.VIN.n1 Transmission_Gate_Layout_2.VIN.n0 1.3109
R5850 Transmission_Gate_Layout_2.VIN.n3 Transmission_Gate_Layout_2.VIN.t12 1.3109
R5851 Transmission_Gate_Layout_2.VIN.n3 Transmission_Gate_Layout_2.VIN.n2 1.3109
R5852 Transmission_Gate_Layout_2.VIN.n5 Transmission_Gate_Layout_2.VIN.t28 1.3109
R5853 Transmission_Gate_Layout_2.VIN.n5 Transmission_Gate_Layout_2.VIN.n4 1.3109
R5854 Transmission_Gate_Layout_2.VIN.n95 Transmission_Gate_Layout_2.VIN.t102 1.3109
R5855 Transmission_Gate_Layout_2.VIN.n95 Transmission_Gate_Layout_2.VIN.n94 1.3109
R5856 Transmission_Gate_Layout_2.VIN.n92 Transmission_Gate_Layout_2.VIN.t109 1.3109
R5857 Transmission_Gate_Layout_2.VIN.n92 Transmission_Gate_Layout_2.VIN.n91 1.3109
R5858 Transmission_Gate_Layout_2.VIN.n90 Transmission_Gate_Layout_2.VIN.t106 1.3109
R5859 Transmission_Gate_Layout_2.VIN.n90 Transmission_Gate_Layout_2.VIN.n89 1.3109
R5860 Transmission_Gate_Layout_2.VIN.n103 Transmission_Gate_Layout_2.VIN.t104 1.3109
R5861 Transmission_Gate_Layout_2.VIN.n103 Transmission_Gate_Layout_2.VIN.n102 1.3109
R5862 Transmission_Gate_Layout_2.VIN.n100 Transmission_Gate_Layout_2.VIN.t105 1.3109
R5863 Transmission_Gate_Layout_2.VIN.n100 Transmission_Gate_Layout_2.VIN.n99 1.3109
R5864 Transmission_Gate_Layout_2.VIN.n98 Transmission_Gate_Layout_2.VIN.t103 1.3109
R5865 Transmission_Gate_Layout_2.VIN.n98 Transmission_Gate_Layout_2.VIN.n97 1.3109
R5866 Transmission_Gate_Layout_2.VIN.n106 Transmission_Gate_Layout_2.VIN.t110 1.3109
R5867 Transmission_Gate_Layout_2.VIN.n106 Transmission_Gate_Layout_2.VIN.n105 1.3109
R5868 Transmission_Gate_Layout_2.VIN.n108 Transmission_Gate_Layout_2.VIN.t101 1.3109
R5869 Transmission_Gate_Layout_2.VIN.n108 Transmission_Gate_Layout_2.VIN.n107 1.3109
R5870 Transmission_Gate_Layout_2.VIN.n110 Transmission_Gate_Layout_2.VIN.t100 1.3109
R5871 Transmission_Gate_Layout_2.VIN.n110 Transmission_Gate_Layout_2.VIN.n109 1.3109
R5872 Transmission_Gate_Layout_2.VIN.n166 Transmission_Gate_Layout_2.VIN.t136 1.3109
R5873 Transmission_Gate_Layout_2.VIN.n166 Transmission_Gate_Layout_2.VIN.n165 1.3109
R5874 Transmission_Gate_Layout_2.VIN.n163 Transmission_Gate_Layout_2.VIN.t140 1.3109
R5875 Transmission_Gate_Layout_2.VIN.n163 Transmission_Gate_Layout_2.VIN.n162 1.3109
R5876 Transmission_Gate_Layout_2.VIN.n161 Transmission_Gate_Layout_2.VIN.t138 1.3109
R5877 Transmission_Gate_Layout_2.VIN.n161 Transmission_Gate_Layout_2.VIN.n160 1.3109
R5878 Transmission_Gate_Layout_2.VIN.n177 Transmission_Gate_Layout_2.VIN.t135 1.3109
R5879 Transmission_Gate_Layout_2.VIN.n177 Transmission_Gate_Layout_2.VIN.n176 1.3109
R5880 Transmission_Gate_Layout_2.VIN.n179 Transmission_Gate_Layout_2.VIN.t137 1.3109
R5881 Transmission_Gate_Layout_2.VIN.n179 Transmission_Gate_Layout_2.VIN.n178 1.3109
R5882 Transmission_Gate_Layout_2.VIN.n181 Transmission_Gate_Layout_2.VIN.t139 1.3109
R5883 Transmission_Gate_Layout_2.VIN.n181 Transmission_Gate_Layout_2.VIN.n180 1.3109
R5884 Transmission_Gate_Layout_2.VIN.n174 Transmission_Gate_Layout_2.VIN.t134 1.3109
R5885 Transmission_Gate_Layout_2.VIN.n174 Transmission_Gate_Layout_2.VIN.n173 1.3109
R5886 Transmission_Gate_Layout_2.VIN.n171 Transmission_Gate_Layout_2.VIN.t132 1.3109
R5887 Transmission_Gate_Layout_2.VIN.n171 Transmission_Gate_Layout_2.VIN.n170 1.3109
R5888 Transmission_Gate_Layout_2.VIN.n169 Transmission_Gate_Layout_2.VIN.t141 1.3109
R5889 Transmission_Gate_Layout_2.VIN.n169 Transmission_Gate_Layout_2.VIN.n168 1.3109
R5890 Transmission_Gate_Layout_2.VIN.n35 Transmission_Gate_Layout_2.VIN.t24 1.3109
R5891 Transmission_Gate_Layout_2.VIN.n35 Transmission_Gate_Layout_2.VIN.n34 1.3109
R5892 Transmission_Gate_Layout_2.VIN.n37 Transmission_Gate_Layout_2.VIN.t18 1.3109
R5893 Transmission_Gate_Layout_2.VIN.n37 Transmission_Gate_Layout_2.VIN.n36 1.3109
R5894 Transmission_Gate_Layout_2.VIN.n39 Transmission_Gate_Layout_2.VIN.t9 1.3109
R5895 Transmission_Gate_Layout_2.VIN.n39 Transmission_Gate_Layout_2.VIN.n38 1.3109
R5896 Transmission_Gate_Layout_2.VIN.n54 Transmission_Gate_Layout_2.VIN.t27 1.3109
R5897 Transmission_Gate_Layout_2.VIN.n54 Transmission_Gate_Layout_2.VIN.n53 1.3109
R5898 Transmission_Gate_Layout_2.VIN.n51 Transmission_Gate_Layout_2.VIN.t11 1.3109
R5899 Transmission_Gate_Layout_2.VIN.n51 Transmission_Gate_Layout_2.VIN.n50 1.3109
R5900 Transmission_Gate_Layout_2.VIN.n49 Transmission_Gate_Layout_2.VIN.t17 1.3109
R5901 Transmission_Gate_Layout_2.VIN.n49 Transmission_Gate_Layout_2.VIN.n48 1.3109
R5902 Transmission_Gate_Layout_2.VIN.n46 Transmission_Gate_Layout_2.VIN.t23 1.3109
R5903 Transmission_Gate_Layout_2.VIN.n46 Transmission_Gate_Layout_2.VIN.n45 1.3109
R5904 Transmission_Gate_Layout_2.VIN.n43 Transmission_Gate_Layout_2.VIN.t7 1.3109
R5905 Transmission_Gate_Layout_2.VIN.n43 Transmission_Gate_Layout_2.VIN.n42 1.3109
R5906 Transmission_Gate_Layout_2.VIN.n41 Transmission_Gate_Layout_2.VIN.t15 1.3109
R5907 Transmission_Gate_Layout_2.VIN.n41 Transmission_Gate_Layout_2.VIN.n40 1.3109
R5908 Transmission_Gate_Layout_2.VIN.n131 Transmission_Gate_Layout_2.VIN.n130 1.24485
R5909 Transmission_Gate_Layout_2.VIN.n88 Transmission_Gate_Layout_2.VIN.n87 1.24485
R5910 Transmission_Gate_Layout_2.VIN.n135 Transmission_Gate_Layout_2.VIN.n134 1.24485
R5911 Transmission_Gate_Layout_2.VIN.n136 Transmission_Gate_Layout_2.VIN.n135 1.24485
R5912 Transmission_Gate_Layout_2.VIN.n80 Transmission_Gate_Layout_2.VIN.n77 1.24485
R5913 Transmission_Gate_Layout_2.VIN.n140 Transmission_Gate_Layout_2.VIN.n139 1.24485
R5914 Transmission_Gate_Layout_2.VIN.n139 Transmission_Gate_Layout_2.VIN.n138 1.24485
R5915 Transmission_Gate_Layout_2.VIN.n142 Transmission_Gate_Layout_2.VIN.n141 1.24485
R5916 Transmission_Gate_Layout_2.VIN.n143 Transmission_Gate_Layout_2.VIN.n142 1.24485
R5917 Transmission_Gate_Layout_2.VIN.n202 Transmission_Gate_Layout_2.VIN.n201 1.24485
R5918 Transmission_Gate_Layout_2.VIN.n159 Transmission_Gate_Layout_2.VIN.n158 1.24485
R5919 Transmission_Gate_Layout_2.VIN.n208 Transmission_Gate_Layout_2.VIN.n206 1.24485
R5920 Transmission_Gate_Layout_2.VIN.n210 Transmission_Gate_Layout_2.VIN.n208 1.24485
R5921 Transmission_Gate_Layout_2.VIN.n151 Transmission_Gate_Layout_2.VIN.n148 1.24485
R5922 Transmission_Gate_Layout_2.VIN.n15 Transmission_Gate_Layout_2.VIN.n14 1.24485
R5923 Transmission_Gate_Layout_2.VIN.n23 Transmission_Gate_Layout_2.VIN.n22 1.24485
R5924 Transmission_Gate_Layout_2.VIN.n30 Transmission_Gate_Layout_2.VIN.n27 1.24485
R5925 Transmission_Gate_Layout_2.VIN.n33 Transmission_Gate_Layout_2.VIN.n30 1.24485
R5926 Transmission_Gate_Layout_2.VIN.n68 Transmission_Gate_Layout_2.VIN.n65 1.24485
R5927 Transmission_Gate_Layout_2.VIN.n134 Transmission_Gate_Layout_2.VIN.n133 1.2018
R5928 Transmission_Gate_Layout_2.VIN.n138 Transmission_Gate_Layout_2.VIN.n137 1.2018
R5929 Transmission_Gate_Layout_2.VIN.n206 Transmission_Gate_Layout_2.VIN.n204 1.2018
R5930 Transmission_Gate_Layout_2.VIN.n24 Transmission_Gate_Layout_2.VIN.n23 1.2018
R5931 Transmission_Gate_Layout_2.VIN.n27 Transmission_Gate_Layout_2.VIN.n24 1.2018
R5932 Transmission_Gate_Layout_2.VIN.n118 Transmission_Gate_Layout_2.VIN.n117 0.957239
R5933 Transmission_Gate_Layout_2.VIN.n122 Transmission_Gate_Layout_2.VIN.n121 0.957239
R5934 Transmission_Gate_Layout_2.VIN.n186 Transmission_Gate_Layout_2.VIN.n185 0.957239
R5935 Transmission_Gate_Layout_2.VIN.n193 Transmission_Gate_Layout_2.VIN.n192 0.957239
R5936 Transmission_Gate_Layout_2.VIN.n56 Transmission_Gate_Layout_2.VIN.n55 0.957239
R5937 Transmission_Gate_Layout_2.VIN.n57 Transmission_Gate_Layout_2.VIN.n56 0.957239
R5938 Transmission_Gate_Layout_2.VIN.n60 Transmission_Gate_Layout_2.VIN.n33 0.806587
R5939 Transmission_Gate_Layout_2.VIN.n69 Transmission_Gate_Layout_2.VIN.n68 0.806587
R5940 Transmission_Gate_Layout_2.VIN.n7 Transmission_Gate_Layout_2.VIN.n6 0.755717
R5941 Transmission_Gate_Layout_2.VIN.n96 Transmission_Gate_Layout_2.VIN.n93 0.755717
R5942 Transmission_Gate_Layout_2.VIN.n104 Transmission_Gate_Layout_2.VIN.n101 0.755717
R5943 Transmission_Gate_Layout_2.VIN.n112 Transmission_Gate_Layout_2.VIN.n111 0.755717
R5944 Transmission_Gate_Layout_2.VIN.n117 Transmission_Gate_Layout_2.VIN.n116 0.755717
R5945 Transmission_Gate_Layout_2.VIN.n120 Transmission_Gate_Layout_2.VIN.n119 0.755717
R5946 Transmission_Gate_Layout_2.VIN.n121 Transmission_Gate_Layout_2.VIN.n120 0.755717
R5947 Transmission_Gate_Layout_2.VIN.n167 Transmission_Gate_Layout_2.VIN.n164 0.755717
R5948 Transmission_Gate_Layout_2.VIN.n183 Transmission_Gate_Layout_2.VIN.n182 0.755717
R5949 Transmission_Gate_Layout_2.VIN.n185 Transmission_Gate_Layout_2.VIN.n184 0.755717
R5950 Transmission_Gate_Layout_2.VIN.n190 Transmission_Gate_Layout_2.VIN.n188 0.755717
R5951 Transmission_Gate_Layout_2.VIN.n192 Transmission_Gate_Layout_2.VIN.n190 0.755717
R5952 Transmission_Gate_Layout_2.VIN.n175 Transmission_Gate_Layout_2.VIN.n172 0.755717
R5953 Transmission_Gate_Layout_2.VIN.n55 Transmission_Gate_Layout_2.VIN.n52 0.755717
R5954 Transmission_Gate_Layout_2.VIN.n47 Transmission_Gate_Layout_2.VIN.n44 0.755717
R5955 Transmission_Gate_Layout_2.VIN.n59 Transmission_Gate_Layout_2.VIN.n58 0.755717
R5956 Transmission_Gate_Layout_2.VIN.n58 Transmission_Gate_Layout_2.VIN.n57 0.755717
R5957 Transmission_Gate_Layout_2.VIN.n67 Transmission_Gate_Layout_2.VIN.t77 0.7285
R5958 Transmission_Gate_Layout_2.VIN.n67 Transmission_Gate_Layout_2.VIN.n66 0.7285
R5959 Transmission_Gate_Layout_2.VIN.n62 Transmission_Gate_Layout_2.VIN.t72 0.7285
R5960 Transmission_Gate_Layout_2.VIN.n62 Transmission_Gate_Layout_2.VIN.n61 0.7285
R5961 Transmission_Gate_Layout_2.VIN.n125 Transmission_Gate_Layout_2.VIN.t61 0.7285
R5962 Transmission_Gate_Layout_2.VIN.n125 Transmission_Gate_Layout_2.VIN.n124 0.7285
R5963 Transmission_Gate_Layout_2.VIN.n127 Transmission_Gate_Layout_2.VIN.t5 0.7285
R5964 Transmission_Gate_Layout_2.VIN.n127 Transmission_Gate_Layout_2.VIN.n126 0.7285
R5965 Transmission_Gate_Layout_2.VIN.n129 Transmission_Gate_Layout_2.VIN.t54 0.7285
R5966 Transmission_Gate_Layout_2.VIN.n129 Transmission_Gate_Layout_2.VIN.n128 0.7285
R5967 Transmission_Gate_Layout_2.VIN.n82 Transmission_Gate_Layout_2.VIN.t60 0.7285
R5968 Transmission_Gate_Layout_2.VIN.n82 Transmission_Gate_Layout_2.VIN.n81 0.7285
R5969 Transmission_Gate_Layout_2.VIN.n84 Transmission_Gate_Layout_2.VIN.t3 0.7285
R5970 Transmission_Gate_Layout_2.VIN.n84 Transmission_Gate_Layout_2.VIN.n83 0.7285
R5971 Transmission_Gate_Layout_2.VIN.n86 Transmission_Gate_Layout_2.VIN.t118 0.7285
R5972 Transmission_Gate_Layout_2.VIN.n86 Transmission_Gate_Layout_2.VIN.n85 0.7285
R5973 Transmission_Gate_Layout_2.VIN.n79 Transmission_Gate_Layout_2.VIN.t59 0.7285
R5974 Transmission_Gate_Layout_2.VIN.n79 Transmission_Gate_Layout_2.VIN.n78 0.7285
R5975 Transmission_Gate_Layout_2.VIN.n76 Transmission_Gate_Layout_2.VIN.t117 0.7285
R5976 Transmission_Gate_Layout_2.VIN.n76 Transmission_Gate_Layout_2.VIN.n75 0.7285
R5977 Transmission_Gate_Layout_2.VIN.n74 Transmission_Gate_Layout_2.VIN.t4 0.7285
R5978 Transmission_Gate_Layout_2.VIN.n74 Transmission_Gate_Layout_2.VIN.n73 0.7285
R5979 Transmission_Gate_Layout_2.VIN.n196 Transmission_Gate_Layout_2.VIN.t32 0.7285
R5980 Transmission_Gate_Layout_2.VIN.n196 Transmission_Gate_Layout_2.VIN.n195 0.7285
R5981 Transmission_Gate_Layout_2.VIN.n198 Transmission_Gate_Layout_2.VIN.t40 0.7285
R5982 Transmission_Gate_Layout_2.VIN.n198 Transmission_Gate_Layout_2.VIN.n197 0.7285
R5983 Transmission_Gate_Layout_2.VIN.n200 Transmission_Gate_Layout_2.VIN.t48 0.7285
R5984 Transmission_Gate_Layout_2.VIN.n200 Transmission_Gate_Layout_2.VIN.n199 0.7285
R5985 Transmission_Gate_Layout_2.VIN.n153 Transmission_Gate_Layout_2.VIN.t39 0.7285
R5986 Transmission_Gate_Layout_2.VIN.n153 Transmission_Gate_Layout_2.VIN.n152 0.7285
R5987 Transmission_Gate_Layout_2.VIN.n155 Transmission_Gate_Layout_2.VIN.t44 0.7285
R5988 Transmission_Gate_Layout_2.VIN.n155 Transmission_Gate_Layout_2.VIN.n154 0.7285
R5989 Transmission_Gate_Layout_2.VIN.n157 Transmission_Gate_Layout_2.VIN.t53 0.7285
R5990 Transmission_Gate_Layout_2.VIN.n157 Transmission_Gate_Layout_2.VIN.n156 0.7285
R5991 Transmission_Gate_Layout_2.VIN.n150 Transmission_Gate_Layout_2.VIN.t41 0.7285
R5992 Transmission_Gate_Layout_2.VIN.n150 Transmission_Gate_Layout_2.VIN.n149 0.7285
R5993 Transmission_Gate_Layout_2.VIN.n147 Transmission_Gate_Layout_2.VIN.t33 0.7285
R5994 Transmission_Gate_Layout_2.VIN.n147 Transmission_Gate_Layout_2.VIN.n146 0.7285
R5995 Transmission_Gate_Layout_2.VIN.n145 Transmission_Gate_Layout_2.VIN.t49 0.7285
R5996 Transmission_Gate_Layout_2.VIN.n145 Transmission_Gate_Layout_2.VIN.n144 0.7285
R5997 Transmission_Gate_Layout_2.VIN.n32 Transmission_Gate_Layout_2.VIN.t75 0.7285
R5998 Transmission_Gate_Layout_2.VIN.n32 Transmission_Gate_Layout_2.VIN.n31 0.7285
R5999 Transmission_Gate_Layout_2.VIN.n29 Transmission_Gate_Layout_2.VIN.t80 0.7285
R6000 Transmission_Gate_Layout_2.VIN.n29 Transmission_Gate_Layout_2.VIN.n28 0.7285
R6001 Transmission_Gate_Layout_2.VIN.n26 Transmission_Gate_Layout_2.VIN.t81 0.7285
R6002 Transmission_Gate_Layout_2.VIN.n26 Transmission_Gate_Layout_2.VIN.n25 0.7285
R6003 Transmission_Gate_Layout_2.VIN.n9 Transmission_Gate_Layout_2.VIN.t76 0.7285
R6004 Transmission_Gate_Layout_2.VIN.n9 Transmission_Gate_Layout_2.VIN.n8 0.7285
R6005 Transmission_Gate_Layout_2.VIN.n11 Transmission_Gate_Layout_2.VIN.t74 0.7285
R6006 Transmission_Gate_Layout_2.VIN.n11 Transmission_Gate_Layout_2.VIN.n10 0.7285
R6007 Transmission_Gate_Layout_2.VIN.n13 Transmission_Gate_Layout_2.VIN.t79 0.7285
R6008 Transmission_Gate_Layout_2.VIN.n13 Transmission_Gate_Layout_2.VIN.n12 0.7285
R6009 Transmission_Gate_Layout_2.VIN.n17 Transmission_Gate_Layout_2.VIN.t73 0.7285
R6010 Transmission_Gate_Layout_2.VIN.n17 Transmission_Gate_Layout_2.VIN.n16 0.7285
R6011 Transmission_Gate_Layout_2.VIN.n19 Transmission_Gate_Layout_2.VIN.t71 0.7285
R6012 Transmission_Gate_Layout_2.VIN.n19 Transmission_Gate_Layout_2.VIN.n18 0.7285
R6013 Transmission_Gate_Layout_2.VIN.n21 Transmission_Gate_Layout_2.VIN.t78 0.7285
R6014 Transmission_Gate_Layout_2.VIN.n21 Transmission_Gate_Layout_2.VIN.n20 0.7285
R6015 Transmission_Gate_Layout_2.VIN.n64 Transmission_Gate_Layout_2.VIN.t82 0.7285
R6016 Transmission_Gate_Layout_2.VIN.n64 Transmission_Gate_Layout_2.VIN.n63 0.7285
R6017 Transmission_Gate_Layout_2.VIN.n123 Transmission_Gate_Layout_2.VIN.n122 0.626587
R6018 Transmission_Gate_Layout_2.VIN.n133 Transmission_Gate_Layout_2.VIN.n132 0.626587
R6019 Transmission_Gate_Layout_2.VIN.n194 Transmission_Gate_Layout_2.VIN.n193 0.626587
R6020 Transmission_Gate_Layout_2.VIN.n204 Transmission_Gate_Layout_2.VIN.n203 0.626587
R6021 Transmission_Gate_Layout_2.VIN.n69 Transmission_Gate_Layout_2.VIN.n60 0.626587
R6022 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.VIN.n140 0.607022
R6023 Transmission_Gate_Layout_2.VIN.n141 Transmission_Gate_Layout_2.VIN 0.607022
R6024 Transmission_Gate_Layout_2.VIN.n212 Transmission_Gate_Layout_2.VIN.n211 0.597239
R6025 Transmission_Gate_Layout_2.VIN.n132 Transmission_Gate_Layout_2.VIN.n131 0.575717
R6026 Transmission_Gate_Layout_2.VIN.n133 Transmission_Gate_Layout_2.VIN.n88 0.575717
R6027 Transmission_Gate_Layout_2.VIN.n137 Transmission_Gate_Layout_2.VIN.n80 0.575717
R6028 Transmission_Gate_Layout_2.VIN.n203 Transmission_Gate_Layout_2.VIN.n202 0.575717
R6029 Transmission_Gate_Layout_2.VIN.n204 Transmission_Gate_Layout_2.VIN.n159 0.575717
R6030 Transmission_Gate_Layout_2.VIN.n211 Transmission_Gate_Layout_2.VIN.n151 0.575717
R6031 Transmission_Gate_Layout_2.VIN.n24 Transmission_Gate_Layout_2.VIN.n15 0.575717
R6032 Transmission_Gate_Layout_2.VIN.n212 Transmission_Gate_Layout_2.VIN.n143 0.54637
R6033 Transmission_Gate_Layout_2.VIN.n69 Transmission_Gate_Layout_2.VIN.n7 0.428978
R6034 Transmission_Gate_Layout_2.VIN.n60 Transmission_Gate_Layout_2.VIN.n59 0.428978
R6035 Transmission_Gate_Layout_2.VIN.n123 Transmission_Gate_Layout_2.VIN.n96 0.331152
R6036 Transmission_Gate_Layout_2.VIN.n122 Transmission_Gate_Layout_2.VIN.n104 0.331152
R6037 Transmission_Gate_Layout_2.VIN.n118 Transmission_Gate_Layout_2.VIN.n112 0.331152
R6038 Transmission_Gate_Layout_2.VIN.n194 Transmission_Gate_Layout_2.VIN.n167 0.331152
R6039 Transmission_Gate_Layout_2.VIN.n186 Transmission_Gate_Layout_2.VIN.n183 0.331152
R6040 Transmission_Gate_Layout_2.VIN.n193 Transmission_Gate_Layout_2.VIN.n175 0.331152
R6041 Transmission_Gate_Layout_2.VIN.n56 Transmission_Gate_Layout_2.VIN.n47 0.331152
R6042 Transmission_Gate_Layout_2.VIN.n132 Transmission_Gate_Layout_2.VIN.n123 0.239196
R6043 Transmission_Gate_Layout_2.VIN.n203 Transmission_Gate_Layout_2.VIN.n194 0.239196
R6044 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.VIN.n69 0.192239
R6045 Transmission_Gate_Layout_13.VIN.n188 Transmission_Gate_Layout_13.VIN.n173 11.4073
R6046 Transmission_Gate_Layout_13.VIN.n46 Transmission_Gate_Layout_13.VIN.t17 5.21612
R6047 Transmission_Gate_Layout_13.VIN.n184 Transmission_Gate_Layout_13.VIN.n182 5.21612
R6048 Transmission_Gate_Layout_13.VIN.n51 Transmission_Gate_Layout_13.VIN.n35 4.4609
R6049 Transmission_Gate_Layout_13.VIN.n50 Transmission_Gate_Layout_13.VIN.n36 4.4609
R6050 Transmission_Gate_Layout_13.VIN.n49 Transmission_Gate_Layout_13.VIN.n37 4.4609
R6051 Transmission_Gate_Layout_13.VIN.n47 Transmission_Gate_Layout_13.VIN.t25 4.4609
R6052 Transmission_Gate_Layout_13.VIN.n46 Transmission_Gate_Layout_13.VIN.t34 4.4609
R6053 Transmission_Gate_Layout_13.VIN.n189 Transmission_Gate_Layout_13.VIN.t116 4.4609
R6054 Transmission_Gate_Layout_13.VIN.n190 Transmission_Gate_Layout_13.VIN.t112 4.4609
R6055 Transmission_Gate_Layout_13.VIN.n191 Transmission_Gate_Layout_13.VIN.t103 4.4609
R6056 Transmission_Gate_Layout_13.VIN.n186 Transmission_Gate_Layout_13.VIN.n185 4.4609
R6057 Transmission_Gate_Layout_13.VIN.n184 Transmission_Gate_Layout_13.VIN.n183 4.4609
R6058 Transmission_Gate_Layout_13.VIN.n25 Transmission_Gate_Layout_13.VIN.n24 3.90572
R6059 Transmission_Gate_Layout_13.VIN.n33 Transmission_Gate_Layout_13.VIN.n32 3.90572
R6060 Transmission_Gate_Layout_13.VIN.n42 Transmission_Gate_Layout_13.VIN.n39 3.90572
R6061 Transmission_Gate_Layout_13.VIN.n93 Transmission_Gate_Layout_13.VIN.n92 3.90572
R6062 Transmission_Gate_Layout_13.VIN.n160 Transmission_Gate_Layout_13.VIN.n157 3.90572
R6063 Transmission_Gate_Layout_13.VIN.n168 Transmission_Gate_Layout_13.VIN.n165 3.90572
R6064 Transmission_Gate_Layout_13.VIN.n143 Transmission_Gate_Layout_13.VIN.n142 3.90572
R6065 Transmission_Gate_Layout_13.VIN.n178 Transmission_Gate_Layout_13.VIN.n175 3.90572
R6066 Transmission_Gate_Layout_13.VIN.n101 Transmission_Gate_Layout_13.VIN.n100 3.90572
R6067 Transmission_Gate_Layout_13.VIN.n7 Transmission_Gate_Layout_13.VIN.n4 3.84485
R6068 Transmission_Gate_Layout_13.VIN.n15 Transmission_Gate_Layout_13.VIN.n12 3.84485
R6069 Transmission_Gate_Layout_13.VIN.n117 Transmission_Gate_Layout_13.VIN.n116 3.84485
R6070 Transmission_Gate_Layout_13.VIN.n109 Transmission_Gate_Layout_13.VIN.n108 3.84485
R6071 Transmission_Gate_Layout_13.VIN.n133 Transmission_Gate_Layout_13.VIN.n130 3.84485
R6072 Transmission_Gate_Layout_13.VIN.n83 Transmission_Gate_Layout_13.VIN.n80 3.84485
R6073 Transmission_Gate_Layout_13.VIN.n75 Transmission_Gate_Layout_13.VIN.n72 3.84485
R6074 Transmission_Gate_Layout_13.VIN.n205 Transmission_Gate_Layout_13.VIN.n204 3.84485
R6075 Transmission_Gate_Layout_13.VIN.n65 Transmission_Gate_Layout_13.VIN.n62 3.84485
R6076 Transmission_Gate_Layout_13.VIN.n58 Transmission_Gate_Layout_13.VIN.n0 3.3285
R6077 Transmission_Gate_Layout_13.VIN.n57 Transmission_Gate_Layout_13.VIN.n1 3.3285
R6078 Transmission_Gate_Layout_13.VIN.n56 Transmission_Gate_Layout_13.VIN.n2 3.3285
R6079 Transmission_Gate_Layout_13.VIN.n70 Transmission_Gate_Layout_13.VIN.t96 3.3285
R6080 Transmission_Gate_Layout_13.VIN.n69 Transmission_Gate_Layout_13.VIN.t87 3.3285
R6081 Transmission_Gate_Layout_13.VIN.n68 Transmission_Gate_Layout_13.VIN.t89 3.3285
R6082 Transmission_Gate_Layout_13.VIN.n209 Transmission_Gate_Layout_13.VIN.n208 3.3285
R6083 Transmission_Gate_Layout_13.VIN.n211 Transmission_Gate_Layout_13.VIN.n210 3.3285
R6084 Transmission_Gate_Layout_13.VIN.n213 Transmission_Gate_Layout_13.VIN.n212 3.3285
R6085 Transmission_Gate_Layout_13.VIN.n196 Transmission_Gate_Layout_13.VIN.t125 3.3285
R6086 Transmission_Gate_Layout_13.VIN.n197 Transmission_Gate_Layout_13.VIN.t138 3.3285
R6087 Transmission_Gate_Layout_13.VIN.n198 Transmission_Gate_Layout_13.VIN.t136 3.3285
R6088 Transmission_Gate_Layout_13.VIN.n25 Transmission_Gate_Layout_13.VIN.n22 3.1505
R6089 Transmission_Gate_Layout_13.VIN.n26 Transmission_Gate_Layout_13.VIN.n20 3.1505
R6090 Transmission_Gate_Layout_13.VIN.n33 Transmission_Gate_Layout_13.VIN.n30 3.1505
R6091 Transmission_Gate_Layout_13.VIN.n34 Transmission_Gate_Layout_13.VIN.n28 3.1505
R6092 Transmission_Gate_Layout_13.VIN.n42 Transmission_Gate_Layout_13.VIN.n41 3.1505
R6093 Transmission_Gate_Layout_13.VIN.n45 Transmission_Gate_Layout_13.VIN.n44 3.1505
R6094 Transmission_Gate_Layout_13.VIN.n93 Transmission_Gate_Layout_13.VIN.n90 3.1505
R6095 Transmission_Gate_Layout_13.VIN.n94 Transmission_Gate_Layout_13.VIN.n88 3.1505
R6096 Transmission_Gate_Layout_13.VIN.n160 Transmission_Gate_Layout_13.VIN.n159 3.1505
R6097 Transmission_Gate_Layout_13.VIN.n163 Transmission_Gate_Layout_13.VIN.n162 3.1505
R6098 Transmission_Gate_Layout_13.VIN.n168 Transmission_Gate_Layout_13.VIN.n167 3.1505
R6099 Transmission_Gate_Layout_13.VIN.n171 Transmission_Gate_Layout_13.VIN.n170 3.1505
R6100 Transmission_Gate_Layout_13.VIN.n143 Transmission_Gate_Layout_13.VIN.n140 3.1505
R6101 Transmission_Gate_Layout_13.VIN.n144 Transmission_Gate_Layout_13.VIN.n138 3.1505
R6102 Transmission_Gate_Layout_13.VIN.n155 Transmission_Gate_Layout_13.VIN.n154 3.1505
R6103 Transmission_Gate_Layout_13.VIN.n152 Transmission_Gate_Layout_13.VIN.n151 3.1505
R6104 Transmission_Gate_Layout_13.VIN.n149 Transmission_Gate_Layout_13.VIN.n148 3.1505
R6105 Transmission_Gate_Layout_13.VIN.n178 Transmission_Gate_Layout_13.VIN.n177 3.1505
R6106 Transmission_Gate_Layout_13.VIN.n181 Transmission_Gate_Layout_13.VIN.n180 3.1505
R6107 Transmission_Gate_Layout_13.VIN.n101 Transmission_Gate_Layout_13.VIN.n98 3.1505
R6108 Transmission_Gate_Layout_13.VIN.n102 Transmission_Gate_Layout_13.VIN.n96 3.1505
R6109 Transmission_Gate_Layout_13.VIN.n67 Transmission_Gate_Layout_13.VIN.n58 2.72398
R6110 Transmission_Gate_Layout_13.VIN.n207 Transmission_Gate_Layout_13.VIN.n198 2.72398
R6111 Transmission_Gate_Layout_13.VIN.n7 Transmission_Gate_Layout_13.VIN.n6 2.6005
R6112 Transmission_Gate_Layout_13.VIN.n10 Transmission_Gate_Layout_13.VIN.n9 2.6005
R6113 Transmission_Gate_Layout_13.VIN.n15 Transmission_Gate_Layout_13.VIN.n14 2.6005
R6114 Transmission_Gate_Layout_13.VIN.n18 Transmission_Gate_Layout_13.VIN.n17 2.6005
R6115 Transmission_Gate_Layout_13.VIN.n117 Transmission_Gate_Layout_13.VIN.n114 2.6005
R6116 Transmission_Gate_Layout_13.VIN.n118 Transmission_Gate_Layout_13.VIN.n112 2.6005
R6117 Transmission_Gate_Layout_13.VIN.n109 Transmission_Gate_Layout_13.VIN.n106 2.6005
R6118 Transmission_Gate_Layout_13.VIN.n110 Transmission_Gate_Layout_13.VIN.n104 2.6005
R6119 Transmission_Gate_Layout_13.VIN.n128 Transmission_Gate_Layout_13.VIN.n127 2.6005
R6120 Transmission_Gate_Layout_13.VIN.n125 Transmission_Gate_Layout_13.VIN.n124 2.6005
R6121 Transmission_Gate_Layout_13.VIN.n122 Transmission_Gate_Layout_13.VIN.n121 2.6005
R6122 Transmission_Gate_Layout_13.VIN.n133 Transmission_Gate_Layout_13.VIN.n132 2.6005
R6123 Transmission_Gate_Layout_13.VIN.n136 Transmission_Gate_Layout_13.VIN.n135 2.6005
R6124 Transmission_Gate_Layout_13.VIN.n83 Transmission_Gate_Layout_13.VIN.n82 2.6005
R6125 Transmission_Gate_Layout_13.VIN.n86 Transmission_Gate_Layout_13.VIN.n85 2.6005
R6126 Transmission_Gate_Layout_13.VIN.n75 Transmission_Gate_Layout_13.VIN.n74 2.6005
R6127 Transmission_Gate_Layout_13.VIN.n78 Transmission_Gate_Layout_13.VIN.n77 2.6005
R6128 Transmission_Gate_Layout_13.VIN.n205 Transmission_Gate_Layout_13.VIN.n202 2.6005
R6129 Transmission_Gate_Layout_13.VIN.n206 Transmission_Gate_Layout_13.VIN.n200 2.6005
R6130 Transmission_Gate_Layout_13.VIN.n66 Transmission_Gate_Layout_13.VIN.n60 2.6005
R6131 Transmission_Gate_Layout_13.VIN.n65 Transmission_Gate_Layout_13.VIN.n64 2.6005
R6132 Transmission_Gate_Layout_13.VIN.n49 Transmission_Gate_Layout_13.VIN.n48 2.47941
R6133 Transmission_Gate_Layout_13.VIN.n188 Transmission_Gate_Layout_13.VIN.n187 2.10376
R6134 Transmission_Gate_Layout_13.VIN.n20 Transmission_Gate_Layout_13.VIN.t30 1.3109
R6135 Transmission_Gate_Layout_13.VIN.n20 Transmission_Gate_Layout_13.VIN.n19 1.3109
R6136 Transmission_Gate_Layout_13.VIN.n22 Transmission_Gate_Layout_13.VIN.t22 1.3109
R6137 Transmission_Gate_Layout_13.VIN.n22 Transmission_Gate_Layout_13.VIN.n21 1.3109
R6138 Transmission_Gate_Layout_13.VIN.n24 Transmission_Gate_Layout_13.VIN.t38 1.3109
R6139 Transmission_Gate_Layout_13.VIN.n24 Transmission_Gate_Layout_13.VIN.n23 1.3109
R6140 Transmission_Gate_Layout_13.VIN.n28 Transmission_Gate_Layout_13.VIN.t35 1.3109
R6141 Transmission_Gate_Layout_13.VIN.n28 Transmission_Gate_Layout_13.VIN.n27 1.3109
R6142 Transmission_Gate_Layout_13.VIN.n30 Transmission_Gate_Layout_13.VIN.t28 1.3109
R6143 Transmission_Gate_Layout_13.VIN.n30 Transmission_Gate_Layout_13.VIN.n29 1.3109
R6144 Transmission_Gate_Layout_13.VIN.n32 Transmission_Gate_Layout_13.VIN.t19 1.3109
R6145 Transmission_Gate_Layout_13.VIN.n32 Transmission_Gate_Layout_13.VIN.n31 1.3109
R6146 Transmission_Gate_Layout_13.VIN.n44 Transmission_Gate_Layout_13.VIN.t31 1.3109
R6147 Transmission_Gate_Layout_13.VIN.n44 Transmission_Gate_Layout_13.VIN.n43 1.3109
R6148 Transmission_Gate_Layout_13.VIN.n41 Transmission_Gate_Layout_13.VIN.t15 1.3109
R6149 Transmission_Gate_Layout_13.VIN.n41 Transmission_Gate_Layout_13.VIN.n40 1.3109
R6150 Transmission_Gate_Layout_13.VIN.n39 Transmission_Gate_Layout_13.VIN.t23 1.3109
R6151 Transmission_Gate_Layout_13.VIN.n39 Transmission_Gate_Layout_13.VIN.n38 1.3109
R6152 Transmission_Gate_Layout_13.VIN.n88 Transmission_Gate_Layout_13.VIN.t143 1.3109
R6153 Transmission_Gate_Layout_13.VIN.n88 Transmission_Gate_Layout_13.VIN.n87 1.3109
R6154 Transmission_Gate_Layout_13.VIN.n90 Transmission_Gate_Layout_13.VIN.t115 1.3109
R6155 Transmission_Gate_Layout_13.VIN.n90 Transmission_Gate_Layout_13.VIN.n89 1.3109
R6156 Transmission_Gate_Layout_13.VIN.n92 Transmission_Gate_Layout_13.VIN.t104 1.3109
R6157 Transmission_Gate_Layout_13.VIN.n92 Transmission_Gate_Layout_13.VIN.n91 1.3109
R6158 Transmission_Gate_Layout_13.VIN.n162 Transmission_Gate_Layout_13.VIN.t8 1.3109
R6159 Transmission_Gate_Layout_13.VIN.n162 Transmission_Gate_Layout_13.VIN.n161 1.3109
R6160 Transmission_Gate_Layout_13.VIN.n159 Transmission_Gate_Layout_13.VIN.t46 1.3109
R6161 Transmission_Gate_Layout_13.VIN.n159 Transmission_Gate_Layout_13.VIN.n158 1.3109
R6162 Transmission_Gate_Layout_13.VIN.n157 Transmission_Gate_Layout_13.VIN.t53 1.3109
R6163 Transmission_Gate_Layout_13.VIN.n157 Transmission_Gate_Layout_13.VIN.n156 1.3109
R6164 Transmission_Gate_Layout_13.VIN.n170 Transmission_Gate_Layout_13.VIN.t44 1.3109
R6165 Transmission_Gate_Layout_13.VIN.n170 Transmission_Gate_Layout_13.VIN.n169 1.3109
R6166 Transmission_Gate_Layout_13.VIN.n167 Transmission_Gate_Layout_13.VIN.t52 1.3109
R6167 Transmission_Gate_Layout_13.VIN.n167 Transmission_Gate_Layout_13.VIN.n166 1.3109
R6168 Transmission_Gate_Layout_13.VIN.n165 Transmission_Gate_Layout_13.VIN.t5 1.3109
R6169 Transmission_Gate_Layout_13.VIN.n165 Transmission_Gate_Layout_13.VIN.n164 1.3109
R6170 Transmission_Gate_Layout_13.VIN.n148 Transmission_Gate_Layout_13.VIN.t50 1.3109
R6171 Transmission_Gate_Layout_13.VIN.n148 Transmission_Gate_Layout_13.VIN.n147 1.3109
R6172 Transmission_Gate_Layout_13.VIN.n151 Transmission_Gate_Layout_13.VIN.t43 1.3109
R6173 Transmission_Gate_Layout_13.VIN.n151 Transmission_Gate_Layout_13.VIN.n150 1.3109
R6174 Transmission_Gate_Layout_13.VIN.n154 Transmission_Gate_Layout_13.VIN.t6 1.3109
R6175 Transmission_Gate_Layout_13.VIN.n154 Transmission_Gate_Layout_13.VIN.n153 1.3109
R6176 Transmission_Gate_Layout_13.VIN.n138 Transmission_Gate_Layout_13.VIN.t7 1.3109
R6177 Transmission_Gate_Layout_13.VIN.n138 Transmission_Gate_Layout_13.VIN.n137 1.3109
R6178 Transmission_Gate_Layout_13.VIN.n140 Transmission_Gate_Layout_13.VIN.t54 1.3109
R6179 Transmission_Gate_Layout_13.VIN.n140 Transmission_Gate_Layout_13.VIN.n139 1.3109
R6180 Transmission_Gate_Layout_13.VIN.n142 Transmission_Gate_Layout_13.VIN.t45 1.3109
R6181 Transmission_Gate_Layout_13.VIN.n142 Transmission_Gate_Layout_13.VIN.n141 1.3109
R6182 Transmission_Gate_Layout_13.VIN.n180 Transmission_Gate_Layout_13.VIN.t109 1.3109
R6183 Transmission_Gate_Layout_13.VIN.n180 Transmission_Gate_Layout_13.VIN.n179 1.3109
R6184 Transmission_Gate_Layout_13.VIN.n177 Transmission_Gate_Layout_13.VIN.t1 1.3109
R6185 Transmission_Gate_Layout_13.VIN.n177 Transmission_Gate_Layout_13.VIN.n176 1.3109
R6186 Transmission_Gate_Layout_13.VIN.n175 Transmission_Gate_Layout_13.VIN.t101 1.3109
R6187 Transmission_Gate_Layout_13.VIN.n175 Transmission_Gate_Layout_13.VIN.n174 1.3109
R6188 Transmission_Gate_Layout_13.VIN.n96 Transmission_Gate_Layout_13.VIN.t0 1.3109
R6189 Transmission_Gate_Layout_13.VIN.n96 Transmission_Gate_Layout_13.VIN.n95 1.3109
R6190 Transmission_Gate_Layout_13.VIN.n98 Transmission_Gate_Layout_13.VIN.t110 1.3109
R6191 Transmission_Gate_Layout_13.VIN.n98 Transmission_Gate_Layout_13.VIN.n97 1.3109
R6192 Transmission_Gate_Layout_13.VIN.n100 Transmission_Gate_Layout_13.VIN.t102 1.3109
R6193 Transmission_Gate_Layout_13.VIN.n100 Transmission_Gate_Layout_13.VIN.n99 1.3109
R6194 Transmission_Gate_Layout_13.VIN.n10 Transmission_Gate_Layout_13.VIN.n7 1.24485
R6195 Transmission_Gate_Layout_13.VIN.n18 Transmission_Gate_Layout_13.VIN.n15 1.24485
R6196 Transmission_Gate_Layout_13.VIN.n58 Transmission_Gate_Layout_13.VIN.n57 1.24485
R6197 Transmission_Gate_Layout_13.VIN.n57 Transmission_Gate_Layout_13.VIN.n56 1.24485
R6198 Transmission_Gate_Layout_13.VIN.n118 Transmission_Gate_Layout_13.VIN.n117 1.24485
R6199 Transmission_Gate_Layout_13.VIN.n110 Transmission_Gate_Layout_13.VIN.n109 1.24485
R6200 Transmission_Gate_Layout_13.VIN.n125 Transmission_Gate_Layout_13.VIN.n122 1.24485
R6201 Transmission_Gate_Layout_13.VIN.n128 Transmission_Gate_Layout_13.VIN.n125 1.24485
R6202 Transmission_Gate_Layout_13.VIN.n136 Transmission_Gate_Layout_13.VIN.n133 1.24485
R6203 Transmission_Gate_Layout_13.VIN.n86 Transmission_Gate_Layout_13.VIN.n83 1.24485
R6204 Transmission_Gate_Layout_13.VIN.n78 Transmission_Gate_Layout_13.VIN.n75 1.24485
R6205 Transmission_Gate_Layout_13.VIN.n198 Transmission_Gate_Layout_13.VIN.n197 1.24485
R6206 Transmission_Gate_Layout_13.VIN.n197 Transmission_Gate_Layout_13.VIN.n196 1.24485
R6207 Transmission_Gate_Layout_13.VIN.n206 Transmission_Gate_Layout_13.VIN.n205 1.24485
R6208 Transmission_Gate_Layout_13.VIN.n211 Transmission_Gate_Layout_13.VIN.n209 1.24485
R6209 Transmission_Gate_Layout_13.VIN.n213 Transmission_Gate_Layout_13.VIN.n211 1.24485
R6210 Transmission_Gate_Layout_13.VIN.n69 Transmission_Gate_Layout_13.VIN.n68 1.24485
R6211 Transmission_Gate_Layout_13.VIN.n70 Transmission_Gate_Layout_13.VIN.n69 1.24485
R6212 Transmission_Gate_Layout_13.VIN.n66 Transmission_Gate_Layout_13.VIN.n65 1.24485
R6213 Transmission_Gate_Layout_13.VIN.n56 Transmission_Gate_Layout_13.VIN.n55 1.2018
R6214 Transmission_Gate_Layout_13.VIN.n119 Transmission_Gate_Layout_13.VIN.n118 1.2018
R6215 Transmission_Gate_Layout_13.VIN.n122 Transmission_Gate_Layout_13.VIN.n119 1.2018
R6216 Transmission_Gate_Layout_13.VIN.n196 Transmission_Gate_Layout_13.VIN.n195 1.2018
R6217 Transmission_Gate_Layout_13.VIN.n209 Transmission_Gate_Layout_13.VIN.n207 1.2018
R6218 Transmission_Gate_Layout_13.VIN.n68 Transmission_Gate_Layout_13.VIN.n67 1.2018
R6219 Transmission_Gate_Layout_13.VIN.n48 Transmission_Gate_Layout_13.VIN.n47 0.957239
R6220 Transmission_Gate_Layout_13.VIN.n52 Transmission_Gate_Layout_13.VIN.n51 0.957239
R6221 Transmission_Gate_Layout_13.VIN.n172 Transmission_Gate_Layout_13.VIN.n171 0.957239
R6222 Transmission_Gate_Layout_13.VIN.n187 Transmission_Gate_Layout_13.VIN.n186 0.957239
R6223 Transmission_Gate_Layout_13.VIN.n192 Transmission_Gate_Layout_13.VIN.n191 0.957239
R6224 Transmission_Gate_Layout_13.VIN.n146 Transmission_Gate_Layout_13.VIN.n128 0.806587
R6225 Transmission_Gate_Layout_13.VIN.n145 Transmission_Gate_Layout_13.VIN.n136 0.806587
R6226 Transmission_Gate_Layout_13.VIN.n26 Transmission_Gate_Layout_13.VIN.n25 0.755717
R6227 Transmission_Gate_Layout_13.VIN.n34 Transmission_Gate_Layout_13.VIN.n33 0.755717
R6228 Transmission_Gate_Layout_13.VIN.n45 Transmission_Gate_Layout_13.VIN.n42 0.755717
R6229 Transmission_Gate_Layout_13.VIN.n47 Transmission_Gate_Layout_13.VIN.n46 0.755717
R6230 Transmission_Gate_Layout_13.VIN.n51 Transmission_Gate_Layout_13.VIN.n50 0.755717
R6231 Transmission_Gate_Layout_13.VIN.n50 Transmission_Gate_Layout_13.VIN.n49 0.755717
R6232 Transmission_Gate_Layout_13.VIN.n94 Transmission_Gate_Layout_13.VIN.n93 0.755717
R6233 Transmission_Gate_Layout_13.VIN.n163 Transmission_Gate_Layout_13.VIN.n160 0.755717
R6234 Transmission_Gate_Layout_13.VIN.n171 Transmission_Gate_Layout_13.VIN.n168 0.755717
R6235 Transmission_Gate_Layout_13.VIN.n144 Transmission_Gate_Layout_13.VIN.n143 0.755717
R6236 Transmission_Gate_Layout_13.VIN.n152 Transmission_Gate_Layout_13.VIN.n149 0.755717
R6237 Transmission_Gate_Layout_13.VIN.n155 Transmission_Gate_Layout_13.VIN.n152 0.755717
R6238 Transmission_Gate_Layout_13.VIN.n181 Transmission_Gate_Layout_13.VIN.n178 0.755717
R6239 Transmission_Gate_Layout_13.VIN.n186 Transmission_Gate_Layout_13.VIN.n184 0.755717
R6240 Transmission_Gate_Layout_13.VIN.n191 Transmission_Gate_Layout_13.VIN.n190 0.755717
R6241 Transmission_Gate_Layout_13.VIN.n190 Transmission_Gate_Layout_13.VIN.n189 0.755717
R6242 Transmission_Gate_Layout_13.VIN.n102 Transmission_Gate_Layout_13.VIN.n101 0.755717
R6243 Transmission_Gate_Layout_13.VIN.n60 Transmission_Gate_Layout_13.VIN.t84 0.7285
R6244 Transmission_Gate_Layout_13.VIN.n60 Transmission_Gate_Layout_13.VIN.n59 0.7285
R6245 Transmission_Gate_Layout_13.VIN.n62 Transmission_Gate_Layout_13.VIN.t91 0.7285
R6246 Transmission_Gate_Layout_13.VIN.n62 Transmission_Gate_Layout_13.VIN.n61 0.7285
R6247 Transmission_Gate_Layout_13.VIN.n9 Transmission_Gate_Layout_13.VIN.t79 0.7285
R6248 Transmission_Gate_Layout_13.VIN.n9 Transmission_Gate_Layout_13.VIN.n8 0.7285
R6249 Transmission_Gate_Layout_13.VIN.n6 Transmission_Gate_Layout_13.VIN.t92 0.7285
R6250 Transmission_Gate_Layout_13.VIN.n6 Transmission_Gate_Layout_13.VIN.n5 0.7285
R6251 Transmission_Gate_Layout_13.VIN.n4 Transmission_Gate_Layout_13.VIN.t94 0.7285
R6252 Transmission_Gate_Layout_13.VIN.n4 Transmission_Gate_Layout_13.VIN.n3 0.7285
R6253 Transmission_Gate_Layout_13.VIN.n17 Transmission_Gate_Layout_13.VIN.t85 0.7285
R6254 Transmission_Gate_Layout_13.VIN.n17 Transmission_Gate_Layout_13.VIN.n16 0.7285
R6255 Transmission_Gate_Layout_13.VIN.n14 Transmission_Gate_Layout_13.VIN.t97 0.7285
R6256 Transmission_Gate_Layout_13.VIN.n14 Transmission_Gate_Layout_13.VIN.n13 0.7285
R6257 Transmission_Gate_Layout_13.VIN.n12 Transmission_Gate_Layout_13.VIN.t75 0.7285
R6258 Transmission_Gate_Layout_13.VIN.n12 Transmission_Gate_Layout_13.VIN.n11 0.7285
R6259 Transmission_Gate_Layout_13.VIN.n200 Transmission_Gate_Layout_13.VIN.t134 0.7285
R6260 Transmission_Gate_Layout_13.VIN.n200 Transmission_Gate_Layout_13.VIN.n199 0.7285
R6261 Transmission_Gate_Layout_13.VIN.n202 Transmission_Gate_Layout_13.VIN.t135 0.7285
R6262 Transmission_Gate_Layout_13.VIN.n202 Transmission_Gate_Layout_13.VIN.n201 0.7285
R6263 Transmission_Gate_Layout_13.VIN.n204 Transmission_Gate_Layout_13.VIN.t74 0.7285
R6264 Transmission_Gate_Layout_13.VIN.n204 Transmission_Gate_Layout_13.VIN.n203 0.7285
R6265 Transmission_Gate_Layout_13.VIN.n121 Transmission_Gate_Layout_13.VIN.t40 0.7285
R6266 Transmission_Gate_Layout_13.VIN.n121 Transmission_Gate_Layout_13.VIN.n120 0.7285
R6267 Transmission_Gate_Layout_13.VIN.n124 Transmission_Gate_Layout_13.VIN.t70 0.7285
R6268 Transmission_Gate_Layout_13.VIN.n124 Transmission_Gate_Layout_13.VIN.n123 0.7285
R6269 Transmission_Gate_Layout_13.VIN.n127 Transmission_Gate_Layout_13.VIN.t120 0.7285
R6270 Transmission_Gate_Layout_13.VIN.n127 Transmission_Gate_Layout_13.VIN.n126 0.7285
R6271 Transmission_Gate_Layout_13.VIN.n112 Transmission_Gate_Layout_13.VIN.t12 0.7285
R6272 Transmission_Gate_Layout_13.VIN.n112 Transmission_Gate_Layout_13.VIN.n111 0.7285
R6273 Transmission_Gate_Layout_13.VIN.n114 Transmission_Gate_Layout_13.VIN.t66 0.7285
R6274 Transmission_Gate_Layout_13.VIN.n114 Transmission_Gate_Layout_13.VIN.n113 0.7285
R6275 Transmission_Gate_Layout_13.VIN.n116 Transmission_Gate_Layout_13.VIN.t41 0.7285
R6276 Transmission_Gate_Layout_13.VIN.n116 Transmission_Gate_Layout_13.VIN.n115 0.7285
R6277 Transmission_Gate_Layout_13.VIN.n104 Transmission_Gate_Layout_13.VIN.t60 0.7285
R6278 Transmission_Gate_Layout_13.VIN.n104 Transmission_Gate_Layout_13.VIN.n103 0.7285
R6279 Transmission_Gate_Layout_13.VIN.n106 Transmission_Gate_Layout_13.VIN.t64 0.7285
R6280 Transmission_Gate_Layout_13.VIN.n106 Transmission_Gate_Layout_13.VIN.n105 0.7285
R6281 Transmission_Gate_Layout_13.VIN.n108 Transmission_Gate_Layout_13.VIN.t2 0.7285
R6282 Transmission_Gate_Layout_13.VIN.n108 Transmission_Gate_Layout_13.VIN.n107 0.7285
R6283 Transmission_Gate_Layout_13.VIN.n135 Transmission_Gate_Layout_13.VIN.t69 0.7285
R6284 Transmission_Gate_Layout_13.VIN.n135 Transmission_Gate_Layout_13.VIN.n134 0.7285
R6285 Transmission_Gate_Layout_13.VIN.n132 Transmission_Gate_Layout_13.VIN.t67 0.7285
R6286 Transmission_Gate_Layout_13.VIN.n132 Transmission_Gate_Layout_13.VIN.n131 0.7285
R6287 Transmission_Gate_Layout_13.VIN.n130 Transmission_Gate_Layout_13.VIN.t14 0.7285
R6288 Transmission_Gate_Layout_13.VIN.n130 Transmission_Gate_Layout_13.VIN.n129 0.7285
R6289 Transmission_Gate_Layout_13.VIN.n85 Transmission_Gate_Layout_13.VIN.t71 0.7285
R6290 Transmission_Gate_Layout_13.VIN.n85 Transmission_Gate_Layout_13.VIN.n84 0.7285
R6291 Transmission_Gate_Layout_13.VIN.n82 Transmission_Gate_Layout_13.VIN.t129 0.7285
R6292 Transmission_Gate_Layout_13.VIN.n82 Transmission_Gate_Layout_13.VIN.n81 0.7285
R6293 Transmission_Gate_Layout_13.VIN.n80 Transmission_Gate_Layout_13.VIN.t124 0.7285
R6294 Transmission_Gate_Layout_13.VIN.n80 Transmission_Gate_Layout_13.VIN.n79 0.7285
R6295 Transmission_Gate_Layout_13.VIN.n77 Transmission_Gate_Layout_13.VIN.t142 0.7285
R6296 Transmission_Gate_Layout_13.VIN.n77 Transmission_Gate_Layout_13.VIN.n76 0.7285
R6297 Transmission_Gate_Layout_13.VIN.n74 Transmission_Gate_Layout_13.VIN.t126 0.7285
R6298 Transmission_Gate_Layout_13.VIN.n74 Transmission_Gate_Layout_13.VIN.n73 0.7285
R6299 Transmission_Gate_Layout_13.VIN.n72 Transmission_Gate_Layout_13.VIN.t39 0.7285
R6300 Transmission_Gate_Layout_13.VIN.n72 Transmission_Gate_Layout_13.VIN.n71 0.7285
R6301 Transmission_Gate_Layout_13.VIN.n64 Transmission_Gate_Layout_13.VIN.t82 0.7285
R6302 Transmission_Gate_Layout_13.VIN.n64 Transmission_Gate_Layout_13.VIN.n63 0.7285
R6303 Transmission_Gate_Layout_13.VIN.n53 Transmission_Gate_Layout_13.VIN.n52 0.626587
R6304 Transmission_Gate_Layout_13.VIN.n55 Transmission_Gate_Layout_13.VIN.n54 0.626587
R6305 Transmission_Gate_Layout_13.VIN.n146 Transmission_Gate_Layout_13.VIN.n145 0.626587
R6306 Transmission_Gate_Layout_13.VIN.n193 Transmission_Gate_Layout_13.VIN.n192 0.626587
R6307 Transmission_Gate_Layout_13.VIN.n195 Transmission_Gate_Layout_13.VIN.n194 0.626587
R6308 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.VIN.n213 0.607022
R6309 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_13.VIN.n70 0.607022
R6310 Transmission_Gate_Layout_13.VIN.n55 Transmission_Gate_Layout_13.VIN.n10 0.575717
R6311 Transmission_Gate_Layout_13.VIN.n54 Transmission_Gate_Layout_13.VIN.n18 0.575717
R6312 Transmission_Gate_Layout_13.VIN.n119 Transmission_Gate_Layout_13.VIN.n110 0.575717
R6313 Transmission_Gate_Layout_13.VIN.n194 Transmission_Gate_Layout_13.VIN.n86 0.575717
R6314 Transmission_Gate_Layout_13.VIN.n195 Transmission_Gate_Layout_13.VIN.n78 0.575717
R6315 Transmission_Gate_Layout_13.VIN.n207 Transmission_Gate_Layout_13.VIN.n206 0.575717
R6316 Transmission_Gate_Layout_13.VIN.n67 Transmission_Gate_Layout_13.VIN.n66 0.575717
R6317 Transmission_Gate_Layout_13.VIN.n173 Transmission_Gate_Layout_13.VIN.n172 0.570002
R6318 Transmission_Gate_Layout_13.VIN.n145 Transmission_Gate_Layout_13.VIN.n144 0.428978
R6319 Transmission_Gate_Layout_13.VIN.n149 Transmission_Gate_Layout_13.VIN.n146 0.428978
R6320 Transmission_Gate_Layout_13.VIN.n53 Transmission_Gate_Layout_13.VIN.n26 0.331152
R6321 Transmission_Gate_Layout_13.VIN.n52 Transmission_Gate_Layout_13.VIN.n34 0.331152
R6322 Transmission_Gate_Layout_13.VIN.n48 Transmission_Gate_Layout_13.VIN.n45 0.331152
R6323 Transmission_Gate_Layout_13.VIN.n193 Transmission_Gate_Layout_13.VIN.n94 0.331152
R6324 Transmission_Gate_Layout_13.VIN.n172 Transmission_Gate_Layout_13.VIN.n163 0.331152
R6325 Transmission_Gate_Layout_13.VIN.n187 Transmission_Gate_Layout_13.VIN.n181 0.331152
R6326 Transmission_Gate_Layout_13.VIN.n192 Transmission_Gate_Layout_13.VIN.n102 0.331152
R6327 Transmission_Gate_Layout_13.VIN.n173 Transmission_Gate_Layout_13.VIN.n155 0.317457
R6328 Transmission_Gate_Layout_13.VIN.n189 Transmission_Gate_Layout_13.VIN.n188 0.317457
R6329 Transmission_Gate_Layout_13.VIN.n54 Transmission_Gate_Layout_13.VIN.n53 0.239196
R6330 Transmission_Gate_Layout_13.VIN.n194 Transmission_Gate_Layout_13.VIN.n193 0.239196
R6331 Transmission_Gate_Layout_13.VIN.n145 Transmission_Gate_Layout_13.VIN 0.192239
R6332 Transmission_Gate_Layout_13.CLK.t4 Transmission_Gate_Layout_13.CLK.t34 82.9076
R6333 Transmission_Gate_Layout_13.CLK.t23 Transmission_Gate_Layout_13.CLK.t4 82.9076
R6334 Transmission_Gate_Layout_13.CLK.n25 Transmission_Gate_Layout_13.CLK.t23 49.7969
R6335 Transmission_Gate_Layout_13.CLK.n24 Transmission_Gate_Layout_13.CLK.n23 35.0405
R6336 Transmission_Gate_Layout_13.CLK.n25 Transmission_Gate_Layout_13.CLK.t2 31.1559
R6337 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_13.CLK.n27 24.3453
R6338 Transmission_Gate_Layout_13.CLK.n26 Transmission_Gate_Layout_13.CLK.t11 22.0309
R6339 Transmission_Gate_Layout_13.CLK.t25 Transmission_Gate_Layout_13.CLK.n0 21.9005
R6340 Transmission_Gate_Layout_13.CLK.t12 Transmission_Gate_Layout_13.CLK.n15 21.9005
R6341 Transmission_Gate_Layout_13.CLK.n16 Transmission_Gate_Layout_13.CLK.t20 21.5094
R6342 Transmission_Gate_Layout_13.CLK.n17 Transmission_Gate_Layout_13.CLK.t13 21.5094
R6343 Transmission_Gate_Layout_13.CLK.n18 Transmission_Gate_Layout_13.CLK.t6 21.5094
R6344 Transmission_Gate_Layout_13.CLK.n19 Transmission_Gate_Layout_13.CLK.t17 21.5094
R6345 Transmission_Gate_Layout_13.CLK.n20 Transmission_Gate_Layout_13.CLK.t10 21.5094
R6346 Transmission_Gate_Layout_13.CLK.n21 Transmission_Gate_Layout_13.CLK.t24 21.5094
R6347 Transmission_Gate_Layout_13.CLK.n22 Transmission_Gate_Layout_13.CLK.t18 21.5094
R6348 Transmission_Gate_Layout_13.CLK.n24 Transmission_Gate_Layout_13.CLK.t25 21.5094
R6349 Transmission_Gate_Layout_13.CLK.n23 Transmission_Gate_Layout_13.CLK.t12 21.5094
R6350 Transmission_Gate_Layout_13.CLK.n27 Transmission_Gate_Layout_13.CLK.t3 21.3791
R6351 Transmission_Gate_Layout_13.CLK.n26 Transmission_Gate_Layout_13.CLK.t8 21.3791
R6352 Transmission_Gate_Layout_13.CLK.n16 Transmission_Gate_Layout_13.CLK.t29 20.988
R6353 Transmission_Gate_Layout_13.CLK.n17 Transmission_Gate_Layout_13.CLK.t22 20.988
R6354 Transmission_Gate_Layout_13.CLK.n18 Transmission_Gate_Layout_13.CLK.t16 20.988
R6355 Transmission_Gate_Layout_13.CLK.n19 Transmission_Gate_Layout_13.CLK.t26 20.988
R6356 Transmission_Gate_Layout_13.CLK.n20 Transmission_Gate_Layout_13.CLK.t19 20.988
R6357 Transmission_Gate_Layout_13.CLK.n21 Transmission_Gate_Layout_13.CLK.t32 20.988
R6358 Transmission_Gate_Layout_13.CLK.n22 Transmission_Gate_Layout_13.CLK.t27 20.988
R6359 Transmission_Gate_Layout_13.CLK.n23 Transmission_Gate_Layout_13.CLK.t21 20.988
R6360 Transmission_Gate_Layout_13.CLK.t2 Transmission_Gate_Layout_13.CLK.n24 20.988
R6361 Transmission_Gate_Layout_13.CLK.n27 Transmission_Gate_Layout_13.CLK.n26 20.8576
R6362 Transmission_Gate_Layout_13.CLK.n8 Transmission_Gate_Layout_13.CLK.t9 20.5969
R6363 Transmission_Gate_Layout_13.CLK.n9 Transmission_Gate_Layout_13.CLK.t33 20.5969
R6364 Transmission_Gate_Layout_13.CLK.n10 Transmission_Gate_Layout_13.CLK.t28 20.5969
R6365 Transmission_Gate_Layout_13.CLK.n11 Transmission_Gate_Layout_13.CLK.t5 20.5969
R6366 Transmission_Gate_Layout_13.CLK.n12 Transmission_Gate_Layout_13.CLK.t30 20.5969
R6367 Transmission_Gate_Layout_13.CLK.n13 Transmission_Gate_Layout_13.CLK.t14 20.5969
R6368 Transmission_Gate_Layout_13.CLK.n14 Transmission_Gate_Layout_13.CLK.t7 20.5969
R6369 Transmission_Gate_Layout_13.CLK.n15 Transmission_Gate_Layout_13.CLK.t31 20.5969
R6370 Transmission_Gate_Layout_13.CLK.n0 Transmission_Gate_Layout_13.CLK.t15 20.5969
R6371 Transmission_Gate_Layout_13.CLK.n9 Transmission_Gate_Layout_13.CLK.n8 19.4672
R6372 Transmission_Gate_Layout_13.CLK.n10 Transmission_Gate_Layout_13.CLK.n9 19.4672
R6373 Transmission_Gate_Layout_13.CLK.n11 Transmission_Gate_Layout_13.CLK.n10 19.4672
R6374 Transmission_Gate_Layout_13.CLK.n12 Transmission_Gate_Layout_13.CLK.n11 19.4672
R6375 Transmission_Gate_Layout_13.CLK.n13 Transmission_Gate_Layout_13.CLK.n12 19.4672
R6376 Transmission_Gate_Layout_13.CLK.n14 Transmission_Gate_Layout_13.CLK.n13 19.4672
R6377 Transmission_Gate_Layout_13.CLK.n15 Transmission_Gate_Layout_13.CLK.n14 19.4672
R6378 Transmission_Gate_Layout_13.CLK.n17 Transmission_Gate_Layout_13.CLK.n16 19.4672
R6379 Transmission_Gate_Layout_13.CLK.n18 Transmission_Gate_Layout_13.CLK.n17 19.4672
R6380 Transmission_Gate_Layout_13.CLK.n19 Transmission_Gate_Layout_13.CLK.n18 19.4672
R6381 Transmission_Gate_Layout_13.CLK.n20 Transmission_Gate_Layout_13.CLK.n19 19.4672
R6382 Transmission_Gate_Layout_13.CLK.n21 Transmission_Gate_Layout_13.CLK.n20 19.4672
R6383 Transmission_Gate_Layout_13.CLK.n22 Transmission_Gate_Layout_13.CLK.n21 19.4672
R6384 Transmission_Gate_Layout_13.CLK.n23 Transmission_Gate_Layout_13.CLK.n22 19.4672
R6385 Transmission_Gate_Layout_13.CLK.t33 Transmission_Gate_Layout_13.CLK.n7 18.9023
R6386 Transmission_Gate_Layout_13.CLK.t28 Transmission_Gate_Layout_13.CLK.n6 18.9023
R6387 Transmission_Gate_Layout_13.CLK.t5 Transmission_Gate_Layout_13.CLK.n5 18.9023
R6388 Transmission_Gate_Layout_13.CLK.t30 Transmission_Gate_Layout_13.CLK.n4 18.9023
R6389 Transmission_Gate_Layout_13.CLK.t14 Transmission_Gate_Layout_13.CLK.n3 18.9023
R6390 Transmission_Gate_Layout_13.CLK.t7 Transmission_Gate_Layout_13.CLK.n2 18.9023
R6391 Transmission_Gate_Layout_13.CLK.t31 Transmission_Gate_Layout_13.CLK.n1 18.9023
R6392 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_13.CLK.n25 16.4436
R6393 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_13.CLK.n28 7.70137
R6394 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_13.CLK.n29 4.70224
R6395 Transmission_Gate_Layout_13.CLKB.n27 Transmission_Gate_Layout_13.CLKB.t10 54.5477
R6396 Transmission_Gate_Layout_13.CLKB.n27 Transmission_Gate_Layout_13.CLKB.t6 38.3255
R6397 Transmission_Gate_Layout_13.CLKB.n28 Transmission_Gate_Layout_13.CLKB.t11 38.3255
R6398 Transmission_Gate_Layout_13.CLKB.n29 Transmission_Gate_Layout_13.CLKB.t8 38.3255
R6399 Transmission_Gate_Layout_13.CLKB.n30 Transmission_Gate_Layout_13.CLKB.t20 38.3255
R6400 Transmission_Gate_Layout_13.CLKB.n32 Transmission_Gate_Layout_13.CLKB.t9 38.3255
R6401 Transmission_Gate_Layout_13.CLKB.n31 Transmission_Gate_Layout_13.CLKB.t13 38.3255
R6402 Transmission_Gate_Layout_13.CLKB.t28 Transmission_Gate_Layout_13.CLKB.n24 37.9344
R6403 Transmission_Gate_Layout_13.CLKB.t22 Transmission_Gate_Layout_13.CLKB.n23 37.9344
R6404 Transmission_Gate_Layout_13.CLKB.t15 Transmission_Gate_Layout_13.CLKB.n20 37.9344
R6405 Transmission_Gate_Layout_13.CLKB.t25 Transmission_Gate_Layout_13.CLKB.n17 37.9344
R6406 Transmission_Gate_Layout_13.CLKB.t18 Transmission_Gate_Layout_13.CLKB.n14 37.9344
R6407 Transmission_Gate_Layout_13.CLKB.t7 Transmission_Gate_Layout_13.CLKB.n11 37.9344
R6408 Transmission_Gate_Layout_13.CLKB.t27 Transmission_Gate_Layout_13.CLKB.n8 37.9344
R6409 Transmission_Gate_Layout_13.CLKB.t21 Transmission_Gate_Layout_13.CLKB.n5 37.9344
R6410 Transmission_Gate_Layout_13.CLKB.n25 Transmission_Gate_Layout_13.CLKB.t28 37.5434
R6411 Transmission_Gate_Layout_13.CLKB.n26 Transmission_Gate_Layout_13.CLKB.t22 37.5434
R6412 Transmission_Gate_Layout_13.CLKB.n21 Transmission_Gate_Layout_13.CLKB.t15 37.5434
R6413 Transmission_Gate_Layout_13.CLKB.n18 Transmission_Gate_Layout_13.CLKB.t25 37.5434
R6414 Transmission_Gate_Layout_13.CLKB.n15 Transmission_Gate_Layout_13.CLKB.t18 37.5434
R6415 Transmission_Gate_Layout_13.CLKB.n12 Transmission_Gate_Layout_13.CLKB.t7 37.5434
R6416 Transmission_Gate_Layout_13.CLKB.n9 Transmission_Gate_Layout_13.CLKB.t27 37.5434
R6417 Transmission_Gate_Layout_13.CLKB.n6 Transmission_Gate_Layout_13.CLKB.t21 37.5434
R6418 Transmission_Gate_Layout_13.CLKB.n25 Transmission_Gate_Layout_13.CLKB.t14 37.413
R6419 Transmission_Gate_Layout_13.CLKB.t10 Transmission_Gate_Layout_13.CLKB.n26 37.413
R6420 Transmission_Gate_Layout_13.CLKB.t6 Transmission_Gate_Layout_13.CLKB.n21 37.413
R6421 Transmission_Gate_Layout_13.CLKB.t11 Transmission_Gate_Layout_13.CLKB.n18 37.413
R6422 Transmission_Gate_Layout_13.CLKB.t8 Transmission_Gate_Layout_13.CLKB.n15 37.413
R6423 Transmission_Gate_Layout_13.CLKB.t20 Transmission_Gate_Layout_13.CLKB.n12 37.413
R6424 Transmission_Gate_Layout_13.CLKB.t9 Transmission_Gate_Layout_13.CLKB.n6 37.413
R6425 Transmission_Gate_Layout_13.CLKB.t13 Transmission_Gate_Layout_13.CLKB.n9 37.413
R6426 Transmission_Gate_Layout_13.CLKB.n5 Transmission_Gate_Layout_13.CLKB.t17 37.0219
R6427 Transmission_Gate_Layout_13.CLKB.n11 Transmission_Gate_Layout_13.CLKB.t29 37.0219
R6428 Transmission_Gate_Layout_13.CLKB.n14 Transmission_Gate_Layout_13.CLKB.t16 37.0219
R6429 Transmission_Gate_Layout_13.CLKB.n17 Transmission_Gate_Layout_13.CLKB.t23 37.0219
R6430 Transmission_Gate_Layout_13.CLKB.n20 Transmission_Gate_Layout_13.CLKB.t12 37.0219
R6431 Transmission_Gate_Layout_13.CLKB.n23 Transmission_Gate_Layout_13.CLKB.t19 37.0219
R6432 Transmission_Gate_Layout_13.CLKB.n24 Transmission_Gate_Layout_13.CLKB.t26 37.0219
R6433 Transmission_Gate_Layout_13.CLKB.n8 Transmission_Gate_Layout_13.CLKB.t24 37.0219
R6434 Transmission_Gate_Layout_13.CLKB.t29 Transmission_Gate_Layout_13.CLKB.n10 35.1969
R6435 Transmission_Gate_Layout_13.CLKB.t16 Transmission_Gate_Layout_13.CLKB.n13 35.1969
R6436 Transmission_Gate_Layout_13.CLKB.t23 Transmission_Gate_Layout_13.CLKB.n16 35.1969
R6437 Transmission_Gate_Layout_13.CLKB.t12 Transmission_Gate_Layout_13.CLKB.n19 35.1969
R6438 Transmission_Gate_Layout_13.CLKB.t19 Transmission_Gate_Layout_13.CLKB.n22 35.1969
R6439 Transmission_Gate_Layout_13.CLKB.t24 Transmission_Gate_Layout_13.CLKB.n7 35.1969
R6440 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLKB.n32 26.6826
R6441 Transmission_Gate_Layout_13.CLKB.n26 Transmission_Gate_Layout_13.CLKB.n25 19.148
R6442 Transmission_Gate_Layout_13.CLKB.n28 Transmission_Gate_Layout_13.CLKB.n27 16.2227
R6443 Transmission_Gate_Layout_13.CLKB.n29 Transmission_Gate_Layout_13.CLKB.n28 16.2227
R6444 Transmission_Gate_Layout_13.CLKB.n30 Transmission_Gate_Layout_13.CLKB.n29 16.2227
R6445 Transmission_Gate_Layout_13.CLKB.n31 Transmission_Gate_Layout_13.CLKB.n30 16.2227
R6446 Transmission_Gate_Layout_13.CLKB.n32 Transmission_Gate_Layout_13.CLKB.n31 16.2227
R6447 Transmission_Gate_Layout_13.CLKB.n36 Transmission_Gate_Layout_13.CLKB.n35 5.21612
R6448 Transmission_Gate_Layout_13.CLKB.n2 Transmission_Gate_Layout_13.CLKB.n0 4.57285
R6449 Transmission_Gate_Layout_13.CLKB.n37 Transmission_Gate_Layout_13.CLKB.n33 4.4609
R6450 Transmission_Gate_Layout_13.CLKB.n36 Transmission_Gate_Layout_13.CLKB.n34 4.4609
R6451 Transmission_Gate_Layout_13.CLKB.n4 Transmission_Gate_Layout_13.CLKB.n3 3.3285
R6452 Transmission_Gate_Layout_13.CLKB.n2 Transmission_Gate_Layout_13.CLKB.n1 3.3285
R6453 Transmission_Gate_Layout_13.CLKB.n4 Transmission_Gate_Layout_13.CLKB.n2 1.24485
R6454 Transmission_Gate_Layout_13.CLKB.n37 Transmission_Gate_Layout_13.CLKB.n36 0.755717
R6455 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLKB.n4 0.750969
R6456 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.CLKB.n37 0.510317
R6457 OUT.n136 OUT 8.9529
R6458 OUT.n46 OUT.t86 5.21612
R6459 OUT.n113 OUT.n111 5.21612
R6460 OUT.n51 OUT.n35 4.4609
R6461 OUT.n50 OUT.n36 4.4609
R6462 OUT.n49 OUT.n37 4.4609
R6463 OUT.n47 OUT.t95 4.4609
R6464 OUT.n46 OUT.t79 4.4609
R6465 OUT.n119 OUT.t58 4.4609
R6466 OUT.n118 OUT.t66 4.4609
R6467 OUT.n117 OUT.t50 4.4609
R6468 OUT.n115 OUT.n114 4.4609
R6469 OUT.n113 OUT.n112 4.4609
R6470 OUT.n25 OUT.n24 3.90572
R6471 OUT.n33 OUT.n32 3.90572
R6472 OUT.n42 OUT.n39 3.90572
R6473 OUT.n93 OUT.n92 3.90572
R6474 OUT.n107 OUT.n104 3.90572
R6475 OUT.n101 OUT.n100 3.90572
R6476 OUT.n7 OUT.n4 3.84485
R6477 OUT.n15 OUT.n12 3.84485
R6478 OUT.n65 OUT.n64 3.84485
R6479 OUT.n83 OUT.n80 3.84485
R6480 OUT.n75 OUT.n72 3.84485
R6481 OUT.n133 OUT.n132 3.84485
R6482 OUT.n138 OUT.n137 3.3285
R6483 OUT.n140 OUT.n139 3.3285
R6484 OUT.n142 OUT.n141 3.3285
R6485 OUT.n70 OUT.t39 3.3285
R6486 OUT.n69 OUT.t26 3.3285
R6487 OUT.n68 OUT.t46 3.3285
R6488 OUT.n58 OUT.n0 3.3285
R6489 OUT.n57 OUT.n1 3.3285
R6490 OUT.n56 OUT.n2 3.3285
R6491 OUT.n126 OUT.t12 3.3285
R6492 OUT.n125 OUT.t8 3.3285
R6493 OUT.n124 OUT.t20 3.3285
R6494 OUT.n25 OUT.n22 3.1505
R6495 OUT.n26 OUT.n20 3.1505
R6496 OUT.n33 OUT.n30 3.1505
R6497 OUT.n34 OUT.n28 3.1505
R6498 OUT.n42 OUT.n41 3.1505
R6499 OUT.n45 OUT.n44 3.1505
R6500 OUT.n93 OUT.n90 3.1505
R6501 OUT.n94 OUT.n88 3.1505
R6502 OUT.n107 OUT.n106 3.1505
R6503 OUT.n110 OUT.n109 3.1505
R6504 OUT.n101 OUT.n98 3.1505
R6505 OUT.n102 OUT.n96 3.1505
R6506 OUT.n67 OUT.n58 2.72398
R6507 OUT.n135 OUT.n126 2.72398
R6508 OUT.n7 OUT.n6 2.6005
R6509 OUT.n10 OUT.n9 2.6005
R6510 OUT.n15 OUT.n14 2.6005
R6511 OUT.n18 OUT.n17 2.6005
R6512 OUT.n65 OUT.n62 2.6005
R6513 OUT.n66 OUT.n60 2.6005
R6514 OUT.n83 OUT.n82 2.6005
R6515 OUT.n86 OUT.n85 2.6005
R6516 OUT.n75 OUT.n74 2.6005
R6517 OUT.n78 OUT.n77 2.6005
R6518 OUT.n133 OUT.n130 2.6005
R6519 OUT.n134 OUT.n128 2.6005
R6520 OUT.n49 OUT.n48 2.47941
R6521 OUT.n117 OUT.n116 2.47941
R6522 OUT.n20 OUT.t78 1.3109
R6523 OUT.n20 OUT.n19 1.3109
R6524 OUT.n22 OUT.t94 1.3109
R6525 OUT.n22 OUT.n21 1.3109
R6526 OUT.n24 OUT.t87 1.3109
R6527 OUT.n24 OUT.n23 1.3109
R6528 OUT.n28 OUT.t72 1.3109
R6529 OUT.n28 OUT.n27 1.3109
R6530 OUT.n30 OUT.t88 1.3109
R6531 OUT.n30 OUT.n29 1.3109
R6532 OUT.n32 OUT.t80 1.3109
R6533 OUT.n32 OUT.n31 1.3109
R6534 OUT.n44 OUT.t91 1.3109
R6535 OUT.n44 OUT.n43 1.3109
R6536 OUT.n41 OUT.t76 1.3109
R6537 OUT.n41 OUT.n40 1.3109
R6538 OUT.n39 OUT.t83 1.3109
R6539 OUT.n39 OUT.n38 1.3109
R6540 OUT.n88 OUT.t55 1.3109
R6541 OUT.n88 OUT.n87 1.3109
R6542 OUT.n90 OUT.t62 1.3109
R6543 OUT.n90 OUT.n89 1.3109
R6544 OUT.n92 OUT.t71 1.3109
R6545 OUT.n92 OUT.n91 1.3109
R6546 OUT.n109 OUT.t48 1.3109
R6547 OUT.n109 OUT.n108 1.3109
R6548 OUT.n106 OUT.t65 1.3109
R6549 OUT.n106 OUT.n105 1.3109
R6550 OUT.n104 OUT.t57 1.3109
R6551 OUT.n104 OUT.n103 1.3109
R6552 OUT.n96 OUT.t49 1.3109
R6553 OUT.n96 OUT.n95 1.3109
R6554 OUT.n98 OUT.t56 1.3109
R6555 OUT.n98 OUT.n97 1.3109
R6556 OUT.n100 OUT.t64 1.3109
R6557 OUT.n100 OUT.n99 1.3109
R6558 OUT.n10 OUT.n7 1.24485
R6559 OUT.n18 OUT.n15 1.24485
R6560 OUT.n58 OUT.n57 1.24485
R6561 OUT.n57 OUT.n56 1.24485
R6562 OUT.n66 OUT.n65 1.24485
R6563 OUT.n69 OUT.n68 1.24485
R6564 OUT.n70 OUT.n69 1.24485
R6565 OUT.n140 OUT.n138 1.24485
R6566 OUT.n142 OUT.n140 1.24485
R6567 OUT.n86 OUT.n83 1.24485
R6568 OUT.n78 OUT.n75 1.24485
R6569 OUT.n126 OUT.n125 1.24485
R6570 OUT.n125 OUT.n124 1.24485
R6571 OUT.n134 OUT.n133 1.24485
R6572 OUT.n56 OUT.n55 1.2018
R6573 OUT.n68 OUT.n67 1.2018
R6574 OUT.n124 OUT.n123 1.2018
R6575 OUT.n48 OUT.n47 0.957239
R6576 OUT.n52 OUT.n51 0.957239
R6577 OUT.n116 OUT.n115 0.957239
R6578 OUT.n120 OUT.n119 0.957239
R6579 OUT.n26 OUT.n25 0.755717
R6580 OUT.n34 OUT.n33 0.755717
R6581 OUT.n45 OUT.n42 0.755717
R6582 OUT.n47 OUT.n46 0.755717
R6583 OUT.n51 OUT.n50 0.755717
R6584 OUT.n50 OUT.n49 0.755717
R6585 OUT.n94 OUT.n93 0.755717
R6586 OUT.n110 OUT.n107 0.755717
R6587 OUT.n115 OUT.n113 0.755717
R6588 OUT.n119 OUT.n118 0.755717
R6589 OUT.n118 OUT.n117 0.755717
R6590 OUT.n102 OUT.n101 0.755717
R6591 OUT.n60 OUT.t43 0.7285
R6592 OUT.n60 OUT.n59 0.7285
R6593 OUT.n62 OUT.t45 0.7285
R6594 OUT.n62 OUT.n61 0.7285
R6595 OUT.n64 OUT.t34 0.7285
R6596 OUT.n64 OUT.n63 0.7285
R6597 OUT.n9 OUT.t24 0.7285
R6598 OUT.n9 OUT.n8 0.7285
R6599 OUT.n6 OUT.t31 0.7285
R6600 OUT.n6 OUT.n5 0.7285
R6601 OUT.n4 OUT.t30 0.7285
R6602 OUT.n4 OUT.n3 0.7285
R6603 OUT.n17 OUT.t29 0.7285
R6604 OUT.n17 OUT.n16 0.7285
R6605 OUT.n14 OUT.t41 0.7285
R6606 OUT.n14 OUT.n13 0.7285
R6607 OUT.n12 OUT.t38 0.7285
R6608 OUT.n12 OUT.n11 0.7285
R6609 OUT.n128 OUT.t10 0.7285
R6610 OUT.n128 OUT.n127 0.7285
R6611 OUT.n130 OUT.t7 0.7285
R6612 OUT.n130 OUT.n129 0.7285
R6613 OUT.n132 OUT.t19 0.7285
R6614 OUT.n132 OUT.n131 0.7285
R6615 OUT.n85 OUT.t18 0.7285
R6616 OUT.n85 OUT.n84 0.7285
R6617 OUT.n82 OUT.t4 0.7285
R6618 OUT.n82 OUT.n81 0.7285
R6619 OUT.n80 OUT.t6 0.7285
R6620 OUT.n80 OUT.n79 0.7285
R6621 OUT.n77 OUT.t9 0.7285
R6622 OUT.n77 OUT.n76 0.7285
R6623 OUT.n74 OUT.t22 0.7285
R6624 OUT.n74 OUT.n73 0.7285
R6625 OUT.n72 OUT.t0 0.7285
R6626 OUT.n72 OUT.n71 0.7285
R6627 OUT.n53 OUT.n52 0.626587
R6628 OUT.n55 OUT.n54 0.626587
R6629 OUT.n121 OUT.n120 0.626587
R6630 OUT.n123 OUT.n122 0.626587
R6631 OUT OUT.n70 0.607022
R6632 OUT OUT.n142 0.607022
R6633 OUT.n136 OUT.n135 0.597239
R6634 OUT.n55 OUT.n10 0.575717
R6635 OUT.n54 OUT.n18 0.575717
R6636 OUT.n67 OUT.n66 0.575717
R6637 OUT.n122 OUT.n86 0.575717
R6638 OUT.n123 OUT.n78 0.575717
R6639 OUT.n135 OUT.n134 0.575717
R6640 OUT.n138 OUT.n136 0.54637
R6641 OUT.n53 OUT.n26 0.331152
R6642 OUT.n52 OUT.n34 0.331152
R6643 OUT.n48 OUT.n45 0.331152
R6644 OUT.n121 OUT.n94 0.331152
R6645 OUT.n116 OUT.n110 0.331152
R6646 OUT.n120 OUT.n102 0.331152
R6647 OUT.n54 OUT.n53 0.239196
R6648 OUT.n122 OUT.n121 0.239196
R6649 Transmission_Gate_Layout_0.CLKB.n24 Transmission_Gate_Layout_0.CLKB.t7 54.5477
R6650 Transmission_Gate_Layout_0.CLKB.n29 Transmission_Gate_Layout_0.CLKB.t29 38.3255
R6651 Transmission_Gate_Layout_0.CLKB.n28 Transmission_Gate_Layout_0.CLKB.t11 38.3255
R6652 Transmission_Gate_Layout_0.CLKB.n27 Transmission_Gate_Layout_0.CLKB.t23 38.3255
R6653 Transmission_Gate_Layout_0.CLKB.n26 Transmission_Gate_Layout_0.CLKB.t28 38.3255
R6654 Transmission_Gate_Layout_0.CLKB.n25 Transmission_Gate_Layout_0.CLKB.t19 38.3255
R6655 Transmission_Gate_Layout_0.CLKB.n24 Transmission_Gate_Layout_0.CLKB.t24 38.3255
R6656 Transmission_Gate_Layout_0.CLKB.t17 Transmission_Gate_Layout_0.CLKB.n2 37.9344
R6657 Transmission_Gate_Layout_0.CLKB.t22 Transmission_Gate_Layout_0.CLKB.n5 37.9344
R6658 Transmission_Gate_Layout_0.CLKB.t9 Transmission_Gate_Layout_0.CLKB.n8 37.9344
R6659 Transmission_Gate_Layout_0.CLKB.t15 Transmission_Gate_Layout_0.CLKB.n11 37.9344
R6660 Transmission_Gate_Layout_0.CLKB.t26 Transmission_Gate_Layout_0.CLKB.n14 37.9344
R6661 Transmission_Gate_Layout_0.CLKB.t12 Transmission_Gate_Layout_0.CLKB.n17 37.9344
R6662 Transmission_Gate_Layout_0.CLKB.t18 Transmission_Gate_Layout_0.CLKB.n20 37.9344
R6663 Transmission_Gate_Layout_0.CLKB.t6 Transmission_Gate_Layout_0.CLKB.n21 37.9344
R6664 Transmission_Gate_Layout_0.CLKB.n3 Transmission_Gate_Layout_0.CLKB.t17 37.5434
R6665 Transmission_Gate_Layout_0.CLKB.n6 Transmission_Gate_Layout_0.CLKB.t22 37.5434
R6666 Transmission_Gate_Layout_0.CLKB.n9 Transmission_Gate_Layout_0.CLKB.t9 37.5434
R6667 Transmission_Gate_Layout_0.CLKB.n12 Transmission_Gate_Layout_0.CLKB.t15 37.5434
R6668 Transmission_Gate_Layout_0.CLKB.n15 Transmission_Gate_Layout_0.CLKB.t26 37.5434
R6669 Transmission_Gate_Layout_0.CLKB.n18 Transmission_Gate_Layout_0.CLKB.t12 37.5434
R6670 Transmission_Gate_Layout_0.CLKB.n23 Transmission_Gate_Layout_0.CLKB.t18 37.5434
R6671 Transmission_Gate_Layout_0.CLKB.n22 Transmission_Gate_Layout_0.CLKB.t6 37.5434
R6672 Transmission_Gate_Layout_0.CLKB.t29 Transmission_Gate_Layout_0.CLKB.n3 37.413
R6673 Transmission_Gate_Layout_0.CLKB.t11 Transmission_Gate_Layout_0.CLKB.n6 37.413
R6674 Transmission_Gate_Layout_0.CLKB.t23 Transmission_Gate_Layout_0.CLKB.n9 37.413
R6675 Transmission_Gate_Layout_0.CLKB.t28 Transmission_Gate_Layout_0.CLKB.n12 37.413
R6676 Transmission_Gate_Layout_0.CLKB.t19 Transmission_Gate_Layout_0.CLKB.n15 37.413
R6677 Transmission_Gate_Layout_0.CLKB.t24 Transmission_Gate_Layout_0.CLKB.n18 37.413
R6678 Transmission_Gate_Layout_0.CLKB.n22 Transmission_Gate_Layout_0.CLKB.t21 37.413
R6679 Transmission_Gate_Layout_0.CLKB.t7 Transmission_Gate_Layout_0.CLKB.n23 37.413
R6680 Transmission_Gate_Layout_0.CLKB.n21 Transmission_Gate_Layout_0.CLKB.t27 37.0219
R6681 Transmission_Gate_Layout_0.CLKB.n17 Transmission_Gate_Layout_0.CLKB.t10 37.0219
R6682 Transmission_Gate_Layout_0.CLKB.n14 Transmission_Gate_Layout_0.CLKB.t25 37.0219
R6683 Transmission_Gate_Layout_0.CLKB.n11 Transmission_Gate_Layout_0.CLKB.t13 37.0219
R6684 Transmission_Gate_Layout_0.CLKB.n8 Transmission_Gate_Layout_0.CLKB.t8 37.0219
R6685 Transmission_Gate_Layout_0.CLKB.n5 Transmission_Gate_Layout_0.CLKB.t20 37.0219
R6686 Transmission_Gate_Layout_0.CLKB.n2 Transmission_Gate_Layout_0.CLKB.t14 37.0219
R6687 Transmission_Gate_Layout_0.CLKB.n20 Transmission_Gate_Layout_0.CLKB.t16 37.0219
R6688 Transmission_Gate_Layout_0.CLKB.t10 Transmission_Gate_Layout_0.CLKB.n16 35.1969
R6689 Transmission_Gate_Layout_0.CLKB.t25 Transmission_Gate_Layout_0.CLKB.n13 35.1969
R6690 Transmission_Gate_Layout_0.CLKB.t13 Transmission_Gate_Layout_0.CLKB.n10 35.1969
R6691 Transmission_Gate_Layout_0.CLKB.t8 Transmission_Gate_Layout_0.CLKB.n7 35.1969
R6692 Transmission_Gate_Layout_0.CLKB.t20 Transmission_Gate_Layout_0.CLKB.n4 35.1969
R6693 Transmission_Gate_Layout_0.CLKB.t16 Transmission_Gate_Layout_0.CLKB.n19 35.1969
R6694 Transmission_Gate_Layout_0.CLKB Transmission_Gate_Layout_0.CLKB.n29 26.6826
R6695 Transmission_Gate_Layout_0.CLKB.n23 Transmission_Gate_Layout_0.CLKB.n22 19.148
R6696 Transmission_Gate_Layout_0.CLKB.n29 Transmission_Gate_Layout_0.CLKB.n28 16.2227
R6697 Transmission_Gate_Layout_0.CLKB.n28 Transmission_Gate_Layout_0.CLKB.n27 16.2227
R6698 Transmission_Gate_Layout_0.CLKB.n27 Transmission_Gate_Layout_0.CLKB.n26 16.2227
R6699 Transmission_Gate_Layout_0.CLKB.n26 Transmission_Gate_Layout_0.CLKB.n25 16.2227
R6700 Transmission_Gate_Layout_0.CLKB.n25 Transmission_Gate_Layout_0.CLKB.n24 16.2227
R6701 Transmission_Gate_Layout_0.CLKB.n30 Transmission_Gate_Layout_0.CLKB.t4 5.21612
R6702 Transmission_Gate_Layout_0.CLKB.n0 Transmission_Gate_Layout_0.CLKB.t2 4.57285
R6703 Transmission_Gate_Layout_0.CLKB.n31 Transmission_Gate_Layout_0.CLKB.t3 4.4609
R6704 Transmission_Gate_Layout_0.CLKB.n30 Transmission_Gate_Layout_0.CLKB.t1 4.4609
R6705 Transmission_Gate_Layout_0.CLKB.n0 Transmission_Gate_Layout_0.CLKB.t5 3.3285
R6706 Transmission_Gate_Layout_0.CLKB.n1 Transmission_Gate_Layout_0.CLKB.t0 3.3285
R6707 Transmission_Gate_Layout_0.CLKB.n1 Transmission_Gate_Layout_0.CLKB.n0 1.24485
R6708 Transmission_Gate_Layout_0.CLKB.n31 Transmission_Gate_Layout_0.CLKB.n30 0.755717
R6709 Transmission_Gate_Layout_0.CLKB Transmission_Gate_Layout_0.CLKB.n1 0.750969
R6710 Transmission_Gate_Layout_0.CLKB Transmission_Gate_Layout_0.CLKB.n31 0.510317
R6711 Transmission_Gate_Layout_12.VIN.n198 Transmission_Gate_Layout_12.VIN.n141 14.268
R6712 Transmission_Gate_Layout_12.VIN.n46 Transmission_Gate_Layout_12.VIN.t116 5.21612
R6713 Transmission_Gate_Layout_12.VIN.n184 Transmission_Gate_Layout_12.VIN.n182 5.21612
R6714 Transmission_Gate_Layout_12.VIN.n51 Transmission_Gate_Layout_12.VIN.n35 4.4609
R6715 Transmission_Gate_Layout_12.VIN.n50 Transmission_Gate_Layout_12.VIN.n36 4.4609
R6716 Transmission_Gate_Layout_12.VIN.n49 Transmission_Gate_Layout_12.VIN.n37 4.4609
R6717 Transmission_Gate_Layout_12.VIN.n47 Transmission_Gate_Layout_12.VIN.t74 4.4609
R6718 Transmission_Gate_Layout_12.VIN.n46 Transmission_Gate_Layout_12.VIN.t81 4.4609
R6719 Transmission_Gate_Layout_12.VIN.n190 Transmission_Gate_Layout_12.VIN.t1 4.4609
R6720 Transmission_Gate_Layout_12.VIN.n189 Transmission_Gate_Layout_12.VIN.t18 4.4609
R6721 Transmission_Gate_Layout_12.VIN.n188 Transmission_Gate_Layout_12.VIN.t9 4.4609
R6722 Transmission_Gate_Layout_12.VIN.n186 Transmission_Gate_Layout_12.VIN.n185 4.4609
R6723 Transmission_Gate_Layout_12.VIN.n184 Transmission_Gate_Layout_12.VIN.n183 4.4609
R6724 Transmission_Gate_Layout_12.VIN.n25 Transmission_Gate_Layout_12.VIN.n24 3.90572
R6725 Transmission_Gate_Layout_12.VIN.n33 Transmission_Gate_Layout_12.VIN.n32 3.90572
R6726 Transmission_Gate_Layout_12.VIN.n42 Transmission_Gate_Layout_12.VIN.n39 3.90572
R6727 Transmission_Gate_Layout_12.VIN.n103 Transmission_Gate_Layout_12.VIN.n100 3.90572
R6728 Transmission_Gate_Layout_12.VIN.n95 Transmission_Gate_Layout_12.VIN.n92 3.90572
R6729 Transmission_Gate_Layout_12.VIN.n125 Transmission_Gate_Layout_12.VIN.n124 3.90572
R6730 Transmission_Gate_Layout_12.VIN.n164 Transmission_Gate_Layout_12.VIN.n163 3.90572
R6731 Transmission_Gate_Layout_12.VIN.n178 Transmission_Gate_Layout_12.VIN.n175 3.90572
R6732 Transmission_Gate_Layout_12.VIN.n172 Transmission_Gate_Layout_12.VIN.n171 3.90572
R6733 Transmission_Gate_Layout_12.VIN.n7 Transmission_Gate_Layout_12.VIN.n4 3.84485
R6734 Transmission_Gate_Layout_12.VIN.n15 Transmission_Gate_Layout_12.VIN.n12 3.84485
R6735 Transmission_Gate_Layout_12.VIN.n65 Transmission_Gate_Layout_12.VIN.n64 3.84485
R6736 Transmission_Gate_Layout_12.VIN.n115 Transmission_Gate_Layout_12.VIN.n112 3.84485
R6737 Transmission_Gate_Layout_12.VIN.n77 Transmission_Gate_Layout_12.VIN.n76 3.84485
R6738 Transmission_Gate_Layout_12.VIN.n139 Transmission_Gate_Layout_12.VIN.n138 3.84485
R6739 Transmission_Gate_Layout_12.VIN.n154 Transmission_Gate_Layout_12.VIN.n151 3.84485
R6740 Transmission_Gate_Layout_12.VIN.n146 Transmission_Gate_Layout_12.VIN.n143 3.84485
R6741 Transmission_Gate_Layout_12.VIN.n205 Transmission_Gate_Layout_12.VIN.n204 3.84485
R6742 Transmission_Gate_Layout_12.VIN.n70 Transmission_Gate_Layout_12.VIN.t133 3.3285
R6743 Transmission_Gate_Layout_12.VIN.n68 Transmission_Gate_Layout_12.VIN.t130 3.3285
R6744 Transmission_Gate_Layout_12.VIN.n58 Transmission_Gate_Layout_12.VIN.n0 3.3285
R6745 Transmission_Gate_Layout_12.VIN.n57 Transmission_Gate_Layout_12.VIN.n1 3.3285
R6746 Transmission_Gate_Layout_12.VIN.n56 Transmission_Gate_Layout_12.VIN.n2 3.3285
R6747 Transmission_Gate_Layout_12.VIN.n209 Transmission_Gate_Layout_12.VIN.n208 3.3285
R6748 Transmission_Gate_Layout_12.VIN.n211 Transmission_Gate_Layout_12.VIN.n210 3.3285
R6749 Transmission_Gate_Layout_12.VIN.n213 Transmission_Gate_Layout_12.VIN.n212 3.3285
R6750 Transmission_Gate_Layout_12.VIN.n197 Transmission_Gate_Layout_12.VIN.t54 3.3285
R6751 Transmission_Gate_Layout_12.VIN.n196 Transmission_Gate_Layout_12.VIN.t56 3.3285
R6752 Transmission_Gate_Layout_12.VIN.n195 Transmission_Gate_Layout_12.VIN.t72 3.3285
R6753 Transmission_Gate_Layout_12.VIN.n69 Transmission_Gate_Layout_12.VIN.t140 3.3285
R6754 Transmission_Gate_Layout_12.VIN.n25 Transmission_Gate_Layout_12.VIN.n22 3.1505
R6755 Transmission_Gate_Layout_12.VIN.n26 Transmission_Gate_Layout_12.VIN.n20 3.1505
R6756 Transmission_Gate_Layout_12.VIN.n33 Transmission_Gate_Layout_12.VIN.n30 3.1505
R6757 Transmission_Gate_Layout_12.VIN.n34 Transmission_Gate_Layout_12.VIN.n28 3.1505
R6758 Transmission_Gate_Layout_12.VIN.n42 Transmission_Gate_Layout_12.VIN.n41 3.1505
R6759 Transmission_Gate_Layout_12.VIN.n45 Transmission_Gate_Layout_12.VIN.n44 3.1505
R6760 Transmission_Gate_Layout_12.VIN.n103 Transmission_Gate_Layout_12.VIN.n102 3.1505
R6761 Transmission_Gate_Layout_12.VIN.n106 Transmission_Gate_Layout_12.VIN.n105 3.1505
R6762 Transmission_Gate_Layout_12.VIN.n95 Transmission_Gate_Layout_12.VIN.n94 3.1505
R6763 Transmission_Gate_Layout_12.VIN.n98 Transmission_Gate_Layout_12.VIN.n97 3.1505
R6764 Transmission_Gate_Layout_12.VIN.n108 Transmission_Gate_Layout_12.VIN.n90 3.1505
R6765 Transmission_Gate_Layout_12.VIN.n109 Transmission_Gate_Layout_12.VIN.n88 3.1505
R6766 Transmission_Gate_Layout_12.VIN.n110 Transmission_Gate_Layout_12.VIN.n86 3.1505
R6767 Transmission_Gate_Layout_12.VIN.n125 Transmission_Gate_Layout_12.VIN.n122 3.1505
R6768 Transmission_Gate_Layout_12.VIN.n126 Transmission_Gate_Layout_12.VIN.n120 3.1505
R6769 Transmission_Gate_Layout_12.VIN.n164 Transmission_Gate_Layout_12.VIN.n161 3.1505
R6770 Transmission_Gate_Layout_12.VIN.n165 Transmission_Gate_Layout_12.VIN.n159 3.1505
R6771 Transmission_Gate_Layout_12.VIN.n178 Transmission_Gate_Layout_12.VIN.n177 3.1505
R6772 Transmission_Gate_Layout_12.VIN.n181 Transmission_Gate_Layout_12.VIN.n180 3.1505
R6773 Transmission_Gate_Layout_12.VIN.n172 Transmission_Gate_Layout_12.VIN.n169 3.1505
R6774 Transmission_Gate_Layout_12.VIN.n173 Transmission_Gate_Layout_12.VIN.n167 3.1505
R6775 Transmission_Gate_Layout_12.VIN.n67 Transmission_Gate_Layout_12.VIN.n58 2.72398
R6776 Transmission_Gate_Layout_12.VIN.n7 Transmission_Gate_Layout_12.VIN.n6 2.6005
R6777 Transmission_Gate_Layout_12.VIN.n10 Transmission_Gate_Layout_12.VIN.n9 2.6005
R6778 Transmission_Gate_Layout_12.VIN.n15 Transmission_Gate_Layout_12.VIN.n14 2.6005
R6779 Transmission_Gate_Layout_12.VIN.n18 Transmission_Gate_Layout_12.VIN.n17 2.6005
R6780 Transmission_Gate_Layout_12.VIN.n65 Transmission_Gate_Layout_12.VIN.n62 2.6005
R6781 Transmission_Gate_Layout_12.VIN.n66 Transmission_Gate_Layout_12.VIN.n60 2.6005
R6782 Transmission_Gate_Layout_12.VIN.n118 Transmission_Gate_Layout_12.VIN.n117 2.6005
R6783 Transmission_Gate_Layout_12.VIN.n115 Transmission_Gate_Layout_12.VIN.n114 2.6005
R6784 Transmission_Gate_Layout_12.VIN.n131 Transmission_Gate_Layout_12.VIN.n80 2.6005
R6785 Transmission_Gate_Layout_12.VIN.n130 Transmission_Gate_Layout_12.VIN.n82 2.6005
R6786 Transmission_Gate_Layout_12.VIN.n129 Transmission_Gate_Layout_12.VIN.n84 2.6005
R6787 Transmission_Gate_Layout_12.VIN.n77 Transmission_Gate_Layout_12.VIN.n74 2.6005
R6788 Transmission_Gate_Layout_12.VIN.n78 Transmission_Gate_Layout_12.VIN.n72 2.6005
R6789 Transmission_Gate_Layout_12.VIN.n139 Transmission_Gate_Layout_12.VIN.n136 2.6005
R6790 Transmission_Gate_Layout_12.VIN.n140 Transmission_Gate_Layout_12.VIN.n134 2.6005
R6791 Transmission_Gate_Layout_12.VIN.n154 Transmission_Gate_Layout_12.VIN.n153 2.6005
R6792 Transmission_Gate_Layout_12.VIN.n157 Transmission_Gate_Layout_12.VIN.n156 2.6005
R6793 Transmission_Gate_Layout_12.VIN.n146 Transmission_Gate_Layout_12.VIN.n145 2.6005
R6794 Transmission_Gate_Layout_12.VIN.n149 Transmission_Gate_Layout_12.VIN.n148 2.6005
R6795 Transmission_Gate_Layout_12.VIN.n205 Transmission_Gate_Layout_12.VIN.n202 2.6005
R6796 Transmission_Gate_Layout_12.VIN.n206 Transmission_Gate_Layout_12.VIN.n200 2.6005
R6797 Transmission_Gate_Layout_12.VIN.n49 Transmission_Gate_Layout_12.VIN.n48 2.47941
R6798 Transmission_Gate_Layout_12.VIN.n188 Transmission_Gate_Layout_12.VIN.n187 2.47941
R6799 Transmission_Gate_Layout_12.VIN.n207 Transmission_Gate_Layout_12.VIN.n198 2.10376
R6800 Transmission_Gate_Layout_12.VIN.n20 Transmission_Gate_Layout_12.VIN.t73 1.3109
R6801 Transmission_Gate_Layout_12.VIN.n20 Transmission_Gate_Layout_12.VIN.n19 1.3109
R6802 Transmission_Gate_Layout_12.VIN.n22 Transmission_Gate_Layout_12.VIN.t0 1.3109
R6803 Transmission_Gate_Layout_12.VIN.n22 Transmission_Gate_Layout_12.VIN.n21 1.3109
R6804 Transmission_Gate_Layout_12.VIN.n24 Transmission_Gate_Layout_12.VIN.t82 1.3109
R6805 Transmission_Gate_Layout_12.VIN.n24 Transmission_Gate_Layout_12.VIN.n23 1.3109
R6806 Transmission_Gate_Layout_12.VIN.n28 Transmission_Gate_Layout_12.VIN.t79 1.3109
R6807 Transmission_Gate_Layout_12.VIN.n28 Transmission_Gate_Layout_12.VIN.n27 1.3109
R6808 Transmission_Gate_Layout_12.VIN.n30 Transmission_Gate_Layout_12.VIN.t87 1.3109
R6809 Transmission_Gate_Layout_12.VIN.n30 Transmission_Gate_Layout_12.VIN.n29 1.3109
R6810 Transmission_Gate_Layout_12.VIN.n32 Transmission_Gate_Layout_12.VIN.t115 1.3109
R6811 Transmission_Gate_Layout_12.VIN.n32 Transmission_Gate_Layout_12.VIN.n31 1.3109
R6812 Transmission_Gate_Layout_12.VIN.n44 Transmission_Gate_Layout_12.VIN.t78 1.3109
R6813 Transmission_Gate_Layout_12.VIN.n44 Transmission_Gate_Layout_12.VIN.n43 1.3109
R6814 Transmission_Gate_Layout_12.VIN.n41 Transmission_Gate_Layout_12.VIN.t114 1.3109
R6815 Transmission_Gate_Layout_12.VIN.n41 Transmission_Gate_Layout_12.VIN.n40 1.3109
R6816 Transmission_Gate_Layout_12.VIN.n39 Transmission_Gate_Layout_12.VIN.t85 1.3109
R6817 Transmission_Gate_Layout_12.VIN.n39 Transmission_Gate_Layout_12.VIN.n38 1.3109
R6818 Transmission_Gate_Layout_12.VIN.n86 Transmission_Gate_Layout_12.VIN.t89 1.3109
R6819 Transmission_Gate_Layout_12.VIN.n86 Transmission_Gate_Layout_12.VIN.n85 1.3109
R6820 Transmission_Gate_Layout_12.VIN.n88 Transmission_Gate_Layout_12.VIN.t105 1.3109
R6821 Transmission_Gate_Layout_12.VIN.n88 Transmission_Gate_Layout_12.VIN.n87 1.3109
R6822 Transmission_Gate_Layout_12.VIN.n90 Transmission_Gate_Layout_12.VIN.t97 1.3109
R6823 Transmission_Gate_Layout_12.VIN.n90 Transmission_Gate_Layout_12.VIN.n89 1.3109
R6824 Transmission_Gate_Layout_12.VIN.n105 Transmission_Gate_Layout_12.VIN.t101 1.3109
R6825 Transmission_Gate_Layout_12.VIN.n105 Transmission_Gate_Layout_12.VIN.n104 1.3109
R6826 Transmission_Gate_Layout_12.VIN.n102 Transmission_Gate_Layout_12.VIN.t109 1.3109
R6827 Transmission_Gate_Layout_12.VIN.n102 Transmission_Gate_Layout_12.VIN.n101 1.3109
R6828 Transmission_Gate_Layout_12.VIN.n100 Transmission_Gate_Layout_12.VIN.t93 1.3109
R6829 Transmission_Gate_Layout_12.VIN.n100 Transmission_Gate_Layout_12.VIN.n99 1.3109
R6830 Transmission_Gate_Layout_12.VIN.n97 Transmission_Gate_Layout_12.VIN.t106 1.3109
R6831 Transmission_Gate_Layout_12.VIN.n97 Transmission_Gate_Layout_12.VIN.n96 1.3109
R6832 Transmission_Gate_Layout_12.VIN.n94 Transmission_Gate_Layout_12.VIN.t91 1.3109
R6833 Transmission_Gate_Layout_12.VIN.n94 Transmission_Gate_Layout_12.VIN.n93 1.3109
R6834 Transmission_Gate_Layout_12.VIN.n92 Transmission_Gate_Layout_12.VIN.t98 1.3109
R6835 Transmission_Gate_Layout_12.VIN.n92 Transmission_Gate_Layout_12.VIN.n91 1.3109
R6836 Transmission_Gate_Layout_12.VIN.n120 Transmission_Gate_Layout_12.VIN.t90 1.3109
R6837 Transmission_Gate_Layout_12.VIN.n120 Transmission_Gate_Layout_12.VIN.n119 1.3109
R6838 Transmission_Gate_Layout_12.VIN.n122 Transmission_Gate_Layout_12.VIN.t108 1.3109
R6839 Transmission_Gate_Layout_12.VIN.n122 Transmission_Gate_Layout_12.VIN.n121 1.3109
R6840 Transmission_Gate_Layout_12.VIN.n124 Transmission_Gate_Layout_12.VIN.t100 1.3109
R6841 Transmission_Gate_Layout_12.VIN.n124 Transmission_Gate_Layout_12.VIN.n123 1.3109
R6842 Transmission_Gate_Layout_12.VIN.n159 Transmission_Gate_Layout_12.VIN.t13 1.3109
R6843 Transmission_Gate_Layout_12.VIN.n159 Transmission_Gate_Layout_12.VIN.n158 1.3109
R6844 Transmission_Gate_Layout_12.VIN.n161 Transmission_Gate_Layout_12.VIN.t5 1.3109
R6845 Transmission_Gate_Layout_12.VIN.n161 Transmission_Gate_Layout_12.VIN.n160 1.3109
R6846 Transmission_Gate_Layout_12.VIN.n163 Transmission_Gate_Layout_12.VIN.t21 1.3109
R6847 Transmission_Gate_Layout_12.VIN.n163 Transmission_Gate_Layout_12.VIN.n162 1.3109
R6848 Transmission_Gate_Layout_12.VIN.n180 Transmission_Gate_Layout_12.VIN.t23 1.3109
R6849 Transmission_Gate_Layout_12.VIN.n180 Transmission_Gate_Layout_12.VIN.n179 1.3109
R6850 Transmission_Gate_Layout_12.VIN.n177 Transmission_Gate_Layout_12.VIN.t8 1.3109
R6851 Transmission_Gate_Layout_12.VIN.n177 Transmission_Gate_Layout_12.VIN.n176 1.3109
R6852 Transmission_Gate_Layout_12.VIN.n175 Transmission_Gate_Layout_12.VIN.t14 1.3109
R6853 Transmission_Gate_Layout_12.VIN.n175 Transmission_Gate_Layout_12.VIN.n174 1.3109
R6854 Transmission_Gate_Layout_12.VIN.n167 Transmission_Gate_Layout_12.VIN.t6 1.3109
R6855 Transmission_Gate_Layout_12.VIN.n167 Transmission_Gate_Layout_12.VIN.n166 1.3109
R6856 Transmission_Gate_Layout_12.VIN.n169 Transmission_Gate_Layout_12.VIN.t22 1.3109
R6857 Transmission_Gate_Layout_12.VIN.n169 Transmission_Gate_Layout_12.VIN.n168 1.3109
R6858 Transmission_Gate_Layout_12.VIN.n171 Transmission_Gate_Layout_12.VIN.t15 1.3109
R6859 Transmission_Gate_Layout_12.VIN.n171 Transmission_Gate_Layout_12.VIN.n170 1.3109
R6860 Transmission_Gate_Layout_12.VIN.n10 Transmission_Gate_Layout_12.VIN.n7 1.24485
R6861 Transmission_Gate_Layout_12.VIN.n18 Transmission_Gate_Layout_12.VIN.n15 1.24485
R6862 Transmission_Gate_Layout_12.VIN.n58 Transmission_Gate_Layout_12.VIN.n57 1.24485
R6863 Transmission_Gate_Layout_12.VIN.n57 Transmission_Gate_Layout_12.VIN.n56 1.24485
R6864 Transmission_Gate_Layout_12.VIN.n66 Transmission_Gate_Layout_12.VIN.n65 1.24485
R6865 Transmission_Gate_Layout_12.VIN.n118 Transmission_Gate_Layout_12.VIN.n115 1.24485
R6866 Transmission_Gate_Layout_12.VIN.n131 Transmission_Gate_Layout_12.VIN.n130 1.24485
R6867 Transmission_Gate_Layout_12.VIN.n130 Transmission_Gate_Layout_12.VIN.n129 1.24485
R6868 Transmission_Gate_Layout_12.VIN.n78 Transmission_Gate_Layout_12.VIN.n77 1.24485
R6869 Transmission_Gate_Layout_12.VIN.n140 Transmission_Gate_Layout_12.VIN.n139 1.24485
R6870 Transmission_Gate_Layout_12.VIN.n157 Transmission_Gate_Layout_12.VIN.n154 1.24485
R6871 Transmission_Gate_Layout_12.VIN.n149 Transmission_Gate_Layout_12.VIN.n146 1.24485
R6872 Transmission_Gate_Layout_12.VIN.n197 Transmission_Gate_Layout_12.VIN.n196 1.24485
R6873 Transmission_Gate_Layout_12.VIN.n196 Transmission_Gate_Layout_12.VIN.n195 1.24485
R6874 Transmission_Gate_Layout_12.VIN.n206 Transmission_Gate_Layout_12.VIN.n205 1.24485
R6875 Transmission_Gate_Layout_12.VIN.n211 Transmission_Gate_Layout_12.VIN.n209 1.24485
R6876 Transmission_Gate_Layout_12.VIN.n213 Transmission_Gate_Layout_12.VIN.n211 1.24485
R6877 Transmission_Gate_Layout_12.VIN.n69 Transmission_Gate_Layout_12.VIN.n68 1.24485
R6878 Transmission_Gate_Layout_12.VIN.n70 Transmission_Gate_Layout_12.VIN.n69 1.24485
R6879 Transmission_Gate_Layout_12.VIN.n56 Transmission_Gate_Layout_12.VIN.n55 1.2018
R6880 Transmission_Gate_Layout_12.VIN.n68 Transmission_Gate_Layout_12.VIN.n67 1.2018
R6881 Transmission_Gate_Layout_12.VIN.n132 Transmission_Gate_Layout_12.VIN.n131 1.2018
R6882 Transmission_Gate_Layout_12.VIN.n195 Transmission_Gate_Layout_12.VIN.n194 1.2018
R6883 Transmission_Gate_Layout_12.VIN.n209 Transmission_Gate_Layout_12.VIN.n207 1.2018
R6884 Transmission_Gate_Layout_12.VIN.n48 Transmission_Gate_Layout_12.VIN.n47 0.957239
R6885 Transmission_Gate_Layout_12.VIN.n52 Transmission_Gate_Layout_12.VIN.n51 0.957239
R6886 Transmission_Gate_Layout_12.VIN.n107 Transmission_Gate_Layout_12.VIN.n106 0.957239
R6887 Transmission_Gate_Layout_12.VIN.n108 Transmission_Gate_Layout_12.VIN.n107 0.957239
R6888 Transmission_Gate_Layout_12.VIN.n187 Transmission_Gate_Layout_12.VIN.n186 0.957239
R6889 Transmission_Gate_Layout_12.VIN.n191 Transmission_Gate_Layout_12.VIN.n190 0.957239
R6890 Transmission_Gate_Layout_12.VIN.n127 Transmission_Gate_Layout_12.VIN.n118 0.806587
R6891 Transmission_Gate_Layout_12.VIN.n129 Transmission_Gate_Layout_12.VIN.n128 0.806587
R6892 Transmission_Gate_Layout_12.VIN.n26 Transmission_Gate_Layout_12.VIN.n25 0.755717
R6893 Transmission_Gate_Layout_12.VIN.n34 Transmission_Gate_Layout_12.VIN.n33 0.755717
R6894 Transmission_Gate_Layout_12.VIN.n45 Transmission_Gate_Layout_12.VIN.n42 0.755717
R6895 Transmission_Gate_Layout_12.VIN.n47 Transmission_Gate_Layout_12.VIN.n46 0.755717
R6896 Transmission_Gate_Layout_12.VIN.n51 Transmission_Gate_Layout_12.VIN.n50 0.755717
R6897 Transmission_Gate_Layout_12.VIN.n50 Transmission_Gate_Layout_12.VIN.n49 0.755717
R6898 Transmission_Gate_Layout_12.VIN.n106 Transmission_Gate_Layout_12.VIN.n103 0.755717
R6899 Transmission_Gate_Layout_12.VIN.n98 Transmission_Gate_Layout_12.VIN.n95 0.755717
R6900 Transmission_Gate_Layout_12.VIN.n110 Transmission_Gate_Layout_12.VIN.n109 0.755717
R6901 Transmission_Gate_Layout_12.VIN.n109 Transmission_Gate_Layout_12.VIN.n108 0.755717
R6902 Transmission_Gate_Layout_12.VIN.n126 Transmission_Gate_Layout_12.VIN.n125 0.755717
R6903 Transmission_Gate_Layout_12.VIN.n165 Transmission_Gate_Layout_12.VIN.n164 0.755717
R6904 Transmission_Gate_Layout_12.VIN.n181 Transmission_Gate_Layout_12.VIN.n178 0.755717
R6905 Transmission_Gate_Layout_12.VIN.n186 Transmission_Gate_Layout_12.VIN.n184 0.755717
R6906 Transmission_Gate_Layout_12.VIN.n190 Transmission_Gate_Layout_12.VIN.n189 0.755717
R6907 Transmission_Gate_Layout_12.VIN.n189 Transmission_Gate_Layout_12.VIN.n188 0.755717
R6908 Transmission_Gate_Layout_12.VIN.n173 Transmission_Gate_Layout_12.VIN.n172 0.755717
R6909 Transmission_Gate_Layout_12.VIN.n60 Transmission_Gate_Layout_12.VIN.t139 0.7285
R6910 Transmission_Gate_Layout_12.VIN.n60 Transmission_Gate_Layout_12.VIN.n59 0.7285
R6911 Transmission_Gate_Layout_12.VIN.n62 Transmission_Gate_Layout_12.VIN.t137 0.7285
R6912 Transmission_Gate_Layout_12.VIN.n62 Transmission_Gate_Layout_12.VIN.n61 0.7285
R6913 Transmission_Gate_Layout_12.VIN.n64 Transmission_Gate_Layout_12.VIN.t131 0.7285
R6914 Transmission_Gate_Layout_12.VIN.n64 Transmission_Gate_Layout_12.VIN.n63 0.7285
R6915 Transmission_Gate_Layout_12.VIN.n9 Transmission_Gate_Layout_12.VIN.t138 0.7285
R6916 Transmission_Gate_Layout_12.VIN.n9 Transmission_Gate_Layout_12.VIN.n8 0.7285
R6917 Transmission_Gate_Layout_12.VIN.n6 Transmission_Gate_Layout_12.VIN.t132 0.7285
R6918 Transmission_Gate_Layout_12.VIN.n6 Transmission_Gate_Layout_12.VIN.n5 0.7285
R6919 Transmission_Gate_Layout_12.VIN.n4 Transmission_Gate_Layout_12.VIN.t134 0.7285
R6920 Transmission_Gate_Layout_12.VIN.n4 Transmission_Gate_Layout_12.VIN.n3 0.7285
R6921 Transmission_Gate_Layout_12.VIN.n17 Transmission_Gate_Layout_12.VIN.t129 0.7285
R6922 Transmission_Gate_Layout_12.VIN.n17 Transmission_Gate_Layout_12.VIN.n16 0.7285
R6923 Transmission_Gate_Layout_12.VIN.n14 Transmission_Gate_Layout_12.VIN.t135 0.7285
R6924 Transmission_Gate_Layout_12.VIN.n14 Transmission_Gate_Layout_12.VIN.n13 0.7285
R6925 Transmission_Gate_Layout_12.VIN.n12 Transmission_Gate_Layout_12.VIN.t136 0.7285
R6926 Transmission_Gate_Layout_12.VIN.n12 Transmission_Gate_Layout_12.VIN.n11 0.7285
R6927 Transmission_Gate_Layout_12.VIN.n200 Transmission_Gate_Layout_12.VIN.t71 0.7285
R6928 Transmission_Gate_Layout_12.VIN.n200 Transmission_Gate_Layout_12.VIN.n199 0.7285
R6929 Transmission_Gate_Layout_12.VIN.n202 Transmission_Gate_Layout_12.VIN.t49 0.7285
R6930 Transmission_Gate_Layout_12.VIN.n202 Transmission_Gate_Layout_12.VIN.n201 0.7285
R6931 Transmission_Gate_Layout_12.VIN.n204 Transmission_Gate_Layout_12.VIN.t60 0.7285
R6932 Transmission_Gate_Layout_12.VIN.n204 Transmission_Gate_Layout_12.VIN.n203 0.7285
R6933 Transmission_Gate_Layout_12.VIN.n84 Transmission_Gate_Layout_12.VIN.t26 0.7285
R6934 Transmission_Gate_Layout_12.VIN.n84 Transmission_Gate_Layout_12.VIN.n83 0.7285
R6935 Transmission_Gate_Layout_12.VIN.n82 Transmission_Gate_Layout_12.VIN.t34 0.7285
R6936 Transmission_Gate_Layout_12.VIN.n82 Transmission_Gate_Layout_12.VIN.n81 0.7285
R6937 Transmission_Gate_Layout_12.VIN.n80 Transmission_Gate_Layout_12.VIN.t48 0.7285
R6938 Transmission_Gate_Layout_12.VIN.n80 Transmission_Gate_Layout_12.VIN.n79 0.7285
R6939 Transmission_Gate_Layout_12.VIN.n112 Transmission_Gate_Layout_12.VIN.t36 0.7285
R6940 Transmission_Gate_Layout_12.VIN.n112 Transmission_Gate_Layout_12.VIN.n111 0.7285
R6941 Transmission_Gate_Layout_12.VIN.n114 Transmission_Gate_Layout_12.VIN.t38 0.7285
R6942 Transmission_Gate_Layout_12.VIN.n114 Transmission_Gate_Layout_12.VIN.n113 0.7285
R6943 Transmission_Gate_Layout_12.VIN.n117 Transmission_Gate_Layout_12.VIN.t28 0.7285
R6944 Transmission_Gate_Layout_12.VIN.n117 Transmission_Gate_Layout_12.VIN.n116 0.7285
R6945 Transmission_Gate_Layout_12.VIN.n72 Transmission_Gate_Layout_12.VIN.t43 0.7285
R6946 Transmission_Gate_Layout_12.VIN.n72 Transmission_Gate_Layout_12.VIN.n71 0.7285
R6947 Transmission_Gate_Layout_12.VIN.n74 Transmission_Gate_Layout_12.VIN.t45 0.7285
R6948 Transmission_Gate_Layout_12.VIN.n74 Transmission_Gate_Layout_12.VIN.n73 0.7285
R6949 Transmission_Gate_Layout_12.VIN.n76 Transmission_Gate_Layout_12.VIN.t33 0.7285
R6950 Transmission_Gate_Layout_12.VIN.n76 Transmission_Gate_Layout_12.VIN.n75 0.7285
R6951 Transmission_Gate_Layout_12.VIN.n134 Transmission_Gate_Layout_12.VIN.t37 0.7285
R6952 Transmission_Gate_Layout_12.VIN.n134 Transmission_Gate_Layout_12.VIN.n133 0.7285
R6953 Transmission_Gate_Layout_12.VIN.n136 Transmission_Gate_Layout_12.VIN.t41 0.7285
R6954 Transmission_Gate_Layout_12.VIN.n136 Transmission_Gate_Layout_12.VIN.n135 0.7285
R6955 Transmission_Gate_Layout_12.VIN.n138 Transmission_Gate_Layout_12.VIN.t29 0.7285
R6956 Transmission_Gate_Layout_12.VIN.n138 Transmission_Gate_Layout_12.VIN.n137 0.7285
R6957 Transmission_Gate_Layout_12.VIN.n156 Transmission_Gate_Layout_12.VIN.t58 0.7285
R6958 Transmission_Gate_Layout_12.VIN.n156 Transmission_Gate_Layout_12.VIN.n155 0.7285
R6959 Transmission_Gate_Layout_12.VIN.n153 Transmission_Gate_Layout_12.VIN.t70 0.7285
R6960 Transmission_Gate_Layout_12.VIN.n153 Transmission_Gate_Layout_12.VIN.n152 0.7285
R6961 Transmission_Gate_Layout_12.VIN.n151 Transmission_Gate_Layout_12.VIN.t68 0.7285
R6962 Transmission_Gate_Layout_12.VIN.n151 Transmission_Gate_Layout_12.VIN.n150 0.7285
R6963 Transmission_Gate_Layout_12.VIN.n148 Transmission_Gate_Layout_12.VIN.t52 0.7285
R6964 Transmission_Gate_Layout_12.VIN.n148 Transmission_Gate_Layout_12.VIN.n147 0.7285
R6965 Transmission_Gate_Layout_12.VIN.n145 Transmission_Gate_Layout_12.VIN.t62 0.7285
R6966 Transmission_Gate_Layout_12.VIN.n145 Transmission_Gate_Layout_12.VIN.n144 0.7285
R6967 Transmission_Gate_Layout_12.VIN.n143 Transmission_Gate_Layout_12.VIN.t59 0.7285
R6968 Transmission_Gate_Layout_12.VIN.n143 Transmission_Gate_Layout_12.VIN.n142 0.7285
R6969 Transmission_Gate_Layout_12.VIN.n53 Transmission_Gate_Layout_12.VIN.n52 0.626587
R6970 Transmission_Gate_Layout_12.VIN.n55 Transmission_Gate_Layout_12.VIN.n54 0.626587
R6971 Transmission_Gate_Layout_12.VIN.n128 Transmission_Gate_Layout_12.VIN.n127 0.626587
R6972 Transmission_Gate_Layout_12.VIN.n192 Transmission_Gate_Layout_12.VIN.n191 0.626587
R6973 Transmission_Gate_Layout_12.VIN.n194 Transmission_Gate_Layout_12.VIN.n193 0.626587
R6974 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.VIN.n213 0.607022
R6975 Transmission_Gate_Layout_12.VIN Transmission_Gate_Layout_12.VIN.n70 0.607022
R6976 Transmission_Gate_Layout_12.VIN.n55 Transmission_Gate_Layout_12.VIN.n10 0.575717
R6977 Transmission_Gate_Layout_12.VIN.n54 Transmission_Gate_Layout_12.VIN.n18 0.575717
R6978 Transmission_Gate_Layout_12.VIN.n67 Transmission_Gate_Layout_12.VIN.n66 0.575717
R6979 Transmission_Gate_Layout_12.VIN.n132 Transmission_Gate_Layout_12.VIN.n78 0.575717
R6980 Transmission_Gate_Layout_12.VIN.n193 Transmission_Gate_Layout_12.VIN.n157 0.575717
R6981 Transmission_Gate_Layout_12.VIN.n194 Transmission_Gate_Layout_12.VIN.n149 0.575717
R6982 Transmission_Gate_Layout_12.VIN.n207 Transmission_Gate_Layout_12.VIN.n206 0.575717
R6983 Transmission_Gate_Layout_12.VIN.n141 Transmission_Gate_Layout_12.VIN.n132 0.570002
R6984 Transmission_Gate_Layout_12.VIN.n141 Transmission_Gate_Layout_12.VIN.n140 0.562022
R6985 Transmission_Gate_Layout_12.VIN.n198 Transmission_Gate_Layout_12.VIN.n197 0.562022
R6986 Transmission_Gate_Layout_12.VIN.n128 Transmission_Gate_Layout_12.VIN.n110 0.428978
R6987 Transmission_Gate_Layout_12.VIN.n127 Transmission_Gate_Layout_12.VIN.n126 0.428978
R6988 Transmission_Gate_Layout_12.VIN.n53 Transmission_Gate_Layout_12.VIN.n26 0.331152
R6989 Transmission_Gate_Layout_12.VIN.n52 Transmission_Gate_Layout_12.VIN.n34 0.331152
R6990 Transmission_Gate_Layout_12.VIN.n48 Transmission_Gate_Layout_12.VIN.n45 0.331152
R6991 Transmission_Gate_Layout_12.VIN.n107 Transmission_Gate_Layout_12.VIN.n98 0.331152
R6992 Transmission_Gate_Layout_12.VIN.n192 Transmission_Gate_Layout_12.VIN.n165 0.331152
R6993 Transmission_Gate_Layout_12.VIN.n187 Transmission_Gate_Layout_12.VIN.n181 0.331152
R6994 Transmission_Gate_Layout_12.VIN.n191 Transmission_Gate_Layout_12.VIN.n173 0.331152
R6995 Transmission_Gate_Layout_12.VIN.n54 Transmission_Gate_Layout_12.VIN.n53 0.239196
R6996 Transmission_Gate_Layout_12.VIN.n193 Transmission_Gate_Layout_12.VIN.n192 0.239196
R6997 Transmission_Gate_Layout_12.VIN.n127 Transmission_Gate_Layout_12.VIN 0.192239
R6998 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.VOUT.n212 8.51067
R6999 Transmission_Gate_Layout_9.VOUT.n116 Transmission_Gate_Layout_9.VOUT.n115 5.21612
R7000 Transmission_Gate_Layout_9.VOUT.n184 Transmission_Gate_Layout_9.VOUT.t15 5.21612
R7001 Transmission_Gate_Layout_9.VOUT.n119 Transmission_Gate_Layout_9.VOUT.t92 4.4609
R7002 Transmission_Gate_Layout_9.VOUT.n120 Transmission_Gate_Layout_9.VOUT.t95 4.4609
R7003 Transmission_Gate_Layout_9.VOUT.n121 Transmission_Gate_Layout_9.VOUT.t89 4.4609
R7004 Transmission_Gate_Layout_9.VOUT.n117 Transmission_Gate_Layout_9.VOUT.n113 4.4609
R7005 Transmission_Gate_Layout_9.VOUT.n116 Transmission_Gate_Layout_9.VOUT.n114 4.4609
R7006 Transmission_Gate_Layout_9.VOUT.n192 Transmission_Gate_Layout_9.VOUT.n191 4.4609
R7007 Transmission_Gate_Layout_9.VOUT.n190 Transmission_Gate_Layout_9.VOUT.n189 4.4609
R7008 Transmission_Gate_Layout_9.VOUT.n188 Transmission_Gate_Layout_9.VOUT.n187 4.4609
R7009 Transmission_Gate_Layout_9.VOUT.n185 Transmission_Gate_Layout_9.VOUT.t21 4.4609
R7010 Transmission_Gate_Layout_9.VOUT.n184 Transmission_Gate_Layout_9.VOUT.t12 4.4609
R7011 Transmission_Gate_Layout_9.VOUT.n6 Transmission_Gate_Layout_9.VOUT.n5 3.90572
R7012 Transmission_Gate_Layout_9.VOUT.n93 Transmission_Gate_Layout_9.VOUT.n90 3.90572
R7013 Transmission_Gate_Layout_9.VOUT.n101 Transmission_Gate_Layout_9.VOUT.n98 3.90572
R7014 Transmission_Gate_Layout_9.VOUT.n111 Transmission_Gate_Layout_9.VOUT.n110 3.90572
R7015 Transmission_Gate_Layout_9.VOUT.n164 Transmission_Gate_Layout_9.VOUT.n161 3.90572
R7016 Transmission_Gate_Layout_9.VOUT.n182 Transmission_Gate_Layout_9.VOUT.n181 3.90572
R7017 Transmission_Gate_Layout_9.VOUT.n172 Transmission_Gate_Layout_9.VOUT.n169 3.90572
R7018 Transmission_Gate_Layout_9.VOUT.n52 Transmission_Gate_Layout_9.VOUT.n49 3.90572
R7019 Transmission_Gate_Layout_9.VOUT.n44 Transmission_Gate_Layout_9.VOUT.n41 3.90572
R7020 Transmission_Gate_Layout_9.VOUT.n130 Transmission_Gate_Layout_9.VOUT.n129 3.84485
R7021 Transmission_Gate_Layout_9.VOUT.n87 Transmission_Gate_Layout_9.VOUT.n86 3.84485
R7022 Transmission_Gate_Layout_9.VOUT.n77 Transmission_Gate_Layout_9.VOUT.n74 3.84485
R7023 Transmission_Gate_Layout_9.VOUT.n201 Transmission_Gate_Layout_9.VOUT.n200 3.84485
R7024 Transmission_Gate_Layout_9.VOUT.n158 Transmission_Gate_Layout_9.VOUT.n157 3.84485
R7025 Transmission_Gate_Layout_9.VOUT.n148 Transmission_Gate_Layout_9.VOUT.n145 3.84485
R7026 Transmission_Gate_Layout_9.VOUT.n14 Transmission_Gate_Layout_9.VOUT.n13 3.84485
R7027 Transmission_Gate_Layout_9.VOUT.n22 Transmission_Gate_Layout_9.VOUT.n21 3.84485
R7028 Transmission_Gate_Layout_9.VOUT.n65 Transmission_Gate_Layout_9.VOUT.n62 3.84485
R7029 Transmission_Gate_Layout_9.VOUT.n141 Transmission_Gate_Layout_9.VOUT.t52 3.3285
R7030 Transmission_Gate_Layout_9.VOUT.n142 Transmission_Gate_Layout_9.VOUT.t60 3.3285
R7031 Transmission_Gate_Layout_9.VOUT.n143 Transmission_Gate_Layout_9.VOUT.t69 3.3285
R7032 Transmission_Gate_Layout_9.VOUT.n138 Transmission_Gate_Layout_9.VOUT.n72 3.3285
R7033 Transmission_Gate_Layout_9.VOUT.n139 Transmission_Gate_Layout_9.VOUT.n71 3.3285
R7034 Transmission_Gate_Layout_9.VOUT.n140 Transmission_Gate_Layout_9.VOUT.n70 3.3285
R7035 Transmission_Gate_Layout_9.VOUT.n134 Transmission_Gate_Layout_9.VOUT.t115 3.3285
R7036 Transmission_Gate_Layout_9.VOUT.n135 Transmission_Gate_Layout_9.VOUT.t5 3.3285
R7037 Transmission_Gate_Layout_9.VOUT.n136 Transmission_Gate_Layout_9.VOUT.t77 3.3285
R7038 Transmission_Gate_Layout_9.VOUT.n210 Transmission_Gate_Layout_9.VOUT.n209 3.3285
R7039 Transmission_Gate_Layout_9.VOUT.n208 Transmission_Gate_Layout_9.VOUT.n207 3.3285
R7040 Transmission_Gate_Layout_9.VOUT.n206 Transmission_Gate_Layout_9.VOUT.n205 3.3285
R7041 Transmission_Gate_Layout_9.VOUT.n6 Transmission_Gate_Layout_9.VOUT.n3 3.1505
R7042 Transmission_Gate_Layout_9.VOUT.n7 Transmission_Gate_Layout_9.VOUT.n1 3.1505
R7043 Transmission_Gate_Layout_9.VOUT.n93 Transmission_Gate_Layout_9.VOUT.n92 3.1505
R7044 Transmission_Gate_Layout_9.VOUT.n96 Transmission_Gate_Layout_9.VOUT.n95 3.1505
R7045 Transmission_Gate_Layout_9.VOUT.n101 Transmission_Gate_Layout_9.VOUT.n100 3.1505
R7046 Transmission_Gate_Layout_9.VOUT.n104 Transmission_Gate_Layout_9.VOUT.n103 3.1505
R7047 Transmission_Gate_Layout_9.VOUT.n111 Transmission_Gate_Layout_9.VOUT.n108 3.1505
R7048 Transmission_Gate_Layout_9.VOUT.n112 Transmission_Gate_Layout_9.VOUT.n106 3.1505
R7049 Transmission_Gate_Layout_9.VOUT.n164 Transmission_Gate_Layout_9.VOUT.n163 3.1505
R7050 Transmission_Gate_Layout_9.VOUT.n167 Transmission_Gate_Layout_9.VOUT.n166 3.1505
R7051 Transmission_Gate_Layout_9.VOUT.n182 Transmission_Gate_Layout_9.VOUT.n179 3.1505
R7052 Transmission_Gate_Layout_9.VOUT.n183 Transmission_Gate_Layout_9.VOUT.n177 3.1505
R7053 Transmission_Gate_Layout_9.VOUT.n172 Transmission_Gate_Layout_9.VOUT.n171 3.1505
R7054 Transmission_Gate_Layout_9.VOUT.n175 Transmission_Gate_Layout_9.VOUT.n174 3.1505
R7055 Transmission_Gate_Layout_9.VOUT.n52 Transmission_Gate_Layout_9.VOUT.n51 3.1505
R7056 Transmission_Gate_Layout_9.VOUT.n55 Transmission_Gate_Layout_9.VOUT.n54 3.1505
R7057 Transmission_Gate_Layout_9.VOUT.n44 Transmission_Gate_Layout_9.VOUT.n43 3.1505
R7058 Transmission_Gate_Layout_9.VOUT.n47 Transmission_Gate_Layout_9.VOUT.n46 3.1505
R7059 Transmission_Gate_Layout_9.VOUT.n57 Transmission_Gate_Layout_9.VOUT.n39 3.1505
R7060 Transmission_Gate_Layout_9.VOUT.n58 Transmission_Gate_Layout_9.VOUT.n37 3.1505
R7061 Transmission_Gate_Layout_9.VOUT.n59 Transmission_Gate_Layout_9.VOUT.n35 3.1505
R7062 Transmission_Gate_Layout_9.VOUT.n137 Transmission_Gate_Layout_9.VOUT.n136 2.72398
R7063 Transmission_Gate_Layout_9.VOUT.n211 Transmission_Gate_Layout_9.VOUT.n210 2.72398
R7064 Transmission_Gate_Layout_9.VOUT.n130 Transmission_Gate_Layout_9.VOUT.n127 2.6005
R7065 Transmission_Gate_Layout_9.VOUT.n131 Transmission_Gate_Layout_9.VOUT.n125 2.6005
R7066 Transmission_Gate_Layout_9.VOUT.n87 Transmission_Gate_Layout_9.VOUT.n84 2.6005
R7067 Transmission_Gate_Layout_9.VOUT.n88 Transmission_Gate_Layout_9.VOUT.n82 2.6005
R7068 Transmission_Gate_Layout_9.VOUT.n77 Transmission_Gate_Layout_9.VOUT.n76 2.6005
R7069 Transmission_Gate_Layout_9.VOUT.n80 Transmission_Gate_Layout_9.VOUT.n79 2.6005
R7070 Transmission_Gate_Layout_9.VOUT.n201 Transmission_Gate_Layout_9.VOUT.n198 2.6005
R7071 Transmission_Gate_Layout_9.VOUT.n202 Transmission_Gate_Layout_9.VOUT.n196 2.6005
R7072 Transmission_Gate_Layout_9.VOUT.n158 Transmission_Gate_Layout_9.VOUT.n155 2.6005
R7073 Transmission_Gate_Layout_9.VOUT.n159 Transmission_Gate_Layout_9.VOUT.n153 2.6005
R7074 Transmission_Gate_Layout_9.VOUT.n148 Transmission_Gate_Layout_9.VOUT.n147 2.6005
R7075 Transmission_Gate_Layout_9.VOUT.n151 Transmission_Gate_Layout_9.VOUT.n150 2.6005
R7076 Transmission_Gate_Layout_9.VOUT.n14 Transmission_Gate_Layout_9.VOUT.n11 2.6005
R7077 Transmission_Gate_Layout_9.VOUT.n15 Transmission_Gate_Layout_9.VOUT.n9 2.6005
R7078 Transmission_Gate_Layout_9.VOUT.n22 Transmission_Gate_Layout_9.VOUT.n19 2.6005
R7079 Transmission_Gate_Layout_9.VOUT.n23 Transmission_Gate_Layout_9.VOUT.n17 2.6005
R7080 Transmission_Gate_Layout_9.VOUT.n27 Transmission_Gate_Layout_9.VOUT.n26 2.6005
R7081 Transmission_Gate_Layout_9.VOUT.n30 Transmission_Gate_Layout_9.VOUT.n29 2.6005
R7082 Transmission_Gate_Layout_9.VOUT.n33 Transmission_Gate_Layout_9.VOUT.n32 2.6005
R7083 Transmission_Gate_Layout_9.VOUT.n68 Transmission_Gate_Layout_9.VOUT.n67 2.6005
R7084 Transmission_Gate_Layout_9.VOUT.n65 Transmission_Gate_Layout_9.VOUT.n64 2.6005
R7085 Transmission_Gate_Layout_9.VOUT.n119 Transmission_Gate_Layout_9.VOUT.n118 2.47941
R7086 Transmission_Gate_Layout_9.VOUT.n188 Transmission_Gate_Layout_9.VOUT.n186 2.47941
R7087 Transmission_Gate_Layout_9.VOUT.n1 Transmission_Gate_Layout_9.VOUT.t37 1.3109
R7088 Transmission_Gate_Layout_9.VOUT.n1 Transmission_Gate_Layout_9.VOUT.n0 1.3109
R7089 Transmission_Gate_Layout_9.VOUT.n3 Transmission_Gate_Layout_9.VOUT.t142 1.3109
R7090 Transmission_Gate_Layout_9.VOUT.n3 Transmission_Gate_Layout_9.VOUT.n2 1.3109
R7091 Transmission_Gate_Layout_9.VOUT.n5 Transmission_Gate_Layout_9.VOUT.t45 1.3109
R7092 Transmission_Gate_Layout_9.VOUT.n5 Transmission_Gate_Layout_9.VOUT.n4 1.3109
R7093 Transmission_Gate_Layout_9.VOUT.n95 Transmission_Gate_Layout_9.VOUT.t94 1.3109
R7094 Transmission_Gate_Layout_9.VOUT.n95 Transmission_Gate_Layout_9.VOUT.n94 1.3109
R7095 Transmission_Gate_Layout_9.VOUT.n92 Transmission_Gate_Layout_9.VOUT.t91 1.3109
R7096 Transmission_Gate_Layout_9.VOUT.n92 Transmission_Gate_Layout_9.VOUT.n91 1.3109
R7097 Transmission_Gate_Layout_9.VOUT.n90 Transmission_Gate_Layout_9.VOUT.t100 1.3109
R7098 Transmission_Gate_Layout_9.VOUT.n90 Transmission_Gate_Layout_9.VOUT.n89 1.3109
R7099 Transmission_Gate_Layout_9.VOUT.n103 Transmission_Gate_Layout_9.VOUT.t97 1.3109
R7100 Transmission_Gate_Layout_9.VOUT.n103 Transmission_Gate_Layout_9.VOUT.n102 1.3109
R7101 Transmission_Gate_Layout_9.VOUT.n100 Transmission_Gate_Layout_9.VOUT.t98 1.3109
R7102 Transmission_Gate_Layout_9.VOUT.n100 Transmission_Gate_Layout_9.VOUT.n99 1.3109
R7103 Transmission_Gate_Layout_9.VOUT.n98 Transmission_Gate_Layout_9.VOUT.t96 1.3109
R7104 Transmission_Gate_Layout_9.VOUT.n98 Transmission_Gate_Layout_9.VOUT.n97 1.3109
R7105 Transmission_Gate_Layout_9.VOUT.n106 Transmission_Gate_Layout_9.VOUT.t99 1.3109
R7106 Transmission_Gate_Layout_9.VOUT.n106 Transmission_Gate_Layout_9.VOUT.n105 1.3109
R7107 Transmission_Gate_Layout_9.VOUT.n108 Transmission_Gate_Layout_9.VOUT.t90 1.3109
R7108 Transmission_Gate_Layout_9.VOUT.n108 Transmission_Gate_Layout_9.VOUT.n107 1.3109
R7109 Transmission_Gate_Layout_9.VOUT.n110 Transmission_Gate_Layout_9.VOUT.t93 1.3109
R7110 Transmission_Gate_Layout_9.VOUT.n110 Transmission_Gate_Layout_9.VOUT.n109 1.3109
R7111 Transmission_Gate_Layout_9.VOUT.n166 Transmission_Gate_Layout_9.VOUT.t10 1.3109
R7112 Transmission_Gate_Layout_9.VOUT.n166 Transmission_Gate_Layout_9.VOUT.n165 1.3109
R7113 Transmission_Gate_Layout_9.VOUT.n163 Transmission_Gate_Layout_9.VOUT.t16 1.3109
R7114 Transmission_Gate_Layout_9.VOUT.n163 Transmission_Gate_Layout_9.VOUT.n162 1.3109
R7115 Transmission_Gate_Layout_9.VOUT.n161 Transmission_Gate_Layout_9.VOUT.t13 1.3109
R7116 Transmission_Gate_Layout_9.VOUT.n161 Transmission_Gate_Layout_9.VOUT.n160 1.3109
R7117 Transmission_Gate_Layout_9.VOUT.n177 Transmission_Gate_Layout_9.VOUT.t14 1.3109
R7118 Transmission_Gate_Layout_9.VOUT.n177 Transmission_Gate_Layout_9.VOUT.n176 1.3109
R7119 Transmission_Gate_Layout_9.VOUT.n179 Transmission_Gate_Layout_9.VOUT.t17 1.3109
R7120 Transmission_Gate_Layout_9.VOUT.n179 Transmission_Gate_Layout_9.VOUT.n178 1.3109
R7121 Transmission_Gate_Layout_9.VOUT.n181 Transmission_Gate_Layout_9.VOUT.t11 1.3109
R7122 Transmission_Gate_Layout_9.VOUT.n181 Transmission_Gate_Layout_9.VOUT.n180 1.3109
R7123 Transmission_Gate_Layout_9.VOUT.n174 Transmission_Gate_Layout_9.VOUT.t19 1.3109
R7124 Transmission_Gate_Layout_9.VOUT.n174 Transmission_Gate_Layout_9.VOUT.n173 1.3109
R7125 Transmission_Gate_Layout_9.VOUT.n171 Transmission_Gate_Layout_9.VOUT.t20 1.3109
R7126 Transmission_Gate_Layout_9.VOUT.n171 Transmission_Gate_Layout_9.VOUT.n170 1.3109
R7127 Transmission_Gate_Layout_9.VOUT.n169 Transmission_Gate_Layout_9.VOUT.t18 1.3109
R7128 Transmission_Gate_Layout_9.VOUT.n169 Transmission_Gate_Layout_9.VOUT.n168 1.3109
R7129 Transmission_Gate_Layout_9.VOUT.n35 Transmission_Gate_Layout_9.VOUT.t80 1.3109
R7130 Transmission_Gate_Layout_9.VOUT.n35 Transmission_Gate_Layout_9.VOUT.n34 1.3109
R7131 Transmission_Gate_Layout_9.VOUT.n37 Transmission_Gate_Layout_9.VOUT.t41 1.3109
R7132 Transmission_Gate_Layout_9.VOUT.n37 Transmission_Gate_Layout_9.VOUT.n36 1.3109
R7133 Transmission_Gate_Layout_9.VOUT.n39 Transmission_Gate_Layout_9.VOUT.t47 1.3109
R7134 Transmission_Gate_Layout_9.VOUT.n39 Transmission_Gate_Layout_9.VOUT.n38 1.3109
R7135 Transmission_Gate_Layout_9.VOUT.n54 Transmission_Gate_Layout_9.VOUT.t44 1.3109
R7136 Transmission_Gate_Layout_9.VOUT.n54 Transmission_Gate_Layout_9.VOUT.n53 1.3109
R7137 Transmission_Gate_Layout_9.VOUT.n51 Transmission_Gate_Layout_9.VOUT.t143 1.3109
R7138 Transmission_Gate_Layout_9.VOUT.n51 Transmission_Gate_Layout_9.VOUT.n50 1.3109
R7139 Transmission_Gate_Layout_9.VOUT.n49 Transmission_Gate_Layout_9.VOUT.t36 1.3109
R7140 Transmission_Gate_Layout_9.VOUT.n49 Transmission_Gate_Layout_9.VOUT.n48 1.3109
R7141 Transmission_Gate_Layout_9.VOUT.n46 Transmission_Gate_Layout_9.VOUT.t38 1.3109
R7142 Transmission_Gate_Layout_9.VOUT.n46 Transmission_Gate_Layout_9.VOUT.n45 1.3109
R7143 Transmission_Gate_Layout_9.VOUT.n43 Transmission_Gate_Layout_9.VOUT.t79 1.3109
R7144 Transmission_Gate_Layout_9.VOUT.n43 Transmission_Gate_Layout_9.VOUT.n42 1.3109
R7145 Transmission_Gate_Layout_9.VOUT.n41 Transmission_Gate_Layout_9.VOUT.t141 1.3109
R7146 Transmission_Gate_Layout_9.VOUT.n41 Transmission_Gate_Layout_9.VOUT.n40 1.3109
R7147 Transmission_Gate_Layout_9.VOUT.n131 Transmission_Gate_Layout_9.VOUT.n130 1.24485
R7148 Transmission_Gate_Layout_9.VOUT.n88 Transmission_Gate_Layout_9.VOUT.n87 1.24485
R7149 Transmission_Gate_Layout_9.VOUT.n135 Transmission_Gate_Layout_9.VOUT.n134 1.24485
R7150 Transmission_Gate_Layout_9.VOUT.n136 Transmission_Gate_Layout_9.VOUT.n135 1.24485
R7151 Transmission_Gate_Layout_9.VOUT.n80 Transmission_Gate_Layout_9.VOUT.n77 1.24485
R7152 Transmission_Gate_Layout_9.VOUT.n140 Transmission_Gate_Layout_9.VOUT.n139 1.24485
R7153 Transmission_Gate_Layout_9.VOUT.n139 Transmission_Gate_Layout_9.VOUT.n138 1.24485
R7154 Transmission_Gate_Layout_9.VOUT.n142 Transmission_Gate_Layout_9.VOUT.n141 1.24485
R7155 Transmission_Gate_Layout_9.VOUT.n143 Transmission_Gate_Layout_9.VOUT.n142 1.24485
R7156 Transmission_Gate_Layout_9.VOUT.n202 Transmission_Gate_Layout_9.VOUT.n201 1.24485
R7157 Transmission_Gate_Layout_9.VOUT.n159 Transmission_Gate_Layout_9.VOUT.n158 1.24485
R7158 Transmission_Gate_Layout_9.VOUT.n208 Transmission_Gate_Layout_9.VOUT.n206 1.24485
R7159 Transmission_Gate_Layout_9.VOUT.n210 Transmission_Gate_Layout_9.VOUT.n208 1.24485
R7160 Transmission_Gate_Layout_9.VOUT.n151 Transmission_Gate_Layout_9.VOUT.n148 1.24485
R7161 Transmission_Gate_Layout_9.VOUT.n15 Transmission_Gate_Layout_9.VOUT.n14 1.24485
R7162 Transmission_Gate_Layout_9.VOUT.n23 Transmission_Gate_Layout_9.VOUT.n22 1.24485
R7163 Transmission_Gate_Layout_9.VOUT.n30 Transmission_Gate_Layout_9.VOUT.n27 1.24485
R7164 Transmission_Gate_Layout_9.VOUT.n33 Transmission_Gate_Layout_9.VOUT.n30 1.24485
R7165 Transmission_Gate_Layout_9.VOUT.n68 Transmission_Gate_Layout_9.VOUT.n65 1.24485
R7166 Transmission_Gate_Layout_9.VOUT.n134 Transmission_Gate_Layout_9.VOUT.n133 1.2018
R7167 Transmission_Gate_Layout_9.VOUT.n138 Transmission_Gate_Layout_9.VOUT.n137 1.2018
R7168 Transmission_Gate_Layout_9.VOUT.n206 Transmission_Gate_Layout_9.VOUT.n204 1.2018
R7169 Transmission_Gate_Layout_9.VOUT.n24 Transmission_Gate_Layout_9.VOUT.n23 1.2018
R7170 Transmission_Gate_Layout_9.VOUT.n27 Transmission_Gate_Layout_9.VOUT.n24 1.2018
R7171 Transmission_Gate_Layout_9.VOUT.n118 Transmission_Gate_Layout_9.VOUT.n117 0.957239
R7172 Transmission_Gate_Layout_9.VOUT.n122 Transmission_Gate_Layout_9.VOUT.n121 0.957239
R7173 Transmission_Gate_Layout_9.VOUT.n186 Transmission_Gate_Layout_9.VOUT.n185 0.957239
R7174 Transmission_Gate_Layout_9.VOUT.n193 Transmission_Gate_Layout_9.VOUT.n192 0.957239
R7175 Transmission_Gate_Layout_9.VOUT.n56 Transmission_Gate_Layout_9.VOUT.n55 0.957239
R7176 Transmission_Gate_Layout_9.VOUT.n57 Transmission_Gate_Layout_9.VOUT.n56 0.957239
R7177 Transmission_Gate_Layout_9.VOUT.n60 Transmission_Gate_Layout_9.VOUT.n33 0.806587
R7178 Transmission_Gate_Layout_9.VOUT.n69 Transmission_Gate_Layout_9.VOUT.n68 0.806587
R7179 Transmission_Gate_Layout_9.VOUT.n7 Transmission_Gate_Layout_9.VOUT.n6 0.755717
R7180 Transmission_Gate_Layout_9.VOUT.n96 Transmission_Gate_Layout_9.VOUT.n93 0.755717
R7181 Transmission_Gate_Layout_9.VOUT.n104 Transmission_Gate_Layout_9.VOUT.n101 0.755717
R7182 Transmission_Gate_Layout_9.VOUT.n112 Transmission_Gate_Layout_9.VOUT.n111 0.755717
R7183 Transmission_Gate_Layout_9.VOUT.n117 Transmission_Gate_Layout_9.VOUT.n116 0.755717
R7184 Transmission_Gate_Layout_9.VOUT.n120 Transmission_Gate_Layout_9.VOUT.n119 0.755717
R7185 Transmission_Gate_Layout_9.VOUT.n121 Transmission_Gate_Layout_9.VOUT.n120 0.755717
R7186 Transmission_Gate_Layout_9.VOUT.n167 Transmission_Gate_Layout_9.VOUT.n164 0.755717
R7187 Transmission_Gate_Layout_9.VOUT.n183 Transmission_Gate_Layout_9.VOUT.n182 0.755717
R7188 Transmission_Gate_Layout_9.VOUT.n185 Transmission_Gate_Layout_9.VOUT.n184 0.755717
R7189 Transmission_Gate_Layout_9.VOUT.n190 Transmission_Gate_Layout_9.VOUT.n188 0.755717
R7190 Transmission_Gate_Layout_9.VOUT.n192 Transmission_Gate_Layout_9.VOUT.n190 0.755717
R7191 Transmission_Gate_Layout_9.VOUT.n175 Transmission_Gate_Layout_9.VOUT.n172 0.755717
R7192 Transmission_Gate_Layout_9.VOUT.n55 Transmission_Gate_Layout_9.VOUT.n52 0.755717
R7193 Transmission_Gate_Layout_9.VOUT.n47 Transmission_Gate_Layout_9.VOUT.n44 0.755717
R7194 Transmission_Gate_Layout_9.VOUT.n59 Transmission_Gate_Layout_9.VOUT.n58 0.755717
R7195 Transmission_Gate_Layout_9.VOUT.n58 Transmission_Gate_Layout_9.VOUT.n57 0.755717
R7196 Transmission_Gate_Layout_9.VOUT.n67 Transmission_Gate_Layout_9.VOUT.t139 0.7285
R7197 Transmission_Gate_Layout_9.VOUT.n67 Transmission_Gate_Layout_9.VOUT.n66 0.7285
R7198 Transmission_Gate_Layout_9.VOUT.n62 Transmission_Gate_Layout_9.VOUT.t130 0.7285
R7199 Transmission_Gate_Layout_9.VOUT.n62 Transmission_Gate_Layout_9.VOUT.n61 0.7285
R7200 Transmission_Gate_Layout_9.VOUT.n125 Transmission_Gate_Layout_9.VOUT.t73 0.7285
R7201 Transmission_Gate_Layout_9.VOUT.n125 Transmission_Gate_Layout_9.VOUT.n124 0.7285
R7202 Transmission_Gate_Layout_9.VOUT.n127 Transmission_Gate_Layout_9.VOUT.t110 0.7285
R7203 Transmission_Gate_Layout_9.VOUT.n127 Transmission_Gate_Layout_9.VOUT.n126 0.7285
R7204 Transmission_Gate_Layout_9.VOUT.n129 Transmission_Gate_Layout_9.VOUT.t2 0.7285
R7205 Transmission_Gate_Layout_9.VOUT.n129 Transmission_Gate_Layout_9.VOUT.n128 0.7285
R7206 Transmission_Gate_Layout_9.VOUT.n82 Transmission_Gate_Layout_9.VOUT.t3 0.7285
R7207 Transmission_Gate_Layout_9.VOUT.n82 Transmission_Gate_Layout_9.VOUT.n81 0.7285
R7208 Transmission_Gate_Layout_9.VOUT.n84 Transmission_Gate_Layout_9.VOUT.t74 0.7285
R7209 Transmission_Gate_Layout_9.VOUT.n84 Transmission_Gate_Layout_9.VOUT.n83 0.7285
R7210 Transmission_Gate_Layout_9.VOUT.n86 Transmission_Gate_Layout_9.VOUT.t112 0.7285
R7211 Transmission_Gate_Layout_9.VOUT.n86 Transmission_Gate_Layout_9.VOUT.n85 0.7285
R7212 Transmission_Gate_Layout_9.VOUT.n79 Transmission_Gate_Layout_9.VOUT.t4 0.7285
R7213 Transmission_Gate_Layout_9.VOUT.n79 Transmission_Gate_Layout_9.VOUT.n78 0.7285
R7214 Transmission_Gate_Layout_9.VOUT.n76 Transmission_Gate_Layout_9.VOUT.t111 0.7285
R7215 Transmission_Gate_Layout_9.VOUT.n76 Transmission_Gate_Layout_9.VOUT.n75 0.7285
R7216 Transmission_Gate_Layout_9.VOUT.n74 Transmission_Gate_Layout_9.VOUT.t76 0.7285
R7217 Transmission_Gate_Layout_9.VOUT.n74 Transmission_Gate_Layout_9.VOUT.n73 0.7285
R7218 Transmission_Gate_Layout_9.VOUT.n196 Transmission_Gate_Layout_9.VOUT.t61 0.7285
R7219 Transmission_Gate_Layout_9.VOUT.n196 Transmission_Gate_Layout_9.VOUT.n195 0.7285
R7220 Transmission_Gate_Layout_9.VOUT.n198 Transmission_Gate_Layout_9.VOUT.t68 0.7285
R7221 Transmission_Gate_Layout_9.VOUT.n198 Transmission_Gate_Layout_9.VOUT.n197 0.7285
R7222 Transmission_Gate_Layout_9.VOUT.n200 Transmission_Gate_Layout_9.VOUT.t53 0.7285
R7223 Transmission_Gate_Layout_9.VOUT.n200 Transmission_Gate_Layout_9.VOUT.n199 0.7285
R7224 Transmission_Gate_Layout_9.VOUT.n153 Transmission_Gate_Layout_9.VOUT.t67 0.7285
R7225 Transmission_Gate_Layout_9.VOUT.n153 Transmission_Gate_Layout_9.VOUT.n152 0.7285
R7226 Transmission_Gate_Layout_9.VOUT.n155 Transmission_Gate_Layout_9.VOUT.t49 0.7285
R7227 Transmission_Gate_Layout_9.VOUT.n155 Transmission_Gate_Layout_9.VOUT.n154 0.7285
R7228 Transmission_Gate_Layout_9.VOUT.n157 Transmission_Gate_Layout_9.VOUT.t59 0.7285
R7229 Transmission_Gate_Layout_9.VOUT.n157 Transmission_Gate_Layout_9.VOUT.n156 0.7285
R7230 Transmission_Gate_Layout_9.VOUT.n150 Transmission_Gate_Layout_9.VOUT.t50 0.7285
R7231 Transmission_Gate_Layout_9.VOUT.n150 Transmission_Gate_Layout_9.VOUT.n149 0.7285
R7232 Transmission_Gate_Layout_9.VOUT.n147 Transmission_Gate_Layout_9.VOUT.t65 0.7285
R7233 Transmission_Gate_Layout_9.VOUT.n147 Transmission_Gate_Layout_9.VOUT.n146 0.7285
R7234 Transmission_Gate_Layout_9.VOUT.n145 Transmission_Gate_Layout_9.VOUT.t58 0.7285
R7235 Transmission_Gate_Layout_9.VOUT.n145 Transmission_Gate_Layout_9.VOUT.n144 0.7285
R7236 Transmission_Gate_Layout_9.VOUT.n32 Transmission_Gate_Layout_9.VOUT.t127 0.7285
R7237 Transmission_Gate_Layout_9.VOUT.n32 Transmission_Gate_Layout_9.VOUT.n31 0.7285
R7238 Transmission_Gate_Layout_9.VOUT.n29 Transmission_Gate_Layout_9.VOUT.t120 0.7285
R7239 Transmission_Gate_Layout_9.VOUT.n29 Transmission_Gate_Layout_9.VOUT.n28 0.7285
R7240 Transmission_Gate_Layout_9.VOUT.n26 Transmission_Gate_Layout_9.VOUT.t121 0.7285
R7241 Transmission_Gate_Layout_9.VOUT.n26 Transmission_Gate_Layout_9.VOUT.n25 0.7285
R7242 Transmission_Gate_Layout_9.VOUT.n9 Transmission_Gate_Layout_9.VOUT.t138 0.7285
R7243 Transmission_Gate_Layout_9.VOUT.n9 Transmission_Gate_Layout_9.VOUT.n8 0.7285
R7244 Transmission_Gate_Layout_9.VOUT.n11 Transmission_Gate_Layout_9.VOUT.t137 0.7285
R7245 Transmission_Gate_Layout_9.VOUT.n11 Transmission_Gate_Layout_9.VOUT.n10 0.7285
R7246 Transmission_Gate_Layout_9.VOUT.n13 Transmission_Gate_Layout_9.VOUT.t123 0.7285
R7247 Transmission_Gate_Layout_9.VOUT.n13 Transmission_Gate_Layout_9.VOUT.n12 0.7285
R7248 Transmission_Gate_Layout_9.VOUT.n17 Transmission_Gate_Layout_9.VOUT.t132 0.7285
R7249 Transmission_Gate_Layout_9.VOUT.n17 Transmission_Gate_Layout_9.VOUT.n16 0.7285
R7250 Transmission_Gate_Layout_9.VOUT.n19 Transmission_Gate_Layout_9.VOUT.t129 0.7285
R7251 Transmission_Gate_Layout_9.VOUT.n19 Transmission_Gate_Layout_9.VOUT.n18 0.7285
R7252 Transmission_Gate_Layout_9.VOUT.n21 Transmission_Gate_Layout_9.VOUT.t117 0.7285
R7253 Transmission_Gate_Layout_9.VOUT.n21 Transmission_Gate_Layout_9.VOUT.n20 0.7285
R7254 Transmission_Gate_Layout_9.VOUT.n64 Transmission_Gate_Layout_9.VOUT.t128 0.7285
R7255 Transmission_Gate_Layout_9.VOUT.n64 Transmission_Gate_Layout_9.VOUT.n63 0.7285
R7256 Transmission_Gate_Layout_9.VOUT.n123 Transmission_Gate_Layout_9.VOUT.n122 0.626587
R7257 Transmission_Gate_Layout_9.VOUT.n133 Transmission_Gate_Layout_9.VOUT.n132 0.626587
R7258 Transmission_Gate_Layout_9.VOUT.n194 Transmission_Gate_Layout_9.VOUT.n193 0.626587
R7259 Transmission_Gate_Layout_9.VOUT.n204 Transmission_Gate_Layout_9.VOUT.n203 0.626587
R7260 Transmission_Gate_Layout_9.VOUT.n69 Transmission_Gate_Layout_9.VOUT.n60 0.626587
R7261 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.VOUT.n140 0.607022
R7262 Transmission_Gate_Layout_9.VOUT.n141 Transmission_Gate_Layout_9.VOUT 0.607022
R7263 Transmission_Gate_Layout_9.VOUT.n212 Transmission_Gate_Layout_9.VOUT.n211 0.597239
R7264 Transmission_Gate_Layout_9.VOUT.n132 Transmission_Gate_Layout_9.VOUT.n131 0.575717
R7265 Transmission_Gate_Layout_9.VOUT.n133 Transmission_Gate_Layout_9.VOUT.n88 0.575717
R7266 Transmission_Gate_Layout_9.VOUT.n137 Transmission_Gate_Layout_9.VOUT.n80 0.575717
R7267 Transmission_Gate_Layout_9.VOUT.n203 Transmission_Gate_Layout_9.VOUT.n202 0.575717
R7268 Transmission_Gate_Layout_9.VOUT.n204 Transmission_Gate_Layout_9.VOUT.n159 0.575717
R7269 Transmission_Gate_Layout_9.VOUT.n211 Transmission_Gate_Layout_9.VOUT.n151 0.575717
R7270 Transmission_Gate_Layout_9.VOUT.n24 Transmission_Gate_Layout_9.VOUT.n15 0.575717
R7271 Transmission_Gate_Layout_9.VOUT.n212 Transmission_Gate_Layout_9.VOUT.n143 0.54637
R7272 Transmission_Gate_Layout_9.VOUT.n69 Transmission_Gate_Layout_9.VOUT.n7 0.428978
R7273 Transmission_Gate_Layout_9.VOUT.n60 Transmission_Gate_Layout_9.VOUT.n59 0.428978
R7274 Transmission_Gate_Layout_9.VOUT.n123 Transmission_Gate_Layout_9.VOUT.n96 0.331152
R7275 Transmission_Gate_Layout_9.VOUT.n122 Transmission_Gate_Layout_9.VOUT.n104 0.331152
R7276 Transmission_Gate_Layout_9.VOUT.n118 Transmission_Gate_Layout_9.VOUT.n112 0.331152
R7277 Transmission_Gate_Layout_9.VOUT.n194 Transmission_Gate_Layout_9.VOUT.n167 0.331152
R7278 Transmission_Gate_Layout_9.VOUT.n186 Transmission_Gate_Layout_9.VOUT.n183 0.331152
R7279 Transmission_Gate_Layout_9.VOUT.n193 Transmission_Gate_Layout_9.VOUT.n175 0.331152
R7280 Transmission_Gate_Layout_9.VOUT.n56 Transmission_Gate_Layout_9.VOUT.n47 0.331152
R7281 Transmission_Gate_Layout_9.VOUT.n132 Transmission_Gate_Layout_9.VOUT.n123 0.239196
R7282 Transmission_Gate_Layout_9.VOUT.n203 Transmission_Gate_Layout_9.VOUT.n194 0.239196
R7283 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_9.VOUT.n69 0.192239
R7284 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.t5 17.8546
R7285 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n0 14.0337
R7286 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.t4 13.5862
R7287 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n2 3.76289
R7288 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n2 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.t3 3.2765
R7289 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n2 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n1 3.2765
R7290 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n4 2.88224
R7291 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n4 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.t2 1.8205
R7292 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n4 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT.n3 1.8205
R7293 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT.t3 17.8546
R7294 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT.n0 14.0337
R7295 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT.t2 13.5862
R7296 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT.n1 9.5898
R7297 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_1.OUT.n2 7.76208
R7298 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT.t3 17.8546
R7299 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT.n0 14.0337
R7300 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT.t2 13.5862
R7301 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT.n1 9.5898
R7302 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_1.OUT.n2 7.76208
R7303 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT.t3 17.8546
R7304 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT.n0 14.0337
R7305 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT.t2 13.5862
R7306 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT.n1 9.5898
R7307 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_2.OUT.n2 7.76208
R7308 Transmission_Gate_Layout_11.CLKB.n27 Transmission_Gate_Layout_11.CLKB.t19 54.5477
R7309 Transmission_Gate_Layout_11.CLKB.n27 Transmission_Gate_Layout_11.CLKB.t25 38.3255
R7310 Transmission_Gate_Layout_11.CLKB.n28 Transmission_Gate_Layout_11.CLKB.t12 38.3255
R7311 Transmission_Gate_Layout_11.CLKB.n29 Transmission_Gate_Layout_11.CLKB.t23 38.3255
R7312 Transmission_Gate_Layout_11.CLKB.n30 Transmission_Gate_Layout_11.CLKB.t11 38.3255
R7313 Transmission_Gate_Layout_11.CLKB.n31 Transmission_Gate_Layout_11.CLKB.t17 38.3255
R7314 Transmission_Gate_Layout_11.CLKB.n32 Transmission_Gate_Layout_11.CLKB.t22 38.3255
R7315 Transmission_Gate_Layout_11.CLKB.t21 Transmission_Gate_Layout_11.CLKB.n24 37.9344
R7316 Transmission_Gate_Layout_11.CLKB.t26 Transmission_Gate_Layout_11.CLKB.n23 37.9344
R7317 Transmission_Gate_Layout_11.CLKB.t8 Transmission_Gate_Layout_11.CLKB.n20 37.9344
R7318 Transmission_Gate_Layout_11.CLKB.t20 Transmission_Gate_Layout_11.CLKB.n17 37.9344
R7319 Transmission_Gate_Layout_11.CLKB.t6 Transmission_Gate_Layout_11.CLKB.n14 37.9344
R7320 Transmission_Gate_Layout_11.CLKB.t18 Transmission_Gate_Layout_11.CLKB.n11 37.9344
R7321 Transmission_Gate_Layout_11.CLKB.t24 Transmission_Gate_Layout_11.CLKB.n8 37.9344
R7322 Transmission_Gate_Layout_11.CLKB.t28 Transmission_Gate_Layout_11.CLKB.n5 37.9344
R7323 Transmission_Gate_Layout_11.CLKB.n25 Transmission_Gate_Layout_11.CLKB.t21 37.5434
R7324 Transmission_Gate_Layout_11.CLKB.n26 Transmission_Gate_Layout_11.CLKB.t26 37.5434
R7325 Transmission_Gate_Layout_11.CLKB.n21 Transmission_Gate_Layout_11.CLKB.t8 37.5434
R7326 Transmission_Gate_Layout_11.CLKB.n18 Transmission_Gate_Layout_11.CLKB.t20 37.5434
R7327 Transmission_Gate_Layout_11.CLKB.n15 Transmission_Gate_Layout_11.CLKB.t6 37.5434
R7328 Transmission_Gate_Layout_11.CLKB.n12 Transmission_Gate_Layout_11.CLKB.t18 37.5434
R7329 Transmission_Gate_Layout_11.CLKB.n9 Transmission_Gate_Layout_11.CLKB.t24 37.5434
R7330 Transmission_Gate_Layout_11.CLKB.n6 Transmission_Gate_Layout_11.CLKB.t28 37.5434
R7331 Transmission_Gate_Layout_11.CLKB.n25 Transmission_Gate_Layout_11.CLKB.t14 37.413
R7332 Transmission_Gate_Layout_11.CLKB.t25 Transmission_Gate_Layout_11.CLKB.n21 37.413
R7333 Transmission_Gate_Layout_11.CLKB.t12 Transmission_Gate_Layout_11.CLKB.n18 37.413
R7334 Transmission_Gate_Layout_11.CLKB.t23 Transmission_Gate_Layout_11.CLKB.n15 37.413
R7335 Transmission_Gate_Layout_11.CLKB.t11 Transmission_Gate_Layout_11.CLKB.n12 37.413
R7336 Transmission_Gate_Layout_11.CLKB.t17 Transmission_Gate_Layout_11.CLKB.n9 37.413
R7337 Transmission_Gate_Layout_11.CLKB.t22 Transmission_Gate_Layout_11.CLKB.n6 37.413
R7338 Transmission_Gate_Layout_11.CLKB.t19 Transmission_Gate_Layout_11.CLKB.n26 37.413
R7339 Transmission_Gate_Layout_11.CLKB.n24 Transmission_Gate_Layout_11.CLKB.t7 37.0219
R7340 Transmission_Gate_Layout_11.CLKB.n23 Transmission_Gate_Layout_11.CLKB.t10 37.0219
R7341 Transmission_Gate_Layout_11.CLKB.n20 Transmission_Gate_Layout_11.CLKB.t16 37.0219
R7342 Transmission_Gate_Layout_11.CLKB.n17 Transmission_Gate_Layout_11.CLKB.t29 37.0219
R7343 Transmission_Gate_Layout_11.CLKB.n14 Transmission_Gate_Layout_11.CLKB.t15 37.0219
R7344 Transmission_Gate_Layout_11.CLKB.n11 Transmission_Gate_Layout_11.CLKB.t27 37.0219
R7345 Transmission_Gate_Layout_11.CLKB.n5 Transmission_Gate_Layout_11.CLKB.t13 37.0219
R7346 Transmission_Gate_Layout_11.CLKB.n8 Transmission_Gate_Layout_11.CLKB.t9 37.0219
R7347 Transmission_Gate_Layout_11.CLKB.t10 Transmission_Gate_Layout_11.CLKB.n22 35.1969
R7348 Transmission_Gate_Layout_11.CLKB.t16 Transmission_Gate_Layout_11.CLKB.n19 35.1969
R7349 Transmission_Gate_Layout_11.CLKB.t29 Transmission_Gate_Layout_11.CLKB.n16 35.1969
R7350 Transmission_Gate_Layout_11.CLKB.t15 Transmission_Gate_Layout_11.CLKB.n13 35.1969
R7351 Transmission_Gate_Layout_11.CLKB.t27 Transmission_Gate_Layout_11.CLKB.n10 35.1969
R7352 Transmission_Gate_Layout_11.CLKB.t9 Transmission_Gate_Layout_11.CLKB.n7 35.1969
R7353 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLKB.n32 26.6826
R7354 Transmission_Gate_Layout_11.CLKB.n26 Transmission_Gate_Layout_11.CLKB.n25 19.148
R7355 Transmission_Gate_Layout_11.CLKB.n28 Transmission_Gate_Layout_11.CLKB.n27 16.2227
R7356 Transmission_Gate_Layout_11.CLKB.n29 Transmission_Gate_Layout_11.CLKB.n28 16.2227
R7357 Transmission_Gate_Layout_11.CLKB.n30 Transmission_Gate_Layout_11.CLKB.n29 16.2227
R7358 Transmission_Gate_Layout_11.CLKB.n31 Transmission_Gate_Layout_11.CLKB.n30 16.2227
R7359 Transmission_Gate_Layout_11.CLKB.n32 Transmission_Gate_Layout_11.CLKB.n31 16.2227
R7360 Transmission_Gate_Layout_11.CLKB.n2 Transmission_Gate_Layout_11.CLKB.n0 5.21612
R7361 Transmission_Gate_Layout_11.CLKB.n35 Transmission_Gate_Layout_11.CLKB.n34 4.57285
R7362 Transmission_Gate_Layout_11.CLKB.n2 Transmission_Gate_Layout_11.CLKB.n1 4.4609
R7363 Transmission_Gate_Layout_11.CLKB.n4 Transmission_Gate_Layout_11.CLKB.n3 4.4609
R7364 Transmission_Gate_Layout_11.CLKB.n35 Transmission_Gate_Layout_11.CLKB.n33 3.3285
R7365 Transmission_Gate_Layout_11.CLKB.n37 Transmission_Gate_Layout_11.CLKB.n36 3.3285
R7366 Transmission_Gate_Layout_11.CLKB.n37 Transmission_Gate_Layout_11.CLKB.n35 1.24485
R7367 Transmission_Gate_Layout_11.CLKB.n4 Transmission_Gate_Layout_11.CLKB.n2 0.755717
R7368 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLKB.n37 0.750969
R7369 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_11.CLKB.n4 0.510317
R7370 Transmission_Gate_Layout_11.VIN.n104 Transmission_Gate_Layout_11.VIN.n95 32.6807
R7371 Transmission_Gate_Layout_11.VIN.n27 Transmission_Gate_Layout_11.VIN.n26 5.21612
R7372 Transmission_Gate_Layout_11.VIN.n28 Transmission_Gate_Layout_11.VIN.n24 4.4609
R7373 Transmission_Gate_Layout_11.VIN.n27 Transmission_Gate_Layout_11.VIN.n25 4.4609
R7374 Transmission_Gate_Layout_11.VIN.n85 Transmission_Gate_Layout_11.VIN.t82 4.4609
R7375 Transmission_Gate_Layout_11.VIN.n84 Transmission_Gate_Layout_11.VIN.t79 4.4609
R7376 Transmission_Gate_Layout_11.VIN.n83 Transmission_Gate_Layout_11.VIN.t76 4.4609
R7377 Transmission_Gate_Layout_11.VIN.n41 Transmission_Gate_Layout_11.VIN.n38 3.90572
R7378 Transmission_Gate_Layout_11.VIN.n33 Transmission_Gate_Layout_11.VIN.n30 3.90572
R7379 Transmission_Gate_Layout_11.VIN.n92 Transmission_Gate_Layout_11.VIN.n91 3.90572
R7380 Transmission_Gate_Layout_11.VIN.n102 Transmission_Gate_Layout_11.VIN.n101 3.90572
R7381 Transmission_Gate_Layout_11.VIN.n22 Transmission_Gate_Layout_11.VIN.n21 3.90572
R7382 Transmission_Gate_Layout_11.VIN.n4 Transmission_Gate_Layout_11.VIN.n1 3.90572
R7383 Transmission_Gate_Layout_11.VIN.n51 Transmission_Gate_Layout_11.VIN.n50 3.84485
R7384 Transmission_Gate_Layout_11.VIN.n65 Transmission_Gate_Layout_11.VIN.n62 3.84485
R7385 Transmission_Gate_Layout_11.VIN.n59 Transmission_Gate_Layout_11.VIN.n58 3.84485
R7386 Transmission_Gate_Layout_11.VIN.n14 Transmission_Gate_Layout_11.VIN.n13 3.84485
R7387 Transmission_Gate_Layout_11.VIN.n125 Transmission_Gate_Layout_11.VIN.n122 3.84485
R7388 Transmission_Gate_Layout_11.VIN.n133 Transmission_Gate_Layout_11.VIN.n130 3.84485
R7389 Transmission_Gate_Layout_11.VIN.n78 Transmission_Gate_Layout_11.VIN.t61 3.3285
R7390 Transmission_Gate_Layout_11.VIN.n77 Transmission_Gate_Layout_11.VIN.t6 3.3285
R7391 Transmission_Gate_Layout_11.VIN.n76 Transmission_Gate_Layout_11.VIN.t67 3.3285
R7392 Transmission_Gate_Layout_11.VIN.n74 Transmission_Gate_Layout_11.VIN.n73 3.3285
R7393 Transmission_Gate_Layout_11.VIN.n72 Transmission_Gate_Layout_11.VIN.n71 3.3285
R7394 Transmission_Gate_Layout_11.VIN.n70 Transmission_Gate_Layout_11.VIN.n69 3.3285
R7395 Transmission_Gate_Layout_11.VIN.n41 Transmission_Gate_Layout_11.VIN.n40 3.1505
R7396 Transmission_Gate_Layout_11.VIN.n44 Transmission_Gate_Layout_11.VIN.n43 3.1505
R7397 Transmission_Gate_Layout_11.VIN.n33 Transmission_Gate_Layout_11.VIN.n32 3.1505
R7398 Transmission_Gate_Layout_11.VIN.n36 Transmission_Gate_Layout_11.VIN.n35 3.1505
R7399 Transmission_Gate_Layout_11.VIN.n92 Transmission_Gate_Layout_11.VIN.n89 3.1505
R7400 Transmission_Gate_Layout_11.VIN.n93 Transmission_Gate_Layout_11.VIN.n87 3.1505
R7401 Transmission_Gate_Layout_11.VIN.n102 Transmission_Gate_Layout_11.VIN.n99 3.1505
R7402 Transmission_Gate_Layout_11.VIN.n103 Transmission_Gate_Layout_11.VIN.n97 3.1505
R7403 Transmission_Gate_Layout_11.VIN.n22 Transmission_Gate_Layout_11.VIN.n19 3.1505
R7404 Transmission_Gate_Layout_11.VIN.n23 Transmission_Gate_Layout_11.VIN.n17 3.1505
R7405 Transmission_Gate_Layout_11.VIN.n114 Transmission_Gate_Layout_11.VIN.n113 3.1505
R7406 Transmission_Gate_Layout_11.VIN.n111 Transmission_Gate_Layout_11.VIN.n110 3.1505
R7407 Transmission_Gate_Layout_11.VIN.n108 Transmission_Gate_Layout_11.VIN.n107 3.1505
R7408 Transmission_Gate_Layout_11.VIN.n4 Transmission_Gate_Layout_11.VIN.n3 3.1505
R7409 Transmission_Gate_Layout_11.VIN.n7 Transmission_Gate_Layout_11.VIN.n6 3.1505
R7410 Transmission_Gate_Layout_11.VIN.n76 Transmission_Gate_Layout_11.VIN.n75 2.72398
R7411 Transmission_Gate_Layout_11.VIN.n51 Transmission_Gate_Layout_11.VIN.n48 2.6005
R7412 Transmission_Gate_Layout_11.VIN.n52 Transmission_Gate_Layout_11.VIN.n46 2.6005
R7413 Transmission_Gate_Layout_11.VIN.n65 Transmission_Gate_Layout_11.VIN.n64 2.6005
R7414 Transmission_Gate_Layout_11.VIN.n68 Transmission_Gate_Layout_11.VIN.n67 2.6005
R7415 Transmission_Gate_Layout_11.VIN.n59 Transmission_Gate_Layout_11.VIN.n56 2.6005
R7416 Transmission_Gate_Layout_11.VIN.n60 Transmission_Gate_Layout_11.VIN.n54 2.6005
R7417 Transmission_Gate_Layout_11.VIN.n14 Transmission_Gate_Layout_11.VIN.n11 2.6005
R7418 Transmission_Gate_Layout_11.VIN.n15 Transmission_Gate_Layout_11.VIN.n9 2.6005
R7419 Transmission_Gate_Layout_11.VIN.n138 Transmission_Gate_Layout_11.VIN.n120 2.6005
R7420 Transmission_Gate_Layout_11.VIN.n139 Transmission_Gate_Layout_11.VIN.n118 2.6005
R7421 Transmission_Gate_Layout_11.VIN.n140 Transmission_Gate_Layout_11.VIN.n116 2.6005
R7422 Transmission_Gate_Layout_11.VIN.n125 Transmission_Gate_Layout_11.VIN.n124 2.6005
R7423 Transmission_Gate_Layout_11.VIN.n128 Transmission_Gate_Layout_11.VIN.n127 2.6005
R7424 Transmission_Gate_Layout_11.VIN.n136 Transmission_Gate_Layout_11.VIN.n135 2.6005
R7425 Transmission_Gate_Layout_11.VIN.n133 Transmission_Gate_Layout_11.VIN.n132 2.6005
R7426 Transmission_Gate_Layout_11.VIN.n94 Transmission_Gate_Layout_11.VIN.n85 2.47941
R7427 Transmission_Gate_Layout_11.VIN.n107 Transmission_Gate_Layout_11.VIN.t51 1.3109
R7428 Transmission_Gate_Layout_11.VIN.n107 Transmission_Gate_Layout_11.VIN.n106 1.3109
R7429 Transmission_Gate_Layout_11.VIN.n110 Transmission_Gate_Layout_11.VIN.t57 1.3109
R7430 Transmission_Gate_Layout_11.VIN.n110 Transmission_Gate_Layout_11.VIN.n109 1.3109
R7431 Transmission_Gate_Layout_11.VIN.n113 Transmission_Gate_Layout_11.VIN.t53 1.3109
R7432 Transmission_Gate_Layout_11.VIN.n113 Transmission_Gate_Layout_11.VIN.n112 1.3109
R7433 Transmission_Gate_Layout_11.VIN.n87 Transmission_Gate_Layout_11.VIN.t77 1.3109
R7434 Transmission_Gate_Layout_11.VIN.n87 Transmission_Gate_Layout_11.VIN.n86 1.3109
R7435 Transmission_Gate_Layout_11.VIN.n89 Transmission_Gate_Layout_11.VIN.t74 1.3109
R7436 Transmission_Gate_Layout_11.VIN.n89 Transmission_Gate_Layout_11.VIN.n88 1.3109
R7437 Transmission_Gate_Layout_11.VIN.n91 Transmission_Gate_Layout_11.VIN.t84 1.3109
R7438 Transmission_Gate_Layout_11.VIN.n91 Transmission_Gate_Layout_11.VIN.n90 1.3109
R7439 Transmission_Gate_Layout_11.VIN.n43 Transmission_Gate_Layout_11.VIN.t80 1.3109
R7440 Transmission_Gate_Layout_11.VIN.n43 Transmission_Gate_Layout_11.VIN.n42 1.3109
R7441 Transmission_Gate_Layout_11.VIN.n40 Transmission_Gate_Layout_11.VIN.t83 1.3109
R7442 Transmission_Gate_Layout_11.VIN.n40 Transmission_Gate_Layout_11.VIN.n39 1.3109
R7443 Transmission_Gate_Layout_11.VIN.n38 Transmission_Gate_Layout_11.VIN.t73 1.3109
R7444 Transmission_Gate_Layout_11.VIN.n38 Transmission_Gate_Layout_11.VIN.n37 1.3109
R7445 Transmission_Gate_Layout_11.VIN.n35 Transmission_Gate_Layout_11.VIN.t75 1.3109
R7446 Transmission_Gate_Layout_11.VIN.n35 Transmission_Gate_Layout_11.VIN.n34 1.3109
R7447 Transmission_Gate_Layout_11.VIN.n32 Transmission_Gate_Layout_11.VIN.t78 1.3109
R7448 Transmission_Gate_Layout_11.VIN.n32 Transmission_Gate_Layout_11.VIN.n31 1.3109
R7449 Transmission_Gate_Layout_11.VIN.n30 Transmission_Gate_Layout_11.VIN.t81 1.3109
R7450 Transmission_Gate_Layout_11.VIN.n30 Transmission_Gate_Layout_11.VIN.n29 1.3109
R7451 Transmission_Gate_Layout_11.VIN.n97 Transmission_Gate_Layout_11.VIN.t60 1.3109
R7452 Transmission_Gate_Layout_11.VIN.n97 Transmission_Gate_Layout_11.VIN.n96 1.3109
R7453 Transmission_Gate_Layout_11.VIN.n99 Transmission_Gate_Layout_11.VIN.t42 1.3109
R7454 Transmission_Gate_Layout_11.VIN.n99 Transmission_Gate_Layout_11.VIN.n98 1.3109
R7455 Transmission_Gate_Layout_11.VIN.n101 Transmission_Gate_Layout_11.VIN.t38 1.3109
R7456 Transmission_Gate_Layout_11.VIN.n101 Transmission_Gate_Layout_11.VIN.n100 1.3109
R7457 Transmission_Gate_Layout_11.VIN.n17 Transmission_Gate_Layout_11.VIN.t45 1.3109
R7458 Transmission_Gate_Layout_11.VIN.n17 Transmission_Gate_Layout_11.VIN.n16 1.3109
R7459 Transmission_Gate_Layout_11.VIN.n19 Transmission_Gate_Layout_11.VIN.t49 1.3109
R7460 Transmission_Gate_Layout_11.VIN.n19 Transmission_Gate_Layout_11.VIN.n18 1.3109
R7461 Transmission_Gate_Layout_11.VIN.n21 Transmission_Gate_Layout_11.VIN.t54 1.3109
R7462 Transmission_Gate_Layout_11.VIN.n21 Transmission_Gate_Layout_11.VIN.n20 1.3109
R7463 Transmission_Gate_Layout_11.VIN.n6 Transmission_Gate_Layout_11.VIN.t39 1.3109
R7464 Transmission_Gate_Layout_11.VIN.n6 Transmission_Gate_Layout_11.VIN.n5 1.3109
R7465 Transmission_Gate_Layout_11.VIN.n3 Transmission_Gate_Layout_11.VIN.t47 1.3109
R7466 Transmission_Gate_Layout_11.VIN.n3 Transmission_Gate_Layout_11.VIN.n2 1.3109
R7467 Transmission_Gate_Layout_11.VIN.n1 Transmission_Gate_Layout_11.VIN.t41 1.3109
R7468 Transmission_Gate_Layout_11.VIN.n1 Transmission_Gate_Layout_11.VIN.n0 1.3109
R7469 Transmission_Gate_Layout_11.VIN.n52 Transmission_Gate_Layout_11.VIN.n51 1.24485
R7470 Transmission_Gate_Layout_11.VIN.n68 Transmission_Gate_Layout_11.VIN.n65 1.24485
R7471 Transmission_Gate_Layout_11.VIN.n72 Transmission_Gate_Layout_11.VIN.n70 1.24485
R7472 Transmission_Gate_Layout_11.VIN.n74 Transmission_Gate_Layout_11.VIN.n72 1.24485
R7473 Transmission_Gate_Layout_11.VIN.n78 Transmission_Gate_Layout_11.VIN.n77 1.24485
R7474 Transmission_Gate_Layout_11.VIN.n77 Transmission_Gate_Layout_11.VIN.n76 1.24485
R7475 Transmission_Gate_Layout_11.VIN.n60 Transmission_Gate_Layout_11.VIN.n59 1.24485
R7476 Transmission_Gate_Layout_11.VIN.n15 Transmission_Gate_Layout_11.VIN.n14 1.24485
R7477 Transmission_Gate_Layout_11.VIN.n140 Transmission_Gate_Layout_11.VIN.n139 1.24485
R7478 Transmission_Gate_Layout_11.VIN.n139 Transmission_Gate_Layout_11.VIN.n138 1.24485
R7479 Transmission_Gate_Layout_11.VIN.n128 Transmission_Gate_Layout_11.VIN.n125 1.24485
R7480 Transmission_Gate_Layout_11.VIN.n136 Transmission_Gate_Layout_11.VIN.n133 1.24485
R7481 Transmission_Gate_Layout_11.VIN.n75 Transmission_Gate_Layout_11.VIN.n74 1.2018
R7482 Transmission_Gate_Layout_11.VIN.n79 Transmission_Gate_Layout_11.VIN.n78 1.2018
R7483 Transmission_Gate_Layout_11.VIN.n138 Transmission_Gate_Layout_11.VIN.n137 1.2018
R7484 Transmission_Gate_Layout_11.VIN.n137 Transmission_Gate_Layout_11.VIN.n128 1.2018
R7485 Transmission_Gate_Layout_11.VIN.n83 Transmission_Gate_Layout_11.VIN.n82 0.957239
R7486 Transmission_Gate_Layout_11.VIN.n108 Transmission_Gate_Layout_11.VIN.n105 0.957239
R7487 Transmission_Gate_Layout_11.VIN.n142 Transmission_Gate_Layout_11.VIN.n15 0.806587
R7488 Transmission_Gate_Layout_11.VIN.n141 Transmission_Gate_Layout_11.VIN.n140 0.806587
R7489 Transmission_Gate_Layout_11.VIN.n28 Transmission_Gate_Layout_11.VIN.n27 0.755717
R7490 Transmission_Gate_Layout_11.VIN.n44 Transmission_Gate_Layout_11.VIN.n41 0.755717
R7491 Transmission_Gate_Layout_11.VIN.n36 Transmission_Gate_Layout_11.VIN.n33 0.755717
R7492 Transmission_Gate_Layout_11.VIN.n85 Transmission_Gate_Layout_11.VIN.n84 0.755717
R7493 Transmission_Gate_Layout_11.VIN.n84 Transmission_Gate_Layout_11.VIN.n83 0.755717
R7494 Transmission_Gate_Layout_11.VIN.n93 Transmission_Gate_Layout_11.VIN.n92 0.755717
R7495 Transmission_Gate_Layout_11.VIN.n103 Transmission_Gate_Layout_11.VIN.n102 0.755717
R7496 Transmission_Gate_Layout_11.VIN.n23 Transmission_Gate_Layout_11.VIN.n22 0.755717
R7497 Transmission_Gate_Layout_11.VIN.n111 Transmission_Gate_Layout_11.VIN.n108 0.755717
R7498 Transmission_Gate_Layout_11.VIN.n114 Transmission_Gate_Layout_11.VIN.n111 0.755717
R7499 Transmission_Gate_Layout_11.VIN.n7 Transmission_Gate_Layout_11.VIN.n4 0.755717
R7500 Transmission_Gate_Layout_11.VIN.n135 Transmission_Gate_Layout_11.VIN.t27 0.7285
R7501 Transmission_Gate_Layout_11.VIN.n135 Transmission_Gate_Layout_11.VIN.n134 0.7285
R7502 Transmission_Gate_Layout_11.VIN.n130 Transmission_Gate_Layout_11.VIN.t19 0.7285
R7503 Transmission_Gate_Layout_11.VIN.n130 Transmission_Gate_Layout_11.VIN.n129 0.7285
R7504 Transmission_Gate_Layout_11.VIN.n116 Transmission_Gate_Layout_11.VIN.t17 0.7285
R7505 Transmission_Gate_Layout_11.VIN.n116 Transmission_Gate_Layout_11.VIN.n115 0.7285
R7506 Transmission_Gate_Layout_11.VIN.n118 Transmission_Gate_Layout_11.VIN.t34 0.7285
R7507 Transmission_Gate_Layout_11.VIN.n118 Transmission_Gate_Layout_11.VIN.n117 0.7285
R7508 Transmission_Gate_Layout_11.VIN.n120 Transmission_Gate_Layout_11.VIN.t26 0.7285
R7509 Transmission_Gate_Layout_11.VIN.n120 Transmission_Gate_Layout_11.VIN.n119 0.7285
R7510 Transmission_Gate_Layout_11.VIN.n46 Transmission_Gate_Layout_11.VIN.t5 0.7285
R7511 Transmission_Gate_Layout_11.VIN.n46 Transmission_Gate_Layout_11.VIN.n45 0.7285
R7512 Transmission_Gate_Layout_11.VIN.n48 Transmission_Gate_Layout_11.VIN.t71 0.7285
R7513 Transmission_Gate_Layout_11.VIN.n48 Transmission_Gate_Layout_11.VIN.n47 0.7285
R7514 Transmission_Gate_Layout_11.VIN.n50 Transmission_Gate_Layout_11.VIN.t10 0.7285
R7515 Transmission_Gate_Layout_11.VIN.n50 Transmission_Gate_Layout_11.VIN.n49 0.7285
R7516 Transmission_Gate_Layout_11.VIN.n67 Transmission_Gate_Layout_11.VIN.t2 0.7285
R7517 Transmission_Gate_Layout_11.VIN.n67 Transmission_Gate_Layout_11.VIN.n66 0.7285
R7518 Transmission_Gate_Layout_11.VIN.n64 Transmission_Gate_Layout_11.VIN.t63 0.7285
R7519 Transmission_Gate_Layout_11.VIN.n64 Transmission_Gate_Layout_11.VIN.n63 0.7285
R7520 Transmission_Gate_Layout_11.VIN.n62 Transmission_Gate_Layout_11.VIN.t70 0.7285
R7521 Transmission_Gate_Layout_11.VIN.n62 Transmission_Gate_Layout_11.VIN.n61 0.7285
R7522 Transmission_Gate_Layout_11.VIN.n54 Transmission_Gate_Layout_11.VIN.t62 0.7285
R7523 Transmission_Gate_Layout_11.VIN.n54 Transmission_Gate_Layout_11.VIN.n53 0.7285
R7524 Transmission_Gate_Layout_11.VIN.n56 Transmission_Gate_Layout_11.VIN.t7 0.7285
R7525 Transmission_Gate_Layout_11.VIN.n56 Transmission_Gate_Layout_11.VIN.n55 0.7285
R7526 Transmission_Gate_Layout_11.VIN.n58 Transmission_Gate_Layout_11.VIN.t68 0.7285
R7527 Transmission_Gate_Layout_11.VIN.n58 Transmission_Gate_Layout_11.VIN.n57 0.7285
R7528 Transmission_Gate_Layout_11.VIN.n9 Transmission_Gate_Layout_11.VIN.t28 0.7285
R7529 Transmission_Gate_Layout_11.VIN.n9 Transmission_Gate_Layout_11.VIN.n8 0.7285
R7530 Transmission_Gate_Layout_11.VIN.n11 Transmission_Gate_Layout_11.VIN.t21 0.7285
R7531 Transmission_Gate_Layout_11.VIN.n11 Transmission_Gate_Layout_11.VIN.n10 0.7285
R7532 Transmission_Gate_Layout_11.VIN.n13 Transmission_Gate_Layout_11.VIN.t35 0.7285
R7533 Transmission_Gate_Layout_11.VIN.n13 Transmission_Gate_Layout_11.VIN.n12 0.7285
R7534 Transmission_Gate_Layout_11.VIN.n127 Transmission_Gate_Layout_11.VIN.t33 0.7285
R7535 Transmission_Gate_Layout_11.VIN.n127 Transmission_Gate_Layout_11.VIN.n126 0.7285
R7536 Transmission_Gate_Layout_11.VIN.n124 Transmission_Gate_Layout_11.VIN.t18 0.7285
R7537 Transmission_Gate_Layout_11.VIN.n124 Transmission_Gate_Layout_11.VIN.n123 0.7285
R7538 Transmission_Gate_Layout_11.VIN.n122 Transmission_Gate_Layout_11.VIN.t25 0.7285
R7539 Transmission_Gate_Layout_11.VIN.n122 Transmission_Gate_Layout_11.VIN.n121 0.7285
R7540 Transmission_Gate_Layout_11.VIN.n132 Transmission_Gate_Layout_11.VIN.t36 0.7285
R7541 Transmission_Gate_Layout_11.VIN.n132 Transmission_Gate_Layout_11.VIN.n131 0.7285
R7542 Transmission_Gate_Layout_11.VIN.n80 Transmission_Gate_Layout_11.VIN.n79 0.626587
R7543 Transmission_Gate_Layout_11.VIN.n82 Transmission_Gate_Layout_11.VIN.n81 0.626587
R7544 Transmission_Gate_Layout_11.VIN.n142 Transmission_Gate_Layout_11.VIN.n141 0.626587
R7545 Transmission_Gate_Layout_11.VIN.n70 Transmission_Gate_Layout_11.VIN 0.607022
R7546 Transmission_Gate_Layout_11.VIN.n95 Transmission_Gate_Layout_11.VIN.n94 0.597239
R7547 Transmission_Gate_Layout_11.VIN.n80 Transmission_Gate_Layout_11.VIN.n52 0.575717
R7548 Transmission_Gate_Layout_11.VIN.n75 Transmission_Gate_Layout_11.VIN.n68 0.575717
R7549 Transmission_Gate_Layout_11.VIN.n79 Transmission_Gate_Layout_11.VIN.n60 0.575717
R7550 Transmission_Gate_Layout_11.VIN.n137 Transmission_Gate_Layout_11.VIN.n136 0.575717
R7551 Transmission_Gate_Layout_11.VIN.n105 Transmission_Gate_Layout_11.VIN.n104 0.570002
R7552 Transmission_Gate_Layout_11.VIN.n141 Transmission_Gate_Layout_11.VIN.n114 0.428978
R7553 Transmission_Gate_Layout_11.VIN.n142 Transmission_Gate_Layout_11.VIN.n7 0.428978
R7554 Transmission_Gate_Layout_11.VIN.n81 Transmission_Gate_Layout_11.VIN.n44 0.331152
R7555 Transmission_Gate_Layout_11.VIN.n82 Transmission_Gate_Layout_11.VIN.n36 0.331152
R7556 Transmission_Gate_Layout_11.VIN.n94 Transmission_Gate_Layout_11.VIN.n93 0.331152
R7557 Transmission_Gate_Layout_11.VIN.n105 Transmission_Gate_Layout_11.VIN.n23 0.331152
R7558 Transmission_Gate_Layout_11.VIN.n104 Transmission_Gate_Layout_11.VIN.n103 0.317457
R7559 Transmission_Gate_Layout_11.VIN.n95 Transmission_Gate_Layout_11.VIN.n28 0.301804
R7560 Transmission_Gate_Layout_11.VIN.n81 Transmission_Gate_Layout_11.VIN.n80 0.239196
R7561 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.VIN.n142 0.192239
R7562 Transmission_Gate_Layout_1.CLK.t32 Transmission_Gate_Layout_1.CLK.t26 82.9076
R7563 Transmission_Gate_Layout_1.CLK.t6 Transmission_Gate_Layout_1.CLK.t32 82.9076
R7564 Transmission_Gate_Layout_1.CLK.t46 Transmission_Gate_Layout_1.CLK.t40 82.9076
R7565 Transmission_Gate_Layout_1.CLK.t17 Transmission_Gate_Layout_1.CLK.t46 82.9076
R7566 Transmission_Gate_Layout_1.CLK.t3 Transmission_Gate_Layout_1.CLK.n32 56.4451
R7567 Transmission_Gate_Layout_1.CLK.n25 Transmission_Gate_Layout_1.CLK.t6 49.7969
R7568 Transmission_Gate_Layout_1.CLK.n51 Transmission_Gate_Layout_1.CLK.t17 49.7969
R7569 Transmission_Gate_Layout_1.CLK.n26 Transmission_Gate_Layout_1.CLK.t8 39.7594
R7570 Transmission_Gate_Layout_1.CLK.n24 Transmission_Gate_Layout_1.CLK.n23 35.0405
R7571 Transmission_Gate_Layout_1.CLK.n34 Transmission_Gate_Layout_1.CLK.n33 35.0405
R7572 Transmission_Gate_Layout_1.CLK.n50 Transmission_Gate_Layout_1.CLK.n49 35.0405
R7573 Transmission_Gate_Layout_1.CLK.n25 Transmission_Gate_Layout_1.CLK.t28 31.1559
R7574 Transmission_Gate_Layout_1.CLK.n51 Transmission_Gate_Layout_1.CLK.t42 31.1559
R7575 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_1.CLK.n53 24.3453
R7576 Transmission_Gate_Layout_1.CLK.n52 Transmission_Gate_Layout_1.CLK.t34 22.0309
R7577 Transmission_Gate_Layout_1.CLK.t10 Transmission_Gate_Layout_1.CLK.n0 21.9005
R7578 Transmission_Gate_Layout_1.CLK.t39 Transmission_Gate_Layout_1.CLK.n15 21.9005
R7579 Transmission_Gate_Layout_1.CLK.t29 Transmission_Gate_Layout_1.CLK.n41 21.9005
R7580 Transmission_Gate_Layout_1.CLK.n40 Transmission_Gate_Layout_1.CLK.t44 21.9005
R7581 Transmission_Gate_Layout_1.CLK.n39 Transmission_Gate_Layout_1.CLK.t21 21.9005
R7582 Transmission_Gate_Layout_1.CLK.n38 Transmission_Gate_Layout_1.CLK.t35 21.9005
R7583 Transmission_Gate_Layout_1.CLK.n37 Transmission_Gate_Layout_1.CLK.t50 21.9005
R7584 Transmission_Gate_Layout_1.CLK.n36 Transmission_Gate_Layout_1.CLK.t18 21.9005
R7585 Transmission_Gate_Layout_1.CLK.n35 Transmission_Gate_Layout_1.CLK.t33 21.9005
R7586 Transmission_Gate_Layout_1.CLK.n33 Transmission_Gate_Layout_1.CLK.t24 21.9005
R7587 Transmission_Gate_Layout_1.CLK.n34 Transmission_Gate_Layout_1.CLK.t5 21.9005
R7588 Transmission_Gate_Layout_1.CLK.n24 Transmission_Gate_Layout_1.CLK.t10 21.5094
R7589 Transmission_Gate_Layout_1.CLK.n23 Transmission_Gate_Layout_1.CLK.t39 21.5094
R7590 Transmission_Gate_Layout_1.CLK.n22 Transmission_Gate_Layout_1.CLK.t60 21.5094
R7591 Transmission_Gate_Layout_1.CLK.n21 Transmission_Gate_Layout_1.CLK.t30 21.5094
R7592 Transmission_Gate_Layout_1.CLK.n20 Transmission_Gate_Layout_1.CLK.t45 21.5094
R7593 Transmission_Gate_Layout_1.CLK.n19 Transmission_Gate_Layout_1.CLK.t59 21.5094
R7594 Transmission_Gate_Layout_1.CLK.n18 Transmission_Gate_Layout_1.CLK.t27 21.5094
R7595 Transmission_Gate_Layout_1.CLK.n17 Transmission_Gate_Layout_1.CLK.t43 21.5094
R7596 Transmission_Gate_Layout_1.CLK.n16 Transmission_Gate_Layout_1.CLK.t13 21.5094
R7597 Transmission_Gate_Layout_1.CLK.n42 Transmission_Gate_Layout_1.CLK.t29 21.5094
R7598 Transmission_Gate_Layout_1.CLK.n43 Transmission_Gate_Layout_1.CLK.t44 21.5094
R7599 Transmission_Gate_Layout_1.CLK.n44 Transmission_Gate_Layout_1.CLK.t21 21.5094
R7600 Transmission_Gate_Layout_1.CLK.n45 Transmission_Gate_Layout_1.CLK.t35 21.5094
R7601 Transmission_Gate_Layout_1.CLK.n46 Transmission_Gate_Layout_1.CLK.t50 21.5094
R7602 Transmission_Gate_Layout_1.CLK.n47 Transmission_Gate_Layout_1.CLK.t18 21.5094
R7603 Transmission_Gate_Layout_1.CLK.n48 Transmission_Gate_Layout_1.CLK.t33 21.5094
R7604 Transmission_Gate_Layout_1.CLK.n50 Transmission_Gate_Layout_1.CLK.t24 21.5094
R7605 Transmission_Gate_Layout_1.CLK.n49 Transmission_Gate_Layout_1.CLK.t5 21.5094
R7606 Transmission_Gate_Layout_1.CLK.n53 Transmission_Gate_Layout_1.CLK.t57 21.3791
R7607 Transmission_Gate_Layout_1.CLK.n52 Transmission_Gate_Layout_1.CLK.t55 21.3791
R7608 Transmission_Gate_Layout_1.CLK.n23 Transmission_Gate_Layout_1.CLK.t58 20.988
R7609 Transmission_Gate_Layout_1.CLK.n22 Transmission_Gate_Layout_1.CLK.t15 20.988
R7610 Transmission_Gate_Layout_1.CLK.n21 Transmission_Gate_Layout_1.CLK.t51 20.988
R7611 Transmission_Gate_Layout_1.CLK.n20 Transmission_Gate_Layout_1.CLK.t64 20.988
R7612 Transmission_Gate_Layout_1.CLK.n19 Transmission_Gate_Layout_1.CLK.t12 20.988
R7613 Transmission_Gate_Layout_1.CLK.n18 Transmission_Gate_Layout_1.CLK.t48 20.988
R7614 Transmission_Gate_Layout_1.CLK.n17 Transmission_Gate_Layout_1.CLK.t61 20.988
R7615 Transmission_Gate_Layout_1.CLK.n16 Transmission_Gate_Layout_1.CLK.t31 20.988
R7616 Transmission_Gate_Layout_1.CLK.t28 Transmission_Gate_Layout_1.CLK.n24 20.988
R7617 Transmission_Gate_Layout_1.CLK.n42 Transmission_Gate_Layout_1.CLK.t49 20.988
R7618 Transmission_Gate_Layout_1.CLK.n43 Transmission_Gate_Layout_1.CLK.t62 20.988
R7619 Transmission_Gate_Layout_1.CLK.n44 Transmission_Gate_Layout_1.CLK.t41 20.988
R7620 Transmission_Gate_Layout_1.CLK.n45 Transmission_Gate_Layout_1.CLK.t54 20.988
R7621 Transmission_Gate_Layout_1.CLK.n46 Transmission_Gate_Layout_1.CLK.t4 20.988
R7622 Transmission_Gate_Layout_1.CLK.n47 Transmission_Gate_Layout_1.CLK.t38 20.988
R7623 Transmission_Gate_Layout_1.CLK.n48 Transmission_Gate_Layout_1.CLK.t52 20.988
R7624 Transmission_Gate_Layout_1.CLK.n49 Transmission_Gate_Layout_1.CLK.t23 20.988
R7625 Transmission_Gate_Layout_1.CLK.t42 Transmission_Gate_Layout_1.CLK.n50 20.988
R7626 Transmission_Gate_Layout_1.CLK.n27 Transmission_Gate_Layout_1.CLK.n26 20.8576
R7627 Transmission_Gate_Layout_1.CLK.n28 Transmission_Gate_Layout_1.CLK.n27 20.8576
R7628 Transmission_Gate_Layout_1.CLK.n29 Transmission_Gate_Layout_1.CLK.n28 20.8576
R7629 Transmission_Gate_Layout_1.CLK.n30 Transmission_Gate_Layout_1.CLK.n29 20.8576
R7630 Transmission_Gate_Layout_1.CLK.n31 Transmission_Gate_Layout_1.CLK.n30 20.8576
R7631 Transmission_Gate_Layout_1.CLK.n32 Transmission_Gate_Layout_1.CLK.n31 20.8576
R7632 Transmission_Gate_Layout_1.CLK.n53 Transmission_Gate_Layout_1.CLK.n52 20.8576
R7633 Transmission_Gate_Layout_1.CLK.n0 Transmission_Gate_Layout_1.CLK.t53 20.5969
R7634 Transmission_Gate_Layout_1.CLK.n15 Transmission_Gate_Layout_1.CLK.t16 20.5969
R7635 Transmission_Gate_Layout_1.CLK.n14 Transmission_Gate_Layout_1.CLK.t37 20.5969
R7636 Transmission_Gate_Layout_1.CLK.n13 Transmission_Gate_Layout_1.CLK.t9 20.5969
R7637 Transmission_Gate_Layout_1.CLK.n12 Transmission_Gate_Layout_1.CLK.t22 20.5969
R7638 Transmission_Gate_Layout_1.CLK.n11 Transmission_Gate_Layout_1.CLK.t36 20.5969
R7639 Transmission_Gate_Layout_1.CLK.n10 Transmission_Gate_Layout_1.CLK.t7 20.5969
R7640 Transmission_Gate_Layout_1.CLK.n8 Transmission_Gate_Layout_1.CLK.t56 20.5969
R7641 Transmission_Gate_Layout_1.CLK.n9 Transmission_Gate_Layout_1.CLK.t19 20.5969
R7642 Transmission_Gate_Layout_1.CLK.n41 Transmission_Gate_Layout_1.CLK.t8 20.5969
R7643 Transmission_Gate_Layout_1.CLK.n40 Transmission_Gate_Layout_1.CLK.t20 20.5969
R7644 Transmission_Gate_Layout_1.CLK.n39 Transmission_Gate_Layout_1.CLK.t2 20.5969
R7645 Transmission_Gate_Layout_1.CLK.n38 Transmission_Gate_Layout_1.CLK.t14 20.5969
R7646 Transmission_Gate_Layout_1.CLK.n37 Transmission_Gate_Layout_1.CLK.t25 20.5969
R7647 Transmission_Gate_Layout_1.CLK.n36 Transmission_Gate_Layout_1.CLK.t63 20.5969
R7648 Transmission_Gate_Layout_1.CLK.n35 Transmission_Gate_Layout_1.CLK.t11 20.5969
R7649 Transmission_Gate_Layout_1.CLK.n34 Transmission_Gate_Layout_1.CLK.t47 20.5969
R7650 Transmission_Gate_Layout_1.CLK.n33 Transmission_Gate_Layout_1.CLK.t3 20.5969
R7651 Transmission_Gate_Layout_1.CLK.n15 Transmission_Gate_Layout_1.CLK.n14 19.4672
R7652 Transmission_Gate_Layout_1.CLK.n14 Transmission_Gate_Layout_1.CLK.n13 19.4672
R7653 Transmission_Gate_Layout_1.CLK.n13 Transmission_Gate_Layout_1.CLK.n12 19.4672
R7654 Transmission_Gate_Layout_1.CLK.n12 Transmission_Gate_Layout_1.CLK.n11 19.4672
R7655 Transmission_Gate_Layout_1.CLK.n11 Transmission_Gate_Layout_1.CLK.n10 19.4672
R7656 Transmission_Gate_Layout_1.CLK.n10 Transmission_Gate_Layout_1.CLK.n9 19.4672
R7657 Transmission_Gate_Layout_1.CLK.n9 Transmission_Gate_Layout_1.CLK.n8 19.4672
R7658 Transmission_Gate_Layout_1.CLK.n23 Transmission_Gate_Layout_1.CLK.n22 19.4672
R7659 Transmission_Gate_Layout_1.CLK.n22 Transmission_Gate_Layout_1.CLK.n21 19.4672
R7660 Transmission_Gate_Layout_1.CLK.n21 Transmission_Gate_Layout_1.CLK.n20 19.4672
R7661 Transmission_Gate_Layout_1.CLK.n20 Transmission_Gate_Layout_1.CLK.n19 19.4672
R7662 Transmission_Gate_Layout_1.CLK.n19 Transmission_Gate_Layout_1.CLK.n18 19.4672
R7663 Transmission_Gate_Layout_1.CLK.n18 Transmission_Gate_Layout_1.CLK.n17 19.4672
R7664 Transmission_Gate_Layout_1.CLK.n17 Transmission_Gate_Layout_1.CLK.n16 19.4672
R7665 Transmission_Gate_Layout_1.CLK.n41 Transmission_Gate_Layout_1.CLK.n40 19.4672
R7666 Transmission_Gate_Layout_1.CLK.n40 Transmission_Gate_Layout_1.CLK.n39 19.4672
R7667 Transmission_Gate_Layout_1.CLK.n39 Transmission_Gate_Layout_1.CLK.n38 19.4672
R7668 Transmission_Gate_Layout_1.CLK.n38 Transmission_Gate_Layout_1.CLK.n37 19.4672
R7669 Transmission_Gate_Layout_1.CLK.n37 Transmission_Gate_Layout_1.CLK.n36 19.4672
R7670 Transmission_Gate_Layout_1.CLK.n36 Transmission_Gate_Layout_1.CLK.n35 19.4672
R7671 Transmission_Gate_Layout_1.CLK.n35 Transmission_Gate_Layout_1.CLK.n34 19.4672
R7672 Transmission_Gate_Layout_1.CLK.n43 Transmission_Gate_Layout_1.CLK.n42 19.4672
R7673 Transmission_Gate_Layout_1.CLK.n44 Transmission_Gate_Layout_1.CLK.n43 19.4672
R7674 Transmission_Gate_Layout_1.CLK.n45 Transmission_Gate_Layout_1.CLK.n44 19.4672
R7675 Transmission_Gate_Layout_1.CLK.n46 Transmission_Gate_Layout_1.CLK.n45 19.4672
R7676 Transmission_Gate_Layout_1.CLK.n47 Transmission_Gate_Layout_1.CLK.n46 19.4672
R7677 Transmission_Gate_Layout_1.CLK.n48 Transmission_Gate_Layout_1.CLK.n47 19.4672
R7678 Transmission_Gate_Layout_1.CLK.n49 Transmission_Gate_Layout_1.CLK.n48 19.4672
R7679 Transmission_Gate_Layout_1.CLK.t16 Transmission_Gate_Layout_1.CLK.n1 18.9023
R7680 Transmission_Gate_Layout_1.CLK.t37 Transmission_Gate_Layout_1.CLK.n2 18.9023
R7681 Transmission_Gate_Layout_1.CLK.t9 Transmission_Gate_Layout_1.CLK.n3 18.9023
R7682 Transmission_Gate_Layout_1.CLK.t22 Transmission_Gate_Layout_1.CLK.n4 18.9023
R7683 Transmission_Gate_Layout_1.CLK.t36 Transmission_Gate_Layout_1.CLK.n5 18.9023
R7684 Transmission_Gate_Layout_1.CLK.t7 Transmission_Gate_Layout_1.CLK.n6 18.9023
R7685 Transmission_Gate_Layout_1.CLK.t19 Transmission_Gate_Layout_1.CLK.n7 18.9023
R7686 Transmission_Gate_Layout_1.CLK.n26 Transmission_Gate_Layout_1.CLK.t20 18.9023
R7687 Transmission_Gate_Layout_1.CLK.n27 Transmission_Gate_Layout_1.CLK.t2 18.9023
R7688 Transmission_Gate_Layout_1.CLK.n28 Transmission_Gate_Layout_1.CLK.t14 18.9023
R7689 Transmission_Gate_Layout_1.CLK.n29 Transmission_Gate_Layout_1.CLK.t25 18.9023
R7690 Transmission_Gate_Layout_1.CLK.n30 Transmission_Gate_Layout_1.CLK.t63 18.9023
R7691 Transmission_Gate_Layout_1.CLK.n31 Transmission_Gate_Layout_1.CLK.t11 18.9023
R7692 Transmission_Gate_Layout_1.CLK.n32 Transmission_Gate_Layout_1.CLK.t47 18.9023
R7693 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_1.CLK.n51 17.6496
R7694 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_1.CLK.n25 16.6488
R7695 Transmission_Gate_Layout_1.CLK.n56 Transmission_Gate_Layout_1.CLK 9.13953
R7696 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_1.CLK.n54 7.70137
R7697 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_1.CLK.n55 4.70224
R7698 Transmission_Gate_Layout_1.CLK.n56 Transmission_Gate_Layout_1.CLK 0.608978
R7699 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_1.CLK.n56 0.248978
R7700 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.t5 17.8546
R7701 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n0 14.0337
R7702 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.t4 13.5862
R7703 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n2 3.76289
R7704 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n2 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.t0 3.2765
R7705 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n2 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n1 3.2765
R7706 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n4 2.88224
R7707 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n4 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.t2 1.8205
R7708 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n4 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT.n3 1.8205
R7709 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.n3 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.n0 5.61007
R7710 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.t3 5.01528
R7711 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.n3 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.n2 2.6005
R7712 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.n2 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.t0 1.8205
R7713 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.n2 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.n1 1.8205
R7714 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1.n3 0.595283
R7715 IN7.n59 IN7 13.868
R7716 IN7.n56 IN7.n55 3.90572
R7717 IN7.n48 IN7.n47 3.90572
R7718 IN7.n4 IN7.n1 3.90572
R7719 IN7.n26 IN7.n23 3.84485
R7720 IN7.n34 IN7.n31 3.84485
R7721 IN7.n14 IN7.n13 3.84485
R7722 IN7.n56 IN7.n53 3.1505
R7723 IN7.n57 IN7.n51 3.1505
R7724 IN7.n48 IN7.n45 3.1505
R7725 IN7.n49 IN7.n43 3.1505
R7726 IN7.n4 IN7.n3 3.1505
R7727 IN7.n7 IN7.n6 3.1505
R7728 IN7.n68 IN7.n67 3.1505
R7729 IN7.n65 IN7.n64 3.1505
R7730 IN7.n62 IN7.n61 3.1505
R7731 IN7.n26 IN7.n25 2.6005
R7732 IN7.n29 IN7.n28 2.6005
R7733 IN7.n34 IN7.n33 2.6005
R7734 IN7.n37 IN7.n36 2.6005
R7735 IN7.n39 IN7.n21 2.6005
R7736 IN7.n40 IN7.n19 2.6005
R7737 IN7.n41 IN7.n17 2.6005
R7738 IN7.n14 IN7.n11 2.6005
R7739 IN7.n15 IN7.n9 2.6005
R7740 IN7.n51 IN7.t31 1.3109
R7741 IN7.n51 IN7.n50 1.3109
R7742 IN7.n53 IN7.t27 1.3109
R7743 IN7.n53 IN7.n52 1.3109
R7744 IN7.n55 IN7.t24 1.3109
R7745 IN7.n55 IN7.n54 1.3109
R7746 IN7.n43 IN7.t34 1.3109
R7747 IN7.n43 IN7.n42 1.3109
R7748 IN7.n45 IN7.t32 1.3109
R7749 IN7.n45 IN7.n44 1.3109
R7750 IN7.n47 IN7.t28 1.3109
R7751 IN7.n47 IN7.n46 1.3109
R7752 IN7.n61 IN7.t30 1.3109
R7753 IN7.n61 IN7.n60 1.3109
R7754 IN7.n64 IN7.t26 1.3109
R7755 IN7.n64 IN7.n63 1.3109
R7756 IN7.n67 IN7.t35 1.3109
R7757 IN7.n67 IN7.n66 1.3109
R7758 IN7.n6 IN7.t33 1.3109
R7759 IN7.n6 IN7.n5 1.3109
R7760 IN7.n3 IN7.t25 1.3109
R7761 IN7.n3 IN7.n2 1.3109
R7762 IN7.n1 IN7.t29 1.3109
R7763 IN7.n1 IN7.n0 1.3109
R7764 IN7.n29 IN7.n26 1.24485
R7765 IN7.n37 IN7.n34 1.24485
R7766 IN7.n41 IN7.n40 1.24485
R7767 IN7.n40 IN7.n39 1.24485
R7768 IN7.n15 IN7.n14 1.24485
R7769 IN7.n38 IN7.n37 1.2018
R7770 IN7.n39 IN7.n38 1.2018
R7771 IN7.n58 IN7.n57 0.957239
R7772 IN7.n69 IN7.n41 0.806587
R7773 IN7.n70 IN7.n15 0.806587
R7774 IN7.n57 IN7.n56 0.755717
R7775 IN7.n49 IN7.n48 0.755717
R7776 IN7.n7 IN7.n4 0.755717
R7777 IN7.n65 IN7.n62 0.755717
R7778 IN7.n68 IN7.n65 0.755717
R7779 IN7.n17 IN7.t14 0.7285
R7780 IN7.n17 IN7.n16 0.7285
R7781 IN7.n19 IN7.t6 0.7285
R7782 IN7.n19 IN7.n18 0.7285
R7783 IN7.n21 IN7.t18 0.7285
R7784 IN7.n21 IN7.n20 0.7285
R7785 IN7.n28 IN7.t8 0.7285
R7786 IN7.n28 IN7.n27 0.7285
R7787 IN7.n25 IN7.t23 0.7285
R7788 IN7.n25 IN7.n24 0.7285
R7789 IN7.n23 IN7.t2 0.7285
R7790 IN7.n23 IN7.n22 0.7285
R7791 IN7.n36 IN7.t16 0.7285
R7792 IN7.n36 IN7.n35 0.7285
R7793 IN7.n33 IN7.t3 0.7285
R7794 IN7.n33 IN7.n32 0.7285
R7795 IN7.n31 IN7.t10 0.7285
R7796 IN7.n31 IN7.n30 0.7285
R7797 IN7.n9 IN7.t15 0.7285
R7798 IN7.n9 IN7.n8 0.7285
R7799 IN7.n11 IN7.t7 0.7285
R7800 IN7.n11 IN7.n10 0.7285
R7801 IN7.n13 IN7.t19 0.7285
R7802 IN7.n13 IN7.n12 0.7285
R7803 IN7.n70 IN7.n69 0.626587
R7804 IN7.n38 IN7.n29 0.575717
R7805 IN7.n59 IN7.n58 0.570002
R7806 IN7.n70 IN7.n7 0.428978
R7807 IN7.n69 IN7.n68 0.428978
R7808 IN7.n58 IN7.n49 0.331152
R7809 IN7.n62 IN7.n59 0.317457
R7810 IN7 IN7.n70 0.192239
R7811 Transmission_Gate_Layout_4.VIN.n96 Transmission_Gate_Layout_4.VIN.n87 5.27032
R7812 Transmission_Gate_Layout_4.VIN.n51 Transmission_Gate_Layout_4.VIN.n50 5.21612
R7813 Transmission_Gate_Layout_4.VIN.n54 Transmission_Gate_Layout_4.VIN.t84 4.4609
R7814 Transmission_Gate_Layout_4.VIN.n55 Transmission_Gate_Layout_4.VIN.t78 4.4609
R7815 Transmission_Gate_Layout_4.VIN.n56 Transmission_Gate_Layout_4.VIN.t72 4.4609
R7816 Transmission_Gate_Layout_4.VIN.n52 Transmission_Gate_Layout_4.VIN.n48 4.4609
R7817 Transmission_Gate_Layout_4.VIN.n51 Transmission_Gate_Layout_4.VIN.n49 4.4609
R7818 Transmission_Gate_Layout_4.VIN.n117 Transmission_Gate_Layout_4.VIN.n114 3.90572
R7819 Transmission_Gate_Layout_4.VIN.n125 Transmission_Gate_Layout_4.VIN.n122 3.90572
R7820 Transmission_Gate_Layout_4.VIN.n28 Transmission_Gate_Layout_4.VIN.n25 3.90572
R7821 Transmission_Gate_Layout_4.VIN.n36 Transmission_Gate_Layout_4.VIN.n33 3.90572
R7822 Transmission_Gate_Layout_4.VIN.n46 Transmission_Gate_Layout_4.VIN.n45 3.90572
R7823 Transmission_Gate_Layout_4.VIN.n140 Transmission_Gate_Layout_4.VIN.n137 3.90572
R7824 Transmission_Gate_Layout_4.VIN.n4 Transmission_Gate_Layout_4.VIN.n1 3.84485
R7825 Transmission_Gate_Layout_4.VIN.n76 Transmission_Gate_Layout_4.VIN.n73 3.84485
R7826 Transmission_Gate_Layout_4.VIN.n65 Transmission_Gate_Layout_4.VIN.n64 3.84485
R7827 Transmission_Gate_Layout_4.VIN.n22 Transmission_Gate_Layout_4.VIN.n21 3.84485
R7828 Transmission_Gate_Layout_4.VIN.n94 Transmission_Gate_Layout_4.VIN.n93 3.84485
R7829 Transmission_Gate_Layout_4.VIN.n14 Transmission_Gate_Layout_4.VIN.n13 3.84485
R7830 Transmission_Gate_Layout_4.VIN.n85 Transmission_Gate_Layout_4.VIN.n84 3.3285
R7831 Transmission_Gate_Layout_4.VIN.n83 Transmission_Gate_Layout_4.VIN.n82 3.3285
R7832 Transmission_Gate_Layout_4.VIN.n81 Transmission_Gate_Layout_4.VIN.n80 3.3285
R7833 Transmission_Gate_Layout_4.VIN.n69 Transmission_Gate_Layout_4.VIN.t11 3.3285
R7834 Transmission_Gate_Layout_4.VIN.n70 Transmission_Gate_Layout_4.VIN.t5 3.3285
R7835 Transmission_Gate_Layout_4.VIN.n71 Transmission_Gate_Layout_4.VIN.t26 3.3285
R7836 Transmission_Gate_Layout_4.VIN.n117 Transmission_Gate_Layout_4.VIN.n116 3.1505
R7837 Transmission_Gate_Layout_4.VIN.n120 Transmission_Gate_Layout_4.VIN.n119 3.1505
R7838 Transmission_Gate_Layout_4.VIN.n125 Transmission_Gate_Layout_4.VIN.n124 3.1505
R7839 Transmission_Gate_Layout_4.VIN.n128 Transmission_Gate_Layout_4.VIN.n127 3.1505
R7840 Transmission_Gate_Layout_4.VIN.n28 Transmission_Gate_Layout_4.VIN.n27 3.1505
R7841 Transmission_Gate_Layout_4.VIN.n31 Transmission_Gate_Layout_4.VIN.n30 3.1505
R7842 Transmission_Gate_Layout_4.VIN.n36 Transmission_Gate_Layout_4.VIN.n35 3.1505
R7843 Transmission_Gate_Layout_4.VIN.n39 Transmission_Gate_Layout_4.VIN.n38 3.1505
R7844 Transmission_Gate_Layout_4.VIN.n46 Transmission_Gate_Layout_4.VIN.n43 3.1505
R7845 Transmission_Gate_Layout_4.VIN.n47 Transmission_Gate_Layout_4.VIN.n41 3.1505
R7846 Transmission_Gate_Layout_4.VIN.n130 Transmission_Gate_Layout_4.VIN.n112 3.1505
R7847 Transmission_Gate_Layout_4.VIN.n131 Transmission_Gate_Layout_4.VIN.n110 3.1505
R7848 Transmission_Gate_Layout_4.VIN.n132 Transmission_Gate_Layout_4.VIN.n108 3.1505
R7849 Transmission_Gate_Layout_4.VIN.n141 Transmission_Gate_Layout_4.VIN.n135 3.1505
R7850 Transmission_Gate_Layout_4.VIN.n140 Transmission_Gate_Layout_4.VIN.n139 3.1505
R7851 Transmission_Gate_Layout_4.VIN.n4 Transmission_Gate_Layout_4.VIN.n3 2.6005
R7852 Transmission_Gate_Layout_4.VIN.n7 Transmission_Gate_Layout_4.VIN.n6 2.6005
R7853 Transmission_Gate_Layout_4.VIN.n76 Transmission_Gate_Layout_4.VIN.n75 2.6005
R7854 Transmission_Gate_Layout_4.VIN.n79 Transmission_Gate_Layout_4.VIN.n78 2.6005
R7855 Transmission_Gate_Layout_4.VIN.n65 Transmission_Gate_Layout_4.VIN.n62 2.6005
R7856 Transmission_Gate_Layout_4.VIN.n66 Transmission_Gate_Layout_4.VIN.n60 2.6005
R7857 Transmission_Gate_Layout_4.VIN.n22 Transmission_Gate_Layout_4.VIN.n19 2.6005
R7858 Transmission_Gate_Layout_4.VIN.n23 Transmission_Gate_Layout_4.VIN.n17 2.6005
R7859 Transmission_Gate_Layout_4.VIN.n94 Transmission_Gate_Layout_4.VIN.n91 2.6005
R7860 Transmission_Gate_Layout_4.VIN.n95 Transmission_Gate_Layout_4.VIN.n89 2.6005
R7861 Transmission_Gate_Layout_4.VIN.n14 Transmission_Gate_Layout_4.VIN.n11 2.6005
R7862 Transmission_Gate_Layout_4.VIN.n15 Transmission_Gate_Layout_4.VIN.n9 2.6005
R7863 Transmission_Gate_Layout_4.VIN.n106 Transmission_Gate_Layout_4.VIN.n105 2.6005
R7864 Transmission_Gate_Layout_4.VIN.n103 Transmission_Gate_Layout_4.VIN.n102 2.6005
R7865 Transmission_Gate_Layout_4.VIN.n100 Transmission_Gate_Layout_4.VIN.n99 2.6005
R7866 Transmission_Gate_Layout_4.VIN.n54 Transmission_Gate_Layout_4.VIN.n53 2.47941
R7867 Transmission_Gate_Layout_4.VIN.n87 Transmission_Gate_Layout_4.VIN.n86 1.90239
R7868 Transmission_Gate_Layout_4.VIN.n135 Transmission_Gate_Layout_4.VIN.t37 1.3109
R7869 Transmission_Gate_Layout_4.VIN.n135 Transmission_Gate_Layout_4.VIN.n134 1.3109
R7870 Transmission_Gate_Layout_4.VIN.n137 Transmission_Gate_Layout_4.VIN.t51 1.3109
R7871 Transmission_Gate_Layout_4.VIN.n137 Transmission_Gate_Layout_4.VIN.n136 1.3109
R7872 Transmission_Gate_Layout_4.VIN.n108 Transmission_Gate_Layout_4.VIN.t38 1.3109
R7873 Transmission_Gate_Layout_4.VIN.n108 Transmission_Gate_Layout_4.VIN.n107 1.3109
R7874 Transmission_Gate_Layout_4.VIN.n110 Transmission_Gate_Layout_4.VIN.t48 1.3109
R7875 Transmission_Gate_Layout_4.VIN.n110 Transmission_Gate_Layout_4.VIN.n109 1.3109
R7876 Transmission_Gate_Layout_4.VIN.n112 Transmission_Gate_Layout_4.VIN.t32 1.3109
R7877 Transmission_Gate_Layout_4.VIN.n112 Transmission_Gate_Layout_4.VIN.n111 1.3109
R7878 Transmission_Gate_Layout_4.VIN.n119 Transmission_Gate_Layout_4.VIN.t31 1.3109
R7879 Transmission_Gate_Layout_4.VIN.n119 Transmission_Gate_Layout_4.VIN.n118 1.3109
R7880 Transmission_Gate_Layout_4.VIN.n116 Transmission_Gate_Layout_4.VIN.t44 1.3109
R7881 Transmission_Gate_Layout_4.VIN.n116 Transmission_Gate_Layout_4.VIN.n115 1.3109
R7882 Transmission_Gate_Layout_4.VIN.n114 Transmission_Gate_Layout_4.VIN.t47 1.3109
R7883 Transmission_Gate_Layout_4.VIN.n114 Transmission_Gate_Layout_4.VIN.n113 1.3109
R7884 Transmission_Gate_Layout_4.VIN.n127 Transmission_Gate_Layout_4.VIN.t45 1.3109
R7885 Transmission_Gate_Layout_4.VIN.n127 Transmission_Gate_Layout_4.VIN.n126 1.3109
R7886 Transmission_Gate_Layout_4.VIN.n124 Transmission_Gate_Layout_4.VIN.t35 1.3109
R7887 Transmission_Gate_Layout_4.VIN.n124 Transmission_Gate_Layout_4.VIN.n123 1.3109
R7888 Transmission_Gate_Layout_4.VIN.n122 Transmission_Gate_Layout_4.VIN.t41 1.3109
R7889 Transmission_Gate_Layout_4.VIN.n122 Transmission_Gate_Layout_4.VIN.n121 1.3109
R7890 Transmission_Gate_Layout_4.VIN.n30 Transmission_Gate_Layout_4.VIN.t89 1.3109
R7891 Transmission_Gate_Layout_4.VIN.n30 Transmission_Gate_Layout_4.VIN.n29 1.3109
R7892 Transmission_Gate_Layout_4.VIN.n27 Transmission_Gate_Layout_4.VIN.t94 1.3109
R7893 Transmission_Gate_Layout_4.VIN.n27 Transmission_Gate_Layout_4.VIN.n26 1.3109
R7894 Transmission_Gate_Layout_4.VIN.n25 Transmission_Gate_Layout_4.VIN.t76 1.3109
R7895 Transmission_Gate_Layout_4.VIN.n25 Transmission_Gate_Layout_4.VIN.n24 1.3109
R7896 Transmission_Gate_Layout_4.VIN.n38 Transmission_Gate_Layout_4.VIN.t80 1.3109
R7897 Transmission_Gate_Layout_4.VIN.n38 Transmission_Gate_Layout_4.VIN.n37 1.3109
R7898 Transmission_Gate_Layout_4.VIN.n35 Transmission_Gate_Layout_4.VIN.t86 1.3109
R7899 Transmission_Gate_Layout_4.VIN.n35 Transmission_Gate_Layout_4.VIN.n34 1.3109
R7900 Transmission_Gate_Layout_4.VIN.n33 Transmission_Gate_Layout_4.VIN.t90 1.3109
R7901 Transmission_Gate_Layout_4.VIN.n33 Transmission_Gate_Layout_4.VIN.n32 1.3109
R7902 Transmission_Gate_Layout_4.VIN.n41 Transmission_Gate_Layout_4.VIN.t74 1.3109
R7903 Transmission_Gate_Layout_4.VIN.n41 Transmission_Gate_Layout_4.VIN.n40 1.3109
R7904 Transmission_Gate_Layout_4.VIN.n43 Transmission_Gate_Layout_4.VIN.t91 1.3109
R7905 Transmission_Gate_Layout_4.VIN.n43 Transmission_Gate_Layout_4.VIN.n42 1.3109
R7906 Transmission_Gate_Layout_4.VIN.n45 Transmission_Gate_Layout_4.VIN.t87 1.3109
R7907 Transmission_Gate_Layout_4.VIN.n45 Transmission_Gate_Layout_4.VIN.n44 1.3109
R7908 Transmission_Gate_Layout_4.VIN.n139 Transmission_Gate_Layout_4.VIN.t42 1.3109
R7909 Transmission_Gate_Layout_4.VIN.n139 Transmission_Gate_Layout_4.VIN.n138 1.3109
R7910 Transmission_Gate_Layout_4.VIN.n7 Transmission_Gate_Layout_4.VIN.n4 1.24485
R7911 Transmission_Gate_Layout_4.VIN.n79 Transmission_Gate_Layout_4.VIN.n76 1.24485
R7912 Transmission_Gate_Layout_4.VIN.n83 Transmission_Gate_Layout_4.VIN.n81 1.24485
R7913 Transmission_Gate_Layout_4.VIN.n85 Transmission_Gate_Layout_4.VIN.n83 1.24485
R7914 Transmission_Gate_Layout_4.VIN.n66 Transmission_Gate_Layout_4.VIN.n65 1.24485
R7915 Transmission_Gate_Layout_4.VIN.n23 Transmission_Gate_Layout_4.VIN.n22 1.24485
R7916 Transmission_Gate_Layout_4.VIN.n70 Transmission_Gate_Layout_4.VIN.n69 1.24485
R7917 Transmission_Gate_Layout_4.VIN.n71 Transmission_Gate_Layout_4.VIN.n70 1.24485
R7918 Transmission_Gate_Layout_4.VIN.n95 Transmission_Gate_Layout_4.VIN.n94 1.24485
R7919 Transmission_Gate_Layout_4.VIN.n15 Transmission_Gate_Layout_4.VIN.n14 1.24485
R7920 Transmission_Gate_Layout_4.VIN.n103 Transmission_Gate_Layout_4.VIN.n100 1.24485
R7921 Transmission_Gate_Layout_4.VIN.n106 Transmission_Gate_Layout_4.VIN.n103 1.24485
R7922 Transmission_Gate_Layout_4.VIN.n86 Transmission_Gate_Layout_4.VIN.n85 1.2018
R7923 Transmission_Gate_Layout_4.VIN.n69 Transmission_Gate_Layout_4.VIN.n68 1.2018
R7924 Transmission_Gate_Layout_4.VIN.n100 Transmission_Gate_Layout_4.VIN.n97 1.2018
R7925 Transmission_Gate_Layout_4.VIN.n129 Transmission_Gate_Layout_4.VIN.n128 0.957239
R7926 Transmission_Gate_Layout_4.VIN.n130 Transmission_Gate_Layout_4.VIN.n129 0.957239
R7927 Transmission_Gate_Layout_4.VIN.n53 Transmission_Gate_Layout_4.VIN.n52 0.957239
R7928 Transmission_Gate_Layout_4.VIN.n57 Transmission_Gate_Layout_4.VIN.n56 0.957239
R7929 Transmission_Gate_Layout_4.VIN.n142 Transmission_Gate_Layout_4.VIN.n7 0.806587
R7930 Transmission_Gate_Layout_4.VIN.n133 Transmission_Gate_Layout_4.VIN.n106 0.806587
R7931 Transmission_Gate_Layout_4.VIN.n120 Transmission_Gate_Layout_4.VIN.n117 0.755717
R7932 Transmission_Gate_Layout_4.VIN.n128 Transmission_Gate_Layout_4.VIN.n125 0.755717
R7933 Transmission_Gate_Layout_4.VIN.n31 Transmission_Gate_Layout_4.VIN.n28 0.755717
R7934 Transmission_Gate_Layout_4.VIN.n39 Transmission_Gate_Layout_4.VIN.n36 0.755717
R7935 Transmission_Gate_Layout_4.VIN.n47 Transmission_Gate_Layout_4.VIN.n46 0.755717
R7936 Transmission_Gate_Layout_4.VIN.n52 Transmission_Gate_Layout_4.VIN.n51 0.755717
R7937 Transmission_Gate_Layout_4.VIN.n55 Transmission_Gate_Layout_4.VIN.n54 0.755717
R7938 Transmission_Gate_Layout_4.VIN.n56 Transmission_Gate_Layout_4.VIN.n55 0.755717
R7939 Transmission_Gate_Layout_4.VIN.n132 Transmission_Gate_Layout_4.VIN.n131 0.755717
R7940 Transmission_Gate_Layout_4.VIN.n131 Transmission_Gate_Layout_4.VIN.n130 0.755717
R7941 Transmission_Gate_Layout_4.VIN.n141 Transmission_Gate_Layout_4.VIN.n140 0.755717
R7942 Transmission_Gate_Layout_4.VIN.n87 Transmission_Gate_Layout_4.VIN.n71 0.742022
R7943 Transmission_Gate_Layout_4.VIN.n6 Transmission_Gate_Layout_4.VIN.t63 0.7285
R7944 Transmission_Gate_Layout_4.VIN.n6 Transmission_Gate_Layout_4.VIN.n5 0.7285
R7945 Transmission_Gate_Layout_4.VIN.n3 Transmission_Gate_Layout_4.VIN.t16 0.7285
R7946 Transmission_Gate_Layout_4.VIN.n3 Transmission_Gate_Layout_4.VIN.n2 0.7285
R7947 Transmission_Gate_Layout_4.VIN.n1 Transmission_Gate_Layout_4.VIN.t22 0.7285
R7948 Transmission_Gate_Layout_4.VIN.n1 Transmission_Gate_Layout_4.VIN.n0 0.7285
R7949 Transmission_Gate_Layout_4.VIN.n99 Transmission_Gate_Layout_4.VIN.t21 0.7285
R7950 Transmission_Gate_Layout_4.VIN.n99 Transmission_Gate_Layout_4.VIN.n98 0.7285
R7951 Transmission_Gate_Layout_4.VIN.n102 Transmission_Gate_Layout_4.VIN.t70 0.7285
R7952 Transmission_Gate_Layout_4.VIN.n102 Transmission_Gate_Layout_4.VIN.n101 0.7285
R7953 Transmission_Gate_Layout_4.VIN.n105 Transmission_Gate_Layout_4.VIN.t62 0.7285
R7954 Transmission_Gate_Layout_4.VIN.n105 Transmission_Gate_Layout_4.VIN.n104 0.7285
R7955 Transmission_Gate_Layout_4.VIN.n78 Transmission_Gate_Layout_4.VIN.t1 0.7285
R7956 Transmission_Gate_Layout_4.VIN.n78 Transmission_Gate_Layout_4.VIN.n77 0.7285
R7957 Transmission_Gate_Layout_4.VIN.n75 Transmission_Gate_Layout_4.VIN.t13 0.7285
R7958 Transmission_Gate_Layout_4.VIN.n75 Transmission_Gate_Layout_4.VIN.n74 0.7285
R7959 Transmission_Gate_Layout_4.VIN.n73 Transmission_Gate_Layout_4.VIN.t54 0.7285
R7960 Transmission_Gate_Layout_4.VIN.n73 Transmission_Gate_Layout_4.VIN.n72 0.7285
R7961 Transmission_Gate_Layout_4.VIN.n60 Transmission_Gate_Layout_4.VIN.t53 0.7285
R7962 Transmission_Gate_Layout_4.VIN.n60 Transmission_Gate_Layout_4.VIN.n59 0.7285
R7963 Transmission_Gate_Layout_4.VIN.n62 Transmission_Gate_Layout_4.VIN.t12 0.7285
R7964 Transmission_Gate_Layout_4.VIN.n62 Transmission_Gate_Layout_4.VIN.n61 0.7285
R7965 Transmission_Gate_Layout_4.VIN.n64 Transmission_Gate_Layout_4.VIN.t0 0.7285
R7966 Transmission_Gate_Layout_4.VIN.n64 Transmission_Gate_Layout_4.VIN.n63 0.7285
R7967 Transmission_Gate_Layout_4.VIN.n17 Transmission_Gate_Layout_4.VIN.t4 0.7285
R7968 Transmission_Gate_Layout_4.VIN.n17 Transmission_Gate_Layout_4.VIN.n16 0.7285
R7969 Transmission_Gate_Layout_4.VIN.n19 Transmission_Gate_Layout_4.VIN.t55 0.7285
R7970 Transmission_Gate_Layout_4.VIN.n19 Transmission_Gate_Layout_4.VIN.n18 0.7285
R7971 Transmission_Gate_Layout_4.VIN.n21 Transmission_Gate_Layout_4.VIN.t9 0.7285
R7972 Transmission_Gate_Layout_4.VIN.n21 Transmission_Gate_Layout_4.VIN.n20 0.7285
R7973 Transmission_Gate_Layout_4.VIN.n89 Transmission_Gate_Layout_4.VIN.t17 0.7285
R7974 Transmission_Gate_Layout_4.VIN.n89 Transmission_Gate_Layout_4.VIN.n88 0.7285
R7975 Transmission_Gate_Layout_4.VIN.n91 Transmission_Gate_Layout_4.VIN.t66 0.7285
R7976 Transmission_Gate_Layout_4.VIN.n91 Transmission_Gate_Layout_4.VIN.n90 0.7285
R7977 Transmission_Gate_Layout_4.VIN.n93 Transmission_Gate_Layout_4.VIN.t56 0.7285
R7978 Transmission_Gate_Layout_4.VIN.n93 Transmission_Gate_Layout_4.VIN.n92 0.7285
R7979 Transmission_Gate_Layout_4.VIN.n9 Transmission_Gate_Layout_4.VIN.t64 0.7285
R7980 Transmission_Gate_Layout_4.VIN.n9 Transmission_Gate_Layout_4.VIN.n8 0.7285
R7981 Transmission_Gate_Layout_4.VIN.n11 Transmission_Gate_Layout_4.VIN.t60 0.7285
R7982 Transmission_Gate_Layout_4.VIN.n11 Transmission_Gate_Layout_4.VIN.n10 0.7285
R7983 Transmission_Gate_Layout_4.VIN.n13 Transmission_Gate_Layout_4.VIN.t18 0.7285
R7984 Transmission_Gate_Layout_4.VIN.n13 Transmission_Gate_Layout_4.VIN.n12 0.7285
R7985 Transmission_Gate_Layout_4.VIN.n58 Transmission_Gate_Layout_4.VIN.n57 0.626587
R7986 Transmission_Gate_Layout_4.VIN.n68 Transmission_Gate_Layout_4.VIN.n67 0.626587
R7987 Transmission_Gate_Layout_4.VIN.n142 Transmission_Gate_Layout_4.VIN.n133 0.626587
R7988 Transmission_Gate_Layout_4.VIN.n81 Transmission_Gate_Layout_4.VIN 0.607022
R7989 Transmission_Gate_Layout_4.VIN.n86 Transmission_Gate_Layout_4.VIN.n79 0.575717
R7990 Transmission_Gate_Layout_4.VIN.n67 Transmission_Gate_Layout_4.VIN.n66 0.575717
R7991 Transmission_Gate_Layout_4.VIN.n68 Transmission_Gate_Layout_4.VIN.n23 0.575717
R7992 Transmission_Gate_Layout_4.VIN.n97 Transmission_Gate_Layout_4.VIN.n15 0.575717
R7993 Transmission_Gate_Layout_4.VIN.n97 Transmission_Gate_Layout_4.VIN.n96 0.570002
R7994 Transmission_Gate_Layout_4.VIN.n96 Transmission_Gate_Layout_4.VIN.n95 0.562022
R7995 Transmission_Gate_Layout_4.VIN.n133 Transmission_Gate_Layout_4.VIN.n132 0.428978
R7996 Transmission_Gate_Layout_4.VIN.n142 Transmission_Gate_Layout_4.VIN.n141 0.428978
R7997 Transmission_Gate_Layout_4.VIN.n129 Transmission_Gate_Layout_4.VIN.n120 0.331152
R7998 Transmission_Gate_Layout_4.VIN.n58 Transmission_Gate_Layout_4.VIN.n31 0.331152
R7999 Transmission_Gate_Layout_4.VIN.n57 Transmission_Gate_Layout_4.VIN.n39 0.331152
R8000 Transmission_Gate_Layout_4.VIN.n53 Transmission_Gate_Layout_4.VIN.n47 0.331152
R8001 Transmission_Gate_Layout_4.VIN.n67 Transmission_Gate_Layout_4.VIN.n58 0.239196
R8002 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.VIN.n142 0.192239
R8003 Transmission_Gate_Layout_18.CLKB.n24 Transmission_Gate_Layout_18.CLKB.t29 54.5477
R8004 Transmission_Gate_Layout_18.CLKB.n29 Transmission_Gate_Layout_18.CLKB.t24 38.3255
R8005 Transmission_Gate_Layout_18.CLKB.n27 Transmission_Gate_Layout_18.CLKB.t12 38.3255
R8006 Transmission_Gate_Layout_18.CLKB.n26 Transmission_Gate_Layout_18.CLKB.t14 38.3255
R8007 Transmission_Gate_Layout_18.CLKB.n25 Transmission_Gate_Layout_18.CLKB.t20 38.3255
R8008 Transmission_Gate_Layout_18.CLKB.n24 Transmission_Gate_Layout_18.CLKB.t22 38.3255
R8009 Transmission_Gate_Layout_18.CLKB.n28 Transmission_Gate_Layout_18.CLKB.t6 38.3255
R8010 Transmission_Gate_Layout_18.CLKB.t17 Transmission_Gate_Layout_18.CLKB.n2 37.9344
R8011 Transmission_Gate_Layout_18.CLKB.t23 Transmission_Gate_Layout_18.CLKB.n5 37.9344
R8012 Transmission_Gate_Layout_18.CLKB.t7 Transmission_Gate_Layout_18.CLKB.n8 37.9344
R8013 Transmission_Gate_Layout_18.CLKB.t8 Transmission_Gate_Layout_18.CLKB.n11 37.9344
R8014 Transmission_Gate_Layout_18.CLKB.t13 Transmission_Gate_Layout_18.CLKB.n14 37.9344
R8015 Transmission_Gate_Layout_18.CLKB.t15 Transmission_Gate_Layout_18.CLKB.n17 37.9344
R8016 Transmission_Gate_Layout_18.CLKB.t21 Transmission_Gate_Layout_18.CLKB.n20 37.9344
R8017 Transmission_Gate_Layout_18.CLKB.t28 Transmission_Gate_Layout_18.CLKB.n21 37.9344
R8018 Transmission_Gate_Layout_18.CLKB.n3 Transmission_Gate_Layout_18.CLKB.t17 37.5434
R8019 Transmission_Gate_Layout_18.CLKB.n6 Transmission_Gate_Layout_18.CLKB.t23 37.5434
R8020 Transmission_Gate_Layout_18.CLKB.n9 Transmission_Gate_Layout_18.CLKB.t7 37.5434
R8021 Transmission_Gate_Layout_18.CLKB.n12 Transmission_Gate_Layout_18.CLKB.t8 37.5434
R8022 Transmission_Gate_Layout_18.CLKB.n15 Transmission_Gate_Layout_18.CLKB.t13 37.5434
R8023 Transmission_Gate_Layout_18.CLKB.n18 Transmission_Gate_Layout_18.CLKB.t15 37.5434
R8024 Transmission_Gate_Layout_18.CLKB.n23 Transmission_Gate_Layout_18.CLKB.t21 37.5434
R8025 Transmission_Gate_Layout_18.CLKB.n22 Transmission_Gate_Layout_18.CLKB.t28 37.5434
R8026 Transmission_Gate_Layout_18.CLKB.t24 Transmission_Gate_Layout_18.CLKB.n3 37.413
R8027 Transmission_Gate_Layout_18.CLKB.t12 Transmission_Gate_Layout_18.CLKB.n9 37.413
R8028 Transmission_Gate_Layout_18.CLKB.t14 Transmission_Gate_Layout_18.CLKB.n12 37.413
R8029 Transmission_Gate_Layout_18.CLKB.t20 Transmission_Gate_Layout_18.CLKB.n15 37.413
R8030 Transmission_Gate_Layout_18.CLKB.t22 Transmission_Gate_Layout_18.CLKB.n18 37.413
R8031 Transmission_Gate_Layout_18.CLKB.t29 Transmission_Gate_Layout_18.CLKB.n23 37.413
R8032 Transmission_Gate_Layout_18.CLKB.n22 Transmission_Gate_Layout_18.CLKB.t11 37.413
R8033 Transmission_Gate_Layout_18.CLKB.t6 Transmission_Gate_Layout_18.CLKB.n6 37.413
R8034 Transmission_Gate_Layout_18.CLKB.n2 Transmission_Gate_Layout_18.CLKB.t27 37.0219
R8035 Transmission_Gate_Layout_18.CLKB.n5 Transmission_Gate_Layout_18.CLKB.t10 37.0219
R8036 Transmission_Gate_Layout_18.CLKB.n8 Transmission_Gate_Layout_18.CLKB.t18 37.0219
R8037 Transmission_Gate_Layout_18.CLKB.n11 Transmission_Gate_Layout_18.CLKB.t19 37.0219
R8038 Transmission_Gate_Layout_18.CLKB.n14 Transmission_Gate_Layout_18.CLKB.t25 37.0219
R8039 Transmission_Gate_Layout_18.CLKB.n17 Transmission_Gate_Layout_18.CLKB.t26 37.0219
R8040 Transmission_Gate_Layout_18.CLKB.n21 Transmission_Gate_Layout_18.CLKB.t16 37.0219
R8041 Transmission_Gate_Layout_18.CLKB.n20 Transmission_Gate_Layout_18.CLKB.t9 37.0219
R8042 Transmission_Gate_Layout_18.CLKB.t10 Transmission_Gate_Layout_18.CLKB.n4 35.1969
R8043 Transmission_Gate_Layout_18.CLKB.t18 Transmission_Gate_Layout_18.CLKB.n7 35.1969
R8044 Transmission_Gate_Layout_18.CLKB.t19 Transmission_Gate_Layout_18.CLKB.n10 35.1969
R8045 Transmission_Gate_Layout_18.CLKB.t25 Transmission_Gate_Layout_18.CLKB.n13 35.1969
R8046 Transmission_Gate_Layout_18.CLKB.t26 Transmission_Gate_Layout_18.CLKB.n16 35.1969
R8047 Transmission_Gate_Layout_18.CLKB.t9 Transmission_Gate_Layout_18.CLKB.n19 35.1969
R8048 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_18.CLKB.n29 26.6826
R8049 Transmission_Gate_Layout_18.CLKB.n23 Transmission_Gate_Layout_18.CLKB.n22 19.148
R8050 Transmission_Gate_Layout_18.CLKB.n29 Transmission_Gate_Layout_18.CLKB.n28 16.2227
R8051 Transmission_Gate_Layout_18.CLKB.n28 Transmission_Gate_Layout_18.CLKB.n27 16.2227
R8052 Transmission_Gate_Layout_18.CLKB.n27 Transmission_Gate_Layout_18.CLKB.n26 16.2227
R8053 Transmission_Gate_Layout_18.CLKB.n26 Transmission_Gate_Layout_18.CLKB.n25 16.2227
R8054 Transmission_Gate_Layout_18.CLKB.n25 Transmission_Gate_Layout_18.CLKB.n24 16.2227
R8055 Transmission_Gate_Layout_18.CLKB.n0 Transmission_Gate_Layout_18.CLKB.t4 5.21612
R8056 Transmission_Gate_Layout_18.CLKB.n30 Transmission_Gate_Layout_18.CLKB.t0 4.57285
R8057 Transmission_Gate_Layout_18.CLKB.n0 Transmission_Gate_Layout_18.CLKB.t3 4.4609
R8058 Transmission_Gate_Layout_18.CLKB.n1 Transmission_Gate_Layout_18.CLKB.t5 4.4609
R8059 Transmission_Gate_Layout_18.CLKB.n31 Transmission_Gate_Layout_18.CLKB.t1 3.3285
R8060 Transmission_Gate_Layout_18.CLKB.n30 Transmission_Gate_Layout_18.CLKB.t2 3.3285
R8061 Transmission_Gate_Layout_18.CLKB.n31 Transmission_Gate_Layout_18.CLKB.n30 1.24485
R8062 Transmission_Gate_Layout_18.CLKB.n1 Transmission_Gate_Layout_18.CLKB.n0 0.755717
R8063 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_18.CLKB.n31 0.750969
R8064 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_18.CLKB.n1 0.510317
R8065 IN2.n58 IN2 21.2759
R8066 IN2.n4 IN2.n1 3.90572
R8067 IN2.n48 IN2.n47 3.90572
R8068 IN2.n56 IN2.n55 3.90572
R8069 IN2.n34 IN2.n31 3.84485
R8070 IN2.n26 IN2.n23 3.84485
R8071 IN2.n14 IN2.n13 3.84485
R8072 IN2.n7 IN2.n6 3.1505
R8073 IN2.n4 IN2.n3 3.1505
R8074 IN2.n62 IN2.n61 3.1505
R8075 IN2.n65 IN2.n64 3.1505
R8076 IN2.n68 IN2.n67 3.1505
R8077 IN2.n48 IN2.n45 3.1505
R8078 IN2.n49 IN2.n43 3.1505
R8079 IN2.n56 IN2.n53 3.1505
R8080 IN2.n57 IN2.n51 3.1505
R8081 IN2.n34 IN2.n33 2.6005
R8082 IN2.n37 IN2.n36 2.6005
R8083 IN2.n26 IN2.n25 2.6005
R8084 IN2.n29 IN2.n28 2.6005
R8085 IN2.n39 IN2.n21 2.6005
R8086 IN2.n40 IN2.n19 2.6005
R8087 IN2.n41 IN2.n17 2.6005
R8088 IN2.n14 IN2.n11 2.6005
R8089 IN2.n15 IN2.n9 2.6005
R8090 IN2.n67 IN2.t30 1.3109
R8091 IN2.n67 IN2.n66 1.3109
R8092 IN2.n64 IN2.t35 1.3109
R8093 IN2.n64 IN2.n63 1.3109
R8094 IN2.n61 IN2.t41 1.3109
R8095 IN2.n61 IN2.n60 1.3109
R8096 IN2.n1 IN2.t33 1.3109
R8097 IN2.n1 IN2.n0 1.3109
R8098 IN2.n3 IN2.t28 1.3109
R8099 IN2.n3 IN2.n2 1.3109
R8100 IN2.n6 IN2.t46 1.3109
R8101 IN2.n6 IN2.n5 1.3109
R8102 IN2.n43 IN2.t24 1.3109
R8103 IN2.n43 IN2.n42 1.3109
R8104 IN2.n45 IN2.t43 1.3109
R8105 IN2.n45 IN2.n44 1.3109
R8106 IN2.n47 IN2.t37 1.3109
R8107 IN2.n47 IN2.n46 1.3109
R8108 IN2.n51 IN2.t39 1.3109
R8109 IN2.n51 IN2.n50 1.3109
R8110 IN2.n53 IN2.t32 1.3109
R8111 IN2.n53 IN2.n52 1.3109
R8112 IN2.n55 IN2.t26 1.3109
R8113 IN2.n55 IN2.n54 1.3109
R8114 IN2.n37 IN2.n34 1.24485
R8115 IN2.n29 IN2.n26 1.24485
R8116 IN2.n41 IN2.n40 1.24485
R8117 IN2.n40 IN2.n39 1.24485
R8118 IN2.n15 IN2.n14 1.24485
R8119 IN2.n38 IN2.n37 1.2018
R8120 IN2.n39 IN2.n38 1.2018
R8121 IN2.n62 IN2.n59 0.957239
R8122 IN2.n69 IN2.n41 0.806587
R8123 IN2.n70 IN2.n15 0.806587
R8124 IN2.n7 IN2.n4 0.755717
R8125 IN2.n65 IN2.n62 0.755717
R8126 IN2.n68 IN2.n65 0.755717
R8127 IN2.n49 IN2.n48 0.755717
R8128 IN2.n57 IN2.n56 0.755717
R8129 IN2.n17 IN2.t9 0.7285
R8130 IN2.n17 IN2.n16 0.7285
R8131 IN2.n19 IN2.t16 0.7285
R8132 IN2.n19 IN2.n18 0.7285
R8133 IN2.n21 IN2.t4 0.7285
R8134 IN2.n21 IN2.n20 0.7285
R8135 IN2.n36 IN2.t2 0.7285
R8136 IN2.n36 IN2.n35 0.7285
R8137 IN2.n33 IN2.t12 0.7285
R8138 IN2.n33 IN2.n32 0.7285
R8139 IN2.n31 IN2.t5 0.7285
R8140 IN2.n31 IN2.n30 0.7285
R8141 IN2.n28 IN2.t11 0.7285
R8142 IN2.n28 IN2.n27 0.7285
R8143 IN2.n25 IN2.t22 0.7285
R8144 IN2.n25 IN2.n24 0.7285
R8145 IN2.n23 IN2.t17 0.7285
R8146 IN2.n23 IN2.n22 0.7285
R8147 IN2.n9 IN2.t0 0.7285
R8148 IN2.n9 IN2.n8 0.7285
R8149 IN2.n11 IN2.t8 0.7285
R8150 IN2.n11 IN2.n10 0.7285
R8151 IN2.n13 IN2.t20 0.7285
R8152 IN2.n13 IN2.n12 0.7285
R8153 IN2.n70 IN2.n69 0.626587
R8154 IN2.n38 IN2.n29 0.575717
R8155 IN2.n59 IN2.n58 0.570002
R8156 IN2.n70 IN2.n7 0.428978
R8157 IN2.n69 IN2.n68 0.428978
R8158 IN2.n59 IN2.n49 0.331152
R8159 IN2.n58 IN2.n57 0.317457
R8160 IN2 IN2.n70 0.192239
R8161 Transmission_Gate_Layout_8.CLKB.n24 Transmission_Gate_Layout_8.CLKB.t21 54.5477
R8162 Transmission_Gate_Layout_8.CLKB.n29 Transmission_Gate_Layout_8.CLKB.t19 38.3255
R8163 Transmission_Gate_Layout_8.CLKB.n27 Transmission_Gate_Layout_8.CLKB.t13 38.3255
R8164 Transmission_Gate_Layout_8.CLKB.n26 Transmission_Gate_Layout_8.CLKB.t18 38.3255
R8165 Transmission_Gate_Layout_8.CLKB.n25 Transmission_Gate_Layout_8.CLKB.t8 38.3255
R8166 Transmission_Gate_Layout_8.CLKB.n24 Transmission_Gate_Layout_8.CLKB.t15 38.3255
R8167 Transmission_Gate_Layout_8.CLKB.n28 Transmission_Gate_Layout_8.CLKB.t24 38.3255
R8168 Transmission_Gate_Layout_8.CLKB.t27 Transmission_Gate_Layout_8.CLKB.n2 37.9344
R8169 Transmission_Gate_Layout_8.CLKB.t6 Transmission_Gate_Layout_8.CLKB.n5 37.9344
R8170 Transmission_Gate_Layout_8.CLKB.t20 Transmission_Gate_Layout_8.CLKB.n8 37.9344
R8171 Transmission_Gate_Layout_8.CLKB.t25 Transmission_Gate_Layout_8.CLKB.n11 37.9344
R8172 Transmission_Gate_Layout_8.CLKB.t14 Transmission_Gate_Layout_8.CLKB.n14 37.9344
R8173 Transmission_Gate_Layout_8.CLKB.t22 Transmission_Gate_Layout_8.CLKB.n17 37.9344
R8174 Transmission_Gate_Layout_8.CLKB.t28 Transmission_Gate_Layout_8.CLKB.n20 37.9344
R8175 Transmission_Gate_Layout_8.CLKB.t17 Transmission_Gate_Layout_8.CLKB.n21 37.9344
R8176 Transmission_Gate_Layout_8.CLKB.n3 Transmission_Gate_Layout_8.CLKB.t27 37.5434
R8177 Transmission_Gate_Layout_8.CLKB.n6 Transmission_Gate_Layout_8.CLKB.t6 37.5434
R8178 Transmission_Gate_Layout_8.CLKB.n9 Transmission_Gate_Layout_8.CLKB.t20 37.5434
R8179 Transmission_Gate_Layout_8.CLKB.n12 Transmission_Gate_Layout_8.CLKB.t25 37.5434
R8180 Transmission_Gate_Layout_8.CLKB.n15 Transmission_Gate_Layout_8.CLKB.t14 37.5434
R8181 Transmission_Gate_Layout_8.CLKB.n18 Transmission_Gate_Layout_8.CLKB.t22 37.5434
R8182 Transmission_Gate_Layout_8.CLKB.n23 Transmission_Gate_Layout_8.CLKB.t28 37.5434
R8183 Transmission_Gate_Layout_8.CLKB.n22 Transmission_Gate_Layout_8.CLKB.t17 37.5434
R8184 Transmission_Gate_Layout_8.CLKB.t19 Transmission_Gate_Layout_8.CLKB.n3 37.413
R8185 Transmission_Gate_Layout_8.CLKB.t13 Transmission_Gate_Layout_8.CLKB.n9 37.413
R8186 Transmission_Gate_Layout_8.CLKB.t18 Transmission_Gate_Layout_8.CLKB.n12 37.413
R8187 Transmission_Gate_Layout_8.CLKB.t8 Transmission_Gate_Layout_8.CLKB.n15 37.413
R8188 Transmission_Gate_Layout_8.CLKB.t15 Transmission_Gate_Layout_8.CLKB.n18 37.413
R8189 Transmission_Gate_Layout_8.CLKB.t21 Transmission_Gate_Layout_8.CLKB.n23 37.413
R8190 Transmission_Gate_Layout_8.CLKB.n22 Transmission_Gate_Layout_8.CLKB.t9 37.413
R8191 Transmission_Gate_Layout_8.CLKB.t24 Transmission_Gate_Layout_8.CLKB.n6 37.413
R8192 Transmission_Gate_Layout_8.CLKB.n2 Transmission_Gate_Layout_8.CLKB.t11 37.0219
R8193 Transmission_Gate_Layout_8.CLKB.n5 Transmission_Gate_Layout_8.CLKB.t16 37.0219
R8194 Transmission_Gate_Layout_8.CLKB.n8 Transmission_Gate_Layout_8.CLKB.t29 37.0219
R8195 Transmission_Gate_Layout_8.CLKB.n11 Transmission_Gate_Layout_8.CLKB.t10 37.0219
R8196 Transmission_Gate_Layout_8.CLKB.n14 Transmission_Gate_Layout_8.CLKB.t23 37.0219
R8197 Transmission_Gate_Layout_8.CLKB.n17 Transmission_Gate_Layout_8.CLKB.t7 37.0219
R8198 Transmission_Gate_Layout_8.CLKB.n21 Transmission_Gate_Layout_8.CLKB.t26 37.0219
R8199 Transmission_Gate_Layout_8.CLKB.n20 Transmission_Gate_Layout_8.CLKB.t12 37.0219
R8200 Transmission_Gate_Layout_8.CLKB.t16 Transmission_Gate_Layout_8.CLKB.n4 35.1969
R8201 Transmission_Gate_Layout_8.CLKB.t29 Transmission_Gate_Layout_8.CLKB.n7 35.1969
R8202 Transmission_Gate_Layout_8.CLKB.t10 Transmission_Gate_Layout_8.CLKB.n10 35.1969
R8203 Transmission_Gate_Layout_8.CLKB.t23 Transmission_Gate_Layout_8.CLKB.n13 35.1969
R8204 Transmission_Gate_Layout_8.CLKB.t7 Transmission_Gate_Layout_8.CLKB.n16 35.1969
R8205 Transmission_Gate_Layout_8.CLKB.t12 Transmission_Gate_Layout_8.CLKB.n19 35.1969
R8206 Transmission_Gate_Layout_8.CLKB Transmission_Gate_Layout_8.CLKB.n29 26.6826
R8207 Transmission_Gate_Layout_8.CLKB.n23 Transmission_Gate_Layout_8.CLKB.n22 19.148
R8208 Transmission_Gate_Layout_8.CLKB.n29 Transmission_Gate_Layout_8.CLKB.n28 16.2227
R8209 Transmission_Gate_Layout_8.CLKB.n28 Transmission_Gate_Layout_8.CLKB.n27 16.2227
R8210 Transmission_Gate_Layout_8.CLKB.n27 Transmission_Gate_Layout_8.CLKB.n26 16.2227
R8211 Transmission_Gate_Layout_8.CLKB.n26 Transmission_Gate_Layout_8.CLKB.n25 16.2227
R8212 Transmission_Gate_Layout_8.CLKB.n25 Transmission_Gate_Layout_8.CLKB.n24 16.2227
R8213 Transmission_Gate_Layout_8.CLKB.n0 Transmission_Gate_Layout_8.CLKB.t3 5.21612
R8214 Transmission_Gate_Layout_8.CLKB.n30 Transmission_Gate_Layout_8.CLKB.t0 4.57285
R8215 Transmission_Gate_Layout_8.CLKB.n0 Transmission_Gate_Layout_8.CLKB.t5 4.4609
R8216 Transmission_Gate_Layout_8.CLKB.n1 Transmission_Gate_Layout_8.CLKB.t4 4.4609
R8217 Transmission_Gate_Layout_8.CLKB.n30 Transmission_Gate_Layout_8.CLKB.t1 3.3285
R8218 Transmission_Gate_Layout_8.CLKB.n31 Transmission_Gate_Layout_8.CLKB.t2 3.3285
R8219 Transmission_Gate_Layout_8.CLKB.n31 Transmission_Gate_Layout_8.CLKB.n30 1.24485
R8220 Transmission_Gate_Layout_8.CLKB.n1 Transmission_Gate_Layout_8.CLKB.n0 0.755717
R8221 Transmission_Gate_Layout_8.CLKB Transmission_Gate_Layout_8.CLKB.n31 0.750969
R8222 Transmission_Gate_Layout_8.CLKB Transmission_Gate_Layout_8.CLKB.n1 0.510317
R8223 Transmission_Gate_Layout_12.CLK.t18 Transmission_Gate_Layout_12.CLK.t14 82.9076
R8224 Transmission_Gate_Layout_12.CLK.t3 Transmission_Gate_Layout_12.CLK.t18 82.9076
R8225 Transmission_Gate_Layout_12.CLK.n27 Transmission_Gate_Layout_12.CLK.t3 49.7969
R8226 Transmission_Gate_Layout_12.CLK.n26 Transmission_Gate_Layout_12.CLK.n25 35.0405
R8227 Transmission_Gate_Layout_12.CLK.n27 Transmission_Gate_Layout_12.CLK.t16 31.1559
R8228 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_12.CLK.n1 24.3453
R8229 Transmission_Gate_Layout_12.CLK.n0 Transmission_Gate_Layout_12.CLK.t28 22.0309
R8230 Transmission_Gate_Layout_12.CLK.t5 Transmission_Gate_Layout_12.CLK.n2 21.9005
R8231 Transmission_Gate_Layout_12.CLK.t32 Transmission_Gate_Layout_12.CLK.n17 21.9005
R8232 Transmission_Gate_Layout_12.CLK.n26 Transmission_Gate_Layout_12.CLK.t5 21.5094
R8233 Transmission_Gate_Layout_12.CLK.n25 Transmission_Gate_Layout_12.CLK.t32 21.5094
R8234 Transmission_Gate_Layout_12.CLK.n24 Transmission_Gate_Layout_12.CLK.t24 21.5094
R8235 Transmission_Gate_Layout_12.CLK.n23 Transmission_Gate_Layout_12.CLK.t7 21.5094
R8236 Transmission_Gate_Layout_12.CLK.n22 Transmission_Gate_Layout_12.CLK.t33 21.5094
R8237 Transmission_Gate_Layout_12.CLK.n21 Transmission_Gate_Layout_12.CLK.t25 21.5094
R8238 Transmission_Gate_Layout_12.CLK.n20 Transmission_Gate_Layout_12.CLK.t8 21.5094
R8239 Transmission_Gate_Layout_12.CLK.n19 Transmission_Gate_Layout_12.CLK.t31 21.5094
R8240 Transmission_Gate_Layout_12.CLK.n18 Transmission_Gate_Layout_12.CLK.t11 21.5094
R8241 Transmission_Gate_Layout_12.CLK.n0 Transmission_Gate_Layout_12.CLK.t27 21.3791
R8242 Transmission_Gate_Layout_12.CLK.n1 Transmission_Gate_Layout_12.CLK.t12 21.3791
R8243 Transmission_Gate_Layout_12.CLK.n25 Transmission_Gate_Layout_12.CLK.t9 20.988
R8244 Transmission_Gate_Layout_12.CLK.n24 Transmission_Gate_Layout_12.CLK.t2 20.988
R8245 Transmission_Gate_Layout_12.CLK.n23 Transmission_Gate_Layout_12.CLK.t17 20.988
R8246 Transmission_Gate_Layout_12.CLK.n22 Transmission_Gate_Layout_12.CLK.t10 20.988
R8247 Transmission_Gate_Layout_12.CLK.n21 Transmission_Gate_Layout_12.CLK.t4 20.988
R8248 Transmission_Gate_Layout_12.CLK.n20 Transmission_Gate_Layout_12.CLK.t19 20.988
R8249 Transmission_Gate_Layout_12.CLK.n19 Transmission_Gate_Layout_12.CLK.t6 20.988
R8250 Transmission_Gate_Layout_12.CLK.n18 Transmission_Gate_Layout_12.CLK.t22 20.988
R8251 Transmission_Gate_Layout_12.CLK.t16 Transmission_Gate_Layout_12.CLK.n26 20.988
R8252 Transmission_Gate_Layout_12.CLK.n1 Transmission_Gate_Layout_12.CLK.n0 20.8576
R8253 Transmission_Gate_Layout_12.CLK.n2 Transmission_Gate_Layout_12.CLK.t26 20.5969
R8254 Transmission_Gate_Layout_12.CLK.n17 Transmission_Gate_Layout_12.CLK.t21 20.5969
R8255 Transmission_Gate_Layout_12.CLK.n16 Transmission_Gate_Layout_12.CLK.t13 20.5969
R8256 Transmission_Gate_Layout_12.CLK.n15 Transmission_Gate_Layout_12.CLK.t29 20.5969
R8257 Transmission_Gate_Layout_12.CLK.n14 Transmission_Gate_Layout_12.CLK.t23 20.5969
R8258 Transmission_Gate_Layout_12.CLK.n13 Transmission_Gate_Layout_12.CLK.t15 20.5969
R8259 Transmission_Gate_Layout_12.CLK.n12 Transmission_Gate_Layout_12.CLK.t30 20.5969
R8260 Transmission_Gate_Layout_12.CLK.n10 Transmission_Gate_Layout_12.CLK.t34 20.5969
R8261 Transmission_Gate_Layout_12.CLK.n11 Transmission_Gate_Layout_12.CLK.t20 20.5969
R8262 Transmission_Gate_Layout_12.CLK.n17 Transmission_Gate_Layout_12.CLK.n16 19.4672
R8263 Transmission_Gate_Layout_12.CLK.n16 Transmission_Gate_Layout_12.CLK.n15 19.4672
R8264 Transmission_Gate_Layout_12.CLK.n15 Transmission_Gate_Layout_12.CLK.n14 19.4672
R8265 Transmission_Gate_Layout_12.CLK.n14 Transmission_Gate_Layout_12.CLK.n13 19.4672
R8266 Transmission_Gate_Layout_12.CLK.n13 Transmission_Gate_Layout_12.CLK.n12 19.4672
R8267 Transmission_Gate_Layout_12.CLK.n12 Transmission_Gate_Layout_12.CLK.n11 19.4672
R8268 Transmission_Gate_Layout_12.CLK.n11 Transmission_Gate_Layout_12.CLK.n10 19.4672
R8269 Transmission_Gate_Layout_12.CLK.n25 Transmission_Gate_Layout_12.CLK.n24 19.4672
R8270 Transmission_Gate_Layout_12.CLK.n24 Transmission_Gate_Layout_12.CLK.n23 19.4672
R8271 Transmission_Gate_Layout_12.CLK.n23 Transmission_Gate_Layout_12.CLK.n22 19.4672
R8272 Transmission_Gate_Layout_12.CLK.n22 Transmission_Gate_Layout_12.CLK.n21 19.4672
R8273 Transmission_Gate_Layout_12.CLK.n21 Transmission_Gate_Layout_12.CLK.n20 19.4672
R8274 Transmission_Gate_Layout_12.CLK.n20 Transmission_Gate_Layout_12.CLK.n19 19.4672
R8275 Transmission_Gate_Layout_12.CLK.n19 Transmission_Gate_Layout_12.CLK.n18 19.4672
R8276 Transmission_Gate_Layout_12.CLK.t21 Transmission_Gate_Layout_12.CLK.n3 18.9023
R8277 Transmission_Gate_Layout_12.CLK.t13 Transmission_Gate_Layout_12.CLK.n4 18.9023
R8278 Transmission_Gate_Layout_12.CLK.t29 Transmission_Gate_Layout_12.CLK.n5 18.9023
R8279 Transmission_Gate_Layout_12.CLK.t23 Transmission_Gate_Layout_12.CLK.n6 18.9023
R8280 Transmission_Gate_Layout_12.CLK.t15 Transmission_Gate_Layout_12.CLK.n7 18.9023
R8281 Transmission_Gate_Layout_12.CLK.t30 Transmission_Gate_Layout_12.CLK.n8 18.9023
R8282 Transmission_Gate_Layout_12.CLK.t20 Transmission_Gate_Layout_12.CLK.n9 18.9023
R8283 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_12.CLK.n27 16.443
R8284 Transmission_Gate_Layout_12.CLK.n28 Transmission_Gate_Layout_12.CLK 8.76208
R8285 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_12.CLK.n29 7.70137
R8286 Transmission_Gate_Layout_12.CLK.n28 Transmission_Gate_Layout_12.CLK 5.55127
R8287 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_12.CLK.n30 4.70224
R8288 Transmission_Gate_Layout_12.CLK.n31 Transmission_Gate_Layout_12.CLK.n28 3.54376
R8289 Transmission_Gate_Layout_12.CLK.n31 Transmission_Gate_Layout_12.CLK 0.608978
R8290 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_12.CLK.n31 0.248978
R8291 IN4.n65 IN4 7.16364
R8292 IN4.n30 IN4.n29 3.90572
R8293 IN4.n22 IN4.n21 3.90572
R8294 IN4.n4 IN4.n1 3.90572
R8295 IN4.n52 IN4.n49 3.84485
R8296 IN4.n60 IN4.n57 3.84485
R8297 IN4.n14 IN4.n13 3.84485
R8298 IN4.n30 IN4.n27 3.1505
R8299 IN4.n31 IN4.n25 3.1505
R8300 IN4.n22 IN4.n19 3.1505
R8301 IN4.n23 IN4.n17 3.1505
R8302 IN4.n41 IN4.n40 3.1505
R8303 IN4.n38 IN4.n37 3.1505
R8304 IN4.n35 IN4.n34 3.1505
R8305 IN4.n4 IN4.n3 3.1505
R8306 IN4.n7 IN4.n6 3.1505
R8307 IN4.n52 IN4.n51 2.6005
R8308 IN4.n55 IN4.n54 2.6005
R8309 IN4.n60 IN4.n59 2.6005
R8310 IN4.n63 IN4.n62 2.6005
R8311 IN4.n14 IN4.n11 2.6005
R8312 IN4.n15 IN4.n9 2.6005
R8313 IN4.n66 IN4.n47 2.6005
R8314 IN4.n67 IN4.n45 2.6005
R8315 IN4.n68 IN4.n43 2.6005
R8316 IN4.n34 IN4.t31 1.3109
R8317 IN4.n34 IN4.n33 1.3109
R8318 IN4.n37 IN4.t25 1.3109
R8319 IN4.n37 IN4.n36 1.3109
R8320 IN4.n40 IN4.t44 1.3109
R8321 IN4.n40 IN4.n39 1.3109
R8322 IN4.n25 IN4.t45 1.3109
R8323 IN4.n25 IN4.n24 1.3109
R8324 IN4.n27 IN4.t38 1.3109
R8325 IN4.n27 IN4.n26 1.3109
R8326 IN4.n29 IN4.t30 1.3109
R8327 IN4.n29 IN4.n28 1.3109
R8328 IN4.n17 IN4.t47 1.3109
R8329 IN4.n17 IN4.n16 1.3109
R8330 IN4.n19 IN4.t41 1.3109
R8331 IN4.n19 IN4.n18 1.3109
R8332 IN4.n21 IN4.t35 1.3109
R8333 IN4.n21 IN4.n20 1.3109
R8334 IN4.n6 IN4.t27 1.3109
R8335 IN4.n6 IN4.n5 1.3109
R8336 IN4.n3 IN4.t33 1.3109
R8337 IN4.n3 IN4.n2 1.3109
R8338 IN4.n1 IN4.t39 1.3109
R8339 IN4.n1 IN4.n0 1.3109
R8340 IN4.n55 IN4.n52 1.24485
R8341 IN4.n63 IN4.n60 1.24485
R8342 IN4.n15 IN4.n14 1.24485
R8343 IN4.n68 IN4.n67 1.24485
R8344 IN4.n67 IN4.n66 1.24485
R8345 IN4.n64 IN4.n63 1.2018
R8346 IN4.n32 IN4.n31 0.957239
R8347 IN4.n35 IN4.n32 0.957239
R8348 IN4.n70 IN4.n15 0.806587
R8349 IN4.n69 IN4.n68 0.806587
R8350 IN4.n31 IN4.n30 0.755717
R8351 IN4.n23 IN4.n22 0.755717
R8352 IN4.n38 IN4.n35 0.755717
R8353 IN4.n41 IN4.n38 0.755717
R8354 IN4.n7 IN4.n4 0.755717
R8355 IN4.n54 IN4.t11 0.7285
R8356 IN4.n54 IN4.n53 0.7285
R8357 IN4.n51 IN4.t1 0.7285
R8358 IN4.n51 IN4.n50 0.7285
R8359 IN4.n49 IN4.t8 0.7285
R8360 IN4.n49 IN4.n48 0.7285
R8361 IN4.n62 IN4.t18 0.7285
R8362 IN4.n62 IN4.n61 0.7285
R8363 IN4.n59 IN4.t4 0.7285
R8364 IN4.n59 IN4.n58 0.7285
R8365 IN4.n57 IN4.t12 0.7285
R8366 IN4.n57 IN4.n56 0.7285
R8367 IN4.n43 IN4.t0 0.7285
R8368 IN4.n43 IN4.n42 0.7285
R8369 IN4.n45 IN4.t17 0.7285
R8370 IN4.n45 IN4.n44 0.7285
R8371 IN4.n47 IN4.t3 0.7285
R8372 IN4.n47 IN4.n46 0.7285
R8373 IN4.n9 IN4.t16 0.7285
R8374 IN4.n9 IN4.n8 0.7285
R8375 IN4.n11 IN4.t9 0.7285
R8376 IN4.n11 IN4.n10 0.7285
R8377 IN4.n13 IN4.t21 0.7285
R8378 IN4.n13 IN4.n12 0.7285
R8379 IN4.n70 IN4.n69 0.626587
R8380 IN4.n64 IN4.n55 0.575717
R8381 IN4.n65 IN4.n64 0.570002
R8382 IN4.n66 IN4.n65 0.562022
R8383 IN4.n69 IN4.n41 0.428978
R8384 IN4.n70 IN4.n7 0.428978
R8385 IN4.n32 IN4.n23 0.331152
R8386 IN4 IN4.n70 0.192239
R8387 Transmission_Gate_Layout_3.CLK.t64 Transmission_Gate_Layout_3.CLK.t59 82.9076
R8388 Transmission_Gate_Layout_3.CLK.t36 Transmission_Gate_Layout_3.CLK.t64 82.9076
R8389 Transmission_Gate_Layout_3.CLK.t53 Transmission_Gate_Layout_3.CLK.t48 82.9076
R8390 Transmission_Gate_Layout_3.CLK.t28 Transmission_Gate_Layout_3.CLK.t53 82.9076
R8391 Transmission_Gate_Layout_3.CLK.t21 Transmission_Gate_Layout_3.CLK.n6 56.4451
R8392 Transmission_Gate_Layout_3.CLK.t11 Transmission_Gate_Layout_3.CLK.n32 56.4451
R8393 Transmission_Gate_Layout_3.CLK.n25 Transmission_Gate_Layout_3.CLK.t36 49.7969
R8394 Transmission_Gate_Layout_3.CLK.n51 Transmission_Gate_Layout_3.CLK.t28 49.7969
R8395 Transmission_Gate_Layout_3.CLK.n0 Transmission_Gate_Layout_3.CLK.t35 39.7594
R8396 Transmission_Gate_Layout_3.CLK.n26 Transmission_Gate_Layout_3.CLK.t23 39.7594
R8397 Transmission_Gate_Layout_3.CLK.n8 Transmission_Gate_Layout_3.CLK.n7 35.0405
R8398 Transmission_Gate_Layout_3.CLK.n24 Transmission_Gate_Layout_3.CLK.n23 35.0405
R8399 Transmission_Gate_Layout_3.CLK.n34 Transmission_Gate_Layout_3.CLK.n33 35.0405
R8400 Transmission_Gate_Layout_3.CLK.n50 Transmission_Gate_Layout_3.CLK.n49 35.0405
R8401 Transmission_Gate_Layout_3.CLK.n25 Transmission_Gate_Layout_3.CLK.t61 31.1559
R8402 Transmission_Gate_Layout_3.CLK.n51 Transmission_Gate_Layout_3.CLK.t50 31.1559
R8403 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_3.CLK.n53 24.3453
R8404 Transmission_Gate_Layout_3.CLK.n52 Transmission_Gate_Layout_3.CLK.t18 22.0309
R8405 Transmission_Gate_Layout_3.CLK.t56 Transmission_Gate_Layout_3.CLK.n15 21.9005
R8406 Transmission_Gate_Layout_3.CLK.n14 Transmission_Gate_Layout_3.CLK.t6 21.9005
R8407 Transmission_Gate_Layout_3.CLK.n13 Transmission_Gate_Layout_3.CLK.t20 21.9005
R8408 Transmission_Gate_Layout_3.CLK.n12 Transmission_Gate_Layout_3.CLK.t52 21.9005
R8409 Transmission_Gate_Layout_3.CLK.n11 Transmission_Gate_Layout_3.CLK.t16 21.9005
R8410 Transmission_Gate_Layout_3.CLK.n10 Transmission_Gate_Layout_3.CLK.t49 21.9005
R8411 Transmission_Gate_Layout_3.CLK.n9 Transmission_Gate_Layout_3.CLK.t2 21.9005
R8412 Transmission_Gate_Layout_3.CLK.n7 Transmission_Gate_Layout_3.CLK.t41 21.9005
R8413 Transmission_Gate_Layout_3.CLK.n8 Transmission_Gate_Layout_3.CLK.t14 21.9005
R8414 Transmission_Gate_Layout_3.CLK.n33 Transmission_Gate_Layout_3.CLK.t33 21.9005
R8415 Transmission_Gate_Layout_3.CLK.n34 Transmission_Gate_Layout_3.CLK.t4 21.9005
R8416 Transmission_Gate_Layout_3.CLK.n35 Transmission_Gate_Layout_3.CLK.t17 21.9005
R8417 Transmission_Gate_Layout_3.CLK.n36 Transmission_Gate_Layout_3.CLK.t51 21.9005
R8418 Transmission_Gate_Layout_3.CLK.n37 Transmission_Gate_Layout_3.CLK.t3 21.9005
R8419 Transmission_Gate_Layout_3.CLK.n38 Transmission_Gate_Layout_3.CLK.t39 21.9005
R8420 Transmission_Gate_Layout_3.CLK.n39 Transmission_Gate_Layout_3.CLK.t57 21.9005
R8421 Transmission_Gate_Layout_3.CLK.n40 Transmission_Gate_Layout_3.CLK.t8 21.9005
R8422 Transmission_Gate_Layout_3.CLK.t42 Transmission_Gate_Layout_3.CLK.n41 21.9005
R8423 Transmission_Gate_Layout_3.CLK.n16 Transmission_Gate_Layout_3.CLK.t56 21.5094
R8424 Transmission_Gate_Layout_3.CLK.n17 Transmission_Gate_Layout_3.CLK.t6 21.5094
R8425 Transmission_Gate_Layout_3.CLK.n18 Transmission_Gate_Layout_3.CLK.t20 21.5094
R8426 Transmission_Gate_Layout_3.CLK.n19 Transmission_Gate_Layout_3.CLK.t52 21.5094
R8427 Transmission_Gate_Layout_3.CLK.n20 Transmission_Gate_Layout_3.CLK.t16 21.5094
R8428 Transmission_Gate_Layout_3.CLK.n21 Transmission_Gate_Layout_3.CLK.t49 21.5094
R8429 Transmission_Gate_Layout_3.CLK.n22 Transmission_Gate_Layout_3.CLK.t2 21.5094
R8430 Transmission_Gate_Layout_3.CLK.n24 Transmission_Gate_Layout_3.CLK.t41 21.5094
R8431 Transmission_Gate_Layout_3.CLK.n23 Transmission_Gate_Layout_3.CLK.t14 21.5094
R8432 Transmission_Gate_Layout_3.CLK.n50 Transmission_Gate_Layout_3.CLK.t33 21.5094
R8433 Transmission_Gate_Layout_3.CLK.n49 Transmission_Gate_Layout_3.CLK.t4 21.5094
R8434 Transmission_Gate_Layout_3.CLK.n48 Transmission_Gate_Layout_3.CLK.t17 21.5094
R8435 Transmission_Gate_Layout_3.CLK.n47 Transmission_Gate_Layout_3.CLK.t51 21.5094
R8436 Transmission_Gate_Layout_3.CLK.n46 Transmission_Gate_Layout_3.CLK.t3 21.5094
R8437 Transmission_Gate_Layout_3.CLK.n45 Transmission_Gate_Layout_3.CLK.t39 21.5094
R8438 Transmission_Gate_Layout_3.CLK.n44 Transmission_Gate_Layout_3.CLK.t57 21.5094
R8439 Transmission_Gate_Layout_3.CLK.n43 Transmission_Gate_Layout_3.CLK.t8 21.5094
R8440 Transmission_Gate_Layout_3.CLK.n42 Transmission_Gate_Layout_3.CLK.t42 21.5094
R8441 Transmission_Gate_Layout_3.CLK.n52 Transmission_Gate_Layout_3.CLK.t25 21.3791
R8442 Transmission_Gate_Layout_3.CLK.n53 Transmission_Gate_Layout_3.CLK.t12 21.3791
R8443 Transmission_Gate_Layout_3.CLK.n16 Transmission_Gate_Layout_3.CLK.t10 20.988
R8444 Transmission_Gate_Layout_3.CLK.n17 Transmission_Gate_Layout_3.CLK.t26 20.988
R8445 Transmission_Gate_Layout_3.CLK.n18 Transmission_Gate_Layout_3.CLK.t40 20.988
R8446 Transmission_Gate_Layout_3.CLK.n19 Transmission_Gate_Layout_3.CLK.t9 20.988
R8447 Transmission_Gate_Layout_3.CLK.n20 Transmission_Gate_Layout_3.CLK.t34 20.988
R8448 Transmission_Gate_Layout_3.CLK.n21 Transmission_Gate_Layout_3.CLK.t5 20.988
R8449 Transmission_Gate_Layout_3.CLK.n22 Transmission_Gate_Layout_3.CLK.t19 20.988
R8450 Transmission_Gate_Layout_3.CLK.n23 Transmission_Gate_Layout_3.CLK.t31 20.988
R8451 Transmission_Gate_Layout_3.CLK.t61 Transmission_Gate_Layout_3.CLK.n24 20.988
R8452 Transmission_Gate_Layout_3.CLK.n49 Transmission_Gate_Layout_3.CLK.t24 20.988
R8453 Transmission_Gate_Layout_3.CLK.n48 Transmission_Gate_Layout_3.CLK.t38 20.988
R8454 Transmission_Gate_Layout_3.CLK.n47 Transmission_Gate_Layout_3.CLK.t7 20.988
R8455 Transmission_Gate_Layout_3.CLK.n46 Transmission_Gate_Layout_3.CLK.t22 20.988
R8456 Transmission_Gate_Layout_3.CLK.n45 Transmission_Gate_Layout_3.CLK.t54 20.988
R8457 Transmission_Gate_Layout_3.CLK.n44 Transmission_Gate_Layout_3.CLK.t13 20.988
R8458 Transmission_Gate_Layout_3.CLK.n43 Transmission_Gate_Layout_3.CLK.t27 20.988
R8459 Transmission_Gate_Layout_3.CLK.n42 Transmission_Gate_Layout_3.CLK.t62 20.988
R8460 Transmission_Gate_Layout_3.CLK.t50 Transmission_Gate_Layout_3.CLK.n50 20.988
R8461 Transmission_Gate_Layout_3.CLK.n1 Transmission_Gate_Layout_3.CLK.n0 20.8576
R8462 Transmission_Gate_Layout_3.CLK.n2 Transmission_Gate_Layout_3.CLK.n1 20.8576
R8463 Transmission_Gate_Layout_3.CLK.n3 Transmission_Gate_Layout_3.CLK.n2 20.8576
R8464 Transmission_Gate_Layout_3.CLK.n4 Transmission_Gate_Layout_3.CLK.n3 20.8576
R8465 Transmission_Gate_Layout_3.CLK.n5 Transmission_Gate_Layout_3.CLK.n4 20.8576
R8466 Transmission_Gate_Layout_3.CLK.n6 Transmission_Gate_Layout_3.CLK.n5 20.8576
R8467 Transmission_Gate_Layout_3.CLK.n32 Transmission_Gate_Layout_3.CLK.n31 20.8576
R8468 Transmission_Gate_Layout_3.CLK.n31 Transmission_Gate_Layout_3.CLK.n30 20.8576
R8469 Transmission_Gate_Layout_3.CLK.n30 Transmission_Gate_Layout_3.CLK.n29 20.8576
R8470 Transmission_Gate_Layout_3.CLK.n29 Transmission_Gate_Layout_3.CLK.n28 20.8576
R8471 Transmission_Gate_Layout_3.CLK.n28 Transmission_Gate_Layout_3.CLK.n27 20.8576
R8472 Transmission_Gate_Layout_3.CLK.n27 Transmission_Gate_Layout_3.CLK.n26 20.8576
R8473 Transmission_Gate_Layout_3.CLK.n53 Transmission_Gate_Layout_3.CLK.n52 20.8576
R8474 Transmission_Gate_Layout_3.CLK.n15 Transmission_Gate_Layout_3.CLK.t35 20.5969
R8475 Transmission_Gate_Layout_3.CLK.n14 Transmission_Gate_Layout_3.CLK.t46 20.5969
R8476 Transmission_Gate_Layout_3.CLK.n13 Transmission_Gate_Layout_3.CLK.t63 20.5969
R8477 Transmission_Gate_Layout_3.CLK.n12 Transmission_Gate_Layout_3.CLK.t32 20.5969
R8478 Transmission_Gate_Layout_3.CLK.n11 Transmission_Gate_Layout_3.CLK.t58 20.5969
R8479 Transmission_Gate_Layout_3.CLK.n10 Transmission_Gate_Layout_3.CLK.t29 20.5969
R8480 Transmission_Gate_Layout_3.CLK.n9 Transmission_Gate_Layout_3.CLK.t43 20.5969
R8481 Transmission_Gate_Layout_3.CLK.n8 Transmission_Gate_Layout_3.CLK.t55 20.5969
R8482 Transmission_Gate_Layout_3.CLK.n7 Transmission_Gate_Layout_3.CLK.t21 20.5969
R8483 Transmission_Gate_Layout_3.CLK.n33 Transmission_Gate_Layout_3.CLK.t11 20.5969
R8484 Transmission_Gate_Layout_3.CLK.n34 Transmission_Gate_Layout_3.CLK.t45 20.5969
R8485 Transmission_Gate_Layout_3.CLK.n35 Transmission_Gate_Layout_3.CLK.t60 20.5969
R8486 Transmission_Gate_Layout_3.CLK.n36 Transmission_Gate_Layout_3.CLK.t30 20.5969
R8487 Transmission_Gate_Layout_3.CLK.n37 Transmission_Gate_Layout_3.CLK.t44 20.5969
R8488 Transmission_Gate_Layout_3.CLK.n38 Transmission_Gate_Layout_3.CLK.t15 20.5969
R8489 Transmission_Gate_Layout_3.CLK.n39 Transmission_Gate_Layout_3.CLK.t37 20.5969
R8490 Transmission_Gate_Layout_3.CLK.n41 Transmission_Gate_Layout_3.CLK.t23 20.5969
R8491 Transmission_Gate_Layout_3.CLK.n40 Transmission_Gate_Layout_3.CLK.t47 20.5969
R8492 Transmission_Gate_Layout_3.CLK.n15 Transmission_Gate_Layout_3.CLK.n14 19.4672
R8493 Transmission_Gate_Layout_3.CLK.n14 Transmission_Gate_Layout_3.CLK.n13 19.4672
R8494 Transmission_Gate_Layout_3.CLK.n13 Transmission_Gate_Layout_3.CLK.n12 19.4672
R8495 Transmission_Gate_Layout_3.CLK.n12 Transmission_Gate_Layout_3.CLK.n11 19.4672
R8496 Transmission_Gate_Layout_3.CLK.n11 Transmission_Gate_Layout_3.CLK.n10 19.4672
R8497 Transmission_Gate_Layout_3.CLK.n10 Transmission_Gate_Layout_3.CLK.n9 19.4672
R8498 Transmission_Gate_Layout_3.CLK.n9 Transmission_Gate_Layout_3.CLK.n8 19.4672
R8499 Transmission_Gate_Layout_3.CLK.n17 Transmission_Gate_Layout_3.CLK.n16 19.4672
R8500 Transmission_Gate_Layout_3.CLK.n18 Transmission_Gate_Layout_3.CLK.n17 19.4672
R8501 Transmission_Gate_Layout_3.CLK.n19 Transmission_Gate_Layout_3.CLK.n18 19.4672
R8502 Transmission_Gate_Layout_3.CLK.n20 Transmission_Gate_Layout_3.CLK.n19 19.4672
R8503 Transmission_Gate_Layout_3.CLK.n21 Transmission_Gate_Layout_3.CLK.n20 19.4672
R8504 Transmission_Gate_Layout_3.CLK.n22 Transmission_Gate_Layout_3.CLK.n21 19.4672
R8505 Transmission_Gate_Layout_3.CLK.n23 Transmission_Gate_Layout_3.CLK.n22 19.4672
R8506 Transmission_Gate_Layout_3.CLK.n35 Transmission_Gate_Layout_3.CLK.n34 19.4672
R8507 Transmission_Gate_Layout_3.CLK.n36 Transmission_Gate_Layout_3.CLK.n35 19.4672
R8508 Transmission_Gate_Layout_3.CLK.n37 Transmission_Gate_Layout_3.CLK.n36 19.4672
R8509 Transmission_Gate_Layout_3.CLK.n38 Transmission_Gate_Layout_3.CLK.n37 19.4672
R8510 Transmission_Gate_Layout_3.CLK.n39 Transmission_Gate_Layout_3.CLK.n38 19.4672
R8511 Transmission_Gate_Layout_3.CLK.n40 Transmission_Gate_Layout_3.CLK.n39 19.4672
R8512 Transmission_Gate_Layout_3.CLK.n41 Transmission_Gate_Layout_3.CLK.n40 19.4672
R8513 Transmission_Gate_Layout_3.CLK.n49 Transmission_Gate_Layout_3.CLK.n48 19.4672
R8514 Transmission_Gate_Layout_3.CLK.n48 Transmission_Gate_Layout_3.CLK.n47 19.4672
R8515 Transmission_Gate_Layout_3.CLK.n47 Transmission_Gate_Layout_3.CLK.n46 19.4672
R8516 Transmission_Gate_Layout_3.CLK.n46 Transmission_Gate_Layout_3.CLK.n45 19.4672
R8517 Transmission_Gate_Layout_3.CLK.n45 Transmission_Gate_Layout_3.CLK.n44 19.4672
R8518 Transmission_Gate_Layout_3.CLK.n44 Transmission_Gate_Layout_3.CLK.n43 19.4672
R8519 Transmission_Gate_Layout_3.CLK.n43 Transmission_Gate_Layout_3.CLK.n42 19.4672
R8520 Transmission_Gate_Layout_3.CLK.n0 Transmission_Gate_Layout_3.CLK.t46 18.9023
R8521 Transmission_Gate_Layout_3.CLK.n1 Transmission_Gate_Layout_3.CLK.t63 18.9023
R8522 Transmission_Gate_Layout_3.CLK.n2 Transmission_Gate_Layout_3.CLK.t32 18.9023
R8523 Transmission_Gate_Layout_3.CLK.n3 Transmission_Gate_Layout_3.CLK.t58 18.9023
R8524 Transmission_Gate_Layout_3.CLK.n4 Transmission_Gate_Layout_3.CLK.t29 18.9023
R8525 Transmission_Gate_Layout_3.CLK.n5 Transmission_Gate_Layout_3.CLK.t43 18.9023
R8526 Transmission_Gate_Layout_3.CLK.n6 Transmission_Gate_Layout_3.CLK.t55 18.9023
R8527 Transmission_Gate_Layout_3.CLK.n32 Transmission_Gate_Layout_3.CLK.t45 18.9023
R8528 Transmission_Gate_Layout_3.CLK.n31 Transmission_Gate_Layout_3.CLK.t60 18.9023
R8529 Transmission_Gate_Layout_3.CLK.n30 Transmission_Gate_Layout_3.CLK.t30 18.9023
R8530 Transmission_Gate_Layout_3.CLK.n29 Transmission_Gate_Layout_3.CLK.t44 18.9023
R8531 Transmission_Gate_Layout_3.CLK.n28 Transmission_Gate_Layout_3.CLK.t15 18.9023
R8532 Transmission_Gate_Layout_3.CLK.n27 Transmission_Gate_Layout_3.CLK.t37 18.9023
R8533 Transmission_Gate_Layout_3.CLK.n26 Transmission_Gate_Layout_3.CLK.t47 18.9023
R8534 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_3.CLK.n25 16.4436
R8535 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_3.CLK.n51 16.4434
R8536 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_3.CLK.n54 7.70137
R8537 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_3.CLK.n55 4.70224
R8538 Transmission_Gate_Layout_14.CLKB.n24 Transmission_Gate_Layout_14.CLKB.t24 54.5477
R8539 Transmission_Gate_Layout_14.CLKB.n29 Transmission_Gate_Layout_14.CLKB.t15 38.3255
R8540 Transmission_Gate_Layout_14.CLKB.n28 Transmission_Gate_Layout_14.CLKB.t27 38.3255
R8541 Transmission_Gate_Layout_14.CLKB.n27 Transmission_Gate_Layout_14.CLKB.t7 38.3255
R8542 Transmission_Gate_Layout_14.CLKB.n26 Transmission_Gate_Layout_14.CLKB.t12 38.3255
R8543 Transmission_Gate_Layout_14.CLKB.n25 Transmission_Gate_Layout_14.CLKB.t29 38.3255
R8544 Transmission_Gate_Layout_14.CLKB.n24 Transmission_Gate_Layout_14.CLKB.t9 38.3255
R8545 Transmission_Gate_Layout_14.CLKB.t26 Transmission_Gate_Layout_14.CLKB.n2 37.9344
R8546 Transmission_Gate_Layout_14.CLKB.t13 Transmission_Gate_Layout_14.CLKB.n5 37.9344
R8547 Transmission_Gate_Layout_14.CLKB.t19 Transmission_Gate_Layout_14.CLKB.n8 37.9344
R8548 Transmission_Gate_Layout_14.CLKB.t25 Transmission_Gate_Layout_14.CLKB.n11 37.9344
R8549 Transmission_Gate_Layout_14.CLKB.t17 Transmission_Gate_Layout_14.CLKB.n14 37.9344
R8550 Transmission_Gate_Layout_14.CLKB.t21 Transmission_Gate_Layout_14.CLKB.n17 37.9344
R8551 Transmission_Gate_Layout_14.CLKB.t8 Transmission_Gate_Layout_14.CLKB.n20 37.9344
R8552 Transmission_Gate_Layout_14.CLKB.t16 Transmission_Gate_Layout_14.CLKB.n21 37.9344
R8553 Transmission_Gate_Layout_14.CLKB.n3 Transmission_Gate_Layout_14.CLKB.t26 37.5434
R8554 Transmission_Gate_Layout_14.CLKB.n6 Transmission_Gate_Layout_14.CLKB.t13 37.5434
R8555 Transmission_Gate_Layout_14.CLKB.n9 Transmission_Gate_Layout_14.CLKB.t19 37.5434
R8556 Transmission_Gate_Layout_14.CLKB.n12 Transmission_Gate_Layout_14.CLKB.t25 37.5434
R8557 Transmission_Gate_Layout_14.CLKB.n15 Transmission_Gate_Layout_14.CLKB.t17 37.5434
R8558 Transmission_Gate_Layout_14.CLKB.n18 Transmission_Gate_Layout_14.CLKB.t21 37.5434
R8559 Transmission_Gate_Layout_14.CLKB.n23 Transmission_Gate_Layout_14.CLKB.t8 37.5434
R8560 Transmission_Gate_Layout_14.CLKB.n22 Transmission_Gate_Layout_14.CLKB.t16 37.5434
R8561 Transmission_Gate_Layout_14.CLKB.t15 Transmission_Gate_Layout_14.CLKB.n3 37.413
R8562 Transmission_Gate_Layout_14.CLKB.t27 Transmission_Gate_Layout_14.CLKB.n6 37.413
R8563 Transmission_Gate_Layout_14.CLKB.t7 Transmission_Gate_Layout_14.CLKB.n9 37.413
R8564 Transmission_Gate_Layout_14.CLKB.t12 Transmission_Gate_Layout_14.CLKB.n12 37.413
R8565 Transmission_Gate_Layout_14.CLKB.t29 Transmission_Gate_Layout_14.CLKB.n15 37.413
R8566 Transmission_Gate_Layout_14.CLKB.t9 Transmission_Gate_Layout_14.CLKB.n18 37.413
R8567 Transmission_Gate_Layout_14.CLKB.n22 Transmission_Gate_Layout_14.CLKB.t28 37.413
R8568 Transmission_Gate_Layout_14.CLKB.t24 Transmission_Gate_Layout_14.CLKB.n23 37.413
R8569 Transmission_Gate_Layout_14.CLKB.n21 Transmission_Gate_Layout_14.CLKB.t11 37.0219
R8570 Transmission_Gate_Layout_14.CLKB.n17 Transmission_Gate_Layout_14.CLKB.t20 37.0219
R8571 Transmission_Gate_Layout_14.CLKB.n14 Transmission_Gate_Layout_14.CLKB.t14 37.0219
R8572 Transmission_Gate_Layout_14.CLKB.n11 Transmission_Gate_Layout_14.CLKB.t22 37.0219
R8573 Transmission_Gate_Layout_14.CLKB.n8 Transmission_Gate_Layout_14.CLKB.t18 37.0219
R8574 Transmission_Gate_Layout_14.CLKB.n5 Transmission_Gate_Layout_14.CLKB.t10 37.0219
R8575 Transmission_Gate_Layout_14.CLKB.n2 Transmission_Gate_Layout_14.CLKB.t23 37.0219
R8576 Transmission_Gate_Layout_14.CLKB.n20 Transmission_Gate_Layout_14.CLKB.t6 37.0219
R8577 Transmission_Gate_Layout_14.CLKB.t20 Transmission_Gate_Layout_14.CLKB.n16 35.1969
R8578 Transmission_Gate_Layout_14.CLKB.t14 Transmission_Gate_Layout_14.CLKB.n13 35.1969
R8579 Transmission_Gate_Layout_14.CLKB.t22 Transmission_Gate_Layout_14.CLKB.n10 35.1969
R8580 Transmission_Gate_Layout_14.CLKB.t18 Transmission_Gate_Layout_14.CLKB.n7 35.1969
R8581 Transmission_Gate_Layout_14.CLKB.t10 Transmission_Gate_Layout_14.CLKB.n4 35.1969
R8582 Transmission_Gate_Layout_14.CLKB.t6 Transmission_Gate_Layout_14.CLKB.n19 35.1969
R8583 Transmission_Gate_Layout_14.CLKB Transmission_Gate_Layout_14.CLKB.n29 26.6826
R8584 Transmission_Gate_Layout_14.CLKB.n23 Transmission_Gate_Layout_14.CLKB.n22 19.148
R8585 Transmission_Gate_Layout_14.CLKB.n29 Transmission_Gate_Layout_14.CLKB.n28 16.2227
R8586 Transmission_Gate_Layout_14.CLKB.n28 Transmission_Gate_Layout_14.CLKB.n27 16.2227
R8587 Transmission_Gate_Layout_14.CLKB.n27 Transmission_Gate_Layout_14.CLKB.n26 16.2227
R8588 Transmission_Gate_Layout_14.CLKB.n26 Transmission_Gate_Layout_14.CLKB.n25 16.2227
R8589 Transmission_Gate_Layout_14.CLKB.n25 Transmission_Gate_Layout_14.CLKB.n24 16.2227
R8590 Transmission_Gate_Layout_14.CLKB.n30 Transmission_Gate_Layout_14.CLKB.t4 5.21612
R8591 Transmission_Gate_Layout_14.CLKB.n0 Transmission_Gate_Layout_14.CLKB.t2 4.57285
R8592 Transmission_Gate_Layout_14.CLKB.n31 Transmission_Gate_Layout_14.CLKB.t5 4.4609
R8593 Transmission_Gate_Layout_14.CLKB.n30 Transmission_Gate_Layout_14.CLKB.t3 4.4609
R8594 Transmission_Gate_Layout_14.CLKB.n0 Transmission_Gate_Layout_14.CLKB.t1 3.3285
R8595 Transmission_Gate_Layout_14.CLKB.n1 Transmission_Gate_Layout_14.CLKB.t0 3.3285
R8596 Transmission_Gate_Layout_14.CLKB.n1 Transmission_Gate_Layout_14.CLKB.n0 1.24485
R8597 Transmission_Gate_Layout_14.CLKB.n31 Transmission_Gate_Layout_14.CLKB.n30 0.755717
R8598 Transmission_Gate_Layout_14.CLKB Transmission_Gate_Layout_14.CLKB.n1 0.750969
R8599 Transmission_Gate_Layout_14.CLKB Transmission_Gate_Layout_14.CLKB.n31 0.510317
R8600 IN3.n68 IN3 8.12709
R8601 IN3.n14 IN3.n13 3.90572
R8602 IN3.n60 IN3.n57 3.90572
R8603 IN3.n52 IN3.n49 3.90572
R8604 IN3.n4 IN3.n1 3.84485
R8605 IN3.n22 IN3.n21 3.84485
R8606 IN3.n30 IN3.n29 3.84485
R8607 IN3.n14 IN3.n11 3.1505
R8608 IN3.n15 IN3.n9 3.1505
R8609 IN3.n60 IN3.n59 3.1505
R8610 IN3.n63 IN3.n62 3.1505
R8611 IN3.n52 IN3.n51 3.1505
R8612 IN3.n55 IN3.n54 3.1505
R8613 IN3.n65 IN3.n47 3.1505
R8614 IN3.n66 IN3.n45 3.1505
R8615 IN3.n67 IN3.n43 3.1505
R8616 IN3.n7 IN3.n6 2.6005
R8617 IN3.n4 IN3.n3 2.6005
R8618 IN3.n22 IN3.n19 2.6005
R8619 IN3.n23 IN3.n17 2.6005
R8620 IN3.n30 IN3.n27 2.6005
R8621 IN3.n31 IN3.n25 2.6005
R8622 IN3.n35 IN3.n34 2.6005
R8623 IN3.n38 IN3.n37 2.6005
R8624 IN3.n41 IN3.n40 2.6005
R8625 IN3.n9 IN3.t46 1.3109
R8626 IN3.n9 IN3.n8 1.3109
R8627 IN3.n11 IN3.t38 1.3109
R8628 IN3.n11 IN3.n10 1.3109
R8629 IN3.n13 IN3.t41 1.3109
R8630 IN3.n13 IN3.n12 1.3109
R8631 IN3.n43 IN3.t44 1.3109
R8632 IN3.n43 IN3.n42 1.3109
R8633 IN3.n45 IN3.t36 1.3109
R8634 IN3.n45 IN3.n44 1.3109
R8635 IN3.n47 IN3.t39 1.3109
R8636 IN3.n47 IN3.n46 1.3109
R8637 IN3.n62 IN3.t47 1.3109
R8638 IN3.n62 IN3.n61 1.3109
R8639 IN3.n59 IN3.t43 1.3109
R8640 IN3.n59 IN3.n58 1.3109
R8641 IN3.n57 IN3.t40 1.3109
R8642 IN3.n57 IN3.n56 1.3109
R8643 IN3.n54 IN3.t37 1.3109
R8644 IN3.n54 IN3.n53 1.3109
R8645 IN3.n51 IN3.t45 1.3109
R8646 IN3.n51 IN3.n50 1.3109
R8647 IN3.n49 IN3.t42 1.3109
R8648 IN3.n49 IN3.n48 1.3109
R8649 IN3.n7 IN3.n4 1.24485
R8650 IN3.n23 IN3.n22 1.24485
R8651 IN3.n31 IN3.n30 1.24485
R8652 IN3.n38 IN3.n35 1.24485
R8653 IN3.n41 IN3.n38 1.24485
R8654 IN3.n32 IN3.n31 1.2018
R8655 IN3.n35 IN3.n32 1.2018
R8656 IN3.n64 IN3.n63 0.957239
R8657 IN3.n65 IN3.n64 0.957239
R8658 IN3.n68 IN3.n41 0.822239
R8659 IN3.n69 IN3.n7 0.806587
R8660 IN3.n15 IN3.n14 0.755717
R8661 IN3.n63 IN3.n60 0.755717
R8662 IN3.n55 IN3.n52 0.755717
R8663 IN3.n67 IN3.n66 0.755717
R8664 IN3.n66 IN3.n65 0.755717
R8665 IN3.n1 IN3.t23 0.7285
R8666 IN3.n1 IN3.n0 0.7285
R8667 IN3.n3 IN3.t21 0.7285
R8668 IN3.n3 IN3.n2 0.7285
R8669 IN3.n6 IN3.t14 0.7285
R8670 IN3.n6 IN3.n5 0.7285
R8671 IN3.n40 IN3.t12 0.7285
R8672 IN3.n40 IN3.n39 0.7285
R8673 IN3.n37 IN3.t18 0.7285
R8674 IN3.n37 IN3.n36 0.7285
R8675 IN3.n34 IN3.t20 0.7285
R8676 IN3.n34 IN3.n33 0.7285
R8677 IN3.n17 IN3.t17 0.7285
R8678 IN3.n17 IN3.n16 0.7285
R8679 IN3.n19 IN3.t16 0.7285
R8680 IN3.n19 IN3.n18 0.7285
R8681 IN3.n21 IN3.t22 0.7285
R8682 IN3.n21 IN3.n20 0.7285
R8683 IN3.n25 IN3.t15 0.7285
R8684 IN3.n25 IN3.n24 0.7285
R8685 IN3.n27 IN3.t13 0.7285
R8686 IN3.n27 IN3.n26 0.7285
R8687 IN3.n29 IN3.t19 0.7285
R8688 IN3.n29 IN3.n28 0.7285
R8689 IN3.n32 IN3.n23 0.575717
R8690 IN3.n69 IN3.n68 0.552239
R8691 IN3.n68 IN3.n67 0.44463
R8692 IN3.n69 IN3.n15 0.428978
R8693 IN3.n64 IN3.n55 0.331152
R8694 IN3 IN3.n69 0.192239
R8695 Transmission_Gate_Layout_10.VIN.n119 Transmission_Gate_Layout_10.VIN.n118 25.4203
R8696 Transmission_Gate_Layout_10.VIN.n46 Transmission_Gate_Layout_10.VIN.t90 5.21612
R8697 Transmission_Gate_Layout_10.VIN.n121 Transmission_Gate_Layout_10.VIN.n37 4.4609
R8698 Transmission_Gate_Layout_10.VIN.n122 Transmission_Gate_Layout_10.VIN.n36 4.4609
R8699 Transmission_Gate_Layout_10.VIN.n123 Transmission_Gate_Layout_10.VIN.n35 4.4609
R8700 Transmission_Gate_Layout_10.VIN.n47 Transmission_Gate_Layout_10.VIN.t81 4.4609
R8701 Transmission_Gate_Layout_10.VIN.n46 Transmission_Gate_Layout_10.VIN.t74 4.4609
R8702 Transmission_Gate_Layout_10.VIN.n25 Transmission_Gate_Layout_10.VIN.n24 3.90572
R8703 Transmission_Gate_Layout_10.VIN.n33 Transmission_Gate_Layout_10.VIN.n32 3.90572
R8704 Transmission_Gate_Layout_10.VIN.n42 Transmission_Gate_Layout_10.VIN.n39 3.90572
R8705 Transmission_Gate_Layout_10.VIN.n92 Transmission_Gate_Layout_10.VIN.n89 3.90572
R8706 Transmission_Gate_Layout_10.VIN.n54 Transmission_Gate_Layout_10.VIN.n53 3.90572
R8707 Transmission_Gate_Layout_10.VIN.n116 Transmission_Gate_Layout_10.VIN.n115 3.90572
R8708 Transmission_Gate_Layout_10.VIN.n7 Transmission_Gate_Layout_10.VIN.n4 3.84485
R8709 Transmission_Gate_Layout_10.VIN.n80 Transmission_Gate_Layout_10.VIN.n77 3.84485
R8710 Transmission_Gate_Layout_10.VIN.n72 Transmission_Gate_Layout_10.VIN.n69 3.84485
R8711 Transmission_Gate_Layout_10.VIN.n102 Transmission_Gate_Layout_10.VIN.n101 3.84485
R8712 Transmission_Gate_Layout_10.VIN.n15 Transmission_Gate_Layout_10.VIN.n12 3.84485
R8713 Transmission_Gate_Layout_10.VIN.n135 Transmission_Gate_Layout_10.VIN.n134 3.84485
R8714 Transmission_Gate_Layout_10.VIN.n128 Transmission_Gate_Layout_10.VIN.n2 3.3285
R8715 Transmission_Gate_Layout_10.VIN.n129 Transmission_Gate_Layout_10.VIN.n1 3.3285
R8716 Transmission_Gate_Layout_10.VIN.n130 Transmission_Gate_Layout_10.VIN.n0 3.3285
R8717 Transmission_Gate_Layout_10.VIN.n140 Transmission_Gate_Layout_10.VIN.t18 3.3285
R8718 Transmission_Gate_Layout_10.VIN.n141 Transmission_Gate_Layout_10.VIN.t13 3.3285
R8719 Transmission_Gate_Layout_10.VIN.n142 Transmission_Gate_Layout_10.VIN.t1 3.3285
R8720 Transmission_Gate_Layout_10.VIN.n25 Transmission_Gate_Layout_10.VIN.n22 3.1505
R8721 Transmission_Gate_Layout_10.VIN.n26 Transmission_Gate_Layout_10.VIN.n20 3.1505
R8722 Transmission_Gate_Layout_10.VIN.n33 Transmission_Gate_Layout_10.VIN.n30 3.1505
R8723 Transmission_Gate_Layout_10.VIN.n34 Transmission_Gate_Layout_10.VIN.n28 3.1505
R8724 Transmission_Gate_Layout_10.VIN.n42 Transmission_Gate_Layout_10.VIN.n41 3.1505
R8725 Transmission_Gate_Layout_10.VIN.n45 Transmission_Gate_Layout_10.VIN.n44 3.1505
R8726 Transmission_Gate_Layout_10.VIN.n95 Transmission_Gate_Layout_10.VIN.n94 3.1505
R8727 Transmission_Gate_Layout_10.VIN.n92 Transmission_Gate_Layout_10.VIN.n91 3.1505
R8728 Transmission_Gate_Layout_10.VIN.n108 Transmission_Gate_Layout_10.VIN.n57 3.1505
R8729 Transmission_Gate_Layout_10.VIN.n107 Transmission_Gate_Layout_10.VIN.n59 3.1505
R8730 Transmission_Gate_Layout_10.VIN.n106 Transmission_Gate_Layout_10.VIN.n61 3.1505
R8731 Transmission_Gate_Layout_10.VIN.n54 Transmission_Gate_Layout_10.VIN.n51 3.1505
R8732 Transmission_Gate_Layout_10.VIN.n55 Transmission_Gate_Layout_10.VIN.n49 3.1505
R8733 Transmission_Gate_Layout_10.VIN.n116 Transmission_Gate_Layout_10.VIN.n113 3.1505
R8734 Transmission_Gate_Layout_10.VIN.n117 Transmission_Gate_Layout_10.VIN.n111 3.1505
R8735 Transmission_Gate_Layout_10.VIN.n139 Transmission_Gate_Layout_10.VIN.n130 2.72398
R8736 Transmission_Gate_Layout_10.VIN.n7 Transmission_Gate_Layout_10.VIN.n6 2.6005
R8737 Transmission_Gate_Layout_10.VIN.n10 Transmission_Gate_Layout_10.VIN.n9 2.6005
R8738 Transmission_Gate_Layout_10.VIN.n80 Transmission_Gate_Layout_10.VIN.n79 2.6005
R8739 Transmission_Gate_Layout_10.VIN.n83 Transmission_Gate_Layout_10.VIN.n82 2.6005
R8740 Transmission_Gate_Layout_10.VIN.n72 Transmission_Gate_Layout_10.VIN.n71 2.6005
R8741 Transmission_Gate_Layout_10.VIN.n75 Transmission_Gate_Layout_10.VIN.n74 2.6005
R8742 Transmission_Gate_Layout_10.VIN.n85 Transmission_Gate_Layout_10.VIN.n67 2.6005
R8743 Transmission_Gate_Layout_10.VIN.n86 Transmission_Gate_Layout_10.VIN.n65 2.6005
R8744 Transmission_Gate_Layout_10.VIN.n87 Transmission_Gate_Layout_10.VIN.n63 2.6005
R8745 Transmission_Gate_Layout_10.VIN.n102 Transmission_Gate_Layout_10.VIN.n99 2.6005
R8746 Transmission_Gate_Layout_10.VIN.n103 Transmission_Gate_Layout_10.VIN.n97 2.6005
R8747 Transmission_Gate_Layout_10.VIN.n15 Transmission_Gate_Layout_10.VIN.n14 2.6005
R8748 Transmission_Gate_Layout_10.VIN.n18 Transmission_Gate_Layout_10.VIN.n17 2.6005
R8749 Transmission_Gate_Layout_10.VIN.n135 Transmission_Gate_Layout_10.VIN.n132 2.6005
R8750 Transmission_Gate_Layout_10.VIN.n138 Transmission_Gate_Layout_10.VIN.n137 2.6005
R8751 Transmission_Gate_Layout_10.VIN.n121 Transmission_Gate_Layout_10.VIN.n120 2.47941
R8752 Transmission_Gate_Layout_10.VIN.n20 Transmission_Gate_Layout_10.VIN.t82 1.3109
R8753 Transmission_Gate_Layout_10.VIN.n20 Transmission_Gate_Layout_10.VIN.n19 1.3109
R8754 Transmission_Gate_Layout_10.VIN.n22 Transmission_Gate_Layout_10.VIN.t88 1.3109
R8755 Transmission_Gate_Layout_10.VIN.n22 Transmission_Gate_Layout_10.VIN.n21 1.3109
R8756 Transmission_Gate_Layout_10.VIN.n24 Transmission_Gate_Layout_10.VIN.t73 1.3109
R8757 Transmission_Gate_Layout_10.VIN.n24 Transmission_Gate_Layout_10.VIN.n23 1.3109
R8758 Transmission_Gate_Layout_10.VIN.n28 Transmission_Gate_Layout_10.VIN.t92 1.3109
R8759 Transmission_Gate_Layout_10.VIN.n28 Transmission_Gate_Layout_10.VIN.n27 1.3109
R8760 Transmission_Gate_Layout_10.VIN.n30 Transmission_Gate_Layout_10.VIN.t75 1.3109
R8761 Transmission_Gate_Layout_10.VIN.n30 Transmission_Gate_Layout_10.VIN.n29 1.3109
R8762 Transmission_Gate_Layout_10.VIN.n32 Transmission_Gate_Layout_10.VIN.t83 1.3109
R8763 Transmission_Gate_Layout_10.VIN.n32 Transmission_Gate_Layout_10.VIN.n31 1.3109
R8764 Transmission_Gate_Layout_10.VIN.n44 Transmission_Gate_Layout_10.VIN.t76 1.3109
R8765 Transmission_Gate_Layout_10.VIN.n44 Transmission_Gate_Layout_10.VIN.n43 1.3109
R8766 Transmission_Gate_Layout_10.VIN.n41 Transmission_Gate_Layout_10.VIN.t91 1.3109
R8767 Transmission_Gate_Layout_10.VIN.n41 Transmission_Gate_Layout_10.VIN.n40 1.3109
R8768 Transmission_Gate_Layout_10.VIN.n39 Transmission_Gate_Layout_10.VIN.t84 1.3109
R8769 Transmission_Gate_Layout_10.VIN.n39 Transmission_Gate_Layout_10.VIN.n38 1.3109
R8770 Transmission_Gate_Layout_10.VIN.n61 Transmission_Gate_Layout_10.VIN.t53 1.3109
R8771 Transmission_Gate_Layout_10.VIN.n61 Transmission_Gate_Layout_10.VIN.n60 1.3109
R8772 Transmission_Gate_Layout_10.VIN.n59 Transmission_Gate_Layout_10.VIN.t61 1.3109
R8773 Transmission_Gate_Layout_10.VIN.n59 Transmission_Gate_Layout_10.VIN.n58 1.3109
R8774 Transmission_Gate_Layout_10.VIN.n57 Transmission_Gate_Layout_10.VIN.t56 1.3109
R8775 Transmission_Gate_Layout_10.VIN.n57 Transmission_Gate_Layout_10.VIN.n56 1.3109
R8776 Transmission_Gate_Layout_10.VIN.n89 Transmission_Gate_Layout_10.VIN.t71 1.3109
R8777 Transmission_Gate_Layout_10.VIN.n89 Transmission_Gate_Layout_10.VIN.n88 1.3109
R8778 Transmission_Gate_Layout_10.VIN.n91 Transmission_Gate_Layout_10.VIN.t54 1.3109
R8779 Transmission_Gate_Layout_10.VIN.n91 Transmission_Gate_Layout_10.VIN.n90 1.3109
R8780 Transmission_Gate_Layout_10.VIN.n94 Transmission_Gate_Layout_10.VIN.t58 1.3109
R8781 Transmission_Gate_Layout_10.VIN.n94 Transmission_Gate_Layout_10.VIN.n93 1.3109
R8782 Transmission_Gate_Layout_10.VIN.n49 Transmission_Gate_Layout_10.VIN.t67 1.3109
R8783 Transmission_Gate_Layout_10.VIN.n49 Transmission_Gate_Layout_10.VIN.n48 1.3109
R8784 Transmission_Gate_Layout_10.VIN.n51 Transmission_Gate_Layout_10.VIN.t49 1.3109
R8785 Transmission_Gate_Layout_10.VIN.n51 Transmission_Gate_Layout_10.VIN.n50 1.3109
R8786 Transmission_Gate_Layout_10.VIN.n53 Transmission_Gate_Layout_10.VIN.t63 1.3109
R8787 Transmission_Gate_Layout_10.VIN.n53 Transmission_Gate_Layout_10.VIN.n52 1.3109
R8788 Transmission_Gate_Layout_10.VIN.n111 Transmission_Gate_Layout_10.VIN.t65 1.3109
R8789 Transmission_Gate_Layout_10.VIN.n111 Transmission_Gate_Layout_10.VIN.n110 1.3109
R8790 Transmission_Gate_Layout_10.VIN.n113 Transmission_Gate_Layout_10.VIN.t48 1.3109
R8791 Transmission_Gate_Layout_10.VIN.n113 Transmission_Gate_Layout_10.VIN.n112 1.3109
R8792 Transmission_Gate_Layout_10.VIN.n115 Transmission_Gate_Layout_10.VIN.t59 1.3109
R8793 Transmission_Gate_Layout_10.VIN.n115 Transmission_Gate_Layout_10.VIN.n114 1.3109
R8794 Transmission_Gate_Layout_10.VIN.n10 Transmission_Gate_Layout_10.VIN.n7 1.24485
R8795 Transmission_Gate_Layout_10.VIN.n83 Transmission_Gate_Layout_10.VIN.n80 1.24485
R8796 Transmission_Gate_Layout_10.VIN.n75 Transmission_Gate_Layout_10.VIN.n72 1.24485
R8797 Transmission_Gate_Layout_10.VIN.n87 Transmission_Gate_Layout_10.VIN.n86 1.24485
R8798 Transmission_Gate_Layout_10.VIN.n86 Transmission_Gate_Layout_10.VIN.n85 1.24485
R8799 Transmission_Gate_Layout_10.VIN.n103 Transmission_Gate_Layout_10.VIN.n102 1.24485
R8800 Transmission_Gate_Layout_10.VIN.n18 Transmission_Gate_Layout_10.VIN.n15 1.24485
R8801 Transmission_Gate_Layout_10.VIN.n130 Transmission_Gate_Layout_10.VIN.n129 1.24485
R8802 Transmission_Gate_Layout_10.VIN.n129 Transmission_Gate_Layout_10.VIN.n128 1.24485
R8803 Transmission_Gate_Layout_10.VIN.n141 Transmission_Gate_Layout_10.VIN.n140 1.24485
R8804 Transmission_Gate_Layout_10.VIN.n142 Transmission_Gate_Layout_10.VIN.n141 1.24485
R8805 Transmission_Gate_Layout_10.VIN.n138 Transmission_Gate_Layout_10.VIN.n135 1.24485
R8806 Transmission_Gate_Layout_10.VIN.n84 Transmission_Gate_Layout_10.VIN.n83 1.2018
R8807 Transmission_Gate_Layout_10.VIN.n85 Transmission_Gate_Layout_10.VIN.n84 1.2018
R8808 Transmission_Gate_Layout_10.VIN.n128 Transmission_Gate_Layout_10.VIN.n127 1.2018
R8809 Transmission_Gate_Layout_10.VIN.n140 Transmission_Gate_Layout_10.VIN.n139 1.2018
R8810 Transmission_Gate_Layout_10.VIN.n109 Transmission_Gate_Layout_10.VIN.n108 0.957239
R8811 Transmission_Gate_Layout_10.VIN.n124 Transmission_Gate_Layout_10.VIN.n123 0.957239
R8812 Transmission_Gate_Layout_10.VIN.n105 Transmission_Gate_Layout_10.VIN.n87 0.806587
R8813 Transmission_Gate_Layout_10.VIN.n104 Transmission_Gate_Layout_10.VIN.n103 0.806587
R8814 Transmission_Gate_Layout_10.VIN.n26 Transmission_Gate_Layout_10.VIN.n25 0.755717
R8815 Transmission_Gate_Layout_10.VIN.n34 Transmission_Gate_Layout_10.VIN.n33 0.755717
R8816 Transmission_Gate_Layout_10.VIN.n45 Transmission_Gate_Layout_10.VIN.n42 0.755717
R8817 Transmission_Gate_Layout_10.VIN.n95 Transmission_Gate_Layout_10.VIN.n92 0.755717
R8818 Transmission_Gate_Layout_10.VIN.n108 Transmission_Gate_Layout_10.VIN.n107 0.755717
R8819 Transmission_Gate_Layout_10.VIN.n107 Transmission_Gate_Layout_10.VIN.n106 0.755717
R8820 Transmission_Gate_Layout_10.VIN.n55 Transmission_Gate_Layout_10.VIN.n54 0.755717
R8821 Transmission_Gate_Layout_10.VIN.n117 Transmission_Gate_Layout_10.VIN.n116 0.755717
R8822 Transmission_Gate_Layout_10.VIN.n47 Transmission_Gate_Layout_10.VIN.n46 0.755717
R8823 Transmission_Gate_Layout_10.VIN.n123 Transmission_Gate_Layout_10.VIN.n122 0.755717
R8824 Transmission_Gate_Layout_10.VIN.n122 Transmission_Gate_Layout_10.VIN.n121 0.755717
R8825 Transmission_Gate_Layout_10.VIN.n132 Transmission_Gate_Layout_10.VIN.t8 0.7285
R8826 Transmission_Gate_Layout_10.VIN.n132 Transmission_Gate_Layout_10.VIN.n131 0.7285
R8827 Transmission_Gate_Layout_10.VIN.n134 Transmission_Gate_Layout_10.VIN.t20 0.7285
R8828 Transmission_Gate_Layout_10.VIN.n134 Transmission_Gate_Layout_10.VIN.n133 0.7285
R8829 Transmission_Gate_Layout_10.VIN.n9 Transmission_Gate_Layout_10.VIN.t2 0.7285
R8830 Transmission_Gate_Layout_10.VIN.n9 Transmission_Gate_Layout_10.VIN.n8 0.7285
R8831 Transmission_Gate_Layout_10.VIN.n6 Transmission_Gate_Layout_10.VIN.t16 0.7285
R8832 Transmission_Gate_Layout_10.VIN.n6 Transmission_Gate_Layout_10.VIN.n5 0.7285
R8833 Transmission_Gate_Layout_10.VIN.n4 Transmission_Gate_Layout_10.VIN.t19 0.7285
R8834 Transmission_Gate_Layout_10.VIN.n4 Transmission_Gate_Layout_10.VIN.n3 0.7285
R8835 Transmission_Gate_Layout_10.VIN.n63 Transmission_Gate_Layout_10.VIN.t31 0.7285
R8836 Transmission_Gate_Layout_10.VIN.n63 Transmission_Gate_Layout_10.VIN.n62 0.7285
R8837 Transmission_Gate_Layout_10.VIN.n65 Transmission_Gate_Layout_10.VIN.t37 0.7285
R8838 Transmission_Gate_Layout_10.VIN.n65 Transmission_Gate_Layout_10.VIN.n64 0.7285
R8839 Transmission_Gate_Layout_10.VIN.n67 Transmission_Gate_Layout_10.VIN.t46 0.7285
R8840 Transmission_Gate_Layout_10.VIN.n67 Transmission_Gate_Layout_10.VIN.n66 0.7285
R8841 Transmission_Gate_Layout_10.VIN.n82 Transmission_Gate_Layout_10.VIN.t40 0.7285
R8842 Transmission_Gate_Layout_10.VIN.n82 Transmission_Gate_Layout_10.VIN.n81 0.7285
R8843 Transmission_Gate_Layout_10.VIN.n79 Transmission_Gate_Layout_10.VIN.t30 0.7285
R8844 Transmission_Gate_Layout_10.VIN.n79 Transmission_Gate_Layout_10.VIN.n78 0.7285
R8845 Transmission_Gate_Layout_10.VIN.n77 Transmission_Gate_Layout_10.VIN.t24 0.7285
R8846 Transmission_Gate_Layout_10.VIN.n77 Transmission_Gate_Layout_10.VIN.n76 0.7285
R8847 Transmission_Gate_Layout_10.VIN.n74 Transmission_Gate_Layout_10.VIN.t36 0.7285
R8848 Transmission_Gate_Layout_10.VIN.n74 Transmission_Gate_Layout_10.VIN.n73 0.7285
R8849 Transmission_Gate_Layout_10.VIN.n71 Transmission_Gate_Layout_10.VIN.t28 0.7285
R8850 Transmission_Gate_Layout_10.VIN.n71 Transmission_Gate_Layout_10.VIN.n70 0.7285
R8851 Transmission_Gate_Layout_10.VIN.n69 Transmission_Gate_Layout_10.VIN.t45 0.7285
R8852 Transmission_Gate_Layout_10.VIN.n69 Transmission_Gate_Layout_10.VIN.n68 0.7285
R8853 Transmission_Gate_Layout_10.VIN.n97 Transmission_Gate_Layout_10.VIN.t25 0.7285
R8854 Transmission_Gate_Layout_10.VIN.n97 Transmission_Gate_Layout_10.VIN.n96 0.7285
R8855 Transmission_Gate_Layout_10.VIN.n99 Transmission_Gate_Layout_10.VIN.t32 0.7285
R8856 Transmission_Gate_Layout_10.VIN.n99 Transmission_Gate_Layout_10.VIN.n98 0.7285
R8857 Transmission_Gate_Layout_10.VIN.n101 Transmission_Gate_Layout_10.VIN.t41 0.7285
R8858 Transmission_Gate_Layout_10.VIN.n101 Transmission_Gate_Layout_10.VIN.n100 0.7285
R8859 Transmission_Gate_Layout_10.VIN.n17 Transmission_Gate_Layout_10.VIN.t17 0.7285
R8860 Transmission_Gate_Layout_10.VIN.n17 Transmission_Gate_Layout_10.VIN.n16 0.7285
R8861 Transmission_Gate_Layout_10.VIN.n14 Transmission_Gate_Layout_10.VIN.t4 0.7285
R8862 Transmission_Gate_Layout_10.VIN.n14 Transmission_Gate_Layout_10.VIN.n13 0.7285
R8863 Transmission_Gate_Layout_10.VIN.n12 Transmission_Gate_Layout_10.VIN.t7 0.7285
R8864 Transmission_Gate_Layout_10.VIN.n12 Transmission_Gate_Layout_10.VIN.n11 0.7285
R8865 Transmission_Gate_Layout_10.VIN.n137 Transmission_Gate_Layout_10.VIN.t9 0.7285
R8866 Transmission_Gate_Layout_10.VIN.n137 Transmission_Gate_Layout_10.VIN.n136 0.7285
R8867 Transmission_Gate_Layout_10.VIN.n105 Transmission_Gate_Layout_10.VIN.n104 0.626587
R8868 Transmission_Gate_Layout_10.VIN.n125 Transmission_Gate_Layout_10.VIN.n124 0.626587
R8869 Transmission_Gate_Layout_10.VIN.n127 Transmission_Gate_Layout_10.VIN.n126 0.626587
R8870 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.VIN.n142 0.607022
R8871 Transmission_Gate_Layout_10.VIN.n127 Transmission_Gate_Layout_10.VIN.n10 0.575717
R8872 Transmission_Gate_Layout_10.VIN.n84 Transmission_Gate_Layout_10.VIN.n75 0.575717
R8873 Transmission_Gate_Layout_10.VIN.n126 Transmission_Gate_Layout_10.VIN.n18 0.575717
R8874 Transmission_Gate_Layout_10.VIN.n139 Transmission_Gate_Layout_10.VIN.n138 0.575717
R8875 Transmission_Gate_Layout_10.VIN.n118 Transmission_Gate_Layout_10.VIN.n109 0.570002
R8876 Transmission_Gate_Layout_10.VIN.n120 Transmission_Gate_Layout_10.VIN.n119 0.553423
R8877 Transmission_Gate_Layout_10.VIN.n104 Transmission_Gate_Layout_10.VIN.n95 0.428978
R8878 Transmission_Gate_Layout_10.VIN.n106 Transmission_Gate_Layout_10.VIN.n105 0.428978
R8879 Transmission_Gate_Layout_10.VIN.n119 Transmission_Gate_Layout_10.VIN.n47 0.344848
R8880 Transmission_Gate_Layout_10.VIN.n125 Transmission_Gate_Layout_10.VIN.n26 0.331152
R8881 Transmission_Gate_Layout_10.VIN.n124 Transmission_Gate_Layout_10.VIN.n34 0.331152
R8882 Transmission_Gate_Layout_10.VIN.n120 Transmission_Gate_Layout_10.VIN.n45 0.331152
R8883 Transmission_Gate_Layout_10.VIN.n109 Transmission_Gate_Layout_10.VIN.n55 0.331152
R8884 Transmission_Gate_Layout_10.VIN.n118 Transmission_Gate_Layout_10.VIN.n117 0.317457
R8885 Transmission_Gate_Layout_10.VIN.n126 Transmission_Gate_Layout_10.VIN.n125 0.239196
R8886 Transmission_Gate_Layout_10.VIN.n104 Transmission_Gate_Layout_10.VIN 0.192239
R8887 Transmission_Gate_Layout_9.CLKB.n27 Transmission_Gate_Layout_9.CLKB.t10 54.5477
R8888 Transmission_Gate_Layout_9.CLKB.n27 Transmission_Gate_Layout_9.CLKB.t27 38.3255
R8889 Transmission_Gate_Layout_9.CLKB.n28 Transmission_Gate_Layout_9.CLKB.t7 38.3255
R8890 Transmission_Gate_Layout_9.CLKB.n29 Transmission_Gate_Layout_9.CLKB.t13 38.3255
R8891 Transmission_Gate_Layout_9.CLKB.n30 Transmission_Gate_Layout_9.CLKB.t24 38.3255
R8892 Transmission_Gate_Layout_9.CLKB.n31 Transmission_Gate_Layout_9.CLKB.t6 38.3255
R8893 Transmission_Gate_Layout_9.CLKB.n32 Transmission_Gate_Layout_9.CLKB.t20 38.3255
R8894 Transmission_Gate_Layout_9.CLKB.t12 Transmission_Gate_Layout_9.CLKB.n24 37.9344
R8895 Transmission_Gate_Layout_9.CLKB.t16 Transmission_Gate_Layout_9.CLKB.n23 37.9344
R8896 Transmission_Gate_Layout_9.CLKB.t9 Transmission_Gate_Layout_9.CLKB.n20 37.9344
R8897 Transmission_Gate_Layout_9.CLKB.t15 Transmission_Gate_Layout_9.CLKB.n17 37.9344
R8898 Transmission_Gate_Layout_9.CLKB.t19 Transmission_Gate_Layout_9.CLKB.n14 37.9344
R8899 Transmission_Gate_Layout_9.CLKB.t8 Transmission_Gate_Layout_9.CLKB.n11 37.9344
R8900 Transmission_Gate_Layout_9.CLKB.t14 Transmission_Gate_Layout_9.CLKB.n8 37.9344
R8901 Transmission_Gate_Layout_9.CLKB.t26 Transmission_Gate_Layout_9.CLKB.n5 37.9344
R8902 Transmission_Gate_Layout_9.CLKB.n25 Transmission_Gate_Layout_9.CLKB.t12 37.5434
R8903 Transmission_Gate_Layout_9.CLKB.n26 Transmission_Gate_Layout_9.CLKB.t16 37.5434
R8904 Transmission_Gate_Layout_9.CLKB.n21 Transmission_Gate_Layout_9.CLKB.t9 37.5434
R8905 Transmission_Gate_Layout_9.CLKB.n18 Transmission_Gate_Layout_9.CLKB.t15 37.5434
R8906 Transmission_Gate_Layout_9.CLKB.n15 Transmission_Gate_Layout_9.CLKB.t19 37.5434
R8907 Transmission_Gate_Layout_9.CLKB.n12 Transmission_Gate_Layout_9.CLKB.t8 37.5434
R8908 Transmission_Gate_Layout_9.CLKB.n9 Transmission_Gate_Layout_9.CLKB.t14 37.5434
R8909 Transmission_Gate_Layout_9.CLKB.n6 Transmission_Gate_Layout_9.CLKB.t26 37.5434
R8910 Transmission_Gate_Layout_9.CLKB.n25 Transmission_Gate_Layout_9.CLKB.t29 37.413
R8911 Transmission_Gate_Layout_9.CLKB.t27 Transmission_Gate_Layout_9.CLKB.n21 37.413
R8912 Transmission_Gate_Layout_9.CLKB.t7 Transmission_Gate_Layout_9.CLKB.n18 37.413
R8913 Transmission_Gate_Layout_9.CLKB.t13 Transmission_Gate_Layout_9.CLKB.n15 37.413
R8914 Transmission_Gate_Layout_9.CLKB.t24 Transmission_Gate_Layout_9.CLKB.n12 37.413
R8915 Transmission_Gate_Layout_9.CLKB.t6 Transmission_Gate_Layout_9.CLKB.n9 37.413
R8916 Transmission_Gate_Layout_9.CLKB.t20 Transmission_Gate_Layout_9.CLKB.n6 37.413
R8917 Transmission_Gate_Layout_9.CLKB.t10 Transmission_Gate_Layout_9.CLKB.n26 37.413
R8918 Transmission_Gate_Layout_9.CLKB.n24 Transmission_Gate_Layout_9.CLKB.t21 37.0219
R8919 Transmission_Gate_Layout_9.CLKB.n23 Transmission_Gate_Layout_9.CLKB.t25 37.0219
R8920 Transmission_Gate_Layout_9.CLKB.n20 Transmission_Gate_Layout_9.CLKB.t18 37.0219
R8921 Transmission_Gate_Layout_9.CLKB.n17 Transmission_Gate_Layout_9.CLKB.t23 37.0219
R8922 Transmission_Gate_Layout_9.CLKB.n14 Transmission_Gate_Layout_9.CLKB.t28 37.0219
R8923 Transmission_Gate_Layout_9.CLKB.n11 Transmission_Gate_Layout_9.CLKB.t17 37.0219
R8924 Transmission_Gate_Layout_9.CLKB.n5 Transmission_Gate_Layout_9.CLKB.t11 37.0219
R8925 Transmission_Gate_Layout_9.CLKB.n8 Transmission_Gate_Layout_9.CLKB.t22 37.0219
R8926 Transmission_Gate_Layout_9.CLKB.t25 Transmission_Gate_Layout_9.CLKB.n22 35.1969
R8927 Transmission_Gate_Layout_9.CLKB.t18 Transmission_Gate_Layout_9.CLKB.n19 35.1969
R8928 Transmission_Gate_Layout_9.CLKB.t23 Transmission_Gate_Layout_9.CLKB.n16 35.1969
R8929 Transmission_Gate_Layout_9.CLKB.t28 Transmission_Gate_Layout_9.CLKB.n13 35.1969
R8930 Transmission_Gate_Layout_9.CLKB.t17 Transmission_Gate_Layout_9.CLKB.n10 35.1969
R8931 Transmission_Gate_Layout_9.CLKB.t22 Transmission_Gate_Layout_9.CLKB.n7 35.1969
R8932 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLKB.n32 26.6826
R8933 Transmission_Gate_Layout_9.CLKB.n26 Transmission_Gate_Layout_9.CLKB.n25 19.148
R8934 Transmission_Gate_Layout_9.CLKB.n28 Transmission_Gate_Layout_9.CLKB.n27 16.2227
R8935 Transmission_Gate_Layout_9.CLKB.n29 Transmission_Gate_Layout_9.CLKB.n28 16.2227
R8936 Transmission_Gate_Layout_9.CLKB.n30 Transmission_Gate_Layout_9.CLKB.n29 16.2227
R8937 Transmission_Gate_Layout_9.CLKB.n31 Transmission_Gate_Layout_9.CLKB.n30 16.2227
R8938 Transmission_Gate_Layout_9.CLKB.n32 Transmission_Gate_Layout_9.CLKB.n31 16.2227
R8939 Transmission_Gate_Layout_9.CLKB.n2 Transmission_Gate_Layout_9.CLKB.n0 5.21612
R8940 Transmission_Gate_Layout_9.CLKB.n36 Transmission_Gate_Layout_9.CLKB.n34 4.57285
R8941 Transmission_Gate_Layout_9.CLKB.n2 Transmission_Gate_Layout_9.CLKB.n1 4.4609
R8942 Transmission_Gate_Layout_9.CLKB.n4 Transmission_Gate_Layout_9.CLKB.n3 4.4609
R8943 Transmission_Gate_Layout_9.CLKB.n37 Transmission_Gate_Layout_9.CLKB.n33 3.3285
R8944 Transmission_Gate_Layout_9.CLKB.n36 Transmission_Gate_Layout_9.CLKB.n35 3.3285
R8945 Transmission_Gate_Layout_9.CLKB.n37 Transmission_Gate_Layout_9.CLKB.n36 1.24485
R8946 Transmission_Gate_Layout_9.CLKB.n4 Transmission_Gate_Layout_9.CLKB.n2 0.755717
R8947 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLKB.n37 0.750969
R8948 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.CLKB.n4 0.510317
R8949 Transmission_Gate_Layout_9.VIN.n105 Transmission_Gate_Layout_9.VIN.n104 15.5517
R8950 Transmission_Gate_Layout_9.VIN.n68 Transmission_Gate_Layout_9.VIN.n67 5.21612
R8951 Transmission_Gate_Layout_9.VIN.n71 Transmission_Gate_Layout_9.VIN.t49 4.4609
R8952 Transmission_Gate_Layout_9.VIN.n72 Transmission_Gate_Layout_9.VIN.t58 4.4609
R8953 Transmission_Gate_Layout_9.VIN.n73 Transmission_Gate_Layout_9.VIN.t55 4.4609
R8954 Transmission_Gate_Layout_9.VIN.n69 Transmission_Gate_Layout_9.VIN.n65 4.4609
R8955 Transmission_Gate_Layout_9.VIN.n68 Transmission_Gate_Layout_9.VIN.n66 4.4609
R8956 Transmission_Gate_Layout_9.VIN.n45 Transmission_Gate_Layout_9.VIN.n42 3.90572
R8957 Transmission_Gate_Layout_9.VIN.n53 Transmission_Gate_Layout_9.VIN.n50 3.90572
R8958 Transmission_Gate_Layout_9.VIN.n63 Transmission_Gate_Layout_9.VIN.n62 3.90572
R8959 Transmission_Gate_Layout_9.VIN.n30 Transmission_Gate_Layout_9.VIN.n29 3.90572
R8960 Transmission_Gate_Layout_9.VIN.n22 Transmission_Gate_Layout_9.VIN.n21 3.90572
R8961 Transmission_Gate_Layout_9.VIN.n4 Transmission_Gate_Layout_9.VIN.n1 3.90572
R8962 Transmission_Gate_Layout_9.VIN.n93 Transmission_Gate_Layout_9.VIN.n90 3.84485
R8963 Transmission_Gate_Layout_9.VIN.n82 Transmission_Gate_Layout_9.VIN.n81 3.84485
R8964 Transmission_Gate_Layout_9.VIN.n39 Transmission_Gate_Layout_9.VIN.n38 3.84485
R8965 Transmission_Gate_Layout_9.VIN.n14 Transmission_Gate_Layout_9.VIN.n13 3.84485
R8966 Transmission_Gate_Layout_9.VIN.n125 Transmission_Gate_Layout_9.VIN.n122 3.84485
R8967 Transmission_Gate_Layout_9.VIN.n133 Transmission_Gate_Layout_9.VIN.n130 3.84485
R8968 Transmission_Gate_Layout_9.VIN.n102 Transmission_Gate_Layout_9.VIN.n101 3.3285
R8969 Transmission_Gate_Layout_9.VIN.n100 Transmission_Gate_Layout_9.VIN.n99 3.3285
R8970 Transmission_Gate_Layout_9.VIN.n98 Transmission_Gate_Layout_9.VIN.n97 3.3285
R8971 Transmission_Gate_Layout_9.VIN.n86 Transmission_Gate_Layout_9.VIN.t87 3.3285
R8972 Transmission_Gate_Layout_9.VIN.n87 Transmission_Gate_Layout_9.VIN.t78 3.3285
R8973 Transmission_Gate_Layout_9.VIN.n88 Transmission_Gate_Layout_9.VIN.t84 3.3285
R8974 Transmission_Gate_Layout_9.VIN.n45 Transmission_Gate_Layout_9.VIN.n44 3.1505
R8975 Transmission_Gate_Layout_9.VIN.n48 Transmission_Gate_Layout_9.VIN.n47 3.1505
R8976 Transmission_Gate_Layout_9.VIN.n53 Transmission_Gate_Layout_9.VIN.n52 3.1505
R8977 Transmission_Gate_Layout_9.VIN.n56 Transmission_Gate_Layout_9.VIN.n55 3.1505
R8978 Transmission_Gate_Layout_9.VIN.n63 Transmission_Gate_Layout_9.VIN.n60 3.1505
R8979 Transmission_Gate_Layout_9.VIN.n64 Transmission_Gate_Layout_9.VIN.n58 3.1505
R8980 Transmission_Gate_Layout_9.VIN.n30 Transmission_Gate_Layout_9.VIN.n27 3.1505
R8981 Transmission_Gate_Layout_9.VIN.n31 Transmission_Gate_Layout_9.VIN.n25 3.1505
R8982 Transmission_Gate_Layout_9.VIN.n22 Transmission_Gate_Layout_9.VIN.n19 3.1505
R8983 Transmission_Gate_Layout_9.VIN.n23 Transmission_Gate_Layout_9.VIN.n17 3.1505
R8984 Transmission_Gate_Layout_9.VIN.n114 Transmission_Gate_Layout_9.VIN.n113 3.1505
R8985 Transmission_Gate_Layout_9.VIN.n111 Transmission_Gate_Layout_9.VIN.n110 3.1505
R8986 Transmission_Gate_Layout_9.VIN.n108 Transmission_Gate_Layout_9.VIN.n107 3.1505
R8987 Transmission_Gate_Layout_9.VIN.n4 Transmission_Gate_Layout_9.VIN.n3 3.1505
R8988 Transmission_Gate_Layout_9.VIN.n7 Transmission_Gate_Layout_9.VIN.n6 3.1505
R8989 Transmission_Gate_Layout_9.VIN.n93 Transmission_Gate_Layout_9.VIN.n92 2.6005
R8990 Transmission_Gate_Layout_9.VIN.n96 Transmission_Gate_Layout_9.VIN.n95 2.6005
R8991 Transmission_Gate_Layout_9.VIN.n82 Transmission_Gate_Layout_9.VIN.n79 2.6005
R8992 Transmission_Gate_Layout_9.VIN.n83 Transmission_Gate_Layout_9.VIN.n77 2.6005
R8993 Transmission_Gate_Layout_9.VIN.n39 Transmission_Gate_Layout_9.VIN.n36 2.6005
R8994 Transmission_Gate_Layout_9.VIN.n40 Transmission_Gate_Layout_9.VIN.n34 2.6005
R8995 Transmission_Gate_Layout_9.VIN.n14 Transmission_Gate_Layout_9.VIN.n11 2.6005
R8996 Transmission_Gate_Layout_9.VIN.n15 Transmission_Gate_Layout_9.VIN.n9 2.6005
R8997 Transmission_Gate_Layout_9.VIN.n138 Transmission_Gate_Layout_9.VIN.n120 2.6005
R8998 Transmission_Gate_Layout_9.VIN.n139 Transmission_Gate_Layout_9.VIN.n118 2.6005
R8999 Transmission_Gate_Layout_9.VIN.n140 Transmission_Gate_Layout_9.VIN.n116 2.6005
R9000 Transmission_Gate_Layout_9.VIN.n125 Transmission_Gate_Layout_9.VIN.n124 2.6005
R9001 Transmission_Gate_Layout_9.VIN.n128 Transmission_Gate_Layout_9.VIN.n127 2.6005
R9002 Transmission_Gate_Layout_9.VIN.n133 Transmission_Gate_Layout_9.VIN.n132 2.6005
R9003 Transmission_Gate_Layout_9.VIN.n136 Transmission_Gate_Layout_9.VIN.n135 2.6005
R9004 Transmission_Gate_Layout_9.VIN.n71 Transmission_Gate_Layout_9.VIN.n70 2.47941
R9005 Transmission_Gate_Layout_9.VIN.n104 Transmission_Gate_Layout_9.VIN.n103 1.90239
R9006 Transmission_Gate_Layout_9.VIN.n107 Transmission_Gate_Layout_9.VIN.t28 1.3109
R9007 Transmission_Gate_Layout_9.VIN.n107 Transmission_Gate_Layout_9.VIN.n106 1.3109
R9008 Transmission_Gate_Layout_9.VIN.n110 Transmission_Gate_Layout_9.VIN.t34 1.3109
R9009 Transmission_Gate_Layout_9.VIN.n110 Transmission_Gate_Layout_9.VIN.n109 1.3109
R9010 Transmission_Gate_Layout_9.VIN.n113 Transmission_Gate_Layout_9.VIN.t42 1.3109
R9011 Transmission_Gate_Layout_9.VIN.n113 Transmission_Gate_Layout_9.VIN.n112 1.3109
R9012 Transmission_Gate_Layout_9.VIN.n47 Transmission_Gate_Layout_9.VIN.t59 1.3109
R9013 Transmission_Gate_Layout_9.VIN.n47 Transmission_Gate_Layout_9.VIN.n46 1.3109
R9014 Transmission_Gate_Layout_9.VIN.n44 Transmission_Gate_Layout_9.VIN.t50 1.3109
R9015 Transmission_Gate_Layout_9.VIN.n44 Transmission_Gate_Layout_9.VIN.n43 1.3109
R9016 Transmission_Gate_Layout_9.VIN.n42 Transmission_Gate_Layout_9.VIN.t52 1.3109
R9017 Transmission_Gate_Layout_9.VIN.n42 Transmission_Gate_Layout_9.VIN.n41 1.3109
R9018 Transmission_Gate_Layout_9.VIN.n55 Transmission_Gate_Layout_9.VIN.t54 1.3109
R9019 Transmission_Gate_Layout_9.VIN.n55 Transmission_Gate_Layout_9.VIN.n54 1.3109
R9020 Transmission_Gate_Layout_9.VIN.n52 Transmission_Gate_Layout_9.VIN.t57 1.3109
R9021 Transmission_Gate_Layout_9.VIN.n52 Transmission_Gate_Layout_9.VIN.n51 1.3109
R9022 Transmission_Gate_Layout_9.VIN.n50 Transmission_Gate_Layout_9.VIN.t48 1.3109
R9023 Transmission_Gate_Layout_9.VIN.n50 Transmission_Gate_Layout_9.VIN.n49 1.3109
R9024 Transmission_Gate_Layout_9.VIN.n58 Transmission_Gate_Layout_9.VIN.t56 1.3109
R9025 Transmission_Gate_Layout_9.VIN.n58 Transmission_Gate_Layout_9.VIN.n57 1.3109
R9026 Transmission_Gate_Layout_9.VIN.n60 Transmission_Gate_Layout_9.VIN.t53 1.3109
R9027 Transmission_Gate_Layout_9.VIN.n60 Transmission_Gate_Layout_9.VIN.n59 1.3109
R9028 Transmission_Gate_Layout_9.VIN.n62 Transmission_Gate_Layout_9.VIN.t51 1.3109
R9029 Transmission_Gate_Layout_9.VIN.n62 Transmission_Gate_Layout_9.VIN.n61 1.3109
R9030 Transmission_Gate_Layout_9.VIN.n25 Transmission_Gate_Layout_9.VIN.t31 1.3109
R9031 Transmission_Gate_Layout_9.VIN.n25 Transmission_Gate_Layout_9.VIN.n24 1.3109
R9032 Transmission_Gate_Layout_9.VIN.n27 Transmission_Gate_Layout_9.VIN.t39 1.3109
R9033 Transmission_Gate_Layout_9.VIN.n27 Transmission_Gate_Layout_9.VIN.n26 1.3109
R9034 Transmission_Gate_Layout_9.VIN.n29 Transmission_Gate_Layout_9.VIN.t36 1.3109
R9035 Transmission_Gate_Layout_9.VIN.n29 Transmission_Gate_Layout_9.VIN.n28 1.3109
R9036 Transmission_Gate_Layout_9.VIN.n17 Transmission_Gate_Layout_9.VIN.t41 1.3109
R9037 Transmission_Gate_Layout_9.VIN.n17 Transmission_Gate_Layout_9.VIN.n16 1.3109
R9038 Transmission_Gate_Layout_9.VIN.n19 Transmission_Gate_Layout_9.VIN.t46 1.3109
R9039 Transmission_Gate_Layout_9.VIN.n19 Transmission_Gate_Layout_9.VIN.n18 1.3109
R9040 Transmission_Gate_Layout_9.VIN.n21 Transmission_Gate_Layout_9.VIN.t30 1.3109
R9041 Transmission_Gate_Layout_9.VIN.n21 Transmission_Gate_Layout_9.VIN.n20 1.3109
R9042 Transmission_Gate_Layout_9.VIN.n6 Transmission_Gate_Layout_9.VIN.t38 1.3109
R9043 Transmission_Gate_Layout_9.VIN.n6 Transmission_Gate_Layout_9.VIN.n5 1.3109
R9044 Transmission_Gate_Layout_9.VIN.n3 Transmission_Gate_Layout_9.VIN.t33 1.3109
R9045 Transmission_Gate_Layout_9.VIN.n3 Transmission_Gate_Layout_9.VIN.n2 1.3109
R9046 Transmission_Gate_Layout_9.VIN.n1 Transmission_Gate_Layout_9.VIN.t26 1.3109
R9047 Transmission_Gate_Layout_9.VIN.n1 Transmission_Gate_Layout_9.VIN.n0 1.3109
R9048 Transmission_Gate_Layout_9.VIN.n96 Transmission_Gate_Layout_9.VIN.n93 1.24485
R9049 Transmission_Gate_Layout_9.VIN.n100 Transmission_Gate_Layout_9.VIN.n98 1.24485
R9050 Transmission_Gate_Layout_9.VIN.n102 Transmission_Gate_Layout_9.VIN.n100 1.24485
R9051 Transmission_Gate_Layout_9.VIN.n83 Transmission_Gate_Layout_9.VIN.n82 1.24485
R9052 Transmission_Gate_Layout_9.VIN.n40 Transmission_Gate_Layout_9.VIN.n39 1.24485
R9053 Transmission_Gate_Layout_9.VIN.n87 Transmission_Gate_Layout_9.VIN.n86 1.24485
R9054 Transmission_Gate_Layout_9.VIN.n88 Transmission_Gate_Layout_9.VIN.n87 1.24485
R9055 Transmission_Gate_Layout_9.VIN.n15 Transmission_Gate_Layout_9.VIN.n14 1.24485
R9056 Transmission_Gate_Layout_9.VIN.n140 Transmission_Gate_Layout_9.VIN.n139 1.24485
R9057 Transmission_Gate_Layout_9.VIN.n139 Transmission_Gate_Layout_9.VIN.n138 1.24485
R9058 Transmission_Gate_Layout_9.VIN.n128 Transmission_Gate_Layout_9.VIN.n125 1.24485
R9059 Transmission_Gate_Layout_9.VIN.n136 Transmission_Gate_Layout_9.VIN.n133 1.24485
R9060 Transmission_Gate_Layout_9.VIN.n103 Transmission_Gate_Layout_9.VIN.n102 1.2018
R9061 Transmission_Gate_Layout_9.VIN.n86 Transmission_Gate_Layout_9.VIN.n85 1.2018
R9062 Transmission_Gate_Layout_9.VIN.n138 Transmission_Gate_Layout_9.VIN.n137 1.2018
R9063 Transmission_Gate_Layout_9.VIN.n137 Transmission_Gate_Layout_9.VIN.n136 1.2018
R9064 Transmission_Gate_Layout_9.VIN.n70 Transmission_Gate_Layout_9.VIN.n69 0.957239
R9065 Transmission_Gate_Layout_9.VIN.n74 Transmission_Gate_Layout_9.VIN.n73 0.957239
R9066 Transmission_Gate_Layout_9.VIN.n32 Transmission_Gate_Layout_9.VIN.n31 0.957239
R9067 Transmission_Gate_Layout_9.VIN.n142 Transmission_Gate_Layout_9.VIN.n15 0.806587
R9068 Transmission_Gate_Layout_9.VIN.n141 Transmission_Gate_Layout_9.VIN.n140 0.806587
R9069 Transmission_Gate_Layout_9.VIN.n48 Transmission_Gate_Layout_9.VIN.n45 0.755717
R9070 Transmission_Gate_Layout_9.VIN.n56 Transmission_Gate_Layout_9.VIN.n53 0.755717
R9071 Transmission_Gate_Layout_9.VIN.n64 Transmission_Gate_Layout_9.VIN.n63 0.755717
R9072 Transmission_Gate_Layout_9.VIN.n69 Transmission_Gate_Layout_9.VIN.n68 0.755717
R9073 Transmission_Gate_Layout_9.VIN.n72 Transmission_Gate_Layout_9.VIN.n71 0.755717
R9074 Transmission_Gate_Layout_9.VIN.n73 Transmission_Gate_Layout_9.VIN.n72 0.755717
R9075 Transmission_Gate_Layout_9.VIN.n31 Transmission_Gate_Layout_9.VIN.n30 0.755717
R9076 Transmission_Gate_Layout_9.VIN.n23 Transmission_Gate_Layout_9.VIN.n22 0.755717
R9077 Transmission_Gate_Layout_9.VIN.n111 Transmission_Gate_Layout_9.VIN.n108 0.755717
R9078 Transmission_Gate_Layout_9.VIN.n114 Transmission_Gate_Layout_9.VIN.n111 0.755717
R9079 Transmission_Gate_Layout_9.VIN.n7 Transmission_Gate_Layout_9.VIN.n4 0.755717
R9080 Transmission_Gate_Layout_9.VIN.n104 Transmission_Gate_Layout_9.VIN.n88 0.742022
R9081 Transmission_Gate_Layout_9.VIN.n135 Transmission_Gate_Layout_9.VIN.t7 0.7285
R9082 Transmission_Gate_Layout_9.VIN.n135 Transmission_Gate_Layout_9.VIN.n134 0.7285
R9083 Transmission_Gate_Layout_9.VIN.n132 Transmission_Gate_Layout_9.VIN.t15 0.7285
R9084 Transmission_Gate_Layout_9.VIN.n132 Transmission_Gate_Layout_9.VIN.n131 0.7285
R9085 Transmission_Gate_Layout_9.VIN.n116 Transmission_Gate_Layout_9.VIN.t2 0.7285
R9086 Transmission_Gate_Layout_9.VIN.n116 Transmission_Gate_Layout_9.VIN.n115 0.7285
R9087 Transmission_Gate_Layout_9.VIN.n118 Transmission_Gate_Layout_9.VIN.t20 0.7285
R9088 Transmission_Gate_Layout_9.VIN.n118 Transmission_Gate_Layout_9.VIN.n117 0.7285
R9089 Transmission_Gate_Layout_9.VIN.n120 Transmission_Gate_Layout_9.VIN.t11 0.7285
R9090 Transmission_Gate_Layout_9.VIN.n120 Transmission_Gate_Layout_9.VIN.n119 0.7285
R9091 Transmission_Gate_Layout_9.VIN.n95 Transmission_Gate_Layout_9.VIN.t80 0.7285
R9092 Transmission_Gate_Layout_9.VIN.n95 Transmission_Gate_Layout_9.VIN.n94 0.7285
R9093 Transmission_Gate_Layout_9.VIN.n92 Transmission_Gate_Layout_9.VIN.t85 0.7285
R9094 Transmission_Gate_Layout_9.VIN.n92 Transmission_Gate_Layout_9.VIN.n91 0.7285
R9095 Transmission_Gate_Layout_9.VIN.n90 Transmission_Gate_Layout_9.VIN.t82 0.7285
R9096 Transmission_Gate_Layout_9.VIN.n90 Transmission_Gate_Layout_9.VIN.n89 0.7285
R9097 Transmission_Gate_Layout_9.VIN.n77 Transmission_Gate_Layout_9.VIN.t79 0.7285
R9098 Transmission_Gate_Layout_9.VIN.n77 Transmission_Gate_Layout_9.VIN.n76 0.7285
R9099 Transmission_Gate_Layout_9.VIN.n79 Transmission_Gate_Layout_9.VIN.t81 0.7285
R9100 Transmission_Gate_Layout_9.VIN.n79 Transmission_Gate_Layout_9.VIN.n78 0.7285
R9101 Transmission_Gate_Layout_9.VIN.n81 Transmission_Gate_Layout_9.VIN.t76 0.7285
R9102 Transmission_Gate_Layout_9.VIN.n81 Transmission_Gate_Layout_9.VIN.n80 0.7285
R9103 Transmission_Gate_Layout_9.VIN.n34 Transmission_Gate_Layout_9.VIN.t86 0.7285
R9104 Transmission_Gate_Layout_9.VIN.n34 Transmission_Gate_Layout_9.VIN.n33 0.7285
R9105 Transmission_Gate_Layout_9.VIN.n36 Transmission_Gate_Layout_9.VIN.t77 0.7285
R9106 Transmission_Gate_Layout_9.VIN.n36 Transmission_Gate_Layout_9.VIN.n35 0.7285
R9107 Transmission_Gate_Layout_9.VIN.n38 Transmission_Gate_Layout_9.VIN.t83 0.7285
R9108 Transmission_Gate_Layout_9.VIN.n38 Transmission_Gate_Layout_9.VIN.n37 0.7285
R9109 Transmission_Gate_Layout_9.VIN.n9 Transmission_Gate_Layout_9.VIN.t0 0.7285
R9110 Transmission_Gate_Layout_9.VIN.n9 Transmission_Gate_Layout_9.VIN.n8 0.7285
R9111 Transmission_Gate_Layout_9.VIN.n11 Transmission_Gate_Layout_9.VIN.t17 0.7285
R9112 Transmission_Gate_Layout_9.VIN.n11 Transmission_Gate_Layout_9.VIN.n10 0.7285
R9113 Transmission_Gate_Layout_9.VIN.n13 Transmission_Gate_Layout_9.VIN.t8 0.7285
R9114 Transmission_Gate_Layout_9.VIN.n13 Transmission_Gate_Layout_9.VIN.n12 0.7285
R9115 Transmission_Gate_Layout_9.VIN.n127 Transmission_Gate_Layout_9.VIN.t1 0.7285
R9116 Transmission_Gate_Layout_9.VIN.n127 Transmission_Gate_Layout_9.VIN.n126 0.7285
R9117 Transmission_Gate_Layout_9.VIN.n124 Transmission_Gate_Layout_9.VIN.t10 0.7285
R9118 Transmission_Gate_Layout_9.VIN.n124 Transmission_Gate_Layout_9.VIN.n123 0.7285
R9119 Transmission_Gate_Layout_9.VIN.n122 Transmission_Gate_Layout_9.VIN.t16 0.7285
R9120 Transmission_Gate_Layout_9.VIN.n122 Transmission_Gate_Layout_9.VIN.n121 0.7285
R9121 Transmission_Gate_Layout_9.VIN.n130 Transmission_Gate_Layout_9.VIN.t23 0.7285
R9122 Transmission_Gate_Layout_9.VIN.n130 Transmission_Gate_Layout_9.VIN.n129 0.7285
R9123 Transmission_Gate_Layout_9.VIN.n75 Transmission_Gate_Layout_9.VIN.n74 0.626587
R9124 Transmission_Gate_Layout_9.VIN.n85 Transmission_Gate_Layout_9.VIN.n84 0.626587
R9125 Transmission_Gate_Layout_9.VIN.n142 Transmission_Gate_Layout_9.VIN.n141 0.626587
R9126 Transmission_Gate_Layout_9.VIN.n98 Transmission_Gate_Layout_9.VIN 0.607022
R9127 Transmission_Gate_Layout_9.VIN.n103 Transmission_Gate_Layout_9.VIN.n96 0.575717
R9128 Transmission_Gate_Layout_9.VIN.n84 Transmission_Gate_Layout_9.VIN.n83 0.575717
R9129 Transmission_Gate_Layout_9.VIN.n85 Transmission_Gate_Layout_9.VIN.n40 0.575717
R9130 Transmission_Gate_Layout_9.VIN.n137 Transmission_Gate_Layout_9.VIN.n128 0.575717
R9131 Transmission_Gate_Layout_9.VIN.n105 Transmission_Gate_Layout_9.VIN.n32 0.570002
R9132 Transmission_Gate_Layout_9.VIN.n141 Transmission_Gate_Layout_9.VIN.n114 0.428978
R9133 Transmission_Gate_Layout_9.VIN.n142 Transmission_Gate_Layout_9.VIN.n7 0.428978
R9134 Transmission_Gate_Layout_9.VIN.n75 Transmission_Gate_Layout_9.VIN.n48 0.331152
R9135 Transmission_Gate_Layout_9.VIN.n74 Transmission_Gate_Layout_9.VIN.n56 0.331152
R9136 Transmission_Gate_Layout_9.VIN.n70 Transmission_Gate_Layout_9.VIN.n64 0.331152
R9137 Transmission_Gate_Layout_9.VIN.n32 Transmission_Gate_Layout_9.VIN.n23 0.331152
R9138 Transmission_Gate_Layout_9.VIN.n108 Transmission_Gate_Layout_9.VIN.n105 0.317457
R9139 Transmission_Gate_Layout_9.VIN.n84 Transmission_Gate_Layout_9.VIN.n75 0.239196
R9140 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.VIN.n142 0.192239
R9141 Transmission_Gate_Layout_6.CLKB.n24 Transmission_Gate_Layout_6.CLKB.t20 54.5477
R9142 Transmission_Gate_Layout_6.CLKB.n29 Transmission_Gate_Layout_6.CLKB.t27 38.3255
R9143 Transmission_Gate_Layout_6.CLKB.n28 Transmission_Gate_Layout_6.CLKB.t24 38.3255
R9144 Transmission_Gate_Layout_6.CLKB.n27 Transmission_Gate_Layout_6.CLKB.t26 38.3255
R9145 Transmission_Gate_Layout_6.CLKB.n26 Transmission_Gate_Layout_6.CLKB.t7 38.3255
R9146 Transmission_Gate_Layout_6.CLKB.n25 Transmission_Gate_Layout_6.CLKB.t13 38.3255
R9147 Transmission_Gate_Layout_6.CLKB.n24 Transmission_Gate_Layout_6.CLKB.t16 38.3255
R9148 Transmission_Gate_Layout_6.CLKB.t11 Transmission_Gate_Layout_6.CLKB.n2 37.9344
R9149 Transmission_Gate_Layout_6.CLKB.t9 Transmission_Gate_Layout_6.CLKB.n5 37.9344
R9150 Transmission_Gate_Layout_6.CLKB.t10 Transmission_Gate_Layout_6.CLKB.n8 37.9344
R9151 Transmission_Gate_Layout_6.CLKB.t19 Transmission_Gate_Layout_6.CLKB.n11 37.9344
R9152 Transmission_Gate_Layout_6.CLKB.t23 Transmission_Gate_Layout_6.CLKB.n14 37.9344
R9153 Transmission_Gate_Layout_6.CLKB.t25 Transmission_Gate_Layout_6.CLKB.n17 37.9344
R9154 Transmission_Gate_Layout_6.CLKB.t6 Transmission_Gate_Layout_6.CLKB.n20 37.9344
R9155 Transmission_Gate_Layout_6.CLKB.t8 Transmission_Gate_Layout_6.CLKB.n21 37.9344
R9156 Transmission_Gate_Layout_6.CLKB.n3 Transmission_Gate_Layout_6.CLKB.t11 37.5434
R9157 Transmission_Gate_Layout_6.CLKB.n6 Transmission_Gate_Layout_6.CLKB.t9 37.5434
R9158 Transmission_Gate_Layout_6.CLKB.n9 Transmission_Gate_Layout_6.CLKB.t10 37.5434
R9159 Transmission_Gate_Layout_6.CLKB.n12 Transmission_Gate_Layout_6.CLKB.t19 37.5434
R9160 Transmission_Gate_Layout_6.CLKB.n15 Transmission_Gate_Layout_6.CLKB.t23 37.5434
R9161 Transmission_Gate_Layout_6.CLKB.n18 Transmission_Gate_Layout_6.CLKB.t25 37.5434
R9162 Transmission_Gate_Layout_6.CLKB.n23 Transmission_Gate_Layout_6.CLKB.t6 37.5434
R9163 Transmission_Gate_Layout_6.CLKB.n22 Transmission_Gate_Layout_6.CLKB.t8 37.5434
R9164 Transmission_Gate_Layout_6.CLKB.t27 Transmission_Gate_Layout_6.CLKB.n3 37.413
R9165 Transmission_Gate_Layout_6.CLKB.t24 Transmission_Gate_Layout_6.CLKB.n6 37.413
R9166 Transmission_Gate_Layout_6.CLKB.t26 Transmission_Gate_Layout_6.CLKB.n9 37.413
R9167 Transmission_Gate_Layout_6.CLKB.t7 Transmission_Gate_Layout_6.CLKB.n12 37.413
R9168 Transmission_Gate_Layout_6.CLKB.t13 Transmission_Gate_Layout_6.CLKB.n15 37.413
R9169 Transmission_Gate_Layout_6.CLKB.t16 Transmission_Gate_Layout_6.CLKB.n18 37.413
R9170 Transmission_Gate_Layout_6.CLKB.n22 Transmission_Gate_Layout_6.CLKB.t22 37.413
R9171 Transmission_Gate_Layout_6.CLKB.t20 Transmission_Gate_Layout_6.CLKB.n23 37.413
R9172 Transmission_Gate_Layout_6.CLKB.n21 Transmission_Gate_Layout_6.CLKB.t14 37.0219
R9173 Transmission_Gate_Layout_6.CLKB.n17 Transmission_Gate_Layout_6.CLKB.t29 37.0219
R9174 Transmission_Gate_Layout_6.CLKB.n14 Transmission_Gate_Layout_6.CLKB.t28 37.0219
R9175 Transmission_Gate_Layout_6.CLKB.n11 Transmission_Gate_Layout_6.CLKB.t21 37.0219
R9176 Transmission_Gate_Layout_6.CLKB.n8 Transmission_Gate_Layout_6.CLKB.t17 37.0219
R9177 Transmission_Gate_Layout_6.CLKB.n5 Transmission_Gate_Layout_6.CLKB.t15 37.0219
R9178 Transmission_Gate_Layout_6.CLKB.n2 Transmission_Gate_Layout_6.CLKB.t18 37.0219
R9179 Transmission_Gate_Layout_6.CLKB.n20 Transmission_Gate_Layout_6.CLKB.t12 37.0219
R9180 Transmission_Gate_Layout_6.CLKB.t29 Transmission_Gate_Layout_6.CLKB.n16 35.1969
R9181 Transmission_Gate_Layout_6.CLKB.t28 Transmission_Gate_Layout_6.CLKB.n13 35.1969
R9182 Transmission_Gate_Layout_6.CLKB.t21 Transmission_Gate_Layout_6.CLKB.n10 35.1969
R9183 Transmission_Gate_Layout_6.CLKB.t17 Transmission_Gate_Layout_6.CLKB.n7 35.1969
R9184 Transmission_Gate_Layout_6.CLKB.t15 Transmission_Gate_Layout_6.CLKB.n4 35.1969
R9185 Transmission_Gate_Layout_6.CLKB.t12 Transmission_Gate_Layout_6.CLKB.n19 35.1969
R9186 Transmission_Gate_Layout_6.CLKB Transmission_Gate_Layout_6.CLKB.n29 26.6826
R9187 Transmission_Gate_Layout_6.CLKB.n23 Transmission_Gate_Layout_6.CLKB.n22 19.148
R9188 Transmission_Gate_Layout_6.CLKB.n29 Transmission_Gate_Layout_6.CLKB.n28 16.2227
R9189 Transmission_Gate_Layout_6.CLKB.n28 Transmission_Gate_Layout_6.CLKB.n27 16.2227
R9190 Transmission_Gate_Layout_6.CLKB.n27 Transmission_Gate_Layout_6.CLKB.n26 16.2227
R9191 Transmission_Gate_Layout_6.CLKB.n26 Transmission_Gate_Layout_6.CLKB.n25 16.2227
R9192 Transmission_Gate_Layout_6.CLKB.n25 Transmission_Gate_Layout_6.CLKB.n24 16.2227
R9193 Transmission_Gate_Layout_6.CLKB.n30 Transmission_Gate_Layout_6.CLKB.t3 5.21612
R9194 Transmission_Gate_Layout_6.CLKB.n0 Transmission_Gate_Layout_6.CLKB.t1 4.57285
R9195 Transmission_Gate_Layout_6.CLKB.n31 Transmission_Gate_Layout_6.CLKB.t5 4.4609
R9196 Transmission_Gate_Layout_6.CLKB.n30 Transmission_Gate_Layout_6.CLKB.t4 4.4609
R9197 Transmission_Gate_Layout_6.CLKB.n1 Transmission_Gate_Layout_6.CLKB.t0 3.3285
R9198 Transmission_Gate_Layout_6.CLKB.n0 Transmission_Gate_Layout_6.CLKB.t2 3.3285
R9199 Transmission_Gate_Layout_6.CLKB.n1 Transmission_Gate_Layout_6.CLKB.n0 1.24485
R9200 Transmission_Gate_Layout_6.CLKB.n31 Transmission_Gate_Layout_6.CLKB.n30 0.755717
R9201 Transmission_Gate_Layout_6.CLKB Transmission_Gate_Layout_6.CLKB.n1 0.750969
R9202 Transmission_Gate_Layout_6.CLKB Transmission_Gate_Layout_6.CLKB.n31 0.510317
R9203 Transmission_Gate_Layout_8.VIN.n104 Transmission_Gate_Layout_8.VIN.n95 7.05901
R9204 Transmission_Gate_Layout_8.VIN.n93 Transmission_Gate_Layout_8.VIN.t86 5.21612
R9205 Transmission_Gate_Layout_8.VIN.n83 Transmission_Gate_Layout_8.VIN.n24 4.4609
R9206 Transmission_Gate_Layout_8.VIN.n82 Transmission_Gate_Layout_8.VIN.n25 4.4609
R9207 Transmission_Gate_Layout_8.VIN.n81 Transmission_Gate_Layout_8.VIN.n26 4.4609
R9208 Transmission_Gate_Layout_8.VIN.n94 Transmission_Gate_Layout_8.VIN.t89 4.4609
R9209 Transmission_Gate_Layout_8.VIN.n93 Transmission_Gate_Layout_8.VIN.t91 4.4609
R9210 Transmission_Gate_Layout_8.VIN.n31 Transmission_Gate_Layout_8.VIN.n28 3.90572
R9211 Transmission_Gate_Layout_8.VIN.n39 Transmission_Gate_Layout_8.VIN.n36 3.90572
R9212 Transmission_Gate_Layout_8.VIN.n90 Transmission_Gate_Layout_8.VIN.n89 3.90572
R9213 Transmission_Gate_Layout_8.VIN.n102 Transmission_Gate_Layout_8.VIN.n101 3.90572
R9214 Transmission_Gate_Layout_8.VIN.n22 Transmission_Gate_Layout_8.VIN.n21 3.90572
R9215 Transmission_Gate_Layout_8.VIN.n4 Transmission_Gate_Layout_8.VIN.n1 3.90572
R9216 Transmission_Gate_Layout_8.VIN.n125 Transmission_Gate_Layout_8.VIN.n122 3.84485
R9217 Transmission_Gate_Layout_8.VIN.n49 Transmission_Gate_Layout_8.VIN.n48 3.84485
R9218 Transmission_Gate_Layout_8.VIN.n57 Transmission_Gate_Layout_8.VIN.n56 3.84485
R9219 Transmission_Gate_Layout_8.VIN.n66 Transmission_Gate_Layout_8.VIN.n63 3.84485
R9220 Transmission_Gate_Layout_8.VIN.n14 Transmission_Gate_Layout_8.VIN.n13 3.84485
R9221 Transmission_Gate_Layout_8.VIN.n133 Transmission_Gate_Layout_8.VIN.n130 3.84485
R9222 Transmission_Gate_Layout_8.VIN.n76 Transmission_Gate_Layout_8.VIN.n59 3.3285
R9223 Transmission_Gate_Layout_8.VIN.n75 Transmission_Gate_Layout_8.VIN.n60 3.3285
R9224 Transmission_Gate_Layout_8.VIN.n74 Transmission_Gate_Layout_8.VIN.n61 3.3285
R9225 Transmission_Gate_Layout_8.VIN.n72 Transmission_Gate_Layout_8.VIN.t10 3.3285
R9226 Transmission_Gate_Layout_8.VIN.n71 Transmission_Gate_Layout_8.VIN.t1 3.3285
R9227 Transmission_Gate_Layout_8.VIN.n70 Transmission_Gate_Layout_8.VIN.t17 3.3285
R9228 Transmission_Gate_Layout_8.VIN.n31 Transmission_Gate_Layout_8.VIN.n30 3.1505
R9229 Transmission_Gate_Layout_8.VIN.n34 Transmission_Gate_Layout_8.VIN.n33 3.1505
R9230 Transmission_Gate_Layout_8.VIN.n39 Transmission_Gate_Layout_8.VIN.n38 3.1505
R9231 Transmission_Gate_Layout_8.VIN.n42 Transmission_Gate_Layout_8.VIN.n41 3.1505
R9232 Transmission_Gate_Layout_8.VIN.n90 Transmission_Gate_Layout_8.VIN.n87 3.1505
R9233 Transmission_Gate_Layout_8.VIN.n91 Transmission_Gate_Layout_8.VIN.n85 3.1505
R9234 Transmission_Gate_Layout_8.VIN.n102 Transmission_Gate_Layout_8.VIN.n99 3.1505
R9235 Transmission_Gate_Layout_8.VIN.n103 Transmission_Gate_Layout_8.VIN.n97 3.1505
R9236 Transmission_Gate_Layout_8.VIN.n22 Transmission_Gate_Layout_8.VIN.n19 3.1505
R9237 Transmission_Gate_Layout_8.VIN.n23 Transmission_Gate_Layout_8.VIN.n17 3.1505
R9238 Transmission_Gate_Layout_8.VIN.n108 Transmission_Gate_Layout_8.VIN.n107 3.1505
R9239 Transmission_Gate_Layout_8.VIN.n111 Transmission_Gate_Layout_8.VIN.n110 3.1505
R9240 Transmission_Gate_Layout_8.VIN.n114 Transmission_Gate_Layout_8.VIN.n113 3.1505
R9241 Transmission_Gate_Layout_8.VIN.n7 Transmission_Gate_Layout_8.VIN.n6 3.1505
R9242 Transmission_Gate_Layout_8.VIN.n4 Transmission_Gate_Layout_8.VIN.n3 3.1505
R9243 Transmission_Gate_Layout_8.VIN.n74 Transmission_Gate_Layout_8.VIN.n73 2.72398
R9244 Transmission_Gate_Layout_8.VIN.n125 Transmission_Gate_Layout_8.VIN.n124 2.6005
R9245 Transmission_Gate_Layout_8.VIN.n128 Transmission_Gate_Layout_8.VIN.n127 2.6005
R9246 Transmission_Gate_Layout_8.VIN.n49 Transmission_Gate_Layout_8.VIN.n46 2.6005
R9247 Transmission_Gate_Layout_8.VIN.n50 Transmission_Gate_Layout_8.VIN.n44 2.6005
R9248 Transmission_Gate_Layout_8.VIN.n57 Transmission_Gate_Layout_8.VIN.n54 2.6005
R9249 Transmission_Gate_Layout_8.VIN.n58 Transmission_Gate_Layout_8.VIN.n52 2.6005
R9250 Transmission_Gate_Layout_8.VIN.n66 Transmission_Gate_Layout_8.VIN.n65 2.6005
R9251 Transmission_Gate_Layout_8.VIN.n69 Transmission_Gate_Layout_8.VIN.n68 2.6005
R9252 Transmission_Gate_Layout_8.VIN.n14 Transmission_Gate_Layout_8.VIN.n11 2.6005
R9253 Transmission_Gate_Layout_8.VIN.n15 Transmission_Gate_Layout_8.VIN.n9 2.6005
R9254 Transmission_Gate_Layout_8.VIN.n138 Transmission_Gate_Layout_8.VIN.n120 2.6005
R9255 Transmission_Gate_Layout_8.VIN.n139 Transmission_Gate_Layout_8.VIN.n118 2.6005
R9256 Transmission_Gate_Layout_8.VIN.n140 Transmission_Gate_Layout_8.VIN.n116 2.6005
R9257 Transmission_Gate_Layout_8.VIN.n136 Transmission_Gate_Layout_8.VIN.n135 2.6005
R9258 Transmission_Gate_Layout_8.VIN.n133 Transmission_Gate_Layout_8.VIN.n132 2.6005
R9259 Transmission_Gate_Layout_8.VIN.n92 Transmission_Gate_Layout_8.VIN.n83 2.47941
R9260 Transmission_Gate_Layout_8.VIN.n113 Transmission_Gate_Layout_8.VIN.t60 1.3109
R9261 Transmission_Gate_Layout_8.VIN.n113 Transmission_Gate_Layout_8.VIN.n112 1.3109
R9262 Transmission_Gate_Layout_8.VIN.n110 Transmission_Gate_Layout_8.VIN.t61 1.3109
R9263 Transmission_Gate_Layout_8.VIN.n110 Transmission_Gate_Layout_8.VIN.n109 1.3109
R9264 Transmission_Gate_Layout_8.VIN.n107 Transmission_Gate_Layout_8.VIN.t53 1.3109
R9265 Transmission_Gate_Layout_8.VIN.n107 Transmission_Gate_Layout_8.VIN.n106 1.3109
R9266 Transmission_Gate_Layout_8.VIN.n85 Transmission_Gate_Layout_8.VIN.t94 1.3109
R9267 Transmission_Gate_Layout_8.VIN.n85 Transmission_Gate_Layout_8.VIN.n84 1.3109
R9268 Transmission_Gate_Layout_8.VIN.n87 Transmission_Gate_Layout_8.VIN.t85 1.3109
R9269 Transmission_Gate_Layout_8.VIN.n87 Transmission_Gate_Layout_8.VIN.n86 1.3109
R9270 Transmission_Gate_Layout_8.VIN.n89 Transmission_Gate_Layout_8.VIN.t95 1.3109
R9271 Transmission_Gate_Layout_8.VIN.n89 Transmission_Gate_Layout_8.VIN.n88 1.3109
R9272 Transmission_Gate_Layout_8.VIN.n33 Transmission_Gate_Layout_8.VIN.t87 1.3109
R9273 Transmission_Gate_Layout_8.VIN.n33 Transmission_Gate_Layout_8.VIN.n32 1.3109
R9274 Transmission_Gate_Layout_8.VIN.n30 Transmission_Gate_Layout_8.VIN.t90 1.3109
R9275 Transmission_Gate_Layout_8.VIN.n30 Transmission_Gate_Layout_8.VIN.n29 1.3109
R9276 Transmission_Gate_Layout_8.VIN.n28 Transmission_Gate_Layout_8.VIN.t88 1.3109
R9277 Transmission_Gate_Layout_8.VIN.n28 Transmission_Gate_Layout_8.VIN.n27 1.3109
R9278 Transmission_Gate_Layout_8.VIN.n41 Transmission_Gate_Layout_8.VIN.t92 1.3109
R9279 Transmission_Gate_Layout_8.VIN.n41 Transmission_Gate_Layout_8.VIN.n40 1.3109
R9280 Transmission_Gate_Layout_8.VIN.n38 Transmission_Gate_Layout_8.VIN.t84 1.3109
R9281 Transmission_Gate_Layout_8.VIN.n38 Transmission_Gate_Layout_8.VIN.n37 1.3109
R9282 Transmission_Gate_Layout_8.VIN.n36 Transmission_Gate_Layout_8.VIN.t93 1.3109
R9283 Transmission_Gate_Layout_8.VIN.n36 Transmission_Gate_Layout_8.VIN.n35 1.3109
R9284 Transmission_Gate_Layout_8.VIN.n97 Transmission_Gate_Layout_8.VIN.t69 1.3109
R9285 Transmission_Gate_Layout_8.VIN.n97 Transmission_Gate_Layout_8.VIN.n96 1.3109
R9286 Transmission_Gate_Layout_8.VIN.n99 Transmission_Gate_Layout_8.VIN.t51 1.3109
R9287 Transmission_Gate_Layout_8.VIN.n99 Transmission_Gate_Layout_8.VIN.n98 1.3109
R9288 Transmission_Gate_Layout_8.VIN.n101 Transmission_Gate_Layout_8.VIN.t49 1.3109
R9289 Transmission_Gate_Layout_8.VIN.n101 Transmission_Gate_Layout_8.VIN.n100 1.3109
R9290 Transmission_Gate_Layout_8.VIN.n17 Transmission_Gate_Layout_8.VIN.t63 1.3109
R9291 Transmission_Gate_Layout_8.VIN.n17 Transmission_Gate_Layout_8.VIN.n16 1.3109
R9292 Transmission_Gate_Layout_8.VIN.n19 Transmission_Gate_Layout_8.VIN.t67 1.3109
R9293 Transmission_Gate_Layout_8.VIN.n19 Transmission_Gate_Layout_8.VIN.n18 1.3109
R9294 Transmission_Gate_Layout_8.VIN.n21 Transmission_Gate_Layout_8.VIN.t55 1.3109
R9295 Transmission_Gate_Layout_8.VIN.n21 Transmission_Gate_Layout_8.VIN.n20 1.3109
R9296 Transmission_Gate_Layout_8.VIN.n1 Transmission_Gate_Layout_8.VIN.t48 1.3109
R9297 Transmission_Gate_Layout_8.VIN.n1 Transmission_Gate_Layout_8.VIN.n0 1.3109
R9298 Transmission_Gate_Layout_8.VIN.n3 Transmission_Gate_Layout_8.VIN.t57 1.3109
R9299 Transmission_Gate_Layout_8.VIN.n3 Transmission_Gate_Layout_8.VIN.n2 1.3109
R9300 Transmission_Gate_Layout_8.VIN.n6 Transmission_Gate_Layout_8.VIN.t71 1.3109
R9301 Transmission_Gate_Layout_8.VIN.n6 Transmission_Gate_Layout_8.VIN.n5 1.3109
R9302 Transmission_Gate_Layout_8.VIN.n128 Transmission_Gate_Layout_8.VIN.n125 1.24485
R9303 Transmission_Gate_Layout_8.VIN.n50 Transmission_Gate_Layout_8.VIN.n49 1.24485
R9304 Transmission_Gate_Layout_8.VIN.n58 Transmission_Gate_Layout_8.VIN.n57 1.24485
R9305 Transmission_Gate_Layout_8.VIN.n69 Transmission_Gate_Layout_8.VIN.n66 1.24485
R9306 Transmission_Gate_Layout_8.VIN.n71 Transmission_Gate_Layout_8.VIN.n70 1.24485
R9307 Transmission_Gate_Layout_8.VIN.n72 Transmission_Gate_Layout_8.VIN.n71 1.24485
R9308 Transmission_Gate_Layout_8.VIN.n76 Transmission_Gate_Layout_8.VIN.n75 1.24485
R9309 Transmission_Gate_Layout_8.VIN.n75 Transmission_Gate_Layout_8.VIN.n74 1.24485
R9310 Transmission_Gate_Layout_8.VIN.n15 Transmission_Gate_Layout_8.VIN.n14 1.24485
R9311 Transmission_Gate_Layout_8.VIN.n140 Transmission_Gate_Layout_8.VIN.n139 1.24485
R9312 Transmission_Gate_Layout_8.VIN.n139 Transmission_Gate_Layout_8.VIN.n138 1.24485
R9313 Transmission_Gate_Layout_8.VIN.n136 Transmission_Gate_Layout_8.VIN.n133 1.24485
R9314 Transmission_Gate_Layout_8.VIN.n73 Transmission_Gate_Layout_8.VIN.n72 1.2018
R9315 Transmission_Gate_Layout_8.VIN.n77 Transmission_Gate_Layout_8.VIN.n76 1.2018
R9316 Transmission_Gate_Layout_8.VIN.n138 Transmission_Gate_Layout_8.VIN.n137 1.2018
R9317 Transmission_Gate_Layout_8.VIN.n137 Transmission_Gate_Layout_8.VIN.n136 1.2018
R9318 Transmission_Gate_Layout_8.VIN.n81 Transmission_Gate_Layout_8.VIN.n80 0.957239
R9319 Transmission_Gate_Layout_8.VIN.n108 Transmission_Gate_Layout_8.VIN.n105 0.957239
R9320 Transmission_Gate_Layout_8.VIN.n142 Transmission_Gate_Layout_8.VIN.n15 0.806587
R9321 Transmission_Gate_Layout_8.VIN.n141 Transmission_Gate_Layout_8.VIN.n140 0.806587
R9322 Transmission_Gate_Layout_8.VIN.n34 Transmission_Gate_Layout_8.VIN.n31 0.755717
R9323 Transmission_Gate_Layout_8.VIN.n42 Transmission_Gate_Layout_8.VIN.n39 0.755717
R9324 Transmission_Gate_Layout_8.VIN.n83 Transmission_Gate_Layout_8.VIN.n82 0.755717
R9325 Transmission_Gate_Layout_8.VIN.n82 Transmission_Gate_Layout_8.VIN.n81 0.755717
R9326 Transmission_Gate_Layout_8.VIN.n91 Transmission_Gate_Layout_8.VIN.n90 0.755717
R9327 Transmission_Gate_Layout_8.VIN.n94 Transmission_Gate_Layout_8.VIN.n93 0.755717
R9328 Transmission_Gate_Layout_8.VIN.n103 Transmission_Gate_Layout_8.VIN.n102 0.755717
R9329 Transmission_Gate_Layout_8.VIN.n23 Transmission_Gate_Layout_8.VIN.n22 0.755717
R9330 Transmission_Gate_Layout_8.VIN.n111 Transmission_Gate_Layout_8.VIN.n108 0.755717
R9331 Transmission_Gate_Layout_8.VIN.n114 Transmission_Gate_Layout_8.VIN.n111 0.755717
R9332 Transmission_Gate_Layout_8.VIN.n7 Transmission_Gate_Layout_8.VIN.n4 0.755717
R9333 Transmission_Gate_Layout_8.VIN.n135 Transmission_Gate_Layout_8.VIN.t42 0.7285
R9334 Transmission_Gate_Layout_8.VIN.n135 Transmission_Gate_Layout_8.VIN.n134 0.7285
R9335 Transmission_Gate_Layout_8.VIN.n130 Transmission_Gate_Layout_8.VIN.t34 0.7285
R9336 Transmission_Gate_Layout_8.VIN.n130 Transmission_Gate_Layout_8.VIN.n129 0.7285
R9337 Transmission_Gate_Layout_8.VIN.n127 Transmission_Gate_Layout_8.VIN.t24 0.7285
R9338 Transmission_Gate_Layout_8.VIN.n127 Transmission_Gate_Layout_8.VIN.n126 0.7285
R9339 Transmission_Gate_Layout_8.VIN.n124 Transmission_Gate_Layout_8.VIN.t33 0.7285
R9340 Transmission_Gate_Layout_8.VIN.n124 Transmission_Gate_Layout_8.VIN.n123 0.7285
R9341 Transmission_Gate_Layout_8.VIN.n122 Transmission_Gate_Layout_8.VIN.t40 0.7285
R9342 Transmission_Gate_Layout_8.VIN.n122 Transmission_Gate_Layout_8.VIN.n121 0.7285
R9343 Transmission_Gate_Layout_8.VIN.n116 Transmission_Gate_Layout_8.VIN.t45 0.7285
R9344 Transmission_Gate_Layout_8.VIN.n116 Transmission_Gate_Layout_8.VIN.n115 0.7285
R9345 Transmission_Gate_Layout_8.VIN.n118 Transmission_Gate_Layout_8.VIN.t39 0.7285
R9346 Transmission_Gate_Layout_8.VIN.n118 Transmission_Gate_Layout_8.VIN.n117 0.7285
R9347 Transmission_Gate_Layout_8.VIN.n120 Transmission_Gate_Layout_8.VIN.t30 0.7285
R9348 Transmission_Gate_Layout_8.VIN.n120 Transmission_Gate_Layout_8.VIN.n119 0.7285
R9349 Transmission_Gate_Layout_8.VIN.n44 Transmission_Gate_Layout_8.VIN.t3 0.7285
R9350 Transmission_Gate_Layout_8.VIN.n44 Transmission_Gate_Layout_8.VIN.n43 0.7285
R9351 Transmission_Gate_Layout_8.VIN.n46 Transmission_Gate_Layout_8.VIN.t9 0.7285
R9352 Transmission_Gate_Layout_8.VIN.n46 Transmission_Gate_Layout_8.VIN.n45 0.7285
R9353 Transmission_Gate_Layout_8.VIN.n48 Transmission_Gate_Layout_8.VIN.t18 0.7285
R9354 Transmission_Gate_Layout_8.VIN.n48 Transmission_Gate_Layout_8.VIN.n47 0.7285
R9355 Transmission_Gate_Layout_8.VIN.n52 Transmission_Gate_Layout_8.VIN.t16 0.7285
R9356 Transmission_Gate_Layout_8.VIN.n52 Transmission_Gate_Layout_8.VIN.n51 0.7285
R9357 Transmission_Gate_Layout_8.VIN.n54 Transmission_Gate_Layout_8.VIN.t23 0.7285
R9358 Transmission_Gate_Layout_8.VIN.n54 Transmission_Gate_Layout_8.VIN.n53 0.7285
R9359 Transmission_Gate_Layout_8.VIN.n56 Transmission_Gate_Layout_8.VIN.t8 0.7285
R9360 Transmission_Gate_Layout_8.VIN.n56 Transmission_Gate_Layout_8.VIN.n55 0.7285
R9361 Transmission_Gate_Layout_8.VIN.n68 Transmission_Gate_Layout_8.VIN.t15 0.7285
R9362 Transmission_Gate_Layout_8.VIN.n68 Transmission_Gate_Layout_8.VIN.n67 0.7285
R9363 Transmission_Gate_Layout_8.VIN.n65 Transmission_Gate_Layout_8.VIN.t7 0.7285
R9364 Transmission_Gate_Layout_8.VIN.n65 Transmission_Gate_Layout_8.VIN.n64 0.7285
R9365 Transmission_Gate_Layout_8.VIN.n63 Transmission_Gate_Layout_8.VIN.t0 0.7285
R9366 Transmission_Gate_Layout_8.VIN.n63 Transmission_Gate_Layout_8.VIN.n62 0.7285
R9367 Transmission_Gate_Layout_8.VIN.n9 Transmission_Gate_Layout_8.VIN.t32 0.7285
R9368 Transmission_Gate_Layout_8.VIN.n9 Transmission_Gate_Layout_8.VIN.n8 0.7285
R9369 Transmission_Gate_Layout_8.VIN.n11 Transmission_Gate_Layout_8.VIN.t25 0.7285
R9370 Transmission_Gate_Layout_8.VIN.n11 Transmission_Gate_Layout_8.VIN.n10 0.7285
R9371 Transmission_Gate_Layout_8.VIN.n13 Transmission_Gate_Layout_8.VIN.t41 0.7285
R9372 Transmission_Gate_Layout_8.VIN.n13 Transmission_Gate_Layout_8.VIN.n12 0.7285
R9373 Transmission_Gate_Layout_8.VIN.n132 Transmission_Gate_Layout_8.VIN.t26 0.7285
R9374 Transmission_Gate_Layout_8.VIN.n132 Transmission_Gate_Layout_8.VIN.n131 0.7285
R9375 Transmission_Gate_Layout_8.VIN.n78 Transmission_Gate_Layout_8.VIN.n77 0.626587
R9376 Transmission_Gate_Layout_8.VIN.n80 Transmission_Gate_Layout_8.VIN.n79 0.626587
R9377 Transmission_Gate_Layout_8.VIN.n142 Transmission_Gate_Layout_8.VIN.n141 0.626587
R9378 Transmission_Gate_Layout_8.VIN.n70 Transmission_Gate_Layout_8.VIN 0.607022
R9379 Transmission_Gate_Layout_8.VIN.n95 Transmission_Gate_Layout_8.VIN.n92 0.579785
R9380 Transmission_Gate_Layout_8.VIN.n137 Transmission_Gate_Layout_8.VIN.n128 0.575717
R9381 Transmission_Gate_Layout_8.VIN.n78 Transmission_Gate_Layout_8.VIN.n50 0.575717
R9382 Transmission_Gate_Layout_8.VIN.n77 Transmission_Gate_Layout_8.VIN.n58 0.575717
R9383 Transmission_Gate_Layout_8.VIN.n73 Transmission_Gate_Layout_8.VIN.n69 0.575717
R9384 Transmission_Gate_Layout_8.VIN.n105 Transmission_Gate_Layout_8.VIN.n104 0.570002
R9385 Transmission_Gate_Layout_8.VIN.n141 Transmission_Gate_Layout_8.VIN.n114 0.428978
R9386 Transmission_Gate_Layout_8.VIN.n142 Transmission_Gate_Layout_8.VIN.n7 0.428978
R9387 Transmission_Gate_Layout_8.VIN.n80 Transmission_Gate_Layout_8.VIN.n34 0.331152
R9388 Transmission_Gate_Layout_8.VIN.n79 Transmission_Gate_Layout_8.VIN.n42 0.331152
R9389 Transmission_Gate_Layout_8.VIN.n92 Transmission_Gate_Layout_8.VIN.n91 0.331152
R9390 Transmission_Gate_Layout_8.VIN.n105 Transmission_Gate_Layout_8.VIN.n23 0.331152
R9391 Transmission_Gate_Layout_8.VIN.n95 Transmission_Gate_Layout_8.VIN.n94 0.317457
R9392 Transmission_Gate_Layout_8.VIN.n104 Transmission_Gate_Layout_8.VIN.n103 0.317457
R9393 Transmission_Gate_Layout_8.VIN.n79 Transmission_Gate_Layout_8.VIN.n78 0.239196
R9394 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.VIN.n142 0.192239
R9395 B1.n2 B1.t0 34.6755
R9396 B1.n1 B1.t3 34.6599
R9397 B1.n0 B1.t4 32.1987
R9398 B1 B1.n2 17.6692
R9399 B1.n1 B1.n0 17.2076
R9400 B1.n2 B1.t1 13.1666
R9401 B1.n0 B1.t2 11.2112
R9402 B1 B1.n1 4.11202
R9403 B1.n3 B1 2.15659
R9404 B1 B1.n3 0.297891
R9405 B1.n3 B1 0.0768043
R9406 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.n1 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.t4 34.6599
R9407 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.t3 32.1987
R9408 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.n1 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.n0 17.2076
R9409 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.t2 11.2112
R9410 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.n2 7.70137
R9411 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.n3 4.70224
R9412 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT.n1 4.11202
R9413 Transmission_Gate_Layout_12.CLKB.n24 Transmission_Gate_Layout_12.CLKB.t26 54.5477
R9414 Transmission_Gate_Layout_12.CLKB.n29 Transmission_Gate_Layout_12.CLKB.t27 38.3255
R9415 Transmission_Gate_Layout_12.CLKB.n28 Transmission_Gate_Layout_12.CLKB.t23 38.3255
R9416 Transmission_Gate_Layout_12.CLKB.n27 Transmission_Gate_Layout_12.CLKB.t8 38.3255
R9417 Transmission_Gate_Layout_12.CLKB.n26 Transmission_Gate_Layout_12.CLKB.t28 38.3255
R9418 Transmission_Gate_Layout_12.CLKB.n25 Transmission_Gate_Layout_12.CLKB.t24 38.3255
R9419 Transmission_Gate_Layout_12.CLKB.n24 Transmission_Gate_Layout_12.CLKB.t10 38.3255
R9420 Transmission_Gate_Layout_12.CLKB.t16 Transmission_Gate_Layout_12.CLKB.n2 37.9344
R9421 Transmission_Gate_Layout_12.CLKB.t7 Transmission_Gate_Layout_12.CLKB.n5 37.9344
R9422 Transmission_Gate_Layout_12.CLKB.t20 Transmission_Gate_Layout_12.CLKB.n8 37.9344
R9423 Transmission_Gate_Layout_12.CLKB.t17 Transmission_Gate_Layout_12.CLKB.n11 37.9344
R9424 Transmission_Gate_Layout_12.CLKB.t9 Transmission_Gate_Layout_12.CLKB.n14 37.9344
R9425 Transmission_Gate_Layout_12.CLKB.t21 Transmission_Gate_Layout_12.CLKB.n17 37.9344
R9426 Transmission_Gate_Layout_12.CLKB.t13 Transmission_Gate_Layout_12.CLKB.n20 37.9344
R9427 Transmission_Gate_Layout_12.CLKB.t25 Transmission_Gate_Layout_12.CLKB.n21 37.9344
R9428 Transmission_Gate_Layout_12.CLKB.n3 Transmission_Gate_Layout_12.CLKB.t16 37.5434
R9429 Transmission_Gate_Layout_12.CLKB.n6 Transmission_Gate_Layout_12.CLKB.t7 37.5434
R9430 Transmission_Gate_Layout_12.CLKB.n9 Transmission_Gate_Layout_12.CLKB.t20 37.5434
R9431 Transmission_Gate_Layout_12.CLKB.n12 Transmission_Gate_Layout_12.CLKB.t17 37.5434
R9432 Transmission_Gate_Layout_12.CLKB.n15 Transmission_Gate_Layout_12.CLKB.t9 37.5434
R9433 Transmission_Gate_Layout_12.CLKB.n18 Transmission_Gate_Layout_12.CLKB.t21 37.5434
R9434 Transmission_Gate_Layout_12.CLKB.n23 Transmission_Gate_Layout_12.CLKB.t13 37.5434
R9435 Transmission_Gate_Layout_12.CLKB.n22 Transmission_Gate_Layout_12.CLKB.t25 37.5434
R9436 Transmission_Gate_Layout_12.CLKB.t27 Transmission_Gate_Layout_12.CLKB.n3 37.413
R9437 Transmission_Gate_Layout_12.CLKB.t23 Transmission_Gate_Layout_12.CLKB.n6 37.413
R9438 Transmission_Gate_Layout_12.CLKB.t8 Transmission_Gate_Layout_12.CLKB.n9 37.413
R9439 Transmission_Gate_Layout_12.CLKB.t28 Transmission_Gate_Layout_12.CLKB.n12 37.413
R9440 Transmission_Gate_Layout_12.CLKB.t24 Transmission_Gate_Layout_12.CLKB.n15 37.413
R9441 Transmission_Gate_Layout_12.CLKB.t10 Transmission_Gate_Layout_12.CLKB.n18 37.413
R9442 Transmission_Gate_Layout_12.CLKB.n22 Transmission_Gate_Layout_12.CLKB.t15 37.413
R9443 Transmission_Gate_Layout_12.CLKB.t26 Transmission_Gate_Layout_12.CLKB.n23 37.413
R9444 Transmission_Gate_Layout_12.CLKB.n21 Transmission_Gate_Layout_12.CLKB.t22 37.0219
R9445 Transmission_Gate_Layout_12.CLKB.n17 Transmission_Gate_Layout_12.CLKB.t19 37.0219
R9446 Transmission_Gate_Layout_12.CLKB.n14 Transmission_Gate_Layout_12.CLKB.t6 37.0219
R9447 Transmission_Gate_Layout_12.CLKB.n11 Transmission_Gate_Layout_12.CLKB.t14 37.0219
R9448 Transmission_Gate_Layout_12.CLKB.n8 Transmission_Gate_Layout_12.CLKB.t18 37.0219
R9449 Transmission_Gate_Layout_12.CLKB.n5 Transmission_Gate_Layout_12.CLKB.t29 37.0219
R9450 Transmission_Gate_Layout_12.CLKB.n2 Transmission_Gate_Layout_12.CLKB.t12 37.0219
R9451 Transmission_Gate_Layout_12.CLKB.n20 Transmission_Gate_Layout_12.CLKB.t11 37.0219
R9452 Transmission_Gate_Layout_12.CLKB.t19 Transmission_Gate_Layout_12.CLKB.n16 35.1969
R9453 Transmission_Gate_Layout_12.CLKB.t6 Transmission_Gate_Layout_12.CLKB.n13 35.1969
R9454 Transmission_Gate_Layout_12.CLKB.t14 Transmission_Gate_Layout_12.CLKB.n10 35.1969
R9455 Transmission_Gate_Layout_12.CLKB.t18 Transmission_Gate_Layout_12.CLKB.n7 35.1969
R9456 Transmission_Gate_Layout_12.CLKB.t29 Transmission_Gate_Layout_12.CLKB.n4 35.1969
R9457 Transmission_Gate_Layout_12.CLKB.t11 Transmission_Gate_Layout_12.CLKB.n19 35.1969
R9458 Transmission_Gate_Layout_12.CLKB Transmission_Gate_Layout_12.CLKB.n29 26.6826
R9459 Transmission_Gate_Layout_12.CLKB.n23 Transmission_Gate_Layout_12.CLKB.n22 19.148
R9460 Transmission_Gate_Layout_12.CLKB.n29 Transmission_Gate_Layout_12.CLKB.n28 16.2227
R9461 Transmission_Gate_Layout_12.CLKB.n28 Transmission_Gate_Layout_12.CLKB.n27 16.2227
R9462 Transmission_Gate_Layout_12.CLKB.n27 Transmission_Gate_Layout_12.CLKB.n26 16.2227
R9463 Transmission_Gate_Layout_12.CLKB.n26 Transmission_Gate_Layout_12.CLKB.n25 16.2227
R9464 Transmission_Gate_Layout_12.CLKB.n25 Transmission_Gate_Layout_12.CLKB.n24 16.2227
R9465 Transmission_Gate_Layout_12.CLKB.n30 Transmission_Gate_Layout_12.CLKB.t3 5.21612
R9466 Transmission_Gate_Layout_12.CLKB.n0 Transmission_Gate_Layout_12.CLKB.t1 4.57285
R9467 Transmission_Gate_Layout_12.CLKB.n31 Transmission_Gate_Layout_12.CLKB.t4 4.4609
R9468 Transmission_Gate_Layout_12.CLKB.n30 Transmission_Gate_Layout_12.CLKB.t5 4.4609
R9469 Transmission_Gate_Layout_12.CLKB.n0 Transmission_Gate_Layout_12.CLKB.t0 3.3285
R9470 Transmission_Gate_Layout_12.CLKB.n1 Transmission_Gate_Layout_12.CLKB.t2 3.3285
R9471 Transmission_Gate_Layout_12.CLKB.n1 Transmission_Gate_Layout_12.CLKB.n0 1.24485
R9472 Transmission_Gate_Layout_12.CLKB.n31 Transmission_Gate_Layout_12.CLKB.n30 0.755717
R9473 Transmission_Gate_Layout_12.CLKB Transmission_Gate_Layout_12.CLKB.n1 0.750969
R9474 Transmission_Gate_Layout_12.CLKB Transmission_Gate_Layout_12.CLKB.n31 0.510317
R9475 Transmission_Gate_Layout_16.CLKB.n27 Transmission_Gate_Layout_16.CLKB.t18 54.5477
R9476 Transmission_Gate_Layout_16.CLKB.n27 Transmission_Gate_Layout_16.CLKB.t24 38.3255
R9477 Transmission_Gate_Layout_16.CLKB.n28 Transmission_Gate_Layout_16.CLKB.t17 38.3255
R9478 Transmission_Gate_Layout_16.CLKB.n29 Transmission_Gate_Layout_16.CLKB.t23 38.3255
R9479 Transmission_Gate_Layout_16.CLKB.n30 Transmission_Gate_Layout_16.CLKB.t26 38.3255
R9480 Transmission_Gate_Layout_16.CLKB.n31 Transmission_Gate_Layout_16.CLKB.t8 38.3255
R9481 Transmission_Gate_Layout_16.CLKB.n32 Transmission_Gate_Layout_16.CLKB.t14 38.3255
R9482 Transmission_Gate_Layout_16.CLKB.t27 Transmission_Gate_Layout_16.CLKB.n24 37.9344
R9483 Transmission_Gate_Layout_16.CLKB.t10 Transmission_Gate_Layout_16.CLKB.n23 37.9344
R9484 Transmission_Gate_Layout_16.CLKB.t16 Transmission_Gate_Layout_16.CLKB.n20 37.9344
R9485 Transmission_Gate_Layout_16.CLKB.t9 Transmission_Gate_Layout_16.CLKB.n17 37.9344
R9486 Transmission_Gate_Layout_16.CLKB.t15 Transmission_Gate_Layout_16.CLKB.n14 37.9344
R9487 Transmission_Gate_Layout_16.CLKB.t19 Transmission_Gate_Layout_16.CLKB.n11 37.9344
R9488 Transmission_Gate_Layout_16.CLKB.t25 Transmission_Gate_Layout_16.CLKB.n8 37.9344
R9489 Transmission_Gate_Layout_16.CLKB.t7 Transmission_Gate_Layout_16.CLKB.n5 37.9344
R9490 Transmission_Gate_Layout_16.CLKB.n25 Transmission_Gate_Layout_16.CLKB.t27 37.5434
R9491 Transmission_Gate_Layout_16.CLKB.n26 Transmission_Gate_Layout_16.CLKB.t10 37.5434
R9492 Transmission_Gate_Layout_16.CLKB.n21 Transmission_Gate_Layout_16.CLKB.t16 37.5434
R9493 Transmission_Gate_Layout_16.CLKB.n18 Transmission_Gate_Layout_16.CLKB.t9 37.5434
R9494 Transmission_Gate_Layout_16.CLKB.n15 Transmission_Gate_Layout_16.CLKB.t15 37.5434
R9495 Transmission_Gate_Layout_16.CLKB.n12 Transmission_Gate_Layout_16.CLKB.t19 37.5434
R9496 Transmission_Gate_Layout_16.CLKB.n9 Transmission_Gate_Layout_16.CLKB.t25 37.5434
R9497 Transmission_Gate_Layout_16.CLKB.n6 Transmission_Gate_Layout_16.CLKB.t7 37.5434
R9498 Transmission_Gate_Layout_16.CLKB.n25 Transmission_Gate_Layout_16.CLKB.t11 37.413
R9499 Transmission_Gate_Layout_16.CLKB.t24 Transmission_Gate_Layout_16.CLKB.n21 37.413
R9500 Transmission_Gate_Layout_16.CLKB.t17 Transmission_Gate_Layout_16.CLKB.n18 37.413
R9501 Transmission_Gate_Layout_16.CLKB.t23 Transmission_Gate_Layout_16.CLKB.n15 37.413
R9502 Transmission_Gate_Layout_16.CLKB.t26 Transmission_Gate_Layout_16.CLKB.n12 37.413
R9503 Transmission_Gate_Layout_16.CLKB.t8 Transmission_Gate_Layout_16.CLKB.n9 37.413
R9504 Transmission_Gate_Layout_16.CLKB.t14 Transmission_Gate_Layout_16.CLKB.n6 37.413
R9505 Transmission_Gate_Layout_16.CLKB.t18 Transmission_Gate_Layout_16.CLKB.n26 37.413
R9506 Transmission_Gate_Layout_16.CLKB.n24 Transmission_Gate_Layout_16.CLKB.t13 37.0219
R9507 Transmission_Gate_Layout_16.CLKB.n23 Transmission_Gate_Layout_16.CLKB.t22 37.0219
R9508 Transmission_Gate_Layout_16.CLKB.n20 Transmission_Gate_Layout_16.CLKB.t29 37.0219
R9509 Transmission_Gate_Layout_16.CLKB.n17 Transmission_Gate_Layout_16.CLKB.t21 37.0219
R9510 Transmission_Gate_Layout_16.CLKB.n14 Transmission_Gate_Layout_16.CLKB.t28 37.0219
R9511 Transmission_Gate_Layout_16.CLKB.n11 Transmission_Gate_Layout_16.CLKB.t6 37.0219
R9512 Transmission_Gate_Layout_16.CLKB.n5 Transmission_Gate_Layout_16.CLKB.t20 37.0219
R9513 Transmission_Gate_Layout_16.CLKB.n8 Transmission_Gate_Layout_16.CLKB.t12 37.0219
R9514 Transmission_Gate_Layout_16.CLKB.t22 Transmission_Gate_Layout_16.CLKB.n22 35.1969
R9515 Transmission_Gate_Layout_16.CLKB.t29 Transmission_Gate_Layout_16.CLKB.n19 35.1969
R9516 Transmission_Gate_Layout_16.CLKB.t21 Transmission_Gate_Layout_16.CLKB.n16 35.1969
R9517 Transmission_Gate_Layout_16.CLKB.t28 Transmission_Gate_Layout_16.CLKB.n13 35.1969
R9518 Transmission_Gate_Layout_16.CLKB.t6 Transmission_Gate_Layout_16.CLKB.n10 35.1969
R9519 Transmission_Gate_Layout_16.CLKB.t12 Transmission_Gate_Layout_16.CLKB.n7 35.1969
R9520 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_16.CLKB.n32 26.6826
R9521 Transmission_Gate_Layout_16.CLKB.n26 Transmission_Gate_Layout_16.CLKB.n25 19.148
R9522 Transmission_Gate_Layout_16.CLKB.n28 Transmission_Gate_Layout_16.CLKB.n27 16.2227
R9523 Transmission_Gate_Layout_16.CLKB.n29 Transmission_Gate_Layout_16.CLKB.n28 16.2227
R9524 Transmission_Gate_Layout_16.CLKB.n30 Transmission_Gate_Layout_16.CLKB.n29 16.2227
R9525 Transmission_Gate_Layout_16.CLKB.n31 Transmission_Gate_Layout_16.CLKB.n30 16.2227
R9526 Transmission_Gate_Layout_16.CLKB.n32 Transmission_Gate_Layout_16.CLKB.n31 16.2227
R9527 Transmission_Gate_Layout_16.CLKB.n2 Transmission_Gate_Layout_16.CLKB.n0 5.21612
R9528 Transmission_Gate_Layout_16.CLKB.n35 Transmission_Gate_Layout_16.CLKB.n34 4.57285
R9529 Transmission_Gate_Layout_16.CLKB.n2 Transmission_Gate_Layout_16.CLKB.n1 4.4609
R9530 Transmission_Gate_Layout_16.CLKB.n4 Transmission_Gate_Layout_16.CLKB.n3 4.4609
R9531 Transmission_Gate_Layout_16.CLKB.n35 Transmission_Gate_Layout_16.CLKB.n33 3.3285
R9532 Transmission_Gate_Layout_16.CLKB.n37 Transmission_Gate_Layout_16.CLKB.n36 3.3285
R9533 Transmission_Gate_Layout_16.CLKB.n37 Transmission_Gate_Layout_16.CLKB.n35 1.24485
R9534 Transmission_Gate_Layout_16.CLKB.n4 Transmission_Gate_Layout_16.CLKB.n2 0.755717
R9535 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_16.CLKB.n37 0.750969
R9536 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_16.CLKB.n4 0.510317
R9537 IN1.n59 IN1 17.6647
R9538 IN1.n56 IN1.n55 3.90572
R9539 IN1.n48 IN1.n47 3.90572
R9540 IN1.n4 IN1.n1 3.90572
R9541 IN1.n26 IN1.n23 3.84485
R9542 IN1.n34 IN1.n31 3.84485
R9543 IN1.n14 IN1.n13 3.84485
R9544 IN1.n56 IN1.n53 3.1505
R9545 IN1.n57 IN1.n51 3.1505
R9546 IN1.n48 IN1.n45 3.1505
R9547 IN1.n49 IN1.n43 3.1505
R9548 IN1.n4 IN1.n3 3.1505
R9549 IN1.n7 IN1.n6 3.1505
R9550 IN1.n68 IN1.n67 3.1505
R9551 IN1.n65 IN1.n64 3.1505
R9552 IN1.n62 IN1.n61 3.1505
R9553 IN1.n26 IN1.n25 2.6005
R9554 IN1.n29 IN1.n28 2.6005
R9555 IN1.n34 IN1.n33 2.6005
R9556 IN1.n37 IN1.n36 2.6005
R9557 IN1.n39 IN1.n21 2.6005
R9558 IN1.n40 IN1.n19 2.6005
R9559 IN1.n41 IN1.n17 2.6005
R9560 IN1.n14 IN1.n11 2.6005
R9561 IN1.n15 IN1.n9 2.6005
R9562 IN1.n51 IN1.t25 1.3109
R9563 IN1.n51 IN1.n50 1.3109
R9564 IN1.n53 IN1.t44 1.3109
R9565 IN1.n53 IN1.n52 1.3109
R9566 IN1.n55 IN1.t39 1.3109
R9567 IN1.n55 IN1.n54 1.3109
R9568 IN1.n43 IN1.t36 1.3109
R9569 IN1.n43 IN1.n42 1.3109
R9570 IN1.n45 IN1.t29 1.3109
R9571 IN1.n45 IN1.n44 1.3109
R9572 IN1.n47 IN1.t47 1.3109
R9573 IN1.n47 IN1.n46 1.3109
R9574 IN1.n61 IN1.t33 1.3109
R9575 IN1.n61 IN1.n60 1.3109
R9576 IN1.n64 IN1.t27 1.3109
R9577 IN1.n64 IN1.n63 1.3109
R9578 IN1.n67 IN1.t46 1.3109
R9579 IN1.n67 IN1.n66 1.3109
R9580 IN1.n6 IN1.t35 1.3109
R9581 IN1.n6 IN1.n5 1.3109
R9582 IN1.n3 IN1.t41 1.3109
R9583 IN1.n3 IN1.n2 1.3109
R9584 IN1.n1 IN1.t24 1.3109
R9585 IN1.n1 IN1.n0 1.3109
R9586 IN1.n29 IN1.n26 1.24485
R9587 IN1.n37 IN1.n34 1.24485
R9588 IN1.n41 IN1.n40 1.24485
R9589 IN1.n40 IN1.n39 1.24485
R9590 IN1.n15 IN1.n14 1.24485
R9591 IN1.n38 IN1.n37 1.2018
R9592 IN1.n39 IN1.n38 1.2018
R9593 IN1.n58 IN1.n57 0.957239
R9594 IN1.n69 IN1.n41 0.806587
R9595 IN1.n70 IN1.n15 0.806587
R9596 IN1.n57 IN1.n56 0.755717
R9597 IN1.n49 IN1.n48 0.755717
R9598 IN1.n7 IN1.n4 0.755717
R9599 IN1.n65 IN1.n62 0.755717
R9600 IN1.n68 IN1.n65 0.755717
R9601 IN1.n17 IN1.t5 0.7285
R9602 IN1.n17 IN1.n16 0.7285
R9603 IN1.n19 IN1.t13 0.7285
R9604 IN1.n19 IN1.n18 0.7285
R9605 IN1.n21 IN1.t0 0.7285
R9606 IN1.n21 IN1.n20 0.7285
R9607 IN1.n28 IN1.t1 0.7285
R9608 IN1.n28 IN1.n27 0.7285
R9609 IN1.n25 IN1.t14 0.7285
R9610 IN1.n25 IN1.n24 0.7285
R9611 IN1.n23 IN1.t6 0.7285
R9612 IN1.n23 IN1.n22 0.7285
R9613 IN1.n36 IN1.t17 0.7285
R9614 IN1.n36 IN1.n35 0.7285
R9615 IN1.n33 IN1.t4 0.7285
R9616 IN1.n33 IN1.n32 0.7285
R9617 IN1.n31 IN1.t21 0.7285
R9618 IN1.n31 IN1.n30 0.7285
R9619 IN1.n9 IN1.t18 0.7285
R9620 IN1.n9 IN1.n8 0.7285
R9621 IN1.n11 IN1.t2 0.7285
R9622 IN1.n11 IN1.n10 0.7285
R9623 IN1.n13 IN1.t16 0.7285
R9624 IN1.n13 IN1.n12 0.7285
R9625 IN1.n70 IN1.n69 0.626587
R9626 IN1.n38 IN1.n29 0.575717
R9627 IN1.n59 IN1.n58 0.570002
R9628 IN1.n70 IN1.n7 0.428978
R9629 IN1.n69 IN1.n68 0.428978
R9630 IN1.n58 IN1.n49 0.331152
R9631 IN1.n62 IN1.n59 0.317457
R9632 IN1 IN1.n70 0.192239
R9633 IN6.n68 IN6 8.15448
R9634 IN6.n4 IN6.n1 3.90572
R9635 IN6.n22 IN6.n21 3.90572
R9636 IN6.n30 IN6.n29 3.90572
R9637 IN6.n14 IN6.n13 3.84485
R9638 IN6.n60 IN6.n57 3.84485
R9639 IN6.n52 IN6.n49 3.84485
R9640 IN6.n7 IN6.n6 3.1505
R9641 IN6.n4 IN6.n3 3.1505
R9642 IN6.n22 IN6.n19 3.1505
R9643 IN6.n23 IN6.n17 3.1505
R9644 IN6.n30 IN6.n27 3.1505
R9645 IN6.n31 IN6.n25 3.1505
R9646 IN6.n35 IN6.n34 3.1505
R9647 IN6.n38 IN6.n37 3.1505
R9648 IN6.n41 IN6.n40 3.1505
R9649 IN6.n14 IN6.n11 2.6005
R9650 IN6.n15 IN6.n9 2.6005
R9651 IN6.n60 IN6.n59 2.6005
R9652 IN6.n63 IN6.n62 2.6005
R9653 IN6.n52 IN6.n51 2.6005
R9654 IN6.n55 IN6.n54 2.6005
R9655 IN6.n65 IN6.n47 2.6005
R9656 IN6.n66 IN6.n45 2.6005
R9657 IN6.n67 IN6.n43 2.6005
R9658 IN6.n1 IN6.t42 1.3109
R9659 IN6.n1 IN6.n0 1.3109
R9660 IN6.n3 IN6.t24 1.3109
R9661 IN6.n3 IN6.n2 1.3109
R9662 IN6.n6 IN6.t32 1.3109
R9663 IN6.n6 IN6.n5 1.3109
R9664 IN6.n40 IN6.t29 1.3109
R9665 IN6.n40 IN6.n39 1.3109
R9666 IN6.n37 IN6.t35 1.3109
R9667 IN6.n37 IN6.n36 1.3109
R9668 IN6.n34 IN6.t28 1.3109
R9669 IN6.n34 IN6.n33 1.3109
R9670 IN6.n17 IN6.t26 1.3109
R9671 IN6.n17 IN6.n16 1.3109
R9672 IN6.n19 IN6.t33 1.3109
R9673 IN6.n19 IN6.n18 1.3109
R9674 IN6.n21 IN6.t47 1.3109
R9675 IN6.n21 IN6.n20 1.3109
R9676 IN6.n25 IN6.t36 1.3109
R9677 IN6.n25 IN6.n24 1.3109
R9678 IN6.n27 IN6.t39 1.3109
R9679 IN6.n27 IN6.n26 1.3109
R9680 IN6.n29 IN6.t40 1.3109
R9681 IN6.n29 IN6.n28 1.3109
R9682 IN6.n15 IN6.n14 1.24485
R9683 IN6.n63 IN6.n60 1.24485
R9684 IN6.n55 IN6.n52 1.24485
R9685 IN6.n67 IN6.n66 1.24485
R9686 IN6.n66 IN6.n65 1.24485
R9687 IN6.n64 IN6.n63 1.2018
R9688 IN6.n65 IN6.n64 1.2018
R9689 IN6.n32 IN6.n31 0.957239
R9690 IN6.n35 IN6.n32 0.957239
R9691 IN6.n68 IN6.n67 0.822239
R9692 IN6.n69 IN6.n15 0.806587
R9693 IN6.n7 IN6.n4 0.755717
R9694 IN6.n23 IN6.n22 0.755717
R9695 IN6.n31 IN6.n30 0.755717
R9696 IN6.n38 IN6.n35 0.755717
R9697 IN6.n41 IN6.n38 0.755717
R9698 IN6.n9 IN6.t13 0.7285
R9699 IN6.n9 IN6.n8 0.7285
R9700 IN6.n11 IN6.t21 0.7285
R9701 IN6.n11 IN6.n10 0.7285
R9702 IN6.n13 IN6.t6 0.7285
R9703 IN6.n13 IN6.n12 0.7285
R9704 IN6.n43 IN6.t19 0.7285
R9705 IN6.n43 IN6.n42 0.7285
R9706 IN6.n45 IN6.t2 0.7285
R9707 IN6.n45 IN6.n44 0.7285
R9708 IN6.n47 IN6.t12 0.7285
R9709 IN6.n47 IN6.n46 0.7285
R9710 IN6.n62 IN6.t20 0.7285
R9711 IN6.n62 IN6.n61 0.7285
R9712 IN6.n59 IN6.t11 0.7285
R9713 IN6.n59 IN6.n58 0.7285
R9714 IN6.n57 IN6.t4 0.7285
R9715 IN6.n57 IN6.n56 0.7285
R9716 IN6.n54 IN6.t14 0.7285
R9717 IN6.n54 IN6.n53 0.7285
R9718 IN6.n51 IN6.t5 0.7285
R9719 IN6.n51 IN6.n50 0.7285
R9720 IN6.n49 IN6.t22 0.7285
R9721 IN6.n49 IN6.n48 0.7285
R9722 IN6.n64 IN6.n55 0.575717
R9723 IN6.n69 IN6.n68 0.552239
R9724 IN6.n68 IN6.n41 0.44463
R9725 IN6.n69 IN6.n7 0.428978
R9726 IN6.n32 IN6.n23 0.331152
R9727 IN6 IN6.n69 0.192239
R9728 Transmission_Gate_Layout_19.CLKB.n27 Transmission_Gate_Layout_19.CLKB.t28 54.5477
R9729 Transmission_Gate_Layout_19.CLKB.n27 Transmission_Gate_Layout_19.CLKB.t6 38.3255
R9730 Transmission_Gate_Layout_19.CLKB.n28 Transmission_Gate_Layout_19.CLKB.t11 38.3255
R9731 Transmission_Gate_Layout_19.CLKB.n29 Transmission_Gate_Layout_19.CLKB.t14 38.3255
R9732 Transmission_Gate_Layout_19.CLKB.n30 Transmission_Gate_Layout_19.CLKB.t20 38.3255
R9733 Transmission_Gate_Layout_19.CLKB.n31 Transmission_Gate_Layout_19.CLKB.t18 38.3255
R9734 Transmission_Gate_Layout_19.CLKB.n32 Transmission_Gate_Layout_19.CLKB.t19 38.3255
R9735 Transmission_Gate_Layout_19.CLKB.t15 Transmission_Gate_Layout_19.CLKB.n24 37.9344
R9736 Transmission_Gate_Layout_19.CLKB.t21 Transmission_Gate_Layout_19.CLKB.n23 37.9344
R9737 Transmission_Gate_Layout_19.CLKB.t23 Transmission_Gate_Layout_19.CLKB.n20 37.9344
R9738 Transmission_Gate_Layout_19.CLKB.t29 Transmission_Gate_Layout_19.CLKB.n17 37.9344
R9739 Transmission_Gate_Layout_19.CLKB.t7 Transmission_Gate_Layout_19.CLKB.n14 37.9344
R9740 Transmission_Gate_Layout_19.CLKB.t13 Transmission_Gate_Layout_19.CLKB.n11 37.9344
R9741 Transmission_Gate_Layout_19.CLKB.t10 Transmission_Gate_Layout_19.CLKB.n8 37.9344
R9742 Transmission_Gate_Layout_19.CLKB.t12 Transmission_Gate_Layout_19.CLKB.n5 37.9344
R9743 Transmission_Gate_Layout_19.CLKB.n25 Transmission_Gate_Layout_19.CLKB.t15 37.5434
R9744 Transmission_Gate_Layout_19.CLKB.n26 Transmission_Gate_Layout_19.CLKB.t21 37.5434
R9745 Transmission_Gate_Layout_19.CLKB.n21 Transmission_Gate_Layout_19.CLKB.t23 37.5434
R9746 Transmission_Gate_Layout_19.CLKB.n18 Transmission_Gate_Layout_19.CLKB.t29 37.5434
R9747 Transmission_Gate_Layout_19.CLKB.n15 Transmission_Gate_Layout_19.CLKB.t7 37.5434
R9748 Transmission_Gate_Layout_19.CLKB.n12 Transmission_Gate_Layout_19.CLKB.t13 37.5434
R9749 Transmission_Gate_Layout_19.CLKB.n9 Transmission_Gate_Layout_19.CLKB.t10 37.5434
R9750 Transmission_Gate_Layout_19.CLKB.n6 Transmission_Gate_Layout_19.CLKB.t12 37.5434
R9751 Transmission_Gate_Layout_19.CLKB.n25 Transmission_Gate_Layout_19.CLKB.t22 37.413
R9752 Transmission_Gate_Layout_19.CLKB.t6 Transmission_Gate_Layout_19.CLKB.n21 37.413
R9753 Transmission_Gate_Layout_19.CLKB.t11 Transmission_Gate_Layout_19.CLKB.n18 37.413
R9754 Transmission_Gate_Layout_19.CLKB.t14 Transmission_Gate_Layout_19.CLKB.n15 37.413
R9755 Transmission_Gate_Layout_19.CLKB.t20 Transmission_Gate_Layout_19.CLKB.n12 37.413
R9756 Transmission_Gate_Layout_19.CLKB.t18 Transmission_Gate_Layout_19.CLKB.n9 37.413
R9757 Transmission_Gate_Layout_19.CLKB.t19 Transmission_Gate_Layout_19.CLKB.n6 37.413
R9758 Transmission_Gate_Layout_19.CLKB.t28 Transmission_Gate_Layout_19.CLKB.n26 37.413
R9759 Transmission_Gate_Layout_19.CLKB.n24 Transmission_Gate_Layout_19.CLKB.t27 37.0219
R9760 Transmission_Gate_Layout_19.CLKB.n23 Transmission_Gate_Layout_19.CLKB.t8 37.0219
R9761 Transmission_Gate_Layout_19.CLKB.n20 Transmission_Gate_Layout_19.CLKB.t9 37.0219
R9762 Transmission_Gate_Layout_19.CLKB.n17 Transmission_Gate_Layout_19.CLKB.t16 37.0219
R9763 Transmission_Gate_Layout_19.CLKB.n14 Transmission_Gate_Layout_19.CLKB.t17 37.0219
R9764 Transmission_Gate_Layout_19.CLKB.n11 Transmission_Gate_Layout_19.CLKB.t26 37.0219
R9765 Transmission_Gate_Layout_19.CLKB.n5 Transmission_Gate_Layout_19.CLKB.t25 37.0219
R9766 Transmission_Gate_Layout_19.CLKB.n8 Transmission_Gate_Layout_19.CLKB.t24 37.0219
R9767 Transmission_Gate_Layout_19.CLKB.t8 Transmission_Gate_Layout_19.CLKB.n22 35.1969
R9768 Transmission_Gate_Layout_19.CLKB.t9 Transmission_Gate_Layout_19.CLKB.n19 35.1969
R9769 Transmission_Gate_Layout_19.CLKB.t16 Transmission_Gate_Layout_19.CLKB.n16 35.1969
R9770 Transmission_Gate_Layout_19.CLKB.t17 Transmission_Gate_Layout_19.CLKB.n13 35.1969
R9771 Transmission_Gate_Layout_19.CLKB.t26 Transmission_Gate_Layout_19.CLKB.n10 35.1969
R9772 Transmission_Gate_Layout_19.CLKB.t24 Transmission_Gate_Layout_19.CLKB.n7 35.1969
R9773 Transmission_Gate_Layout_19.CLKB Transmission_Gate_Layout_19.CLKB.n32 26.6826
R9774 Transmission_Gate_Layout_19.CLKB.n26 Transmission_Gate_Layout_19.CLKB.n25 19.148
R9775 Transmission_Gate_Layout_19.CLKB.n28 Transmission_Gate_Layout_19.CLKB.n27 16.2227
R9776 Transmission_Gate_Layout_19.CLKB.n29 Transmission_Gate_Layout_19.CLKB.n28 16.2227
R9777 Transmission_Gate_Layout_19.CLKB.n30 Transmission_Gate_Layout_19.CLKB.n29 16.2227
R9778 Transmission_Gate_Layout_19.CLKB.n31 Transmission_Gate_Layout_19.CLKB.n30 16.2227
R9779 Transmission_Gate_Layout_19.CLKB.n32 Transmission_Gate_Layout_19.CLKB.n31 16.2227
R9780 Transmission_Gate_Layout_19.CLKB.n2 Transmission_Gate_Layout_19.CLKB.n0 5.21612
R9781 Transmission_Gate_Layout_19.CLKB.n36 Transmission_Gate_Layout_19.CLKB.n34 4.57285
R9782 Transmission_Gate_Layout_19.CLKB.n2 Transmission_Gate_Layout_19.CLKB.n1 4.4609
R9783 Transmission_Gate_Layout_19.CLKB.n4 Transmission_Gate_Layout_19.CLKB.n3 4.4609
R9784 Transmission_Gate_Layout_19.CLKB.n37 Transmission_Gate_Layout_19.CLKB.n33 3.3285
R9785 Transmission_Gate_Layout_19.CLKB.n36 Transmission_Gate_Layout_19.CLKB.n35 3.3285
R9786 Transmission_Gate_Layout_19.CLKB.n37 Transmission_Gate_Layout_19.CLKB.n36 1.24485
R9787 Transmission_Gate_Layout_19.CLKB.n4 Transmission_Gate_Layout_19.CLKB.n2 0.755717
R9788 Transmission_Gate_Layout_19.CLKB Transmission_Gate_Layout_19.CLKB.n37 0.750969
R9789 Transmission_Gate_Layout_19.CLKB Transmission_Gate_Layout_19.CLKB.n4 0.510317
R9790 Transmission_Gate_Layout_1.CLKB.n27 Transmission_Gate_Layout_1.CLKB.t17 54.5477
R9791 Transmission_Gate_Layout_1.CLKB.n27 Transmission_Gate_Layout_1.CLKB.t10 38.3255
R9792 Transmission_Gate_Layout_1.CLKB.n28 Transmission_Gate_Layout_1.CLKB.t15 38.3255
R9793 Transmission_Gate_Layout_1.CLKB.n29 Transmission_Gate_Layout_1.CLKB.t20 38.3255
R9794 Transmission_Gate_Layout_1.CLKB.n30 Transmission_Gate_Layout_1.CLKB.t9 38.3255
R9795 Transmission_Gate_Layout_1.CLKB.n32 Transmission_Gate_Layout_1.CLKB.t29 38.3255
R9796 Transmission_Gate_Layout_1.CLKB.n31 Transmission_Gate_Layout_1.CLKB.t14 38.3255
R9797 Transmission_Gate_Layout_1.CLKB.t24 Transmission_Gate_Layout_1.CLKB.n24 37.9344
R9798 Transmission_Gate_Layout_1.CLKB.t6 Transmission_Gate_Layout_1.CLKB.n23 37.9344
R9799 Transmission_Gate_Layout_1.CLKB.t21 Transmission_Gate_Layout_1.CLKB.n20 37.9344
R9800 Transmission_Gate_Layout_1.CLKB.t27 Transmission_Gate_Layout_1.CLKB.n17 37.9344
R9801 Transmission_Gate_Layout_1.CLKB.t8 Transmission_Gate_Layout_1.CLKB.n14 37.9344
R9802 Transmission_Gate_Layout_1.CLKB.t19 Transmission_Gate_Layout_1.CLKB.n11 37.9344
R9803 Transmission_Gate_Layout_1.CLKB.t26 Transmission_Gate_Layout_1.CLKB.n8 37.9344
R9804 Transmission_Gate_Layout_1.CLKB.t13 Transmission_Gate_Layout_1.CLKB.n5 37.9344
R9805 Transmission_Gate_Layout_1.CLKB.n25 Transmission_Gate_Layout_1.CLKB.t24 37.5434
R9806 Transmission_Gate_Layout_1.CLKB.n26 Transmission_Gate_Layout_1.CLKB.t6 37.5434
R9807 Transmission_Gate_Layout_1.CLKB.n21 Transmission_Gate_Layout_1.CLKB.t21 37.5434
R9808 Transmission_Gate_Layout_1.CLKB.n18 Transmission_Gate_Layout_1.CLKB.t27 37.5434
R9809 Transmission_Gate_Layout_1.CLKB.n15 Transmission_Gate_Layout_1.CLKB.t8 37.5434
R9810 Transmission_Gate_Layout_1.CLKB.n12 Transmission_Gate_Layout_1.CLKB.t19 37.5434
R9811 Transmission_Gate_Layout_1.CLKB.n9 Transmission_Gate_Layout_1.CLKB.t26 37.5434
R9812 Transmission_Gate_Layout_1.CLKB.n6 Transmission_Gate_Layout_1.CLKB.t13 37.5434
R9813 Transmission_Gate_Layout_1.CLKB.n25 Transmission_Gate_Layout_1.CLKB.t12 37.413
R9814 Transmission_Gate_Layout_1.CLKB.t17 Transmission_Gate_Layout_1.CLKB.n26 37.413
R9815 Transmission_Gate_Layout_1.CLKB.t10 Transmission_Gate_Layout_1.CLKB.n21 37.413
R9816 Transmission_Gate_Layout_1.CLKB.t15 Transmission_Gate_Layout_1.CLKB.n18 37.413
R9817 Transmission_Gate_Layout_1.CLKB.t20 Transmission_Gate_Layout_1.CLKB.n15 37.413
R9818 Transmission_Gate_Layout_1.CLKB.t9 Transmission_Gate_Layout_1.CLKB.n12 37.413
R9819 Transmission_Gate_Layout_1.CLKB.t29 Transmission_Gate_Layout_1.CLKB.n6 37.413
R9820 Transmission_Gate_Layout_1.CLKB.t14 Transmission_Gate_Layout_1.CLKB.n9 37.413
R9821 Transmission_Gate_Layout_1.CLKB.n5 Transmission_Gate_Layout_1.CLKB.t11 37.0219
R9822 Transmission_Gate_Layout_1.CLKB.n11 Transmission_Gate_Layout_1.CLKB.t16 37.0219
R9823 Transmission_Gate_Layout_1.CLKB.n14 Transmission_Gate_Layout_1.CLKB.t7 37.0219
R9824 Transmission_Gate_Layout_1.CLKB.n17 Transmission_Gate_Layout_1.CLKB.t25 37.0219
R9825 Transmission_Gate_Layout_1.CLKB.n20 Transmission_Gate_Layout_1.CLKB.t18 37.0219
R9826 Transmission_Gate_Layout_1.CLKB.n23 Transmission_Gate_Layout_1.CLKB.t28 37.0219
R9827 Transmission_Gate_Layout_1.CLKB.n24 Transmission_Gate_Layout_1.CLKB.t22 37.0219
R9828 Transmission_Gate_Layout_1.CLKB.n8 Transmission_Gate_Layout_1.CLKB.t23 37.0219
R9829 Transmission_Gate_Layout_1.CLKB.t16 Transmission_Gate_Layout_1.CLKB.n10 35.1969
R9830 Transmission_Gate_Layout_1.CLKB.t7 Transmission_Gate_Layout_1.CLKB.n13 35.1969
R9831 Transmission_Gate_Layout_1.CLKB.t25 Transmission_Gate_Layout_1.CLKB.n16 35.1969
R9832 Transmission_Gate_Layout_1.CLKB.t18 Transmission_Gate_Layout_1.CLKB.n19 35.1969
R9833 Transmission_Gate_Layout_1.CLKB.t28 Transmission_Gate_Layout_1.CLKB.n22 35.1969
R9834 Transmission_Gate_Layout_1.CLKB.t23 Transmission_Gate_Layout_1.CLKB.n7 35.1969
R9835 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLKB.n32 26.6826
R9836 Transmission_Gate_Layout_1.CLKB.n26 Transmission_Gate_Layout_1.CLKB.n25 19.148
R9837 Transmission_Gate_Layout_1.CLKB.n28 Transmission_Gate_Layout_1.CLKB.n27 16.2227
R9838 Transmission_Gate_Layout_1.CLKB.n29 Transmission_Gate_Layout_1.CLKB.n28 16.2227
R9839 Transmission_Gate_Layout_1.CLKB.n30 Transmission_Gate_Layout_1.CLKB.n29 16.2227
R9840 Transmission_Gate_Layout_1.CLKB.n31 Transmission_Gate_Layout_1.CLKB.n30 16.2227
R9841 Transmission_Gate_Layout_1.CLKB.n32 Transmission_Gate_Layout_1.CLKB.n31 16.2227
R9842 Transmission_Gate_Layout_1.CLKB.n36 Transmission_Gate_Layout_1.CLKB.n35 5.21612
R9843 Transmission_Gate_Layout_1.CLKB.n2 Transmission_Gate_Layout_1.CLKB.n0 4.57285
R9844 Transmission_Gate_Layout_1.CLKB.n37 Transmission_Gate_Layout_1.CLKB.n33 4.4609
R9845 Transmission_Gate_Layout_1.CLKB.n36 Transmission_Gate_Layout_1.CLKB.n34 4.4609
R9846 Transmission_Gate_Layout_1.CLKB.n2 Transmission_Gate_Layout_1.CLKB.n1 3.3285
R9847 Transmission_Gate_Layout_1.CLKB.n4 Transmission_Gate_Layout_1.CLKB.n3 3.3285
R9848 Transmission_Gate_Layout_1.CLKB.n4 Transmission_Gate_Layout_1.CLKB.n2 1.24485
R9849 Transmission_Gate_Layout_1.CLKB.n37 Transmission_Gate_Layout_1.CLKB.n36 0.755717
R9850 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLKB.n4 0.750969
R9851 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_1.CLKB.n37 0.510317
R9852 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT.t2 17.8546
R9853 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT.n0 14.0337
R9854 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT.t3 13.5862
R9855 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT.n1 9.5898
R9856 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_5.OUT.n2 7.76208
R9857 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT.t3 17.8546
R9858 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT.n0 14.0337
R9859 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT.t2 13.5862
R9860 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT.n1 9.5898
R9861 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_4.OUT.n2 7.76208
R9862 Transmission_Gate_Layout_5.CLKB.n24 Transmission_Gate_Layout_5.CLKB.t15 54.5477
R9863 Transmission_Gate_Layout_5.CLKB.n29 Transmission_Gate_Layout_5.CLKB.t21 38.3255
R9864 Transmission_Gate_Layout_5.CLKB.n28 Transmission_Gate_Layout_5.CLKB.t26 38.3255
R9865 Transmission_Gate_Layout_5.CLKB.n27 Transmission_Gate_Layout_5.CLKB.t29 38.3255
R9866 Transmission_Gate_Layout_5.CLKB.n26 Transmission_Gate_Layout_5.CLKB.t10 38.3255
R9867 Transmission_Gate_Layout_5.CLKB.n25 Transmission_Gate_Layout_5.CLKB.t12 38.3255
R9868 Transmission_Gate_Layout_5.CLKB.n24 Transmission_Gate_Layout_5.CLKB.t9 38.3255
R9869 Transmission_Gate_Layout_5.CLKB.t6 Transmission_Gate_Layout_5.CLKB.n2 37.9344
R9870 Transmission_Gate_Layout_5.CLKB.t13 Transmission_Gate_Layout_5.CLKB.n5 37.9344
R9871 Transmission_Gate_Layout_5.CLKB.t14 Transmission_Gate_Layout_5.CLKB.n8 37.9344
R9872 Transmission_Gate_Layout_5.CLKB.t20 Transmission_Gate_Layout_5.CLKB.n11 37.9344
R9873 Transmission_Gate_Layout_5.CLKB.t22 Transmission_Gate_Layout_5.CLKB.n14 37.9344
R9874 Transmission_Gate_Layout_5.CLKB.t19 Transmission_Gate_Layout_5.CLKB.n17 37.9344
R9875 Transmission_Gate_Layout_5.CLKB.t25 Transmission_Gate_Layout_5.CLKB.n20 37.9344
R9876 Transmission_Gate_Layout_5.CLKB.t28 Transmission_Gate_Layout_5.CLKB.n21 37.9344
R9877 Transmission_Gate_Layout_5.CLKB.n3 Transmission_Gate_Layout_5.CLKB.t6 37.5434
R9878 Transmission_Gate_Layout_5.CLKB.n6 Transmission_Gate_Layout_5.CLKB.t13 37.5434
R9879 Transmission_Gate_Layout_5.CLKB.n9 Transmission_Gate_Layout_5.CLKB.t14 37.5434
R9880 Transmission_Gate_Layout_5.CLKB.n12 Transmission_Gate_Layout_5.CLKB.t20 37.5434
R9881 Transmission_Gate_Layout_5.CLKB.n15 Transmission_Gate_Layout_5.CLKB.t22 37.5434
R9882 Transmission_Gate_Layout_5.CLKB.n18 Transmission_Gate_Layout_5.CLKB.t19 37.5434
R9883 Transmission_Gate_Layout_5.CLKB.n23 Transmission_Gate_Layout_5.CLKB.t25 37.5434
R9884 Transmission_Gate_Layout_5.CLKB.n22 Transmission_Gate_Layout_5.CLKB.t28 37.5434
R9885 Transmission_Gate_Layout_5.CLKB.t21 Transmission_Gate_Layout_5.CLKB.n3 37.413
R9886 Transmission_Gate_Layout_5.CLKB.t26 Transmission_Gate_Layout_5.CLKB.n6 37.413
R9887 Transmission_Gate_Layout_5.CLKB.t29 Transmission_Gate_Layout_5.CLKB.n9 37.413
R9888 Transmission_Gate_Layout_5.CLKB.t10 Transmission_Gate_Layout_5.CLKB.n12 37.413
R9889 Transmission_Gate_Layout_5.CLKB.t12 Transmission_Gate_Layout_5.CLKB.n15 37.413
R9890 Transmission_Gate_Layout_5.CLKB.t9 Transmission_Gate_Layout_5.CLKB.n18 37.413
R9891 Transmission_Gate_Layout_5.CLKB.n22 Transmission_Gate_Layout_5.CLKB.t17 37.413
R9892 Transmission_Gate_Layout_5.CLKB.t15 Transmission_Gate_Layout_5.CLKB.n23 37.413
R9893 Transmission_Gate_Layout_5.CLKB.n21 Transmission_Gate_Layout_5.CLKB.t8 37.0219
R9894 Transmission_Gate_Layout_5.CLKB.n17 Transmission_Gate_Layout_5.CLKB.t23 37.0219
R9895 Transmission_Gate_Layout_5.CLKB.n14 Transmission_Gate_Layout_5.CLKB.t27 37.0219
R9896 Transmission_Gate_Layout_5.CLKB.n11 Transmission_Gate_Layout_5.CLKB.t24 37.0219
R9897 Transmission_Gate_Layout_5.CLKB.n8 Transmission_Gate_Layout_5.CLKB.t18 37.0219
R9898 Transmission_Gate_Layout_5.CLKB.n5 Transmission_Gate_Layout_5.CLKB.t16 37.0219
R9899 Transmission_Gate_Layout_5.CLKB.n2 Transmission_Gate_Layout_5.CLKB.t11 37.0219
R9900 Transmission_Gate_Layout_5.CLKB.n20 Transmission_Gate_Layout_5.CLKB.t7 37.0219
R9901 Transmission_Gate_Layout_5.CLKB.t23 Transmission_Gate_Layout_5.CLKB.n16 35.1969
R9902 Transmission_Gate_Layout_5.CLKB.t27 Transmission_Gate_Layout_5.CLKB.n13 35.1969
R9903 Transmission_Gate_Layout_5.CLKB.t24 Transmission_Gate_Layout_5.CLKB.n10 35.1969
R9904 Transmission_Gate_Layout_5.CLKB.t18 Transmission_Gate_Layout_5.CLKB.n7 35.1969
R9905 Transmission_Gate_Layout_5.CLKB.t16 Transmission_Gate_Layout_5.CLKB.n4 35.1969
R9906 Transmission_Gate_Layout_5.CLKB.t7 Transmission_Gate_Layout_5.CLKB.n19 35.1969
R9907 Transmission_Gate_Layout_5.CLKB Transmission_Gate_Layout_5.CLKB.n29 26.6826
R9908 Transmission_Gate_Layout_5.CLKB.n23 Transmission_Gate_Layout_5.CLKB.n22 19.148
R9909 Transmission_Gate_Layout_5.CLKB.n29 Transmission_Gate_Layout_5.CLKB.n28 16.2227
R9910 Transmission_Gate_Layout_5.CLKB.n28 Transmission_Gate_Layout_5.CLKB.n27 16.2227
R9911 Transmission_Gate_Layout_5.CLKB.n27 Transmission_Gate_Layout_5.CLKB.n26 16.2227
R9912 Transmission_Gate_Layout_5.CLKB.n26 Transmission_Gate_Layout_5.CLKB.n25 16.2227
R9913 Transmission_Gate_Layout_5.CLKB.n25 Transmission_Gate_Layout_5.CLKB.n24 16.2227
R9914 Transmission_Gate_Layout_5.CLKB.n30 Transmission_Gate_Layout_5.CLKB.t5 5.21612
R9915 Transmission_Gate_Layout_5.CLKB.n0 Transmission_Gate_Layout_5.CLKB.t0 4.57285
R9916 Transmission_Gate_Layout_5.CLKB.n31 Transmission_Gate_Layout_5.CLKB.t4 4.4609
R9917 Transmission_Gate_Layout_5.CLKB.n30 Transmission_Gate_Layout_5.CLKB.t3 4.4609
R9918 Transmission_Gate_Layout_5.CLKB.n0 Transmission_Gate_Layout_5.CLKB.t1 3.3285
R9919 Transmission_Gate_Layout_5.CLKB.n1 Transmission_Gate_Layout_5.CLKB.t2 3.3285
R9920 Transmission_Gate_Layout_5.CLKB.n1 Transmission_Gate_Layout_5.CLKB.n0 1.24485
R9921 Transmission_Gate_Layout_5.CLKB.n31 Transmission_Gate_Layout_5.CLKB.n30 0.755717
R9922 Transmission_Gate_Layout_5.CLKB Transmission_Gate_Layout_5.CLKB.n1 0.750969
R9923 Transmission_Gate_Layout_5.CLKB Transmission_Gate_Layout_5.CLKB.n31 0.510317
R9924 Transmission_Gate_Layout_10.CLKB.n24 Transmission_Gate_Layout_10.CLKB.t9 54.5477
R9925 Transmission_Gate_Layout_10.CLKB.n29 Transmission_Gate_Layout_10.CLKB.t8 38.3255
R9926 Transmission_Gate_Layout_10.CLKB.n27 Transmission_Gate_Layout_10.CLKB.t29 38.3255
R9927 Transmission_Gate_Layout_10.CLKB.n26 Transmission_Gate_Layout_10.CLKB.t10 38.3255
R9928 Transmission_Gate_Layout_10.CLKB.n25 Transmission_Gate_Layout_10.CLKB.t15 38.3255
R9929 Transmission_Gate_Layout_10.CLKB.n24 Transmission_Gate_Layout_10.CLKB.t27 38.3255
R9930 Transmission_Gate_Layout_10.CLKB.n28 Transmission_Gate_Layout_10.CLKB.t17 38.3255
R9931 Transmission_Gate_Layout_10.CLKB.t14 Transmission_Gate_Layout_10.CLKB.n2 37.9344
R9932 Transmission_Gate_Layout_10.CLKB.t22 Transmission_Gate_Layout_10.CLKB.n5 37.9344
R9933 Transmission_Gate_Layout_10.CLKB.t12 Transmission_Gate_Layout_10.CLKB.n8 37.9344
R9934 Transmission_Gate_Layout_10.CLKB.t18 Transmission_Gate_Layout_10.CLKB.n11 37.9344
R9935 Transmission_Gate_Layout_10.CLKB.t21 Transmission_Gate_Layout_10.CLKB.n14 37.9344
R9936 Transmission_Gate_Layout_10.CLKB.t11 Transmission_Gate_Layout_10.CLKB.n17 37.9344
R9937 Transmission_Gate_Layout_10.CLKB.t16 Transmission_Gate_Layout_10.CLKB.n20 37.9344
R9938 Transmission_Gate_Layout_10.CLKB.t28 Transmission_Gate_Layout_10.CLKB.n21 37.9344
R9939 Transmission_Gate_Layout_10.CLKB.n3 Transmission_Gate_Layout_10.CLKB.t14 37.5434
R9940 Transmission_Gate_Layout_10.CLKB.n6 Transmission_Gate_Layout_10.CLKB.t22 37.5434
R9941 Transmission_Gate_Layout_10.CLKB.n9 Transmission_Gate_Layout_10.CLKB.t12 37.5434
R9942 Transmission_Gate_Layout_10.CLKB.n12 Transmission_Gate_Layout_10.CLKB.t18 37.5434
R9943 Transmission_Gate_Layout_10.CLKB.n15 Transmission_Gate_Layout_10.CLKB.t21 37.5434
R9944 Transmission_Gate_Layout_10.CLKB.n18 Transmission_Gate_Layout_10.CLKB.t11 37.5434
R9945 Transmission_Gate_Layout_10.CLKB.n23 Transmission_Gate_Layout_10.CLKB.t16 37.5434
R9946 Transmission_Gate_Layout_10.CLKB.n22 Transmission_Gate_Layout_10.CLKB.t28 37.5434
R9947 Transmission_Gate_Layout_10.CLKB.t8 Transmission_Gate_Layout_10.CLKB.n3 37.413
R9948 Transmission_Gate_Layout_10.CLKB.t29 Transmission_Gate_Layout_10.CLKB.n9 37.413
R9949 Transmission_Gate_Layout_10.CLKB.t10 Transmission_Gate_Layout_10.CLKB.n12 37.413
R9950 Transmission_Gate_Layout_10.CLKB.t15 Transmission_Gate_Layout_10.CLKB.n15 37.413
R9951 Transmission_Gate_Layout_10.CLKB.t27 Transmission_Gate_Layout_10.CLKB.n18 37.413
R9952 Transmission_Gate_Layout_10.CLKB.t9 Transmission_Gate_Layout_10.CLKB.n23 37.413
R9953 Transmission_Gate_Layout_10.CLKB.n22 Transmission_Gate_Layout_10.CLKB.t23 37.413
R9954 Transmission_Gate_Layout_10.CLKB.t17 Transmission_Gate_Layout_10.CLKB.n6 37.413
R9955 Transmission_Gate_Layout_10.CLKB.n2 Transmission_Gate_Layout_10.CLKB.t24 37.0219
R9956 Transmission_Gate_Layout_10.CLKB.n5 Transmission_Gate_Layout_10.CLKB.t7 37.0219
R9957 Transmission_Gate_Layout_10.CLKB.n8 Transmission_Gate_Layout_10.CLKB.t20 37.0219
R9958 Transmission_Gate_Layout_10.CLKB.n11 Transmission_Gate_Layout_10.CLKB.t26 37.0219
R9959 Transmission_Gate_Layout_10.CLKB.n14 Transmission_Gate_Layout_10.CLKB.t6 37.0219
R9960 Transmission_Gate_Layout_10.CLKB.n17 Transmission_Gate_Layout_10.CLKB.t19 37.0219
R9961 Transmission_Gate_Layout_10.CLKB.n21 Transmission_Gate_Layout_10.CLKB.t13 37.0219
R9962 Transmission_Gate_Layout_10.CLKB.n20 Transmission_Gate_Layout_10.CLKB.t25 37.0219
R9963 Transmission_Gate_Layout_10.CLKB.t7 Transmission_Gate_Layout_10.CLKB.n4 35.1969
R9964 Transmission_Gate_Layout_10.CLKB.t20 Transmission_Gate_Layout_10.CLKB.n7 35.1969
R9965 Transmission_Gate_Layout_10.CLKB.t26 Transmission_Gate_Layout_10.CLKB.n10 35.1969
R9966 Transmission_Gate_Layout_10.CLKB.t6 Transmission_Gate_Layout_10.CLKB.n13 35.1969
R9967 Transmission_Gate_Layout_10.CLKB.t19 Transmission_Gate_Layout_10.CLKB.n16 35.1969
R9968 Transmission_Gate_Layout_10.CLKB.t25 Transmission_Gate_Layout_10.CLKB.n19 35.1969
R9969 Transmission_Gate_Layout_10.CLKB Transmission_Gate_Layout_10.CLKB.n29 26.6826
R9970 Transmission_Gate_Layout_10.CLKB.n23 Transmission_Gate_Layout_10.CLKB.n22 19.148
R9971 Transmission_Gate_Layout_10.CLKB.n29 Transmission_Gate_Layout_10.CLKB.n28 16.2227
R9972 Transmission_Gate_Layout_10.CLKB.n28 Transmission_Gate_Layout_10.CLKB.n27 16.2227
R9973 Transmission_Gate_Layout_10.CLKB.n27 Transmission_Gate_Layout_10.CLKB.n26 16.2227
R9974 Transmission_Gate_Layout_10.CLKB.n26 Transmission_Gate_Layout_10.CLKB.n25 16.2227
R9975 Transmission_Gate_Layout_10.CLKB.n25 Transmission_Gate_Layout_10.CLKB.n24 16.2227
R9976 Transmission_Gate_Layout_10.CLKB.n0 Transmission_Gate_Layout_10.CLKB.t4 5.21612
R9977 Transmission_Gate_Layout_10.CLKB.n30 Transmission_Gate_Layout_10.CLKB.t2 4.57285
R9978 Transmission_Gate_Layout_10.CLKB.n0 Transmission_Gate_Layout_10.CLKB.t3 4.4609
R9979 Transmission_Gate_Layout_10.CLKB.n1 Transmission_Gate_Layout_10.CLKB.t5 4.4609
R9980 Transmission_Gate_Layout_10.CLKB.n31 Transmission_Gate_Layout_10.CLKB.t1 3.3285
R9981 Transmission_Gate_Layout_10.CLKB.n30 Transmission_Gate_Layout_10.CLKB.t0 3.3285
R9982 Transmission_Gate_Layout_10.CLKB.n31 Transmission_Gate_Layout_10.CLKB.n30 1.24485
R9983 Transmission_Gate_Layout_10.CLKB.n1 Transmission_Gate_Layout_10.CLKB.n0 0.755717
R9984 Transmission_Gate_Layout_10.CLKB Transmission_Gate_Layout_10.CLKB.n31 0.750969
R9985 Transmission_Gate_Layout_10.CLKB Transmission_Gate_Layout_10.CLKB.n1 0.510317
R9986 Transmission_Gate_Layout_21.CLKB.n24 Transmission_Gate_Layout_21.CLKB.t11 54.5477
R9987 Transmission_Gate_Layout_21.CLKB.n29 Transmission_Gate_Layout_21.CLKB.t26 38.3255
R9988 Transmission_Gate_Layout_21.CLKB.n27 Transmission_Gate_Layout_21.CLKB.t20 38.3255
R9989 Transmission_Gate_Layout_21.CLKB.n26 Transmission_Gate_Layout_21.CLKB.t25 38.3255
R9990 Transmission_Gate_Layout_21.CLKB.n25 Transmission_Gate_Layout_21.CLKB.t17 38.3255
R9991 Transmission_Gate_Layout_21.CLKB.n24 Transmission_Gate_Layout_21.CLKB.t22 38.3255
R9992 Transmission_Gate_Layout_21.CLKB.n28 Transmission_Gate_Layout_21.CLKB.t14 38.3255
R9993 Transmission_Gate_Layout_21.CLKB.t9 Transmission_Gate_Layout_21.CLKB.n2 37.9344
R9994 Transmission_Gate_Layout_21.CLKB.t21 Transmission_Gate_Layout_21.CLKB.n5 37.9344
R9995 Transmission_Gate_Layout_21.CLKB.t27 Transmission_Gate_Layout_21.CLKB.n8 37.9344
R9996 Transmission_Gate_Layout_21.CLKB.t7 Transmission_Gate_Layout_21.CLKB.n11 37.9344
R9997 Transmission_Gate_Layout_21.CLKB.t24 Transmission_Gate_Layout_21.CLKB.n14 37.9344
R9998 Transmission_Gate_Layout_21.CLKB.t29 Transmission_Gate_Layout_21.CLKB.n17 37.9344
R9999 Transmission_Gate_Layout_21.CLKB.t19 Transmission_Gate_Layout_21.CLKB.n20 37.9344
R10000 Transmission_Gate_Layout_21.CLKB.t23 Transmission_Gate_Layout_21.CLKB.n21 37.9344
R10001 Transmission_Gate_Layout_21.CLKB.n3 Transmission_Gate_Layout_21.CLKB.t9 37.5434
R10002 Transmission_Gate_Layout_21.CLKB.n6 Transmission_Gate_Layout_21.CLKB.t21 37.5434
R10003 Transmission_Gate_Layout_21.CLKB.n9 Transmission_Gate_Layout_21.CLKB.t27 37.5434
R10004 Transmission_Gate_Layout_21.CLKB.n12 Transmission_Gate_Layout_21.CLKB.t7 37.5434
R10005 Transmission_Gate_Layout_21.CLKB.n15 Transmission_Gate_Layout_21.CLKB.t24 37.5434
R10006 Transmission_Gate_Layout_21.CLKB.n18 Transmission_Gate_Layout_21.CLKB.t29 37.5434
R10007 Transmission_Gate_Layout_21.CLKB.n23 Transmission_Gate_Layout_21.CLKB.t19 37.5434
R10008 Transmission_Gate_Layout_21.CLKB.n22 Transmission_Gate_Layout_21.CLKB.t23 37.5434
R10009 Transmission_Gate_Layout_21.CLKB.t26 Transmission_Gate_Layout_21.CLKB.n3 37.413
R10010 Transmission_Gate_Layout_21.CLKB.t20 Transmission_Gate_Layout_21.CLKB.n9 37.413
R10011 Transmission_Gate_Layout_21.CLKB.t25 Transmission_Gate_Layout_21.CLKB.n12 37.413
R10012 Transmission_Gate_Layout_21.CLKB.t17 Transmission_Gate_Layout_21.CLKB.n15 37.413
R10013 Transmission_Gate_Layout_21.CLKB.t22 Transmission_Gate_Layout_21.CLKB.n18 37.413
R10014 Transmission_Gate_Layout_21.CLKB.t11 Transmission_Gate_Layout_21.CLKB.n23 37.413
R10015 Transmission_Gate_Layout_21.CLKB.n22 Transmission_Gate_Layout_21.CLKB.t15 37.413
R10016 Transmission_Gate_Layout_21.CLKB.t14 Transmission_Gate_Layout_21.CLKB.n6 37.413
R10017 Transmission_Gate_Layout_21.CLKB.n2 Transmission_Gate_Layout_21.CLKB.t18 37.0219
R10018 Transmission_Gate_Layout_21.CLKB.n5 Transmission_Gate_Layout_21.CLKB.t6 37.0219
R10019 Transmission_Gate_Layout_21.CLKB.n8 Transmission_Gate_Layout_21.CLKB.t12 37.0219
R10020 Transmission_Gate_Layout_21.CLKB.n11 Transmission_Gate_Layout_21.CLKB.t16 37.0219
R10021 Transmission_Gate_Layout_21.CLKB.n14 Transmission_Gate_Layout_21.CLKB.t10 37.0219
R10022 Transmission_Gate_Layout_21.CLKB.n17 Transmission_Gate_Layout_21.CLKB.t13 37.0219
R10023 Transmission_Gate_Layout_21.CLKB.n21 Transmission_Gate_Layout_21.CLKB.t8 37.0219
R10024 Transmission_Gate_Layout_21.CLKB.n20 Transmission_Gate_Layout_21.CLKB.t28 37.0219
R10025 Transmission_Gate_Layout_21.CLKB.t6 Transmission_Gate_Layout_21.CLKB.n4 35.1969
R10026 Transmission_Gate_Layout_21.CLKB.t12 Transmission_Gate_Layout_21.CLKB.n7 35.1969
R10027 Transmission_Gate_Layout_21.CLKB.t16 Transmission_Gate_Layout_21.CLKB.n10 35.1969
R10028 Transmission_Gate_Layout_21.CLKB.t10 Transmission_Gate_Layout_21.CLKB.n13 35.1969
R10029 Transmission_Gate_Layout_21.CLKB.t13 Transmission_Gate_Layout_21.CLKB.n16 35.1969
R10030 Transmission_Gate_Layout_21.CLKB.t28 Transmission_Gate_Layout_21.CLKB.n19 35.1969
R10031 Transmission_Gate_Layout_21.CLKB Transmission_Gate_Layout_21.CLKB.n29 26.6826
R10032 Transmission_Gate_Layout_21.CLKB.n23 Transmission_Gate_Layout_21.CLKB.n22 19.148
R10033 Transmission_Gate_Layout_21.CLKB.n29 Transmission_Gate_Layout_21.CLKB.n28 16.2227
R10034 Transmission_Gate_Layout_21.CLKB.n28 Transmission_Gate_Layout_21.CLKB.n27 16.2227
R10035 Transmission_Gate_Layout_21.CLKB.n27 Transmission_Gate_Layout_21.CLKB.n26 16.2227
R10036 Transmission_Gate_Layout_21.CLKB.n26 Transmission_Gate_Layout_21.CLKB.n25 16.2227
R10037 Transmission_Gate_Layout_21.CLKB.n25 Transmission_Gate_Layout_21.CLKB.n24 16.2227
R10038 Transmission_Gate_Layout_21.CLKB.n0 Transmission_Gate_Layout_21.CLKB.t4 5.21612
R10039 Transmission_Gate_Layout_21.CLKB.n30 Transmission_Gate_Layout_21.CLKB.t2 4.57285
R10040 Transmission_Gate_Layout_21.CLKB.n0 Transmission_Gate_Layout_21.CLKB.t5 4.4609
R10041 Transmission_Gate_Layout_21.CLKB.n1 Transmission_Gate_Layout_21.CLKB.t3 4.4609
R10042 Transmission_Gate_Layout_21.CLKB.n31 Transmission_Gate_Layout_21.CLKB.t1 3.3285
R10043 Transmission_Gate_Layout_21.CLKB.n30 Transmission_Gate_Layout_21.CLKB.t0 3.3285
R10044 Transmission_Gate_Layout_21.CLKB.n31 Transmission_Gate_Layout_21.CLKB.n30 1.24485
R10045 Transmission_Gate_Layout_21.CLKB.n1 Transmission_Gate_Layout_21.CLKB.n0 0.755717
R10046 Transmission_Gate_Layout_21.CLKB Transmission_Gate_Layout_21.CLKB.n31 0.750969
R10047 Transmission_Gate_Layout_21.CLKB Transmission_Gate_Layout_21.CLKB.n1 0.510317
R10048 Transmission_Gate_Layout_17.CLKB.n27 Transmission_Gate_Layout_17.CLKB.t8 54.5477
R10049 Transmission_Gate_Layout_17.CLKB.n27 Transmission_Gate_Layout_17.CLKB.t24 38.3255
R10050 Transmission_Gate_Layout_17.CLKB.n28 Transmission_Gate_Layout_17.CLKB.t7 38.3255
R10051 Transmission_Gate_Layout_17.CLKB.n29 Transmission_Gate_Layout_17.CLKB.t12 38.3255
R10052 Transmission_Gate_Layout_17.CLKB.n30 Transmission_Gate_Layout_17.CLKB.t14 38.3255
R10053 Transmission_Gate_Layout_17.CLKB.n31 Transmission_Gate_Layout_17.CLKB.t20 38.3255
R10054 Transmission_Gate_Layout_17.CLKB.n32 Transmission_Gate_Layout_17.CLKB.t21 38.3255
R10055 Transmission_Gate_Layout_17.CLKB.t17 Transmission_Gate_Layout_17.CLKB.n24 37.9344
R10056 Transmission_Gate_Layout_17.CLKB.t23 Transmission_Gate_Layout_17.CLKB.n23 37.9344
R10057 Transmission_Gate_Layout_17.CLKB.t16 Transmission_Gate_Layout_17.CLKB.n20 37.9344
R10058 Transmission_Gate_Layout_17.CLKB.t22 Transmission_Gate_Layout_17.CLKB.n17 37.9344
R10059 Transmission_Gate_Layout_17.CLKB.t6 Transmission_Gate_Layout_17.CLKB.n14 37.9344
R10060 Transmission_Gate_Layout_17.CLKB.t9 Transmission_Gate_Layout_17.CLKB.n11 37.9344
R10061 Transmission_Gate_Layout_17.CLKB.t13 Transmission_Gate_Layout_17.CLKB.n8 37.9344
R10062 Transmission_Gate_Layout_17.CLKB.t15 Transmission_Gate_Layout_17.CLKB.n5 37.9344
R10063 Transmission_Gate_Layout_17.CLKB.n25 Transmission_Gate_Layout_17.CLKB.t17 37.5434
R10064 Transmission_Gate_Layout_17.CLKB.n26 Transmission_Gate_Layout_17.CLKB.t23 37.5434
R10065 Transmission_Gate_Layout_17.CLKB.n21 Transmission_Gate_Layout_17.CLKB.t16 37.5434
R10066 Transmission_Gate_Layout_17.CLKB.n18 Transmission_Gate_Layout_17.CLKB.t22 37.5434
R10067 Transmission_Gate_Layout_17.CLKB.n15 Transmission_Gate_Layout_17.CLKB.t6 37.5434
R10068 Transmission_Gate_Layout_17.CLKB.n12 Transmission_Gate_Layout_17.CLKB.t9 37.5434
R10069 Transmission_Gate_Layout_17.CLKB.n9 Transmission_Gate_Layout_17.CLKB.t13 37.5434
R10070 Transmission_Gate_Layout_17.CLKB.n6 Transmission_Gate_Layout_17.CLKB.t15 37.5434
R10071 Transmission_Gate_Layout_17.CLKB.n25 Transmission_Gate_Layout_17.CLKB.t25 37.413
R10072 Transmission_Gate_Layout_17.CLKB.t24 Transmission_Gate_Layout_17.CLKB.n21 37.413
R10073 Transmission_Gate_Layout_17.CLKB.t7 Transmission_Gate_Layout_17.CLKB.n18 37.413
R10074 Transmission_Gate_Layout_17.CLKB.t12 Transmission_Gate_Layout_17.CLKB.n15 37.413
R10075 Transmission_Gate_Layout_17.CLKB.t14 Transmission_Gate_Layout_17.CLKB.n12 37.413
R10076 Transmission_Gate_Layout_17.CLKB.t20 Transmission_Gate_Layout_17.CLKB.n9 37.413
R10077 Transmission_Gate_Layout_17.CLKB.t21 Transmission_Gate_Layout_17.CLKB.n6 37.413
R10078 Transmission_Gate_Layout_17.CLKB.t8 Transmission_Gate_Layout_17.CLKB.n26 37.413
R10079 Transmission_Gate_Layout_17.CLKB.n24 Transmission_Gate_Layout_17.CLKB.t29 37.0219
R10080 Transmission_Gate_Layout_17.CLKB.n23 Transmission_Gate_Layout_17.CLKB.t11 37.0219
R10081 Transmission_Gate_Layout_17.CLKB.n20 Transmission_Gate_Layout_17.CLKB.t28 37.0219
R10082 Transmission_Gate_Layout_17.CLKB.n17 Transmission_Gate_Layout_17.CLKB.t10 37.0219
R10083 Transmission_Gate_Layout_17.CLKB.n14 Transmission_Gate_Layout_17.CLKB.t18 37.0219
R10084 Transmission_Gate_Layout_17.CLKB.n11 Transmission_Gate_Layout_17.CLKB.t19 37.0219
R10085 Transmission_Gate_Layout_17.CLKB.n5 Transmission_Gate_Layout_17.CLKB.t27 37.0219
R10086 Transmission_Gate_Layout_17.CLKB.n8 Transmission_Gate_Layout_17.CLKB.t26 37.0219
R10087 Transmission_Gate_Layout_17.CLKB.t11 Transmission_Gate_Layout_17.CLKB.n22 35.1969
R10088 Transmission_Gate_Layout_17.CLKB.t28 Transmission_Gate_Layout_17.CLKB.n19 35.1969
R10089 Transmission_Gate_Layout_17.CLKB.t10 Transmission_Gate_Layout_17.CLKB.n16 35.1969
R10090 Transmission_Gate_Layout_17.CLKB.t18 Transmission_Gate_Layout_17.CLKB.n13 35.1969
R10091 Transmission_Gate_Layout_17.CLKB.t19 Transmission_Gate_Layout_17.CLKB.n10 35.1969
R10092 Transmission_Gate_Layout_17.CLKB.t26 Transmission_Gate_Layout_17.CLKB.n7 35.1969
R10093 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_17.CLKB.n32 26.6826
R10094 Transmission_Gate_Layout_17.CLKB.n26 Transmission_Gate_Layout_17.CLKB.n25 19.148
R10095 Transmission_Gate_Layout_17.CLKB.n28 Transmission_Gate_Layout_17.CLKB.n27 16.2227
R10096 Transmission_Gate_Layout_17.CLKB.n29 Transmission_Gate_Layout_17.CLKB.n28 16.2227
R10097 Transmission_Gate_Layout_17.CLKB.n30 Transmission_Gate_Layout_17.CLKB.n29 16.2227
R10098 Transmission_Gate_Layout_17.CLKB.n31 Transmission_Gate_Layout_17.CLKB.n30 16.2227
R10099 Transmission_Gate_Layout_17.CLKB.n32 Transmission_Gate_Layout_17.CLKB.n31 16.2227
R10100 Transmission_Gate_Layout_17.CLKB.n2 Transmission_Gate_Layout_17.CLKB.n0 5.21612
R10101 Transmission_Gate_Layout_17.CLKB.n36 Transmission_Gate_Layout_17.CLKB.n34 4.57285
R10102 Transmission_Gate_Layout_17.CLKB.n2 Transmission_Gate_Layout_17.CLKB.n1 4.4609
R10103 Transmission_Gate_Layout_17.CLKB.n4 Transmission_Gate_Layout_17.CLKB.n3 4.4609
R10104 Transmission_Gate_Layout_17.CLKB.n37 Transmission_Gate_Layout_17.CLKB.n33 3.3285
R10105 Transmission_Gate_Layout_17.CLKB.n36 Transmission_Gate_Layout_17.CLKB.n35 3.3285
R10106 Transmission_Gate_Layout_17.CLKB.n37 Transmission_Gate_Layout_17.CLKB.n36 1.24485
R10107 Transmission_Gate_Layout_17.CLKB.n4 Transmission_Gate_Layout_17.CLKB.n2 0.755717
R10108 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_17.CLKB.n37 0.750969
R10109 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_17.CLKB.n4 0.510317
R10110 IN8.n68 IN8 8.14861
R10111 IN8.n14 IN8.n13 3.90572
R10112 IN8.n60 IN8.n57 3.90572
R10113 IN8.n52 IN8.n49 3.90572
R10114 IN8.n4 IN8.n1 3.84485
R10115 IN8.n22 IN8.n21 3.84485
R10116 IN8.n30 IN8.n29 3.84485
R10117 IN8.n14 IN8.n11 3.1505
R10118 IN8.n15 IN8.n9 3.1505
R10119 IN8.n60 IN8.n59 3.1505
R10120 IN8.n63 IN8.n62 3.1505
R10121 IN8.n52 IN8.n51 3.1505
R10122 IN8.n55 IN8.n54 3.1505
R10123 IN8.n65 IN8.n47 3.1505
R10124 IN8.n66 IN8.n45 3.1505
R10125 IN8.n67 IN8.n43 3.1505
R10126 IN8.n7 IN8.n6 2.6005
R10127 IN8.n4 IN8.n3 2.6005
R10128 IN8.n22 IN8.n19 2.6005
R10129 IN8.n23 IN8.n17 2.6005
R10130 IN8.n30 IN8.n27 2.6005
R10131 IN8.n31 IN8.n25 2.6005
R10132 IN8.n35 IN8.n34 2.6005
R10133 IN8.n38 IN8.n37 2.6005
R10134 IN8.n41 IN8.n40 2.6005
R10135 IN8.n9 IN8.t44 1.3109
R10136 IN8.n9 IN8.n8 1.3109
R10137 IN8.n11 IN8.t31 1.3109
R10138 IN8.n11 IN8.n10 1.3109
R10139 IN8.n13 IN8.t39 1.3109
R10140 IN8.n13 IN8.n12 1.3109
R10141 IN8.n43 IN8.t28 1.3109
R10142 IN8.n43 IN8.n42 1.3109
R10143 IN8.n45 IN8.t38 1.3109
R10144 IN8.n45 IN8.n44 1.3109
R10145 IN8.n47 IN8.t24 1.3109
R10146 IN8.n47 IN8.n46 1.3109
R10147 IN8.n62 IN8.t29 1.3109
R10148 IN8.n62 IN8.n61 1.3109
R10149 IN8.n59 IN8.t41 1.3109
R10150 IN8.n59 IN8.n58 1.3109
R10151 IN8.n57 IN8.t35 1.3109
R10152 IN8.n57 IN8.n56 1.3109
R10153 IN8.n54 IN8.t42 1.3109
R10154 IN8.n54 IN8.n53 1.3109
R10155 IN8.n51 IN8.t33 1.3109
R10156 IN8.n51 IN8.n50 1.3109
R10157 IN8.n49 IN8.t27 1.3109
R10158 IN8.n49 IN8.n48 1.3109
R10159 IN8.n7 IN8.n4 1.24485
R10160 IN8.n23 IN8.n22 1.24485
R10161 IN8.n31 IN8.n30 1.24485
R10162 IN8.n38 IN8.n35 1.24485
R10163 IN8.n41 IN8.n38 1.24485
R10164 IN8.n32 IN8.n31 1.2018
R10165 IN8.n35 IN8.n32 1.2018
R10166 IN8.n64 IN8.n63 0.957239
R10167 IN8.n65 IN8.n64 0.957239
R10168 IN8.n68 IN8.n41 0.822239
R10169 IN8.n69 IN8.n7 0.806587
R10170 IN8.n15 IN8.n14 0.755717
R10171 IN8.n63 IN8.n60 0.755717
R10172 IN8.n55 IN8.n52 0.755717
R10173 IN8.n67 IN8.n66 0.755717
R10174 IN8.n66 IN8.n65 0.755717
R10175 IN8.n1 IN8.t14 0.7285
R10176 IN8.n1 IN8.n0 0.7285
R10177 IN8.n3 IN8.t6 0.7285
R10178 IN8.n3 IN8.n2 0.7285
R10179 IN8.n6 IN8.t9 0.7285
R10180 IN8.n6 IN8.n5 0.7285
R10181 IN8.n40 IN8.t16 0.7285
R10182 IN8.n40 IN8.n39 0.7285
R10183 IN8.n37 IN8.t11 0.7285
R10184 IN8.n37 IN8.n36 0.7285
R10185 IN8.n34 IN8.t1 0.7285
R10186 IN8.n34 IN8.n33 0.7285
R10187 IN8.n17 IN8.t2 0.7285
R10188 IN8.n17 IN8.n16 0.7285
R10189 IN8.n19 IN8.t12 0.7285
R10190 IN8.n19 IN8.n18 0.7285
R10191 IN8.n21 IN8.t17 0.7285
R10192 IN8.n21 IN8.n20 0.7285
R10193 IN8.n25 IN8.t23 0.7285
R10194 IN8.n25 IN8.n24 0.7285
R10195 IN8.n27 IN8.t18 0.7285
R10196 IN8.n27 IN8.n26 0.7285
R10197 IN8.n29 IN8.t5 0.7285
R10198 IN8.n29 IN8.n28 0.7285
R10199 IN8.n32 IN8.n23 0.575717
R10200 IN8.n69 IN8.n68 0.552239
R10201 IN8.n68 IN8.n67 0.44463
R10202 IN8.n69 IN8.n15 0.428978
R10203 IN8.n64 IN8.n55 0.331152
R10204 IN8 IN8.n69 0.192239
R10205 IN5.n59 IN5 10.19
R10206 IN5.n56 IN5.n55 3.90572
R10207 IN5.n48 IN5.n47 3.90572
R10208 IN5.n4 IN5.n1 3.90572
R10209 IN5.n26 IN5.n23 3.84485
R10210 IN5.n34 IN5.n31 3.84485
R10211 IN5.n14 IN5.n13 3.84485
R10212 IN5.n56 IN5.n53 3.1505
R10213 IN5.n57 IN5.n51 3.1505
R10214 IN5.n48 IN5.n45 3.1505
R10215 IN5.n49 IN5.n43 3.1505
R10216 IN5.n4 IN5.n3 3.1505
R10217 IN5.n7 IN5.n6 3.1505
R10218 IN5.n68 IN5.n67 3.1505
R10219 IN5.n65 IN5.n64 3.1505
R10220 IN5.n62 IN5.n61 3.1505
R10221 IN5.n26 IN5.n25 2.6005
R10222 IN5.n29 IN5.n28 2.6005
R10223 IN5.n34 IN5.n33 2.6005
R10224 IN5.n37 IN5.n36 2.6005
R10225 IN5.n39 IN5.n21 2.6005
R10226 IN5.n40 IN5.n19 2.6005
R10227 IN5.n41 IN5.n17 2.6005
R10228 IN5.n14 IN5.n11 2.6005
R10229 IN5.n15 IN5.n9 2.6005
R10230 IN5.n51 IN5.t19 1.3109
R10231 IN5.n51 IN5.n50 1.3109
R10232 IN5.n53 IN5.t13 1.3109
R10233 IN5.n53 IN5.n52 1.3109
R10234 IN5.n55 IN5.t7 1.3109
R10235 IN5.n55 IN5.n54 1.3109
R10236 IN5.n43 IN5.t8 1.3109
R10237 IN5.n43 IN5.n42 1.3109
R10238 IN5.n45 IN5.t1 1.3109
R10239 IN5.n45 IN5.n44 1.3109
R10240 IN5.n47 IN5.t21 1.3109
R10241 IN5.n47 IN5.n46 1.3109
R10242 IN5.n61 IN5.t17 1.3109
R10243 IN5.n61 IN5.n60 1.3109
R10244 IN5.n64 IN5.t11 1.3109
R10245 IN5.n64 IN5.n63 1.3109
R10246 IN5.n67 IN5.t5 1.3109
R10247 IN5.n67 IN5.n66 1.3109
R10248 IN5.n6 IN5.t3 1.3109
R10249 IN5.n6 IN5.n5 1.3109
R10250 IN5.n3 IN5.t9 1.3109
R10251 IN5.n3 IN5.n2 1.3109
R10252 IN5.n1 IN5.t16 1.3109
R10253 IN5.n1 IN5.n0 1.3109
R10254 IN5.n29 IN5.n26 1.24485
R10255 IN5.n37 IN5.n34 1.24485
R10256 IN5.n41 IN5.n40 1.24485
R10257 IN5.n40 IN5.n39 1.24485
R10258 IN5.n15 IN5.n14 1.24485
R10259 IN5.n38 IN5.n37 1.2018
R10260 IN5.n39 IN5.n38 1.2018
R10261 IN5.n58 IN5.n57 0.957239
R10262 IN5.n69 IN5.n41 0.806587
R10263 IN5.n70 IN5.n15 0.806587
R10264 IN5.n57 IN5.n56 0.755717
R10265 IN5.n49 IN5.n48 0.755717
R10266 IN5.n7 IN5.n4 0.755717
R10267 IN5.n65 IN5.n62 0.755717
R10268 IN5.n68 IN5.n65 0.755717
R10269 IN5.n17 IN5.t36 0.7285
R10270 IN5.n17 IN5.n16 0.7285
R10271 IN5.n19 IN5.t43 0.7285
R10272 IN5.n19 IN5.n18 0.7285
R10273 IN5.n21 IN5.t31 0.7285
R10274 IN5.n21 IN5.n20 0.7285
R10275 IN5.n28 IN5.t24 0.7285
R10276 IN5.n28 IN5.n27 0.7285
R10277 IN5.n25 IN5.t34 0.7285
R10278 IN5.n25 IN5.n24 0.7285
R10279 IN5.n23 IN5.t26 0.7285
R10280 IN5.n23 IN5.n22 0.7285
R10281 IN5.n36 IN5.t33 0.7285
R10282 IN5.n36 IN5.n35 0.7285
R10283 IN5.n33 IN5.t47 0.7285
R10284 IN5.n33 IN5.n32 0.7285
R10285 IN5.n31 IN5.t39 0.7285
R10286 IN5.n31 IN5.n30 0.7285
R10287 IN5.n9 IN5.t35 0.7285
R10288 IN5.n9 IN5.n8 0.7285
R10289 IN5.n11 IN5.t42 0.7285
R10290 IN5.n11 IN5.n10 0.7285
R10291 IN5.n13 IN5.t30 0.7285
R10292 IN5.n13 IN5.n12 0.7285
R10293 IN5.n70 IN5.n69 0.626587
R10294 IN5.n38 IN5.n29 0.575717
R10295 IN5.n59 IN5.n58 0.570002
R10296 IN5.n70 IN5.n7 0.428978
R10297 IN5.n69 IN5.n68 0.428978
R10298 IN5.n58 IN5.n49 0.331152
R10299 IN5.n62 IN5.n59 0.317457
R10300 IN5 IN5.n70 0.192239
R10301 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.t5 17.8546
R10302 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n0 14.0337
R10303 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.t4 13.5862
R10304 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n2 3.76289
R10305 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n2 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.t3 3.2765
R10306 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n2 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n1 3.2765
R10307 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n4 2.88224
R10308 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n4 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.t2 1.8205
R10309 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n4 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT.n3 1.8205
R10310 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.t4 17.8546
R10311 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n0 14.0337
R10312 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.t5 13.5862
R10313 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n2 3.76289
R10314 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n2 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.t2 3.2765
R10315 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n2 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n1 3.2765
R10316 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n4 2.88224
R10317 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n4 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.t0 1.8205
R10318 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n4 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT.n3 1.8205
R10319 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT.t2 17.8546
R10320 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT.n0 14.0337
R10321 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT.t3 13.5862
R10322 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT.n1 9.5898
R10323 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_5.OUT.n2 7.76208
R10324 Transmission_Gate_Layout_3.CLKB.n27 Transmission_Gate_Layout_3.CLKB.t29 54.5477
R10325 Transmission_Gate_Layout_3.CLKB.n27 Transmission_Gate_Layout_3.CLKB.t13 38.3255
R10326 Transmission_Gate_Layout_3.CLKB.n28 Transmission_Gate_Layout_3.CLKB.t26 38.3255
R10327 Transmission_Gate_Layout_3.CLKB.n29 Transmission_Gate_Layout_3.CLKB.t11 38.3255
R10328 Transmission_Gate_Layout_3.CLKB.n30 Transmission_Gate_Layout_3.CLKB.t25 38.3255
R10329 Transmission_Gate_Layout_3.CLKB.n32 Transmission_Gate_Layout_3.CLKB.t8 38.3255
R10330 Transmission_Gate_Layout_3.CLKB.n31 Transmission_Gate_Layout_3.CLKB.t28 38.3255
R10331 Transmission_Gate_Layout_3.CLKB.t14 Transmission_Gate_Layout_3.CLKB.n24 37.9344
R10332 Transmission_Gate_Layout_3.CLKB.t18 Transmission_Gate_Layout_3.CLKB.n23 37.9344
R10333 Transmission_Gate_Layout_3.CLKB.t24 Transmission_Gate_Layout_3.CLKB.n20 37.9344
R10334 Transmission_Gate_Layout_3.CLKB.t12 Transmission_Gate_Layout_3.CLKB.n17 37.9344
R10335 Transmission_Gate_Layout_3.CLKB.t23 Transmission_Gate_Layout_3.CLKB.n14 37.9344
R10336 Transmission_Gate_Layout_3.CLKB.t9 Transmission_Gate_Layout_3.CLKB.n11 37.9344
R10337 Transmission_Gate_Layout_3.CLKB.t16 Transmission_Gate_Layout_3.CLKB.n8 37.9344
R10338 Transmission_Gate_Layout_3.CLKB.t21 Transmission_Gate_Layout_3.CLKB.n5 37.9344
R10339 Transmission_Gate_Layout_3.CLKB.n25 Transmission_Gate_Layout_3.CLKB.t14 37.5434
R10340 Transmission_Gate_Layout_3.CLKB.n26 Transmission_Gate_Layout_3.CLKB.t18 37.5434
R10341 Transmission_Gate_Layout_3.CLKB.n21 Transmission_Gate_Layout_3.CLKB.t24 37.5434
R10342 Transmission_Gate_Layout_3.CLKB.n18 Transmission_Gate_Layout_3.CLKB.t12 37.5434
R10343 Transmission_Gate_Layout_3.CLKB.n15 Transmission_Gate_Layout_3.CLKB.t23 37.5434
R10344 Transmission_Gate_Layout_3.CLKB.n12 Transmission_Gate_Layout_3.CLKB.t9 37.5434
R10345 Transmission_Gate_Layout_3.CLKB.n9 Transmission_Gate_Layout_3.CLKB.t16 37.5434
R10346 Transmission_Gate_Layout_3.CLKB.n6 Transmission_Gate_Layout_3.CLKB.t21 37.5434
R10347 Transmission_Gate_Layout_3.CLKB.n25 Transmission_Gate_Layout_3.CLKB.t27 37.413
R10348 Transmission_Gate_Layout_3.CLKB.t29 Transmission_Gate_Layout_3.CLKB.n26 37.413
R10349 Transmission_Gate_Layout_3.CLKB.t13 Transmission_Gate_Layout_3.CLKB.n21 37.413
R10350 Transmission_Gate_Layout_3.CLKB.t26 Transmission_Gate_Layout_3.CLKB.n18 37.413
R10351 Transmission_Gate_Layout_3.CLKB.t11 Transmission_Gate_Layout_3.CLKB.n15 37.413
R10352 Transmission_Gate_Layout_3.CLKB.t25 Transmission_Gate_Layout_3.CLKB.n12 37.413
R10353 Transmission_Gate_Layout_3.CLKB.t8 Transmission_Gate_Layout_3.CLKB.n6 37.413
R10354 Transmission_Gate_Layout_3.CLKB.t28 Transmission_Gate_Layout_3.CLKB.n9 37.413
R10355 Transmission_Gate_Layout_3.CLKB.n5 Transmission_Gate_Layout_3.CLKB.t19 37.0219
R10356 Transmission_Gate_Layout_3.CLKB.n11 Transmission_Gate_Layout_3.CLKB.t6 37.0219
R10357 Transmission_Gate_Layout_3.CLKB.n14 Transmission_Gate_Layout_3.CLKB.t20 37.0219
R10358 Transmission_Gate_Layout_3.CLKB.n17 Transmission_Gate_Layout_3.CLKB.t7 37.0219
R10359 Transmission_Gate_Layout_3.CLKB.n20 Transmission_Gate_Layout_3.CLKB.t22 37.0219
R10360 Transmission_Gate_Layout_3.CLKB.n23 Transmission_Gate_Layout_3.CLKB.t17 37.0219
R10361 Transmission_Gate_Layout_3.CLKB.n24 Transmission_Gate_Layout_3.CLKB.t10 37.0219
R10362 Transmission_Gate_Layout_3.CLKB.n8 Transmission_Gate_Layout_3.CLKB.t15 37.0219
R10363 Transmission_Gate_Layout_3.CLKB.t6 Transmission_Gate_Layout_3.CLKB.n10 35.1969
R10364 Transmission_Gate_Layout_3.CLKB.t20 Transmission_Gate_Layout_3.CLKB.n13 35.1969
R10365 Transmission_Gate_Layout_3.CLKB.t7 Transmission_Gate_Layout_3.CLKB.n16 35.1969
R10366 Transmission_Gate_Layout_3.CLKB.t22 Transmission_Gate_Layout_3.CLKB.n19 35.1969
R10367 Transmission_Gate_Layout_3.CLKB.t17 Transmission_Gate_Layout_3.CLKB.n22 35.1969
R10368 Transmission_Gate_Layout_3.CLKB.t15 Transmission_Gate_Layout_3.CLKB.n7 35.1969
R10369 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLKB.n32 26.6826
R10370 Transmission_Gate_Layout_3.CLKB.n26 Transmission_Gate_Layout_3.CLKB.n25 19.148
R10371 Transmission_Gate_Layout_3.CLKB.n28 Transmission_Gate_Layout_3.CLKB.n27 16.2227
R10372 Transmission_Gate_Layout_3.CLKB.n29 Transmission_Gate_Layout_3.CLKB.n28 16.2227
R10373 Transmission_Gate_Layout_3.CLKB.n30 Transmission_Gate_Layout_3.CLKB.n29 16.2227
R10374 Transmission_Gate_Layout_3.CLKB.n31 Transmission_Gate_Layout_3.CLKB.n30 16.2227
R10375 Transmission_Gate_Layout_3.CLKB.n32 Transmission_Gate_Layout_3.CLKB.n31 16.2227
R10376 Transmission_Gate_Layout_3.CLKB.n36 Transmission_Gate_Layout_3.CLKB.n35 5.21612
R10377 Transmission_Gate_Layout_3.CLKB.n2 Transmission_Gate_Layout_3.CLKB.n0 4.57285
R10378 Transmission_Gate_Layout_3.CLKB.n37 Transmission_Gate_Layout_3.CLKB.n33 4.4609
R10379 Transmission_Gate_Layout_3.CLKB.n36 Transmission_Gate_Layout_3.CLKB.n34 4.4609
R10380 Transmission_Gate_Layout_3.CLKB.n2 Transmission_Gate_Layout_3.CLKB.n1 3.3285
R10381 Transmission_Gate_Layout_3.CLKB.n4 Transmission_Gate_Layout_3.CLKB.n3 3.3285
R10382 Transmission_Gate_Layout_3.CLKB.n4 Transmission_Gate_Layout_3.CLKB.n2 1.24485
R10383 Transmission_Gate_Layout_3.CLKB.n37 Transmission_Gate_Layout_3.CLKB.n36 0.755717
R10384 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLKB.n4 0.750969
R10385 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_3.CLKB.n37 0.510317
R10386 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.t3 34.6755
R10387 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.n0 17.6692
R10388 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.t2 13.1666
R10389 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.n1 9.5898
R10390 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_0.OUT.n2 7.50578
R10391 A1.n2 A1.t4 34.6755
R10392 A1.n1 A1.t0 34.6599
R10393 A1.n0 A1.t1 32.1987
R10394 A1 A1.n2 17.6692
R10395 A1.n1 A1.n0 17.2076
R10396 A1.n2 A1.t2 13.1666
R10397 A1.n0 A1.t3 11.2112
R10398 A1 A1.n1 4.11202
R10399 A1.n3 A1 2.15659
R10400 A1 A1.n3 0.297891
R10401 A1.n3 A1 0.0768043
R10402 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.n3 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.n0 5.61007
R10403 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.t3 5.01528
R10404 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.n3 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.n2 2.6005
R10405 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.n2 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.t1 1.8205
R10406 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.n2 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.n1 1.8205
R10407 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1.n3 0.595283
R10408 Transmission_Gate_Layout_20.CLKB.n24 Transmission_Gate_Layout_20.CLKB.t26 54.5477
R10409 Transmission_Gate_Layout_20.CLKB.n29 Transmission_Gate_Layout_20.CLKB.t11 38.3255
R10410 Transmission_Gate_Layout_20.CLKB.n28 Transmission_Gate_Layout_20.CLKB.t13 38.3255
R10411 Transmission_Gate_Layout_20.CLKB.n27 Transmission_Gate_Layout_20.CLKB.t19 38.3255
R10412 Transmission_Gate_Layout_20.CLKB.n26 Transmission_Gate_Layout_20.CLKB.t24 38.3255
R10413 Transmission_Gate_Layout_20.CLKB.n25 Transmission_Gate_Layout_20.CLKB.t18 38.3255
R10414 Transmission_Gate_Layout_20.CLKB.n24 Transmission_Gate_Layout_20.CLKB.t23 38.3255
R10415 Transmission_Gate_Layout_20.CLKB.t20 Transmission_Gate_Layout_20.CLKB.n2 37.9344
R10416 Transmission_Gate_Layout_20.CLKB.t21 Transmission_Gate_Layout_20.CLKB.n5 37.9344
R10417 Transmission_Gate_Layout_20.CLKB.t29 Transmission_Gate_Layout_20.CLKB.n8 37.9344
R10418 Transmission_Gate_Layout_20.CLKB.t10 Transmission_Gate_Layout_20.CLKB.n11 37.9344
R10419 Transmission_Gate_Layout_20.CLKB.t28 Transmission_Gate_Layout_20.CLKB.n14 37.9344
R10420 Transmission_Gate_Layout_20.CLKB.t9 Transmission_Gate_Layout_20.CLKB.n17 37.9344
R10421 Transmission_Gate_Layout_20.CLKB.t12 Transmission_Gate_Layout_20.CLKB.n20 37.9344
R10422 Transmission_Gate_Layout_20.CLKB.t17 Transmission_Gate_Layout_20.CLKB.n21 37.9344
R10423 Transmission_Gate_Layout_20.CLKB.n3 Transmission_Gate_Layout_20.CLKB.t20 37.5434
R10424 Transmission_Gate_Layout_20.CLKB.n6 Transmission_Gate_Layout_20.CLKB.t21 37.5434
R10425 Transmission_Gate_Layout_20.CLKB.n9 Transmission_Gate_Layout_20.CLKB.t29 37.5434
R10426 Transmission_Gate_Layout_20.CLKB.n12 Transmission_Gate_Layout_20.CLKB.t10 37.5434
R10427 Transmission_Gate_Layout_20.CLKB.n15 Transmission_Gate_Layout_20.CLKB.t28 37.5434
R10428 Transmission_Gate_Layout_20.CLKB.n18 Transmission_Gate_Layout_20.CLKB.t9 37.5434
R10429 Transmission_Gate_Layout_20.CLKB.n23 Transmission_Gate_Layout_20.CLKB.t12 37.5434
R10430 Transmission_Gate_Layout_20.CLKB.n22 Transmission_Gate_Layout_20.CLKB.t17 37.5434
R10431 Transmission_Gate_Layout_20.CLKB.t11 Transmission_Gate_Layout_20.CLKB.n3 37.413
R10432 Transmission_Gate_Layout_20.CLKB.t13 Transmission_Gate_Layout_20.CLKB.n6 37.413
R10433 Transmission_Gate_Layout_20.CLKB.t19 Transmission_Gate_Layout_20.CLKB.n9 37.413
R10434 Transmission_Gate_Layout_20.CLKB.t24 Transmission_Gate_Layout_20.CLKB.n12 37.413
R10435 Transmission_Gate_Layout_20.CLKB.t18 Transmission_Gate_Layout_20.CLKB.n15 37.413
R10436 Transmission_Gate_Layout_20.CLKB.t23 Transmission_Gate_Layout_20.CLKB.n18 37.413
R10437 Transmission_Gate_Layout_20.CLKB.n22 Transmission_Gate_Layout_20.CLKB.t6 37.413
R10438 Transmission_Gate_Layout_20.CLKB.t26 Transmission_Gate_Layout_20.CLKB.n23 37.413
R10439 Transmission_Gate_Layout_20.CLKB.n21 Transmission_Gate_Layout_20.CLKB.t22 37.0219
R10440 Transmission_Gate_Layout_20.CLKB.n17 Transmission_Gate_Layout_20.CLKB.t14 37.0219
R10441 Transmission_Gate_Layout_20.CLKB.n14 Transmission_Gate_Layout_20.CLKB.t7 37.0219
R10442 Transmission_Gate_Layout_20.CLKB.n11 Transmission_Gate_Layout_20.CLKB.t15 37.0219
R10443 Transmission_Gate_Layout_20.CLKB.n8 Transmission_Gate_Layout_20.CLKB.t8 37.0219
R10444 Transmission_Gate_Layout_20.CLKB.n5 Transmission_Gate_Layout_20.CLKB.t27 37.0219
R10445 Transmission_Gate_Layout_20.CLKB.n2 Transmission_Gate_Layout_20.CLKB.t25 37.0219
R10446 Transmission_Gate_Layout_20.CLKB.n20 Transmission_Gate_Layout_20.CLKB.t16 37.0219
R10447 Transmission_Gate_Layout_20.CLKB.t14 Transmission_Gate_Layout_20.CLKB.n16 35.1969
R10448 Transmission_Gate_Layout_20.CLKB.t7 Transmission_Gate_Layout_20.CLKB.n13 35.1969
R10449 Transmission_Gate_Layout_20.CLKB.t15 Transmission_Gate_Layout_20.CLKB.n10 35.1969
R10450 Transmission_Gate_Layout_20.CLKB.t8 Transmission_Gate_Layout_20.CLKB.n7 35.1969
R10451 Transmission_Gate_Layout_20.CLKB.t27 Transmission_Gate_Layout_20.CLKB.n4 35.1969
R10452 Transmission_Gate_Layout_20.CLKB.t16 Transmission_Gate_Layout_20.CLKB.n19 35.1969
R10453 Transmission_Gate_Layout_20.CLKB Transmission_Gate_Layout_20.CLKB.n29 26.6826
R10454 Transmission_Gate_Layout_20.CLKB.n23 Transmission_Gate_Layout_20.CLKB.n22 19.148
R10455 Transmission_Gate_Layout_20.CLKB.n29 Transmission_Gate_Layout_20.CLKB.n28 16.2227
R10456 Transmission_Gate_Layout_20.CLKB.n28 Transmission_Gate_Layout_20.CLKB.n27 16.2227
R10457 Transmission_Gate_Layout_20.CLKB.n27 Transmission_Gate_Layout_20.CLKB.n26 16.2227
R10458 Transmission_Gate_Layout_20.CLKB.n26 Transmission_Gate_Layout_20.CLKB.n25 16.2227
R10459 Transmission_Gate_Layout_20.CLKB.n25 Transmission_Gate_Layout_20.CLKB.n24 16.2227
R10460 Transmission_Gate_Layout_20.CLKB.n30 Transmission_Gate_Layout_20.CLKB.t3 5.21612
R10461 Transmission_Gate_Layout_20.CLKB.n0 Transmission_Gate_Layout_20.CLKB.t0 4.57285
R10462 Transmission_Gate_Layout_20.CLKB.n31 Transmission_Gate_Layout_20.CLKB.t4 4.4609
R10463 Transmission_Gate_Layout_20.CLKB.n30 Transmission_Gate_Layout_20.CLKB.t5 4.4609
R10464 Transmission_Gate_Layout_20.CLKB.n0 Transmission_Gate_Layout_20.CLKB.t1 3.3285
R10465 Transmission_Gate_Layout_20.CLKB.n1 Transmission_Gate_Layout_20.CLKB.t2 3.3285
R10466 Transmission_Gate_Layout_20.CLKB.n1 Transmission_Gate_Layout_20.CLKB.n0 1.24485
R10467 Transmission_Gate_Layout_20.CLKB.n31 Transmission_Gate_Layout_20.CLKB.n30 0.755717
R10468 Transmission_Gate_Layout_20.CLKB Transmission_Gate_Layout_20.CLKB.n1 0.750969
R10469 Transmission_Gate_Layout_20.CLKB Transmission_Gate_Layout_20.CLKB.n31 0.510317
R10470 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.t3 34.6755
R10471 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.n0 17.6692
R10472 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.t2 13.1666
R10473 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.n1 9.5898
R10474 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_3.OUT.n2 7.50578
R10475 Transmission_Gate_Layout_4.CLKB.n27 Transmission_Gate_Layout_4.CLKB.t18 54.5477
R10476 Transmission_Gate_Layout_4.CLKB.n27 Transmission_Gate_Layout_4.CLKB.t12 38.3255
R10477 Transmission_Gate_Layout_4.CLKB.n28 Transmission_Gate_Layout_4.CLKB.t17 38.3255
R10478 Transmission_Gate_Layout_4.CLKB.n29 Transmission_Gate_Layout_4.CLKB.t23 38.3255
R10479 Transmission_Gate_Layout_4.CLKB.n30 Transmission_Gate_Layout_4.CLKB.t25 38.3255
R10480 Transmission_Gate_Layout_4.CLKB.n32 Transmission_Gate_Layout_4.CLKB.t9 38.3255
R10481 Transmission_Gate_Layout_4.CLKB.n31 Transmission_Gate_Layout_4.CLKB.t6 38.3255
R10482 Transmission_Gate_Layout_4.CLKB.t21 Transmission_Gate_Layout_4.CLKB.n24 37.9344
R10483 Transmission_Gate_Layout_4.CLKB.t29 Transmission_Gate_Layout_4.CLKB.n23 37.9344
R10484 Transmission_Gate_Layout_4.CLKB.t20 Transmission_Gate_Layout_4.CLKB.n20 37.9344
R10485 Transmission_Gate_Layout_4.CLKB.t28 Transmission_Gate_Layout_4.CLKB.n17 37.9344
R10486 Transmission_Gate_Layout_4.CLKB.t10 Transmission_Gate_Layout_4.CLKB.n14 37.9344
R10487 Transmission_Gate_Layout_4.CLKB.t11 Transmission_Gate_Layout_4.CLKB.n11 37.9344
R10488 Transmission_Gate_Layout_4.CLKB.t16 Transmission_Gate_Layout_4.CLKB.n8 37.9344
R10489 Transmission_Gate_Layout_4.CLKB.t19 Transmission_Gate_Layout_4.CLKB.n5 37.9344
R10490 Transmission_Gate_Layout_4.CLKB.n25 Transmission_Gate_Layout_4.CLKB.t21 37.5434
R10491 Transmission_Gate_Layout_4.CLKB.n26 Transmission_Gate_Layout_4.CLKB.t29 37.5434
R10492 Transmission_Gate_Layout_4.CLKB.n21 Transmission_Gate_Layout_4.CLKB.t20 37.5434
R10493 Transmission_Gate_Layout_4.CLKB.n18 Transmission_Gate_Layout_4.CLKB.t28 37.5434
R10494 Transmission_Gate_Layout_4.CLKB.n15 Transmission_Gate_Layout_4.CLKB.t10 37.5434
R10495 Transmission_Gate_Layout_4.CLKB.n12 Transmission_Gate_Layout_4.CLKB.t11 37.5434
R10496 Transmission_Gate_Layout_4.CLKB.n9 Transmission_Gate_Layout_4.CLKB.t16 37.5434
R10497 Transmission_Gate_Layout_4.CLKB.n6 Transmission_Gate_Layout_4.CLKB.t19 37.5434
R10498 Transmission_Gate_Layout_4.CLKB.n25 Transmission_Gate_Layout_4.CLKB.t13 37.413
R10499 Transmission_Gate_Layout_4.CLKB.t18 Transmission_Gate_Layout_4.CLKB.n26 37.413
R10500 Transmission_Gate_Layout_4.CLKB.t12 Transmission_Gate_Layout_4.CLKB.n21 37.413
R10501 Transmission_Gate_Layout_4.CLKB.t17 Transmission_Gate_Layout_4.CLKB.n18 37.413
R10502 Transmission_Gate_Layout_4.CLKB.t23 Transmission_Gate_Layout_4.CLKB.n15 37.413
R10503 Transmission_Gate_Layout_4.CLKB.t25 Transmission_Gate_Layout_4.CLKB.n12 37.413
R10504 Transmission_Gate_Layout_4.CLKB.t9 Transmission_Gate_Layout_4.CLKB.n6 37.413
R10505 Transmission_Gate_Layout_4.CLKB.t6 Transmission_Gate_Layout_4.CLKB.n9 37.413
R10506 Transmission_Gate_Layout_4.CLKB.n5 Transmission_Gate_Layout_4.CLKB.t24 37.0219
R10507 Transmission_Gate_Layout_4.CLKB.n11 Transmission_Gate_Layout_4.CLKB.t15 37.0219
R10508 Transmission_Gate_Layout_4.CLKB.n14 Transmission_Gate_Layout_4.CLKB.t14 37.0219
R10509 Transmission_Gate_Layout_4.CLKB.n17 Transmission_Gate_Layout_4.CLKB.t7 37.0219
R10510 Transmission_Gate_Layout_4.CLKB.n20 Transmission_Gate_Layout_4.CLKB.t26 37.0219
R10511 Transmission_Gate_Layout_4.CLKB.n23 Transmission_Gate_Layout_4.CLKB.t8 37.0219
R10512 Transmission_Gate_Layout_4.CLKB.n24 Transmission_Gate_Layout_4.CLKB.t27 37.0219
R10513 Transmission_Gate_Layout_4.CLKB.n8 Transmission_Gate_Layout_4.CLKB.t22 37.0219
R10514 Transmission_Gate_Layout_4.CLKB.t15 Transmission_Gate_Layout_4.CLKB.n10 35.1969
R10515 Transmission_Gate_Layout_4.CLKB.t14 Transmission_Gate_Layout_4.CLKB.n13 35.1969
R10516 Transmission_Gate_Layout_4.CLKB.t7 Transmission_Gate_Layout_4.CLKB.n16 35.1969
R10517 Transmission_Gate_Layout_4.CLKB.t26 Transmission_Gate_Layout_4.CLKB.n19 35.1969
R10518 Transmission_Gate_Layout_4.CLKB.t8 Transmission_Gate_Layout_4.CLKB.n22 35.1969
R10519 Transmission_Gate_Layout_4.CLKB.t22 Transmission_Gate_Layout_4.CLKB.n7 35.1969
R10520 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_4.CLKB.n32 26.6826
R10521 Transmission_Gate_Layout_4.CLKB.n26 Transmission_Gate_Layout_4.CLKB.n25 19.148
R10522 Transmission_Gate_Layout_4.CLKB.n28 Transmission_Gate_Layout_4.CLKB.n27 16.2227
R10523 Transmission_Gate_Layout_4.CLKB.n29 Transmission_Gate_Layout_4.CLKB.n28 16.2227
R10524 Transmission_Gate_Layout_4.CLKB.n30 Transmission_Gate_Layout_4.CLKB.n29 16.2227
R10525 Transmission_Gate_Layout_4.CLKB.n31 Transmission_Gate_Layout_4.CLKB.n30 16.2227
R10526 Transmission_Gate_Layout_4.CLKB.n32 Transmission_Gate_Layout_4.CLKB.n31 16.2227
R10527 Transmission_Gate_Layout_4.CLKB.n36 Transmission_Gate_Layout_4.CLKB.n35 5.21612
R10528 Transmission_Gate_Layout_4.CLKB.n2 Transmission_Gate_Layout_4.CLKB.n0 4.57285
R10529 Transmission_Gate_Layout_4.CLKB.n37 Transmission_Gate_Layout_4.CLKB.n33 4.4609
R10530 Transmission_Gate_Layout_4.CLKB.n36 Transmission_Gate_Layout_4.CLKB.n34 4.4609
R10531 Transmission_Gate_Layout_4.CLKB.n2 Transmission_Gate_Layout_4.CLKB.n1 3.3285
R10532 Transmission_Gate_Layout_4.CLKB.n4 Transmission_Gate_Layout_4.CLKB.n3 3.3285
R10533 Transmission_Gate_Layout_4.CLKB.n4 Transmission_Gate_Layout_4.CLKB.n2 1.24485
R10534 Transmission_Gate_Layout_4.CLKB.n37 Transmission_Gate_Layout_4.CLKB.n36 0.755717
R10535 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_4.CLKB.n4 0.750969
R10536 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_4.CLKB.n37 0.510317
R10537 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.t3 34.6755
R10538 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.n0 17.6692
R10539 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.t2 13.1666
R10540 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.n1 9.5898
R10541 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_3.OUT.n2 7.50578
R10542 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.n1 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.t3 34.6599
R10543 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.t4 32.1987
R10544 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.n1 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.n0 17.2076
R10545 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.t2 11.2112
R10546 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.n2 7.70137
R10547 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.n3 4.70224
R10548 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT.n1 4.11202
R10549 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT.t2 17.8546
R10550 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT.n0 14.0337
R10551 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT.t3 13.5862
R10552 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT.n1 9.5898
R10553 Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_2.Inv_16x_Layout_4.OUT.n2 7.76208
R10554 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.n3 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.n0 5.61007
R10555 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.t1 5.01528
R10556 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.n3 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.n2 2.6005
R10557 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.n2 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.t3 1.8205
R10558 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.n2 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.n1 1.8205
R10559 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1.n3 0.595283
R10560 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.n3 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.n2 5.61007
R10561 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.t2 5.01528
R10562 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.n3 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.n1 2.6005
R10563 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.n1 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.t0 1.8205
R10564 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.n1 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.n0 1.8205
R10565 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1.n3 0.595283
R10566 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT.t3 17.8546
R10567 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT.n0 14.0337
R10568 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT.t2 13.5862
R10569 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT.n1 9.5898
R10570 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_5.OUT.n2 7.76208
R10571 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT.t2 17.8546
R10572 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT.n0 14.0337
R10573 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT.t3 13.5862
R10574 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT.n1 9.5898
R10575 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_4.OUT.n2 7.76208
R10576 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT.t2 17.8546
R10577 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT.n0 14.0337
R10578 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT.t3 13.5862
R10579 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT.n1 9.5898
R10580 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_2.OUT.n2 7.76208
R10581 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.t2 34.6755
R10582 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.n0 17.6692
R10583 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.t3 13.1666
R10584 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.n1 9.5898
R10585 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_0.OUT.n2 7.50578
R10586 C1.n2 C1.t3 34.6755
R10587 C1.n1 C1.t0 34.6599
R10588 C1.n0 C1.t1 32.1987
R10589 C1 C1.n2 17.6692
R10590 C1.n1 C1.n0 17.2076
R10591 C1.n2 C1.t2 13.1666
R10592 C1.n0 C1.t4 11.2112
R10593 C1 C1.n1 4.11202
R10594 C1.n3 C1 2.15659
R10595 C1 C1.n3 0.297891
R10596 C1.n3 C1 0.0768043
R10597 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.n3 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.n0 5.61007
R10598 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.t3 5.01528
R10599 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.n3 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.n2 2.6005
R10600 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.n2 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.t1 1.8205
R10601 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.n2 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.n1 1.8205
R10602 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1.n3 0.595283
R10603 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT.t2 17.8546
R10604 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT.n0 14.0337
R10605 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT.t3 13.5862
R10606 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT.n1 9.5898
R10607 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_2.OUT.n2 7.76208
R10608 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.n1 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.t4 34.6599
R10609 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.t3 32.1987
R10610 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.n1 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.n0 17.2076
R10611 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.t2 11.2112
R10612 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.n2 7.70137
R10613 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.n3 4.70224
R10614 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT.n1 4.11202
R10615 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.t5 17.8546
R10616 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n0 14.0337
R10617 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.t4 13.5862
R10618 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n5 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n2 3.76289
R10619 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n2 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.t2 3.2765
R10620 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n2 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n1 3.2765
R10621 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n5 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n4 2.88224
R10622 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n4 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.t1 1.8205
R10623 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n4 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n3 1.8205
R10624 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT.n5 0.155065
R10625 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT.t3 17.8546
R10626 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT.n0 14.0337
R10627 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT.t2 13.5862
R10628 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT.n1 9.5898
R10629 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_1.OUT.n2 7.76208
R10630 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.t2 34.6755
R10631 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.n0 17.6692
R10632 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.t3 13.1666
R10633 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.n1 9.5898
R10634 Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_1.Inv_16x_Layout_0.OUT.n2 7.50578
R10635 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.t2 34.6755
R10636 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.n0 17.6692
R10637 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.n0 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.t3 13.1666
R10638 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.n1 9.5898
R10639 Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT Non_Ovl_CLK_Gen_Layout_0.Inv_16x_Layout_3.OUT.n2 7.50578
R10640 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.t5 17.8546
R10641 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n0 14.0337
R10642 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n0 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.t4 13.5862
R10643 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n2 3.76289
R10644 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n2 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.t3 3.2765
R10645 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n2 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n1 3.2765
R10646 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n4 2.88224
R10647 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n4 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.t2 1.8205
R10648 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n4 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT.n3 1.8205
R10649 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.n3 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.n0 5.61007
R10650 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.t1 5.01528
R10651 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.n3 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.n2 2.6005
R10652 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.n2 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.t3 1.8205
R10653 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.n2 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.n1 1.8205
R10654 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1.n3 0.595283
C0 Transmission_Gate_Layout_5.CLKB IN5 5.2e-19
C1 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_10.CLKB 0.653f
C2 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_3.CLK 0.00887f
C3 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_5.VIN 11.3f
C4 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_9.VOUT 0.482f
C5 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 0.371f
C6 Transmission_Gate_Layout_13.CLK Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT 0.237f
C7 Transmission_Gate_Layout_5.CLKB IN8 0.0182f
C8 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT VDD 0.481f
C9 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_9.CLKB 2.05e-20
C10 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT Transmission_Gate_Layout_9.CLK 0.0404f
C11 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_13.CLK 0.00172f
C12 Transmission_Gate_Layout_13.CLK OUT 0.672f
C13 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT 6.1e-20
C14 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_6.CLKB 0.00272f
C15 Transmission_Gate_Layout_19.CLKB VDD 3.74f
C16 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_12.VIN 0.0673f
C17 Transmission_Gate_Layout_3.CLK Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 0.00134f
C18 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_5.CLKB 3.1e-19
C19 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_13.CLK 0.00152f
C20 Transmission_Gate_Layout_11.VIN IN2 0.434f
C21 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_16.CLKB 0.0188f
C22 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_3.VIN 11.3f
C23 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_6.VIN 0.0402f
C24 Transmission_Gate_Layout_6.VIN EN 0.562f
C25 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_11.CLKB 8.17e-19
C26 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT Transmission_Gate_Layout_12.CLK 0.00892f
C27 Transmission_Gate_Layout_2.CLKB Transmission_Gate_Layout_13.VIN 2.18f
C28 Transmission_Gate_Layout_4.CLKB IN7 5.2e-19
C29 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_2.VIN 11.3f
C30 Transmission_Gate_Layout_6.VIN IN1 11.3f
C31 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_12.CLK 0.00352f
C32 Transmission_Gate_Layout_12.CLK OUT 0.492f
C33 Transmission_Gate_Layout_9.CLK Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT 0.00895f
C34 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 0.371f
C35 Transmission_Gate_Layout_12.VIN VDD 3.7f
C36 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_2.CLKB 6.63e-19
C37 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_12.CLK 0.00185f
C38 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_12.VIN 0.209f
C39 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_11.VIN 0.00876f
C40 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_19.CLKB 0.00265f
C41 Transmission_Gate_Layout_11.CLK Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT 0.237f
C42 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_0.CLKB 0.578f
C43 Transmission_Gate_Layout_10.CLKB Transmission_Gate_Layout_13.VIN 0.00356f
C44 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_11.CLKB 2.79e-19
C45 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_7.CLKB 0.0256f
C46 Transmission_Gate_Layout_1.VIN VDD 3.55f
C47 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_1.CLK 0.00415f
C48 Transmission_Gate_Layout_6.CLKB Transmission_Gate_Layout_3.VIN 2.19f
C49 Transmission_Gate_Layout_21.CLKB VDD 3.75f
C50 Transmission_Gate_Layout_12.CLKB Transmission_Gate_Layout_3.CLKB 0.00887f
C51 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_6.CLKB 7.47e-19
C52 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_10.VIN 0.063f
C53 Transmission_Gate_Layout_6.CLKB EN 0.00142f
C54 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT A1 0.0691f
C55 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.CLK 0.433f
C56 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_8.VIN 3.1e-19
C57 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_21.CLKB 0.00356f
C58 Transmission_Gate_Layout_11.VIN IN7 0.119f
C59 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_3.CLKB 0.323f
C60 Transmission_Gate_Layout_18.CLKB VDD 3.74f
C61 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_10.CLKB 0.0668f
C62 Transmission_Gate_Layout_6.CLKB IN1 5.2e-19
C63 Transmission_Gate_Layout_1.CLK VDD 2.03f
C64 Transmission_Gate_Layout_11.CLK Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT 0.00752f
C65 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_10.VIN 0.571f
C66 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_11.CLK 0.0948f
C67 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_5.VIN 0.0286f
C68 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_3.CLK 0.00886f
C69 Transmission_Gate_Layout_5.VIN IN6 8.72e-19
C70 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT Transmission_Gate_Layout_13.CLK 0.00751f
C71 Transmission_Gate_Layout_12.CLKB VDD 3.72f
C72 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_1.VIN 0.633f
C73 Transmission_Gate_Layout_3.CLK VDD 1.65f
C74 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_10.VIN 0.351f
C75 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_20.CLKB 0.00432f
C76 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT A1 0.0264f
C77 Transmission_Gate_Layout_19.CLKB EN 0.37f
C78 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_1.CLK 0.00394f
C79 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_6.CLKB 0.247f
C80 Transmission_Gate_Layout_3.CLK Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 0.0365f
C81 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_3.CLKB 0.00422f
C82 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_4.VIN 0.00307f
C83 Transmission_Gate_Layout_13.VIN Transmission_Gate_Layout_12.VIN 0.23f
C84 Transmission_Gate_Layout_7.CLKB IN2 5.2e-19
C85 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_10.CLKB 0.329f
C86 Transmission_Gate_Layout_11.VIN IN4 11.3f
C87 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 C1 0.00102f
C88 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT 0.0311f
C89 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_6.CLKB 0.0819f
C90 Transmission_Gate_Layout_8.CLKB Transmission_Gate_Layout_12.VIN 0.00356f
C91 VDD IN2 0.115f
C92 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_12.VIN 0.0978f
C93 Transmission_Gate_Layout_5.VIN Transmission_Gate_Layout_8.VIN 0.0157f
C94 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_10.CLKB 0.0141f
C95 Transmission_Gate_Layout_20.CLKB Transmission_Gate_Layout_5.VIN 2.19f
C96 Transmission_Gate_Layout_2.VIN VDD 3.46f
C97 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_8.CLKB 0.0706f
C98 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT C1 0.0264f
C99 Transmission_Gate_Layout_8.CLKB Transmission_Gate_Layout_21.CLKB 7.68e-19
C100 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.VIN 12f
C101 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_13.VIN 0.485f
C102 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT 0.0323f
C103 Transmission_Gate_Layout_5.VIN IN4 0.00819f
C104 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_12.VIN 3.88e-19
C105 Transmission_Gate_Layout_1.VIN EN 3.75e-20
C106 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_4.CLKB 0.0321f
C107 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_6.CLKB 5.56e-19
C108 Transmission_Gate_Layout_21.CLKB EN 0.333f
C109 Transmission_Gate_Layout_15.CLKB VDD 3.76f
C110 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_3.VIN 0.00432f
C111 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 Transmission_Gate_Layout_1.CLK 0.00134f
C112 Transmission_Gate_Layout_19.CLKB IN5 0.0173f
C113 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_18.CLKB 2.19f
C114 Transmission_Gate_Layout_18.CLKB EN 0.216f
C115 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_1.CLK 0.0475f
C116 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_12.CLK 2.96f
C117 VDD IN6 0.143f
C118 Transmission_Gate_Layout_12.CLKB Transmission_Gate_Layout_13.VIN 0.0092f
C119 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_13.VIN 0.725f
C120 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT 0.0311f
C121 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1 0.371f
C122 Transmission_Gate_Layout_19.CLKB IN8 5.2e-19
C123 VDD IN7 0.119f
C124 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_12.VIN 0.00378f
C125 Transmission_Gate_Layout_12.VIN OUT 11.3f
C126 Transmission_Gate_Layout_1.CLK Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 0.0366f
C127 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLK 0.533f
C128 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_12.VIN 3.27e-19
C129 Transmission_Gate_Layout_3.CLK EN 0.0129f
C130 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_1.CLKB 0.0321f
C131 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_11.VIN 0.00872f
C132 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_9.VIN 2.19f
C133 Transmission_Gate_Layout_14.CLKB VDD 3.75f
C134 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_1.VIN 0.532f
C135 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_14.CLKB 2.18f
C136 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_12.VIN 0.00404f
C137 VDD C1 0.476f
C138 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_12.CLKB 0.0141f
C139 Transmission_Gate_Layout_8.VIN VDD 2.12f
C140 VDD IN3 0.143f
C141 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_1.VIN 0.772f
C142 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_1.CLK 0.0205f
C143 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_13.VIN 11.5f
C144 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_21.CLKB 0.014f
C145 Transmission_Gate_Layout_10.VIN IN3 11.3f
C146 Transmission_Gate_Layout_9.VIN IN7 0.0353f
C147 Transmission_Gate_Layout_20.CLKB VDD 3.75f
C148 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_11.CLK 0.00142f
C149 Transmission_Gate_Layout_10.CLKB Transmission_Gate_Layout_9.VOUT 2.05e-20
C150 Transmission_Gate_Layout_7.VIN IN2 11.3f
C151 EN IN2 0.425f
C152 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_1.CLK 0.141f
C153 Transmission_Gate_Layout_1.VIN IN8 2.33e-19
C154 Transmission_Gate_Layout_3.CLK Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT 0.00751f
C155 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT 0.0189f
C156 IN2 IN1 4.9f
C157 VDD IN4 0.176f
C158 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_11.CLKB 0.0748f
C159 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_2.VIN 1f
C160 Transmission_Gate_Layout_12.CLKB OUT 2.18f
C161 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_3.CLK 1.28f
C162 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1 VDD 0.85f
C163 VDD B1 0.479f
C164 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_1.VIN 11.3f
C165 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_8.VIN 0.0257f
C166 Transmission_Gate_Layout_8.CLKB IN6 0.0187f
C167 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_3.CLK 0.0306f
C168 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 0.371f
C169 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_17.CLKB 7.68e-19
C170 Transmission_Gate_Layout_15.CLKB EN 0.314f
C171 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 B1 0.00102f
C172 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_11.CLKB 0.031f
C173 Transmission_Gate_Layout_0.CLKB Transmission_Gate_Layout_12.VIN 2.18f
C174 EN IN6 0.605f
C175 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT Transmission_Gate_Layout_13.CLK 0.0404f
C176 Transmission_Gate_Layout_9.VIN IN4 4.29e-19
C177 EN IN7 0.541f
C178 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 VDD 0.847f
C179 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_0.CLKB 6.63e-19
C180 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_2.VIN 0.69f
C181 IN2 IN5 8.14e-19
C182 IN1 IN7 3.58f
C183 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_5.VIN 0.00197f
C184 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_12.VIN 11.5f
C185 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_2.VIN 0.472f
C186 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_8.CLKB 0.48f
C187 Transmission_Gate_Layout_14.CLKB EN 0.304f
C188 Transmission_Gate_Layout_5.CLKB Transmission_Gate_Layout_1.VIN 2.18f
C189 Transmission_Gate_Layout_1.CLK Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT 0.00892f
C190 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_2.VIN 2.18f
C191 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.VOUT 1.02f
C192 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_6.CLKB 0.484f
C193 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_21.CLKB 4.32e-20
C194 EN IN3 0.57f
C195 Transmission_Gate_Layout_8.VIN EN 0.525f
C196 Transmission_Gate_Layout_17.CLKB VDD 3.75f
C197 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_11.CLK 0.00142f
C198 Transmission_Gate_Layout_20.CLKB EN 0.334f
C199 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_12.VIN 0.125f
C200 Transmission_Gate_Layout_15.CLKB IN5 0.466f
C201 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_0.CLKB 0.297f
C202 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_9.VOUT 0.00626f
C203 Transmission_Gate_Layout_11.CLK IN6 0.0496f
C204 Transmission_Gate_Layout_3.CLK Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT 0.237f
C205 EN IN4 0.675f
C206 IN8 IN6 3.12e-19
C207 IN7 IN5 2.21f
C208 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT C1 5.36e-19
C209 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 B1 6.1e-20
C210 Transmission_Gate_Layout_10.CLKB Transmission_Gate_Layout_2.CLKB 0.0321f
C211 Transmission_Gate_Layout_1.CLKB VDD 3.75f
C212 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_9.VOUT 0.544f
C213 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_13.CLK 0.979f
C214 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_12.VIN 0.494f
C215 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_1.CLKB 0.0127f
C216 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_9.VIN 0.0205f
C217 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_15.CLKB 0.00265f
C218 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_11.VIN 0.00872f
C219 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT 0.00563f
C220 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_8.VIN 4.74e-19
C221 Transmission_Gate_Layout_4.CLKB VDD 3.75f
C222 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 B1 0.167f
C223 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_8.VIN 0.588f
C224 Transmission_Gate_Layout_4.VIN IN7 11.3f
C225 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_12.CLKB 0.0708f
C226 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_20.CLKB 0.0142f
C227 Transmission_Gate_Layout_9.CLKB VDD 3.75f
C228 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_13.CLK 0.642f
C229 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_3.CLKB 5.2e-19
C230 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.CLKB 0.0211f
C231 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_12.CLK 0.0846f
C232 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_1.CLKB 5.2e-19
C233 Transmission_Gate_Layout_8.VIN IN8 8.72e-19
C234 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT Transmission_Gate_Layout_1.CLK 0.00752f
C235 Transmission_Gate_Layout_20.CLKB IN8 0.528f
C236 IN5 IN4 2.88e-19
C237 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_7.CLKB 0.121f
C238 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_5.CLKB 0.0256f
C239 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_1.VIN 6.05e-20
C240 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_4.CLKB 0.181f
C241 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_12.CLKB 0.316f
C242 IN4 IN8 0.00961f
C243 Transmission_Gate_Layout_11.VIN VDD 1.87f
C244 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_12.CLK 0.0322f
C245 Transmission_Gate_Layout_2.CLKB Transmission_Gate_Layout_12.VIN 0.0716f
C246 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLKB 0.466f
C247 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_6.VIN 2.05e-20
C248 Transmission_Gate_Layout_1.CLK Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT 0.237f
C249 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_10.VIN 0.0257f
C250 Transmission_Gate_Layout_17.CLKB EN 0.314f
C251 Transmission_Gate_Layout_9.VOUT IN6 2.42e-19
C252 Transmission_Gate_Layout_17.CLKB IN1 0.0174f
C253 Transmission_Gate_Layout_0.CLKB Transmission_Gate_Layout_14.CLKB 7.68e-19
C254 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_13.VIN 2.05e-20
C255 Transmission_Gate_Layout_9.CLK Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 0.0365f
C256 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 VDD 0.847f
C257 Transmission_Gate_Layout_0.CLKB IN3 0.0182f
C258 Transmission_Gate_Layout_10.CLKB Transmission_Gate_Layout_12.VIN 0.00426f
C259 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_0.CLKB 5.2e-19
C260 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT Transmission_Gate_Layout_3.CLK 0.00895f
C261 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_2.CLKB 0.289f
C262 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_11.VIN 0.0751f
C263 Transmission_Gate_Layout_5.VIN VDD 2.29f
C264 Transmission_Gate_Layout_6.CLKB Transmission_Gate_Layout_1.VIN 2.05e-20
C265 Transmission_Gate_Layout_5.CLKB Transmission_Gate_Layout_8.VIN 0.0043f
C266 A1 B1 0.0224f
C267 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_8.CLKB 0.0141f
C268 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_3.VIN 2.05e-20
C269 Transmission_Gate_Layout_5.CLKB Transmission_Gate_Layout_20.CLKB 7.68e-19
C270 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT VDD 0.564f
C271 Transmission_Gate_Layout_3.CLK Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT 0.0404f
C272 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.VIN 11.3f
C273 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_2.CLKB 0.0812f
C274 Transmission_Gate_Layout_16.CLKB VDD 3.76f
C275 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_10.CLKB 0.0836f
C276 Transmission_Gate_Layout_6.VIN IN2 6.78e-19
C277 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT B1 5.36e-19
C278 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_5.VIN 0.0664f
C279 Transmission_Gate_Layout_13.CLK C1 1.06e-21
C280 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 A1 0.00102f
C281 Transmission_Gate_Layout_3.CLKB VDD 3.75f
C282 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT VDD 0.547f
C283 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_3.VIN 0.443f
C284 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.VIN 0.592f
C285 Transmission_Gate_Layout_11.VIN EN 1.49f
C286 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_4.VIN 2.19f
C287 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_4.CLKB 0.228f
C288 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_2.CLKB 0.571f
C289 Transmission_Gate_Layout_11.VIN IN1 0.123f
C290 Transmission_Gate_Layout_7.CLKB VDD 3.75f
C291 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.CLKB 0.23f
C292 Transmission_Gate_Layout_12.CLK C1 0.0401f
C293 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_12.VIN 11.5f
C294 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_4.CLKB 0.0818f
C295 Transmission_Gate_Layout_6.VIN IN7 2.12e-19
C296 Transmission_Gate_Layout_10.VIN VDD 2.39f
C297 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_12.VIN 1.02f
C298 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 VDD 0.847f
C299 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_10.CLKB 2.19f
C300 Transmission_Gate_Layout_5.VIN EN 0.519f
C301 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_9.CLK 0.0833f
C302 Transmission_Gate_Layout_12.CLK Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1 0.0366f
C303 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLK 0.438f
C304 Transmission_Gate_Layout_12.CLKB Transmission_Gate_Layout_12.VIN 0.491f
C305 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_4.CLKB 0.479f
C306 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.SD1 0.254f
C307 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_12.VIN 0.717f
C308 Transmission_Gate_Layout_9.VIN VDD 2.47f
C309 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_3.VIN 0.00432f
C310 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLK 0.803f
C311 Transmission_Gate_Layout_11.VIN IN5 0.111f
C312 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_10.VIN 0.00819f
C313 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_16.CLKB 2.05e-20
C314 Transmission_Gate_Layout_16.CLKB EN 0.315f
C315 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 0.371f
C316 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_0.CLKB 0.0141f
C317 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_13.VIN 2.19f
C318 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_11.CLKB 0.466f
C319 Transmission_Gate_Layout_16.CLKB IN1 0.466f
C320 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_3.CLK 0.129f
C321 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_5.VIN 2.98e-19
C322 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT B1 0.0264f
C323 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_3.CLKB 0.555f
C324 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_3.CLK 2.89f
C325 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_19.CLKB 7.68e-19
C326 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT 0.0323f
C327 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_1.CLKB 0.00422f
C328 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_11.VIN 0.0751f
C329 Transmission_Gate_Layout_13.VIN VDD 3.3f
C330 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_5.VIN 0.588f
C331 Transmission_Gate_Layout_5.VIN IN5 0.0278f
C332 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_13.VIN 0.349f
C333 Transmission_Gate_Layout_2.VIN Transmission_Gate_Layout_12.VIN 0.124f
C334 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_3.VIN 2.19f
C335 Transmission_Gate_Layout_8.CLKB VDD 3.75f
C336 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_5.CLKB 0.0141f
C337 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_7.CLKB 0.483f
C338 Transmission_Gate_Layout_7.CLKB EN 0.00142f
C339 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_9.CLK 0.00142f
C340 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_12.CLKB 7.37e-19
C341 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT B1 0.0691f
C342 Transmission_Gate_Layout_5.VIN IN8 11.3f
C343 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 VDD 0.847f
C344 Transmission_Gate_Layout_3.VIN VDD 3.54f
C345 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT C1 0.0691f
C346 Transmission_Gate_Layout_18.CLKB IN2 0.466f
C347 Transmission_Gate_Layout_7.VIN VDD 1.81f
C348 VDD EN 3.84f
C349 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_10.VIN 0.186f
C350 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_9.VOUT 2.18f
C351 Transmission_Gate_Layout_10.VIN EN 0.49f
C352 VDD IN1 0.119f
C353 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_5.VIN 0.0263f
C354 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_2.VIN 0.595f
C355 Transmission_Gate_Layout_3.CLKB OUT 7.69e-21
C356 Transmission_Gate_Layout_13.CLKB VDD 3.76f
C357 Transmission_Gate_Layout_15.CLKB Transmission_Gate_Layout_1.VIN 0.00432f
C358 Transmission_Gate_Layout_9.CLK Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT 0.237f
C359 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 VDD 0.847f
C360 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_8.CLKB 3.1e-19
C361 Transmission_Gate_Layout_19.CLKB Transmission_Gate_Layout_20.CLKB 0.0256f
C362 Transmission_Gate_Layout_21.CLKB IN6 0.528f
C363 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_7.CLKB 0.00145f
C364 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT VDD 0.554f
C365 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT Transmission_Gate_Layout_11.CLK 0.00892f
C366 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_3.VIN 0.00104f
C367 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_3.CLKB 0.0321f
C368 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_17.CLKB 0.00265f
C369 Transmission_Gate_Layout_9.VIN EN 0.567f
C370 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_4.VIN 4.32e-20
C371 Transmission_Gate_Layout_14.CLKB Transmission_Gate_Layout_12.VIN 4.32e-20
C372 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_2.VIN 0.136f
C373 Transmission_Gate_Layout_19.CLKB IN4 0.497f
C374 Transmission_Gate_Layout_9.CLK VDD 2.1f
C375 VDD OUT 3.4f
C376 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_7.CLKB 0.349f
C377 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_10.VIN 0.79f
C378 Transmission_Gate_Layout_12.VIN IN3 3.52e-19
C379 Transmission_Gate_Layout_11.CLK VDD 2.38f
C380 VDD IN5 0.119f
C381 Transmission_Gate_Layout_21.CLKB Transmission_Gate_Layout_14.CLKB 0.0321f
C382 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_10.VIN 2.98e-19
C383 Transmission_Gate_Layout_5.CLKB Transmission_Gate_Layout_5.VIN 0.527f
C384 Transmission_Gate_Layout_11.CLKB VDD 3.75f
C385 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_10.VIN 3.1e-19
C386 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_13.VIN 11.5f
C387 VDD IN8 0.143f
C388 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_8.VIN 0.0873f
C389 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_21.CLKB 2.18f
C390 Transmission_Gate_Layout_21.CLKB IN3 5.2e-19
C391 Transmission_Gate_Layout_20.CLKB Transmission_Gate_Layout_1.VIN 4.32e-20
C392 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.CLK 0.605f
C393 Transmission_Gate_Layout_8.CLKB EN 2.98e-19
C394 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT A1 5.36e-19
C395 Transmission_Gate_Layout_13.CLK Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 0.0365f
C396 Transmission_Gate_Layout_4.VIN VDD 2.26f
C397 Transmission_Gate_Layout_13.CLKB Transmission_Gate_Layout_13.VIN 0.466f
C398 Transmission_Gate_Layout_2.CLKB Transmission_Gate_Layout_1.CLKB 0.0188f
C399 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_11.CLK 0.0657f
C400 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_3.VIN 11.4f
C401 Transmission_Gate_Layout_3.VIN EN 7.5e-20
C402 Transmission_Gate_Layout_9.VIN IN5 11.3f
C403 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_14.CLKB 0.0142f
C404 Transmission_Gate_Layout_7.VIN EN 0.437f
C405 Transmission_Gate_Layout_7.VIN IN1 6.05e-20
C406 EN IN1 0.541f
C407 IN2 IN7 0.00148f
C408 Transmission_Gate_Layout_3.CLK IN3 0.0308f
C409 VDD A1 0.477f
C410 Transmission_Gate_Layout_13.CLK Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT 0.00895f
C411 Transmission_Gate_Layout_1.CLK B1 0.0401f
C412 Transmission_Gate_Layout_13.VIN OUT 11.4f
C413 Transmission_Gate_Layout_0.CLKB VDD 3.75f
C414 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_0.CLKB 0.0114f
C415 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.VIN 0.522f
C416 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_11.VIN 0.0751f
C417 Transmission_Gate_Layout_6.CLKB Transmission_Gate_Layout_4.CLKB 0.0194f
C418 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT VDD 0.553f
C419 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_3.VIN 0.616f
C420 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_8.CLKB 0.246f
C421 Transmission_Gate_Layout_11.CLKB Transmission_Gate_Layout_13.VIN 0.00356f
C422 Transmission_Gate_Layout_15.CLKB IN7 0.0174f
C423 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_9.CLK 3.58e-19
C424 Transmission_Gate_Layout_9.CLK EN 0.00132f
C425 Transmission_Gate_Layout_5.CLKB VDD 3.76f
C426 Transmission_Gate_Layout_3.CLK B1 1.06e-21
C427 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 0.371f
C428 Transmission_Gate_Layout_10.CLKB Transmission_Gate_Layout_9.CLKB 0.0194f
C429 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_3.CLKB 2.05e-19
C430 Transmission_Gate_Layout_12.CLK Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.OUT 0.237f
C431 Transmission_Gate_Layout_11.CLK Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 0.0366f
C432 Transmission_Gate_Layout_9.VOUT VDD 3.47f
C433 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_3.VIN 0.855f
C434 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT 0.0311f
C435 Transmission_Gate_Layout_7.VIN Transmission_Gate_Layout_11.CLK 0.482f
C436 Transmission_Gate_Layout_11.CLK EN 0.1f
C437 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_9.VOUT 0.0704f
C438 EN IN5 0.544f
C439 Transmission_Gate_Layout_3.VIN Transmission_Gate_Layout_11.CLKB 0.0887f
C440 Transmission_Gate_Layout_13.CLKB OUT 2.26f
C441 IN1 IN5 0.0015f
C442 Transmission_Gate_Layout_14.CLKB IN6 5.2e-19
C443 EN IN8 0.605f
C444 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_1.VIN 0.00356f
C445 Transmission_Gate_Layout_11.CLK Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 0.00134f
C446 Non_Ovl_CLK_Gen_Layout_1.Inverter_Layout_2.OUT VDD 0.478f
C447 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 6.1e-20
C448 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_5.CLKB 0.0423f
C449 Transmission_Gate_Layout_13.CLK VDD 1.06f
C450 Transmission_Gate_Layout_8.VIN IN6 11.3f
C451 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_3.CLKB 4.84e-19
C452 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_10.CLKB 3.1e-19
C453 Transmission_Gate_Layout_1.CLKB Transmission_Gate_Layout_12.VIN 2.2f
C454 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_3.VIN 6.78e-19
C455 Transmission_Gate_Layout_9.VIN Transmission_Gate_Layout_9.VOUT 11.3f
C456 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_6.VIN 2.19f
C457 Transmission_Gate_Layout_4.VIN EN 0.562f
C458 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 Transmission_Gate_Layout_13.CLK 0.00134f
C459 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT 0.0323f
C460 Transmission_Gate_Layout_4.VIN IN1 6.27e-19
C461 Transmission_Gate_Layout_15.CLKB IN4 1.97e-19
C462 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_11.CLK 2.43f
C463 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_1.CLKB 0.575f
C464 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.SD1 A1 0.167f
C465 Transmission_Gate_Layout_8.CLKB Transmission_Gate_Layout_0.CLKB 0.0321f
C466 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_11.CLKB 0.0781f
C467 Transmission_Gate_Layout_12.CLK VDD 1.2f
C468 Transmission_Gate_Layout_14.CLKB IN3 0.528f
C469 Transmission_Gate_Layout_8.VIN Transmission_Gate_Layout_14.CLKB 0.00356f
C470 Transmission_Gate_Layout_9.CLKB Transmission_Gate_Layout_12.VIN 0.00828f
C471 Transmission_Gate_Layout_19.CLKB Transmission_Gate_Layout_11.VIN 2.19f
C472 Non_Ovl_CLK_Gen_Layout_1.NOR_Layout_0.OUT VDD 0.553f
C473 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_1.CLKB 0.282f
C474 Transmission_Gate_Layout_0.CLKB EN 2.98e-19
C475 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_11.CLKB 0.246f
C476 Transmission_Gate_Layout_4.CLKB Transmission_Gate_Layout_1.VIN 2.18f
C477 Non_Ovl_CLK_Gen_Layout_0.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.SD1 0.254f
C478 Transmission_Gate_Layout_11.CLK IN8 0.0572f
C479 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.SD1 A1 6.1e-20
C480 Transmission_Gate_Layout_1.VIN Transmission_Gate_Layout_9.CLKB 0.11f
C481 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_7.CLKB 7.47e-19
C482 Transmission_Gate_Layout_16.CLKB Transmission_Gate_Layout_6.CLKB 0.0256f
C483 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_9.CLK 0.422f
C484 Transmission_Gate_Layout_9.VOUT Transmission_Gate_Layout_8.CLKB 2.19f
C485 Transmission_Gate_Layout_3.CLKB Transmission_Gate_Layout_2.CLKB 0.0141f
C486 Transmission_Gate_Layout_5.CLKB EN 0.00172f
C487 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_0.OUT VDD 0.553f
C488 Transmission_Gate_Layout_3.CLK Transmission_Gate_Layout_1.CLKB 0.0819f
C489 Transmission_Gate_Layout_1.CLK Transmission_Gate_Layout_9.CLKB 0.00717f
C490 Transmission_Gate_Layout_6.VIN VDD 2.27f
C491 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_12.VIN 0.00455f
C492 Transmission_Gate_Layout_4.VIN Transmission_Gate_Layout_11.CLK 0.079f
C493 Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_0.SD1 C1 0.167f
C494 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_10.VIN 0.00347f
C495 Transmission_Gate_Layout_4.VIN IN5 2.12e-19
C496 Transmission_Gate_Layout_19.CLKB Transmission_Gate_Layout_5.VIN 0.00432f
C497 Transmission_Gate_Layout_20.CLKB IN4 0.0117f
C498 B1 C1 0.0135f
C499 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_13.VIN 0.678f
C500 Transmission_Gate_Layout_9.CLK A1 1.06e-21
C501 Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.OUT Non_Ovl_CLK_Gen_Layout_0.NOR_Layout_1.OUT 0.0189f
C502 Transmission_Gate_Layout_11.CLK A1 0.0401f
C503 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT VDD 0.481f
C504 Transmission_Gate_Layout_2.CLKB VDD 3.75f
C505 Transmission_Gate_Layout_10.VIN Transmission_Gate_Layout_2.CLKB 0.196f
C506 Transmission_Gate_Layout_17.CLKB Transmission_Gate_Layout_15.CLKB 7.68e-19
C507 Transmission_Gate_Layout_18.CLKB Transmission_Gate_Layout_11.VIN 0.12f
C508 Transmission_Gate_Layout_11.VIN Transmission_Gate_Layout_1.CLK 0.0556f
C509 Transmission_Gate_Layout_7.CLKB Transmission_Gate_Layout_6.CLKB 0.0141f
C510 Non_Ovl_CLK_Gen_Layout_2.Inverter_Layout_2.OUT Non_Ovl_CLK_Gen_Layout_2.NOR_Layout_1.SD1 0.254f
C511 Transmission_Gate_Layout_6.VIN Transmission_Gate_Layout_9.VIN 1.41e-20
C512 Transmission_Gate_Layout_12.CLK Transmission_Gate_Layout_13.VIN 0.0545f
C513 Transmission_Gate_Layout_6.CLKB VDD 3.76f
C514 Transmission_Gate_Layout_9.CLK Transmission_Gate_Layout_9.VOUT 0.464f
C515 Transmission_Gate_Layout_13.CLK Transmission_Gate_Layout_13.CLKB 0.297f
C516 Transmission_Gate_Layout_17.CLKB IN7 0.466f
C517 Transmission_Gate_Layout_10.CLKB VDD 3.75f
C518 Transmission_Gate_Layout_11.CLK Transmission_Gate_Layout_5.CLKB 0.328f
.ends

