magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1019 -1409 1019 1409
<< metal1 >>
rect -19 403 19 409
rect -19 -403 -13 403
rect 13 -403 19 403
rect -19 -409 19 -403
<< via1 >>
rect -13 -403 13 403
<< metal2 >>
rect -19 403 19 409
rect -19 -403 -13 403
rect 13 -403 19 403
rect -19 -409 19 -403
<< end >>
