magic
tech gf180mcuC
magscale 1 10
timestamp 1695206022
<< nwell >>
rect 3181 4618 3351 4783
rect 3181 4547 6156 4618
rect 3181 4481 6634 4547
rect 3181 4375 3216 4481
rect 6003 4477 6634 4481
rect 6003 4375 6244 4477
rect 6003 4374 6291 4375
rect 2523 3501 2575 3560
rect 74 2187 3045 2518
<< metal1 >>
rect 2690 6570 5918 6783
rect 2275 6181 2457 6233
rect 2275 6120 2313 6181
rect 2403 6120 2457 6181
rect 2275 6077 2457 6120
rect 2696 4537 2805 6570
rect 5627 6245 5701 6265
rect 5627 6188 5633 6245
rect 5688 6188 5701 6245
rect 5627 6175 5701 6188
rect 5623 5745 5704 5759
rect 5623 5687 5638 5745
rect 5690 5687 5704 5745
rect 5623 5672 5704 5687
rect 6824 5507 8983 5679
rect 8634 5409 8983 5507
rect 5619 5172 5700 5186
rect 5619 5113 5632 5172
rect 5688 5113 5700 5172
rect 6492 5121 6607 5158
rect 5619 5099 5700 5113
rect 6045 5049 6607 5121
rect 6492 5028 6607 5049
rect 8924 4919 9125 4977
rect 72 4367 2805 4537
rect 3181 4618 3351 4783
rect 3181 4547 6156 4618
rect 3181 4481 6634 4547
rect 3181 4375 3216 4481
rect 6003 4477 6634 4481
rect 6003 4375 6244 4477
rect 6003 4374 6291 4375
rect 2696 4353 2805 4367
rect 2506 4044 2581 4059
rect 2506 3985 2518 4044
rect 2570 3985 2581 4044
rect 2506 3973 2581 3985
rect 2514 3560 2580 3568
rect 2514 3501 2523 3560
rect 2575 3501 2580 3560
rect 2514 3487 2580 3501
rect 3155 3221 3287 3227
rect 2929 3218 3534 3221
rect 2929 3117 3172 3218
rect 3273 3117 3534 3218
rect 2929 3112 3534 3117
rect 3155 3097 3287 3112
rect 2515 2962 2581 2974
rect 2515 2905 2517 2962
rect 2569 2905 2581 2962
rect 2515 2893 2581 2905
rect 2992 2909 3063 2925
rect 2992 2850 3006 2909
rect 3058 2850 3063 2909
rect 2992 2838 3063 2850
rect 74 2287 3045 2518
rect 74 2187 3702 2287
rect 3043 2131 3702 2187
rect 6183 2127 6800 2292
rect 70 1856 154 1863
rect 70 1801 82 1856
rect 147 1801 154 1856
rect 70 1789 154 1801
rect 529 1799 611 1813
rect 529 1741 545 1799
rect 597 1741 611 1799
rect 529 1727 611 1741
rect 3250 1791 3348 1803
rect 3250 1724 3263 1791
rect 3335 1724 3348 1791
rect 6365 1788 6448 1797
rect 3250 1717 3348 1724
rect 3752 1734 3829 1749
rect 3752 1680 3764 1734
rect 3823 1680 3829 1734
rect 6365 1727 6377 1788
rect 6436 1727 6448 1788
rect 6365 1722 6448 1727
rect 6845 1734 6928 1748
rect 3752 1668 3829 1680
rect 6845 1666 6858 1734
rect 6916 1666 6928 1734
rect 6845 1653 6928 1666
rect 3156 1521 3316 1536
rect 3156 1436 3174 1521
rect 3259 1436 3316 1521
rect 3156 1416 3316 1436
rect 526 1203 604 1211
rect 526 1140 534 1203
rect 595 1140 604 1203
rect 526 1134 604 1140
rect 531 733 609 745
rect 531 681 545 733
rect 597 681 609 733
rect 531 668 609 681
rect 3744 654 3837 664
rect 3744 589 3759 654
rect 3825 589 3837 654
rect 6853 659 6923 668
rect 6853 604 6861 659
rect 6914 604 6923 659
rect 6853 595 6923 604
rect 3744 577 3837 589
rect 313 105 9354 294
<< via1 >>
rect 2313 6120 2403 6181
rect 5633 6188 5688 6245
rect 4619 6104 4671 6156
rect 5638 5687 5690 5745
rect 5632 5113 5688 5172
rect 2518 3985 2570 4044
rect 1489 3896 1541 3948
rect 2523 3501 2575 3560
rect 3172 3117 3273 3218
rect 2517 2905 2569 2962
rect 3006 2850 3058 2909
rect 4254 2190 4332 2246
rect 82 1801 147 1856
rect 545 1741 597 1799
rect 3263 1724 3335 1791
rect 3764 1680 3823 1734
rect 6377 1727 6436 1788
rect 6858 1666 6916 1734
rect 3174 1436 3259 1521
rect 534 1140 595 1203
rect 3760 1086 3826 1151
rect 6855 1082 6920 1156
rect 1573 759 1625 811
rect 545 681 597 733
rect 4785 690 4841 744
rect 7879 692 7931 744
rect 3759 589 3825 654
rect 6861 604 6914 659
<< metal2 >>
rect 5627 6245 5701 6265
rect 2275 6205 2457 6233
rect 2275 6110 2307 6205
rect 2431 6110 2457 6205
rect 5627 6188 5633 6245
rect 5688 6188 5701 6245
rect 5627 6175 5701 6188
rect 2275 6077 2457 6110
rect 4603 6162 4700 6169
rect 4603 6104 4615 6162
rect 4679 6104 4700 6162
rect 4603 6092 4700 6104
rect 5627 5759 5693 6175
rect 5623 5745 5704 5759
rect 5623 5687 5638 5745
rect 5690 5687 5704 5745
rect 5623 5672 5704 5687
rect 3356 5171 3412 5247
rect 5627 5186 5693 5672
rect 3003 5115 3412 5171
rect 5619 5172 5700 5186
rect 2506 4044 2581 4059
rect 2506 3985 2518 4044
rect 2570 3985 2581 4044
rect 2506 3973 2581 3985
rect 1481 3951 1617 3956
rect 1481 3948 1498 3951
rect 1481 3896 1489 3948
rect 1481 3887 1498 3896
rect 1603 3887 1617 3951
rect 1481 3883 1617 3887
rect 2515 3568 2575 3973
rect 2514 3560 2580 3568
rect 2514 3501 2523 3560
rect 2575 3501 2580 3560
rect 2514 3487 2580 3501
rect 245 2969 301 3041
rect 97 2913 301 2969
rect 2515 2974 2575 3487
rect 2515 2962 2581 2974
rect 97 1863 153 2913
rect 2515 2905 2517 2962
rect 2569 2905 2581 2962
rect 3003 2925 3059 5115
rect 5619 5113 5632 5172
rect 5688 5113 5700 5172
rect 5619 5099 5700 5113
rect 3155 3218 3287 3227
rect 3155 3117 3164 3218
rect 3273 3117 3287 3218
rect 3155 3097 3287 3117
rect 2515 2893 2581 2905
rect 2992 2909 3063 2925
rect 2992 2850 3006 2909
rect 3058 2850 3063 2909
rect 2992 2838 3063 2850
rect 4267 2255 4323 2545
rect 6964 2259 7020 3012
rect 4233 2246 4346 2255
rect 4233 2190 4254 2246
rect 4332 2190 4346 2246
rect 6964 2203 9342 2259
rect 4233 2178 4346 2190
rect 70 1856 154 1863
rect 70 1801 82 1856
rect 147 1801 154 1856
rect 70 1789 154 1801
rect 529 1799 611 1813
rect 529 1741 545 1799
rect 597 1741 611 1799
rect 3250 1796 3348 1803
rect 529 1727 611 1741
rect 2818 1791 3348 1796
rect 2818 1740 3263 1791
rect 534 1211 603 1727
rect 2818 1685 2874 1740
rect 3250 1724 3263 1740
rect 3335 1724 3348 1791
rect 6365 1788 6449 1797
rect 3250 1717 3348 1724
rect 3758 1734 3829 1747
rect 3758 1680 3764 1734
rect 3823 1680 3829 1734
rect 6365 1727 6377 1788
rect 6436 1727 6449 1788
rect 6365 1723 6449 1727
rect 3156 1521 3316 1536
rect 3156 1436 3174 1521
rect 3259 1436 3316 1521
rect 3156 1416 3316 1436
rect 526 1203 604 1211
rect 526 1140 534 1203
rect 595 1140 604 1203
rect 526 1134 604 1140
rect 3758 1151 3829 1680
rect 6044 1667 6449 1723
rect 6853 1734 6923 1746
rect 6044 1600 6100 1667
rect 6853 1666 6858 1734
rect 6916 1666 6923 1734
rect 9286 1726 9342 2203
rect 534 745 603 1134
rect 3758 1086 3760 1151
rect 3826 1086 3829 1151
rect 1545 813 1637 820
rect 1545 757 1555 813
rect 1625 757 1637 813
rect 1545 753 1637 757
rect 531 733 609 745
rect 531 681 545 733
rect 597 681 609 733
rect 531 668 609 681
rect 3758 664 3829 1086
rect 6853 1156 6923 1666
rect 9137 1670 9342 1726
rect 9137 1598 9193 1670
rect 6853 1082 6855 1156
rect 6920 1082 6923 1156
rect 4766 748 4857 760
rect 4766 682 4776 748
rect 4848 682 4857 748
rect 4766 671 4857 682
rect 3744 654 3837 664
rect 3744 589 3759 654
rect 3825 589 3837 654
rect 6853 659 6923 1082
rect 7855 745 7946 754
rect 7855 678 7867 745
rect 7936 678 7946 745
rect 7855 665 7946 678
rect 6853 604 6861 659
rect 6914 604 6923 659
rect 6853 595 6923 604
rect 3744 577 3837 589
<< via2 >>
rect 2307 6181 2431 6205
rect 2307 6120 2313 6181
rect 2313 6120 2403 6181
rect 2403 6120 2431 6181
rect 2307 6110 2431 6120
rect 4615 6156 4679 6162
rect 4615 6104 4619 6156
rect 4619 6104 4671 6156
rect 4671 6104 4679 6156
rect 1498 3948 1603 3951
rect 1498 3896 1541 3948
rect 1541 3896 1603 3948
rect 1498 3887 1603 3896
rect 3164 3117 3172 3218
rect 3172 3117 3270 3218
rect 3174 1436 3259 1521
rect 1555 811 1625 813
rect 1555 759 1573 811
rect 1573 759 1625 811
rect 1555 757 1625 759
rect 4776 744 4848 748
rect 4776 690 4785 744
rect 4785 690 4841 744
rect 4841 690 4848 744
rect 4776 682 4848 690
rect 7867 744 7936 745
rect 7867 692 7879 744
rect 7879 692 7931 744
rect 7931 692 7936 744
rect 7867 678 7936 692
<< metal3 >>
rect 2275 6205 2457 6233
rect 2275 6110 2307 6205
rect 2431 6195 2457 6205
rect 2431 6162 6411 6195
rect 2431 6110 4615 6162
rect 2275 6104 4615 6110
rect 4679 6104 6411 6162
rect 2275 6099 6411 6104
rect 2275 6077 2457 6099
rect 1481 3951 1617 3956
rect 1481 3887 1498 3951
rect 1603 3887 1617 3951
rect 1481 3883 1617 3887
rect 1547 823 1617 3883
rect 3155 3218 3287 3227
rect 3155 3117 3164 3218
rect 3270 3117 3287 3218
rect 3155 3097 3287 3117
rect 3169 1536 3266 3097
rect 6314 2895 6410 6099
rect 6303 2821 6419 2895
rect 3156 1521 3316 1536
rect 3156 1436 3174 1521
rect 3259 1436 3316 1521
rect 3156 1416 3316 1436
rect 1547 820 1659 823
rect 1545 813 1659 820
rect 1545 757 1555 813
rect 1625 757 1659 813
rect 1545 753 1659 757
rect 1547 752 1659 753
rect 6314 752 6410 2821
rect 1547 748 7967 752
rect 1547 682 4776 748
rect 4848 745 7967 748
rect 4848 682 7867 745
rect 1547 678 7867 682
rect 7936 678 7967 745
rect 1547 656 7967 678
use CLK_div_3_mag  CLK_div_3_mag_0
timestamp 1695206022
transform 1 0 3185 0 1 2392
box -34 -1 6461 3249
use JK_FF_mag  JK_FF_mag_0
timestamp 1695127730
transform 1 0 464 0 1 205
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_2
timestamp 1695127730
transform 1 0 3690 0 1 139
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_3
timestamp 1695127730
transform 1 0 6783 0 1 139
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_4
timestamp 1695127730
transform -1 0 5766 0 -1 6707
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_5
timestamp 1695127730
transform -1 0 2655 0 -1 4501
box -390 0 2603 2148
<< labels >>
flabel metal1 6545 5099 6545 5099 0 FreeSans 640 0 0 0 CLK
port 0 nsew
flabel metal1 3295 4568 3295 4568 0 FreeSans 640 0 0 0 VDD
port 2 nsew
flabel metal1 3335 190 3335 190 0 FreeSans 640 0 0 0 VSS
port 3 nsew
flabel metal1 9093 4945 9093 4945 0 FreeSans 640 0 0 0 Vdiv96
port 4 nsew
flabel via2 2360 6164 2360 6164 0 FreeSans 960 0 0 0 RST
port 5 nsew
<< end >>
