magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2000 -2000 9344 2160
<< polysilicon >>
rect 0 103 102 160
rect 0 57 13 103
rect 59 57 102 103
rect 0 0 102 57
rect 7242 103 7344 160
rect 7242 57 7285 103
rect 7331 57 7344 103
rect 7242 0 7344 57
<< polycontact >>
rect 13 57 59 103
rect 7285 57 7331 103
<< ppolyres >>
rect 102 0 7242 160
<< metal1 >>
rect 2 103 70 158
rect 2 57 13 103
rect 59 57 70 103
rect 2 2 70 57
rect 7274 103 7342 158
rect 7274 57 7285 103
rect 7331 57 7342 103
rect 7274 2 7342 57
<< labels >>
rlabel polycontact 7308 80 7308 80 4 MINUS
rlabel polycontact 36 80 36 80 4 PLUS
<< end >>
