magic
tech gf180mcuC
magscale 1 10
timestamp 1694711135
<< nwell >>
rect -89 5603 10119 5761
rect -89 4643 111 5603
rect -89 4642 165 4643
rect -89 4636 168 4642
rect 9919 4637 10119 5603
rect 9897 4636 10119 4637
rect -89 4570 111 4636
rect 9667 4570 10119 4636
rect -89 4564 167 4570
rect -89 4563 165 4564
rect -89 4256 111 4563
rect 9919 4372 10119 4570
rect -89 4196 581 4256
rect 9720 4247 10119 4372
rect -89 4195 580 4196
rect -89 4145 291 4195
rect 350 4194 580 4195
rect 350 4145 581 4194
rect -89 4027 581 4145
rect -89 3527 111 4027
rect 9919 3991 10119 4247
rect 9887 3990 10119 3991
rect 9907 3924 10119 3990
rect 9919 3617 10119 3924
rect 9891 3550 10119 3617
rect 9919 3527 10119 3550
rect -89 3321 10119 3527
<< nsubdiff >>
rect -39 5698 10069 5715
rect -39 5648 -22 5698
rect 24 5652 76 5698
rect 122 5652 174 5698
rect 220 5652 272 5698
rect 318 5652 370 5698
rect 416 5652 468 5698
rect 514 5652 566 5698
rect 612 5652 664 5698
rect 710 5652 762 5698
rect 808 5652 860 5698
rect 906 5652 958 5698
rect 1004 5652 1056 5698
rect 1102 5652 1154 5698
rect 1200 5652 1252 5698
rect 1298 5652 1350 5698
rect 1396 5652 1448 5698
rect 1494 5652 1546 5698
rect 1592 5652 1644 5698
rect 1690 5652 1742 5698
rect 1788 5652 1840 5698
rect 1886 5652 1938 5698
rect 1984 5652 2036 5698
rect 2082 5652 2134 5698
rect 2180 5652 2232 5698
rect 2278 5652 2330 5698
rect 2376 5652 2428 5698
rect 2474 5652 2526 5698
rect 2572 5652 2624 5698
rect 2670 5652 2722 5698
rect 2768 5652 2820 5698
rect 2866 5652 2918 5698
rect 2964 5652 3016 5698
rect 3062 5652 3114 5698
rect 3160 5652 3212 5698
rect 3258 5652 3310 5698
rect 3356 5652 3408 5698
rect 3454 5652 3506 5698
rect 3552 5652 3604 5698
rect 3650 5652 3702 5698
rect 3748 5652 3800 5698
rect 3846 5652 3898 5698
rect 3944 5652 3996 5698
rect 4042 5652 4094 5698
rect 4140 5652 4192 5698
rect 4238 5652 4290 5698
rect 4336 5652 4388 5698
rect 4434 5652 4486 5698
rect 4532 5652 4584 5698
rect 4630 5652 4682 5698
rect 4728 5652 4780 5698
rect 4826 5652 4878 5698
rect 4924 5652 4976 5698
rect 5022 5652 5074 5698
rect 5120 5652 5172 5698
rect 5218 5652 5270 5698
rect 5316 5652 5368 5698
rect 5414 5652 5466 5698
rect 5512 5652 5564 5698
rect 5610 5652 5662 5698
rect 5708 5652 5760 5698
rect 5806 5652 5858 5698
rect 5904 5652 5956 5698
rect 6002 5652 6054 5698
rect 6100 5652 6152 5698
rect 6198 5652 6250 5698
rect 6296 5652 6348 5698
rect 6394 5652 6446 5698
rect 6492 5652 6544 5698
rect 6590 5652 6642 5698
rect 6688 5652 6740 5698
rect 6786 5652 6838 5698
rect 6884 5652 6936 5698
rect 6982 5652 7034 5698
rect 7080 5652 7132 5698
rect 7178 5652 7230 5698
rect 7276 5652 7328 5698
rect 7374 5652 7426 5698
rect 7472 5652 7524 5698
rect 7570 5652 7622 5698
rect 7668 5652 7720 5698
rect 7766 5652 7818 5698
rect 7864 5652 7916 5698
rect 7962 5652 8014 5698
rect 8060 5652 8112 5698
rect 8158 5652 8210 5698
rect 8256 5652 8308 5698
rect 8354 5652 8406 5698
rect 8452 5652 8504 5698
rect 8550 5652 8602 5698
rect 8648 5652 8700 5698
rect 8746 5652 8798 5698
rect 8844 5652 8896 5698
rect 8942 5652 8994 5698
rect 9040 5652 9092 5698
rect 9138 5652 9190 5698
rect 9236 5652 9288 5698
rect 9334 5652 9386 5698
rect 9432 5652 9484 5698
rect 9530 5652 9582 5698
rect 9628 5652 9680 5698
rect 9726 5652 9778 5698
rect 9824 5652 9876 5698
rect 9922 5652 10006 5698
rect 24 5648 10006 5652
rect 10052 5648 10069 5698
rect -39 5635 10069 5648
rect -39 5596 41 5635
rect -39 5550 -22 5596
rect 24 5550 41 5596
rect -39 5498 41 5550
rect -39 5452 -22 5498
rect 24 5452 41 5498
rect -39 5400 41 5452
rect -39 5354 -22 5400
rect 24 5354 41 5400
rect -39 5302 41 5354
rect -39 5256 -22 5302
rect 24 5256 41 5302
rect -39 5204 41 5256
rect -39 5158 -22 5204
rect 24 5158 41 5204
rect -39 5106 41 5158
rect -39 5060 -22 5106
rect 24 5060 41 5106
rect -39 5008 41 5060
rect -39 4962 -22 5008
rect 24 4962 41 5008
rect -39 4910 41 4962
rect -39 4864 -22 4910
rect 24 4864 41 4910
rect -39 4812 41 4864
rect -39 4766 -22 4812
rect 24 4766 41 4812
rect -39 4714 41 4766
rect -39 4668 -22 4714
rect 24 4668 41 4714
rect 9989 5596 10069 5635
rect 9989 5550 10006 5596
rect 10052 5550 10069 5596
rect 9989 5498 10069 5550
rect 9989 5452 10006 5498
rect 10052 5452 10069 5498
rect 9989 5400 10069 5452
rect 9989 5354 10006 5400
rect 10052 5354 10069 5400
rect 9989 5302 10069 5354
rect 9989 5256 10006 5302
rect 10052 5256 10069 5302
rect 9989 5204 10069 5256
rect 9989 5158 10006 5204
rect 10052 5158 10069 5204
rect 9989 5106 10069 5158
rect 9989 5060 10006 5106
rect 10052 5060 10069 5106
rect 9989 5008 10069 5060
rect 9989 4962 10006 5008
rect 10052 4962 10069 5008
rect 9989 4910 10069 4962
rect 9989 4864 10006 4910
rect 10052 4864 10069 4910
rect 9989 4812 10069 4864
rect 9989 4766 10006 4812
rect 10052 4766 10069 4812
rect 9989 4714 10069 4766
rect -39 4616 41 4668
rect 9989 4668 10006 4714
rect 10052 4668 10069 4714
rect -39 4570 -22 4616
rect 24 4570 41 4616
rect -39 4518 41 4570
rect -39 4472 -22 4518
rect 24 4472 41 4518
rect -39 4420 41 4472
rect -39 4374 -22 4420
rect 24 4374 41 4420
rect -39 4322 41 4374
rect -39 4276 -22 4322
rect 24 4276 41 4322
rect -39 4224 41 4276
rect -39 4178 -22 4224
rect 24 4178 41 4224
rect -39 4126 41 4178
rect -39 4080 -22 4126
rect 24 4080 41 4126
rect -39 4028 41 4080
rect -39 3982 -22 4028
rect 24 3982 41 4028
rect -39 3930 41 3982
rect -39 3884 -22 3930
rect 24 3884 41 3930
rect -39 3832 41 3884
rect -39 3786 -22 3832
rect 24 3786 41 3832
rect -39 3734 41 3786
rect -39 3688 -22 3734
rect 24 3688 41 3734
rect -39 3636 41 3688
rect -39 3590 -22 3636
rect 24 3590 41 3636
rect -39 3538 41 3590
rect -39 3492 -22 3538
rect 24 3492 41 3538
rect -39 3457 41 3492
rect 9989 4616 10069 4668
rect 9989 4570 10006 4616
rect 10052 4570 10069 4616
rect 9989 4518 10069 4570
rect 9989 4472 10006 4518
rect 10052 4472 10069 4518
rect 9989 4420 10069 4472
rect 9989 4374 10006 4420
rect 10052 4374 10069 4420
rect 9989 4322 10069 4374
rect 9989 4276 10006 4322
rect 10052 4276 10069 4322
rect 9989 4224 10069 4276
rect 9989 4178 10006 4224
rect 10052 4178 10069 4224
rect 9989 4126 10069 4178
rect 9989 4080 10006 4126
rect 10052 4080 10069 4126
rect 9989 4028 10069 4080
rect 9989 3982 10006 4028
rect 10052 3982 10069 4028
rect 9989 3930 10069 3982
rect 9989 3884 10006 3930
rect 10052 3884 10069 3930
rect 9989 3832 10069 3884
rect 9989 3786 10006 3832
rect 10052 3786 10069 3832
rect 9989 3734 10069 3786
rect 9989 3688 10006 3734
rect 10052 3688 10069 3734
rect 9989 3636 10069 3688
rect 9989 3590 10006 3636
rect 10052 3590 10069 3636
rect 9989 3538 10069 3590
rect 9989 3492 10006 3538
rect 10052 3492 10069 3538
rect 9989 3457 10069 3492
rect -39 3440 10069 3457
rect -39 3394 -22 3440
rect 24 3394 76 3440
rect 122 3394 174 3440
rect 220 3394 272 3440
rect 318 3394 370 3440
rect 416 3394 468 3440
rect 514 3394 566 3440
rect 612 3394 664 3440
rect 710 3394 762 3440
rect 808 3394 860 3440
rect 906 3394 958 3440
rect 1004 3394 1056 3440
rect 1102 3394 1154 3440
rect 1200 3394 1252 3440
rect 1298 3394 1350 3440
rect 1396 3394 1448 3440
rect 1494 3394 1546 3440
rect 1592 3394 1644 3440
rect 1690 3394 1742 3440
rect 1788 3394 1840 3440
rect 1886 3394 1938 3440
rect 1984 3394 2036 3440
rect 2082 3394 2134 3440
rect 2180 3394 2232 3440
rect 2278 3394 2330 3440
rect 2376 3394 2428 3440
rect 2474 3394 2526 3440
rect 2572 3394 2624 3440
rect 2670 3394 2722 3440
rect 2768 3394 2820 3440
rect 2866 3394 2918 3440
rect 2964 3394 3016 3440
rect 3062 3394 3114 3440
rect 3160 3394 3212 3440
rect 3258 3394 3310 3440
rect 3356 3394 3408 3440
rect 3454 3394 3506 3440
rect 3552 3394 3604 3440
rect 3650 3394 3702 3440
rect 3748 3394 3800 3440
rect 3846 3394 3898 3440
rect 3944 3394 3996 3440
rect 4042 3394 4094 3440
rect 4140 3394 4192 3440
rect 4238 3394 4290 3440
rect 4336 3394 4388 3440
rect 4434 3394 4486 3440
rect 4532 3394 4584 3440
rect 4630 3394 4682 3440
rect 4728 3394 4780 3440
rect 4826 3394 4878 3440
rect 4924 3394 4976 3440
rect 5022 3394 5074 3440
rect 5120 3394 5172 3440
rect 5218 3394 5270 3440
rect 5316 3394 5368 3440
rect 5414 3394 5466 3440
rect 5512 3394 5564 3440
rect 5610 3394 5662 3440
rect 5708 3394 5760 3440
rect 5806 3394 5858 3440
rect 5904 3394 5956 3440
rect 6002 3394 6054 3440
rect 6100 3394 6152 3440
rect 6198 3394 6250 3440
rect 6296 3394 6348 3440
rect 6394 3394 6446 3440
rect 6492 3394 6544 3440
rect 6590 3394 6642 3440
rect 6688 3394 6740 3440
rect 6786 3394 6838 3440
rect 6884 3394 6936 3440
rect 6982 3394 7034 3440
rect 7080 3394 7132 3440
rect 7178 3394 7230 3440
rect 7276 3394 7328 3440
rect 7374 3394 7426 3440
rect 7472 3394 7524 3440
rect 7570 3394 7622 3440
rect 7668 3394 7720 3440
rect 7766 3394 7818 3440
rect 7864 3394 7916 3440
rect 7962 3394 8014 3440
rect 8060 3394 8112 3440
rect 8158 3394 8210 3440
rect 8256 3394 8308 3440
rect 8354 3394 8406 3440
rect 8452 3394 8504 3440
rect 8550 3394 8602 3440
rect 8648 3394 8700 3440
rect 8746 3394 8798 3440
rect 8844 3394 8896 3440
rect 8942 3394 8994 3440
rect 9040 3394 9092 3440
rect 9138 3394 9190 3440
rect 9236 3394 9288 3440
rect 9334 3394 9386 3440
rect 9432 3394 9484 3440
rect 9530 3394 9582 3440
rect 9628 3394 9680 3440
rect 9726 3394 9778 3440
rect 9824 3394 9876 3440
rect 9922 3394 10006 3440
rect 10052 3394 10069 3440
rect -39 3377 10069 3394
<< nsubdiffcont >>
rect -22 5648 24 5698
rect 76 5652 122 5698
rect 174 5652 220 5698
rect 272 5652 318 5698
rect 370 5652 416 5698
rect 468 5652 514 5698
rect 566 5652 612 5698
rect 664 5652 710 5698
rect 762 5652 808 5698
rect 860 5652 906 5698
rect 958 5652 1004 5698
rect 1056 5652 1102 5698
rect 1154 5652 1200 5698
rect 1252 5652 1298 5698
rect 1350 5652 1396 5698
rect 1448 5652 1494 5698
rect 1546 5652 1592 5698
rect 1644 5652 1690 5698
rect 1742 5652 1788 5698
rect 1840 5652 1886 5698
rect 1938 5652 1984 5698
rect 2036 5652 2082 5698
rect 2134 5652 2180 5698
rect 2232 5652 2278 5698
rect 2330 5652 2376 5698
rect 2428 5652 2474 5698
rect 2526 5652 2572 5698
rect 2624 5652 2670 5698
rect 2722 5652 2768 5698
rect 2820 5652 2866 5698
rect 2918 5652 2964 5698
rect 3016 5652 3062 5698
rect 3114 5652 3160 5698
rect 3212 5652 3258 5698
rect 3310 5652 3356 5698
rect 3408 5652 3454 5698
rect 3506 5652 3552 5698
rect 3604 5652 3650 5698
rect 3702 5652 3748 5698
rect 3800 5652 3846 5698
rect 3898 5652 3944 5698
rect 3996 5652 4042 5698
rect 4094 5652 4140 5698
rect 4192 5652 4238 5698
rect 4290 5652 4336 5698
rect 4388 5652 4434 5698
rect 4486 5652 4532 5698
rect 4584 5652 4630 5698
rect 4682 5652 4728 5698
rect 4780 5652 4826 5698
rect 4878 5652 4924 5698
rect 4976 5652 5022 5698
rect 5074 5652 5120 5698
rect 5172 5652 5218 5698
rect 5270 5652 5316 5698
rect 5368 5652 5414 5698
rect 5466 5652 5512 5698
rect 5564 5652 5610 5698
rect 5662 5652 5708 5698
rect 5760 5652 5806 5698
rect 5858 5652 5904 5698
rect 5956 5652 6002 5698
rect 6054 5652 6100 5698
rect 6152 5652 6198 5698
rect 6250 5652 6296 5698
rect 6348 5652 6394 5698
rect 6446 5652 6492 5698
rect 6544 5652 6590 5698
rect 6642 5652 6688 5698
rect 6740 5652 6786 5698
rect 6838 5652 6884 5698
rect 6936 5652 6982 5698
rect 7034 5652 7080 5698
rect 7132 5652 7178 5698
rect 7230 5652 7276 5698
rect 7328 5652 7374 5698
rect 7426 5652 7472 5698
rect 7524 5652 7570 5698
rect 7622 5652 7668 5698
rect 7720 5652 7766 5698
rect 7818 5652 7864 5698
rect 7916 5652 7962 5698
rect 8014 5652 8060 5698
rect 8112 5652 8158 5698
rect 8210 5652 8256 5698
rect 8308 5652 8354 5698
rect 8406 5652 8452 5698
rect 8504 5652 8550 5698
rect 8602 5652 8648 5698
rect 8700 5652 8746 5698
rect 8798 5652 8844 5698
rect 8896 5652 8942 5698
rect 8994 5652 9040 5698
rect 9092 5652 9138 5698
rect 9190 5652 9236 5698
rect 9288 5652 9334 5698
rect 9386 5652 9432 5698
rect 9484 5652 9530 5698
rect 9582 5652 9628 5698
rect 9680 5652 9726 5698
rect 9778 5652 9824 5698
rect 9876 5652 9922 5698
rect 10006 5648 10052 5698
rect -22 5550 24 5596
rect -22 5452 24 5498
rect -22 5354 24 5400
rect -22 5256 24 5302
rect -22 5158 24 5204
rect -22 5060 24 5106
rect -22 4962 24 5008
rect -22 4864 24 4910
rect -22 4766 24 4812
rect -22 4668 24 4714
rect 10006 5550 10052 5596
rect 10006 5452 10052 5498
rect 10006 5354 10052 5400
rect 10006 5256 10052 5302
rect 10006 5158 10052 5204
rect 10006 5060 10052 5106
rect 10006 4962 10052 5008
rect 10006 4864 10052 4910
rect 10006 4766 10052 4812
rect 10006 4668 10052 4714
rect -22 4570 24 4616
rect -22 4472 24 4518
rect -22 4374 24 4420
rect -22 4276 24 4322
rect -22 4178 24 4224
rect -22 4080 24 4126
rect -22 3982 24 4028
rect -22 3884 24 3930
rect -22 3786 24 3832
rect -22 3688 24 3734
rect -22 3590 24 3636
rect -22 3492 24 3538
rect 10006 4570 10052 4616
rect 10006 4472 10052 4518
rect 10006 4374 10052 4420
rect 10006 4276 10052 4322
rect 10006 4178 10052 4224
rect 10006 4080 10052 4126
rect 10006 3982 10052 4028
rect 10006 3884 10052 3930
rect 10006 3786 10052 3832
rect 10006 3688 10052 3734
rect 10006 3590 10052 3636
rect 10006 3492 10052 3538
rect -22 3394 24 3440
rect 76 3394 122 3440
rect 174 3394 220 3440
rect 272 3394 318 3440
rect 370 3394 416 3440
rect 468 3394 514 3440
rect 566 3394 612 3440
rect 664 3394 710 3440
rect 762 3394 808 3440
rect 860 3394 906 3440
rect 958 3394 1004 3440
rect 1056 3394 1102 3440
rect 1154 3394 1200 3440
rect 1252 3394 1298 3440
rect 1350 3394 1396 3440
rect 1448 3394 1494 3440
rect 1546 3394 1592 3440
rect 1644 3394 1690 3440
rect 1742 3394 1788 3440
rect 1840 3394 1886 3440
rect 1938 3394 1984 3440
rect 2036 3394 2082 3440
rect 2134 3394 2180 3440
rect 2232 3394 2278 3440
rect 2330 3394 2376 3440
rect 2428 3394 2474 3440
rect 2526 3394 2572 3440
rect 2624 3394 2670 3440
rect 2722 3394 2768 3440
rect 2820 3394 2866 3440
rect 2918 3394 2964 3440
rect 3016 3394 3062 3440
rect 3114 3394 3160 3440
rect 3212 3394 3258 3440
rect 3310 3394 3356 3440
rect 3408 3394 3454 3440
rect 3506 3394 3552 3440
rect 3604 3394 3650 3440
rect 3702 3394 3748 3440
rect 3800 3394 3846 3440
rect 3898 3394 3944 3440
rect 3996 3394 4042 3440
rect 4094 3394 4140 3440
rect 4192 3394 4238 3440
rect 4290 3394 4336 3440
rect 4388 3394 4434 3440
rect 4486 3394 4532 3440
rect 4584 3394 4630 3440
rect 4682 3394 4728 3440
rect 4780 3394 4826 3440
rect 4878 3394 4924 3440
rect 4976 3394 5022 3440
rect 5074 3394 5120 3440
rect 5172 3394 5218 3440
rect 5270 3394 5316 3440
rect 5368 3394 5414 3440
rect 5466 3394 5512 3440
rect 5564 3394 5610 3440
rect 5662 3394 5708 3440
rect 5760 3394 5806 3440
rect 5858 3394 5904 3440
rect 5956 3394 6002 3440
rect 6054 3394 6100 3440
rect 6152 3394 6198 3440
rect 6250 3394 6296 3440
rect 6348 3394 6394 3440
rect 6446 3394 6492 3440
rect 6544 3394 6590 3440
rect 6642 3394 6688 3440
rect 6740 3394 6786 3440
rect 6838 3394 6884 3440
rect 6936 3394 6982 3440
rect 7034 3394 7080 3440
rect 7132 3394 7178 3440
rect 7230 3394 7276 3440
rect 7328 3394 7374 3440
rect 7426 3394 7472 3440
rect 7524 3394 7570 3440
rect 7622 3394 7668 3440
rect 7720 3394 7766 3440
rect 7818 3394 7864 3440
rect 7916 3394 7962 3440
rect 8014 3394 8060 3440
rect 8112 3394 8158 3440
rect 8210 3394 8256 3440
rect 8308 3394 8354 3440
rect 8406 3394 8452 3440
rect 8504 3394 8550 3440
rect 8602 3394 8648 3440
rect 8700 3394 8746 3440
rect 8798 3394 8844 3440
rect 8896 3394 8942 3440
rect 8994 3394 9040 3440
rect 9092 3394 9138 3440
rect 9190 3394 9236 3440
rect 9288 3394 9334 3440
rect 9386 3394 9432 3440
rect 9484 3394 9530 3440
rect 9582 3394 9628 3440
rect 9680 3394 9726 3440
rect 9778 3394 9824 3440
rect 9876 3394 9922 3440
rect 10006 3394 10052 3440
<< polysilicon >>
rect 5435 4665 5524 4708
<< metal1 >>
rect -39 5698 10069 5715
rect -39 5648 -22 5698
rect 24 5652 76 5698
rect 122 5652 174 5698
rect 220 5652 272 5698
rect 318 5652 370 5698
rect 416 5652 468 5698
rect 514 5652 566 5698
rect 612 5652 664 5698
rect 710 5652 762 5698
rect 808 5652 860 5698
rect 906 5652 958 5698
rect 1004 5652 1056 5698
rect 1102 5652 1154 5698
rect 1200 5652 1252 5698
rect 1298 5652 1350 5698
rect 1396 5652 1448 5698
rect 1494 5652 1546 5698
rect 1592 5652 1644 5698
rect 1690 5652 1742 5698
rect 1788 5652 1840 5698
rect 1886 5652 1938 5698
rect 1984 5652 2036 5698
rect 2082 5652 2134 5698
rect 2180 5652 2232 5698
rect 2278 5652 2330 5698
rect 2376 5652 2428 5698
rect 2474 5652 2526 5698
rect 2572 5652 2624 5698
rect 2670 5652 2722 5698
rect 2768 5652 2820 5698
rect 2866 5652 2918 5698
rect 2964 5652 3016 5698
rect 3062 5652 3114 5698
rect 3160 5652 3212 5698
rect 3258 5652 3310 5698
rect 3356 5652 3408 5698
rect 3454 5652 3506 5698
rect 3552 5652 3604 5698
rect 3650 5652 3702 5698
rect 3748 5652 3800 5698
rect 3846 5652 3898 5698
rect 3944 5652 3996 5698
rect 4042 5652 4094 5698
rect 4140 5652 4192 5698
rect 4238 5652 4290 5698
rect 4336 5652 4388 5698
rect 4434 5652 4486 5698
rect 4532 5652 4584 5698
rect 4630 5652 4682 5698
rect 4728 5652 4780 5698
rect 4826 5652 4878 5698
rect 4924 5652 4976 5698
rect 5022 5652 5074 5698
rect 5120 5652 5172 5698
rect 5218 5652 5270 5698
rect 5316 5652 5368 5698
rect 5414 5652 5466 5698
rect 5512 5652 5564 5698
rect 5610 5652 5662 5698
rect 5708 5652 5760 5698
rect 5806 5652 5858 5698
rect 5904 5652 5956 5698
rect 6002 5652 6054 5698
rect 6100 5652 6152 5698
rect 6198 5652 6250 5698
rect 6296 5652 6348 5698
rect 6394 5652 6446 5698
rect 6492 5652 6544 5698
rect 6590 5652 6642 5698
rect 6688 5652 6740 5698
rect 6786 5652 6838 5698
rect 6884 5652 6936 5698
rect 6982 5652 7034 5698
rect 7080 5652 7132 5698
rect 7178 5652 7230 5698
rect 7276 5652 7328 5698
rect 7374 5652 7426 5698
rect 7472 5652 7524 5698
rect 7570 5652 7622 5698
rect 7668 5652 7720 5698
rect 7766 5652 7818 5698
rect 7864 5652 7916 5698
rect 7962 5652 8014 5698
rect 8060 5652 8112 5698
rect 8158 5652 8210 5698
rect 8256 5652 8308 5698
rect 8354 5652 8406 5698
rect 8452 5652 8504 5698
rect 8550 5652 8602 5698
rect 8648 5652 8700 5698
rect 8746 5652 8798 5698
rect 8844 5652 8896 5698
rect 8942 5652 8994 5698
rect 9040 5652 9092 5698
rect 9138 5652 9190 5698
rect 9236 5652 9288 5698
rect 9334 5652 9386 5698
rect 9432 5652 9484 5698
rect 9530 5652 9582 5698
rect 9628 5652 9680 5698
rect 9726 5652 9778 5698
rect 9824 5652 9876 5698
rect 9922 5652 10006 5698
rect 24 5648 10006 5652
rect 10052 5648 10069 5698
rect -39 5635 10069 5648
rect -39 5596 41 5635
rect -39 5550 -22 5596
rect 24 5550 41 5596
rect -39 5498 41 5550
rect -39 5452 -22 5498
rect 24 5452 41 5498
rect -39 5400 41 5452
rect -39 5354 -22 5400
rect 24 5354 41 5400
rect -39 5302 41 5354
rect -39 5256 -22 5302
rect 24 5256 41 5302
rect -39 5204 41 5256
rect -39 5158 -22 5204
rect 24 5158 41 5204
rect -39 5106 41 5158
rect -39 5060 -22 5106
rect 24 5060 41 5106
rect -39 5008 41 5060
rect 369 5030 438 5635
rect 9989 5596 10069 5635
rect 9989 5550 10006 5596
rect 10052 5550 10069 5596
rect 2454 5512 2644 5516
rect 2454 5503 2466 5512
rect 1556 5457 2466 5503
rect 1556 5406 1602 5457
rect 2454 5456 2466 5457
rect 2522 5456 2576 5512
rect 2632 5456 2644 5512
rect 2454 5452 2644 5456
rect 2906 5512 3096 5516
rect 2906 5456 2918 5512
rect 2974 5456 3028 5512
rect 3084 5503 3096 5512
rect 6934 5512 7124 5516
rect 6934 5503 6946 5512
rect 3084 5457 3994 5503
rect 3084 5456 3096 5457
rect 2906 5452 3096 5456
rect 577 5360 1064 5406
rect 1137 5360 1148 5406
rect 588 5074 669 5360
rect 1192 5208 1249 5406
rect 1322 5360 1333 5406
rect 1417 5360 1428 5406
rect 1556 5360 1613 5406
rect 1695 5401 1895 5410
rect 1695 5345 1709 5401
rect 1765 5345 1819 5401
rect 1875 5345 1895 5401
rect 1977 5360 1988 5406
rect 1695 5333 1895 5345
rect 2052 5304 2102 5408
rect 2162 5360 2173 5406
rect 2257 5360 2733 5406
rect 2817 5360 3293 5406
rect 3377 5360 3388 5406
rect 3448 5304 3498 5408
rect 3562 5360 3573 5406
rect 3655 5401 3855 5410
rect 3948 5406 3994 5457
rect 6036 5457 6946 5503
rect 6036 5406 6082 5457
rect 6934 5456 6946 5457
rect 7002 5456 7056 5512
rect 7112 5456 7124 5512
rect 6934 5452 7124 5456
rect 7386 5512 7576 5516
rect 7386 5456 7398 5512
rect 7454 5456 7508 5512
rect 7564 5503 7576 5512
rect 7564 5457 8474 5503
rect 7564 5456 7576 5457
rect 7386 5452 7576 5456
rect 3655 5345 3675 5401
rect 3731 5345 3785 5401
rect 3841 5345 3855 5401
rect 3937 5360 3994 5406
rect 4122 5360 4133 5406
rect 4217 5360 4228 5406
rect 3655 5333 3855 5345
rect 2052 5254 3498 5304
rect 4301 5208 4358 5406
rect 4402 5360 4413 5406
rect 4486 5360 4973 5406
rect 5057 5360 5544 5406
rect 5617 5360 5628 5406
rect 1192 5151 4358 5208
rect 5672 5208 5729 5406
rect 5802 5360 5813 5406
rect 5897 5360 5908 5406
rect 6036 5360 6093 5406
rect 6175 5401 6375 5410
rect 6175 5345 6189 5401
rect 6245 5345 6299 5401
rect 6355 5345 6375 5401
rect 6457 5360 6468 5406
rect 6175 5333 6375 5345
rect 6532 5304 6582 5408
rect 6642 5360 6653 5406
rect 6737 5360 7213 5406
rect 7297 5360 7773 5406
rect 7857 5360 7868 5406
rect 7928 5304 7978 5408
rect 8042 5360 8053 5406
rect 8135 5401 8335 5410
rect 8428 5406 8474 5457
rect 9989 5498 10069 5550
rect 9989 5452 10006 5498
rect 10052 5452 10069 5498
rect 9989 5412 10069 5452
rect 8135 5345 8155 5401
rect 8211 5345 8265 5401
rect 8321 5345 8335 5401
rect 8417 5360 8474 5406
rect 8602 5360 8613 5406
rect 8697 5360 8708 5406
rect 8135 5333 8335 5345
rect 6532 5254 7978 5304
rect 8781 5208 8838 5406
rect 8882 5360 8893 5406
rect 8966 5360 9453 5406
rect 9537 5360 9548 5406
rect 9720 5400 10069 5412
rect 9720 5355 10006 5400
rect 5672 5151 8838 5208
rect 9989 5354 10006 5355
rect 10052 5354 10069 5400
rect 9989 5302 10069 5354
rect 9989 5256 10006 5302
rect 10052 5256 10069 5302
rect 9989 5204 10069 5256
rect 9989 5158 10006 5204
rect 10052 5158 10069 5204
rect 9989 5106 10069 5158
rect 577 5038 669 5074
rect 855 5086 1055 5100
rect 577 5028 634 5038
rect -39 4962 -22 5008
rect 24 4962 41 5008
rect -39 4910 41 4962
rect -39 4864 -22 4910
rect 24 4864 41 4910
rect 333 4967 530 4972
rect 333 4911 349 4967
rect 405 4911 459 4967
rect 515 4962 530 4967
rect 588 4962 634 5028
rect 855 5030 867 5086
rect 923 5030 975 5086
rect 1031 5030 1055 5086
rect 1415 5093 1615 5101
rect 855 5023 1055 5030
rect 1137 5028 1148 5074
rect 515 4916 634 4962
rect 515 4911 530 4916
rect 333 4906 530 4911
rect -39 4812 41 4864
rect -236 4752 -170 4767
rect -236 4696 -231 4752
rect -175 4696 -170 4752
rect -236 4642 -170 4696
rect -236 4586 -231 4642
rect -175 4586 -170 4642
rect -236 4570 -170 4586
rect -39 4766 -22 4812
rect 24 4766 41 4812
rect -39 4763 41 4766
rect 714 4900 1029 4904
rect 714 4844 851 4900
rect 907 4844 961 4900
rect 1017 4844 1029 4900
rect 714 4838 1029 4844
rect 1155 4857 1201 5073
rect 1322 5028 1333 5074
rect 1415 5037 1428 5093
rect 1484 5037 1538 5093
rect 1594 5037 1615 5093
rect 1415 5024 1615 5037
rect 1695 5090 1895 5101
rect 1695 5034 1709 5090
rect 1765 5034 1819 5090
rect 1875 5034 1895 5090
rect 2255 5087 2455 5101
rect 1695 5024 1895 5034
rect 1977 5028 2038 5074
rect 2162 5028 2173 5074
rect 2255 5031 2267 5087
rect 2323 5031 2377 5087
rect 2433 5031 2455 5087
rect 3095 5087 3295 5101
rect 1250 4966 1442 4968
rect 1988 4966 2038 5028
rect 2255 5024 2455 5031
rect 2537 5028 3013 5074
rect 3095 5031 3117 5087
rect 3173 5031 3227 5087
rect 3283 5031 3295 5087
rect 3655 5090 3855 5101
rect 3095 5024 3295 5031
rect 3377 5028 3388 5074
rect 3512 5028 3573 5074
rect 3655 5034 3675 5090
rect 3731 5034 3785 5090
rect 3841 5034 3855 5090
rect 1250 4965 2038 4966
rect 1250 4909 1262 4965
rect 1318 4909 1372 4965
rect 1428 4920 2038 4965
rect 3512 4966 3562 5028
rect 3655 5024 3855 5034
rect 3935 5093 4135 5101
rect 3935 5037 3956 5093
rect 4012 5037 4066 5093
rect 4122 5037 4135 5093
rect 4495 5086 4695 5100
rect 3935 5024 4135 5037
rect 4217 5028 4228 5074
rect 4108 4966 4300 4968
rect 3512 4965 4300 4966
rect 3512 4920 4122 4965
rect 1428 4909 1442 4920
rect 1250 4906 1442 4909
rect 4108 4909 4122 4920
rect 4178 4909 4232 4965
rect 4288 4909 4300 4965
rect 4108 4906 4300 4909
rect 4349 4857 4395 5073
rect 4402 5028 4413 5074
rect 4495 5030 4519 5086
rect 4575 5030 4627 5086
rect 4683 5030 4695 5086
rect 5335 5086 5535 5100
rect 4495 5023 4695 5030
rect 4916 5028 4973 5074
rect 5057 5028 5114 5074
rect 5242 5028 5253 5074
rect 5335 5030 5347 5086
rect 5403 5030 5455 5086
rect 5511 5030 5535 5086
rect 5895 5093 6095 5101
rect 4916 4982 4962 5028
rect 5068 4982 5114 5028
rect 5335 5023 5535 5030
rect 5617 5028 5628 5074
rect 4884 4936 5114 4982
rect -39 4714 348 4763
rect -39 4668 -22 4714
rect 24 4697 348 4714
rect 714 4708 762 4838
rect 1155 4811 2038 4857
rect 855 4744 1055 4756
rect 24 4668 41 4697
rect 855 4688 870 4744
rect 926 4688 980 4744
rect 1036 4688 1055 4744
rect 855 4678 1055 4688
rect 1135 4750 1335 4758
rect 1135 4694 1150 4750
rect 1206 4694 1260 4750
rect 1316 4694 1335 4750
rect 1417 4708 1428 4754
rect 1135 4681 1335 4694
rect -39 4616 41 4668
rect -39 4570 -22 4616
rect 24 4570 41 4616
rect 96 4632 293 4636
rect 1491 4632 1541 4755
rect 1602 4708 1613 4754
rect 1697 4708 1708 4754
rect 96 4631 1541 4632
rect 96 4575 109 4631
rect 165 4575 219 4631
rect 275 4582 1541 4631
rect 1775 4630 1825 4755
rect 1988 4754 2038 4811
rect 3512 4811 4395 4857
rect 4519 4899 4836 4904
rect 4519 4843 4531 4899
rect 4587 4843 4641 4899
rect 4697 4843 4836 4899
rect 4519 4838 4836 4843
rect 1882 4708 1893 4754
rect 1977 4708 2038 4754
rect 2162 4708 2173 4754
rect 2255 4743 2455 4757
rect 2255 4687 2269 4743
rect 2325 4687 2379 4743
rect 2435 4687 2455 4743
rect 2255 4677 2455 4687
rect 2535 4745 2735 4758
rect 2535 4689 2548 4745
rect 2604 4689 2658 4745
rect 2714 4689 2735 4745
rect 2535 4681 2735 4689
rect 2815 4745 3015 4758
rect 2815 4689 2836 4745
rect 2892 4689 2946 4745
rect 3002 4689 3015 4745
rect 2815 4681 3015 4689
rect 3095 4743 3295 4757
rect 3512 4754 3562 4811
rect 3095 4687 3115 4743
rect 3171 4687 3225 4743
rect 3281 4687 3295 4743
rect 3377 4708 3388 4754
rect 3512 4708 3573 4754
rect 3657 4708 3668 4754
rect 3095 4677 3295 4687
rect 3725 4630 3775 4755
rect 3842 4708 3853 4754
rect 3937 4708 3948 4754
rect 275 4575 293 4582
rect 1775 4580 3775 4630
rect 4009 4632 4059 4755
rect 4122 4708 4133 4754
rect 4215 4750 4415 4758
rect 4215 4694 4234 4750
rect 4290 4694 4344 4750
rect 4400 4694 4415 4750
rect 4215 4681 4415 4694
rect 4495 4744 4695 4756
rect 4788 4754 4836 4838
rect 5194 4900 5509 4904
rect 5194 4844 5331 4900
rect 5387 4844 5441 4900
rect 5497 4844 5509 4900
rect 5194 4838 5509 4844
rect 5635 4857 5681 5073
rect 5802 5028 5813 5074
rect 5895 5037 5908 5093
rect 5964 5037 6018 5093
rect 6074 5037 6095 5093
rect 5895 5024 6095 5037
rect 6175 5090 6375 5101
rect 6175 5034 6189 5090
rect 6245 5034 6299 5090
rect 6355 5034 6375 5090
rect 6735 5087 6935 5101
rect 6175 5024 6375 5034
rect 6457 5028 6518 5074
rect 6642 5028 6653 5074
rect 6735 5031 6747 5087
rect 6803 5031 6857 5087
rect 6913 5031 6935 5087
rect 7575 5087 7775 5101
rect 5730 4966 5922 4968
rect 6468 4966 6518 5028
rect 6735 5024 6935 5031
rect 7017 5028 7493 5074
rect 7575 5031 7597 5087
rect 7653 5031 7707 5087
rect 7763 5031 7775 5087
rect 8135 5090 8335 5101
rect 7575 5024 7775 5031
rect 7857 5028 7868 5074
rect 7992 5028 8053 5074
rect 8135 5034 8155 5090
rect 8211 5034 8265 5090
rect 8321 5034 8335 5090
rect 5730 4965 6518 4966
rect 5730 4909 5742 4965
rect 5798 4909 5852 4965
rect 5908 4920 6518 4965
rect 7992 4966 8042 5028
rect 8135 5024 8335 5034
rect 8415 5093 8615 5101
rect 8415 5037 8436 5093
rect 8492 5037 8546 5093
rect 8602 5037 8615 5093
rect 8975 5086 9175 5100
rect 9989 5086 10006 5106
rect 8415 5024 8615 5037
rect 8697 5028 8708 5074
rect 8588 4966 8780 4968
rect 7992 4965 8780 4966
rect 7992 4920 8602 4965
rect 5908 4909 5922 4920
rect 5730 4906 5922 4909
rect 8588 4909 8602 4920
rect 8658 4909 8712 4965
rect 8768 4909 8780 4965
rect 8588 4906 8780 4909
rect 8829 4857 8875 5073
rect 8882 5028 8893 5074
rect 8975 5030 8999 5086
rect 9055 5030 9107 5086
rect 9163 5030 9175 5086
rect 8975 5023 9175 5030
rect 9257 5028 9268 5074
rect 9396 5028 9453 5074
rect 9537 5028 9548 5074
rect 9720 5060 10006 5086
rect 10052 5060 10069 5106
rect 9720 5029 10069 5060
rect 9722 5028 9733 5029
rect 9396 4962 9442 5028
rect 9989 5008 10069 5029
rect 9700 4967 9897 4972
rect 9700 4962 9713 4967
rect 9396 4916 9713 4962
rect 9700 4911 9713 4916
rect 9771 4911 9823 4967
rect 9881 4911 9897 4967
rect 9700 4906 9897 4911
rect 9989 4962 10006 5008
rect 10052 4962 10069 5008
rect 9989 4910 10069 4962
rect 5194 4754 5242 4838
rect 5635 4811 6518 4857
rect 4495 4688 4514 4744
rect 4570 4688 4624 4744
rect 4680 4688 4695 4744
rect 4777 4708 4836 4754
rect 4962 4708 4973 4754
rect 5057 4708 5068 4754
rect 5194 4708 5253 4754
rect 5335 4744 5535 4756
rect 4495 4678 4695 4688
rect 5335 4688 5350 4744
rect 5406 4688 5460 4744
rect 5516 4688 5535 4744
rect 5335 4678 5535 4688
rect 5615 4750 5815 4758
rect 5615 4694 5630 4750
rect 5686 4694 5740 4750
rect 5796 4694 5815 4750
rect 5897 4708 5908 4754
rect 5615 4681 5815 4694
rect 5971 4632 6021 4755
rect 6082 4708 6093 4754
rect 6177 4708 6188 4754
rect 4009 4582 6021 4632
rect 6255 4630 6305 4755
rect 6468 4754 6518 4811
rect 7992 4811 8875 4857
rect 8999 4899 9316 4904
rect 8999 4843 9011 4899
rect 9067 4843 9121 4899
rect 9177 4843 9316 4899
rect 8999 4838 9316 4843
rect 6362 4708 6373 4754
rect 6457 4708 6518 4754
rect 6642 4708 6653 4754
rect 6735 4743 6935 4757
rect 6735 4687 6749 4743
rect 6805 4687 6859 4743
rect 6915 4687 6935 4743
rect 6735 4677 6935 4687
rect 7015 4745 7215 4758
rect 7015 4689 7028 4745
rect 7084 4689 7138 4745
rect 7194 4689 7215 4745
rect 7015 4681 7215 4689
rect 7295 4745 7495 4758
rect 7295 4689 7316 4745
rect 7372 4689 7426 4745
rect 7482 4689 7495 4745
rect 7295 4681 7495 4689
rect 7575 4743 7775 4757
rect 7992 4754 8042 4811
rect 7575 4687 7595 4743
rect 7651 4687 7705 4743
rect 7761 4687 7775 4743
rect 7857 4708 7868 4754
rect 7992 4708 8053 4754
rect 8137 4708 8148 4754
rect 7575 4677 7775 4687
rect 8205 4630 8255 4755
rect 8322 4708 8333 4754
rect 8417 4708 8428 4754
rect 6255 4580 8255 4630
rect 8489 4632 8539 4755
rect 8602 4708 8613 4754
rect 8695 4750 8895 4758
rect 8695 4694 8714 4750
rect 8770 4694 8824 4750
rect 8880 4694 8895 4750
rect 8695 4681 8895 4694
rect 8975 4744 9175 4756
rect 9268 4754 9316 4838
rect 9989 4864 10006 4910
rect 10052 4864 10069 4910
rect 9989 4812 10069 4864
rect 9989 4766 10006 4812
rect 10052 4766 10069 4812
rect 9989 4763 10069 4766
rect 8975 4688 8994 4744
rect 9050 4688 9104 4744
rect 9160 4688 9175 4744
rect 9257 4708 9316 4754
rect 9442 4708 9453 4754
rect 9537 4708 9548 4754
rect 9718 4714 10069 4763
rect 9718 4706 10006 4714
rect 8975 4678 9175 4688
rect 9989 4668 10006 4706
rect 10052 4668 10069 4714
rect 9485 4632 9682 4636
rect 8489 4631 9682 4632
rect 8489 4582 9503 4631
rect 96 4570 293 4575
rect -346 4447 -280 4462
rect -346 4391 -341 4447
rect -285 4391 -280 4447
rect -468 4325 -402 4340
rect -468 4269 -463 4325
rect -407 4269 -402 4325
rect -468 4215 -402 4269
rect -468 4159 -463 4215
rect -407 4159 -402 4215
rect -468 4153 -402 4159
rect -469 4143 -402 4153
rect -346 4337 -280 4391
rect -346 4281 -341 4337
rect -285 4281 -280 4337
rect -346 4265 -280 4281
rect -582 3733 -516 3748
rect -582 3677 -577 3733
rect -521 3677 -516 3733
rect -582 3623 -516 3677
rect -582 3567 -577 3623
rect -521 3567 -516 3623
rect -582 3553 -516 3567
rect -582 3551 -517 3553
rect -580 3321 -517 3551
rect -469 3321 -406 4143
rect -346 3321 -283 4265
rect -234 3321 -171 4570
rect -39 4518 41 4570
rect -39 4472 -22 4518
rect 24 4472 41 4518
rect -39 4443 41 4472
rect -39 4420 349 4443
rect 855 4438 1055 4448
rect -39 4374 -22 4420
rect 24 4377 349 4420
rect 24 4374 41 4377
rect 577 4376 634 4422
rect -39 4322 41 4374
rect -39 4276 -22 4322
rect 24 4276 41 4322
rect -39 4224 41 4276
rect 87 4326 284 4331
rect 87 4270 100 4326
rect 156 4270 210 4326
rect 266 4323 284 4326
rect 588 4323 634 4376
rect 855 4382 868 4438
rect 924 4382 978 4438
rect 1034 4382 1055 4438
rect 855 4371 1055 4382
rect 1135 4439 1335 4449
rect 1135 4383 1148 4439
rect 1204 4383 1258 4439
rect 1314 4383 1335 4439
rect 2255 4437 2455 4449
rect 1987 4422 2037 4423
rect 1135 4372 1335 4383
rect 1417 4376 1893 4422
rect 1977 4376 2037 4422
rect 2162 4376 2173 4422
rect 2255 4381 2270 4437
rect 2326 4381 2380 4437
rect 2436 4381 2455 4437
rect 266 4277 634 4323
rect 1987 4320 2037 4376
rect 2255 4371 2455 4381
rect 2537 4437 2734 4442
rect 2537 4381 2553 4437
rect 2609 4381 2663 4437
rect 2719 4422 2734 4437
rect 2817 4437 3014 4442
rect 2817 4422 2833 4437
rect 2719 4381 2833 4422
rect 2889 4381 2943 4437
rect 2999 4381 3014 4437
rect 2537 4376 3014 4381
rect 3095 4437 3295 4449
rect 3095 4381 3114 4437
rect 3170 4381 3224 4437
rect 3280 4381 3295 4437
rect 4215 4439 4415 4449
rect 3513 4422 3563 4423
rect 3095 4371 3295 4381
rect 3377 4376 3388 4422
rect 3513 4376 3573 4422
rect 3657 4376 4133 4422
rect 4215 4383 4236 4439
rect 4292 4383 4346 4439
rect 4402 4383 4415 4439
rect 266 4270 284 4277
rect 87 4265 284 4270
rect 1154 4274 2037 4320
rect 3513 4320 3563 4376
rect 4215 4372 4415 4383
rect 4495 4438 4695 4448
rect 4495 4382 4516 4438
rect 4572 4382 4626 4438
rect 4682 4382 4695 4438
rect 5335 4438 5535 4448
rect 4495 4371 4695 4382
rect 4916 4376 4973 4422
rect 5057 4376 5114 4422
rect 5242 4376 5253 4422
rect 5335 4382 5348 4438
rect 5404 4382 5458 4438
rect 5514 4382 5535 4438
rect 4916 4330 4962 4376
rect 5068 4330 5114 4376
rect 5335 4371 5535 4382
rect 5615 4439 5815 4449
rect 5615 4383 5628 4439
rect 5684 4383 5738 4439
rect 5794 4383 5815 4439
rect 6735 4437 6935 4449
rect 6467 4422 6517 4423
rect 5615 4372 5815 4383
rect 5897 4376 6373 4422
rect 6457 4376 6517 4422
rect 6642 4376 6653 4422
rect 6735 4381 6750 4437
rect 6806 4381 6860 4437
rect 6916 4381 6935 4437
rect 7575 4437 7775 4449
rect 3513 4274 4396 4320
rect 4884 4284 5114 4330
rect 6467 4320 6517 4376
rect 6735 4371 6935 4381
rect 7017 4376 7493 4422
rect 7575 4381 7594 4437
rect 7650 4381 7704 4437
rect 7760 4381 7775 4437
rect 8695 4439 8895 4449
rect 7993 4422 8043 4423
rect 7575 4371 7775 4381
rect 7857 4376 7868 4422
rect 7993 4376 8053 4422
rect 8137 4376 8613 4422
rect 8695 4383 8716 4439
rect 8772 4383 8826 4439
rect 8882 4383 8895 4439
rect -39 4178 -22 4224
rect 24 4178 41 4224
rect -39 4126 41 4178
rect 350 4209 547 4214
rect 350 4153 366 4209
rect 422 4153 476 4209
rect 532 4194 547 4209
rect 532 4153 634 4194
rect 350 4148 634 4153
rect -39 4080 -22 4126
rect 24 4103 41 4126
rect 24 4101 313 4103
rect 588 4102 634 4148
rect 24 4080 315 4101
rect -39 4058 315 4080
rect -39 4056 313 4058
rect 581 4056 634 4102
rect 855 4096 1055 4106
rect -39 4028 41 4056
rect 855 4040 868 4096
rect 924 4040 978 4096
rect 1034 4040 1055 4096
rect 1137 4056 1148 4102
rect 1154 4058 1200 4274
rect 1249 4210 1329 4215
rect 1249 4154 1261 4210
rect 1317 4204 1329 4210
rect 4221 4210 4301 4215
rect 4221 4204 4233 4210
rect 1317 4158 2038 4204
rect 1317 4154 1329 4158
rect 1249 4148 1329 4154
rect 1322 4056 1333 4102
rect 1415 4095 1615 4106
rect 855 4029 1055 4040
rect 1415 4039 1429 4095
rect 1485 4039 1539 4095
rect 1595 4039 1615 4095
rect 1415 4029 1615 4039
rect 1695 4096 1895 4106
rect 1988 4102 2038 4158
rect 3512 4158 4233 4204
rect 3512 4102 3562 4158
rect 4221 4154 4233 4158
rect 4289 4154 4301 4210
rect 4221 4148 4301 4154
rect 1695 4040 1710 4096
rect 1766 4040 1820 4096
rect 1876 4040 1895 4096
rect 1977 4056 2038 4102
rect 2162 4056 2173 4102
rect 2257 4056 2584 4102
rect 2680 4056 2733 4102
rect 2817 4056 2877 4102
rect 2973 4056 3293 4102
rect 3377 4056 3388 4102
rect 3512 4056 3573 4102
rect 3655 4096 3855 4106
rect 1695 4029 1895 4040
rect 3655 4040 3674 4096
rect 3730 4040 3784 4096
rect 3840 4040 3855 4096
rect 3655 4029 3855 4040
rect 3935 4095 4135 4106
rect 3935 4039 3955 4095
rect 4011 4039 4065 4095
rect 4121 4039 4135 4095
rect 4217 4056 4228 4102
rect 4350 4058 4396 4274
rect 5634 4274 6517 4320
rect 7993 4320 8043 4376
rect 8695 4372 8895 4383
rect 8975 4438 9175 4448
rect 8975 4382 8996 4438
rect 9052 4382 9106 4438
rect 9162 4382 9175 4438
rect 9268 4422 9326 4582
rect 9485 4575 9503 4582
rect 9559 4575 9613 4631
rect 9669 4575 9682 4631
rect 9485 4570 9682 4575
rect 9989 4616 10069 4668
rect 9989 4570 10006 4616
rect 10052 4570 10069 4616
rect 9989 4518 10069 4570
rect 9989 4472 10006 4518
rect 10052 4472 10069 4518
rect 9989 4425 10069 4472
rect 8975 4371 9175 4382
rect 9257 4376 9326 4422
rect 9537 4376 9548 4422
rect 9717 4420 10069 4425
rect 9717 4374 10006 4420
rect 10052 4374 10069 4420
rect 9717 4368 10069 4374
rect 9989 4322 10069 4368
rect 7993 4274 8876 4320
rect 4884 4148 5114 4194
rect 4402 4056 4413 4102
rect 4495 4096 4695 4106
rect 3935 4029 4135 4039
rect 4495 4040 4516 4096
rect 4572 4040 4626 4096
rect 4682 4040 4695 4096
rect 4916 4102 4962 4148
rect 5068 4102 5114 4148
rect 4916 4056 4973 4102
rect 5057 4056 5114 4102
rect 5242 4056 5253 4102
rect 5335 4096 5535 4106
rect 4495 4029 4695 4040
rect 5335 4040 5348 4096
rect 5404 4040 5458 4096
rect 5514 4040 5535 4096
rect 5617 4056 5628 4102
rect 5634 4058 5680 4274
rect 5729 4210 5809 4215
rect 5729 4154 5741 4210
rect 5797 4204 5809 4210
rect 8701 4210 8781 4215
rect 8701 4204 8713 4210
rect 5797 4158 6518 4204
rect 5797 4154 5809 4158
rect 5729 4148 5809 4154
rect 5802 4056 5813 4102
rect 5895 4095 6095 4106
rect 5335 4029 5535 4040
rect 5895 4039 5909 4095
rect 5965 4039 6019 4095
rect 6075 4039 6095 4095
rect 5895 4029 6095 4039
rect 6175 4096 6375 4106
rect 6468 4102 6518 4158
rect 7992 4158 8713 4204
rect 7992 4102 8042 4158
rect 8701 4154 8713 4158
rect 8769 4154 8781 4210
rect 8701 4148 8781 4154
rect 6175 4040 6190 4096
rect 6246 4040 6300 4096
rect 6356 4040 6375 4096
rect 6457 4056 6518 4102
rect 6642 4056 6653 4102
rect 6737 4056 7213 4102
rect 7297 4056 7773 4102
rect 7857 4056 7868 4102
rect 7992 4056 8053 4102
rect 8135 4096 8335 4106
rect 6175 4029 6375 4040
rect 8135 4040 8154 4096
rect 8210 4040 8264 4096
rect 8320 4040 8335 4096
rect 8135 4029 8335 4040
rect 8415 4095 8615 4106
rect 8415 4039 8435 4095
rect 8491 4039 8545 4095
rect 8601 4039 8615 4095
rect 8697 4056 8708 4102
rect 8830 4058 8876 4274
rect 9989 4276 10006 4322
rect 10052 4276 10069 4322
rect 9989 4224 10069 4276
rect 9484 4209 9681 4214
rect 9484 4195 9502 4209
rect 9442 4194 9502 4195
rect 9396 4153 9502 4194
rect 9558 4153 9612 4209
rect 9668 4153 9681 4209
rect 9396 4148 9681 4153
rect 9989 4178 10006 4224
rect 10052 4178 10069 4224
rect 8882 4056 8893 4102
rect 8975 4096 9175 4106
rect 9396 4102 9442 4148
rect 9989 4126 10069 4178
rect 9989 4107 10006 4126
rect 8415 4029 8615 4039
rect 8975 4040 8996 4096
rect 9052 4040 9106 4096
rect 9162 4040 9175 4096
rect 9257 4056 9268 4102
rect 9396 4056 9453 4102
rect 9537 4056 9548 4102
rect 9722 4080 10006 4107
rect 10052 4080 10069 4126
rect 9722 4050 10069 4080
rect 8975 4029 9175 4040
rect -39 3982 -22 4028
rect 24 3982 41 4028
rect 9989 4028 10069 4050
rect -39 3930 41 3982
rect -39 3884 -22 3930
rect 24 3884 41 3930
rect 88 3985 285 3990
rect 88 3929 101 3985
rect 157 3929 211 3985
rect 267 3983 285 3985
rect 9733 3985 9935 3990
rect 9733 3983 9751 3985
rect 267 3933 2038 3983
rect 267 3929 285 3933
rect 88 3924 285 3929
rect -39 3832 41 3884
rect -39 3786 -22 3832
rect 24 3786 41 3832
rect -39 3777 41 3786
rect 857 3793 1054 3798
rect -39 3734 327 3777
rect 857 3770 870 3793
rect -39 3688 -22 3734
rect 24 3720 327 3734
rect 577 3737 870 3770
rect 926 3737 980 3793
rect 1036 3737 1054 3793
rect 1415 3795 1612 3800
rect 1322 3767 1333 3770
rect 577 3732 1054 3737
rect 577 3724 1053 3732
rect 1232 3724 1333 3767
rect 1415 3739 1428 3795
rect 1484 3739 1538 3795
rect 1594 3770 1612 3795
rect 1988 3770 2038 3933
rect 3512 3933 6518 3983
rect 2255 3782 2455 3797
rect 1594 3739 1613 3770
rect 1415 3734 1613 3739
rect 1417 3724 1428 3734
rect 24 3688 41 3720
rect -39 3636 41 3688
rect -39 3590 -22 3636
rect 24 3590 41 3636
rect -39 3538 41 3590
rect 92 3612 289 3617
rect 92 3556 105 3612
rect 161 3556 215 3612
rect 271 3610 289 3612
rect 1232 3610 1322 3724
rect 1429 3610 1482 3734
rect 1602 3724 1613 3734
rect 1697 3724 1708 3770
rect 271 3557 1482 3610
rect 271 3556 289 3557
rect 92 3551 289 3556
rect 1429 3550 1482 3557
rect 1827 3605 1880 3769
rect 1882 3724 1893 3770
rect 1977 3726 2038 3770
rect 1977 3724 1988 3726
rect 2162 3724 2173 3770
rect 2255 3726 2267 3782
rect 2323 3726 2377 3782
rect 2433 3726 2455 3782
rect 3095 3782 3295 3797
rect 2255 3720 2455 3726
rect 2537 3724 2584 3770
rect 2680 3724 2877 3770
rect 2973 3724 3013 3770
rect 3095 3726 3117 3782
rect 3173 3726 3227 3782
rect 3283 3726 3295 3782
rect 3512 3770 3562 3933
rect 4333 3822 5697 3872
rect 4333 3796 4402 3822
rect 4332 3770 4402 3796
rect 5628 3796 5697 3822
rect 5628 3770 5698 3796
rect 6468 3770 6518 3933
rect 7992 3933 9751 3983
rect 6735 3782 6935 3797
rect 3095 3720 3295 3726
rect 3377 3724 3388 3770
rect 3512 3726 3573 3770
rect 3562 3724 3573 3726
rect 3657 3724 3668 3770
rect 3670 3605 3723 3769
rect 3842 3724 3853 3770
rect 3937 3724 3948 3770
rect 1827 3552 3723 3605
rect 4068 3610 4121 3767
rect 4122 3724 4133 3770
rect 4217 3724 4228 3770
rect 4332 3726 4413 3770
rect 4402 3724 4413 3726
rect 4497 3724 4973 3770
rect 5057 3724 5533 3770
rect 5617 3726 5698 3770
rect 5617 3724 5628 3726
rect 5802 3724 5813 3770
rect 5897 3724 5908 3770
rect 5909 3610 5962 3767
rect 6082 3724 6093 3770
rect 6177 3724 6188 3770
rect 4068 3557 5962 3610
rect 4068 3550 4121 3557
rect 5909 3550 5962 3557
rect 6307 3605 6360 3769
rect 6362 3724 6373 3770
rect 6457 3726 6518 3770
rect 6457 3724 6468 3726
rect 6642 3724 6653 3770
rect 6735 3726 6747 3782
rect 6803 3726 6857 3782
rect 6913 3726 6935 3782
rect 7575 3782 7775 3797
rect 6735 3720 6935 3726
rect 7017 3724 7493 3770
rect 7575 3726 7597 3782
rect 7653 3726 7707 3782
rect 7763 3726 7775 3782
rect 7992 3770 8042 3933
rect 9733 3929 9751 3933
rect 9807 3929 9861 3985
rect 9917 3929 9935 3985
rect 9733 3924 9935 3929
rect 9989 3982 10006 4028
rect 10052 3982 10069 4028
rect 9989 3930 10069 3982
rect 9483 3882 9680 3887
rect 9483 3872 9501 3882
rect 8813 3826 9501 3872
rect 9557 3826 9611 3882
rect 9667 3826 9680 3882
rect 8813 3822 9680 3826
rect 8813 3796 8882 3822
rect 9483 3821 9680 3822
rect 9989 3884 10006 3930
rect 10052 3884 10069 3930
rect 9989 3832 10069 3884
rect 8812 3770 8882 3796
rect 9989 3786 10006 3832
rect 10052 3786 10069 3832
rect 9989 3777 10069 3786
rect 7575 3720 7775 3726
rect 7857 3724 7868 3770
rect 7992 3726 8053 3770
rect 8042 3724 8053 3726
rect 8137 3724 8148 3770
rect 8150 3605 8203 3769
rect 8322 3724 8333 3770
rect 8417 3724 8428 3770
rect 6307 3552 8203 3605
rect 8548 3610 8601 3767
rect 8602 3724 8613 3770
rect 8697 3724 8708 3770
rect 8812 3726 8893 3770
rect 8882 3724 8893 3726
rect 8977 3724 9453 3770
rect 9537 3724 9548 3770
rect 9710 3734 10069 3777
rect 9710 3720 10006 3734
rect 9989 3688 10006 3720
rect 10052 3688 10069 3734
rect 9989 3636 10069 3688
rect 9713 3612 9910 3617
rect 9713 3610 9731 3612
rect 8548 3557 9731 3610
rect 8548 3550 8601 3557
rect 9713 3556 9731 3557
rect 9787 3556 9841 3612
rect 9897 3556 9910 3612
rect 9713 3551 9910 3556
rect 9989 3590 10006 3636
rect 10052 3590 10069 3636
rect -39 3492 -22 3538
rect 24 3492 41 3538
rect -39 3457 41 3492
rect 9989 3538 10069 3590
rect 9989 3492 10006 3538
rect 10052 3492 10069 3538
rect 9989 3457 10069 3492
rect -39 3440 10069 3457
rect -39 3394 -22 3440
rect 24 3394 76 3440
rect 122 3394 174 3440
rect 220 3394 272 3440
rect 318 3394 370 3440
rect 416 3394 468 3440
rect 514 3394 566 3440
rect 612 3394 664 3440
rect 710 3394 762 3440
rect 808 3394 860 3440
rect 906 3394 958 3440
rect 1004 3394 1056 3440
rect 1102 3394 1154 3440
rect 1200 3394 1252 3440
rect 1298 3394 1350 3440
rect 1396 3394 1448 3440
rect 1494 3394 1546 3440
rect 1592 3394 1644 3440
rect 1690 3394 1742 3440
rect 1788 3394 1840 3440
rect 1886 3394 1938 3440
rect 1984 3394 2036 3440
rect 2082 3394 2134 3440
rect 2180 3394 2232 3440
rect 2278 3394 2330 3440
rect 2376 3394 2428 3440
rect 2474 3394 2526 3440
rect 2572 3394 2624 3440
rect 2670 3394 2722 3440
rect 2768 3394 2820 3440
rect 2866 3394 2918 3440
rect 2964 3394 3016 3440
rect 3062 3394 3114 3440
rect 3160 3394 3212 3440
rect 3258 3394 3310 3440
rect 3356 3394 3408 3440
rect 3454 3394 3506 3440
rect 3552 3394 3604 3440
rect 3650 3394 3702 3440
rect 3748 3394 3800 3440
rect 3846 3394 3898 3440
rect 3944 3394 3996 3440
rect 4042 3394 4094 3440
rect 4140 3394 4192 3440
rect 4238 3394 4290 3440
rect 4336 3394 4388 3440
rect 4434 3394 4486 3440
rect 4532 3394 4584 3440
rect 4630 3394 4682 3440
rect 4728 3394 4780 3440
rect 4826 3394 4878 3440
rect 4924 3394 4976 3440
rect 5022 3394 5074 3440
rect 5120 3394 5172 3440
rect 5218 3394 5270 3440
rect 5316 3394 5368 3440
rect 5414 3394 5466 3440
rect 5512 3394 5564 3440
rect 5610 3394 5662 3440
rect 5708 3394 5760 3440
rect 5806 3394 5858 3440
rect 5904 3394 5956 3440
rect 6002 3394 6054 3440
rect 6100 3394 6152 3440
rect 6198 3394 6250 3440
rect 6296 3394 6348 3440
rect 6394 3394 6446 3440
rect 6492 3394 6544 3440
rect 6590 3394 6642 3440
rect 6688 3394 6740 3440
rect 6786 3394 6838 3440
rect 6884 3394 6936 3440
rect 6982 3394 7034 3440
rect 7080 3394 7132 3440
rect 7178 3394 7230 3440
rect 7276 3394 7328 3440
rect 7374 3394 7426 3440
rect 7472 3394 7524 3440
rect 7570 3394 7622 3440
rect 7668 3394 7720 3440
rect 7766 3394 7818 3440
rect 7864 3394 7916 3440
rect 7962 3394 8014 3440
rect 8060 3394 8112 3440
rect 8158 3394 8210 3440
rect 8256 3394 8308 3440
rect 8354 3394 8406 3440
rect 8452 3394 8504 3440
rect 8550 3394 8602 3440
rect 8648 3394 8700 3440
rect 8746 3394 8798 3440
rect 8844 3394 8896 3440
rect 8942 3394 8994 3440
rect 9040 3394 9092 3440
rect 9138 3394 9190 3440
rect 9236 3394 9288 3440
rect 9334 3394 9386 3440
rect 9432 3394 9484 3440
rect 9530 3394 9582 3440
rect 9628 3394 9680 3440
rect 9726 3394 9778 3440
rect 9824 3394 9876 3440
rect 9922 3394 10006 3440
rect 10052 3394 10069 3440
rect -39 3377 10069 3394
rect 10122 4645 10185 4660
rect 10122 4589 10127 4645
rect 10183 4589 10185 4645
rect 10122 4535 10185 4589
rect 10122 4479 10127 4535
rect 10183 4479 10185 4535
rect 10122 3321 10185 4479
rect 10231 4106 10297 4121
rect 10231 4050 10236 4106
rect 10292 4050 10297 4106
rect 10231 3996 10297 4050
rect 10231 3940 10236 3996
rect 10292 3940 10297 3996
rect 10231 3924 10297 3940
rect 10231 3321 10294 3924
rect 10360 3904 10423 3919
rect 10360 3848 10365 3904
rect 10421 3848 10423 3904
rect 10360 3794 10423 3848
rect 10360 3738 10365 3794
rect 10421 3738 10423 3794
rect 10360 3321 10423 3738
rect 10481 3733 10545 3748
rect 10481 3677 10484 3733
rect 10540 3677 10545 3733
rect 10481 3623 10545 3677
rect 10481 3617 10484 3623
rect 10479 3567 10484 3617
rect 10540 3567 10545 3623
rect 10479 3551 10545 3567
rect 10479 3321 10542 3551
<< via1 >>
rect 2466 5456 2522 5512
rect 2576 5456 2632 5512
rect 2918 5456 2974 5512
rect 3028 5456 3084 5512
rect 1709 5345 1765 5401
rect 1819 5345 1875 5401
rect 6946 5456 7002 5512
rect 7056 5456 7112 5512
rect 7398 5456 7454 5512
rect 7508 5456 7564 5512
rect 3675 5345 3731 5401
rect 3785 5345 3841 5401
rect 6189 5345 6245 5401
rect 6299 5345 6355 5401
rect 8155 5345 8211 5401
rect 8265 5345 8321 5401
rect 349 4911 405 4967
rect 459 4911 515 4967
rect 867 5030 923 5086
rect 975 5030 1031 5086
rect -231 4696 -175 4752
rect -231 4586 -175 4642
rect 851 4844 907 4900
rect 961 4844 1017 4900
rect 1428 5037 1484 5093
rect 1538 5037 1594 5093
rect 1709 5034 1765 5090
rect 1819 5034 1875 5090
rect 2267 5031 2323 5087
rect 2377 5031 2433 5087
rect 3117 5031 3173 5087
rect 3227 5031 3283 5087
rect 3675 5034 3731 5090
rect 3785 5034 3841 5090
rect 1262 4909 1318 4965
rect 1372 4909 1428 4965
rect 3956 5037 4012 5093
rect 4066 5037 4122 5093
rect 4122 4909 4178 4965
rect 4232 4909 4288 4965
rect 4519 5030 4575 5086
rect 4627 5030 4683 5086
rect 5347 5030 5403 5086
rect 5455 5030 5511 5086
rect 870 4688 926 4744
rect 980 4688 1036 4744
rect 1150 4694 1206 4750
rect 1260 4694 1316 4750
rect 109 4575 165 4631
rect 219 4575 275 4631
rect 4531 4843 4587 4899
rect 4641 4843 4697 4899
rect 2269 4687 2325 4743
rect 2379 4687 2435 4743
rect 2548 4689 2604 4745
rect 2658 4689 2714 4745
rect 2836 4689 2892 4745
rect 2946 4689 3002 4745
rect 3115 4687 3171 4743
rect 3225 4687 3281 4743
rect 4234 4694 4290 4750
rect 4344 4694 4400 4750
rect 5331 4844 5387 4900
rect 5441 4844 5497 4900
rect 5908 5037 5964 5093
rect 6018 5037 6074 5093
rect 6189 5034 6245 5090
rect 6299 5034 6355 5090
rect 6747 5031 6803 5087
rect 6857 5031 6913 5087
rect 7597 5031 7653 5087
rect 7707 5031 7763 5087
rect 8155 5034 8211 5090
rect 8265 5034 8321 5090
rect 5742 4909 5798 4965
rect 5852 4909 5908 4965
rect 8436 5037 8492 5093
rect 8546 5037 8602 5093
rect 8602 4909 8658 4965
rect 8712 4909 8768 4965
rect 8999 5030 9055 5086
rect 9107 5030 9163 5086
rect 9713 4911 9771 4967
rect 9823 4911 9881 4967
rect 4514 4688 4570 4744
rect 4624 4688 4680 4744
rect 5350 4688 5406 4744
rect 5460 4688 5516 4744
rect 5630 4694 5686 4750
rect 5740 4694 5796 4750
rect 9011 4843 9067 4899
rect 9121 4843 9177 4899
rect 6749 4687 6805 4743
rect 6859 4687 6915 4743
rect 7028 4689 7084 4745
rect 7138 4689 7194 4745
rect 7316 4689 7372 4745
rect 7426 4689 7482 4745
rect 7595 4687 7651 4743
rect 7705 4687 7761 4743
rect 8714 4694 8770 4750
rect 8824 4694 8880 4750
rect 8994 4688 9050 4744
rect 9104 4688 9160 4744
rect -341 4391 -285 4447
rect -463 4269 -407 4325
rect -463 4159 -407 4215
rect -341 4281 -285 4337
rect -577 3677 -521 3733
rect -577 3567 -521 3623
rect 100 4270 156 4326
rect 210 4270 266 4326
rect 868 4382 924 4438
rect 978 4382 1034 4438
rect 1148 4383 1204 4439
rect 1258 4383 1314 4439
rect 2270 4381 2326 4437
rect 2380 4381 2436 4437
rect 2553 4381 2609 4437
rect 2663 4381 2719 4437
rect 2833 4381 2889 4437
rect 2943 4381 2999 4437
rect 3114 4381 3170 4437
rect 3224 4381 3280 4437
rect 4236 4383 4292 4439
rect 4346 4383 4402 4439
rect 4516 4382 4572 4438
rect 4626 4382 4682 4438
rect 5348 4382 5404 4438
rect 5458 4382 5514 4438
rect 5628 4383 5684 4439
rect 5738 4383 5794 4439
rect 6750 4381 6806 4437
rect 6860 4381 6916 4437
rect 7594 4381 7650 4437
rect 7704 4381 7760 4437
rect 8716 4383 8772 4439
rect 8826 4383 8882 4439
rect 366 4153 422 4209
rect 476 4153 532 4209
rect 868 4040 924 4096
rect 978 4040 1034 4096
rect 1261 4154 1317 4210
rect 1429 4039 1485 4095
rect 1539 4039 1595 4095
rect 4233 4154 4289 4210
rect 1710 4040 1766 4096
rect 1820 4040 1876 4096
rect 3674 4040 3730 4096
rect 3784 4040 3840 4096
rect 3955 4039 4011 4095
rect 4065 4039 4121 4095
rect 8996 4382 9052 4438
rect 9106 4382 9162 4438
rect 9503 4575 9559 4631
rect 9613 4575 9669 4631
rect 4516 4040 4572 4096
rect 4626 4040 4682 4096
rect 5348 4040 5404 4096
rect 5458 4040 5514 4096
rect 5741 4154 5797 4210
rect 5909 4039 5965 4095
rect 6019 4039 6075 4095
rect 8713 4154 8769 4210
rect 6190 4040 6246 4096
rect 6300 4040 6356 4096
rect 8154 4040 8210 4096
rect 8264 4040 8320 4096
rect 8435 4039 8491 4095
rect 8545 4039 8601 4095
rect 9502 4153 9558 4209
rect 9612 4153 9668 4209
rect 8996 4040 9052 4096
rect 9106 4040 9162 4096
rect 101 3929 157 3985
rect 211 3929 267 3985
rect 870 3737 926 3793
rect 980 3737 1036 3793
rect 1428 3739 1484 3795
rect 1538 3739 1594 3795
rect 105 3556 161 3612
rect 215 3556 271 3612
rect 2267 3726 2323 3782
rect 2377 3726 2433 3782
rect 3117 3726 3173 3782
rect 3227 3726 3283 3782
rect 6747 3726 6803 3782
rect 6857 3726 6913 3782
rect 7597 3726 7653 3782
rect 7707 3726 7763 3782
rect 9751 3929 9807 3985
rect 9861 3929 9917 3985
rect 9501 3826 9557 3882
rect 9611 3826 9667 3882
rect 9731 3556 9787 3612
rect 9841 3556 9897 3612
rect 10127 4589 10183 4645
rect 10127 4479 10183 4535
rect 10236 4050 10292 4106
rect 10236 3940 10292 3996
rect 10365 3848 10421 3904
rect 10365 3738 10421 3794
rect 10484 3677 10540 3733
rect 10484 3567 10540 3623
<< metal2 >>
rect 2454 5512 2644 5516
rect 2454 5456 2466 5512
rect 2522 5456 2576 5512
rect 2632 5456 2644 5512
rect 2454 5452 2644 5456
rect 2906 5512 3096 5516
rect 2906 5456 2918 5512
rect 2974 5456 3028 5512
rect 3084 5456 3096 5512
rect 2906 5452 3096 5456
rect 6934 5512 7124 5516
rect 6934 5456 6946 5512
rect 7002 5456 7056 5512
rect 7112 5456 7124 5512
rect 6934 5452 7124 5456
rect 7386 5512 7576 5516
rect 7386 5456 7398 5512
rect 7454 5456 7508 5512
rect 7564 5456 7576 5512
rect 7386 5452 7576 5456
rect 1709 5410 1765 5411
rect 1695 5401 1895 5410
rect 1695 5345 1709 5401
rect 1765 5345 1819 5401
rect 1875 5345 1895 5401
rect 1695 5333 1895 5345
rect 1428 5101 1484 5103
rect 855 5091 1055 5100
rect 603 5086 1055 5091
rect 603 5030 867 5086
rect 923 5030 975 5086
rect 1031 5030 1055 5086
rect 603 5025 1055 5030
rect 333 4967 530 4972
rect 333 4911 349 4967
rect 405 4911 459 4967
rect 515 4911 530 4967
rect 333 4906 530 4911
rect -236 4752 -170 4767
rect -236 4696 -231 4752
rect -175 4696 -170 4752
rect -236 4642 -170 4696
rect -236 4586 -231 4642
rect -175 4636 -170 4642
rect -175 4631 293 4636
rect -175 4586 109 4631
rect -236 4575 109 4586
rect 165 4575 219 4631
rect 275 4575 293 4631
rect -236 4570 293 4575
rect -346 4447 -280 4462
rect -346 4391 -341 4447
rect -285 4391 -280 4447
rect -468 4325 -402 4340
rect -468 4269 -463 4325
rect -407 4269 -402 4325
rect -468 4215 -402 4269
rect -346 4337 -280 4391
rect -346 4281 -341 4337
rect -285 4331 -280 4337
rect -285 4326 284 4331
rect -285 4281 100 4326
rect -346 4270 100 4281
rect 156 4270 210 4326
rect 266 4270 284 4326
rect -346 4265 284 4270
rect -468 4159 -463 4215
rect -407 4209 -402 4215
rect 430 4214 496 4906
rect 350 4209 547 4214
rect -407 4159 366 4209
rect -468 4153 366 4159
rect 422 4153 476 4209
rect 532 4153 547 4209
rect -468 4148 547 4153
rect -468 4143 350 4148
rect 88 3985 285 3990
rect 88 3929 101 3985
rect 157 3929 211 3985
rect 267 3929 285 3985
rect 88 3924 285 3929
rect -582 3733 -516 3748
rect -582 3677 -577 3733
rect -521 3677 -516 3733
rect -582 3623 -516 3677
rect -582 3567 -577 3623
rect -521 3617 -516 3623
rect 603 3676 669 5025
rect 855 5023 1055 5025
rect 1415 5093 1615 5101
rect 1415 5037 1428 5093
rect 1484 5037 1538 5093
rect 1594 5037 1615 5093
rect 1415 5024 1615 5037
rect 1695 5090 1895 5101
rect 1695 5034 1709 5090
rect 1765 5034 1819 5090
rect 1875 5034 1895 5090
rect 1695 5024 1895 5034
rect 2255 5087 2455 5101
rect 2255 5031 2267 5087
rect 2323 5031 2377 5087
rect 2433 5031 2455 5087
rect 2255 5024 2455 5031
rect 865 5020 921 5023
rect 1250 4965 1442 4968
rect 1250 4909 1262 4965
rect 1318 4909 1372 4965
rect 1428 4909 1442 4965
rect 1250 4906 1442 4909
rect 839 4900 1029 4904
rect 839 4844 851 4900
rect 907 4844 961 4900
rect 1017 4844 1029 4900
rect 839 4839 1029 4844
rect 851 4838 1029 4839
rect 1256 4758 1322 4906
rect 855 4744 1055 4756
rect 855 4688 870 4744
rect 926 4688 980 4744
rect 1036 4688 1055 4744
rect 855 4678 1055 4688
rect 1135 4750 1335 4758
rect 1135 4694 1150 4750
rect 1206 4694 1260 4750
rect 1316 4694 1335 4750
rect 1135 4681 1335 4694
rect 1812 4700 1884 5024
rect 2542 4758 2608 5452
rect 2942 4758 3008 5452
rect 3785 5410 3841 5411
rect 6189 5410 6245 5411
rect 3655 5401 3855 5410
rect 3655 5345 3675 5401
rect 3731 5345 3785 5401
rect 3841 5345 3855 5401
rect 3655 5333 3855 5345
rect 6175 5401 6375 5410
rect 6175 5345 6189 5401
rect 6245 5345 6299 5401
rect 6355 5345 6375 5401
rect 6175 5333 6375 5345
rect 4066 5101 4122 5103
rect 5908 5101 5964 5103
rect 3095 5087 3295 5101
rect 3095 5031 3117 5087
rect 3173 5031 3227 5087
rect 3283 5031 3295 5087
rect 3095 5024 3295 5031
rect 3655 5090 3855 5101
rect 3655 5034 3675 5090
rect 3731 5034 3785 5090
rect 3841 5034 3855 5090
rect 3655 5024 3855 5034
rect 3935 5093 4135 5101
rect 3935 5037 3956 5093
rect 4012 5037 4066 5093
rect 4122 5037 4135 5093
rect 3935 5024 4135 5037
rect 4495 5091 4695 5100
rect 5335 5091 5535 5100
rect 4495 5086 4947 5091
rect 4495 5030 4519 5086
rect 4575 5030 4627 5086
rect 4683 5030 4947 5086
rect 4495 5025 4947 5030
rect 2255 4743 2455 4757
rect 2255 4700 2269 4743
rect 1812 4687 2269 4700
rect 2325 4687 2379 4743
rect 2435 4687 2455 4743
rect 1812 4677 2455 4687
rect 2535 4745 2735 4758
rect 2535 4689 2548 4745
rect 2604 4689 2658 4745
rect 2714 4689 2735 4745
rect 2535 4681 2735 4689
rect 2815 4745 3015 4758
rect 2815 4689 2836 4745
rect 2892 4689 2946 4745
rect 3002 4689 3015 4745
rect 2815 4681 3015 4689
rect 3095 4743 3295 4757
rect 3095 4687 3115 4743
rect 3171 4687 3225 4743
rect 3281 4700 3295 4743
rect 3666 4700 3738 5024
rect 4495 5023 4695 5025
rect 4629 5020 4685 5023
rect 4108 4965 4300 4968
rect 4108 4909 4122 4965
rect 4178 4909 4232 4965
rect 4288 4909 4300 4965
rect 4108 4906 4300 4909
rect 4228 4758 4294 4906
rect 4519 4899 4709 4904
rect 4519 4843 4531 4899
rect 4587 4843 4641 4899
rect 4697 4843 4709 4899
rect 4519 4838 4709 4843
rect 3281 4687 3738 4700
rect 2548 4679 2675 4681
rect 1812 4628 2370 4677
rect 855 4438 1055 4448
rect 855 4382 868 4438
rect 924 4382 978 4438
rect 1034 4382 1055 4438
rect 855 4371 1055 4382
rect 1135 4439 1335 4449
rect 1135 4383 1148 4439
rect 1204 4383 1258 4439
rect 1314 4383 1335 4439
rect 1135 4372 1335 4383
rect 2255 4437 2455 4449
rect 2599 4442 2675 4679
rect 2890 4679 3002 4681
rect 2890 4442 2966 4679
rect 3095 4677 3738 4687
rect 4215 4750 4415 4758
rect 4215 4694 4234 4750
rect 4290 4694 4344 4750
rect 4400 4694 4415 4750
rect 4215 4681 4415 4694
rect 4495 4744 4695 4756
rect 4495 4688 4514 4744
rect 4570 4688 4624 4744
rect 4680 4688 4695 4744
rect 4495 4678 4695 4688
rect 3180 4628 3738 4677
rect 2255 4381 2270 4437
rect 2326 4381 2380 4437
rect 2436 4381 2455 4437
rect 1256 4215 1322 4372
rect 2255 4371 2455 4381
rect 2537 4437 2734 4442
rect 2537 4381 2553 4437
rect 2609 4381 2663 4437
rect 2719 4381 2734 4437
rect 2537 4376 2734 4381
rect 2817 4437 3014 4442
rect 2817 4381 2833 4437
rect 2889 4381 2943 4437
rect 2999 4381 3014 4437
rect 2817 4376 3014 4381
rect 3095 4437 3295 4449
rect 3095 4381 3114 4437
rect 3170 4381 3224 4437
rect 3280 4381 3295 4437
rect 3095 4371 3295 4381
rect 4215 4439 4415 4449
rect 4215 4383 4236 4439
rect 4292 4383 4346 4439
rect 4402 4383 4415 4439
rect 4215 4372 4415 4383
rect 4495 4438 4695 4448
rect 4495 4382 4516 4438
rect 4572 4382 4626 4438
rect 4682 4382 4695 4438
rect 2272 4249 2340 4371
rect 1249 4210 1329 4215
rect 1249 4154 1261 4210
rect 1317 4154 1329 4210
rect 1249 4148 1329 4154
rect 1777 4181 2340 4249
rect 3210 4249 3278 4371
rect 3210 4181 3773 4249
rect 4228 4215 4294 4372
rect 4495 4371 4695 4382
rect 1777 4106 1845 4181
rect 3705 4106 3773 4181
rect 4221 4210 4301 4215
rect 4221 4154 4233 4210
rect 4289 4154 4301 4210
rect 4221 4148 4301 4154
rect 855 4096 1055 4106
rect 855 4040 868 4096
rect 924 4040 978 4096
rect 1034 4040 1055 4096
rect 855 4029 1055 4040
rect 1415 4095 1615 4106
rect 1415 4039 1429 4095
rect 1485 4039 1539 4095
rect 1595 4039 1615 4095
rect 1415 4029 1615 4039
rect 1695 4096 1895 4106
rect 1695 4040 1710 4096
rect 1766 4040 1820 4096
rect 1876 4040 1895 4096
rect 1695 4029 1895 4040
rect 3655 4096 3855 4106
rect 3655 4040 3674 4096
rect 3730 4040 3784 4096
rect 3840 4040 3855 4096
rect 3655 4029 3855 4040
rect 3935 4095 4135 4106
rect 3935 4039 3955 4095
rect 4011 4039 4065 4095
rect 4121 4039 4135 4095
rect 3935 4029 4135 4039
rect 4495 4096 4695 4106
rect 4495 4040 4516 4096
rect 4572 4040 4626 4096
rect 4682 4040 4695 4096
rect 4495 4029 4695 4040
rect 1477 3800 1547 4029
rect 857 3793 1054 3798
rect 857 3737 870 3793
rect 926 3737 980 3793
rect 1036 3737 1054 3793
rect 857 3732 1054 3737
rect 1415 3795 1612 3800
rect 1415 3739 1428 3795
rect 1484 3739 1538 3795
rect 1594 3739 1612 3795
rect 1415 3734 1612 3739
rect 2255 3782 2455 3797
rect 2255 3726 2267 3782
rect 2323 3726 2377 3782
rect 2433 3726 2455 3782
rect 2255 3720 2455 3726
rect 3095 3782 3295 3797
rect 3095 3726 3117 3782
rect 3173 3726 3227 3782
rect 3283 3726 3295 3782
rect 3095 3720 3295 3726
rect 2255 3716 2323 3720
rect 3227 3716 3295 3720
rect 2255 3676 2321 3716
rect -521 3612 289 3617
rect -521 3567 105 3612
rect -582 3556 105 3567
rect 161 3556 215 3612
rect 271 3556 289 3612
rect 603 3610 2321 3676
rect 3229 3676 3295 3716
rect 4881 3676 4947 5025
rect 3229 3610 4947 3676
rect 5083 5086 5535 5091
rect 5083 5030 5347 5086
rect 5403 5030 5455 5086
rect 5511 5030 5535 5086
rect 5083 5025 5535 5030
rect 5083 3676 5149 5025
rect 5335 5023 5535 5025
rect 5895 5093 6095 5101
rect 5895 5037 5908 5093
rect 5964 5037 6018 5093
rect 6074 5037 6095 5093
rect 5895 5024 6095 5037
rect 6175 5090 6375 5101
rect 6175 5034 6189 5090
rect 6245 5034 6299 5090
rect 6355 5034 6375 5090
rect 6175 5024 6375 5034
rect 6735 5087 6935 5101
rect 6735 5031 6747 5087
rect 6803 5031 6857 5087
rect 6913 5031 6935 5087
rect 6735 5024 6935 5031
rect 5345 5020 5401 5023
rect 5730 4965 5922 4968
rect 5730 4909 5742 4965
rect 5798 4909 5852 4965
rect 5908 4909 5922 4965
rect 5730 4906 5922 4909
rect 5319 4900 5509 4904
rect 5319 4844 5331 4900
rect 5387 4844 5441 4900
rect 5497 4844 5509 4900
rect 5319 4839 5509 4844
rect 5331 4838 5509 4839
rect 5736 4758 5802 4906
rect 5335 4744 5535 4756
rect 5335 4688 5350 4744
rect 5406 4688 5460 4744
rect 5516 4688 5535 4744
rect 5335 4678 5535 4688
rect 5615 4750 5815 4758
rect 5615 4694 5630 4750
rect 5686 4694 5740 4750
rect 5796 4694 5815 4750
rect 5615 4681 5815 4694
rect 6292 4700 6364 5024
rect 7022 4758 7088 5452
rect 7422 4758 7488 5452
rect 8265 5410 8321 5411
rect 8135 5401 8335 5410
rect 8135 5345 8155 5401
rect 8211 5345 8265 5401
rect 8321 5345 8335 5401
rect 8135 5333 8335 5345
rect 8546 5101 8602 5103
rect 7575 5087 7775 5101
rect 7575 5031 7597 5087
rect 7653 5031 7707 5087
rect 7763 5031 7775 5087
rect 7575 5024 7775 5031
rect 8135 5090 8335 5101
rect 8135 5034 8155 5090
rect 8211 5034 8265 5090
rect 8321 5034 8335 5090
rect 8135 5024 8335 5034
rect 8415 5093 8615 5101
rect 8415 5037 8436 5093
rect 8492 5037 8546 5093
rect 8602 5037 8615 5093
rect 8415 5024 8615 5037
rect 8975 5091 9175 5100
rect 8975 5086 9427 5091
rect 8975 5030 8999 5086
rect 9055 5030 9107 5086
rect 9163 5030 9427 5086
rect 8975 5025 9427 5030
rect 6735 4743 6935 4757
rect 6735 4700 6749 4743
rect 6292 4687 6749 4700
rect 6805 4687 6859 4743
rect 6915 4687 6935 4743
rect 6292 4677 6935 4687
rect 7015 4745 7215 4758
rect 7015 4689 7028 4745
rect 7084 4689 7138 4745
rect 7194 4689 7215 4745
rect 7015 4681 7215 4689
rect 7295 4745 7495 4758
rect 7295 4689 7316 4745
rect 7372 4689 7426 4745
rect 7482 4689 7495 4745
rect 7295 4681 7495 4689
rect 7575 4743 7775 4757
rect 7575 4687 7595 4743
rect 7651 4687 7705 4743
rect 7761 4700 7775 4743
rect 8146 4700 8218 5024
rect 8975 5023 9175 5025
rect 9109 5020 9165 5023
rect 8588 4965 8780 4968
rect 8588 4909 8602 4965
rect 8658 4909 8712 4965
rect 8768 4909 8780 4965
rect 8588 4906 8780 4909
rect 8708 4758 8774 4906
rect 8999 4899 9189 4904
rect 8999 4843 9011 4899
rect 9067 4843 9121 4899
rect 9177 4843 9189 4899
rect 8999 4838 9189 4843
rect 7761 4687 8218 4700
rect 7028 4679 7084 4681
rect 7426 4679 7482 4681
rect 7575 4677 8218 4687
rect 8695 4750 8895 4758
rect 8695 4694 8714 4750
rect 8770 4694 8824 4750
rect 8880 4694 8895 4750
rect 8695 4681 8895 4694
rect 8975 4744 9175 4756
rect 8975 4688 8994 4744
rect 9050 4688 9104 4744
rect 9160 4688 9175 4744
rect 8975 4678 9175 4688
rect 6292 4628 6850 4677
rect 7660 4628 8218 4677
rect 5335 4438 5535 4448
rect 5335 4382 5348 4438
rect 5404 4382 5458 4438
rect 5514 4382 5535 4438
rect 5335 4371 5535 4382
rect 5615 4439 5815 4449
rect 5615 4383 5628 4439
rect 5684 4383 5738 4439
rect 5794 4383 5815 4439
rect 5615 4372 5815 4383
rect 6735 4437 6935 4449
rect 6735 4381 6750 4437
rect 6806 4381 6860 4437
rect 6916 4381 6935 4437
rect 5736 4215 5802 4372
rect 6735 4371 6935 4381
rect 7575 4437 7775 4449
rect 7575 4381 7594 4437
rect 7650 4381 7704 4437
rect 7760 4381 7775 4437
rect 7575 4371 7775 4381
rect 8695 4439 8895 4449
rect 8695 4383 8716 4439
rect 8772 4383 8826 4439
rect 8882 4383 8895 4439
rect 8695 4372 8895 4383
rect 8975 4438 9175 4448
rect 8975 4382 8996 4438
rect 9052 4382 9106 4438
rect 9162 4382 9175 4438
rect 6752 4249 6820 4371
rect 5729 4210 5809 4215
rect 5729 4154 5741 4210
rect 5797 4154 5809 4210
rect 5729 4148 5809 4154
rect 6257 4181 6820 4249
rect 7690 4249 7758 4371
rect 7690 4181 8253 4249
rect 8708 4215 8774 4372
rect 8975 4371 9175 4382
rect 6257 4106 6325 4181
rect 8185 4106 8253 4181
rect 8701 4210 8781 4215
rect 8701 4154 8713 4210
rect 8769 4154 8781 4210
rect 8701 4148 8781 4154
rect 5335 4096 5535 4106
rect 5335 4040 5348 4096
rect 5404 4040 5458 4096
rect 5514 4040 5535 4096
rect 5335 4029 5535 4040
rect 5895 4095 6095 4106
rect 5895 4039 5909 4095
rect 5965 4039 6019 4095
rect 6075 4039 6095 4095
rect 5895 4029 6095 4039
rect 6175 4096 6375 4106
rect 6175 4040 6190 4096
rect 6246 4040 6300 4096
rect 6356 4040 6375 4096
rect 6175 4029 6375 4040
rect 8135 4096 8335 4106
rect 8135 4040 8154 4096
rect 8210 4040 8264 4096
rect 8320 4040 8335 4096
rect 8135 4029 8335 4040
rect 8415 4095 8615 4106
rect 8415 4039 8435 4095
rect 8491 4039 8545 4095
rect 8601 4039 8615 4095
rect 8415 4029 8615 4039
rect 8975 4096 9175 4106
rect 8975 4040 8996 4096
rect 9052 4040 9106 4096
rect 9162 4040 9175 4096
rect 8975 4029 9175 4040
rect 6735 3782 6935 3797
rect 6735 3726 6747 3782
rect 6803 3726 6857 3782
rect 6913 3726 6935 3782
rect 6735 3720 6935 3726
rect 7575 3782 7775 3797
rect 7575 3726 7597 3782
rect 7653 3726 7707 3782
rect 7763 3726 7775 3782
rect 7575 3720 7775 3726
rect 6735 3716 6803 3720
rect 7707 3716 7775 3720
rect 6735 3676 6801 3716
rect 5083 3610 6801 3676
rect 7709 3676 7775 3716
rect 9361 3676 9427 5025
rect 9700 4967 9897 4972
rect 9700 4911 9713 4967
rect 9771 4911 9823 4967
rect 9881 4911 9897 4967
rect 9700 4906 9897 4911
rect 10122 4645 10185 4660
rect 10122 4636 10127 4645
rect 9485 4631 10127 4636
rect 9485 4575 9503 4631
rect 9559 4575 9613 4631
rect 9669 4589 10127 4631
rect 10183 4636 10185 4645
rect 10183 4589 10311 4636
rect 9669 4575 10311 4589
rect 9485 4570 10311 4575
rect 10122 4535 10185 4570
rect 10122 4479 10127 4535
rect 10183 4479 10185 4535
rect 10122 4462 10185 4479
rect 9484 4209 9681 4214
rect 9484 4153 9502 4209
rect 9558 4153 9612 4209
rect 9668 4153 9681 4209
rect 9484 4148 9681 4153
rect 9555 3887 9621 4148
rect 10231 4106 10297 4121
rect 10231 4050 10236 4106
rect 10292 4050 10297 4106
rect 10231 3996 10297 4050
rect 10231 3990 10236 3996
rect 9733 3985 10236 3990
rect 9733 3929 9751 3985
rect 9807 3929 9861 3985
rect 9917 3940 10236 3985
rect 10292 3940 10297 3996
rect 9917 3929 10297 3940
rect 9733 3924 10297 3929
rect 10360 3904 10423 3919
rect 9483 3882 9680 3887
rect 9483 3826 9501 3882
rect 9557 3826 9611 3882
rect 9667 3826 9680 3882
rect 9483 3821 9680 3826
rect 9614 3788 9680 3821
rect 10360 3848 10365 3904
rect 10421 3848 10423 3904
rect 10360 3794 10423 3848
rect 10360 3788 10365 3794
rect 9614 3738 10365 3788
rect 10421 3738 10423 3794
rect 9614 3722 10423 3738
rect 10481 3733 10545 3748
rect 7709 3610 9427 3676
rect 10481 3677 10484 3733
rect 10540 3677 10545 3733
rect 10481 3623 10545 3677
rect 10481 3617 10484 3623
rect 9713 3612 10484 3617
rect -582 3551 289 3556
rect 9713 3556 9731 3612
rect 9787 3556 9841 3612
rect 9897 3567 10484 3612
rect 10540 3567 10545 3623
rect 9897 3556 10545 3567
rect 9713 3551 10545 3556
<< via2 >>
rect 1709 5345 1765 5401
rect 1819 5345 1875 5401
rect 109 4575 165 4631
rect 219 4575 275 4631
rect 101 3929 157 3985
rect 211 3929 267 3985
rect 1428 5037 1484 5093
rect 1538 5037 1594 5093
rect 2267 5031 2323 5087
rect 2377 5031 2433 5087
rect 851 4844 907 4900
rect 961 4844 1017 4900
rect 870 4688 926 4744
rect 980 4688 1036 4744
rect 3675 5345 3731 5401
rect 3785 5345 3841 5401
rect 6189 5345 6245 5401
rect 6299 5345 6355 5401
rect 3117 5031 3173 5087
rect 3227 5031 3283 5087
rect 3956 5037 4012 5093
rect 4066 5037 4122 5093
rect 4531 4843 4587 4899
rect 4641 4843 4697 4899
rect 868 4382 924 4438
rect 978 4382 1034 4438
rect 4514 4688 4570 4744
rect 4624 4688 4680 4744
rect 4516 4382 4572 4438
rect 4626 4382 4682 4438
rect 868 4040 924 4096
rect 978 4040 1034 4096
rect 1429 4039 1485 4095
rect 1539 4039 1595 4095
rect 3955 4039 4011 4095
rect 4065 4039 4121 4095
rect 4516 4040 4572 4096
rect 4626 4040 4682 4096
rect 870 3737 926 3793
rect 980 3737 1036 3793
rect 1428 3739 1484 3795
rect 1538 3739 1594 3795
rect 5908 5037 5964 5093
rect 6018 5037 6074 5093
rect 6747 5031 6803 5087
rect 6857 5031 6913 5087
rect 5331 4844 5387 4900
rect 5441 4844 5497 4900
rect 5350 4688 5406 4744
rect 5460 4688 5516 4744
rect 8155 5345 8211 5401
rect 8265 5345 8321 5401
rect 7597 5031 7653 5087
rect 7707 5031 7763 5087
rect 8436 5037 8492 5093
rect 8546 5037 8602 5093
rect 9011 4843 9067 4899
rect 9121 4843 9177 4899
rect 8994 4688 9050 4744
rect 9104 4688 9160 4744
rect 5348 4382 5404 4438
rect 5458 4382 5514 4438
rect 8996 4382 9052 4438
rect 9106 4382 9162 4438
rect 5348 4040 5404 4096
rect 5458 4040 5514 4096
rect 5909 4039 5965 4095
rect 6019 4039 6075 4095
rect 8435 4039 8491 4095
rect 8545 4039 8601 4095
rect 8996 4040 9052 4096
rect 9106 4040 9162 4096
rect 9713 4911 9769 4967
rect 9823 4911 9879 4967
rect 9751 3929 9807 3985
rect 9861 3929 9917 3985
<< metal3 >>
rect 1695 5401 1895 5410
rect 1695 5345 1709 5401
rect 1765 5345 1819 5401
rect 1875 5345 1895 5401
rect 1695 5333 1895 5345
rect 3655 5401 3855 5410
rect 3655 5345 3675 5401
rect 3731 5345 3785 5401
rect 3841 5345 3855 5401
rect 3655 5333 3855 5345
rect 6175 5401 6375 5410
rect 6175 5345 6189 5401
rect 6245 5345 6299 5401
rect 6355 5345 6375 5401
rect 6175 5333 6375 5345
rect 8135 5401 8335 5410
rect 8135 5345 8155 5401
rect 8211 5345 8265 5401
rect 8321 5345 8335 5401
rect 8135 5333 8335 5345
rect 1415 5093 1615 5101
rect 1415 5037 1428 5093
rect 1484 5037 1538 5093
rect 1594 5037 1615 5093
rect 1415 5024 1615 5037
rect 1460 4904 1526 5024
rect 713 4900 1526 4904
rect 713 4844 851 4900
rect 907 4844 961 4900
rect 1017 4844 1526 4900
rect 713 4838 1526 4844
rect 855 4744 1055 4756
rect 855 4688 870 4744
rect 926 4688 980 4744
rect 1036 4710 1055 4744
rect 1036 4688 1057 4710
rect 855 4678 1057 4688
rect 932 4668 1057 4678
rect 1708 4668 1772 5333
rect 2255 5087 2455 5101
rect 2255 5031 2267 5087
rect 2323 5031 2377 5087
rect 2433 5031 2455 5087
rect 2255 5024 2455 5031
rect 3095 5087 3295 5101
rect 3095 5031 3117 5087
rect 3173 5031 3227 5087
rect 3283 5031 3295 5087
rect 3095 5024 3295 5031
rect 96 4631 293 4636
rect 96 4575 109 4631
rect 165 4575 219 4631
rect 275 4575 293 4631
rect 96 4570 293 4575
rect 932 4604 1772 4668
rect 160 3990 226 4570
rect 932 4448 1016 4604
rect 855 4438 1055 4448
rect 855 4382 868 4438
rect 924 4382 978 4438
rect 1034 4382 1055 4438
rect 855 4371 1055 4382
rect 982 4286 1055 4371
rect 982 4213 1514 4286
rect 1441 4106 1514 4213
rect 855 4096 1055 4106
rect 855 4040 868 4096
rect 924 4040 978 4096
rect 1034 4040 1055 4096
rect 855 4029 1055 4040
rect 1415 4095 1615 4106
rect 1415 4039 1429 4095
rect 1485 4039 1539 4095
rect 1595 4039 1615 4095
rect 1415 4029 1615 4039
rect 88 3985 285 3990
rect 88 3929 101 3985
rect 157 3929 211 3985
rect 267 3929 285 3985
rect 88 3924 285 3929
rect 954 3973 1055 4029
rect 2352 3973 2418 5024
rect 954 3907 2418 3973
rect 3132 3973 3198 5024
rect 3778 4668 3842 5333
rect 3935 5093 4135 5101
rect 3935 5037 3956 5093
rect 4012 5037 4066 5093
rect 4122 5037 4135 5093
rect 3935 5024 4135 5037
rect 5895 5093 6095 5101
rect 5895 5037 5908 5093
rect 5964 5037 6018 5093
rect 6074 5037 6095 5093
rect 5895 5024 6095 5037
rect 4024 4904 4090 5024
rect 5940 4904 6006 5024
rect 4024 4899 4709 4904
rect 4024 4843 4531 4899
rect 4587 4843 4641 4899
rect 4697 4843 4709 4899
rect 4024 4838 4709 4843
rect 5193 4900 6006 4904
rect 5193 4844 5331 4900
rect 5387 4844 5441 4900
rect 5497 4844 6006 4900
rect 5193 4838 6006 4844
rect 4495 4744 4695 4756
rect 4495 4688 4514 4744
rect 4570 4688 4624 4744
rect 4680 4688 4695 4744
rect 4495 4678 4695 4688
rect 5335 4744 5535 4756
rect 5335 4688 5350 4744
rect 5406 4688 5460 4744
rect 5516 4688 5535 4744
rect 5335 4678 5535 4688
rect 4495 4668 4607 4678
rect 3778 4604 4607 4668
rect 5420 4668 5535 4678
rect 6188 4668 6252 5333
rect 6735 5087 6935 5101
rect 6735 5031 6747 5087
rect 6803 5031 6857 5087
rect 6913 5031 6935 5087
rect 6735 5024 6935 5031
rect 7575 5087 7775 5101
rect 7575 5031 7597 5087
rect 7653 5031 7707 5087
rect 7763 5031 7775 5087
rect 7575 5024 7775 5031
rect 5420 4604 6252 4668
rect 4495 4438 4695 4448
rect 4495 4382 4516 4438
rect 4572 4382 4626 4438
rect 4682 4382 4695 4438
rect 4495 4371 4695 4382
rect 5335 4438 5535 4448
rect 5335 4382 5348 4438
rect 5404 4382 5458 4438
rect 5514 4382 5535 4438
rect 5335 4371 5535 4382
rect 4495 4286 4568 4371
rect 4036 4213 4568 4286
rect 5462 4286 5535 4371
rect 5462 4213 5994 4286
rect 4036 4106 4109 4213
rect 5921 4106 5994 4213
rect 3935 4095 4135 4106
rect 3935 4039 3955 4095
rect 4011 4039 4065 4095
rect 4121 4039 4135 4095
rect 3935 4029 4135 4039
rect 4495 4096 4695 4106
rect 4495 4040 4516 4096
rect 4572 4040 4626 4096
rect 4682 4040 4695 4096
rect 4495 4029 4695 4040
rect 5335 4096 5535 4106
rect 5335 4040 5348 4096
rect 5404 4040 5458 4096
rect 5514 4040 5535 4096
rect 5335 4029 5535 4040
rect 5895 4095 6095 4106
rect 5895 4039 5909 4095
rect 5965 4039 6019 4095
rect 6075 4039 6095 4095
rect 5895 4029 6095 4039
rect 4495 3973 4596 4029
rect 3132 3907 4596 3973
rect 5434 3973 5535 4029
rect 6832 3973 6898 5024
rect 5434 3907 6898 3973
rect 7612 3973 7678 5024
rect 8258 4668 8322 5333
rect 8415 5093 8615 5101
rect 8415 5037 8436 5093
rect 8492 5037 8546 5093
rect 8602 5037 8615 5093
rect 8415 5024 8615 5037
rect 8504 4904 8570 5024
rect 9700 4967 9897 4972
rect 9700 4911 9713 4967
rect 9769 4911 9823 4967
rect 9879 4911 9897 4967
rect 9700 4906 9897 4911
rect 8504 4899 9189 4904
rect 8504 4843 9011 4899
rect 9067 4843 9121 4899
rect 9177 4843 9189 4899
rect 8504 4838 9189 4843
rect 8975 4744 9175 4756
rect 8975 4688 8994 4744
rect 9050 4688 9104 4744
rect 9160 4688 9175 4744
rect 8975 4678 9175 4688
rect 8975 4668 9087 4678
rect 8258 4604 9087 4668
rect 8975 4438 9175 4448
rect 8975 4382 8996 4438
rect 9052 4382 9106 4438
rect 9162 4382 9175 4438
rect 8975 4371 9175 4382
rect 8975 4286 9048 4371
rect 8516 4213 9048 4286
rect 8516 4106 8589 4213
rect 8415 4095 8615 4106
rect 8415 4039 8435 4095
rect 8491 4039 8545 4095
rect 8601 4039 8615 4095
rect 8415 4029 8615 4039
rect 8975 4096 9175 4106
rect 8975 4040 8996 4096
rect 9052 4040 9106 4096
rect 9162 4040 9175 4096
rect 8975 4029 9175 4040
rect 8975 3973 9076 4029
rect 9801 3990 9867 4906
rect 7612 3907 9076 3973
rect 9738 3985 9935 3990
rect 9738 3929 9751 3985
rect 9807 3929 9861 3985
rect 9917 3929 9935 3985
rect 9738 3924 9935 3929
rect 954 3798 1055 3907
rect 857 3793 1055 3798
rect 857 3737 870 3793
rect 926 3737 980 3793
rect 1036 3769 1055 3793
rect 1415 3795 1612 3800
rect 1036 3737 1054 3769
rect 857 3732 1054 3737
rect 1415 3739 1428 3795
rect 1484 3739 1538 3795
rect 1594 3739 1612 3795
rect 1415 3734 1612 3739
use ppolyf_u_VRC5QE  ppolyf_u_VRC5QE_0
timestamp 1694610567
transform 1 0 5015 0 1 3913
box -4904 -386 4904 386
use ppolyf_u_VRC5QE  ppolyf_u_VRC5QE_1
timestamp 1694610567
transform 1 0 5015 0 1 5217
box -4904 -386 4904 386
use ppolyf_u_VRC5QE  ppolyf_u_VRC5QE_2
timestamp 1694610567
transform 1 0 5015 0 1 4565
box -4904 -386 4904 386
<< labels >>
flabel metal2 -186 4177 -186 4177 0 FreeSans 800 0 0 0 E
port 7 nsew
flabel metal2 10122 3943 10122 3943 0 FreeSans 800 0 0 0 D
port 13 nsew
flabel metal2 10113 3748 10113 3748 0 FreeSans 800 0 0 0 F
port 12 nsew
flabel metal2 10126 3578 10126 3578 0 FreeSans 800 0 0 0 H
port 11 nsew
flabel via1 -207 4594 -207 4594 0 FreeSans 800 0 0 0 C
port 9 nsew
flabel metal2 -220 3582 -220 3582 0 FreeSans 800 0 0 0 G
port 5 nsew
flabel metal2 10292 4594 10292 4594 0 FreeSans 800 0 0 0 B
port 3 nsew
flabel metal2 -238 4290 -238 4290 0 FreeSans 800 0 0 0 A
port 0 nsew
flabel metal1 4655 5669 4655 5669 0 FreeSans 1280 0 0 0 VDD
port 15 nsew
<< end >>
