magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1331 1045 1331
<< metal1 >>
rect -45 325 45 331
rect -45 -325 -39 325
rect 39 -325 45 325
rect -45 -331 45 -325
<< via1 >>
rect -39 -325 39 325
<< metal2 >>
rect -45 325 45 331
rect -45 -325 -39 325
rect 39 -325 45 325
rect -45 -331 45 -325
<< end >>
