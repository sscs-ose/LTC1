* NGSPICE file created from BIG_CM_MSB_flat.ext - technology: gf180mcuC

.subckt BIG_CM_MSB_flat IM_T IM OUT VSS
X0 VSS IM.t0 a_212_68.t1 VSS.t1 nfet_03v3 ad=16.9p pd=77.7u as=9.98p ps=38.9u w=38.4u l=0.5u
R0 IM_T.n0 IM_T.t0 291.928
R1 IM_T IM_T.n0 4.5185
R2 OUT OUT.t0 10.8529
R3 a_212_68.n0 a_212_68.t1 0.0858125
R4 VSS.n1 VSS.t1 125.394
R5 VSS.t1 VSS.t0 81.8625
R6 VSS VSS.n2 10.9035
R7 VSS VSS.n1 2.60241
R8 VSS.n1 VSS.n0 0.165206
R9 IM.n0 IM.t0 292.219
R10 IM IM.n0 4.9625
C0 IM OUT 0.00216f
C1 OUT IM_T 0.00816f
C2 IM IM_T 0.063f
.ends

