magic
tech gf180mcuD
magscale 1 10
timestamp 1713185578
<< checkpaint >>
rect -2446 -2422 2446 2422
<< nwell >>
rect -446 -422 446 422
<< pmos >>
rect -272 68 -160 292
rect -56 68 56 292
rect 160 68 272 292
rect -272 -292 -160 -68
rect -56 -292 56 -68
rect 160 -292 272 -68
<< pdiff >>
rect -360 250 -272 292
rect -360 110 -347 250
rect -301 110 -272 250
rect -360 68 -272 110
rect -160 250 -56 292
rect -160 110 -131 250
rect -85 110 -56 250
rect -160 68 -56 110
rect 56 250 160 292
rect 56 110 85 250
rect 131 110 160 250
rect 56 68 160 110
rect 272 250 360 292
rect 272 110 301 250
rect 347 110 360 250
rect 272 68 360 110
rect -360 -110 -272 -68
rect -360 -250 -347 -110
rect -301 -250 -272 -110
rect -360 -292 -272 -250
rect -160 -110 -56 -68
rect -160 -250 -131 -110
rect -85 -250 -56 -110
rect -160 -292 -56 -250
rect 56 -110 160 -68
rect 56 -250 85 -110
rect 131 -250 160 -110
rect 56 -292 160 -250
rect 272 -110 360 -68
rect 272 -250 301 -110
rect 347 -250 360 -110
rect 272 -292 360 -250
<< pdiffc >>
rect -347 110 -301 250
rect -131 110 -85 250
rect 85 110 131 250
rect 301 110 347 250
rect -347 -250 -301 -110
rect -131 -250 -85 -110
rect 85 -250 131 -110
rect 301 -250 347 -110
<< polysilicon >>
rect -272 292 -160 336
rect -56 292 56 336
rect 160 292 272 336
rect -272 24 -160 68
rect -56 24 56 68
rect 160 24 272 68
rect -272 -68 -160 -24
rect -56 -68 56 -24
rect 160 -68 272 -24
rect -272 -336 -160 -292
rect -56 -336 56 -292
rect 160 -336 272 -292
<< metal1 >>
rect -347 250 -301 290
rect -347 70 -301 110
rect -131 250 -85 290
rect -131 70 -85 110
rect 85 250 131 290
rect 85 70 131 110
rect 301 250 347 290
rect 301 70 347 110
rect -347 -110 -301 -70
rect -347 -290 -301 -250
rect -131 -110 -85 -70
rect -131 -290 -85 -250
rect 85 -110 131 -70
rect 85 -290 131 -250
rect 301 -110 347 -70
rect 301 -290 347 -250
<< end >>
