magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -2665 -2045 2665 2045
<< psubdiff >>
rect -665 23 665 45
rect -665 -23 -643 23
rect -597 -23 -519 23
rect -473 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 597 23
rect 643 -23 665 23
rect -665 -45 665 -23
<< psubdiffcont >>
rect -643 -23 -597 23
rect -519 -23 -473 23
rect -395 -23 -349 23
rect -271 -23 -225 23
rect -147 -23 -101 23
rect -23 -23 23 23
rect 101 -23 147 23
rect 225 -23 271 23
rect 349 -23 395 23
rect 473 -23 519 23
rect 597 -23 643 23
<< metal1 >>
rect -654 23 654 34
rect -654 -23 -643 23
rect -597 -23 -519 23
rect -473 -23 -395 23
rect -349 -23 -271 23
rect -225 -23 -147 23
rect -101 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 597 23
rect 643 -23 654 23
rect -654 -34 654 -23
<< end >>
