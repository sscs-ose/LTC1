* NGSPICE file created from CLK_div_3_mag_flat.ext - technology: gf180mcuC

.subckt CLK_div_3_mag_flat VSS Q1 Q0 Vdiv3 RST CLK VDD
X0 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 VDD.t46 VDD.t45 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 a_794_1309# CLK.t0 a_634_1309# VSS.t11 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X2 a_4375_1353# JK_FF_mag_0.nand3_mag_0.OUT VSS.t27 VSS.t26 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X3 Q0 JK_FF_mag_1.J.t3 a_5503_1353# VSS.t48 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X4 JK_FF_mag_0.nand3_mag_2.OUT Q0.t3 VDD.t5 VDD.t4 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X5 or_2_mag_0.GF_INV_MAG_1.IN Q0.t4 a_5060_2688# VDD.t109 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X6 Vdiv3 or_2_mag_0.GF_INV_MAG_1.IN VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X7 JK_FF_mag_0.nand2_mag_3.IN1 CLK.t1 VDD.t105 VDD.t104 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X8 JK_FF_mag_0.nand3_mag_0.OUT Q1.t3 VDD.t27 VDD.t26 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X9 a_2076_256# JK_FF_mag_1.nand3_mag_1.OUT VSS.t60 VSS.t59 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X10 a_5060_2688# or_2_mag_0.IN2 VDD.t11 VDD.t10 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X11 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t31 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X12 Q0 JK_FF_mag_0.nand2_mag_1.IN2 VDD.t3 VDD.t2 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X13 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t78 VDD.t77 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X14 a_788_212# CLK.t2 a_628_212# VSS.t10 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X15 JK_FF_mag_0.nand3_mag_2.OUT Q0.t5 a_3805_212# VSS.t63 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X16 VDD JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t89 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X17 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand3_mag_1.IN1 VDD.t9 VDD.t8 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X18 JK_FF_mag_1.nand3_mag_2.OUT Q1.t4 VDD.t101 VDD.t100 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X19 JK_FF_mag_0.nand3_mag_2.OUT VDD.t65 VDD.t67 VDD.t66 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X20 VDD Q0.t6 JK_FF_mag_1.J.t2 VDD.t97 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X21 JK_FF_mag_1.QB Q1.t5 a_2640_256# VSS.t66 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X22 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.QB VDD.t56 VDD.t55 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X23 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT VDD.t42 VDD.t41 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X24 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t18 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X25 VDD RST.t0 JK_FF_mag_1.nand3_mag_1.OUT VDD.t23 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X26 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_2076_256# VSS.t22 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X27 a_5657_256# JK_FF_mag_0.nand2_mag_4.IN2 VSS.t55 VSS.t54 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X28 VDD CLK.t3 JK_FF_mag_1.nand3_mag_0.OUT VDD.t94 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X29 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_2.OUT VDD.t37 VDD.t36 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X30 JK_FF_mag_1.nand3_mag_2.OUT Q1.t6 a_788_212# VSS.t30 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X31 a_3645_212# VDD.t110 VSS.t47 VSS.t46 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X32 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_1.J.t4 a_3811_1309# VSS.t14 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X33 a_4939_1353# JK_FF_mag_0.nand3_mag_1.IN1 VSS.t38 VSS.t37 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X34 VDD JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand2_mag_4.IN2 VDD.t28 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X35 a_1512_212# RST.t1 a_1352_212# VSS.t23 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X36 or_2_mag_0.GF_INV_MAG_1.IN or_2_mag_0.IN2 VSS.t20 VSS.t19 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X37 a_634_1309# JK_FF_mag_1.J.t5 VSS.t32 VSS.t31 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X38 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_4939_1353# VSS.t25 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X39 a_5503_1353# JK_FF_mag_0.nand2_mag_1.IN2 VSS.t13 VSS.t12 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X40 a_5093_256# JK_FF_mag_0.nand3_mag_1.OUT VSS.t51 VSS.t50 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X41 JK_FF_mag_0.nand2_mag_3.IN1 CLK.t4 VSS.t9 VSS.t8 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X42 a_4369_212# JK_FF_mag_0.nand3_mag_2.OUT VSS.t29 VSS.t28 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X43 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_1.OUT a_1358_1353# VSS.t58 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X44 a_1922_1353# JK_FF_mag_1.nand3_mag_1.IN1 VSS.t18 VSS.t17 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X45 a_1358_1353# JK_FF_mag_1.nand3_mag_0.OUT VSS.t35 VSS.t34 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X46 VDD RST.t2 JK_FF_mag_0.nand3_mag_1.OUT VDD.t106 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X47 JK_FF_mag_1.J Q0.t7 a_5657_256# VSS.t15 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X48 Vdiv3 or_2_mag_0.GF_INV_MAG_1.IN VSS.t1 VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X49 VDD JK_FF_mag_1.QB Q1.t1 VDD.t52 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X50 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_3.IN1 a_1922_1353# VSS.t21 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X51 VSS Q0.t8 or_2_mag_0.GF_INV_MAG_1.IN VSS.t67 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
X52 Q1 JK_FF_mag_1.nand2_mag_1.IN2 VDD.t80 VDD.t79 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X53 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_1.J.t6 VDD.t82 VDD.t81 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X54 and2_mag_0.GF_INV_MAG_0.IN Q1.t7 a_4087_2452# VSS.t43 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X55 a_4529_212# RST.t3 a_4369_212# VSS.t33 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X56 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 a_5093_256# VSS.t24 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X57 a_4087_2452# CLK.t5 VSS.t7 VSS.t6 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X58 JK_FF_mag_1.nand2_mag_3.IN1 CLK.t6 VDD.t48 VDD.t47 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X59 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.J.t7 VDD.t103 VDD.t102 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X60 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_4.IN2 VDD.t93 VDD.t92 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X61 a_3811_1309# CLK.t7 a_3651_1309# VSS.t5 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X62 JK_FF_mag_1.nand3_mag_2.OUT VDD.t62 VDD.t64 VDD.t63 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X63 or_2_mag_0.IN2 and2_mag_0.GF_INV_MAG_0.IN VSS.t42 VSS.t41 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X64 VDD CLK.t8 JK_FF_mag_0.nand3_mag_2.OUT VDD.t49 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X65 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 VDD.t7 VDD.t6 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X66 Q1 JK_FF_mag_1.QB a_2486_1353# VSS.t40 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X67 a_628_212# VDD.t111 VSS.t45 VSS.t44 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X68 a_2486_1353# JK_FF_mag_1.nand2_mag_1.IN2 VSS.t53 VSS.t52 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X69 a_3805_212# CLK.t9 a_3645_212# VSS.t4 nfet_03v3 ad=0.172p pd=1.18u as=0.172p ps=1.18u w=0.66u l=0.28u
X70 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 a_1512_212# VSS.t16 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X71 VDD CLK.t10 JK_FF_mag_0.nand3_mag_0.OUT VDD.t68 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X72 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_2.OUT VDD.t86 VDD.t85 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X73 a_2640_256# JK_FF_mag_1.nand2_mag_4.IN2 VSS.t62 VSS.t61 nfet_03v3 ad=0.114p pd=0.96u as=0.194p ps=1.76u w=0.44u l=0.28u
X74 VDD JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t74 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X75 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT VDD.t35 VDD.t34 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X76 VDD JK_FF_mag_1.J.t8 Q0.t2 VDD.t71 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X77 JK_FF_mag_1.nand2_mag_3.IN1 CLK.t11 VSS.t3 VSS.t2 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X78 a_3651_1309# Q1.t8 VSS.t65 VSS.t64 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X79 JK_FF_mag_1.nand2_mag_4.IN2 JK_FF_mag_1.nand3_mag_1.OUT VDD.t88 VDD.t87 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X80 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 VDD.t44 VDD.t43 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X81 a_1352_212# JK_FF_mag_1.nand3_mag_2.OUT VSS.t57 VSS.t56 nfet_03v3 ad=0.172p pd=1.18u as=0.29p ps=2.2u w=0.66u l=0.28u
X82 VDD Q1.t9 JK_FF_mag_1.QB VDD.t59 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X83 JK_FF_mag_0.nand3_mag_1.OUT JK_FF_mag_0.nand3_mag_1.IN1 a_4529_212# VSS.t36 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X84 VDD Q1.t10 and2_mag_0.GF_INV_MAG_0.IN VDD.t38 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X85 or_2_mag_0.IN2 and2_mag_0.GF_INV_MAG_0.IN VDD.t58 VDD.t57 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X86 and2_mag_0.GF_INV_MAG_0.IN CLK.t12 VDD.t22 VDD.t21 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
X87 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.QB a_794_1309# VSS.t39 nfet_03v3 ad=0.29p pd=2.2u as=0.172p ps=1.18u w=0.66u l=0.28u
X88 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT a_4375_1353# VSS.t49 nfet_03v3 ad=0.194p pd=1.76u as=0.114p ps=0.96u w=0.44u l=0.28u
X89 VDD CLK.t13 JK_FF_mag_1.nand3_mag_2.OUT VDD.t12 pfet_03v3 ad=0.208p pd=1.32u as=0.208p ps=1.32u w=0.8u l=0.28u
X90 VDD JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 VDD.t15 pfet_03v3 ad=0.352p pd=2.48u as=0.208p ps=1.32u w=0.8u l=0.28u
X91 JK_FF_mag_1.J JK_FF_mag_0.nand2_mag_4.IN2 VDD.t84 VDD.t83 pfet_03v3 ad=0.208p pd=1.32u as=0.352p ps=2.48u w=0.8u l=0.28u
R0 VDD.n63 VDD.n62 11185.2
R1 VDD.t18 VDD.t79 961.905
R2 VDD.t55 VDD.t41 961.905
R3 VDD.t28 VDD.t83 765.152
R4 VDD.t43 VDD.t77 765.152
R5 VDD.t4 VDD.t36 765.152
R6 VDD.t31 VDD.t2 765.152
R7 VDD.t45 VDD.t74 765.152
R8 VDD.t81 VDD.t34 765.152
R9 VDD.t15 VDD.t92 765.152
R10 VDD.t6 VDD.t87 765.152
R11 VDD.t100 VDD.t85 765.152
R12 VDD.n62 VDD.t8 676.191
R13 VDD.n63 VDD.t102 485.714
R14 VDD.n110 VDD 429.187
R15 VDD VDD.n3 427.092
R16 VDD.t47 VDD.n63 426.44
R17 VDD.n8 VDD 420.935
R18 VDD.t26 VDD.n110 386.365
R19 VDD.t94 VDD.t55 380.952
R20 VDD.t38 VDD.n8 378.788
R21 VDD.n8 VDD.t10 322.223
R22 VDD.n3 VDD.t109 320.635
R23 VDD.t106 VDD.t43 303.031
R24 VDD.t49 VDD.t4 303.031
R25 VDD.t68 VDD.t81 303.031
R26 VDD.t23 VDD.t6 303.031
R27 VDD.t12 VDD.t100 303.031
R28 VDD.n62 VDD.t89 285.714
R29 VDD.n54 VDD.t52 242.857
R30 VDD.n56 VDD.t18 242.857
R31 VDD.t89 VDD.n58 242.857
R32 VDD.n61 VDD.t94 242.857
R33 VDD.n18 VDD.t97 193.183
R34 VDD.n20 VDD.t28 193.183
R35 VDD.n23 VDD.t106 193.183
R36 VDD.n26 VDD.t49 193.183
R37 VDD.n41 VDD.t71 193.183
R38 VDD.n42 VDD.t31 193.183
R39 VDD.n51 VDD.t74 193.183
R40 VDD.n111 VDD.t68 193.183
R41 VDD.n77 VDD.t59 193.183
R42 VDD.n79 VDD.t15 193.183
R43 VDD.n82 VDD.t23 193.183
R44 VDD.n85 VDD.t12 193.183
R45 VDD.n9 VDD.t38 193.183
R46 VDD.n7 VDD.t109 142.857
R47 VDD.t79 VDD.n54 138.095
R48 VDD.t8 VDD.n56 138.095
R49 VDD.t41 VDD.n58 138.095
R50 VDD.t102 VDD.n61 138.095
R51 VDD.t10 VDD.n7 111.112
R52 VDD.t83 VDD.n18 109.849
R53 VDD.t77 VDD.n20 109.849
R54 VDD.t36 VDD.n23 109.849
R55 VDD.n26 VDD.t66 109.849
R56 VDD.t2 VDD.n41 109.849
R57 VDD.n42 VDD.t45 109.849
R58 VDD.t34 VDD.n51 109.849
R59 VDD.n111 VDD.t26 109.849
R60 VDD.t92 VDD.n77 109.849
R61 VDD.t87 VDD.n79 109.849
R62 VDD.t85 VDD.n82 109.849
R63 VDD.n85 VDD.t63 109.849
R64 VDD.n9 VDD.t21 109.849
R65 VDD.n110 VDD.t104 59.702
R66 VDD.n3 VDD.t0 59.4064
R67 VDD.n8 VDD.t57 58.5371
R68 VDD.n88 VDD.t65 30.9379
R69 VDD.n87 VDD.t62 30.0062
R70 VDD.n88 VDD.t110 24.5101
R71 VDD.n93 VDD.t111 24.4392
R72 VDD VDD.t47 10.5649
R73 VDD.n94 VDD.n93 8.0005
R74 VDD.n90 VDD.n89 6.98838
R75 VDD.n27 VDD.n26 6.3005
R76 VDD.n30 VDD.n23 6.3005
R77 VDD.n33 VDD.n20 6.3005
R78 VDD.n36 VDD.n18 6.3005
R79 VDD.n65 VDD.n61 6.3005
R80 VDD.n68 VDD.n58 6.3005
R81 VDD.n71 VDD.n56 6.3005
R82 VDD.n74 VDD.n54 6.3005
R83 VDD.n97 VDD.n85 6.3005
R84 VDD.n100 VDD.n82 6.3005
R85 VDD.n103 VDD.n79 6.3005
R86 VDD.n106 VDD.n77 6.3005
R87 VDD.n51 VDD.n50 6.3005
R88 VDD.n43 VDD.n42 6.3005
R89 VDD.n41 VDD.n40 6.3005
R90 VDD.n7 VDD.n6 6.3005
R91 VDD.n10 VDD.n9 6.3005
R92 VDD.n112 VDD.n111 6.3005
R93 VDD.n27 VDD.t67 5.213
R94 VDD VDD.t48 5.16454
R95 VDD.n49 VDD.t35 5.13287
R96 VDD.n45 VDD.n13 5.13287
R97 VDD.n44 VDD.t46 5.13287
R98 VDD.n15 VDD.n14 5.13287
R99 VDD.n39 VDD.t3 5.13287
R100 VDD.n38 VDD.n16 5.13287
R101 VDD.n29 VDD.t37 5.13287
R102 VDD.n32 VDD.t78 5.13287
R103 VDD.n34 VDD.n19 5.13287
R104 VDD.n35 VDD.t84 5.13287
R105 VDD.n37 VDD.n17 5.13287
R106 VDD.n64 VDD.t103 5.13287
R107 VDD.n67 VDD.t42 5.13287
R108 VDD.n69 VDD.n57 5.13287
R109 VDD.n70 VDD.t9 5.13287
R110 VDD.n72 VDD.n55 5.13287
R111 VDD.n73 VDD.t80 5.13287
R112 VDD.n75 VDD.n53 5.13287
R113 VDD.n99 VDD.t86 5.13287
R114 VDD.n102 VDD.t88 5.13287
R115 VDD.n104 VDD.n78 5.13287
R116 VDD.n105 VDD.t93 5.13287
R117 VDD.n107 VDD.n76 5.13287
R118 VDD.n52 VDD.t27 5.13287
R119 VDD.n11 VDD.t22 5.13287
R120 VDD.n1 VDD.n0 5.13287
R121 VDD.n109 VDD.t105 5.09407
R122 VDD.n4 VDD.t1 5.09407
R123 VDD.n2 VDD.t58 5.09407
R124 VDD.n96 VDD.t64 4.8755
R125 VDD.n90 VDD.n86 4.51383
R126 VDD.n93 VDD.n92 4.5005
R127 VDD.n5 VDD.t11 4.12326
R128 VDD.n91 VDD.n87 3.61662
R129 VDD.n48 VDD.n47 2.85787
R130 VDD.n28 VDD.n25 2.85787
R131 VDD.n31 VDD.n22 2.85787
R132 VDD.n66 VDD.n60 2.85787
R133 VDD.n98 VDD.n84 2.85787
R134 VDD.n101 VDD.n81 2.85787
R135 VDD.n47 VDD.t82 2.2755
R136 VDD.n47 VDD.n46 2.2755
R137 VDD.n25 VDD.t5 2.2755
R138 VDD.n25 VDD.n24 2.2755
R139 VDD.n22 VDD.t44 2.2755
R140 VDD.n22 VDD.n21 2.2755
R141 VDD.n60 VDD.t56 2.2755
R142 VDD.n60 VDD.n59 2.2755
R143 VDD.n84 VDD.t101 2.2755
R144 VDD.n84 VDD.n83 2.2755
R145 VDD.n81 VDD.t7 2.2755
R146 VDD.n81 VDD.n80 2.2755
R147 VDD.n89 VDD.n88 2.11318
R148 VDD.n64 VDD 1.77285
R149 VDD VDD.n52 1.77285
R150 VDD.n92 VDD.n90 1.54785
R151 VDD.n38 VDD.n37 1.16167
R152 VDD.n108 VDD.n107 1.07428
R153 VDD.n93 VDD.n87 0.840632
R154 VDD.n12 VDD 0.468962
R155 VDD.n6 VDD.n4 0.388218
R156 VDD.n97 VDD.n96 0.337997
R157 VDD.n96 VDD.n95 0.328132
R158 VDD VDD.n11 0.273757
R159 VDD.n5 VDD 0.269151
R160 VDD.n32 VDD.n31 0.233919
R161 VDD.n29 VDD.n28 0.233919
R162 VDD.n102 VDD.n101 0.233919
R163 VDD.n99 VDD.n98 0.233919
R164 VDD.n2 VDD.n1 0.170231
R165 VDD.n108 VDD.n75 0.143501
R166 VDD.n35 VDD.n34 0.141016
R167 VDD.n73 VDD.n72 0.141016
R168 VDD.n70 VDD.n69 0.141016
R169 VDD.n105 VDD.n104 0.141016
R170 VDD.n39 VDD.n15 0.141016
R171 VDD.n45 VDD.n44 0.141016
R172 VDD.n109 VDD.n108 0.138896
R173 VDD.n67 VDD 0.122435
R174 VDD.n49 VDD 0.122435
R175 VDD VDD.n66 0.111984
R176 VDD VDD.n48 0.111984
R177 VDD VDD.n5 0.110164
R178 VDD.n37 VDD.n36 0.107339
R179 VDD.n34 VDD.n33 0.107339
R180 VDD.n75 VDD.n74 0.107339
R181 VDD.n72 VDD.n71 0.107339
R182 VDD.n69 VDD.n68 0.107339
R183 VDD.n107 VDD.n106 0.107339
R184 VDD.n104 VDD.n103 0.107339
R185 VDD.n40 VDD.n38 0.107339
R186 VDD.n43 VDD.n15 0.107339
R187 VDD.n50 VDD.n45 0.107339
R188 VDD.n10 VDD.n1 0.107339
R189 VDD.n89 VDD 0.106795
R190 VDD.n31 VDD 0.106177
R191 VDD.n28 VDD 0.106177
R192 VDD.n66 VDD 0.106177
R193 VDD.n101 VDD 0.106177
R194 VDD.n98 VDD 0.106177
R195 VDD.n30 VDD.n29 0.080629
R196 VDD.n65 VDD.n64 0.080629
R197 VDD.n100 VDD.n99 0.080629
R198 VDD VDD.n35 0.0794677
R199 VDD VDD.n32 0.0794677
R200 VDD VDD.n73 0.0794677
R201 VDD VDD.n70 0.0794677
R202 VDD VDD.n67 0.0794677
R203 VDD VDD.n105 0.0794677
R204 VDD VDD.n102 0.0794677
R205 VDD VDD.n39 0.0794677
R206 VDD.n44 VDD 0.0794677
R207 VDD VDD.n49 0.0794677
R208 VDD.n11 VDD 0.0759839
R209 VDD VDD.n109 0.0709717
R210 VDD.n4 VDD 0.0709717
R211 VDD VDD.n2 0.0709717
R212 VDD.n52 VDD.n12 0.0562419
R213 VDD.n95 VDD 0.049022
R214 VDD.n48 VDD.n12 0.0411452
R215 VDD.n94 VDD.n86 0.0358571
R216 VDD.n95 VDD.n94 0.03425
R217 VDD.n112 VDD.n12 0.0201154
R218 VDD.n6 VDD 0.00579412
R219 VDD VDD.n10 0.00514516
R220 VDD.n91 VDD.n86 0.00371429
R221 VDD.n92 VDD.n91 0.00210714
R222 VDD.n36 VDD 0.00166129
R223 VDD.n33 VDD 0.00166129
R224 VDD VDD.n30 0.00166129
R225 VDD VDD.n27 0.00166129
R226 VDD.n74 VDD 0.00166129
R227 VDD.n71 VDD 0.00166129
R228 VDD.n68 VDD 0.00166129
R229 VDD VDD.n65 0.00166129
R230 VDD.n106 VDD 0.00166129
R231 VDD.n103 VDD 0.00166129
R232 VDD VDD.n100 0.00166129
R233 VDD VDD.n97 0.00166129
R234 VDD.n40 VDD 0.00166129
R235 VDD VDD.n43 0.00166129
R236 VDD.n50 VDD 0.00166129
R237 VDD VDD.n112 0.00107692
R238 CLK.n9 CLK.t0 36.935
R239 CLK.n3 CLK.t2 36.935
R240 CLK.n24 CLK.t7 36.935
R241 CLK.n17 CLK.t9 36.935
R242 CLK.n13 CLK.t12 30.6315
R243 CLK.n37 CLK.t6 25.5364
R244 CLK.n29 CLK.t1 25.5364
R245 CLK.n13 CLK.t5 21.7275
R246 CLK.n9 CLK.t3 18.1962
R247 CLK.n3 CLK.t13 18.1962
R248 CLK.n24 CLK.t10 18.1962
R249 CLK.n17 CLK.t8 18.1962
R250 CLK.n29 CLK.t4 14.0749
R251 CLK.n37 CLK.t11 14.0749
R252 CLK.n21 CLK.n14 7.41477
R253 CLK.n35 CLK.n34 5.37352
R254 CLK.n5 CLK.n2 4.5005
R255 CLK.n5 CLK.n4 4.5005
R256 CLK.n8 CLK.n7 4.5005
R257 CLK.n10 CLK.n7 4.5005
R258 CLK.n19 CLK.n16 4.5005
R259 CLK.n19 CLK.n18 4.5005
R260 CLK.n23 CLK.n22 4.5005
R261 CLK.n25 CLK.n22 4.5005
R262 CLK.n30 CLK.n28 4.5005
R263 CLK.n31 CLK.n28 4.5005
R264 CLK.n39 CLK.n38 4.5005
R265 CLK.n40 CLK.n39 4.5005
R266 CLK.n12 CLK.n11 2.25107
R267 CLK.n27 CLK.n26 2.25107
R268 CLK.n33 CLK.n32 2.24385
R269 CLK.n36 CLK.n0 2.24385
R270 CLK.n4 CLK.n3 2.12175
R271 CLK.n18 CLK.n17 2.12175
R272 CLK.n10 CLK.n9 2.12075
R273 CLK.n25 CLK.n24 2.12075
R274 CLK.n14 CLK.n13 1.80496
R275 CLK.n7 CLK.n6 1.74297
R276 CLK.n21 CLK.n20 1.62464
R277 CLK.n6 CLK.n1 1.49778
R278 CLK.n20 CLK.n15 1.49778
R279 CLK.n30 CLK.n29 1.42706
R280 CLK.n38 CLK.n37 1.42706
R281 CLK.n35 CLK.n12 0.882596
R282 CLK.n34 CLK.n27 0.882596
R283 CLK.n31 CLK 0.1605
R284 CLK.n22 CLK.n21 0.118826
R285 CLK.n14 CLK 0.106541
R286 CLK.n34 CLK.n33 0.0726935
R287 CLK.n36 CLK.n35 0.0726935
R288 CLK CLK.n40 0.05925
R289 CLK.n8 CLK 0.0473512
R290 CLK.n2 CLK 0.0473512
R291 CLK.n23 CLK 0.0473512
R292 CLK.n16 CLK 0.0473512
R293 CLK.n11 CLK.n8 0.0361897
R294 CLK.n2 CLK.n1 0.0361897
R295 CLK.n26 CLK.n23 0.0361897
R296 CLK.n16 CLK.n15 0.0361897
R297 CLK.n32 CLK.n31 0.03175
R298 CLK.n40 CLK.n0 0.03175
R299 CLK.n33 CLK.n28 0.0205196
R300 CLK.n39 CLK.n36 0.0205196
R301 CLK.n6 CLK.n5 0.0131772
R302 CLK.n20 CLK.n19 0.0131772
R303 CLK.n12 CLK.n7 0.0122182
R304 CLK.n27 CLK.n22 0.0122182
R305 CLK.n11 CLK.n10 0.00515517
R306 CLK.n4 CLK.n1 0.00515517
R307 CLK.n26 CLK.n25 0.00515517
R308 CLK.n18 CLK.n15 0.00515517
R309 CLK.n32 CLK.n30 0.00175
R310 CLK.n38 CLK.n0 0.00175
R311 VSS.n42 VSS.n9 20976.7
R312 VSS.n26 VSS.t15 12337.5
R313 VSS.n55 VSS.t44 6806.14
R314 VSS.n26 VSS.n25 5448.69
R315 VSS.n41 VSS.n10 3893.61
R316 VSS.n25 VSS.t0 3035.98
R317 VSS.t41 VSS.t19 2781.65
R318 VSS.n10 VSS.t46 2623.57
R319 VSS.n10 VSS.t66 2617.37
R320 VSS.t24 VSS.t54 2505.73
R321 VSS.t63 VSS.t28 2505.73
R322 VSS.t22 VSS.t61 2505.73
R323 VSS.t30 VSS.t56 2505.73
R324 VSS.t25 VSS.t12 2307.56
R325 VSS.t37 VSS.t49 2307.56
R326 VSS.t26 VSS.t14 2307.56
R327 VSS.t8 VSS.t64 2307.56
R328 VSS.t21 VSS.t52 2307.56
R329 VSS.t17 VSS.t58 2307.56
R330 VSS.t39 VSS.t34 2307.56
R331 VSS.t48 VSS.n26 2073.37
R332 VSS.t40 VSS.n42 1713.53
R333 VSS.n42 VSS.n41 1565.03
R334 VSS.t33 VSS.t36 992.366
R335 VSS.t4 VSS.t63 992.366
R336 VSS.t23 VSS.t16 992.366
R337 VSS.t10 VSS.t30 992.366
R338 VSS.t14 VSS.t5 913.885
R339 VSS.t11 VSS.t39 913.885
R340 VSS.n12 VSS.t67 776.83
R341 VSS.t15 VSS.n0 595.42
R342 VSS.n1 VSS.t24 595.42
R343 VSS.n2 VSS.t33 595.42
R344 VSS.n3 VSS.t4 595.42
R345 VSS.t66 VSS.n5 595.42
R346 VSS.n6 VSS.t22 595.42
R347 VSS.n7 VSS.t23 595.42
R348 VSS.n8 VSS.t10 595.42
R349 VSS.t19 VSS.n12 554.879
R350 VSS.n29 VSS.t48 548.331
R351 VSS.n30 VSS.t25 548.331
R352 VSS.n38 VSS.t5 548.331
R353 VSS.n45 VSS.t40 548.331
R354 VSS.n46 VSS.t21 548.331
R355 VSS.n51 VSS.t58 548.331
R356 VSS.n52 VSS.t11 548.331
R357 VSS.n16 VSS.t43 546.41
R358 VSS.t54 VSS.n0 396.947
R359 VSS.n1 VSS.t50 396.947
R360 VSS.t28 VSS.n2 396.947
R361 VSS.t46 VSS.n3 396.947
R362 VSS.t61 VSS.n5 396.947
R363 VSS.n6 VSS.t59 396.947
R364 VSS.t56 VSS.n7 396.947
R365 VSS.t44 VSS.n8 396.947
R366 VSS.t12 VSS.n29 365.555
R367 VSS.n30 VSS.t37 365.555
R368 VSS.n33 VSS.t26 365.555
R369 VSS.t64 VSS.n38 365.555
R370 VSS.t52 VSS.n45 365.555
R371 VSS.n46 VSS.t17 365.555
R372 VSS.t34 VSS.n51 365.555
R373 VSS.n52 VSS.t31 365.555
R374 VSS.n16 VSS.t6 364.274
R375 VSS.n41 VSS.n40 119.948
R376 VSS.t0 VSS.n24 47.5615
R377 VSS.n40 VSS.t8 34.2711
R378 VSS.n13 VSS.t41 34.1511
R379 VSS.n55 VSS.t2 22.8476
R380 VSS.n56 VSS.n55 16.6241
R381 VSS.n56 VSS.t3 9.3736
R382 VSS.n39 VSS.t9 9.3736
R383 VSS.n15 VSS.t42 9.36521
R384 VSS.n21 VSS.n11 9.3221
R385 VSS.n19 VSS.t20 9.3221
R386 VSS.n22 VSS.t1 9.30652
R387 VSS VSS.t7 7.30633
R388 VSS.n73 VSS.t55 7.19156
R389 VSS.n71 VSS.t51 7.19156
R390 VSS.n64 VSS.t62 7.19156
R391 VSS.n62 VSS.t60 7.19156
R392 VSS.n27 VSS.t13 7.19156
R393 VSS.n32 VSS.t38 7.19156
R394 VSS.n35 VSS.t27 7.19156
R395 VSS.n43 VSS.t53 7.19156
R396 VSS.n48 VSS.t18 7.19156
R397 VSS.n49 VSS.t35 7.19156
R398 VSS.n69 VSS.t29 5.91399
R399 VSS.n67 VSS.t47 5.91399
R400 VSS.n60 VSS.t57 5.91399
R401 VSS.n58 VSS.t45 5.91399
R402 VSS.n36 VSS.t65 5.91399
R403 VSS.n54 VSS.t32 5.91399
R404 VSS.n14 VSS.n13 5.2005
R405 VSS.n17 VSS.n16 5.2005
R406 VSS.n24 VSS.n23 5.2005
R407 VSS.n20 VSS.n12 5.2005
R408 VSS.n29 VSS.n28 5.2005
R409 VSS.n31 VSS.n30 5.2005
R410 VSS.n34 VSS.n33 5.2005
R411 VSS.n38 VSS.n37 5.2005
R412 VSS.n40 VSS.n39 5.2005
R413 VSS.n45 VSS.n44 5.2005
R414 VSS.n47 VSS.n46 5.2005
R415 VSS.n51 VSS.n50 5.2005
R416 VSS.n53 VSS.n52 5.2005
R417 VSS.n59 VSS.n8 5.2005
R418 VSS.n61 VSS.n7 5.2005
R419 VSS.n63 VSS.n6 5.2005
R420 VSS.n65 VSS.n5 5.2005
R421 VSS.n68 VSS.n3 5.2005
R422 VSS.n70 VSS.n2 5.2005
R423 VSS.n72 VSS.n1 5.2005
R424 VSS.n74 VSS.n0 5.2005
R425 VSS.n58 VSS.n57 1.03335
R426 VSS.n66 VSS.n4 0.845914
R427 VSS.n71 VSS.n70 0.480225
R428 VSS.n69 VSS.n68 0.480225
R429 VSS.n62 VSS.n61 0.480225
R430 VSS.n60 VSS.n59 0.480225
R431 VSS.n27 VSS 0.343161
R432 VSS VSS.n32 0.343161
R433 VSS.n43 VSS 0.343161
R434 VSS VSS.n48 0.343161
R435 VSS.n73 VSS 0.343161
R436 VSS.n64 VSS 0.343161
R437 VSS.n19 VSS.n18 0.309418
R438 VSS.n37 VSS 0.289491
R439 VSS.n53 VSS 0.289491
R440 VSS.n18 VSS.n17 0.255008
R441 VSS VSS.n35 0.191234
R442 VSS.n49 VSS 0.191234
R443 VSS.n67 VSS.n66 0.187931
R444 VSS.n66 VSS 0.183803
R445 VSS.n22 VSS.n21 0.168119
R446 VSS.n18 VSS.n15 0.141461
R447 VSS.n57 VSS 0.137685
R448 VSS VSS.n4 0.137685
R449 VSS.n21 VSS.n20 0.136634
R450 VSS.n28 VSS.n27 0.118573
R451 VSS.n32 VSS.n31 0.118573
R452 VSS.n35 VSS.n34 0.118573
R453 VSS.n44 VSS.n43 0.118573
R454 VSS.n48 VSS.n47 0.118573
R455 VSS.n50 VSS.n49 0.118573
R456 VSS.n74 VSS.n73 0.118573
R457 VSS.n72 VSS.n71 0.118573
R458 VSS.n65 VSS.n64 0.118573
R459 VSS.n63 VSS.n62 0.118573
R460 VSS VSS.n19 0.115458
R461 VSS VSS.n36 0.115271
R462 VSS.n54 VSS 0.115271
R463 VSS VSS.n69 0.115271
R464 VSS VSS.n67 0.115271
R465 VSS VSS.n60 0.115271
R466 VSS VSS.n58 0.115271
R467 VSS.n36 VSS.n4 0.10206
R468 VSS.n57 VSS.n54 0.10206
R469 VSS.n15 VSS.n14 0.0589274
R470 VSS.n23 VSS.n22 0.0564843
R471 VSS.n28 VSS 0.00545413
R472 VSS.n31 VSS 0.00545413
R473 VSS.n34 VSS 0.00545413
R474 VSS.n44 VSS 0.00545413
R475 VSS.n47 VSS 0.00545413
R476 VSS.n50 VSS 0.00545413
R477 VSS VSS.n74 0.00545413
R478 VSS VSS.n72 0.00545413
R479 VSS VSS.n65 0.00545413
R480 VSS VSS.n63 0.00545413
R481 VSS.n37 VSS 0.00380275
R482 VSS.n17 VSS 0.00380275
R483 VSS VSS.n53 0.00380275
R484 VSS.n70 VSS 0.00380275
R485 VSS.n68 VSS 0.00380275
R486 VSS.n61 VSS 0.00380275
R487 VSS.n59 VSS 0.00380275
R488 VSS.n20 VSS 0.00352521
R489 VSS VSS.n56 0.00219811
R490 VSS.n39 VSS 0.00219811
R491 VSS.n14 VSS 0.00219811
R492 VSS.n23 VSS 0.00191732
R493 JK_FF_mag_1.J.n4 JK_FF_mag_1.J.t4 37.1986
R494 JK_FF_mag_1.J.n3 JK_FF_mag_1.J.t3 31.528
R495 JK_FF_mag_1.J.n2 JK_FF_mag_1.J.t7 30.5184
R496 JK_FF_mag_1.J.n2 JK_FF_mag_1.J.t5 24.7029
R497 JK_FF_mag_1.J.n4 JK_FF_mag_1.J.t6 17.6614
R498 JK_FF_mag_1.J.n3 JK_FF_mag_1.J.t8 15.3826
R499 JK_FF_mag_1.J.n0 JK_FF_mag_1.J 12.0843
R500 JK_FF_mag_1.J.n0 JK_FF_mag_1.J.n3 9.86691
R501 JK_FF_mag_1.J.n5 JK_FF_mag_1.J 6.09789
R502 JK_FF_mag_1.J.n1 JK_FF_mag_1.J.n7 2.99416
R503 JK_FF_mag_1.J.n7 JK_FF_mag_1.J.t2 2.2755
R504 JK_FF_mag_1.J.n7 JK_FF_mag_1.J.n6 2.2755
R505 JK_FF_mag_1.J.n1 JK_FF_mag_1.J.n5 2.2505
R506 JK_FF_mag_1.J.n0 JK_FF_mag_1.J 2.24173
R507 JK_FF_mag_1.J.n5 JK_FF_mag_1.J.n0 1.93723
R508 JK_FF_mag_1.J JK_FF_mag_1.J.n2 1.81225
R509 JK_FF_mag_1.J JK_FF_mag_1.J.n4 1.43709
R510 JK_FF_mag_1.J JK_FF_mag_1.J.n1 0.281955
R511 Q0.n2 Q0.t5 36.935
R512 Q0.n4 Q0.t7 31.528
R513 Q0.n0 Q0.t4 29.8635
R514 Q0.n0 Q0.t8 27.7543
R515 Q0.n2 Q0.t3 18.1962
R516 Q0.n4 Q0.t6 15.3826
R517 Q0.n11 Q0.n8 7.09905
R518 Q0.n5 Q0.n4 6.86134
R519 Q0.n6 Q0.n3 5.01116
R520 Q0.n7 Q0.n1 3.41795
R521 Q0.n11 Q0.n10 3.25085
R522 Q0.n10 Q0.t2 2.2755
R523 Q0.n10 Q0.n9 2.2755
R524 Q0.n12 Q0.n7 2.2505
R525 Q0.n3 Q0.n2 2.13398
R526 Q0.n1 Q0.n0 1.73738
R527 Q0.n7 Q0.n6 1.50498
R528 Q0.n6 Q0.n5 1.12056
R529 Q0.n12 Q0.n11 0.0919062
R530 Q0.n5 Q0 0.0857632
R531 Q0.n3 Q0 0.0810725
R532 Q0 Q0.n12 0.073625
R533 Q0.n1 Q0 0.0694712
R534 Vdiv3.n2 Vdiv3.n1 9.33985
R535 Vdiv3.n2 Vdiv3.n0 5.17836
R536 Vdiv3 Vdiv3.n2 0.0749828
R537 Q1.n11 Q1.t6 36.935
R538 Q1.n4 Q1.t7 31.528
R539 Q1.n9 Q1.t5 31.528
R540 Q1.n0 Q1.t3 30.5184
R541 Q1.n0 Q1.t8 24.7029
R542 Q1.n11 Q1.t4 18.1962
R543 Q1.n4 Q1.t10 15.3826
R544 Q1.n9 Q1.t9 15.3826
R545 Q1.n8 Q1.n7 7.43416
R546 Q1.n18 Q1.n15 7.09905
R547 Q1.n10 Q1.n9 6.86134
R548 Q1.n5 Q1.n4 5.68456
R549 Q1.n13 Q1.n12 5.01109
R550 Q1.n3 Q1.n2 4.5005
R551 Q1.n5 Q1.n2 4.5005
R552 Q1.n18 Q1.n17 3.25085
R553 Q1.n19 Q1.n14 2.34532
R554 Q1.n17 Q1.t1 2.2755
R555 Q1.n17 Q1.n16 2.2755
R556 Q1.n7 Q1.n6 2.2414
R557 Q1.n12 Q1.n11 2.13398
R558 Q1.n1 Q1.n0 1.81206
R559 Q1.n14 Q1.n13 1.49653
R560 Q1.n14 Q1.n8 1.23718
R561 Q1.n13 Q1.n10 1.12725
R562 Q1.n8 Q1.n1 0.977039
R563 Q1.n1 Q1 0.105733
R564 Q1.n19 Q1.n18 0.0919062
R565 Q1.n10 Q1 0.0857632
R566 Q1.n12 Q1 0.0810725
R567 Q1 Q1.n19 0.073625
R568 Q1.n3 Q1 0.0444655
R569 Q1.n6 Q1.n3 0.028431
R570 Q1.n7 Q1.n2 0.0234177
R571 Q1.n6 Q1.n5 0.0129138
R572 RST.n7 RST.t3 37.1991
R573 RST.n0 RST.t1 36.935
R574 RST.n0 RST.t0 18.1962
R575 RST.n7 RST.t2 17.66
R576 RST.n11 RST.n10 9.41757
R577 RST.n11 RST.n4 4.5005
R578 RST.n13 RST.n12 2.24959
R579 RST.n10 RST.n9 2.24157
R580 RST.n2 RST.n0 2.11961
R581 RST.n8 RST.n7 1.41552
R582 RST RST.n13 0.0592509
R583 RST.n6 RST 0.0410354
R584 RST.n9 RST.n6 0.0361897
R585 RST RST.n11 0.0293
R586 RST.n10 RST.n5 0.0230258
R587 RST.n13 RST.n4 0.0188336
R588 RST.n2 RST.n1 0.00556597
R589 RST.n3 RST.n2 0.00546378
R590 RST.n9 RST.n8 0.00515517
R591 RST.n4 RST.n3 0.00332638
R592 RST.n12 RST 0.0017
C0 JK_FF_mag_0.nand2_mag_1.IN2 CLK 7.81e-19
C1 or_2_mag_0.GF_INV_MAG_1.IN JK_FF_mag_1.J 0.00205f
C2 a_5657_256# JK_FF_mag_1.J 0.0811f
C3 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_4.IN2 0.122f
C4 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_1.IN1 0.765f
C5 a_5060_2688# JK_FF_mag_1.J 0.00168f
C6 CLK a_1358_1353# 6.43e-21
C7 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00166f
C8 a_2076_256# JK_FF_mag_1.nand2_mag_3.IN1 0.0036f
C9 JK_FF_mag_0.nand3_mag_2.OUT a_3645_212# 0.0202f
C10 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.nand2_mag_4.IN2 8.59e-20
C11 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C12 Q0 JK_FF_mag_0.nand2_mag_3.IN1 0.0175f
C13 JK_FF_mag_0.nand2_mag_1.IN2 or_2_mag_0.IN2 3.81e-19
C14 RST JK_FF_mag_0.nand3_mag_1.OUT 0.276f
C15 Vdiv3 Q1 2.53e-19
C16 a_2486_1353# JK_FF_mag_1.nand2_mag_3.IN1 0.00118f
C17 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_3.IN1 0.21f
C18 a_1512_212# JK_FF_mag_1.QB 0.00696f
C19 a_4529_212# JK_FF_mag_0.nand3_mag_1.IN1 8.64e-19
C20 JK_FF_mag_0.nand3_mag_1.IN1 CLK 0.00254f
C21 JK_FF_mag_0.nand2_mag_4.IN2 Q0 0.0635f
C22 a_2076_256# RST 5.68e-19
C23 a_5093_256# JK_FF_mag_1.J 0.00964f
C24 a_1922_1353# JK_FF_mag_1.nand2_mag_3.IN1 0.011f
C25 Q0 VDD 1.26f
C26 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_0.OUT 0.0622f
C27 a_4375_1353# RST 1.9e-19
C28 JK_FF_mag_1.nand3_mag_1.OUT a_788_212# 1.5e-20
C29 or_2_mag_0.GF_INV_MAG_1.IN Q0 0.209f
C30 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.J 9.62e-20
C31 Q1 JK_FF_mag_0.nand3_mag_1.OUT 4.33e-19
C32 Q0 a_5657_256# 0.0157f
C33 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand3_mag_2.OUT 0.00183f
C34 JK_FF_mag_1.nand3_mag_2.OUT a_788_212# 0.0731f
C35 a_2486_1353# RST 7.24e-19
C36 JK_FF_mag_1.QB RST 0.584f
C37 or_2_mag_0.IN2 JK_FF_mag_0.nand3_mag_1.IN1 1.82e-19
C38 a_5060_2688# Q0 0.0134f
C39 JK_FF_mag_1.nand2_mag_1.IN2 JK_FF_mag_1.J 8.58e-20
C40 a_2076_256# Q1 0.00859f
C41 JK_FF_mag_1.nand2_mag_3.IN1 VDD 1f
C42 a_1922_1353# RST 3.62e-19
C43 a_5503_1353# JK_FF_mag_1.J 0.012f
C44 JK_FF_mag_0.nand2_mag_3.IN1 RST 0.00941f
C45 a_1512_212# VDD 9.82e-19
C46 and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_0.nand3_mag_1.IN1 6.02e-20
C47 a_4369_212# JK_FF_mag_0.nand3_mag_2.OUT 9.1e-19
C48 a_2486_1353# Q1 0.069f
C49 JK_FF_mag_1.QB Q1 1.94f
C50 JK_FF_mag_0.nand2_mag_4.IN2 RST 0.00239f
C51 a_5093_256# Q0 0.00859f
C52 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand3_mag_0.OUT 0.122f
C53 RST VDD 0.548f
C54 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.J 8.58e-20
C55 JK_FF_mag_0.nand2_mag_3.IN1 Q1 0.104f
C56 a_4529_212# JK_FF_mag_0.nand3_mag_1.OUT 0.0733f
C57 CLK JK_FF_mag_0.nand3_mag_1.OUT 0.00302f
C58 JK_FF_mag_1.nand3_mag_0.OUT a_794_1309# 0.0732f
C59 a_634_1309# a_794_1309# 0.0504f
C60 Q0 a_5503_1353# 0.069f
C61 Vdiv3 and2_mag_0.GF_INV_MAG_0.IN 1e-19
C62 Q1 VDD 2.49f
C63 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_3.IN1 0.159f
C64 or_2_mag_0.GF_INV_MAG_1.IN Q1 0.00139f
C65 RST a_2640_256# 0.00114f
C66 a_4375_1353# CLK 6.43e-21
C67 a_1512_212# JK_FF_mag_1.nand3_mag_1.OUT 0.0733f
C68 or_2_mag_0.IN2 JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C69 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_2.OUT 0.00169f
C70 a_3645_212# JK_FF_mag_0.nand3_mag_1.OUT 1.17e-20
C71 a_634_1309# JK_FF_mag_1.nand3_mag_0.OUT 0.0203f
C72 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand3_mag_2.OUT 0.00118f
C73 a_1512_212# JK_FF_mag_1.nand3_mag_2.OUT 2.88e-20
C74 a_2486_1353# CLK 9.45e-19
C75 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.J 0.0948f
C76 JK_FF_mag_1.QB CLK 0.362f
C77 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.IN1 0.109f
C78 a_634_1309# JK_FF_mag_1.J 8.64e-19
C79 a_4939_1353# or_2_mag_0.IN2 4.9e-20
C80 a_3805_212# Q0 0.00789f
C81 a_5060_2688# Q1 6.83e-19
C82 a_4087_2452# VDD 5.92e-19
C83 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_1.IN2 0.359f
C84 JK_FF_mag_1.QB a_3811_1309# 1.41e-20
C85 JK_FF_mag_1.J JK_FF_mag_0.nand3_mag_0.OUT 0.352f
C86 and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_0.nand3_mag_1.OUT 6.11e-19
C87 a_1922_1353# CLK 6.06e-21
C88 JK_FF_mag_1.nand3_mag_1.OUT RST 0.311f
C89 JK_FF_mag_0.nand2_mag_3.IN1 CLK 0.471f
C90 Q1 a_2640_256# 0.0157f
C91 JK_FF_mag_0.nand2_mag_3.IN1 a_3811_1309# 0.00119f
C92 JK_FF_mag_1.QB a_3651_1309# 1.86e-20
C93 a_628_212# VDD 0.0132f
C94 RST JK_FF_mag_1.nand3_mag_2.OUT 0.0545f
C95 RST JK_FF_mag_1.nand2_mag_1.IN2 6.71e-19
C96 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.nand2_mag_4.IN2 0.313f
C97 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.nand2_mag_3.IN1 0.231f
C98 CLK VDD 2.37f
C99 a_1512_212# JK_FF_mag_1.nand3_mag_1.IN1 8.64e-19
C100 or_2_mag_0.IN2 JK_FF_mag_0.nand2_mag_3.IN1 5.32e-19
C101 JK_FF_mag_1.nand3_mag_1.OUT Q1 0.0343f
C102 or_2_mag_0.GF_INV_MAG_1.IN CLK 7.03e-21
C103 Q1 JK_FF_mag_1.nand3_mag_2.OUT 0.338f
C104 JK_FF_mag_1.nand2_mag_3.IN1 a_794_1309# 0.00119f
C105 and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_0.nand2_mag_3.IN1 3.67e-20
C106 a_3651_1309# VDD 2.21e-19
C107 a_3805_212# RST 0.00218f
C108 Q1 JK_FF_mag_1.nand2_mag_1.IN2 0.109f
C109 Q0 JK_FF_mag_0.nand3_mag_0.OUT 7.24e-19
C110 Q0 JK_FF_mag_1.J 2.37f
C111 a_4369_212# JK_FF_mag_0.nand3_mag_1.OUT 0.0203f
C112 RST JK_FF_mag_1.nand2_mag_4.IN2 0.0562f
C113 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.121f
C114 or_2_mag_0.IN2 VDD 0.49f
C115 JK_FF_mag_1.nand3_mag_1.IN1 RST 0.193f
C116 VDD a_3645_212# 0.00743f
C117 or_2_mag_0.GF_INV_MAG_1.IN or_2_mag_0.IN2 0.0445f
C118 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.00975f
C119 and2_mag_0.GF_INV_MAG_0.IN VDD 0.465f
C120 JK_FF_mag_1.nand3_mag_0.OUT JK_FF_mag_1.nand2_mag_3.IN1 0.0854f
C121 a_628_212# JK_FF_mag_1.nand3_mag_1.OUT 1.17e-20
C122 JK_FF_mag_1.nand2_mag_3.IN1 a_788_212# 1.46e-19
C123 a_3805_212# Q1 1.86e-20
C124 JK_FF_mag_0.nand2_mag_1.IN2 a_4939_1353# 0.069f
C125 a_5060_2688# or_2_mag_0.IN2 8.64e-19
C126 or_2_mag_0.GF_INV_MAG_1.IN and2_mag_0.GF_INV_MAG_0.IN 3.34e-19
C127 JK_FF_mag_1.nand2_mag_3.IN1 JK_FF_mag_1.J 0.0718f
C128 a_628_212# JK_FF_mag_1.nand3_mag_2.OUT 0.0202f
C129 Q1 JK_FF_mag_1.nand2_mag_4.IN2 0.0636f
C130 JK_FF_mag_1.nand3_mag_1.IN1 Q1 0.00335f
C131 a_5060_2688# and2_mag_0.GF_INV_MAG_0.IN 3.25e-19
C132 JK_FF_mag_1.nand3_mag_1.OUT CLK 0.00481f
C133 CLK JK_FF_mag_1.nand3_mag_2.OUT 0.235f
C134 Q1 a_794_1309# 2.79e-20
C135 RST JK_FF_mag_1.J 0.249f
C136 RST JK_FF_mag_0.nand3_mag_0.OUT 0.00412f
C137 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_1.OUT 0.768f
C138 JK_FF_mag_1.nand2_mag_1.IN2 CLK 0.0215f
C139 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_2.OUT 9.52e-19
C140 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.36f
C141 JK_FF_mag_1.QB a_1358_1353# 3.33e-19
C142 a_4939_1353# JK_FF_mag_0.nand3_mag_1.IN1 0.0059f
C143 a_4369_212# VDD 2.21e-19
C144 JK_FF_mag_1.nand3_mag_0.OUT Q1 7.24e-19
C145 a_4375_1353# JK_FF_mag_0.nand3_mag_1.IN1 0.0697f
C146 Q1 a_788_212# 0.00789f
C147 JK_FF_mag_0.nand3_mag_2.OUT VDD 0.739f
C148 a_3805_212# CLK 0.00164f
C149 Q1 JK_FF_mag_1.J 0.363f
C150 Q1 JK_FF_mag_0.nand3_mag_0.OUT 0.101f
C151 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_1.IN2 8.16e-20
C152 CLK JK_FF_mag_1.nand2_mag_4.IN2 5.57e-19
C153 JK_FF_mag_0.nand2_mag_1.IN2 VDD 0.398f
C154 JK_FF_mag_1.nand3_mag_1.IN1 CLK 0.013f
C155 JK_FF_mag_1.QB a_1352_212# 0.00695f
C156 or_2_mag_0.GF_INV_MAG_1.IN JK_FF_mag_0.nand2_mag_1.IN2 1.53e-19
C157 VDD a_1358_1353# 3.14e-19
C158 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand2_mag_3.IN1 0.233f
C159 Q0 RST 0.0447f
C160 CLK a_794_1309# 0.00939f
C161 a_3805_212# a_3645_212# 0.0504f
C162 a_628_212# a_788_212# 0.0504f
C163 JK_FF_mag_0.nand3_mag_1.IN1 VDD 0.652f
C164 a_1352_212# VDD 0.0012f
C165 JK_FF_mag_1.nand3_mag_0.OUT CLK 0.298f
C166 RST JK_FF_mag_1.nand2_mag_3.IN1 0.13f
C167 a_634_1309# CLK 0.0101f
C168 Q0 Q1 0.0285f
C169 CLK a_788_212# 0.00164f
C170 a_4939_1353# JK_FF_mag_0.nand3_mag_1.OUT 4.52e-20
C171 a_1512_212# RST 0.00135f
C172 a_4529_212# JK_FF_mag_1.J 0.00696f
C173 CLK JK_FF_mag_1.J 2.09f
C174 CLK JK_FF_mag_0.nand3_mag_0.OUT 0.272f
C175 a_3811_1309# JK_FF_mag_0.nand3_mag_0.OUT 0.0732f
C176 a_3811_1309# JK_FF_mag_1.J 0.00392f
C177 a_4375_1353# JK_FF_mag_0.nand3_mag_1.OUT 0.0202f
C178 a_3651_1309# JK_FF_mag_0.nand3_mag_0.OUT 0.0203f
C179 Q1 JK_FF_mag_1.nand2_mag_3.IN1 0.0177f
C180 JK_FF_mag_1.nand3_mag_1.OUT a_1358_1353# 0.0202f
C181 or_2_mag_0.IN2 JK_FF_mag_1.J 0.00761f
C182 a_1512_212# Q1 0.0101f
C183 JK_FF_mag_0.nand2_mag_1.IN2 a_5503_1353# 0.00372f
C184 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_1.OUT 0.16f
C185 and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_1.J 0.00384f
C186 and2_mag_0.GF_INV_MAG_0.IN JK_FF_mag_0.nand3_mag_0.OUT 2.34e-19
C187 a_2076_256# JK_FF_mag_1.QB 0.00964f
C188 Vdiv3 VDD 0.152f
C189 a_3805_212# JK_FF_mag_0.nand3_mag_2.OUT 0.0731f
C190 or_2_mag_0.GF_INV_MAG_1.IN Vdiv3 0.126f
C191 a_4939_1353# JK_FF_mag_0.nand2_mag_3.IN1 0.011f
C192 Q1 RST 0.0659f
C193 a_4529_212# Q0 0.0101f
C194 Q0 CLK 0.149f
C195 JK_FF_mag_1.nand3_mag_1.OUT a_1352_212# 0.0203f
C196 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand3_mag_1.OUT 0.122f
C197 Q0 a_3811_1309# 2.79e-20
C198 a_2486_1353# JK_FF_mag_1.QB 0.0112f
C199 JK_FF_mag_1.nand3_mag_2.OUT a_1352_212# 9.1e-19
C200 a_4375_1353# JK_FF_mag_0.nand2_mag_3.IN1 1.43e-19
C201 VDD JK_FF_mag_0.nand3_mag_1.OUT 0.995f
C202 a_4939_1353# VDD 3.14e-19
C203 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_1.QB 7.08e-20
C204 JK_FF_mag_1.nand3_mag_1.IN1 a_1358_1353# 0.0697f
C205 a_2076_256# VDD 0.00149f
C206 Q0 or_2_mag_0.IN2 0.0655f
C207 JK_FF_mag_1.nand2_mag_3.IN1 CLK 1.29f
C208 Q0 a_3645_212# 0.00335f
C209 a_4375_1353# VDD 3.14e-19
C210 Q0 and2_mag_0.GF_INV_MAG_0.IN 8.04e-19
C211 a_4369_212# JK_FF_mag_1.J 0.00695f
C212 a_2486_1353# VDD 3.56e-19
C213 a_4087_2452# Q1 0.01f
C214 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_1.J 0.0881f
C215 JK_FF_mag_0.nand3_mag_2.OUT JK_FF_mag_0.nand3_mag_0.OUT 0.00183f
C216 JK_FF_mag_1.QB VDD 0.875f
C217 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_0.nand2_mag_3.IN1 0.321f
C218 a_4529_212# RST 0.00103f
C219 RST CLK 0.03f
C220 JK_FF_mag_0.nand2_mag_1.IN2 JK_FF_mag_1.J 0.0725f
C221 RST a_3811_1309# 6.43e-19
C222 a_1922_1353# VDD 3.14e-19
C223 a_5093_256# JK_FF_mag_0.nand3_mag_1.OUT 0.00378f
C224 JK_FF_mag_0.nand2_mag_3.IN1 VDD 1.08f
C225 JK_FF_mag_1.nand3_mag_0.OUT a_1358_1353# 0.00378f
C226 a_628_212# Q1 0.00335f
C227 or_2_mag_0.GF_INV_MAG_1.IN JK_FF_mag_0.nand2_mag_3.IN1 1.99e-19
C228 RST a_3651_1309# 7.78e-19
C229 JK_FF_mag_0.nand2_mag_4.IN2 VDD 0.391f
C230 JK_FF_mag_1.QB a_2640_256# 0.0811f
C231 a_5060_2688# JK_FF_mag_0.nand2_mag_3.IN1 1.4e-19
C232 or_2_mag_0.GF_INV_MAG_1.IN JK_FF_mag_0.nand2_mag_4.IN2 4.44e-20
C233 Q1 CLK 1.03f
C234 RST a_3645_212# 0.00218f
C235 a_2076_256# JK_FF_mag_1.nand3_mag_1.OUT 0.00378f
C236 JK_FF_mag_0.nand2_mag_4.IN2 a_5657_256# 0.00372f
C237 or_2_mag_0.GF_INV_MAG_1.IN VDD 0.412f
C238 a_5657_256# VDD 3.14e-19
C239 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_1.J 0.0435f
C240 JK_FF_mag_0.nand3_mag_1.IN1 JK_FF_mag_0.nand3_mag_0.OUT 0.122f
C241 a_4369_212# Q0 0.0102f
C242 Q1 a_3651_1309# 0.00149f
C243 Q0 JK_FF_mag_0.nand3_mag_2.OUT 0.338f
C244 a_4087_2452# CLK 0.0103f
C245 a_5060_2688# VDD 0.165f
C246 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.QB 0.215f
C247 JK_FF_mag_0.nand2_mag_1.IN2 Q0 0.107f
C248 or_2_mag_0.IN2 Q1 0.0138f
C249 a_5060_2688# or_2_mag_0.GF_INV_MAG_1.IN 0.132f
C250 a_5093_256# JK_FF_mag_0.nand2_mag_3.IN1 0.0036f
C251 Q1 a_3645_212# 2.55e-20
C252 a_3805_212# JK_FF_mag_0.nand3_mag_1.OUT 1.5e-20
C253 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_2.OUT 0.103f
C254 a_1922_1353# JK_FF_mag_1.nand3_mag_1.OUT 4.52e-20
C255 VDD a_2640_256# 0.00149f
C256 a_2486_1353# JK_FF_mag_1.nand2_mag_1.IN2 0.00372f
C257 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_1.IN2 0.0576f
C258 and2_mag_0.GF_INV_MAG_0.IN Q1 0.305f
C259 a_628_212# CLK 0.00117f
C260 a_5093_256# JK_FF_mag_0.nand2_mag_4.IN2 0.069f
C261 a_4087_2452# or_2_mag_0.IN2 7.48e-20
C262 a_1922_1353# JK_FF_mag_1.nand2_mag_1.IN2 0.069f
C263 a_5093_256# VDD 3.14e-19
C264 a_2076_256# JK_FF_mag_1.nand2_mag_4.IN2 0.069f
C265 a_3811_1309# CLK 0.00939f
C266 a_4087_2452# and2_mag_0.GF_INV_MAG_0.IN 0.069f
C267 JK_FF_mag_0.nand2_mag_3.IN1 a_5503_1353# 0.00118f
C268 JK_FF_mag_1.nand3_mag_1.OUT VDD 0.999f
C269 Vdiv3 JK_FF_mag_1.J 4.46e-19
C270 Q0 JK_FF_mag_0.nand3_mag_1.IN1 0.00335f
C271 JK_FF_mag_1.nand2_mag_3.IN1 a_1358_1353# 1.43e-19
C272 a_4369_212# RST 0.00119f
C273 JK_FF_mag_1.nand3_mag_2.OUT VDD 0.802f
C274 a_2486_1353# JK_FF_mag_1.nand2_mag_4.IN2 4.52e-20
C275 a_3651_1309# CLK 0.0101f
C276 RST JK_FF_mag_0.nand3_mag_2.OUT 0.0981f
C277 JK_FF_mag_1.QB JK_FF_mag_1.nand2_mag_4.IN2 0.175f
C278 JK_FF_mag_1.nand3_mag_1.IN1 JK_FF_mag_1.QB 0.0147f
C279 a_3651_1309# a_3811_1309# 0.0504f
C280 JK_FF_mag_0.nand2_mag_4.IN2 a_5503_1353# 4.52e-20
C281 JK_FF_mag_1.nand2_mag_1.IN2 VDD 0.397f
C282 a_3805_212# JK_FF_mag_0.nand2_mag_3.IN1 1.46e-19
C283 or_2_mag_0.IN2 CLK 6.62e-20
C284 a_5503_1353# VDD 3.56e-19
C285 JK_FF_mag_1.J JK_FF_mag_0.nand3_mag_1.OUT 0.23f
C286 JK_FF_mag_0.nand3_mag_0.OUT JK_FF_mag_0.nand3_mag_1.OUT 0.0622f
C287 CLK a_3645_212# 0.00117f
C288 a_1922_1353# JK_FF_mag_1.nand3_mag_1.IN1 0.0059f
C289 or_2_mag_0.GF_INV_MAG_1.IN a_5503_1353# 4.94e-20
C290 JK_FF_mag_1.QB a_794_1309# 0.00392f
C291 a_4939_1353# JK_FF_mag_1.J 2.96e-19
C292 a_4369_212# Q1 3.6e-22
C293 and2_mag_0.GF_INV_MAG_0.IN CLK 0.0983f
C294 a_1512_212# a_1352_212# 0.0504f
C295 Q1 JK_FF_mag_0.nand3_mag_2.OUT 9.98e-19
C296 a_3805_212# VDD 0.00305f
C297 JK_FF_mag_0.nand2_mag_1.IN2 Q1 1.12e-19
C298 a_4375_1353# JK_FF_mag_0.nand3_mag_0.OUT 0.00378f
C299 a_4375_1353# JK_FF_mag_1.J 1.75e-19
C300 JK_FF_mag_1.nand2_mag_4.IN2 VDD 0.394f
C301 JK_FF_mag_1.nand3_mag_1.IN1 VDD 0.652f
C302 JK_FF_mag_1.QB JK_FF_mag_1.nand3_mag_0.OUT 0.343f
C303 Q0 Vdiv3 0.0076f
C304 JK_FF_mag_0.nand3_mag_1.IN1 RST 0.143f
C305 JK_FF_mag_1.QB JK_FF_mag_0.nand3_mag_0.OUT 2.81e-20
C306 JK_FF_mag_1.QB JK_FF_mag_1.J 3.28e-19
C307 and2_mag_0.GF_INV_MAG_0.IN or_2_mag_0.IN2 0.124f
C308 RST a_1352_212# 8.64e-19
C309 VDD a_794_1309# 2.65e-19
C310 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand3_mag_2.OUT 0.121f
C311 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_0.nand3_mag_0.OUT 0.0894f
C312 JK_FF_mag_0.nand2_mag_3.IN1 JK_FF_mag_1.J 0.69f
C313 JK_FF_mag_1.nand3_mag_1.OUT JK_FF_mag_1.nand2_mag_1.IN2 0.00975f
C314 Q0 JK_FF_mag_0.nand3_mag_1.OUT 0.0343f
C315 JK_FF_mag_1.nand2_mag_4.IN2 a_2640_256# 0.00372f
C316 JK_FF_mag_0.nand3_mag_1.IN1 Q1 6.7e-19
C317 Q1 a_1352_212# 0.0102f
C318 JK_FF_mag_0.nand2_mag_4.IN2 JK_FF_mag_1.J 0.198f
C319 a_4529_212# a_4369_212# 0.0504f
C320 JK_FF_mag_1.nand3_mag_0.OUT VDD 0.647f
C321 a_4529_212# JK_FF_mag_0.nand3_mag_2.OUT 2.88e-20
C322 CLK JK_FF_mag_0.nand3_mag_2.OUT 0.235f
C323 a_634_1309# VDD 5.99e-19
C324 a_788_212# VDD 0.00888f
C325 VDD JK_FF_mag_1.J 2.22f
C326 VDD JK_FF_mag_0.nand3_mag_0.OUT 0.647f
C327 a_5657_256# VSS 0.0675f
C328 a_5093_256# VSS 0.0676f
C329 a_4529_212# VSS 0.0343f
C330 a_4369_212# VSS 0.0881f
C331 a_3805_212# VSS 0.0343f
C332 a_3645_212# VSS 0.0881f
C333 a_2640_256# VSS 0.0675f
C334 a_2076_256# VSS 0.0676f
C335 a_1512_212# VSS 0.0343f
C336 a_1352_212# VSS 0.0881f
C337 a_788_212# VSS 0.0343f
C338 a_628_212# VSS 0.0881f
C339 JK_FF_mag_0.nand2_mag_4.IN2 VSS 0.415f
C340 JK_FF_mag_0.nand3_mag_2.OUT VSS 0.539f
C341 JK_FF_mag_1.nand2_mag_4.IN2 VSS 0.416f
C342 RST VSS 0.9f
C343 JK_FF_mag_1.nand3_mag_2.OUT VSS 0.519f
C344 a_5503_1353# VSS 0.0676f
C345 a_4939_1353# VSS 0.0676f
C346 a_4375_1353# VSS 0.0676f
C347 a_3811_1309# VSS 0.0343f
C348 a_3651_1309# VSS 0.0881f
C349 a_2486_1353# VSS 0.0676f
C350 a_1922_1353# VSS 0.0676f
C351 a_1358_1353# VSS 0.0676f
C352 a_794_1309# VSS 0.0343f
C353 a_634_1309# VSS 0.0881f
C354 JK_FF_mag_0.nand2_mag_1.IN2 VSS 0.415f
C355 JK_FF_mag_0.nand2_mag_3.IN1 VSS 0.69f
C356 JK_FF_mag_0.nand3_mag_1.IN1 VSS 0.724f
C357 JK_FF_mag_0.nand3_mag_1.OUT VSS 0.809f
C358 JK_FF_mag_0.nand3_mag_0.OUT VSS 0.509f
C359 JK_FF_mag_1.nand2_mag_1.IN2 VSS 0.415f
C360 JK_FF_mag_1.nand2_mag_3.IN1 VSS 0.708f
C361 JK_FF_mag_1.nand3_mag_1.IN1 VSS 0.724f
C362 JK_FF_mag_1.nand3_mag_1.OUT VSS 0.809f
C363 JK_FF_mag_1.nand3_mag_0.OUT VSS 0.509f
C364 JK_FF_mag_1.QB VSS 0.859f
C365 JK_FF_mag_1.J VSS 4.65f
C366 a_4087_2452# VSS 0.0676f
C367 Vdiv3 VSS 0.176f
C368 or_2_mag_0.GF_INV_MAG_1.IN VSS 0.6f
C369 a_5060_2688# VSS 0.0247f
C370 Q0 VSS 2.03f
C371 or_2_mag_0.IN2 VSS 0.418f
C372 and2_mag_0.GF_INV_MAG_0.IN VSS 0.435f
C373 Q1 VSS 1.84f
C374 CLK VSS 2.46f
C375 VDD VSS 33.9f
C376 Q1.t8 VSS 0.0273f
C377 Q1.t3 VSS 0.0352f
C378 Q1.n0 VSS 0.0697f
C379 Q1.n1 VSS 0.0272f
C380 Q1.n2 VSS 0.0111f
C381 Q1.n3 VSS 0.00546f
C382 Q1.t10 VSS 0.0218f
C383 Q1.t7 VSS 0.0274f
C384 Q1.n4 VSS 0.0616f
C385 Q1.n5 VSS 0.0274f
C386 Q1.n6 VSS 0.0031f
C387 Q1.n7 VSS 0.336f
C388 Q1.n8 VSS 0.272f
C389 Q1.t9 VSS 0.0218f
C390 Q1.t5 VSS 0.0274f
C391 Q1.n9 VSS 0.0633f
C392 Q1.n10 VSS 0.0395f
C393 Q1.t4 VSS 0.0251f
C394 Q1.t6 VSS 0.0381f
C395 Q1.n11 VSS 0.0676f
C396 Q1.n12 VSS 0.265f
C397 Q1.n13 VSS 0.496f
C398 Q1.n14 VSS 0.21f
C399 Q1.n15 VSS 0.0207f
C400 Q1.t1 VSS 0.0171f
C401 Q1.n16 VSS 0.0171f
C402 Q1.n17 VSS 0.0469f
C403 Q1.n18 VSS 0.151f
C404 Q1.n19 VSS 0.0157f
C405 Q0.t4 VSS 0.0632f
C406 Q0.t8 VSS 0.0195f
C407 Q0.n0 VSS 0.0665f
C408 Q0.n1 VSS 0.197f
C409 Q0.t3 VSS 0.0298f
C410 Q0.t5 VSS 0.0452f
C411 Q0.n2 VSS 0.0802f
C412 Q0.n3 VSS 0.314f
C413 Q0.t6 VSS 0.0259f
C414 Q0.t7 VSS 0.0325f
C415 Q0.n4 VSS 0.0752f
C416 Q0.n5 VSS 0.0467f
C417 Q0.n6 VSS 0.597f
C418 Q0.n7 VSS 0.441f
C419 Q0.n8 VSS 0.0246f
C420 Q0.t2 VSS 0.0203f
C421 Q0.n9 VSS 0.0203f
C422 Q0.n10 VSS 0.0557f
C423 Q0.n11 VSS 0.18f
C424 Q0.n12 VSS 0.0182f
C425 JK_FF_mag_1.J.n0 VSS 2.03f
C426 JK_FF_mag_1.J.n1 VSS 0.196f
C427 JK_FF_mag_1.J.t7 VSS 0.0683f
C428 JK_FF_mag_1.J.t5 VSS 0.053f
C429 JK_FF_mag_1.J.n2 VSS 0.135f
C430 JK_FF_mag_1.J.t8 VSS 0.0424f
C431 JK_FF_mag_1.J.t3 VSS 0.0531f
C432 JK_FF_mag_1.J.n3 VSS 0.137f
C433 JK_FF_mag_1.J.t4 VSS 0.0745f
C434 JK_FF_mag_1.J.t6 VSS 0.0475f
C435 JK_FF_mag_1.J.n4 VSS 0.132f
C436 JK_FF_mag_1.J.n5 VSS 1.13f
C437 JK_FF_mag_1.J.t2 VSS 0.0332f
C438 JK_FF_mag_1.J.n6 VSS 0.0332f
C439 JK_FF_mag_1.J.n7 VSS 0.0782f
C440 CLK.n0 VSS 0.00561f
C441 CLK.n1 VSS 0.0046f
C442 CLK.n2 VSS 0.00921f
C443 CLK.t13 VSS 0.0366f
C444 CLK.t2 VSS 0.0555f
C445 CLK.n3 VSS 0.0981f
C446 CLK.n4 VSS 0.0126f
C447 CLK.n5 VSS 0.0179f
C448 CLK.n6 VSS 0.181f
C449 CLK.n7 VSS 0.184f
C450 CLK.n8 VSS 0.00921f
C451 CLK.t3 VSS 0.0366f
C452 CLK.t0 VSS 0.0555f
C453 CLK.n9 VSS 0.0981f
C454 CLK.n10 VSS 0.0126f
C455 CLK.n11 VSS 0.00455f
C456 CLK.n12 VSS 0.106f
C457 CLK.t12 VSS 0.0515f
C458 CLK.t5 VSS 0.0287f
C459 CLK.n13 VSS 0.098f
C460 CLK.n14 VSS 0.314f
C461 CLK.n15 VSS 0.0046f
C462 CLK.n16 VSS 0.00921f
C463 CLK.t8 VSS 0.0366f
C464 CLK.t9 VSS 0.0555f
C465 CLK.n17 VSS 0.0981f
C466 CLK.n18 VSS 0.0126f
C467 CLK.n19 VSS 0.0179f
C468 CLK.n20 VSS 0.169f
C469 CLK.n21 VSS 0.381f
C470 CLK.n22 VSS 0.0142f
C471 CLK.n23 VSS 0.00921f
C472 CLK.t10 VSS 0.0366f
C473 CLK.t7 VSS 0.0555f
C474 CLK.n24 VSS 0.0981f
C475 CLK.n25 VSS 0.0126f
C476 CLK.n26 VSS 0.00455f
C477 CLK.n27 VSS 0.106f
C478 CLK.n28 VSS 0.0193f
C479 CLK.t1 VSS 0.0459f
C480 CLK.t4 VSS 0.0117f
C481 CLK.n29 VSS 0.0759f
C482 CLK.n30 VSS 0.0161f
C483 CLK.n31 VSS 0.033f
C484 CLK.n32 VSS 0.00561f
C485 CLK.n33 VSS 0.0122f
C486 CLK.n34 VSS 0.702f
C487 CLK.n35 VSS 0.702f
C488 CLK.n36 VSS 0.0122f
C489 CLK.t6 VSS 0.0459f
C490 CLK.t11 VSS 0.0117f
C491 CLK.n37 VSS 0.0759f
C492 CLK.n38 VSS 0.0161f
C493 CLK.n39 VSS 0.0193f
C494 CLK.n40 VSS 0.0155f
C495 VDD.t22 VSS 0.00641f
C496 VDD.n0 VSS 0.0064f
C497 VDD.n1 VSS 0.0315f
C498 VDD.t58 VSS 0.00638f
C499 VDD.n2 VSS 0.0226f
C500 VDD.t57 VSS 0.0576f
C501 VDD.t109 VSS 0.0573f
C502 VDD.t1 VSS 0.00638f
C503 VDD.t0 VSS 0.0568f
C504 VDD.n3 VSS 0.0658f
C505 VDD.n4 VSS 0.0343f
C506 VDD.t11 VSS 0.0153f
C507 VDD.n5 VSS 0.0347f
C508 VDD.n6 VSS 0.0341f
C509 VDD.n7 VSS 0.0387f
C510 VDD.t10 VSS 0.0545f
C511 VDD.n8 VSS 0.0998f
C512 VDD.t38 VSS 0.0505f
C513 VDD.t21 VSS 0.077f
C514 VDD.n9 VSS 0.0398f
C515 VDD.n10 VSS 0.0224f
C516 VDD.n11 VSS 0.044f
C517 VDD.n12 VSS 0.0499f
C518 VDD.t74 VSS 0.0846f
C519 VDD.n13 VSS 0.0064f
C520 VDD.t46 VSS 0.00641f
C521 VDD.n14 VSS 0.0064f
C522 VDD.n15 VSS 0.0317f
C523 VDD.t71 VSS 0.0834f
C524 VDD.n16 VSS 0.0064f
C525 VDD.n17 VSS 0.0064f
C526 VDD.t97 VSS 0.0834f
C527 VDD.n18 VSS 0.0398f
C528 VDD.t84 VSS 0.00641f
C529 VDD.n19 VSS 0.0064f
C530 VDD.t83 VSS 0.0772f
C531 VDD.t28 VSS 0.0846f
C532 VDD.n20 VSS 0.0398f
C533 VDD.t78 VSS 0.00641f
C534 VDD.t44 VSS 0.00263f
C535 VDD.n21 VSS 0.00263f
C536 VDD.n22 VSS 0.00575f
C537 VDD.t77 VSS 0.0772f
C538 VDD.t43 VSS 0.0943f
C539 VDD.t106 VSS 0.0438f
C540 VDD.n23 VSS 0.0398f
C541 VDD.t37 VSS 0.00641f
C542 VDD.t5 VSS 0.00263f
C543 VDD.n24 VSS 0.00263f
C544 VDD.n25 VSS 0.00575f
C545 VDD.t36 VSS 0.0772f
C546 VDD.t4 VSS 0.0943f
C547 VDD.t49 VSS 0.0438f
C548 VDD.t66 VSS 0.077f
C549 VDD.n26 VSS 0.0398f
C550 VDD.t67 VSS 0.00687f
C551 VDD.n27 VSS 0.0493f
C552 VDD.n28 VSS 0.0365f
C553 VDD.n29 VSS 0.0375f
C554 VDD.n30 VSS 0.0199f
C555 VDD.n31 VSS 0.0365f
C556 VDD.n32 VSS 0.0374f
C557 VDD.n33 VSS 0.0221f
C558 VDD.n34 VSS 0.0317f
C559 VDD.n35 VSS 0.0295f
C560 VDD.n36 VSS 0.0221f
C561 VDD.n37 VSS 0.0604f
C562 VDD.n38 VSS 0.0687f
C563 VDD.t3 VSS 0.00641f
C564 VDD.n39 VSS 0.0295f
C565 VDD.n40 VSS 0.0221f
C566 VDD.n41 VSS 0.0398f
C567 VDD.t2 VSS 0.0772f
C568 VDD.t31 VSS 0.0846f
C569 VDD.t45 VSS 0.0772f
C570 VDD.n42 VSS 0.0398f
C571 VDD.n43 VSS 0.0221f
C572 VDD.n44 VSS 0.0295f
C573 VDD.n45 VSS 0.0317f
C574 VDD.t35 VSS 0.00641f
C575 VDD.t82 VSS 0.00263f
C576 VDD.n46 VSS 0.00263f
C577 VDD.n47 VSS 0.00575f
C578 VDD.n48 VSS 0.0207f
C579 VDD.n49 VSS 0.0279f
C580 VDD.n50 VSS 0.0221f
C581 VDD.n51 VSS 0.0398f
C582 VDD.t34 VSS 0.0772f
C583 VDD.t81 VSS 0.0943f
C584 VDD.t68 VSS 0.0438f
C585 VDD.t27 VSS 0.00641f
C586 VDD.n52 VSS 0.0282f
C587 VDD.t105 VSS 0.00638f
C588 VDD.n53 VSS 0.0064f
C589 VDD.t52 VSS 0.0673f
C590 VDD.n54 VSS 0.0343f
C591 VDD.t80 VSS 0.00641f
C592 VDD.n55 VSS 0.0064f
C593 VDD.t79 VSS 0.0614f
C594 VDD.t18 VSS 0.0673f
C595 VDD.n56 VSS 0.0343f
C596 VDD.t9 VSS 0.00641f
C597 VDD.n57 VSS 0.0064f
C598 VDD.n58 VSS 0.0343f
C599 VDD.t42 VSS 0.00641f
C600 VDD.t56 VSS 0.00263f
C601 VDD.n59 VSS 0.00263f
C602 VDD.n60 VSS 0.00575f
C603 VDD.t41 VSS 0.0614f
C604 VDD.t55 VSS 0.075f
C605 VDD.t94 VSS 0.0348f
C606 VDD.n61 VSS 0.0343f
C607 VDD.t103 VSS 0.00641f
C608 VDD.t8 VSS 0.0455f
C609 VDD.t89 VSS 0.0295f
C610 VDD.n62 VSS 0.178f
C611 VDD.t102 VSS 0.0348f
C612 VDD.n63 VSS 0.0981f
C613 VDD.t47 VSS 0.0706f
C614 VDD.t48 VSS 0.00669f
C615 VDD.n64 VSS 0.0302f
C616 VDD.n65 VSS 0.0199f
C617 VDD.n66 VSS 0.0262f
C618 VDD.n67 VSS 0.0279f
C619 VDD.n68 VSS 0.0221f
C620 VDD.n69 VSS 0.0317f
C621 VDD.n70 VSS 0.0295f
C622 VDD.n71 VSS 0.0221f
C623 VDD.n72 VSS 0.0317f
C624 VDD.n73 VSS 0.0295f
C625 VDD.n74 VSS 0.0221f
C626 VDD.n75 VSS 0.0325f
C627 VDD.n76 VSS 0.0064f
C628 VDD.t59 VSS 0.0834f
C629 VDD.n77 VSS 0.0398f
C630 VDD.t93 VSS 0.00641f
C631 VDD.n78 VSS 0.0064f
C632 VDD.t92 VSS 0.0772f
C633 VDD.t15 VSS 0.0846f
C634 VDD.n79 VSS 0.0398f
C635 VDD.t88 VSS 0.00641f
C636 VDD.t7 VSS 0.00263f
C637 VDD.n80 VSS 0.00263f
C638 VDD.n81 VSS 0.00575f
C639 VDD.t87 VSS 0.0772f
C640 VDD.t6 VSS 0.0943f
C641 VDD.t23 VSS 0.0438f
C642 VDD.n82 VSS 0.0398f
C643 VDD.t86 VSS 0.00641f
C644 VDD.t101 VSS 0.00263f
C645 VDD.n83 VSS 0.00263f
C646 VDD.n84 VSS 0.00575f
C647 VDD.t85 VSS 0.0772f
C648 VDD.t100 VSS 0.0943f
C649 VDD.t12 VSS 0.0438f
C650 VDD.t63 VSS 0.077f
C651 VDD.n85 VSS 0.0398f
C652 VDD.t64 VSS 0.00599f
C653 VDD.n86 VSS 0.00165f
C654 VDD.t62 VSS 0.00534f
C655 VDD.n87 VSS 0.00527f
C656 VDD.t65 VSS 0.0055f
C657 VDD.t110 VSS 0.00417f
C658 VDD.n88 VSS 0.0107f
C659 VDD.n89 VSS 0.0602f
C660 VDD.n90 VSS 0.0787f
C661 VDD.n91 VSS 5.32e-20
C662 VDD.n92 VSS 0.0014f
C663 VDD.t111 VSS 0.00415f
C664 VDD.n93 VSS 0.00563f
C665 VDD.n94 VSS 7.62e-19
C666 VDD.n95 VSS 0.00478f
C667 VDD.n96 VSS 0.0149f
C668 VDD.n97 VSS 0.0366f
C669 VDD.n98 VSS 0.0365f
C670 VDD.n99 VSS 0.0375f
C671 VDD.n100 VSS 0.0199f
C672 VDD.n101 VSS 0.0365f
C673 VDD.n102 VSS 0.0374f
C674 VDD.n103 VSS 0.0221f
C675 VDD.n104 VSS 0.0317f
C676 VDD.n105 VSS 0.0295f
C677 VDD.n106 VSS 0.0221f
C678 VDD.n107 VSS 0.0567f
C679 VDD.n108 VSS 0.0453f
C680 VDD.n109 VSS 0.0201f
C681 VDD.t104 VSS 0.0565f
C682 VDD.n110 VSS 0.0595f
C683 VDD.t26 VSS 0.0438f
C684 VDD.n111 VSS 0.0398f
C685 VDD.n112 VSS 0.0147f
.ends

