magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1045 -1019 1045 1019
<< metal2 >>
rect -45 14 45 19
rect -45 -14 -40 14
rect 40 -14 45 14
rect -45 -19 45 -14
<< via2 >>
rect -40 -14 40 14
<< metal3 >>
rect -45 14 45 19
rect -45 -14 -40 14
rect 40 -14 45 14
rect -45 -19 45 -14
<< end >>
