* NGSPICE file created from or_2_mag_flat.ext - technology: gf180mcuC

.subckt or_2_mag_flat VDD IN2 IN1 OUT VSS
X0 OUT GF_INV_MAG_1.IN VDD.t1 VDD.t0 pfet_03v3 ad=0.352p pd=2.48u as=0.352p ps=2.48u w=0.8u l=0.28u
X1 a_560_998# IN2.t0 VDD.t3 VDD.t2 pfet_03v3 ad=0.416p pd=2.12u as=0.704p ps=4.08u w=1.6u l=0.28u
X2 OUT GF_INV_MAG_1.IN VSS.t6 VSS.t5 nfet_03v3 ad=0.152p pd=1.64u as=0.152p ps=1.64u w=0.22u l=0.28u
X3 GF_INV_MAG_1.IN IN1.t0 a_560_998# VDD.t4 pfet_03v3 ad=0.704p pd=4.08u as=0.416p ps=2.12u w=1.6u l=0.28u
X4 GF_INV_MAG_1.IN IN2.t1 VSS.t4 VSS.t3 nfet_03v3 ad=86.8f pd=0.92u as=0.152p ps=1.64u w=0.22u l=0.28u
X5 VSS IN1.t1 GF_INV_MAG_1.IN VSS.t0 nfet_03v3 ad=0.152p pd=1.64u as=86.8f ps=0.92u w=0.22u l=0.28u
R0 VDD.n2 VDD 427.092
R1 VDD.t4 VDD.n2 309.341
R2 VDD.n3 VDD.t4 137.826
R3 VDD.n3 VDD.t2 107.198
R4 VDD.n2 VDD.t0 59.4064
R5 VDD.n0 VDD.t1 5.09407
R6 VDD VDD.t3 4.23293
R7 VDD.n5 VDD.n4 3.1505
R8 VDD.n4 VDD.n3 3.1505
R9 VDD.n4 VDD.n1 0.474694
R10 VDD.n5 VDD.n0 0.388218
R11 VDD VDD.n0 0.0709717
R12 VDD VDD.n5 0.00579412
R13 OUT.n2 OUT.n1 9.33985
R14 OUT.n2 OUT.n0 5.17836
R15 OUT OUT.n2 0.0749828
R16 IN2.n0 IN2.t0 40.2519
R17 IN2.n0 IN2.t1 15.3826
R18 IN2 IN2.n0 4.07224
R19 VSS.n6 VSS.t0 889.665
R20 VSS.n6 VSS.t3 635.476
R21 VSS.n1 VSS.t5 54.4698
R22 VSS VSS.t4 9.43705
R23 VSS.n4 VSS.n0 9.3221
R24 VSS.n3 VSS.t6 9.30652
R25 VSS.n2 VSS.n1 5.2005
R26 VSS.n8 VSS.n7 2.6005
R27 VSS.n7 VSS.n6 2.6005
R28 VSS.n7 VSS.n5 0.301575
R29 VSS.n4 VSS.n3 0.184546
R30 VSS.n8 VSS.n4 0.136634
R31 VSS.n3 VSS.n2 0.0675755
R32 VSS VSS.n8 0.00352521
R33 VSS.n2 VSS 0.00219811
R34 IN1.n0 IN1.t0 30.6344
R35 IN1.n0 IN1.t1 27.3855
R36 IN1 IN1.n0 4.07551
C0 IN1 OUT 2.11e-19
C1 IN1 IN2 0.0443f
C2 IN1 VDD 0.135f
C3 a_560_998# IN1 0.0129f
C4 GF_INV_MAG_1.IN OUT 0.126f
C5 GF_INV_MAG_1.IN IN2 0.0394f
C6 GF_INV_MAG_1.IN VDD 0.408f
C7 a_560_998# GF_INV_MAG_1.IN 0.132f
C8 VDD OUT 0.152f
C9 IN1 GF_INV_MAG_1.IN 0.162f
C10 IN2 VDD 0.142f
C11 a_560_998# IN2 8.64e-19
C12 a_560_998# VDD 0.165f
C13 IN1 VSS 0.196f
C14 IN2 VSS 0.264f
C15 OUT VSS 0.176f
C16 GF_INV_MAG_1.IN VSS 0.605f
C17 a_560_998# VSS 0.0247f
C18 VDD VSS 2.01f
.ends

