magic
tech gf180mcuC
magscale 1 10
timestamp 1714558796
<< nwell >>
rect 11105 3381 11205 3455
rect 11434 3340 11543 3356
rect 11434 3336 11457 3340
rect 11434 3312 11438 3336
rect 11489 3312 11543 3340
rect 11932 3300 12034 3312
<< nsubdiff >>
rect 11190 3478 11420 3484
rect 11190 3419 12034 3478
rect 11190 3391 11420 3419
rect 11190 3300 11283 3391
rect 140 2192 667 2199
rect 795 2192 867 2199
rect 140 2094 882 2192
rect 140 2037 667 2094
rect 795 2039 882 2094
<< metal1 >>
rect 1453 4969 1466 5014
rect 12029 3912 12188 3981
rect 12063 3909 12188 3912
rect 11108 3392 11224 3490
rect -125 1389 -47 3374
rect 11434 3312 11543 3356
rect 48 2955 91 2994
rect 7157 2497 7274 2724
rect 12119 2627 12188 3909
rect 11927 2558 12188 2627
rect 768 2105 882 2288
rect 12 1600 71 1652
rect -125 1388 28 1389
rect -125 1283 66 1388
<< metal3 >>
rect 1472 622 1530 5018
rect 1473 621 1490 622
use CLK_div_10_mag  CLK_div_10_mag_0
timestamp 1714558667
transform 1 0 0 0 1 0
box -40 0 12197 3533
use CLK_div_10_mag  CLK_div_10_mag_1
timestamp 1714558667
transform -1 0 12072 0 -1 5567
box -40 0 12197 3533
<< labels >>
flabel metal1 -78 2965 -78 2965 0 FreeSans 320 0 0 0 VSS
port 0 nsew
flabel metal1 7204 2612 7204 2612 0 FreeSans 320 0 0 0 VDD
port 1 nsew
flabel metal1 40 1612 40 1612 0 FreeSans 320 0 0 0 CLK
port 2 nsew
flabel metal1 68 2973 68 2973 0 FreeSans 320 0 0 0 Vdiv100
port 3 nsew
flabel metal1 1459 4985 1459 4985 0 FreeSans 320 0 0 0 RST
port 4 nsew
<< end >>
