magic
tech gf180mcuC
magscale 1 10
timestamp 1691673501
<< nwell >>
rect 418 770 1302 828
rect 418 723 1272 770
rect 418 703 1142 723
<< psubdiff >>
rect 24 -228 1695 -215
rect 24 -274 37 -228
rect 83 -274 131 -228
rect 177 -274 225 -228
rect 271 -274 319 -228
rect 365 -274 413 -228
rect 459 -274 507 -228
rect 553 -274 601 -228
rect 647 -274 695 -228
rect 741 -274 789 -228
rect 835 -274 883 -228
rect 929 -274 977 -228
rect 1023 -274 1071 -228
rect 1117 -274 1165 -228
rect 1211 -274 1259 -228
rect 1305 -274 1353 -228
rect 1399 -274 1447 -228
rect 1493 -274 1541 -228
rect 1587 -274 1635 -228
rect 1681 -274 1695 -228
rect 24 -287 1695 -274
<< nsubdiff >>
rect 448 782 1272 795
rect 448 736 461 782
rect 507 736 555 782
rect 601 736 649 782
rect 695 736 743 782
rect 789 736 837 782
rect 883 736 931 782
rect 977 736 1025 782
rect 1071 736 1119 782
rect 1165 736 1213 782
rect 1259 736 1272 782
rect 448 723 1272 736
<< psubdiffcont >>
rect 37 -274 83 -228
rect 131 -274 177 -228
rect 225 -274 271 -228
rect 319 -274 365 -228
rect 413 -274 459 -228
rect 507 -274 553 -228
rect 601 -274 647 -228
rect 695 -274 741 -228
rect 789 -274 835 -228
rect 883 -274 929 -228
rect 977 -274 1023 -228
rect 1071 -274 1117 -228
rect 1165 -274 1211 -228
rect 1259 -274 1305 -228
rect 1353 -274 1399 -228
rect 1447 -274 1493 -228
rect 1541 -274 1587 -228
rect 1635 -274 1681 -228
<< nsubdiffcont >>
rect 461 736 507 782
rect 555 736 601 782
rect 649 736 695 782
rect 743 736 789 782
rect 837 736 883 782
rect 931 736 977 782
rect 1025 736 1071 782
rect 1119 736 1165 782
rect 1213 736 1259 782
<< polysilicon >>
rect 279 396 357 405
rect 279 392 648 396
rect 279 345 292 392
rect 339 345 648 392
rect 279 340 648 345
rect 279 332 357 340
rect 432 162 488 340
rect 752 175 808 430
rect 912 316 968 430
rect 1072 385 1608 420
rect 1072 364 1303 385
rect 1290 339 1303 364
rect 1349 364 1608 385
rect 1349 339 1362 364
rect 1290 326 1362 339
rect 912 260 1128 316
rect 1072 163 1128 260
rect 1552 133 1608 364
rect 112 -8 488 48
rect 592 -8 968 48
rect 1072 -8 1448 48
rect 573 -82 647 -73
rect 695 -82 751 -8
rect 573 -86 751 -82
rect 573 -138 586 -86
rect 634 -138 751 -86
rect 1392 -55 1448 -8
rect 1599 -55 1672 -46
rect 1392 -59 1672 -55
rect 1392 -106 1612 -59
rect 1659 -106 1672 -59
rect 1392 -111 1672 -106
rect 1599 -119 1672 -111
rect 573 -151 647 -138
<< polycontact >>
rect 292 345 339 392
rect 1303 339 1349 385
rect 586 -138 634 -86
rect 1612 -106 1659 -59
<< metal1 >>
rect 418 782 1302 815
rect 418 736 461 782
rect 507 736 555 782
rect 601 736 649 782
rect 695 736 743 782
rect 789 736 837 782
rect 883 736 931 782
rect 977 736 1025 782
rect 1071 736 1119 782
rect 1165 736 1213 782
rect 1259 736 1302 782
rect 418 703 1302 736
rect 675 609 721 703
rect 997 609 1043 703
rect 279 396 350 403
rect 199 392 350 396
rect 199 345 292 392
rect 339 345 350 392
rect 199 340 350 345
rect 279 334 350 340
rect 517 385 563 470
rect 837 385 883 470
rect 1157 442 1783 488
rect 1292 385 1360 396
rect 517 339 1303 385
rect 1349 339 1360 385
rect 517 258 563 339
rect 1292 328 1360 339
rect 37 212 563 258
rect 677 212 1363 258
rect 37 137 83 212
rect 357 137 403 212
rect 677 137 723 212
rect 997 137 1043 212
rect 1317 137 1363 212
rect 1637 137 1683 442
rect 197 24 243 96
rect 517 24 563 98
rect 837 24 883 98
rect 197 -22 883 24
rect 585 -85 645 -75
rect 483 -86 645 -85
rect 483 -138 586 -86
rect 634 -138 645 -86
rect 483 -141 645 -138
rect 585 -149 645 -141
rect 1157 -195 1203 98
rect 1477 -195 1523 98
rect 1601 -56 1659 -48
rect 1601 -59 1780 -56
rect 1601 -106 1612 -59
rect 1659 -106 1780 -59
rect 1601 -112 1780 -106
rect 1601 -117 1659 -112
rect 4 -228 1715 -195
rect 4 -274 37 -228
rect 83 -274 131 -228
rect 177 -274 225 -228
rect 271 -274 319 -228
rect 365 -274 413 -228
rect 459 -274 507 -228
rect 553 -274 601 -228
rect 647 -274 695 -228
rect 741 -274 789 -228
rect 835 -274 883 -228
rect 929 -274 977 -228
rect 1023 -274 1071 -228
rect 1117 -274 1165 -228
rect 1211 -274 1259 -228
rect 1305 -274 1353 -228
rect 1399 -274 1447 -228
rect 1493 -274 1541 -228
rect 1587 -274 1635 -228
rect 1681 -274 1715 -228
rect 4 -307 1715 -274
use nmos_3p3_HZS5UA  nmos_3p3_HZS5UA_0
timestamp 1691478827
transform 1 0 1580 0 1 118
box -140 -118 140 118
use nmos_3p3_JCGST2#0  nmos_3p3_JCGST2_0
timestamp 1691132869
transform 1 0 1260 0 1 118
box -300 -118 300 118
use nmos_3p3_JCGST2#0  nmos_3p3_JCGST2_1
timestamp 1691132869
transform 1 0 300 0 1 118
box -300 -118 300 118
use nmos_3p3_JCGST2#0  nmos_3p3_JCGST2_2
timestamp 1691132869
transform 1 0 780 0 1 118
box -300 -118 300 118
use pmos_3p3_MNVUAR#3  pmos_3p3_MNVUAR_0
timestamp 1691670445
transform 1 0 780 0 1 540
box -202 -230 202 230
use pmos_3p3_MNVUAR#3  pmos_3p3_MNVUAR_1
timestamp 1691670445
transform 1 0 620 0 1 540
box -202 -230 202 230
use pmos_3p3_MNVUAR#3  pmos_3p3_MNVUAR_2
timestamp 1691670445
transform 1 0 1100 0 1 540
box -202 -230 202 230
use pmos_3p3_MNVUAR#3  pmos_3p3_MNVUAR_3
timestamp 1691670445
transform 1 0 940 0 1 540
box -202 -230 202 230
<< labels >>
flabel metal1 493 -115 493 -115 0 FreeSans 320 0 0 0 B
port 2 nsew
flabel metal1 1760 462 1760 462 0 FreeSans 320 0 0 0 OUT
port 5 nsew
flabel nsubdiffcont 860 759 860 759 0 FreeSans 320 0 0 0 VDD
port 6 nsew
flabel psubdiff 858 -251 858 -251 0 FreeSans 320 0 0 0 VSS
port 8 nsew
flabel metal1 1770 -86 1770 -86 0 FreeSans 320 180 0 0 C
port 3 nsew
flabel metal1 213 362 213 362 0 FreeSans 320 0 0 0 A
port 1 nsew
<< end >>
