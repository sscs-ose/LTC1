magic
tech gf180mcuC
magscale 1 10
timestamp 1693916241
<< pwell >>
rect -540 -368 540 368
<< nmos >>
rect -428 -300 -372 300
rect -268 -300 -212 300
rect -108 -300 -52 300
rect 52 -300 108 300
rect 212 -300 268 300
rect 372 -300 428 300
<< ndiff >>
rect -516 287 -428 300
rect -516 -287 -503 287
rect -457 -287 -428 287
rect -516 -300 -428 -287
rect -372 287 -268 300
rect -372 -287 -343 287
rect -297 -287 -268 287
rect -372 -300 -268 -287
rect -212 287 -108 300
rect -212 -287 -183 287
rect -137 -287 -108 287
rect -212 -300 -108 -287
rect -52 287 52 300
rect -52 -287 -23 287
rect 23 -287 52 287
rect -52 -300 52 -287
rect 108 287 212 300
rect 108 -287 137 287
rect 183 -287 212 287
rect 108 -300 212 -287
rect 268 287 372 300
rect 268 -287 297 287
rect 343 -287 372 287
rect 268 -300 372 -287
rect 428 287 516 300
rect 428 -287 457 287
rect 503 -287 516 287
rect 428 -300 516 -287
<< ndiffc >>
rect -503 -287 -457 287
rect -343 -287 -297 287
rect -183 -287 -137 287
rect -23 -287 23 287
rect 137 -287 183 287
rect 297 -287 343 287
rect 457 -287 503 287
<< polysilicon >>
rect -428 300 -372 344
rect -268 300 -212 344
rect -108 300 -52 344
rect 52 300 108 344
rect 212 300 268 344
rect 372 300 428 344
rect -428 -344 -372 -300
rect -268 -344 -212 -300
rect -108 -344 -52 -300
rect 52 -344 108 -300
rect 212 -344 268 -300
rect 372 -344 428 -300
<< metal1 >>
rect -503 287 -457 298
rect -503 -298 -457 -287
rect -343 287 -297 298
rect -343 -298 -297 -287
rect -183 287 -137 298
rect -183 -298 -137 -287
rect -23 287 23 298
rect -23 -298 23 -287
rect 137 287 183 298
rect 137 -298 183 -287
rect 297 287 343 298
rect 297 -298 343 -287
rect 457 287 503 298
rect 457 -298 503 -287
<< properties >>
string gencell nmos_3p3
string library gf180mcu
string parameters w 3 l 0.280 m 1 nf 6 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
