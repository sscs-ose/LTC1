magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1589 -1285 1589 1285
<< metal1 >>
rect -589 279 589 285
rect -589 253 -583 279
rect -557 253 -507 279
rect -481 253 -431 279
rect -405 253 -355 279
rect -329 253 -279 279
rect -253 253 -203 279
rect -177 253 -127 279
rect -101 253 -51 279
rect -25 253 25 279
rect 51 253 101 279
rect 127 253 177 279
rect 203 253 253 279
rect 279 253 329 279
rect 355 253 405 279
rect 431 253 481 279
rect 507 253 557 279
rect 583 253 589 279
rect -589 203 589 253
rect -589 177 -583 203
rect -557 177 -507 203
rect -481 177 -431 203
rect -405 177 -355 203
rect -329 177 -279 203
rect -253 177 -203 203
rect -177 177 -127 203
rect -101 177 -51 203
rect -25 177 25 203
rect 51 177 101 203
rect 127 177 177 203
rect 203 177 253 203
rect 279 177 329 203
rect 355 177 405 203
rect 431 177 481 203
rect 507 177 557 203
rect 583 177 589 203
rect -589 127 589 177
rect -589 101 -583 127
rect -557 101 -507 127
rect -481 101 -431 127
rect -405 101 -355 127
rect -329 101 -279 127
rect -253 101 -203 127
rect -177 101 -127 127
rect -101 101 -51 127
rect -25 101 25 127
rect 51 101 101 127
rect 127 101 177 127
rect 203 101 253 127
rect 279 101 329 127
rect 355 101 405 127
rect 431 101 481 127
rect 507 101 557 127
rect 583 101 589 127
rect -589 51 589 101
rect -589 25 -583 51
rect -557 25 -507 51
rect -481 25 -431 51
rect -405 25 -355 51
rect -329 25 -279 51
rect -253 25 -203 51
rect -177 25 -127 51
rect -101 25 -51 51
rect -25 25 25 51
rect 51 25 101 51
rect 127 25 177 51
rect 203 25 253 51
rect 279 25 329 51
rect 355 25 405 51
rect 431 25 481 51
rect 507 25 557 51
rect 583 25 589 51
rect -589 -25 589 25
rect -589 -51 -583 -25
rect -557 -51 -507 -25
rect -481 -51 -431 -25
rect -405 -51 -355 -25
rect -329 -51 -279 -25
rect -253 -51 -203 -25
rect -177 -51 -127 -25
rect -101 -51 -51 -25
rect -25 -51 25 -25
rect 51 -51 101 -25
rect 127 -51 177 -25
rect 203 -51 253 -25
rect 279 -51 329 -25
rect 355 -51 405 -25
rect 431 -51 481 -25
rect 507 -51 557 -25
rect 583 -51 589 -25
rect -589 -101 589 -51
rect -589 -127 -583 -101
rect -557 -127 -507 -101
rect -481 -127 -431 -101
rect -405 -127 -355 -101
rect -329 -127 -279 -101
rect -253 -127 -203 -101
rect -177 -127 -127 -101
rect -101 -127 -51 -101
rect -25 -127 25 -101
rect 51 -127 101 -101
rect 127 -127 177 -101
rect 203 -127 253 -101
rect 279 -127 329 -101
rect 355 -127 405 -101
rect 431 -127 481 -101
rect 507 -127 557 -101
rect 583 -127 589 -101
rect -589 -177 589 -127
rect -589 -203 -583 -177
rect -557 -203 -507 -177
rect -481 -203 -431 -177
rect -405 -203 -355 -177
rect -329 -203 -279 -177
rect -253 -203 -203 -177
rect -177 -203 -127 -177
rect -101 -203 -51 -177
rect -25 -203 25 -177
rect 51 -203 101 -177
rect 127 -203 177 -177
rect 203 -203 253 -177
rect 279 -203 329 -177
rect 355 -203 405 -177
rect 431 -203 481 -177
rect 507 -203 557 -177
rect 583 -203 589 -177
rect -589 -253 589 -203
rect -589 -279 -583 -253
rect -557 -279 -507 -253
rect -481 -279 -431 -253
rect -405 -279 -355 -253
rect -329 -279 -279 -253
rect -253 -279 -203 -253
rect -177 -279 -127 -253
rect -101 -279 -51 -253
rect -25 -279 25 -253
rect 51 -279 101 -253
rect 127 -279 177 -253
rect 203 -279 253 -253
rect 279 -279 329 -253
rect 355 -279 405 -253
rect 431 -279 481 -253
rect 507 -279 557 -253
rect 583 -279 589 -253
rect -589 -285 589 -279
<< via1 >>
rect -583 253 -557 279
rect -507 253 -481 279
rect -431 253 -405 279
rect -355 253 -329 279
rect -279 253 -253 279
rect -203 253 -177 279
rect -127 253 -101 279
rect -51 253 -25 279
rect 25 253 51 279
rect 101 253 127 279
rect 177 253 203 279
rect 253 253 279 279
rect 329 253 355 279
rect 405 253 431 279
rect 481 253 507 279
rect 557 253 583 279
rect -583 177 -557 203
rect -507 177 -481 203
rect -431 177 -405 203
rect -355 177 -329 203
rect -279 177 -253 203
rect -203 177 -177 203
rect -127 177 -101 203
rect -51 177 -25 203
rect 25 177 51 203
rect 101 177 127 203
rect 177 177 203 203
rect 253 177 279 203
rect 329 177 355 203
rect 405 177 431 203
rect 481 177 507 203
rect 557 177 583 203
rect -583 101 -557 127
rect -507 101 -481 127
rect -431 101 -405 127
rect -355 101 -329 127
rect -279 101 -253 127
rect -203 101 -177 127
rect -127 101 -101 127
rect -51 101 -25 127
rect 25 101 51 127
rect 101 101 127 127
rect 177 101 203 127
rect 253 101 279 127
rect 329 101 355 127
rect 405 101 431 127
rect 481 101 507 127
rect 557 101 583 127
rect -583 25 -557 51
rect -507 25 -481 51
rect -431 25 -405 51
rect -355 25 -329 51
rect -279 25 -253 51
rect -203 25 -177 51
rect -127 25 -101 51
rect -51 25 -25 51
rect 25 25 51 51
rect 101 25 127 51
rect 177 25 203 51
rect 253 25 279 51
rect 329 25 355 51
rect 405 25 431 51
rect 481 25 507 51
rect 557 25 583 51
rect -583 -51 -557 -25
rect -507 -51 -481 -25
rect -431 -51 -405 -25
rect -355 -51 -329 -25
rect -279 -51 -253 -25
rect -203 -51 -177 -25
rect -127 -51 -101 -25
rect -51 -51 -25 -25
rect 25 -51 51 -25
rect 101 -51 127 -25
rect 177 -51 203 -25
rect 253 -51 279 -25
rect 329 -51 355 -25
rect 405 -51 431 -25
rect 481 -51 507 -25
rect 557 -51 583 -25
rect -583 -127 -557 -101
rect -507 -127 -481 -101
rect -431 -127 -405 -101
rect -355 -127 -329 -101
rect -279 -127 -253 -101
rect -203 -127 -177 -101
rect -127 -127 -101 -101
rect -51 -127 -25 -101
rect 25 -127 51 -101
rect 101 -127 127 -101
rect 177 -127 203 -101
rect 253 -127 279 -101
rect 329 -127 355 -101
rect 405 -127 431 -101
rect 481 -127 507 -101
rect 557 -127 583 -101
rect -583 -203 -557 -177
rect -507 -203 -481 -177
rect -431 -203 -405 -177
rect -355 -203 -329 -177
rect -279 -203 -253 -177
rect -203 -203 -177 -177
rect -127 -203 -101 -177
rect -51 -203 -25 -177
rect 25 -203 51 -177
rect 101 -203 127 -177
rect 177 -203 203 -177
rect 253 -203 279 -177
rect 329 -203 355 -177
rect 405 -203 431 -177
rect 481 -203 507 -177
rect 557 -203 583 -177
rect -583 -279 -557 -253
rect -507 -279 -481 -253
rect -431 -279 -405 -253
rect -355 -279 -329 -253
rect -279 -279 -253 -253
rect -203 -279 -177 -253
rect -127 -279 -101 -253
rect -51 -279 -25 -253
rect 25 -279 51 -253
rect 101 -279 127 -253
rect 177 -279 203 -253
rect 253 -279 279 -253
rect 329 -279 355 -253
rect 405 -279 431 -253
rect 481 -279 507 -253
rect 557 -279 583 -253
<< metal2 >>
rect -589 279 589 285
rect -589 253 -583 279
rect -557 253 -507 279
rect -481 253 -431 279
rect -405 253 -355 279
rect -329 253 -279 279
rect -253 253 -203 279
rect -177 253 -127 279
rect -101 253 -51 279
rect -25 253 25 279
rect 51 253 101 279
rect 127 253 177 279
rect 203 253 253 279
rect 279 253 329 279
rect 355 253 405 279
rect 431 253 481 279
rect 507 253 557 279
rect 583 253 589 279
rect -589 203 589 253
rect -589 177 -583 203
rect -557 177 -507 203
rect -481 177 -431 203
rect -405 177 -355 203
rect -329 177 -279 203
rect -253 177 -203 203
rect -177 177 -127 203
rect -101 177 -51 203
rect -25 177 25 203
rect 51 177 101 203
rect 127 177 177 203
rect 203 177 253 203
rect 279 177 329 203
rect 355 177 405 203
rect 431 177 481 203
rect 507 177 557 203
rect 583 177 589 203
rect -589 127 589 177
rect -589 101 -583 127
rect -557 101 -507 127
rect -481 101 -431 127
rect -405 101 -355 127
rect -329 101 -279 127
rect -253 101 -203 127
rect -177 101 -127 127
rect -101 101 -51 127
rect -25 101 25 127
rect 51 101 101 127
rect 127 101 177 127
rect 203 101 253 127
rect 279 101 329 127
rect 355 101 405 127
rect 431 101 481 127
rect 507 101 557 127
rect 583 101 589 127
rect -589 51 589 101
rect -589 25 -583 51
rect -557 25 -507 51
rect -481 25 -431 51
rect -405 25 -355 51
rect -329 25 -279 51
rect -253 25 -203 51
rect -177 25 -127 51
rect -101 25 -51 51
rect -25 25 25 51
rect 51 25 101 51
rect 127 25 177 51
rect 203 25 253 51
rect 279 25 329 51
rect 355 25 405 51
rect 431 25 481 51
rect 507 25 557 51
rect 583 25 589 51
rect -589 -25 589 25
rect -589 -51 -583 -25
rect -557 -51 -507 -25
rect -481 -51 -431 -25
rect -405 -51 -355 -25
rect -329 -51 -279 -25
rect -253 -51 -203 -25
rect -177 -51 -127 -25
rect -101 -51 -51 -25
rect -25 -51 25 -25
rect 51 -51 101 -25
rect 127 -51 177 -25
rect 203 -51 253 -25
rect 279 -51 329 -25
rect 355 -51 405 -25
rect 431 -51 481 -25
rect 507 -51 557 -25
rect 583 -51 589 -25
rect -589 -101 589 -51
rect -589 -127 -583 -101
rect -557 -127 -507 -101
rect -481 -127 -431 -101
rect -405 -127 -355 -101
rect -329 -127 -279 -101
rect -253 -127 -203 -101
rect -177 -127 -127 -101
rect -101 -127 -51 -101
rect -25 -127 25 -101
rect 51 -127 101 -101
rect 127 -127 177 -101
rect 203 -127 253 -101
rect 279 -127 329 -101
rect 355 -127 405 -101
rect 431 -127 481 -101
rect 507 -127 557 -101
rect 583 -127 589 -101
rect -589 -177 589 -127
rect -589 -203 -583 -177
rect -557 -203 -507 -177
rect -481 -203 -431 -177
rect -405 -203 -355 -177
rect -329 -203 -279 -177
rect -253 -203 -203 -177
rect -177 -203 -127 -177
rect -101 -203 -51 -177
rect -25 -203 25 -177
rect 51 -203 101 -177
rect 127 -203 177 -177
rect 203 -203 253 -177
rect 279 -203 329 -177
rect 355 -203 405 -177
rect 431 -203 481 -177
rect 507 -203 557 -177
rect 583 -203 589 -177
rect -589 -253 589 -203
rect -589 -279 -583 -253
rect -557 -279 -507 -253
rect -481 -279 -431 -253
rect -405 -279 -355 -253
rect -329 -279 -279 -253
rect -253 -279 -203 -253
rect -177 -279 -127 -253
rect -101 -279 -51 -253
rect -25 -279 25 -253
rect 51 -279 101 -253
rect 127 -279 177 -253
rect 203 -279 253 -253
rect 279 -279 329 -253
rect 355 -279 405 -253
rect 431 -279 481 -253
rect 507 -279 557 -253
rect 583 -279 589 -253
rect -589 -285 589 -279
<< end >>
