* NGSPICE file created from CP_flat.ext - technology: gf180mcuC

.subckt loop_filter_V1_pex VDD ITAIL ITAIL1 VCTRL UP down VSS
X0 ITAIL ITAIL.t14 VDD.t20 VDD.t5 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X1 VDD a_n638_n190# a_n374_n194.t11 VDD.t21 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X2 VSS ITAIL1.t2 ITAIL1.t3 VSS.t12 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X3 VSS down.t0 a_n166_n835# VSS.t3 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X4 ITAIL ITAIL.t12 VDD.t19 VDD.t13 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X5 VCTRL ITAIL1.t8 a_n166_n835# VSS.t5 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X6 VDD ITAIL.t10 ITAIL.t11 VDD.t12 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X7 VCTRL ITAIL.t19 a_n374_n194.t6 VDD.t5 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X8 a_n638_n190# UP.t0 VSS.t21 VSS.t20 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X9 a_n166_n835# down.t1 VSS.t22 VSS.t3 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X10 VCTRL ITAIL1.t9 a_n166_n835# VSS.t3 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X11 VDD ITAIL.t8 ITAIL.t9 VDD.t12 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X12 VCTRL ITAIL.t20 a_n374_n194.t5 VDD.t5 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X13 VCTRL ITAIL.t21 a_n374_n194.t4 VDD.t13 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X14 a_n166_n835# down.t2 VSS.t4 VSS.t3 nfet_03v3 ad=92.8f pd=0.92u as=92.8f ps=0.92u w=0.28u l=0.56u
X15 VCTRL ITAIL.t22 a_n374_n194.t3 VDD.t13 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X16 a_n638_n190# UP.t1 VDD.t1 VDD.t0 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X17 VSS ITAIL1.t0 ITAIL1.t1 VSS.t7 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X18 VDD a_n638_n190# a_n374_n194.t10 VDD.t21 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X19 VDD a_n638_n190# a_n374_n194.t9 VDD.t21 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X20 a_n638_n190# UP.t2 VDD.t4 VDD.t0 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X21 a_n166_n835# ITAIL1.t10 VCTRL.t9 VSS.t9 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X22 a_n638_n190# UP.t3 VSS.t16 VSS.t15 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X23 ITAIL1 ITAIL1.t6 VSS.t8 VSS.t7 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X24 a_n638_n190# UP.t4 VDD.t3 VDD.t0 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X25 ITAIL ITAIL.t0 VDD.t14 VDD.t13 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X26 a_n638_n190# UP.t5 VDD.t2 VDD.t0 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X27 VDD a_n638_n190# a_n374_n194.t8 VDD.t21 pfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.56u
X28 VSS down.t3 a_n166_n835# VSS.t0 nfet_03v3 ad=0.158p pd=1.64u as=92.8f ps=0.92u w=0.28u l=0.56u
X29 a_n166_n835# down.t4 VSS.t17 VSS.t0 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
X30 VDD ITAIL.t6 ITAIL.t7 VDD.t7 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X31 ITAIL1 ITAIL1.t4 VSS.t6 VSS.t0 nfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X32 VDD ITAIL.t4 ITAIL.t5 VDD.t7 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X33 ITAIL ITAIL.t2 VDD.t6 VDD.t5 pfet_03v3 ad=0.158p pd=1.64u as=0.158p ps=1.64u w=0.28u l=0.56u
X34 a_n166_n835# ITAIL1.t13 VCTRL.t11 VSS.t5 nfet_03v3 ad=92.8f pd=0.92u as=0.158p ps=1.64u w=0.28u l=0.56u
R0 ITAIL.n0 ITAIL.t2 10.9054
R1 ITAIL.n12 ITAIL.t23 10.8613
R2 ITAIL.n12 ITAIL.t4 10.5984
R3 ITAIL.n0 ITAIL.t20 10.5336
R4 ITAIL.n13 ITAIL.t25 10.5334
R5 ITAIL.n25 ITAIL.t10 10.0523
R6 ITAIL.n20 ITAIL.t19 9.85461
R7 ITAIL.n45 ITAIL.t22 9.78943
R8 ITAIL.n31 ITAIL.t8 9.78943
R9 ITAIL.n3 ITAIL.t14 9.72546
R10 ITAIL.n28 ITAIL.t16 9.72425
R11 ITAIL.n36 ITAIL.t26 9.65907
R12 ITAIL.n32 ITAIL.t0 9.65907
R13 ITAIL.n16 ITAIL.t6 9.65907
R14 ITAIL.n55 ITAIL.t12 8.55104
R15 ITAIL.n34 ITAIL.n33 7.7573
R16 ITAIL.n51 ITAIL.n29 7.7433
R17 ITAIL.n9 ITAIL.n8 7.69237
R18 ITAIL.n9 ITAIL.t5 7.66468
R19 ITAIL.n42 ITAIL.t9 7.5883
R20 ITAIL.n10 ITAIL.n7 7.58811
R21 ITAIL.n11 ITAIL.t7 7.39887
R22 ITAIL.n27 ITAIL.t21 7.34965
R23 ITAIL.n61 ITAIL.t11 7.33058
R24 ITAIL ITAIL.n68 4.63009
R25 ITAIL.n63 ITAIL.n27 2.2505
R26 ITAIL.n4 ITAIL.n3 1.50717
R27 ITAIL.n18 ITAIL.n17 1.5029
R28 ITAIL.n56 ITAIL.n55 1.5005
R29 ITAIL.n47 ITAIL.n31 1.5005
R30 ITAIL.n38 ITAIL.n32 1.5005
R31 ITAIL.n46 ITAIL.n45 1.12992
R32 ITAIL.n65 ITAIL.n25 1.12943
R33 ITAIL.n21 ITAIL.n20 1.12721
R34 ITAIL.n37 ITAIL.n36 1.12703
R35 ITAIL.n58 ITAIL.n28 1.1255
R36 ITAIL.n13 ITAIL.n12 0.390708
R37 ITAIL.n14 ITAIL.n13 0.357771
R38 ITAIL.n1 ITAIL.n0 0.341087
R39 ITAIL.n6 ITAIL.n5 0.328487
R40 ITAIL.n10 ITAIL.n9 0.106635
R41 ITAIL.n11 ITAIL.n10 0.106083
R42 ITAIL.n68 ITAIL.n23 0.0746286
R43 ITAIL.n21 ITAIL.n19 0.0444571
R44 ITAIL.n19 ITAIL.n18 0.0425807
R45 ITAIL.n19 ITAIL.n11 0.0323939
R46 ITAIL.n42 ITAIL.n41 0.0323094
R47 ITAIL.n51 ITAIL.n50 0.0321928
R48 ITAIL.n68 ITAIL.n67 0.0320905
R49 ITAIL.n61 ITAIL.n60 0.0320216
R50 ITAIL.n4 ITAIL.n1 0.028981
R51 ITAIL.n62 ITAIL.n61 0.0167151
R52 ITAIL.n5 ITAIL.n4 0.0163348
R53 ITAIL.n43 ITAIL.n42 0.015769
R54 ITAIL.n52 ITAIL.n51 0.0134294
R55 ITAIL.n15 ITAIL.n14 0.0107874
R56 ITAIL.n27 ITAIL.n26 0.00997368
R57 ITAIL.n22 ITAIL.n6 0.0061962
R58 ITAIL.n46 ITAIL.n44 0.00569669
R59 ITAIL.n23 ITAIL.n22 0.00498133
R60 ITAIL.n49 ITAIL.n48 0.00444881
R61 ITAIL.n37 ITAIL.n34 0.00412886
R62 ITAIL.n60 ITAIL.n59 0.00346161
R63 ITAIL.n18 ITAIL.n15 0.00342167
R64 ITAIL.n58 ITAIL.n57 0.00329708
R65 ITAIL.n53 ITAIL.n52 0.00329708
R66 ITAIL.n67 ITAIL.n66 0.00313254
R67 ITAIL.n41 ITAIL.n40 0.00306266
R68 ITAIL.n40 ITAIL.n39 0.00304881
R69 ITAIL.n22 ITAIL.n21 0.00260507
R70 ITAIL.n25 ITAIL.n24 0.00245007
R71 ITAIL.n3 ITAIL.n2 0.00242648
R72 ITAIL.n66 ITAIL.n65 0.00214534
R73 ITAIL.n38 ITAIL.n37 0.00198191
R74 ITAIL.n65 ITAIL.n64 0.0019808
R75 ITAIL.n64 ITAIL.n63 0.00181627
R76 ITAIL.n63 ITAIL.n62 0.00181627
R77 ITAIL.n59 ITAIL.n58 0.00181627
R78 ITAIL.n56 ITAIL.n53 0.00181627
R79 ITAIL.n55 ITAIL.n54 0.00175
R80 ITAIL.n36 ITAIL.n35 0.00168421
R81 ITAIL.n31 ITAIL.n30 0.00166883
R82 ITAIL.n17 ITAIL.n16 0.00155882
R83 ITAIL.n47 ITAIL.n46 0.0014166
R84 ITAIL.n50 ITAIL.n49 0.000829068
R85 ITAIL.n57 ITAIL.n56 0.000664534
R86 ITAIL.n48 ITAIL.n47 0.000664534
R87 ITAIL.n44 ITAIL.n43 0.000664534
R88 ITAIL.n39 ITAIL.n38 0.000664534
R89 VCTRL.n1 VCTRL.n0 9.42182
R90 VCTRL.n6 VCTRL.n5 9.3792
R91 VCTRL.n12 VCTRL.n11 9.07899
R92 VCTRL.n6 VCTRL.t5 8.84311
R93 VCTRL.n9 VCTRL.t2 8.83779
R94 VCTRL.n8 VCTRL.n7 8.83029
R95 VCTRL.n3 VCTRL.n2 8.83029
R96 VCTRL.n1 VCTRL.t3 8.79474
R97 VCTRL.n4 VCTRL.t4 8.76273
R98 VCTRL.n14 VCTRL.n13 8.5505
R99 VCTRL.n12 VCTRL.t11 8.5505
R100 VCTRL.n15 VCTRL.t9 8.03277
R101 VCTRL VCTRL.n15 3.84211
R102 VCTRL.n10 VCTRL.n9 1.92684
R103 VCTRL VCTRL.n10 1.72887
R104 VCTRL.n14 VCTRL.n12 1.1179
R105 VCTRL.n3 VCTRL.n1 0.576883
R106 VCTRL.n4 VCTRL.n3 0.571972
R107 VCTRL.n9 VCTRL.n8 0.550283
R108 VCTRL.n8 VCTRL.n6 0.544413
R109 VCTRL.n15 VCTRL.n14 0.454295
R110 VCTRL.n10 VCTRL.n4 0.112274
R111 a_n374_n194.n5 a_n374_n194.n4 10.0413
R112 a_n374_n194.n10 a_n374_n194.t4 8.81226
R113 a_n374_n194.n5 a_n374_n194.n3 8.80202
R114 a_n374_n194.n11 a_n374_n194.t3 8.78441
R115 a_n374_n194.n8 a_n374_n194.t6 8.6005
R116 a_n374_n194.n0 a_n374_n194.t5 7.89525
R117 a_n374_n194.n0 a_n374_n194.n6 7.89324
R118 a_n374_n194.n0 a_n374_n194.n7 7.72809
R119 a_n374_n194.n1 a_n374_n194.t8 5.72901
R120 a_n374_n194.n1 a_n374_n194.t9 5.2005
R121 a_n374_n194.n2 a_n374_n194.t11 5.2005
R122 a_n374_n194.t10 a_n374_n194.n12 5.2005
R123 a_n374_n194.n8 a_n374_n194.n0 2.56002
R124 a_n374_n194.n9 a_n374_n194.n5 2.34763
R125 a_n374_n194.n10 a_n374_n194.n9 2.1305
R126 a_n374_n194.n12 a_n374_n194.n11 1.88322
R127 a_n374_n194.n11 a_n374_n194.n10 1.10344
R128 a_n374_n194.n2 a_n374_n194.n1 0.529011
R129 a_n374_n194.n12 a_n374_n194.n2 0.529011
R130 a_n374_n194.n9 a_n374_n194.n8 0.294424
R131 VDD.n20 VDD.t7 47.9334
R132 VDD.n35 VDD.t13 45.5368
R133 VDD.n28 VDD.t12 33.5535
R134 VDD.n48 VDD.t0 31.1569
R135 VDD.n5 VDD.n4 9.4133
R136 VDD.n49 VDD.t2 9.02932
R137 VDD.n7 VDD.n6 8.82188
R138 VDD.n5 VDD.t20 8.79795
R139 VDD.n49 VDD.t3 8.6005
R140 VDD.n50 VDD.t1 8.6005
R141 VDD.n51 VDD.t4 8.6005
R142 VDD.n18 VDD.n0 7.5859
R143 VDD.n71 VDD.t14 7.58462
R144 VDD.n70 VDD.t19 7.58462
R145 VDD.n24 VDD.t5 7.19043
R146 VDD.n63 VDD.t21 7.19043
R147 VDD.n14 VDD.n13 6.44895
R148 VDD.n60 VDD.n59 6.3005
R149 VDD.n55 VDD.n47 6.3005
R150 VDD.n53 VDD.n48 6.3005
R151 VDD.n69 VDD.n36 6.3005
R152 VDD.n21 VDD.n20 6.3005
R153 VDD.n23 VDD.n22 6.3005
R154 VDD.n25 VDD.n24 6.3005
R155 VDD.n27 VDD.n26 6.3005
R156 VDD.n29 VDD.n28 6.3005
R157 VDD.n78 VDD.n34 6.3005
R158 VDD.n77 VDD.n35 6.3005
R159 VDD.n8 VDD.t6 6.27989
R160 VDD.n41 VDD.n40 5.7405
R161 VDD.n43 VDD.n37 5.2005
R162 VDD.n42 VDD.n38 5.2005
R163 VDD.n41 VDD.n39 5.2005
R164 VDD.n10 VDD.n1 4.5005
R165 VDD.n16 VDD.n15 4.5005
R166 VDD.n62 VDD.n61 4.5005
R167 VDD.n9 VDD.n8 3.15744
R168 VDD.n65 VDD.n64 3.1505
R169 VDD.n64 VDD.n63 3.1505
R170 VDD.n33 VDD.n32 3.1505
R171 VDD.n32 VDD.n31 3.1505
R172 VDD.n76 VDD.n75 2.55963
R173 VDD.n19 VDD.n18 2.50553
R174 VDD.n57 VDD.n46 2.25076
R175 VDD.n10 VDD.n9 2.2505
R176 VDD.n64 VDD.n60 1.5405
R177 VDD.n64 VDD.n62 1.1905
R178 VDD.n67 VDD.n43 0.845717
R179 VDD.n8 VDD.n7 0.735716
R180 VDD.n75 VDD.n70 0.604129
R181 VDD.n7 VDD.n5 0.576883
R182 VDD.n74 VDD.n72 0.543743
R183 VDD.n43 VDD.n42 0.5405
R184 VDD.n42 VDD.n41 0.5405
R185 VDD.n72 VDD.n71 0.482825
R186 VDD.n52 VDD.n51 0.431971
R187 VDD.n51 VDD.n50 0.429324
R188 VDD.n50 VDD.n49 0.429324
R189 VDD.n18 VDD.n17 0.40301
R190 VDD.n32 VDD.n30 0.2105
R191 VDD.n74 VDD.n73 0.205675
R192 VDD.n46 VDD.n44 0.154098
R193 VDD.n21 VDD.n19 0.08917
R194 VDD.n23 VDD.n21 0.08917
R195 VDD.n25 VDD.n23 0.08917
R196 VDD.n27 VDD.n25 0.08917
R197 VDD.n29 VDD.n27 0.08917
R198 VDD.n33 VDD.n29 0.08917
R199 VDD.n78 VDD.n77 0.08917
R200 VDD VDD.n78 0.0878399
R201 VDD.n53 VDD.n52 0.071122
R202 VDD.n76 VDD.n69 0.0664791
R203 VDD.n56 VDD.n55 0.0646627
R204 VDD.n54 VDD.n53 0.0452847
R205 VDD.n67 VDD.n66 0.042701
R206 VDD.n55 VDD.n54 0.0418397
R207 VDD.n75 VDD.n74 0.0357448
R208 VDD.n46 VDD.n45 0.0347499
R209 VDD.n68 VDD.n67 0.0244531
R210 VDD.n77 VDD.n76 0.0231108
R211 VDD.n17 VDD.n16 0.0168043
R212 VDD.n10 VDD.n2 0.0155
R213 VDD.n69 VDD.n68 0.0114756
R214 VDD.n15 VDD.n14 0.0103544
R215 VDD.n66 VDD.n65 0.00997368
R216 VDD.n57 VDD.n56 0.00997368
R217 VDD.n65 VDD.n58 0.00782057
R218 VDD.n15 VDD.n12 0.00725
R219 VDD.n58 VDD.n57 0.00566746
R220 VDD.n9 VDD.n3 0.00283766
R221 VDD.n16 VDD.n11 0.00245652
R222 VDD VDD.n33 0.00183005
R223 VDD.n11 VDD.n10 0.00180435
R224 ITAIL1.n5 ITAIL1.n4 28.0418
R225 ITAIL1.n3 ITAIL1.n2 14.6005
R226 ITAIL1.n1 ITAIL1.n0 7.61735
R227 ITAIL1.n1 ITAIL1.t1 7.20135
R228 ITAIL1.n8 ITAIL1.n7 6.82463
R229 ITAIL1.n10 ITAIL1.t2 6.77907
R230 ITAIL1.n5 ITAIL1.t4 6.71389
R231 ITAIL1.n2 ITAIL1.t8 6.51836
R232 ITAIL1.n2 ITAIL1.t6 6.51836
R233 ITAIL1.n3 ITAIL1.t13 6.51836
R234 ITAIL1.n10 ITAIL1.t10 6.25764
R235 ITAIL1.n4 ITAIL1.t0 6.25764
R236 ITAIL1.n6 ITAIL1.t9 6.19246
R237 ITAIL1.n11 ITAIL1.t3 5.89613
R238 ITAIL1.n11 ITAIL1.n10 4.23548
R239 ITAIL1.n8 ITAIL1.n6 4.21461
R240 ITAIL1 ITAIL1.n12 2.92243
R241 ITAIL1.n9 ITAIL1.n8 1.42665
R242 ITAIL1.n12 ITAIL1.n11 1.13763
R243 ITAIL1.n12 ITAIL1.n9 0.474918
R244 ITAIL1.n4 ITAIL1.n3 0.261214
R245 ITAIL1.n9 ITAIL1.n1 0.2105
R246 ITAIL1.n6 ITAIL1.n5 0.130857
R247 VSS.n17 VSS.t15 267.033
R248 VSS.t9 VSS.t20 177.706
R249 VSS.n3 VSS.t6 11.3982
R250 VSS.n14 VSS.t21 8.88029
R251 VSS.t20 VSS.t0 8.55313
R252 VSS.n3 VSS.n2 8.5505
R253 VSS.n12 VSS.t17 8.5505
R254 VSS.n13 VSS.t22 8.5505
R255 VSS.n11 VSS.n8 8.5505
R256 VSS.n14 VSS.t16 8.5505
R257 VSS.n1 VSS.n0 5.4005
R258 VSS.n1 VSS.t8 5.4005
R259 VSS.n10 VSS.n9 5.4005
R260 VSS.n10 VSS.t4 5.4005
R261 VSS VSS.n7 5.2005
R262 VSS VSS.n7 5.2005
R263 VSS.n5 VSS.n1 3.48846
R264 VSS.n11 VSS.n10 3.25515
R265 VSS.t5 VSS.t12 2.85138
R266 VSS.t7 VSS.t9 2.85138
R267 VSS.n17 VSS.n7 2.6005
R268 VSS.n18 VSS.n17 1.24621
R269 VSS.n4 VSS.n3 1.04354
R270 VSS.t0 VSS.t5 0.950792
R271 VSS.t3 VSS.t7 0.950792
R272 VSS.t15 VSS.t3 0.950792
R273 VSS.n12 VSS.n11 0.699074
R274 VSS.n13 VSS.n12 0.237342
R275 VSS VSS.n18 0.224988
R276 VSS.n16 VSS.n13 0.217211
R277 VSS.n18 VSS.n16 0.20351
R278 VSS.n5 VSS.n4 0.182946
R279 VSS.n15 VSS.n14 0.168475
R280 VSS.n16 VSS.n15 0.0922128
R281 VSS VSS.n6 0.0914091
R282 VSS.n6 VSS.n5 0.0432273
R283 down.n1 down.n0 14.6005
R284 down.n3 down.n2 12.8446
R285 down down.n3 7.49733
R286 down.n0 down.t4 6.51836
R287 down.n0 down.t1 6.51836
R288 down.n1 down.t0 6.51836
R289 down.n3 down.t2 6.388
R290 down.n2 down.t3 6.19246
R291 down.n2 down.n1 0.326393
R292 UP.t0 UP.t3 12.5148
R293 UP.n3 UP.t0 10.215
R294 UP.n0 UP.t2 10.1117
R295 UP.n1 UP.t4 9.54068
R296 UP.n2 UP.t5 9.4755
R297 UP.n0 UP.t1 9.4755
R298 UP.n2 UP.n1 0.50481
R299 UP.n1 UP.n0 0.501707
R300 UP.n3 UP.n2 0.393086
R301 UP UP.n3 0.287704
C0 ITAIL1 down 0.0774f
C1 VDD ITAIL 6.84f
C2 UP VDD 1.92f
C3 a_n638_n190# VCTRL 5.88e-19
C4 a_n166_n835# VDD 0.00882f
C5 VDD down 0.172f
C6 a_n638_n190# ITAIL 0.0168f
C7 ITAIL1 VDD 0.531f
C8 UP a_n638_n190# 1.4f
C9 a_n638_n190# down 0.0496f
C10 ITAIL1 a_n638_n190# 2.45e-19
C11 VCTRL ITAIL 2.14f
C12 UP VCTRL 1.07e-19
C13 VDD a_n638_n190# 1.23f
C14 a_n166_n835# VCTRL 0.509f
C15 VCTRL down 0.0026f
C16 UP ITAIL 0.0149f
C17 ITAIL1 VCTRL 1.35f
C18 a_n166_n835# ITAIL 0.00187f
C19 down ITAIL 0.0122f
C20 a_n166_n835# UP 2.33e-20
C21 ITAIL1 ITAIL 0.0091f
C22 UP down 0.0605f
C23 VDD VCTRL 1.09f
C24 ITAIL1 UP 4.3e-19
C25 a_n166_n835# down 0.13f
C26 a_n166_n835# ITAIL1 0.655f
.ends

