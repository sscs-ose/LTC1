magic
tech gf180mcuC
magscale 1 10
timestamp 1692805350
<< nwell >>
rect 65 1023 533 1603
rect 61 267 529 847
rect 846 715 1723 1597
rect 61 -488 529 92
rect 846 -232 1405 492
rect 2698 -514 3609 1410
rect 4612 -514 5523 1410
rect 6526 -514 7057 1410
<< pwell >>
rect -163 1023 35 1603
rect -167 267 31 847
rect 1765 715 1963 1597
rect -167 -488 31 92
rect 1511 -190 1709 602
rect 1511 -555 1709 -267
rect 2428 -452 2626 1348
rect 3681 -452 3879 1348
rect 4342 -452 4540 1348
rect 5595 -452 5793 1348
rect 6256 -452 6454 1348
<< nmos >>
rect -89 1369 -39 1425
rect -89 1201 -39 1257
rect 1839 1363 1889 1419
rect 1839 1195 1889 1251
rect 1839 893 1889 949
rect -93 613 -43 669
rect 2502 1176 2552 1232
rect 2502 1008 2552 1064
rect 2502 840 2552 896
rect 3755 1176 3805 1232
rect 4416 1176 4466 1232
rect 3755 1008 3805 1064
rect 4416 1008 4466 1064
rect 3755 840 3805 896
rect 2502 672 2552 728
rect 4416 840 4466 896
rect -93 445 -43 501
rect 1585 430 1635 486
rect 3755 672 3805 728
rect 5669 1176 5719 1232
rect 6330 1176 6380 1232
rect 5669 1008 5719 1064
rect 6330 1008 6380 1064
rect 5669 840 5719 896
rect 2502 504 2552 560
rect 4416 672 4466 728
rect 6330 840 6380 896
rect 3755 504 3805 560
rect 5669 672 5719 728
rect 2502 336 2552 392
rect 1585 262 1635 318
rect 2502 168 2552 224
rect 4416 504 4466 560
rect -93 -142 -43 -86
rect 1585 94 1635 150
rect -93 -310 -43 -254
rect 1585 -74 1635 -18
rect 3755 336 3805 392
rect 6330 672 6380 728
rect 5669 504 5719 560
rect 4416 336 4466 392
rect 3755 168 3805 224
rect 2502 0 2552 56
rect 2502 -168 2552 -112
rect 3755 0 3805 56
rect 3755 -168 3805 -112
rect 4416 168 4466 224
rect 6330 504 6380 560
rect 2502 -336 2552 -280
rect 5669 336 5719 392
rect 6330 336 6380 392
rect 5669 168 5719 224
rect 4416 0 4466 56
rect 4416 -168 4466 -112
rect 5669 0 5719 56
rect 1585 -439 1635 -383
rect 3755 -336 3805 -280
rect 5669 -168 5719 -112
rect 6330 168 6380 224
rect 4416 -336 4466 -280
rect 6330 0 6380 56
rect 6330 -168 6380 -112
rect 5669 -336 5719 -280
rect 6330 -336 6380 -280
<< pmos >>
rect 201 1369 251 1425
rect 201 1201 251 1257
rect 1144 1363 1194 1419
rect 1274 1363 1324 1419
rect 1407 1363 1457 1419
rect 1537 1363 1587 1419
rect 1144 1195 1194 1251
rect 1274 1195 1324 1251
rect 1407 1195 1457 1251
rect 1537 1195 1587 1251
rect 1144 893 1194 949
rect 1407 893 1457 949
rect 1537 893 1587 949
rect 197 613 247 669
rect 2834 1176 2884 1232
rect 2834 1008 2884 1064
rect 2834 840 2884 896
rect 3423 1176 3473 1232
rect 3423 1008 3473 1064
rect 4748 1176 4798 1232
rect 4748 1008 4798 1064
rect 3423 840 3473 896
rect 2834 672 2884 728
rect 4748 840 4798 896
rect 197 445 247 501
rect 3423 672 3473 728
rect 5337 1176 5387 1232
rect 5337 1008 5387 1064
rect 6662 1176 6712 1232
rect 6662 1008 6712 1064
rect 5337 840 5387 896
rect 2834 504 2884 560
rect 4748 672 4798 728
rect 6662 840 6712 896
rect 3423 504 3473 560
rect 5337 672 5387 728
rect 2834 336 2884 392
rect 1175 262 1275 318
rect 1175 102 1275 158
rect 2834 168 2884 224
rect 4748 504 4798 560
rect 197 -142 247 -86
rect 1175 -58 1275 -2
rect 197 -310 247 -254
rect 3423 336 3473 392
rect 6662 672 6712 728
rect 5337 504 5387 560
rect 4748 336 4798 392
rect 3423 168 3473 224
rect 2834 0 2884 56
rect 3423 0 3473 56
rect 2834 -168 2884 -112
rect 3423 -168 3473 -112
rect 4748 168 4798 224
rect 6662 504 6712 560
rect 2834 -336 2884 -280
rect 5337 336 5387 392
rect 6662 336 6712 392
rect 5337 168 5387 224
rect 4748 0 4798 56
rect 5337 0 5387 56
rect 4748 -168 4798 -112
rect 3423 -336 3473 -280
rect 5337 -168 5387 -112
rect 6662 168 6712 224
rect 4748 -336 4798 -280
rect 6662 0 6712 56
rect 6662 -168 6712 -112
rect 5337 -336 5387 -280
rect 6662 -336 6712 -280
<< ndiff >>
rect -100 1504 -28 1517
rect -100 1458 -87 1504
rect -41 1458 -28 1504
rect -100 1445 -28 1458
rect -89 1425 -39 1445
rect -89 1349 -39 1369
rect -100 1336 -28 1349
rect -100 1290 -87 1336
rect -41 1290 -28 1336
rect -100 1277 -28 1290
rect -89 1257 -39 1277
rect -89 1181 -39 1201
rect -100 1168 -28 1181
rect -100 1122 -87 1168
rect -41 1122 -28 1168
rect -100 1109 -28 1122
rect 1828 1498 1900 1511
rect 1828 1452 1841 1498
rect 1887 1452 1900 1498
rect 1828 1439 1900 1452
rect 1839 1419 1889 1439
rect 1839 1343 1889 1363
rect 1828 1330 1900 1343
rect 1828 1284 1841 1330
rect 1887 1284 1900 1330
rect 1828 1271 1900 1284
rect 1839 1251 1889 1271
rect 1839 1175 1889 1195
rect 1828 1162 1900 1175
rect 1828 1116 1841 1162
rect 1887 1116 1900 1162
rect 1828 1103 1900 1116
rect 1828 1028 1900 1041
rect 1828 982 1841 1028
rect 1887 982 1900 1028
rect 1828 969 1900 982
rect 1839 949 1889 969
rect -104 748 -32 761
rect -104 702 -91 748
rect -45 702 -32 748
rect -104 689 -32 702
rect -93 669 -43 689
rect 1839 873 1889 893
rect 1828 860 1900 873
rect 1828 814 1841 860
rect 1887 814 1900 860
rect 1828 801 1900 814
rect 2491 1311 2563 1324
rect 2491 1265 2504 1311
rect 2550 1265 2563 1311
rect 2491 1252 2563 1265
rect 2502 1232 2552 1252
rect 2502 1156 2552 1176
rect 2491 1143 2563 1156
rect 2491 1097 2504 1143
rect 2550 1097 2563 1143
rect 2491 1084 2563 1097
rect 2502 1064 2552 1084
rect 2502 988 2552 1008
rect 2491 975 2563 988
rect 2491 929 2504 975
rect 2550 929 2563 975
rect 2491 916 2563 929
rect 2502 896 2552 916
rect 2502 820 2552 840
rect -93 593 -43 613
rect -104 580 -32 593
rect -104 534 -91 580
rect -45 534 -32 580
rect -104 521 -32 534
rect -93 501 -43 521
rect 2491 807 2563 820
rect 2491 761 2504 807
rect 2550 761 2563 807
rect 2491 748 2563 761
rect 2502 728 2552 748
rect 3744 1311 3816 1324
rect 3744 1265 3757 1311
rect 3803 1265 3816 1311
rect 3744 1252 3816 1265
rect 3755 1232 3805 1252
rect 4405 1311 4477 1324
rect 4405 1265 4418 1311
rect 4464 1265 4477 1311
rect 4405 1252 4477 1265
rect 4416 1232 4466 1252
rect 3755 1156 3805 1176
rect 3744 1143 3816 1156
rect 3744 1097 3757 1143
rect 3803 1097 3816 1143
rect 3744 1084 3816 1097
rect 4416 1156 4466 1176
rect 3755 1064 3805 1084
rect 4405 1143 4477 1156
rect 4405 1097 4418 1143
rect 4464 1097 4477 1143
rect 4405 1084 4477 1097
rect 4416 1064 4466 1084
rect 3755 988 3805 1008
rect 3744 975 3816 988
rect 3744 929 3757 975
rect 3803 929 3816 975
rect 3744 916 3816 929
rect 4416 988 4466 1008
rect 3755 896 3805 916
rect 4405 975 4477 988
rect 4405 929 4418 975
rect 4464 929 4477 975
rect 4405 916 4477 929
rect 4416 896 4466 916
rect 3755 820 3805 840
rect 3744 807 3816 820
rect 3744 761 3757 807
rect 3803 761 3816 807
rect 3744 748 3816 761
rect 4416 820 4466 840
rect 3755 728 3805 748
rect 2502 652 2552 672
rect 1574 565 1646 578
rect -93 425 -43 445
rect -104 412 -32 425
rect -104 366 -91 412
rect -45 366 -32 412
rect -104 353 -32 366
rect 1574 519 1587 565
rect 1633 519 1646 565
rect 1574 506 1646 519
rect 1585 486 1635 506
rect 1585 410 1635 430
rect 1574 397 1646 410
rect 2491 639 2563 652
rect 2491 593 2504 639
rect 2550 593 2563 639
rect 2491 580 2563 593
rect 2502 560 2552 580
rect 4405 807 4477 820
rect 4405 761 4418 807
rect 4464 761 4477 807
rect 4405 748 4477 761
rect 4416 728 4466 748
rect 5658 1311 5730 1324
rect 5658 1265 5671 1311
rect 5717 1265 5730 1311
rect 5658 1252 5730 1265
rect 5669 1232 5719 1252
rect 6319 1311 6391 1324
rect 6319 1265 6332 1311
rect 6378 1265 6391 1311
rect 6319 1252 6391 1265
rect 6330 1232 6380 1252
rect 5669 1156 5719 1176
rect 5658 1143 5730 1156
rect 5658 1097 5671 1143
rect 5717 1097 5730 1143
rect 5658 1084 5730 1097
rect 6330 1156 6380 1176
rect 5669 1064 5719 1084
rect 6319 1143 6391 1156
rect 6319 1097 6332 1143
rect 6378 1097 6391 1143
rect 6319 1084 6391 1097
rect 6330 1064 6380 1084
rect 5669 988 5719 1008
rect 5658 975 5730 988
rect 5658 929 5671 975
rect 5717 929 5730 975
rect 5658 916 5730 929
rect 6330 988 6380 1008
rect 5669 896 5719 916
rect 6319 975 6391 988
rect 6319 929 6332 975
rect 6378 929 6391 975
rect 6319 916 6391 929
rect 6330 896 6380 916
rect 2502 484 2552 504
rect 1574 351 1587 397
rect 1633 351 1646 397
rect 1574 338 1646 351
rect 2491 471 2563 484
rect 2491 425 2504 471
rect 2550 425 2563 471
rect 2491 412 2563 425
rect 2502 392 2552 412
rect 3755 652 3805 672
rect 5669 820 5719 840
rect 5658 807 5730 820
rect 5658 761 5671 807
rect 5717 761 5730 807
rect 5658 748 5730 761
rect 6330 820 6380 840
rect 5669 728 5719 748
rect 3744 639 3816 652
rect 3744 593 3757 639
rect 3803 593 3816 639
rect 3744 580 3816 593
rect 4416 652 4466 672
rect 3755 560 3805 580
rect 4405 639 4477 652
rect 4405 593 4418 639
rect 4464 593 4477 639
rect 4405 580 4477 593
rect 4416 560 4466 580
rect 6319 807 6391 820
rect 6319 761 6332 807
rect 6378 761 6391 807
rect 6319 748 6391 761
rect 6330 728 6380 748
rect 1585 318 1635 338
rect 1585 242 1635 262
rect 1574 229 1646 242
rect 1574 183 1587 229
rect 1633 183 1646 229
rect 1574 170 1646 183
rect 1585 150 1635 170
rect 2502 316 2552 336
rect 2491 303 2563 316
rect 2491 257 2504 303
rect 2550 257 2563 303
rect 2491 244 2563 257
rect 2502 224 2552 244
rect 3755 484 3805 504
rect 3744 471 3816 484
rect 3744 425 3757 471
rect 3803 425 3816 471
rect 3744 412 3816 425
rect 4416 484 4466 504
rect 3755 392 3805 412
rect -104 -7 -32 6
rect -104 -53 -91 -7
rect -45 -53 -32 -7
rect -104 -66 -32 -53
rect -93 -86 -43 -66
rect -93 -162 -43 -142
rect -104 -175 -32 -162
rect -104 -221 -91 -175
rect -45 -221 -32 -175
rect -104 -234 -32 -221
rect -93 -254 -43 -234
rect 1585 74 1635 94
rect 1574 61 1646 74
rect 1574 15 1587 61
rect 1633 15 1646 61
rect 1574 2 1646 15
rect 1585 -18 1635 2
rect -93 -330 -43 -310
rect -104 -343 -32 -330
rect -104 -389 -91 -343
rect -45 -389 -32 -343
rect -104 -402 -32 -389
rect 1585 -94 1635 -74
rect 1574 -107 1646 -94
rect 1574 -153 1587 -107
rect 1633 -153 1646 -107
rect 1574 -166 1646 -153
rect 1574 -304 1646 -291
rect 1574 -350 1587 -304
rect 1633 -350 1646 -304
rect 2502 148 2552 168
rect 4405 471 4477 484
rect 4405 425 4418 471
rect 4464 425 4477 471
rect 4405 412 4477 425
rect 4416 392 4466 412
rect 5669 652 5719 672
rect 5658 639 5730 652
rect 5658 593 5671 639
rect 5717 593 5730 639
rect 5658 580 5730 593
rect 6330 652 6380 672
rect 5669 560 5719 580
rect 6319 639 6391 652
rect 6319 593 6332 639
rect 6378 593 6391 639
rect 6319 580 6391 593
rect 6330 560 6380 580
rect 3755 316 3805 336
rect 3744 303 3816 316
rect 3744 257 3757 303
rect 3803 257 3816 303
rect 3744 244 3816 257
rect 4416 316 4466 336
rect 3755 224 3805 244
rect 4405 303 4477 316
rect 4405 257 4418 303
rect 4464 257 4477 303
rect 4405 244 4477 257
rect 2491 135 2563 148
rect 2491 89 2504 135
rect 2550 89 2563 135
rect 2491 76 2563 89
rect 3755 148 3805 168
rect 2502 56 2552 76
rect 2502 -20 2552 0
rect 3744 135 3816 148
rect 3744 89 3757 135
rect 3803 89 3816 135
rect 3744 76 3816 89
rect 2491 -33 2563 -20
rect 2491 -79 2504 -33
rect 2550 -79 2563 -33
rect 2491 -92 2563 -79
rect 2502 -112 2552 -92
rect 3755 56 3805 76
rect 3755 -20 3805 0
rect 3744 -33 3816 -20
rect 2502 -188 2552 -168
rect 2491 -201 2563 -188
rect 2491 -247 2504 -201
rect 2550 -247 2563 -201
rect 2491 -260 2563 -247
rect 2502 -280 2552 -260
rect 3744 -79 3757 -33
rect 3803 -79 3816 -33
rect 3744 -92 3816 -79
rect 3755 -112 3805 -92
rect 4416 224 4466 244
rect 5669 484 5719 504
rect 5658 471 5730 484
rect 5658 425 5671 471
rect 5717 425 5730 471
rect 5658 412 5730 425
rect 6330 484 6380 504
rect 5669 392 5719 412
rect 1574 -363 1646 -350
rect 3755 -188 3805 -168
rect 4416 148 4466 168
rect 6319 471 6391 484
rect 6319 425 6332 471
rect 6378 425 6391 471
rect 6319 412 6391 425
rect 6330 392 6380 412
rect 5669 316 5719 336
rect 5658 303 5730 316
rect 5658 257 5671 303
rect 5717 257 5730 303
rect 5658 244 5730 257
rect 6330 316 6380 336
rect 5669 224 5719 244
rect 6319 303 6391 316
rect 6319 257 6332 303
rect 6378 257 6391 303
rect 6319 244 6391 257
rect 4405 135 4477 148
rect 4405 89 4418 135
rect 4464 89 4477 135
rect 4405 76 4477 89
rect 5669 148 5719 168
rect 4416 56 4466 76
rect 4416 -20 4466 0
rect 5658 135 5730 148
rect 5658 89 5671 135
rect 5717 89 5730 135
rect 5658 76 5730 89
rect 4405 -33 4477 -20
rect 4405 -79 4418 -33
rect 4464 -79 4477 -33
rect 4405 -92 4477 -79
rect 4416 -112 4466 -92
rect 5669 56 5719 76
rect 5669 -20 5719 0
rect 5658 -33 5730 -20
rect 3744 -201 3816 -188
rect 3744 -247 3757 -201
rect 3803 -247 3816 -201
rect 3744 -260 3816 -247
rect 4416 -188 4466 -168
rect 3755 -280 3805 -260
rect 1585 -383 1635 -363
rect 1585 -459 1635 -439
rect 1574 -472 1646 -459
rect 1574 -518 1587 -472
rect 1633 -518 1646 -472
rect 1574 -531 1646 -518
rect 2502 -356 2552 -336
rect 2491 -369 2563 -356
rect 2491 -415 2504 -369
rect 2550 -415 2563 -369
rect 2491 -428 2563 -415
rect 4405 -201 4477 -188
rect 4405 -247 4418 -201
rect 4464 -247 4477 -201
rect 4405 -260 4477 -247
rect 4416 -280 4466 -260
rect 5658 -79 5671 -33
rect 5717 -79 5730 -33
rect 5658 -92 5730 -79
rect 5669 -112 5719 -92
rect 6330 224 6380 244
rect 5669 -188 5719 -168
rect 6330 148 6380 168
rect 6319 135 6391 148
rect 6319 89 6332 135
rect 6378 89 6391 135
rect 6319 76 6391 89
rect 6330 56 6380 76
rect 6330 -20 6380 0
rect 6319 -33 6391 -20
rect 6319 -79 6332 -33
rect 6378 -79 6391 -33
rect 6319 -92 6391 -79
rect 6330 -112 6380 -92
rect 5658 -201 5730 -188
rect 5658 -247 5671 -201
rect 5717 -247 5730 -201
rect 5658 -260 5730 -247
rect 6330 -188 6380 -168
rect 5669 -280 5719 -260
rect 3755 -356 3805 -336
rect 3744 -369 3816 -356
rect 3744 -415 3757 -369
rect 3803 -415 3816 -369
rect 3744 -428 3816 -415
rect 4416 -356 4466 -336
rect 4405 -369 4477 -356
rect 4405 -415 4418 -369
rect 4464 -415 4477 -369
rect 4405 -428 4477 -415
rect 6319 -201 6391 -188
rect 6319 -247 6332 -201
rect 6378 -247 6391 -201
rect 6319 -260 6391 -247
rect 6330 -280 6380 -260
rect 5669 -356 5719 -336
rect 5658 -369 5730 -356
rect 5658 -415 5671 -369
rect 5717 -415 5730 -369
rect 5658 -428 5730 -415
rect 6330 -356 6380 -336
rect 6319 -369 6391 -356
rect 6319 -415 6332 -369
rect 6378 -415 6391 -369
rect 6319 -428 6391 -415
<< pdiff >>
rect 190 1504 262 1517
rect 190 1458 203 1504
rect 249 1458 262 1504
rect 190 1445 262 1458
rect 201 1425 251 1445
rect 201 1349 251 1369
rect 190 1336 262 1349
rect 190 1290 203 1336
rect 249 1290 262 1336
rect 190 1277 262 1290
rect 201 1257 251 1277
rect 201 1181 251 1201
rect 190 1168 262 1181
rect 190 1122 203 1168
rect 249 1122 262 1168
rect 190 1109 262 1122
rect 1133 1498 1205 1511
rect 1133 1452 1146 1498
rect 1192 1452 1205 1498
rect 1133 1439 1205 1452
rect 1263 1498 1335 1511
rect 1263 1452 1276 1498
rect 1322 1452 1335 1498
rect 1263 1439 1335 1452
rect 1396 1498 1468 1511
rect 1396 1452 1409 1498
rect 1455 1452 1468 1498
rect 1396 1439 1468 1452
rect 1526 1498 1598 1511
rect 1526 1452 1539 1498
rect 1585 1452 1598 1498
rect 1526 1439 1598 1452
rect 1144 1419 1194 1439
rect 1274 1419 1324 1439
rect 1407 1419 1457 1439
rect 1537 1419 1587 1439
rect 1144 1343 1194 1363
rect 1274 1343 1324 1363
rect 1407 1343 1457 1363
rect 1537 1343 1587 1363
rect 1133 1330 1205 1343
rect 1133 1284 1146 1330
rect 1192 1284 1205 1330
rect 1133 1271 1205 1284
rect 1263 1330 1335 1343
rect 1263 1284 1276 1330
rect 1322 1284 1335 1330
rect 1263 1271 1335 1284
rect 1396 1330 1468 1343
rect 1396 1284 1409 1330
rect 1455 1284 1468 1330
rect 1396 1271 1468 1284
rect 1526 1330 1598 1343
rect 1526 1284 1539 1330
rect 1585 1284 1598 1330
rect 1526 1271 1598 1284
rect 1144 1251 1194 1271
rect 1274 1251 1324 1271
rect 1407 1251 1457 1271
rect 1537 1251 1587 1271
rect 1144 1175 1194 1195
rect 1274 1175 1324 1195
rect 1407 1175 1457 1195
rect 1537 1175 1587 1195
rect 1133 1162 1205 1175
rect 1133 1116 1146 1162
rect 1192 1116 1205 1162
rect 1133 1103 1205 1116
rect 1263 1162 1335 1175
rect 1263 1116 1276 1162
rect 1322 1116 1335 1162
rect 1263 1103 1335 1116
rect 1396 1162 1468 1175
rect 1396 1116 1409 1162
rect 1455 1116 1468 1162
rect 1396 1103 1468 1116
rect 1526 1162 1598 1175
rect 1526 1116 1539 1162
rect 1585 1116 1598 1162
rect 1526 1103 1598 1116
rect 1133 1028 1205 1041
rect 1133 982 1146 1028
rect 1192 982 1205 1028
rect 1133 969 1205 982
rect 1396 1028 1468 1041
rect 1396 982 1409 1028
rect 1455 982 1468 1028
rect 1396 969 1468 982
rect 1526 1028 1598 1041
rect 1526 982 1539 1028
rect 1585 982 1598 1028
rect 1526 969 1598 982
rect 1144 949 1194 969
rect 1407 949 1457 969
rect 1537 949 1587 969
rect 186 748 258 761
rect 186 702 199 748
rect 245 702 258 748
rect 186 689 258 702
rect 197 669 247 689
rect 1144 873 1194 893
rect 1407 873 1457 893
rect 1537 873 1587 893
rect 1133 860 1205 873
rect 1133 814 1146 860
rect 1192 814 1205 860
rect 1133 801 1205 814
rect 1396 860 1468 873
rect 1396 814 1409 860
rect 1455 814 1468 860
rect 1396 801 1468 814
rect 1526 860 1598 873
rect 1526 814 1539 860
rect 1585 814 1598 860
rect 1526 801 1598 814
rect 2823 1311 2895 1324
rect 2823 1265 2836 1311
rect 2882 1265 2895 1311
rect 2823 1252 2895 1265
rect 2834 1232 2884 1252
rect 2834 1156 2884 1176
rect 2823 1143 2895 1156
rect 2823 1097 2836 1143
rect 2882 1097 2895 1143
rect 2823 1084 2895 1097
rect 2834 1064 2884 1084
rect 2834 988 2884 1008
rect 2823 975 2895 988
rect 2823 929 2836 975
rect 2882 929 2895 975
rect 2823 916 2895 929
rect 2834 896 2884 916
rect 197 593 247 613
rect 186 580 258 593
rect 186 534 199 580
rect 245 534 258 580
rect 186 521 258 534
rect 2834 820 2884 840
rect 2823 807 2895 820
rect 2823 761 2836 807
rect 2882 761 2895 807
rect 2823 748 2895 761
rect 3412 1311 3484 1324
rect 3412 1265 3425 1311
rect 3471 1265 3484 1311
rect 3412 1252 3484 1265
rect 3423 1232 3473 1252
rect 4737 1311 4809 1324
rect 3423 1156 3473 1176
rect 3412 1143 3484 1156
rect 3412 1097 3425 1143
rect 3471 1097 3484 1143
rect 3412 1084 3484 1097
rect 3423 1064 3473 1084
rect 4737 1265 4750 1311
rect 4796 1265 4809 1311
rect 4737 1252 4809 1265
rect 4748 1232 4798 1252
rect 3423 988 3473 1008
rect 3412 975 3484 988
rect 3412 929 3425 975
rect 3471 929 3484 975
rect 3412 916 3484 929
rect 3423 896 3473 916
rect 4748 1156 4798 1176
rect 4737 1143 4809 1156
rect 4737 1097 4750 1143
rect 4796 1097 4809 1143
rect 4737 1084 4809 1097
rect 4748 1064 4798 1084
rect 4748 988 4798 1008
rect 4737 975 4809 988
rect 4737 929 4750 975
rect 4796 929 4809 975
rect 4737 916 4809 929
rect 4748 896 4798 916
rect 3423 820 3473 840
rect 2834 728 2884 748
rect 3412 807 3484 820
rect 3412 761 3425 807
rect 3471 761 3484 807
rect 3412 748 3484 761
rect 3423 728 3473 748
rect 197 501 247 521
rect 197 425 247 445
rect 186 412 258 425
rect 186 366 199 412
rect 245 366 258 412
rect 186 353 258 366
rect 1175 393 1275 406
rect 1175 347 1188 393
rect 1262 347 1275 393
rect 1175 318 1275 347
rect 2834 652 2884 672
rect 4748 820 4798 840
rect 4737 807 4809 820
rect 4737 761 4750 807
rect 4796 761 4809 807
rect 4737 748 4809 761
rect 5326 1311 5398 1324
rect 5326 1265 5339 1311
rect 5385 1265 5398 1311
rect 5326 1252 5398 1265
rect 5337 1232 5387 1252
rect 6651 1311 6723 1324
rect 5337 1156 5387 1176
rect 5326 1143 5398 1156
rect 5326 1097 5339 1143
rect 5385 1097 5398 1143
rect 5326 1084 5398 1097
rect 5337 1064 5387 1084
rect 6651 1265 6664 1311
rect 6710 1265 6723 1311
rect 6651 1252 6723 1265
rect 6662 1232 6712 1252
rect 5337 988 5387 1008
rect 5326 975 5398 988
rect 5326 929 5339 975
rect 5385 929 5398 975
rect 5326 916 5398 929
rect 5337 896 5387 916
rect 6662 1156 6712 1176
rect 6651 1143 6723 1156
rect 6651 1097 6664 1143
rect 6710 1097 6723 1143
rect 6651 1084 6723 1097
rect 6662 1064 6712 1084
rect 6662 988 6712 1008
rect 6651 975 6723 988
rect 6651 929 6664 975
rect 6710 929 6723 975
rect 6651 916 6723 929
rect 6662 896 6712 916
rect 5337 820 5387 840
rect 4748 728 4798 748
rect 2823 639 2895 652
rect 2823 593 2836 639
rect 2882 593 2895 639
rect 2823 580 2895 593
rect 3423 652 3473 672
rect 2834 560 2884 580
rect 2834 484 2884 504
rect 3412 639 3484 652
rect 3412 593 3425 639
rect 3471 593 3484 639
rect 3412 580 3484 593
rect 3423 560 3473 580
rect 5326 807 5398 820
rect 5326 761 5339 807
rect 5385 761 5398 807
rect 5326 748 5398 761
rect 5337 728 5387 748
rect 4748 652 4798 672
rect 6662 820 6712 840
rect 6651 807 6723 820
rect 6651 761 6664 807
rect 6710 761 6723 807
rect 6651 748 6723 761
rect 6662 728 6712 748
rect 4737 639 4809 652
rect 4737 593 4750 639
rect 4796 593 4809 639
rect 4737 580 4809 593
rect 5337 652 5387 672
rect 4748 560 4798 580
rect 2823 471 2895 484
rect 2823 425 2836 471
rect 2882 425 2895 471
rect 2823 412 2895 425
rect 3423 484 3473 504
rect 2834 392 2884 412
rect 1175 233 1275 262
rect 1175 187 1188 233
rect 1262 187 1275 233
rect 1175 158 1275 187
rect 2834 316 2884 336
rect 2823 303 2895 316
rect 2823 257 2836 303
rect 2882 257 2895 303
rect 2823 244 2895 257
rect 2834 224 2884 244
rect 3412 471 3484 484
rect 3412 425 3425 471
rect 3471 425 3484 471
rect 3412 412 3484 425
rect 3423 392 3473 412
rect 1175 73 1275 102
rect 186 -7 258 6
rect 186 -53 199 -7
rect 245 -53 258 -7
rect 186 -66 258 -53
rect 197 -86 247 -66
rect 1175 27 1188 73
rect 1262 27 1275 73
rect 1175 -2 1275 27
rect 197 -162 247 -142
rect 186 -175 258 -162
rect 186 -221 199 -175
rect 245 -221 258 -175
rect 186 -234 258 -221
rect 1175 -87 1275 -58
rect 1175 -133 1188 -87
rect 1262 -133 1275 -87
rect 1175 -146 1275 -133
rect 197 -254 247 -234
rect 197 -330 247 -310
rect 186 -343 258 -330
rect 186 -389 199 -343
rect 245 -389 258 -343
rect 186 -402 258 -389
rect 2834 148 2884 168
rect 4748 484 4798 504
rect 5326 639 5398 652
rect 5326 593 5339 639
rect 5385 593 5398 639
rect 5326 580 5398 593
rect 5337 560 5387 580
rect 6662 652 6712 672
rect 6651 639 6723 652
rect 6651 593 6664 639
rect 6710 593 6723 639
rect 6651 580 6723 593
rect 6662 560 6712 580
rect 4737 471 4809 484
rect 4737 425 4750 471
rect 4796 425 4809 471
rect 4737 412 4809 425
rect 5337 484 5387 504
rect 4748 392 4798 412
rect 3423 316 3473 336
rect 3412 303 3484 316
rect 3412 257 3425 303
rect 3471 257 3484 303
rect 3412 244 3484 257
rect 4748 316 4798 336
rect 3423 224 3473 244
rect 4737 303 4809 316
rect 4737 257 4750 303
rect 4796 257 4809 303
rect 4737 244 4809 257
rect 2823 135 2895 148
rect 2823 89 2836 135
rect 2882 89 2895 135
rect 2823 76 2895 89
rect 3423 148 3473 168
rect 2834 56 2884 76
rect 2834 -20 2884 0
rect 3412 135 3484 148
rect 3412 89 3425 135
rect 3471 89 3484 135
rect 3412 76 3484 89
rect 2823 -33 2895 -20
rect 2823 -79 2836 -33
rect 2882 -79 2895 -33
rect 2823 -92 2895 -79
rect 3423 56 3473 76
rect 3423 -20 3473 0
rect 2834 -112 2884 -92
rect 3412 -33 3484 -20
rect 3412 -79 3425 -33
rect 3471 -79 3484 -33
rect 3412 -92 3484 -79
rect 3423 -112 3473 -92
rect 2834 -188 2884 -168
rect 4748 224 4798 244
rect 5326 471 5398 484
rect 5326 425 5339 471
rect 5385 425 5398 471
rect 5326 412 5398 425
rect 5337 392 5387 412
rect 2823 -201 2895 -188
rect 2823 -247 2836 -201
rect 2882 -247 2895 -201
rect 2823 -260 2895 -247
rect 3423 -188 3473 -168
rect 2834 -280 2884 -260
rect 3412 -201 3484 -188
rect 3412 -247 3425 -201
rect 3471 -247 3484 -201
rect 3412 -260 3484 -247
rect 3423 -280 3473 -260
rect 4748 148 4798 168
rect 6662 484 6712 504
rect 6651 471 6723 484
rect 6651 425 6664 471
rect 6710 425 6723 471
rect 6651 412 6723 425
rect 6662 392 6712 412
rect 5337 316 5387 336
rect 5326 303 5398 316
rect 5326 257 5339 303
rect 5385 257 5398 303
rect 5326 244 5398 257
rect 6662 316 6712 336
rect 5337 224 5387 244
rect 6651 303 6723 316
rect 6651 257 6664 303
rect 6710 257 6723 303
rect 6651 244 6723 257
rect 4737 135 4809 148
rect 4737 89 4750 135
rect 4796 89 4809 135
rect 4737 76 4809 89
rect 5337 148 5387 168
rect 4748 56 4798 76
rect 4748 -20 4798 0
rect 5326 135 5398 148
rect 5326 89 5339 135
rect 5385 89 5398 135
rect 5326 76 5398 89
rect 4737 -33 4809 -20
rect 4737 -79 4750 -33
rect 4796 -79 4809 -33
rect 4737 -92 4809 -79
rect 5337 56 5387 76
rect 5337 -20 5387 0
rect 4748 -112 4798 -92
rect 5326 -33 5398 -20
rect 5326 -79 5339 -33
rect 5385 -79 5398 -33
rect 5326 -92 5398 -79
rect 5337 -112 5387 -92
rect 2834 -356 2884 -336
rect 2823 -369 2895 -356
rect 2823 -415 2836 -369
rect 2882 -415 2895 -369
rect 2823 -428 2895 -415
rect 4748 -188 4798 -168
rect 6662 224 6712 244
rect 4737 -201 4809 -188
rect 4737 -247 4750 -201
rect 4796 -247 4809 -201
rect 4737 -260 4809 -247
rect 5337 -188 5387 -168
rect 4748 -280 4798 -260
rect 5326 -201 5398 -188
rect 5326 -247 5339 -201
rect 5385 -247 5398 -201
rect 5326 -260 5398 -247
rect 5337 -280 5387 -260
rect 6662 148 6712 168
rect 6651 135 6723 148
rect 6651 89 6664 135
rect 6710 89 6723 135
rect 6651 76 6723 89
rect 6662 56 6712 76
rect 6662 -20 6712 0
rect 6651 -33 6723 -20
rect 6651 -79 6664 -33
rect 6710 -79 6723 -33
rect 6651 -92 6723 -79
rect 6662 -112 6712 -92
rect 3423 -356 3473 -336
rect 3412 -369 3484 -356
rect 3412 -415 3425 -369
rect 3471 -415 3484 -369
rect 3412 -428 3484 -415
rect 4748 -356 4798 -336
rect 4737 -369 4809 -356
rect 4737 -415 4750 -369
rect 4796 -415 4809 -369
rect 4737 -428 4809 -415
rect 6662 -188 6712 -168
rect 6651 -201 6723 -188
rect 6651 -247 6664 -201
rect 6710 -247 6723 -201
rect 6651 -260 6723 -247
rect 6662 -280 6712 -260
rect 5337 -356 5387 -336
rect 5326 -369 5398 -356
rect 5326 -415 5339 -369
rect 5385 -415 5398 -369
rect 5326 -428 5398 -415
rect 6662 -356 6712 -336
rect 6651 -369 6723 -356
rect 6651 -415 6664 -369
rect 6710 -415 6723 -369
rect 6651 -428 6723 -415
<< ndiffc >>
rect -87 1458 -41 1504
rect -87 1290 -41 1336
rect -87 1122 -41 1168
rect 1841 1452 1887 1498
rect 1841 1284 1887 1330
rect 1841 1116 1887 1162
rect 1841 982 1887 1028
rect -91 702 -45 748
rect 1841 814 1887 860
rect 2504 1265 2550 1311
rect 2504 1097 2550 1143
rect 2504 929 2550 975
rect -91 534 -45 580
rect 2504 761 2550 807
rect 3757 1265 3803 1311
rect 4418 1265 4464 1311
rect 3757 1097 3803 1143
rect 4418 1097 4464 1143
rect 3757 929 3803 975
rect 4418 929 4464 975
rect 3757 761 3803 807
rect -91 366 -45 412
rect 1587 519 1633 565
rect 2504 593 2550 639
rect 4418 761 4464 807
rect 5671 1265 5717 1311
rect 6332 1265 6378 1311
rect 5671 1097 5717 1143
rect 6332 1097 6378 1143
rect 5671 929 5717 975
rect 6332 929 6378 975
rect 1587 351 1633 397
rect 2504 425 2550 471
rect 5671 761 5717 807
rect 3757 593 3803 639
rect 4418 593 4464 639
rect 6332 761 6378 807
rect 1587 183 1633 229
rect 2504 257 2550 303
rect 3757 425 3803 471
rect -91 -53 -45 -7
rect -91 -221 -45 -175
rect 1587 15 1633 61
rect -91 -389 -45 -343
rect 1587 -153 1633 -107
rect 1587 -350 1633 -304
rect 4418 425 4464 471
rect 5671 593 5717 639
rect 6332 593 6378 639
rect 3757 257 3803 303
rect 4418 257 4464 303
rect 2504 89 2550 135
rect 3757 89 3803 135
rect 2504 -79 2550 -33
rect 2504 -247 2550 -201
rect 3757 -79 3803 -33
rect 5671 425 5717 471
rect 6332 425 6378 471
rect 5671 257 5717 303
rect 6332 257 6378 303
rect 4418 89 4464 135
rect 5671 89 5717 135
rect 4418 -79 4464 -33
rect 3757 -247 3803 -201
rect 1587 -518 1633 -472
rect 2504 -415 2550 -369
rect 4418 -247 4464 -201
rect 5671 -79 5717 -33
rect 6332 89 6378 135
rect 6332 -79 6378 -33
rect 5671 -247 5717 -201
rect 3757 -415 3803 -369
rect 4418 -415 4464 -369
rect 6332 -247 6378 -201
rect 5671 -415 5717 -369
rect 6332 -415 6378 -369
<< pdiffc >>
rect 203 1458 249 1504
rect 203 1290 249 1336
rect 203 1122 249 1168
rect 1146 1452 1192 1498
rect 1276 1452 1322 1498
rect 1409 1452 1455 1498
rect 1539 1452 1585 1498
rect 1146 1284 1192 1330
rect 1276 1284 1322 1330
rect 1409 1284 1455 1330
rect 1539 1284 1585 1330
rect 1146 1116 1192 1162
rect 1276 1116 1322 1162
rect 1409 1116 1455 1162
rect 1539 1116 1585 1162
rect 1146 982 1192 1028
rect 1409 982 1455 1028
rect 1539 982 1585 1028
rect 199 702 245 748
rect 1146 814 1192 860
rect 1409 814 1455 860
rect 1539 814 1585 860
rect 2836 1265 2882 1311
rect 2836 1097 2882 1143
rect 2836 929 2882 975
rect 199 534 245 580
rect 2836 761 2882 807
rect 3425 1265 3471 1311
rect 3425 1097 3471 1143
rect 4750 1265 4796 1311
rect 3425 929 3471 975
rect 4750 1097 4796 1143
rect 4750 929 4796 975
rect 3425 761 3471 807
rect 199 366 245 412
rect 1188 347 1262 393
rect 4750 761 4796 807
rect 5339 1265 5385 1311
rect 5339 1097 5385 1143
rect 6664 1265 6710 1311
rect 5339 929 5385 975
rect 6664 1097 6710 1143
rect 6664 929 6710 975
rect 2836 593 2882 639
rect 3425 593 3471 639
rect 5339 761 5385 807
rect 6664 761 6710 807
rect 4750 593 4796 639
rect 2836 425 2882 471
rect 1188 187 1262 233
rect 2836 257 2882 303
rect 3425 425 3471 471
rect 199 -53 245 -7
rect 1188 27 1262 73
rect 199 -221 245 -175
rect 1188 -133 1262 -87
rect 199 -389 245 -343
rect 5339 593 5385 639
rect 6664 593 6710 639
rect 4750 425 4796 471
rect 3425 257 3471 303
rect 4750 257 4796 303
rect 2836 89 2882 135
rect 3425 89 3471 135
rect 2836 -79 2882 -33
rect 3425 -79 3471 -33
rect 5339 425 5385 471
rect 2836 -247 2882 -201
rect 3425 -247 3471 -201
rect 6664 425 6710 471
rect 5339 257 5385 303
rect 6664 257 6710 303
rect 4750 89 4796 135
rect 5339 89 5385 135
rect 4750 -79 4796 -33
rect 5339 -79 5385 -33
rect 2836 -415 2882 -369
rect 4750 -247 4796 -201
rect 5339 -247 5385 -201
rect 6664 89 6710 135
rect 6664 -79 6710 -33
rect 3425 -415 3471 -369
rect 4750 -415 4796 -369
rect 6664 -247 6710 -201
rect 5339 -415 5385 -369
rect 6664 -415 6710 -369
<< psubdiff >>
rect -318 1564 -246 1577
rect -318 1518 -305 1564
rect -259 1518 -246 1564
rect -318 1453 -246 1518
rect -318 1407 -305 1453
rect -259 1407 -246 1453
rect -318 1342 -246 1407
rect -318 1296 -305 1342
rect -259 1296 -246 1342
rect -318 1231 -246 1296
rect -318 1185 -305 1231
rect -259 1185 -246 1231
rect -318 1120 -246 1185
rect -318 1074 -305 1120
rect -259 1074 -246 1120
rect -318 1049 -246 1074
rect 1998 1553 2084 1569
rect 1998 1498 2013 1553
rect 2068 1498 2084 1553
rect 1998 1430 2084 1498
rect 1998 1375 2013 1430
rect 2068 1375 2084 1430
rect 1998 1307 2084 1375
rect 1998 1252 2013 1307
rect 2068 1252 2084 1307
rect 1998 1184 2084 1252
rect 1998 1129 2013 1184
rect 2068 1129 2084 1184
rect 1998 1061 2084 1129
rect 1998 1006 2013 1061
rect 2068 1006 2084 1061
rect 1998 938 2084 1006
rect -322 808 -250 821
rect -322 762 -309 808
rect -263 762 -250 808
rect -322 697 -250 762
rect -322 651 -309 697
rect -263 651 -250 697
rect -322 586 -250 651
rect 1998 883 2013 938
rect 2068 883 2084 938
rect 1998 815 2084 883
rect 1998 760 2013 815
rect 2068 760 2084 815
rect 1998 743 2084 760
rect 2160 1366 2234 1379
rect 2160 1314 2173 1366
rect 2220 1314 2234 1366
rect 2160 1256 2234 1314
rect 2160 1204 2173 1256
rect 2220 1204 2234 1256
rect 2160 1146 2234 1204
rect 2160 1094 2173 1146
rect 2220 1094 2234 1146
rect 2160 1036 2234 1094
rect 2160 984 2173 1036
rect 2220 984 2234 1036
rect 2160 926 2234 984
rect 2160 874 2173 926
rect 2220 874 2234 926
rect 2160 816 2234 874
rect 2160 764 2173 816
rect 2220 764 2234 816
rect -322 540 -309 586
rect -263 540 -250 586
rect -322 475 -250 540
rect 2160 706 2234 764
rect 4073 1366 4148 1379
rect 4073 1314 4087 1366
rect 4134 1314 4148 1366
rect 4073 1256 4148 1314
rect 4073 1204 4087 1256
rect 4134 1204 4148 1256
rect 4073 1146 4148 1204
rect 4073 1094 4087 1146
rect 4134 1094 4148 1146
rect 4073 1036 4148 1094
rect 4073 984 4087 1036
rect 4134 984 4148 1036
rect 4073 926 4148 984
rect 4073 874 4087 926
rect 4134 874 4148 926
rect 2160 654 2173 706
rect 2220 654 2234 706
rect 4073 816 4148 874
rect 4073 764 4087 816
rect 4134 764 4148 816
rect 2160 596 2234 654
rect -322 429 -309 475
rect -263 429 -250 475
rect -322 364 -250 429
rect -322 318 -309 364
rect -263 318 -250 364
rect -322 293 -250 318
rect 1790 551 1879 568
rect 1790 422 1805 551
rect 1864 422 1879 551
rect 1790 405 1879 422
rect 2160 544 2173 596
rect 2220 544 2234 596
rect 4073 706 4148 764
rect 5987 1366 6062 1379
rect 5987 1314 6001 1366
rect 6048 1314 6062 1366
rect 5987 1256 6062 1314
rect 5987 1204 6001 1256
rect 6048 1204 6062 1256
rect 5987 1146 6062 1204
rect 5987 1094 6001 1146
rect 6048 1094 6062 1146
rect 5987 1036 6062 1094
rect 5987 984 6001 1036
rect 6048 984 6062 1036
rect 5987 926 6062 984
rect 5987 874 6001 926
rect 6048 874 6062 926
rect 2160 486 2234 544
rect 2160 434 2173 486
rect 2220 434 2234 486
rect 2160 376 2234 434
rect 4073 654 4087 706
rect 4134 654 4148 706
rect 5987 816 6062 874
rect 5987 764 6001 816
rect 6048 764 6062 816
rect 4073 596 4148 654
rect 4073 544 4087 596
rect 4134 544 4148 596
rect 5987 706 6062 764
rect 2160 324 2173 376
rect 2220 324 2234 376
rect 1784 306 1873 323
rect 1784 177 1799 306
rect 1858 177 1873 306
rect 1784 160 1873 177
rect 2160 266 2234 324
rect 2160 214 2173 266
rect 2220 214 2234 266
rect 2160 156 2234 214
rect 4073 486 4148 544
rect 4073 434 4087 486
rect 4134 434 4148 486
rect -322 53 -250 66
rect -322 7 -309 53
rect -263 7 -250 53
rect -322 -58 -250 7
rect -322 -104 -309 -58
rect -263 -104 -250 -58
rect -322 -169 -250 -104
rect 2160 104 2173 156
rect 2220 104 2234 156
rect -322 -215 -309 -169
rect -263 -215 -250 -169
rect -322 -280 -250 -215
rect 1787 74 1876 91
rect -322 -326 -309 -280
rect -263 -326 -250 -280
rect -322 -391 -250 -326
rect -322 -437 -309 -391
rect -263 -437 -250 -391
rect -322 -462 -250 -437
rect 1787 -55 1802 74
rect 1861 -55 1876 74
rect 1787 -72 1876 -55
rect 2160 46 2234 104
rect 2160 -6 2173 46
rect 2220 -6 2234 46
rect 2160 -64 2234 -6
rect 2160 -116 2173 -64
rect 2220 -116 2234 -64
rect 1788 -173 1877 -156
rect 1788 -302 1803 -173
rect 1862 -302 1877 -173
rect 1788 -319 1877 -302
rect 2160 -174 2234 -116
rect 4073 376 4148 434
rect 5987 654 6001 706
rect 6048 654 6062 706
rect 5987 596 6062 654
rect 5987 544 6001 596
rect 6048 544 6062 596
rect 4073 324 4087 376
rect 4134 324 4148 376
rect 4073 266 4148 324
rect 4073 214 4087 266
rect 4134 214 4148 266
rect 2160 -226 2173 -174
rect 2220 -226 2234 -174
rect 2160 -284 2234 -226
rect 4073 156 4148 214
rect 5987 486 6062 544
rect 5987 434 6001 486
rect 6048 434 6062 486
rect 4073 104 4087 156
rect 4134 104 4148 156
rect 4073 46 4148 104
rect 4073 -6 4087 46
rect 4134 -6 4148 46
rect 4073 -64 4148 -6
rect 4073 -116 4087 -64
rect 4134 -116 4148 -64
rect 2160 -336 2173 -284
rect 2220 -336 2234 -284
rect 4073 -174 4148 -116
rect 5987 376 6062 434
rect 5987 324 6001 376
rect 6048 324 6062 376
rect 5987 266 6062 324
rect 5987 214 6001 266
rect 6048 214 6062 266
rect 4073 -226 4087 -174
rect 4134 -226 4148 -174
rect 1788 -397 1877 -380
rect 1788 -526 1803 -397
rect 1862 -526 1877 -397
rect 2160 -394 2234 -336
rect 2160 -446 2173 -394
rect 2220 -446 2234 -394
rect 4073 -284 4148 -226
rect 5987 156 6062 214
rect 5987 104 6001 156
rect 6048 104 6062 156
rect 5987 46 6062 104
rect 5987 -6 6001 46
rect 6048 -6 6062 46
rect 5987 -64 6062 -6
rect 5987 -116 6001 -64
rect 6048 -116 6062 -64
rect 4073 -336 4087 -284
rect 4134 -336 4148 -284
rect 5987 -174 6062 -116
rect 5987 -226 6001 -174
rect 6048 -226 6062 -174
rect 2160 -474 2234 -446
rect 4073 -394 4148 -336
rect 4073 -446 4087 -394
rect 4134 -446 4148 -394
rect 5987 -284 6062 -226
rect 5987 -336 6001 -284
rect 6048 -336 6062 -284
rect 4073 -474 4148 -446
rect 5987 -394 6062 -336
rect 5987 -446 6001 -394
rect 6048 -446 6062 -394
rect 5987 -474 6062 -446
rect 1788 -543 1877 -526
<< nsubdiff >>
rect 437 1564 509 1577
rect 437 1518 450 1564
rect 496 1518 509 1564
rect 437 1453 509 1518
rect 437 1407 450 1453
rect 496 1407 509 1453
rect 437 1342 509 1407
rect 437 1296 450 1342
rect 496 1296 509 1342
rect 437 1231 509 1296
rect 437 1185 450 1231
rect 496 1185 509 1231
rect 437 1120 509 1185
rect 437 1074 450 1120
rect 496 1074 509 1120
rect 437 1049 509 1074
rect 874 1553 960 1569
rect 874 1498 889 1553
rect 944 1498 960 1553
rect 874 1430 960 1498
rect 874 1375 889 1430
rect 944 1375 960 1430
rect 874 1307 960 1375
rect 874 1252 889 1307
rect 944 1252 960 1307
rect 874 1184 960 1252
rect 874 1129 889 1184
rect 944 1129 960 1184
rect 874 1061 960 1129
rect 874 1006 889 1061
rect 944 1006 960 1061
rect 874 938 960 1006
rect 874 883 889 938
rect 944 883 960 938
rect 433 808 505 821
rect 433 762 446 808
rect 492 762 505 808
rect 433 697 505 762
rect 874 815 960 883
rect 874 760 889 815
rect 944 760 960 815
rect 874 743 960 760
rect 3114 1366 3193 1380
rect 3114 1315 3128 1366
rect 3179 1315 3193 1366
rect 3114 1256 3193 1315
rect 3114 1205 3128 1256
rect 3179 1205 3193 1256
rect 3114 1146 3193 1205
rect 3114 1095 3128 1146
rect 3179 1095 3193 1146
rect 3114 1036 3193 1095
rect 3114 985 3128 1036
rect 3179 985 3193 1036
rect 3114 926 3193 985
rect 3114 875 3128 926
rect 3179 875 3193 926
rect 433 651 446 697
rect 492 651 505 697
rect 433 586 505 651
rect 433 540 446 586
rect 492 540 505 586
rect 3114 816 3193 875
rect 3114 765 3128 816
rect 3179 765 3193 816
rect 3114 706 3193 765
rect 5028 1366 5107 1380
rect 5028 1315 5042 1366
rect 5093 1315 5107 1366
rect 5028 1256 5107 1315
rect 5028 1205 5042 1256
rect 5093 1205 5107 1256
rect 5028 1146 5107 1205
rect 5028 1095 5042 1146
rect 5093 1095 5107 1146
rect 5028 1036 5107 1095
rect 5028 985 5042 1036
rect 5093 985 5107 1036
rect 5028 926 5107 985
rect 5028 875 5042 926
rect 5093 875 5107 926
rect 433 475 505 540
rect 433 429 446 475
rect 492 429 505 475
rect 433 364 505 429
rect 433 318 446 364
rect 492 318 505 364
rect 433 293 505 318
rect 876 440 958 456
rect 876 324 891 440
rect 942 324 958 440
rect 876 311 958 324
rect 873 189 954 205
rect 873 73 889 189
rect 940 73 954 189
rect 3114 655 3128 706
rect 3179 655 3193 706
rect 5028 816 5107 875
rect 5028 765 5042 816
rect 5093 765 5107 816
rect 3114 596 3193 655
rect 3114 545 3128 596
rect 3179 545 3193 596
rect 3114 486 3193 545
rect 5028 706 5107 765
rect 6942 1366 7020 1380
rect 6942 1315 6956 1366
rect 7007 1315 7020 1366
rect 6942 1256 7020 1315
rect 6942 1205 6956 1256
rect 7007 1205 7020 1256
rect 6942 1146 7020 1205
rect 6942 1095 6956 1146
rect 7007 1095 7020 1146
rect 6942 1036 7020 1095
rect 6942 985 6956 1036
rect 7007 985 7020 1036
rect 6942 926 7020 985
rect 6942 875 6956 926
rect 7007 875 7020 926
rect 5028 655 5042 706
rect 5093 655 5107 706
rect 6942 816 7020 875
rect 6942 765 6956 816
rect 7007 765 7020 816
rect 5028 596 5107 655
rect 3114 435 3128 486
rect 3179 435 3193 486
rect 3114 376 3193 435
rect 3114 325 3128 376
rect 3179 325 3193 376
rect 3114 266 3193 325
rect 3114 215 3128 266
rect 3179 215 3193 266
rect 433 53 505 66
rect 873 60 954 73
rect 433 7 446 53
rect 492 7 505 53
rect 433 -58 505 7
rect 433 -104 446 -58
rect 492 -104 505 -58
rect 433 -169 505 -104
rect 433 -215 446 -169
rect 492 -215 505 -169
rect 875 -51 956 -35
rect 875 -167 890 -51
rect 941 -167 956 -51
rect 875 -180 956 -167
rect 433 -280 505 -215
rect 433 -326 446 -280
rect 492 -326 505 -280
rect 433 -391 505 -326
rect 433 -437 446 -391
rect 492 -437 505 -391
rect 433 -462 505 -437
rect 3114 156 3193 215
rect 5028 545 5042 596
rect 5093 545 5107 596
rect 5028 486 5107 545
rect 6942 706 7020 765
rect 6942 655 6956 706
rect 7007 655 7020 706
rect 6942 596 7020 655
rect 5028 435 5042 486
rect 5093 435 5107 486
rect 3114 105 3128 156
rect 3179 105 3193 156
rect 3114 46 3193 105
rect 3114 -5 3128 46
rect 3179 -5 3193 46
rect 3114 -64 3193 -5
rect 3114 -115 3128 -64
rect 3179 -115 3193 -64
rect 3114 -174 3193 -115
rect 5028 376 5107 435
rect 5028 325 5042 376
rect 5093 325 5107 376
rect 5028 266 5107 325
rect 5028 215 5042 266
rect 5093 215 5107 266
rect 3114 -225 3128 -174
rect 3179 -225 3193 -174
rect 3114 -284 3193 -225
rect 5028 156 5107 215
rect 6942 545 6956 596
rect 7007 545 7020 596
rect 6942 486 7020 545
rect 6942 435 6956 486
rect 7007 435 7020 486
rect 5028 105 5042 156
rect 5093 105 5107 156
rect 5028 46 5107 105
rect 5028 -5 5042 46
rect 5093 -5 5107 46
rect 5028 -64 5107 -5
rect 5028 -115 5042 -64
rect 5093 -115 5107 -64
rect 3114 -335 3128 -284
rect 3179 -335 3193 -284
rect 3114 -394 3193 -335
rect 5028 -174 5107 -115
rect 6942 376 7020 435
rect 6942 325 6956 376
rect 7007 325 7020 376
rect 6942 266 7020 325
rect 6942 215 6956 266
rect 7007 215 7020 266
rect 5028 -225 5042 -174
rect 5093 -225 5107 -174
rect 5028 -284 5107 -225
rect 6942 156 7020 215
rect 6942 105 6956 156
rect 7007 105 7020 156
rect 6942 46 7020 105
rect 6942 -5 6956 46
rect 7007 -5 7020 46
rect 6942 -64 7020 -5
rect 6942 -115 6956 -64
rect 7007 -115 7020 -64
rect 5028 -335 5042 -284
rect 5093 -335 5107 -284
rect 3114 -445 3128 -394
rect 3179 -445 3193 -394
rect 3114 -477 3193 -445
rect 5028 -394 5107 -335
rect 6942 -174 7020 -115
rect 6942 -225 6956 -174
rect 7007 -225 7020 -174
rect 6942 -284 7020 -225
rect 6942 -335 6956 -284
rect 7007 -335 7020 -284
rect 5028 -445 5042 -394
rect 5093 -445 5107 -394
rect 5028 -477 5107 -445
rect 6942 -394 7020 -335
rect 6942 -445 6956 -394
rect 7007 -445 7020 -394
rect 6942 -477 7020 -445
<< psubdiffcont >>
rect -305 1518 -259 1564
rect -305 1407 -259 1453
rect -305 1296 -259 1342
rect -305 1185 -259 1231
rect -305 1074 -259 1120
rect 2013 1498 2068 1553
rect 2013 1375 2068 1430
rect 2013 1252 2068 1307
rect 2013 1129 2068 1184
rect 2013 1006 2068 1061
rect -309 762 -263 808
rect -309 651 -263 697
rect 2013 883 2068 938
rect 2013 760 2068 815
rect 2173 1314 2220 1366
rect 2173 1204 2220 1256
rect 2173 1094 2220 1146
rect 2173 984 2220 1036
rect 2173 874 2220 926
rect 2173 764 2220 816
rect -309 540 -263 586
rect 4087 1314 4134 1366
rect 4087 1204 4134 1256
rect 4087 1094 4134 1146
rect 4087 984 4134 1036
rect 4087 874 4134 926
rect 2173 654 2220 706
rect 4087 764 4134 816
rect -309 429 -263 475
rect -309 318 -263 364
rect 1805 422 1864 551
rect 2173 544 2220 596
rect 6001 1314 6048 1366
rect 6001 1204 6048 1256
rect 6001 1094 6048 1146
rect 6001 984 6048 1036
rect 6001 874 6048 926
rect 2173 434 2220 486
rect 4087 654 4134 706
rect 6001 764 6048 816
rect 4087 544 4134 596
rect 2173 324 2220 376
rect 1799 177 1858 306
rect 2173 214 2220 266
rect 4087 434 4134 486
rect -309 7 -263 53
rect -309 -104 -263 -58
rect 2173 104 2220 156
rect -309 -215 -263 -169
rect -309 -326 -263 -280
rect -309 -437 -263 -391
rect 1802 -55 1861 74
rect 2173 -6 2220 46
rect 2173 -116 2220 -64
rect 1803 -302 1862 -173
rect 6001 654 6048 706
rect 6001 544 6048 596
rect 4087 324 4134 376
rect 4087 214 4134 266
rect 2173 -226 2220 -174
rect 6001 434 6048 486
rect 4087 104 4134 156
rect 4087 -6 4134 46
rect 4087 -116 4134 -64
rect 2173 -336 2220 -284
rect 6001 324 6048 376
rect 6001 214 6048 266
rect 4087 -226 4134 -174
rect 1803 -526 1862 -397
rect 2173 -446 2220 -394
rect 6001 104 6048 156
rect 6001 -6 6048 46
rect 6001 -116 6048 -64
rect 4087 -336 4134 -284
rect 6001 -226 6048 -174
rect 4087 -446 4134 -394
rect 6001 -336 6048 -284
rect 6001 -446 6048 -394
<< nsubdiffcont >>
rect 450 1518 496 1564
rect 450 1407 496 1453
rect 450 1296 496 1342
rect 450 1185 496 1231
rect 450 1074 496 1120
rect 889 1498 944 1553
rect 889 1375 944 1430
rect 889 1252 944 1307
rect 889 1129 944 1184
rect 889 1006 944 1061
rect 889 883 944 938
rect 446 762 492 808
rect 889 760 944 815
rect 3128 1315 3179 1366
rect 3128 1205 3179 1256
rect 3128 1095 3179 1146
rect 3128 985 3179 1036
rect 3128 875 3179 926
rect 446 651 492 697
rect 446 540 492 586
rect 3128 765 3179 816
rect 5042 1315 5093 1366
rect 5042 1205 5093 1256
rect 5042 1095 5093 1146
rect 5042 985 5093 1036
rect 5042 875 5093 926
rect 446 429 492 475
rect 446 318 492 364
rect 891 324 942 440
rect 889 73 940 189
rect 3128 655 3179 706
rect 5042 765 5093 816
rect 3128 545 3179 596
rect 6956 1315 7007 1366
rect 6956 1205 7007 1256
rect 6956 1095 7007 1146
rect 6956 985 7007 1036
rect 6956 875 7007 926
rect 5042 655 5093 706
rect 6956 765 7007 816
rect 3128 435 3179 486
rect 3128 325 3179 376
rect 3128 215 3179 266
rect 446 7 492 53
rect 446 -104 492 -58
rect 446 -215 492 -169
rect 890 -167 941 -51
rect 446 -326 492 -280
rect 446 -437 492 -391
rect 5042 545 5093 596
rect 6956 655 7007 706
rect 5042 435 5093 486
rect 3128 105 3179 156
rect 3128 -5 3179 46
rect 3128 -115 3179 -64
rect 5042 325 5093 376
rect 5042 215 5093 266
rect 3128 -225 3179 -174
rect 6956 545 7007 596
rect 6956 435 7007 486
rect 5042 105 5093 156
rect 5042 -5 5093 46
rect 5042 -115 5093 -64
rect 3128 -335 3179 -284
rect 6956 325 7007 376
rect 6956 215 7007 266
rect 5042 -225 5093 -174
rect 6956 105 7007 156
rect 6956 -5 7007 46
rect 6956 -115 7007 -64
rect 5042 -335 5093 -284
rect 3128 -445 3179 -394
rect 6956 -225 7007 -174
rect 6956 -335 7007 -284
rect 5042 -445 5093 -394
rect 6956 -445 7007 -394
<< polysilicon >>
rect 1047 1615 1120 1628
rect 1047 1569 1061 1615
rect 1107 1569 1120 1615
rect -205 1425 -133 1433
rect 314 1442 386 1455
rect 314 1425 327 1442
rect -205 1420 -89 1425
rect -205 1374 -192 1420
rect -146 1374 -89 1420
rect -205 1369 -89 1374
rect -39 1369 5 1425
rect 128 1369 201 1425
rect 251 1396 327 1425
rect 373 1396 386 1442
rect 251 1369 386 1396
rect -205 1361 -133 1369
rect 128 1257 167 1369
rect -133 1201 -89 1257
rect -39 1201 201 1257
rect 251 1201 295 1257
rect 1047 1556 1120 1569
rect 1056 1419 1112 1556
rect 1056 1363 1144 1419
rect 1194 1363 1274 1419
rect 1324 1363 1407 1419
rect 1457 1363 1537 1419
rect 1587 1363 1839 1419
rect 1889 1363 1933 1419
rect 2972 1429 3044 1442
rect 2972 1383 2985 1429
rect 3031 1383 3044 1429
rect 1631 1273 1703 1286
rect 1631 1251 1644 1273
rect 1100 1195 1144 1251
rect 1194 1195 1274 1251
rect 1324 1195 1407 1251
rect 1457 1195 1537 1251
rect 1587 1227 1644 1251
rect 1690 1251 1703 1273
rect 1690 1227 1839 1251
rect 1587 1195 1839 1227
rect 1889 1195 1933 1251
rect 1632 977 1704 990
rect 1021 949 1094 957
rect 1632 949 1645 977
rect 1021 944 1144 949
rect 1021 898 1035 944
rect 1081 898 1144 944
rect 1021 893 1144 898
rect 1194 893 1238 949
rect 1363 893 1407 949
rect 1457 893 1537 949
rect 1587 931 1645 949
rect 1691 949 1704 977
rect 1691 931 1839 949
rect 1587 893 1839 931
rect 1889 893 1933 949
rect 1021 885 1094 893
rect -209 669 -137 677
rect 310 686 382 699
rect 310 669 323 686
rect -209 664 -93 669
rect -209 618 -196 664
rect -150 618 -93 664
rect -209 613 -93 618
rect -43 613 1 669
rect 124 613 197 669
rect 247 640 323 669
rect 369 640 382 686
rect 247 613 382 640
rect 2972 1370 3044 1383
rect 3263 1429 3335 1442
rect 3263 1383 3276 1429
rect 3322 1383 3335 1429
rect 2704 1277 2776 1290
rect 2704 1232 2717 1277
rect 2458 1176 2502 1232
rect 2552 1231 2717 1232
rect 2763 1232 2776 1277
rect 2763 1231 2834 1232
rect 2552 1176 2834 1231
rect 2884 1176 2928 1232
rect 2593 1064 2629 1176
rect 2458 1008 2502 1064
rect 2552 1008 2629 1064
rect 2753 1064 2790 1176
rect 2753 1008 2834 1064
rect 2884 1008 2928 1064
rect 2593 896 2629 1008
rect 2980 896 3036 1370
rect 2458 840 2502 896
rect 2552 840 2629 896
rect 2754 840 2834 896
rect 2884 840 3036 896
rect 3263 1370 3335 1383
rect 4886 1429 4958 1442
rect 4886 1383 4899 1429
rect 4945 1383 4958 1429
rect -209 605 -137 613
rect 124 501 163 613
rect 2754 728 2790 840
rect 3271 896 3327 1370
rect 4886 1370 4958 1383
rect 5177 1429 5249 1442
rect 5177 1383 5190 1429
rect 5236 1383 5249 1429
rect 3531 1277 3603 1290
rect 3531 1232 3544 1277
rect 3379 1176 3423 1232
rect 3473 1231 3544 1232
rect 3590 1232 3603 1277
rect 3590 1231 3755 1232
rect 3473 1176 3755 1231
rect 3805 1176 3849 1232
rect 4618 1277 4690 1290
rect 4618 1232 4631 1277
rect 3517 1064 3554 1176
rect 3379 1008 3423 1064
rect 3473 1008 3554 1064
rect 3678 1064 3714 1176
rect 4372 1176 4416 1232
rect 4466 1231 4631 1232
rect 4677 1232 4690 1277
rect 4677 1231 4748 1232
rect 4466 1176 4748 1231
rect 4798 1176 4842 1232
rect 3678 1008 3755 1064
rect 3805 1008 3849 1064
rect 4507 1064 4543 1176
rect 3678 896 3714 1008
rect 4372 1008 4416 1064
rect 4466 1008 4543 1064
rect 4667 1064 4704 1176
rect 4667 1008 4748 1064
rect 4798 1008 4842 1064
rect 3271 840 3423 896
rect 3473 840 3553 896
rect 3678 840 3755 896
rect 3805 840 3849 896
rect 4507 896 4543 1008
rect 4894 896 4950 1370
rect 2458 672 2502 728
rect 2552 672 2834 728
rect 2884 672 2928 728
rect 3517 728 3553 840
rect 4372 840 4416 896
rect 4466 840 4543 896
rect 4668 840 4748 896
rect 4798 840 4950 896
rect 5177 1370 5249 1383
rect 6800 1429 6872 1442
rect 6800 1383 6813 1429
rect 6859 1383 6872 1429
rect -137 445 -93 501
rect -43 445 197 501
rect 247 445 291 501
rect 1456 520 1538 536
rect 1020 505 1095 519
rect 1020 459 1035 505
rect 1081 459 1095 505
rect 1020 445 1095 459
rect 1456 472 1475 520
rect 1524 486 1538 520
rect 1524 472 1585 486
rect 1456 456 1585 472
rect 1035 158 1081 445
rect 1471 430 1585 456
rect 1635 430 1679 486
rect 1471 318 1527 430
rect 2583 560 2619 672
rect 3379 672 3423 728
rect 3473 672 3755 728
rect 3805 672 3849 728
rect 4668 728 4704 840
rect 5185 896 5241 1370
rect 6800 1370 6872 1383
rect 5445 1277 5517 1290
rect 5445 1232 5458 1277
rect 5293 1176 5337 1232
rect 5387 1231 5458 1232
rect 5504 1232 5517 1277
rect 5504 1231 5669 1232
rect 5387 1176 5669 1231
rect 5719 1176 5763 1232
rect 6532 1277 6604 1290
rect 6532 1232 6545 1277
rect 5431 1064 5468 1176
rect 5293 1008 5337 1064
rect 5387 1008 5468 1064
rect 5592 1064 5628 1176
rect 6286 1176 6330 1232
rect 6380 1231 6545 1232
rect 6591 1232 6604 1277
rect 6591 1231 6662 1232
rect 6380 1176 6662 1231
rect 6712 1176 6756 1232
rect 5592 1008 5669 1064
rect 5719 1008 5763 1064
rect 6421 1064 6457 1176
rect 5592 896 5628 1008
rect 6286 1008 6330 1064
rect 6380 1008 6457 1064
rect 6581 1064 6618 1176
rect 6581 1008 6662 1064
rect 6712 1008 6756 1064
rect 5185 840 5337 896
rect 5387 840 5467 896
rect 5592 840 5669 896
rect 5719 840 5763 896
rect 6421 896 6457 1008
rect 6808 896 6864 1370
rect 2942 560 3014 568
rect 2458 504 2502 560
rect 2552 504 2619 560
rect 2790 504 2834 560
rect 2884 555 3014 560
rect 2884 509 2955 555
rect 3001 509 3014 555
rect 2884 504 3014 509
rect 2583 392 2619 504
rect 2942 496 3014 504
rect 3293 560 3365 568
rect 3688 560 3724 672
rect 4372 672 4416 728
rect 4466 672 4748 728
rect 4798 672 4842 728
rect 5431 728 5467 840
rect 6286 840 6330 896
rect 6380 840 6457 896
rect 6582 840 6662 896
rect 6712 840 6864 896
rect 3293 555 3423 560
rect 3293 509 3306 555
rect 3352 509 3423 555
rect 3293 504 3423 509
rect 3473 504 3517 560
rect 3688 504 3755 560
rect 3805 504 3849 560
rect 4497 560 4533 672
rect 5293 672 5337 728
rect 5387 672 5669 728
rect 5719 672 5763 728
rect 6582 728 6618 840
rect 4856 560 4928 568
rect 3293 496 3365 504
rect 2458 336 2502 392
rect 2552 336 2619 392
rect 2790 336 2834 392
rect 2884 336 2964 392
rect 1131 262 1175 318
rect 1275 262 1585 318
rect 1635 262 1679 318
rect 1035 102 1175 158
rect 1275 150 1319 158
rect 2294 227 2366 240
rect 2294 181 2307 227
rect 2353 224 2366 227
rect 2928 224 2964 336
rect 2353 181 2502 224
rect 2294 168 2502 181
rect 2552 168 2834 224
rect 2884 168 2964 224
rect 3688 392 3724 504
rect 4372 504 4416 560
rect 4466 504 4533 560
rect 4704 504 4748 560
rect 4798 555 4928 560
rect 4798 509 4869 555
rect 4915 509 4928 555
rect 4798 504 4928 509
rect 1275 102 1585 150
rect -209 -86 -137 -78
rect 310 -69 382 -56
rect 310 -86 323 -69
rect -209 -91 -93 -86
rect -209 -137 -196 -91
rect -150 -137 -93 -91
rect -209 -142 -93 -137
rect -43 -142 1 -86
rect 124 -142 197 -86
rect 247 -115 323 -86
rect 369 -115 382 -69
rect 247 -142 382 -115
rect 1481 94 1585 102
rect 1635 94 1679 150
rect 1337 15 1415 35
rect 1337 8 1355 15
rect 1327 -2 1355 8
rect -209 -150 -137 -142
rect 124 -254 163 -142
rect 1131 -58 1175 -2
rect 1275 -31 1355 -2
rect 1401 -31 1415 15
rect 1275 -42 1415 -31
rect 1481 -18 1529 94
rect 1275 -58 1408 -42
rect -137 -310 -93 -254
rect -43 -310 197 -254
rect 247 -310 291 -254
rect 1319 -383 1375 -58
rect 1481 -74 1585 -18
rect 1635 -74 1679 -18
rect 2432 56 2468 168
rect 3343 336 3423 392
rect 3473 336 3517 392
rect 3688 336 3755 392
rect 3805 336 3849 392
rect 4497 392 4533 504
rect 4856 496 4928 504
rect 5207 560 5279 568
rect 5602 560 5638 672
rect 6286 672 6330 728
rect 6380 672 6662 728
rect 6712 672 6756 728
rect 5207 555 5337 560
rect 5207 509 5220 555
rect 5266 509 5337 555
rect 5207 504 5337 509
rect 5387 504 5431 560
rect 5602 504 5669 560
rect 5719 504 5763 560
rect 6411 560 6447 672
rect 6770 560 6842 568
rect 5207 496 5279 504
rect 3343 224 3379 336
rect 4372 336 4416 392
rect 4466 336 4533 392
rect 4704 336 4748 392
rect 4798 336 4878 392
rect 3941 227 4013 240
rect 3941 224 3954 227
rect 3343 168 3423 224
rect 3473 168 3755 224
rect 3805 181 3954 224
rect 4000 181 4013 227
rect 3805 168 4013 181
rect 2942 56 3014 64
rect 2432 0 2502 56
rect 2552 0 2596 56
rect 2790 0 2834 56
rect 2884 51 3014 56
rect 2884 5 2955 51
rect 3001 5 3014 51
rect 2884 0 3014 5
rect 2432 -112 2468 0
rect 2942 -8 3014 0
rect 2688 -72 2760 -59
rect 2432 -168 2502 -112
rect 2552 -168 2596 -112
rect 2688 -118 2701 -72
rect 2747 -112 2760 -72
rect 3293 56 3365 64
rect 3839 56 3875 168
rect 3293 51 3423 56
rect 3293 5 3306 51
rect 3352 5 3423 51
rect 3293 0 3423 5
rect 3473 0 3517 56
rect 3711 0 3755 56
rect 3805 0 3875 56
rect 3293 -8 3365 0
rect 2747 -118 2834 -112
rect 2688 -168 2834 -118
rect 2884 -168 2928 -112
rect 3547 -72 3619 -59
rect 3547 -112 3560 -72
rect 2754 -280 2790 -168
rect 3379 -168 3423 -112
rect 3473 -118 3560 -112
rect 3606 -118 3619 -72
rect 3839 -112 3875 0
rect 3473 -168 3619 -118
rect 3711 -168 3755 -112
rect 3805 -168 3875 -112
rect 4208 227 4280 240
rect 4208 181 4221 227
rect 4267 224 4280 227
rect 4842 224 4878 336
rect 4267 181 4416 224
rect 4208 168 4416 181
rect 4466 168 4748 224
rect 4798 168 4878 224
rect 5602 392 5638 504
rect 6286 504 6330 560
rect 6380 504 6447 560
rect 6618 504 6662 560
rect 6712 555 6842 560
rect 6712 509 6783 555
rect 6829 509 6842 555
rect 6712 504 6842 509
rect 2458 -336 2502 -280
rect 2552 -336 2834 -280
rect 2884 -336 2928 -280
rect 3517 -280 3553 -168
rect 4346 56 4382 168
rect 5257 336 5337 392
rect 5387 336 5431 392
rect 5602 336 5669 392
rect 5719 336 5763 392
rect 6411 392 6447 504
rect 6770 496 6842 504
rect 5257 224 5293 336
rect 6286 336 6330 392
rect 6380 336 6447 392
rect 6618 336 6662 392
rect 6712 336 6792 392
rect 5855 227 5927 240
rect 5855 224 5868 227
rect 5257 168 5337 224
rect 5387 168 5669 224
rect 5719 181 5868 224
rect 5914 181 5927 227
rect 5719 168 5927 181
rect 4856 56 4928 64
rect 4346 0 4416 56
rect 4466 0 4510 56
rect 4704 0 4748 56
rect 4798 51 4928 56
rect 4798 5 4869 51
rect 4915 5 4928 51
rect 4798 0 4928 5
rect 4346 -112 4382 0
rect 4856 -8 4928 0
rect 4602 -72 4674 -59
rect 4346 -168 4416 -112
rect 4466 -168 4510 -112
rect 4602 -118 4615 -72
rect 4661 -112 4674 -72
rect 5207 56 5279 64
rect 5753 56 5789 168
rect 5207 51 5337 56
rect 5207 5 5220 51
rect 5266 5 5337 51
rect 5207 0 5337 5
rect 5387 0 5431 56
rect 5625 0 5669 56
rect 5719 0 5789 56
rect 5207 -8 5279 0
rect 4661 -118 4748 -112
rect 4602 -168 4748 -118
rect 4798 -168 4842 -112
rect 5461 -72 5533 -59
rect 5461 -112 5474 -72
rect 1319 -439 1585 -383
rect 1635 -439 1679 -383
rect 3379 -336 3423 -280
rect 3473 -336 3755 -280
rect 3805 -336 3849 -280
rect 4668 -280 4704 -168
rect 5293 -168 5337 -112
rect 5387 -118 5474 -112
rect 5520 -118 5533 -72
rect 5753 -112 5789 0
rect 5387 -168 5533 -118
rect 5625 -168 5669 -112
rect 5719 -168 5789 -112
rect 6122 227 6194 240
rect 6122 181 6135 227
rect 6181 224 6194 227
rect 6756 224 6792 336
rect 6181 181 6330 224
rect 6122 168 6330 181
rect 6380 168 6662 224
rect 6712 168 6792 224
rect 4372 -336 4416 -280
rect 4466 -336 4748 -280
rect 4798 -336 4842 -280
rect 5431 -280 5467 -168
rect 6260 56 6296 168
rect 6770 56 6842 64
rect 6260 0 6330 56
rect 6380 0 6424 56
rect 6618 0 6662 56
rect 6712 51 6842 56
rect 6712 5 6783 51
rect 6829 5 6842 51
rect 6712 0 6842 5
rect 6260 -112 6296 0
rect 6770 -8 6842 0
rect 6516 -72 6588 -59
rect 6260 -168 6330 -112
rect 6380 -168 6424 -112
rect 6516 -118 6529 -72
rect 6575 -112 6588 -72
rect 6575 -118 6662 -112
rect 6516 -168 6662 -118
rect 6712 -168 6756 -112
rect 5293 -336 5337 -280
rect 5387 -336 5669 -280
rect 5719 -336 5763 -280
rect 6582 -280 6618 -168
rect 6286 -336 6330 -280
rect 6380 -336 6662 -280
rect 6712 -336 6756 -280
<< polycontact >>
rect 1061 1569 1107 1615
rect -192 1374 -146 1420
rect 327 1396 373 1442
rect 2985 1383 3031 1429
rect 1644 1227 1690 1273
rect 1035 898 1081 944
rect 1645 931 1691 977
rect -196 618 -150 664
rect 323 640 369 686
rect 3276 1383 3322 1429
rect 2717 1231 2763 1277
rect 4899 1383 4945 1429
rect 5190 1383 5236 1429
rect 3544 1231 3590 1277
rect 4631 1231 4677 1277
rect 6813 1383 6859 1429
rect 1035 459 1081 505
rect 1475 472 1524 520
rect 5458 1231 5504 1277
rect 6545 1231 6591 1277
rect 2955 509 3001 555
rect 3306 509 3352 555
rect 2307 181 2353 227
rect 4869 509 4915 555
rect -196 -137 -150 -91
rect 323 -115 369 -69
rect 1355 -31 1401 15
rect 5220 509 5266 555
rect 3954 181 4000 227
rect 2955 5 3001 51
rect 2701 -118 2747 -72
rect 3306 5 3352 51
rect 3560 -118 3606 -72
rect 4221 181 4267 227
rect 6783 509 6829 555
rect 5868 181 5914 227
rect 4869 5 4915 51
rect 4615 -118 4661 -72
rect 5220 5 5266 51
rect 5474 -118 5520 -72
rect 6135 181 6181 227
rect 6783 5 6829 51
rect 6529 -118 6575 -72
<< metal1 >>
rect -607 2398 -529 2410
rect -607 2344 -595 2398
rect -541 2344 -529 2398
rect -607 2332 -529 2344
rect 2304 2398 2382 2410
rect 2304 2344 2316 2398
rect 2370 2344 2382 2398
rect 2304 2332 2382 2344
rect 4218 2398 4296 2410
rect 4218 2344 4230 2398
rect 4284 2344 4296 2398
rect 4218 2332 4296 2344
rect 6130 2398 6208 2410
rect 6130 2344 6142 2398
rect 6196 2344 6208 2398
rect 6130 2332 6208 2344
rect -607 -533 -560 2332
rect 669 2271 747 2283
rect 669 2217 681 2271
rect 735 2217 747 2271
rect 669 2205 747 2217
rect 1628 2271 1706 2283
rect 1628 2217 1640 2271
rect 1694 2217 1706 2271
rect 1628 2205 1706 2217
rect -511 2143 -433 2155
rect -511 2089 -499 2143
rect -445 2089 -433 2143
rect -511 2077 -433 2089
rect -511 216 -464 2077
rect 544 2006 622 2018
rect 544 1952 556 2006
rect 610 1952 622 2006
rect 544 1940 622 1952
rect -417 1880 -339 1892
rect -417 1826 -405 1880
rect -351 1826 -339 1880
rect -417 1814 -339 1826
rect -417 973 -370 1814
rect 312 1755 390 1767
rect 312 1701 324 1755
rect 378 1701 390 1755
rect 312 1689 390 1701
rect -322 1564 -242 1587
rect -322 1518 -305 1564
rect -259 1518 -242 1564
rect -322 1453 -242 1518
rect -87 1504 -41 1515
rect 203 1504 249 1515
rect -322 1407 -305 1453
rect -259 1420 -242 1453
rect -189 1458 -87 1504
rect -189 1433 -133 1458
rect -87 1447 -41 1458
rect 109 1458 203 1504
rect -196 1420 -133 1433
rect -259 1407 -192 1420
rect -322 1374 -192 1407
rect -146 1374 -133 1420
rect -322 1342 -242 1374
rect -196 1361 -133 1374
rect -322 1296 -305 1342
rect -259 1296 -242 1342
rect -322 1231 -242 1296
rect -189 1336 -133 1361
rect -87 1336 -41 1347
rect -189 1290 -87 1336
rect -87 1279 -41 1290
rect -322 1185 -305 1231
rect -259 1185 -242 1231
rect -322 1120 -242 1185
rect -322 1074 -305 1120
rect -259 1074 -242 1120
rect -87 1168 -41 1179
rect 109 1168 155 1458
rect 203 1447 249 1458
rect 327 1455 373 1689
rect 433 1564 513 1587
rect 433 1518 450 1564
rect 496 1518 513 1564
rect 314 1442 386 1455
rect 314 1396 327 1442
rect 373 1396 386 1442
rect 314 1383 386 1396
rect 433 1453 513 1518
rect 433 1407 450 1453
rect 496 1407 513 1453
rect 203 1336 249 1347
rect 433 1342 513 1407
rect 433 1336 450 1342
rect 249 1296 450 1336
rect 496 1296 513 1342
rect 249 1290 513 1296
rect 203 1279 249 1290
rect 433 1231 513 1290
rect 433 1185 450 1231
rect 496 1185 513 1231
rect 203 1168 249 1179
rect -41 1122 203 1168
rect -87 1111 -41 1122
rect -322 1039 -242 1074
rect -417 961 -339 973
rect -417 907 -405 961
rect -351 907 -339 961
rect -417 895 -339 907
rect -293 831 -246 1039
rect 58 973 104 1122
rect 203 1111 249 1122
rect 433 1120 513 1185
rect 433 1074 450 1120
rect 496 1074 513 1120
rect 433 1039 513 1074
rect 42 961 120 973
rect 42 907 54 961
rect 108 907 120 961
rect 42 895 120 907
rect -326 808 -246 831
rect 303 885 381 897
rect 303 831 315 885
rect 369 831 381 885
rect 441 831 489 1039
rect 559 941 606 1940
rect 545 929 623 941
rect 545 875 557 929
rect 611 875 623 929
rect 545 863 623 875
rect 303 819 381 831
rect -326 762 -309 808
rect -263 762 -246 808
rect -326 697 -246 762
rect -91 748 -45 759
rect 199 748 245 759
rect -326 651 -309 697
rect -263 664 -246 697
rect -193 702 -91 748
rect -193 677 -137 702
rect -91 691 -45 702
rect 105 702 199 748
rect -200 664 -137 677
rect -263 651 -196 664
rect -326 618 -196 651
rect -150 618 -137 664
rect -326 586 -246 618
rect -200 605 -137 618
rect -326 540 -309 586
rect -263 540 -246 586
rect -326 475 -246 540
rect -193 580 -137 605
rect -91 580 -45 591
rect -193 534 -91 580
rect -91 523 -45 534
rect -326 429 -309 475
rect -263 429 -246 475
rect -326 364 -246 429
rect -326 318 -309 364
rect -263 318 -246 364
rect -91 412 -45 423
rect 105 412 151 702
rect 199 691 245 702
rect 323 699 369 819
rect 429 808 509 831
rect 429 762 446 808
rect 492 762 509 808
rect 310 686 382 699
rect 310 640 323 686
rect 369 640 382 686
rect 310 627 382 640
rect 429 697 509 762
rect 429 651 446 697
rect 492 651 509 697
rect 199 580 245 591
rect 429 586 509 651
rect 429 580 446 586
rect 245 540 446 580
rect 492 540 509 586
rect 245 534 509 540
rect 199 523 245 534
rect 429 475 509 534
rect 429 429 446 475
rect 492 429 509 475
rect 199 412 245 423
rect -45 366 199 412
rect -91 355 -45 366
rect -326 283 -246 318
rect -511 204 -433 216
rect -511 150 -499 204
rect -445 150 -433 204
rect -511 138 -433 150
rect -295 76 -247 283
rect 54 216 100 366
rect 199 355 245 366
rect 429 364 509 429
rect 429 318 446 364
rect 492 318 509 364
rect 429 283 509 318
rect 38 204 116 216
rect 38 150 50 204
rect 104 150 116 204
rect 38 138 116 150
rect 310 155 375 167
rect 310 101 319 155
rect 373 101 375 155
rect 310 89 375 101
rect -326 53 -246 76
rect -326 7 -309 53
rect -263 7 -246 53
rect -326 -58 -246 7
rect -91 -7 -45 4
rect 199 -7 245 4
rect -326 -104 -309 -58
rect -263 -91 -246 -58
rect -193 -53 -91 -7
rect -193 -78 -137 -53
rect -91 -64 -45 -53
rect 105 -53 199 -7
rect -200 -91 -137 -78
rect -263 -104 -196 -91
rect -326 -137 -196 -104
rect -150 -137 -137 -91
rect -326 -169 -246 -137
rect -200 -150 -137 -137
rect -326 -215 -309 -169
rect -263 -215 -246 -169
rect -326 -280 -246 -215
rect -193 -175 -137 -150
rect -91 -175 -45 -164
rect -193 -221 -91 -175
rect -91 -232 -45 -221
rect -326 -326 -309 -280
rect -263 -326 -246 -280
rect -326 -391 -246 -326
rect -326 -437 -309 -391
rect -263 -437 -246 -391
rect -91 -343 -45 -332
rect 105 -343 151 -53
rect 199 -64 245 -53
rect 323 -56 369 89
rect 446 76 494 283
rect 669 166 716 2205
rect 1045 2017 1123 2029
rect 1045 1963 1057 2017
rect 1111 1963 1123 2017
rect 1045 1951 1123 1963
rect 762 1755 840 1767
rect 762 1701 774 1755
rect 828 1701 840 1755
rect 762 1689 840 1701
rect 762 643 809 1689
rect 1061 1628 1107 1951
rect 1047 1615 1120 1628
rect 860 1553 974 1583
rect 1047 1569 1061 1615
rect 1107 1569 1120 1615
rect 1047 1556 1120 1569
rect 860 1498 889 1553
rect 944 1498 974 1553
rect 1146 1498 1192 1509
rect 1276 1498 1322 1509
rect 1409 1498 1455 1509
rect 1539 1498 1585 1509
rect 860 1452 1146 1498
rect 1192 1452 1276 1498
rect 1322 1452 1409 1498
rect 1455 1452 1539 1498
rect 860 1430 974 1452
rect 1146 1441 1192 1452
rect 1276 1441 1322 1452
rect 1409 1441 1455 1452
rect 1539 1441 1585 1452
rect 860 1375 889 1430
rect 944 1375 974 1430
rect 860 1307 974 1375
rect 860 1252 889 1307
rect 944 1252 974 1307
rect 1146 1330 1192 1341
rect 1276 1330 1322 1341
rect 1409 1330 1455 1341
rect 1539 1330 1585 1341
rect 1192 1284 1276 1330
rect 1322 1284 1409 1330
rect 1455 1284 1539 1330
rect 1644 1286 1690 2205
rect 1984 1553 2098 1583
rect 1841 1498 1887 1509
rect 1749 1452 1841 1498
rect 1146 1273 1192 1284
rect 1276 1273 1322 1284
rect 1409 1273 1455 1284
rect 1539 1273 1585 1284
rect 1631 1273 1703 1286
rect 860 1184 974 1252
rect 1631 1227 1644 1273
rect 1690 1227 1703 1273
rect 1631 1214 1703 1227
rect 860 1129 889 1184
rect 944 1129 974 1184
rect 860 1061 974 1129
rect 1146 1162 1192 1173
rect 1276 1162 1322 1173
rect 1409 1162 1455 1173
rect 1539 1162 1585 1173
rect 1749 1162 1795 1452
rect 1841 1441 1887 1452
rect 1984 1498 2013 1553
rect 2068 1498 2098 1553
rect 1984 1430 2098 1498
rect 1984 1375 2013 1430
rect 2068 1375 2098 1430
rect 1841 1330 1887 1341
rect 1984 1330 2098 1375
rect 1887 1307 2098 1330
rect 1887 1284 2013 1307
rect 1841 1273 1887 1284
rect 1984 1252 2013 1284
rect 2068 1252 2098 1307
rect 1984 1184 2098 1252
rect 1841 1162 1887 1173
rect 1192 1116 1276 1162
rect 1322 1116 1409 1162
rect 1455 1116 1539 1162
rect 1585 1116 1841 1162
rect 1146 1105 1192 1116
rect 1276 1105 1322 1116
rect 1409 1105 1455 1116
rect 1539 1105 1585 1116
rect 860 1006 889 1061
rect 944 1006 974 1061
rect 1146 1028 1192 1039
rect 1409 1028 1455 1039
rect 1539 1028 1585 1039
rect 860 944 974 1006
rect 1035 982 1146 1028
rect 1192 982 1409 1028
rect 1455 982 1539 1028
rect 1645 990 1691 1116
rect 1841 1105 1887 1116
rect 1984 1129 2013 1184
rect 2068 1129 2098 1184
rect 1984 1061 2098 1129
rect 1841 1028 1887 1039
rect 1984 1028 2013 1061
rect 1035 957 1094 982
rect 1146 971 1192 982
rect 1409 971 1455 982
rect 1539 971 1585 982
rect 1632 977 1704 990
rect 1021 944 1094 957
rect 860 938 1035 944
rect 860 883 889 938
rect 944 898 1035 938
rect 1081 898 1094 944
rect 1632 931 1645 977
rect 1691 931 1704 977
rect 1887 1006 2013 1028
rect 2068 1006 2098 1061
rect 1887 982 2098 1006
rect 1841 971 1887 982
rect 1632 918 1704 931
rect 1984 938 2098 982
rect 944 883 974 898
rect 1021 885 1094 898
rect 860 815 974 883
rect 860 760 889 815
rect 944 760 974 815
rect 1035 860 1094 885
rect 1984 883 2013 938
rect 2068 883 2098 938
rect 1146 860 1192 871
rect 1409 860 1455 871
rect 1539 860 1585 871
rect 1841 860 1887 871
rect 1035 814 1146 860
rect 1146 803 1192 814
rect 1298 814 1409 860
rect 1455 814 1539 860
rect 1585 814 1841 860
rect 860 729 974 760
rect 762 631 840 643
rect 762 577 774 631
rect 828 577 840 631
rect 762 565 840 577
rect 891 492 939 729
rect 1298 652 1344 814
rect 1409 803 1455 814
rect 1539 803 1585 814
rect 1841 803 1887 814
rect 1984 815 2098 883
rect 1984 760 2013 815
rect 2068 760 2098 815
rect 1984 729 2098 760
rect 2146 1366 2248 1393
rect 2146 1314 2173 1366
rect 2220 1314 2248 1366
rect 2146 1256 2248 1314
rect 2146 1204 2173 1256
rect 2220 1204 2248 1256
rect 2146 1146 2248 1204
rect 2146 1094 2173 1146
rect 2220 1094 2248 1146
rect 2146 1036 2248 1094
rect 2146 984 2173 1036
rect 2220 984 2248 1036
rect 2146 926 2248 984
rect 2146 874 2173 926
rect 2220 874 2248 926
rect 2146 816 2248 874
rect 2146 764 2173 816
rect 2220 764 2248 816
rect 1017 631 1095 643
rect 1017 577 1029 631
rect 1083 577 1095 631
rect 1298 606 1523 652
rect 1017 565 1095 577
rect 1033 519 1079 565
rect 1476 536 1523 606
rect 1587 565 1633 576
rect 1456 520 1538 536
rect 1020 505 1095 519
rect 610 154 716 166
rect 610 100 622 154
rect 676 100 716 154
rect 610 88 716 100
rect 846 440 969 492
rect 1020 459 1035 505
rect 1081 459 1095 505
rect 1020 445 1095 459
rect 1456 472 1475 520
rect 1524 472 1538 520
rect 1633 519 1729 565
rect 1587 508 1633 519
rect 1456 456 1538 472
rect 846 324 891 440
rect 942 393 969 440
rect 1587 397 1633 408
rect 942 347 1188 393
rect 1262 347 1273 393
rect 1356 351 1587 397
rect 942 324 969 347
rect 846 189 969 324
rect 1356 233 1402 351
rect 1587 340 1633 351
rect 429 53 509 76
rect 429 7 446 53
rect 492 7 509 53
rect 310 -69 382 -56
rect 310 -115 323 -69
rect 369 -115 382 -69
rect 310 -128 382 -115
rect 429 -58 509 7
rect 429 -104 446 -58
rect 492 -104 509 -58
rect 429 -107 509 -104
rect 846 73 889 189
rect 940 73 969 189
rect 1177 187 1188 233
rect 1262 187 1402 233
rect 1585 229 1633 240
rect 1683 229 1729 519
rect 846 27 1188 73
rect 1262 27 1273 73
rect 1356 35 1402 187
rect 1492 183 1587 229
rect 1633 183 1729 229
rect 1779 551 1893 603
rect 1779 422 1805 551
rect 1864 538 1893 551
rect 2014 538 2062 729
rect 2146 706 2248 764
rect 2146 654 2173 706
rect 2220 654 2248 706
rect 2146 596 2248 654
rect 2146 544 2173 596
rect 2220 544 2248 596
rect 2146 538 2248 544
rect 1864 490 2248 538
rect 1864 422 1893 490
rect 1779 306 1893 422
rect 846 -51 969 27
rect 1337 15 1415 35
rect 1337 -31 1355 15
rect 1401 -31 1415 15
rect 1337 -42 1415 -31
rect 846 -107 890 -51
rect 199 -175 245 -164
rect 429 -167 890 -107
rect 941 -167 969 -51
rect 1177 -133 1188 -87
rect 1262 -133 1319 -87
rect 429 -169 969 -167
rect 429 -175 446 -169
rect 245 -215 446 -175
rect 492 -178 969 -169
rect 492 -215 509 -178
rect 245 -221 509 -215
rect 199 -232 245 -221
rect 429 -280 509 -221
rect 846 -232 969 -178
rect 429 -326 446 -280
rect 492 -326 509 -280
rect 199 -343 245 -332
rect -45 -389 199 -343
rect -91 -400 -45 -389
rect -326 -472 -246 -437
rect -607 -545 -529 -533
rect -607 -599 -595 -545
rect -541 -599 -529 -545
rect -607 -611 -529 -599
rect -309 -687 -263 -472
rect 54 -534 100 -389
rect 199 -400 245 -389
rect 429 -391 509 -326
rect 429 -437 446 -391
rect 492 -437 509 -391
rect 429 -472 509 -437
rect 1272 -471 1319 -133
rect 1492 -107 1538 183
rect 1585 172 1633 183
rect 1779 177 1799 306
rect 1858 177 1893 306
rect 1779 74 1893 177
rect 1587 61 1633 72
rect 1779 61 1802 74
rect 1633 15 1802 61
rect 1587 4 1633 15
rect 1779 -55 1802 15
rect 1861 -55 1893 74
rect 1585 -107 1633 -96
rect 1492 -153 1587 -107
rect 1585 -164 1633 -153
rect 1779 -173 1893 -55
rect 1587 -304 1633 -293
rect 1779 -302 1803 -173
rect 1862 -302 1893 -173
rect 1779 -304 1893 -302
rect 1633 -350 1893 -304
rect 1587 -361 1633 -350
rect 1779 -397 1893 -350
rect 1587 -471 1633 -461
rect 1272 -472 1633 -471
rect 38 -546 116 -534
rect 38 -600 50 -546
rect 104 -600 116 -546
rect 38 -612 116 -600
rect -325 -699 -247 -687
rect -325 -753 -313 -699
rect -259 -753 -247 -699
rect -325 -765 -247 -753
rect 451 -827 497 -472
rect 1272 -518 1587 -472
rect 435 -839 513 -827
rect 435 -893 447 -839
rect 501 -893 513 -839
rect 435 -905 513 -893
rect 1272 -950 1319 -518
rect 1587 -529 1633 -518
rect 1779 -526 1803 -397
rect 1862 -526 1893 -397
rect 2146 486 2248 490
rect 2146 434 2173 486
rect 2220 434 2248 486
rect 2146 376 2248 434
rect 2146 324 2173 376
rect 2220 324 2248 376
rect 2146 266 2248 324
rect 2146 214 2173 266
rect 2220 214 2248 266
rect 2320 240 2366 2332
rect 3925 2271 4003 2283
rect 3925 2217 3937 2271
rect 3991 2217 4003 2271
rect 3925 2205 4003 2217
rect 2969 2144 3047 2156
rect 2969 2090 2981 2144
rect 3035 2090 3047 2144
rect 2969 2078 3047 2090
rect 2701 1755 2779 1767
rect 2701 1701 2713 1755
rect 2767 1701 2779 1755
rect 2701 1689 2779 1701
rect 2504 1311 2550 1322
rect 2550 1265 2642 1311
rect 2717 1290 2763 1689
rect 2985 1442 3031 2078
rect 3260 2017 3338 2029
rect 3260 1963 3272 2017
rect 3326 1963 3338 2017
rect 3260 1951 3338 1963
rect 3276 1442 3322 1951
rect 3528 1880 3606 1892
rect 3528 1826 3540 1880
rect 3594 1826 3606 1880
rect 3528 1814 3606 1826
rect 2972 1429 3044 1442
rect 2972 1383 2985 1429
rect 3031 1383 3044 1429
rect 3263 1429 3335 1442
rect 2972 1370 3044 1383
rect 3102 1366 3205 1392
rect 3263 1383 3276 1429
rect 3322 1383 3335 1429
rect 3263 1370 3335 1383
rect 2836 1311 2882 1322
rect 3102 1315 3128 1366
rect 3179 1315 3205 1366
rect 3102 1311 3205 1315
rect 3425 1311 3471 1322
rect 2504 1254 2550 1265
rect 2504 1143 2550 1154
rect 2412 1097 2504 1143
rect 2412 807 2458 1097
rect 2504 1086 2550 1097
rect 2596 1015 2642 1265
rect 2704 1277 2776 1290
rect 2704 1231 2717 1277
rect 2763 1231 2776 1277
rect 2882 1265 3425 1311
rect 3544 1290 3590 1814
rect 3757 1311 3803 1322
rect 2836 1254 2882 1265
rect 3102 1256 3205 1265
rect 2704 1218 2776 1231
rect 3102 1205 3128 1256
rect 3179 1205 3205 1256
rect 3425 1254 3471 1265
rect 3531 1277 3603 1290
rect 3531 1231 3544 1277
rect 3590 1231 3603 1277
rect 3531 1218 3603 1231
rect 3665 1265 3757 1311
rect 2836 1143 2882 1154
rect 2744 1097 2836 1143
rect 2744 1015 2790 1097
rect 2836 1086 2882 1097
rect 3102 1146 3205 1205
rect 3102 1095 3128 1146
rect 3179 1095 3205 1146
rect 2504 975 2550 986
rect 2596 975 2790 1015
rect 3102 1036 3205 1095
rect 3425 1143 3471 1154
rect 3471 1097 3563 1143
rect 3425 1086 3471 1097
rect 2550 969 2790 975
rect 2550 929 2642 969
rect 2504 918 2550 929
rect 2504 807 2550 818
rect 2744 807 2790 969
rect 2836 975 2882 986
rect 3102 985 3128 1036
rect 3179 985 3205 1036
rect 3517 1015 3563 1097
rect 3665 1015 3711 1265
rect 3757 1254 3803 1265
rect 3757 1143 3803 1154
rect 3803 1097 3895 1143
rect 3757 1086 3803 1097
rect 3102 975 3205 985
rect 3425 975 3471 986
rect 2882 929 3425 975
rect 2836 918 2882 929
rect 3102 926 3205 929
rect 3102 875 3128 926
rect 3179 875 3205 926
rect 3425 918 3471 929
rect 3517 975 3711 1015
rect 3757 975 3803 986
rect 3517 969 3757 975
rect 2836 807 2882 818
rect 2412 761 2504 807
rect 2550 761 2642 807
rect 2504 750 2550 761
rect 2504 639 2550 650
rect 2412 593 2504 639
rect 2412 303 2458 593
rect 2504 582 2550 593
rect 2504 471 2550 482
rect 2596 471 2642 761
rect 2550 425 2642 471
rect 2744 761 2836 807
rect 2504 414 2550 425
rect 2504 303 2550 314
rect 2744 303 2790 761
rect 2836 750 2882 761
rect 3102 816 3205 875
rect 3102 765 3128 816
rect 3179 765 3205 816
rect 3102 706 3205 765
rect 3425 807 3471 818
rect 3517 807 3563 969
rect 3665 929 3757 969
rect 3757 918 3803 929
rect 3757 807 3803 818
rect 3849 807 3895 1097
rect 3471 761 3563 807
rect 3425 750 3471 761
rect 3102 655 3128 706
rect 3179 655 3205 706
rect 2836 639 2882 650
rect 2882 593 3001 639
rect 2836 582 2882 593
rect 2942 568 3001 593
rect 3102 596 3205 655
rect 3425 639 3471 650
rect 2942 555 3014 568
rect 3102 555 3128 596
rect 2942 509 2955 555
rect 3001 545 3128 555
rect 3179 555 3205 596
rect 3306 593 3425 639
rect 3306 568 3365 593
rect 3425 582 3471 593
rect 3293 555 3365 568
rect 3179 545 3306 555
rect 3001 509 3306 545
rect 3352 509 3365 555
rect 2942 496 3014 509
rect 2836 471 2882 482
rect 2942 471 3001 496
rect 2882 425 3001 471
rect 3102 486 3205 509
rect 3293 496 3365 509
rect 3102 435 3128 486
rect 3179 435 3205 486
rect 2836 414 2882 425
rect 3102 376 3205 435
rect 3306 471 3365 496
rect 3425 471 3471 482
rect 3306 425 3425 471
rect 3425 414 3471 425
rect 3102 325 3128 376
rect 3179 325 3205 376
rect 2836 303 2882 314
rect 2412 257 2504 303
rect 2550 257 2642 303
rect 2504 246 2550 257
rect 2146 156 2248 214
rect 2294 227 2366 240
rect 2294 181 2307 227
rect 2353 181 2366 227
rect 2294 168 2366 181
rect 2146 104 2173 156
rect 2220 104 2248 156
rect 2504 135 2550 146
rect 2146 46 2248 104
rect 2146 -6 2173 46
rect 2220 -6 2248 46
rect 2146 -64 2248 -6
rect 2146 -116 2173 -64
rect 2220 -116 2248 -64
rect 2146 -174 2248 -116
rect 2146 -226 2173 -174
rect 2220 -201 2248 -174
rect 2412 89 2504 135
rect 2412 -201 2458 89
rect 2504 78 2550 89
rect 2504 -33 2550 -22
rect 2596 -33 2642 257
rect 2744 257 2836 303
rect 2744 143 2790 257
rect 2836 246 2882 257
rect 3102 266 3205 325
rect 3102 215 3128 266
rect 3179 215 3205 266
rect 3425 303 3471 314
rect 3517 303 3563 761
rect 3665 761 3757 807
rect 3803 761 3895 807
rect 3665 471 3711 761
rect 3757 750 3803 761
rect 3757 639 3803 650
rect 3803 593 3895 639
rect 3757 582 3803 593
rect 3757 471 3803 482
rect 3665 425 3757 471
rect 3757 414 3803 425
rect 3757 303 3803 314
rect 3849 303 3895 593
rect 3471 257 3563 303
rect 3425 246 3471 257
rect 3102 156 3205 215
rect 2550 -79 2642 -33
rect 2701 97 2790 143
rect 2836 135 2882 146
rect 2701 -59 2747 97
rect 2882 89 3001 135
rect 2836 78 2882 89
rect 2942 64 3001 89
rect 3102 105 3128 156
rect 3179 105 3205 156
rect 3425 135 3471 146
rect 2942 51 3014 64
rect 3102 51 3205 105
rect 3306 89 3425 135
rect 3517 143 3563 257
rect 3665 257 3757 303
rect 3803 257 3895 303
rect 3517 97 3606 143
rect 3306 64 3365 89
rect 3425 78 3471 89
rect 3293 51 3365 64
rect 2942 5 2955 51
rect 3001 46 3306 51
rect 3001 5 3128 46
rect 2942 -8 3014 5
rect 3102 -5 3128 5
rect 3179 5 3306 46
rect 3352 5 3365 51
rect 3179 -5 3205 5
rect 2836 -33 2882 -22
rect 2942 -33 3001 -8
rect 2688 -72 2760 -59
rect 2504 -90 2550 -79
rect 2688 -118 2701 -72
rect 2747 -118 2760 -72
rect 2882 -79 3001 -33
rect 3102 -64 3205 -5
rect 3293 -8 3365 5
rect 2836 -90 2882 -79
rect 2688 -129 2760 -118
rect 3102 -115 3128 -64
rect 3179 -115 3205 -64
rect 3306 -33 3365 -8
rect 3425 -33 3471 -22
rect 3306 -79 3425 -33
rect 3560 -59 3606 97
rect 3665 -33 3711 257
rect 3757 246 3803 257
rect 3941 240 3987 2205
rect 4059 1366 4162 1393
rect 4059 1314 4087 1366
rect 4134 1314 4162 1366
rect 4059 1256 4162 1314
rect 4059 1204 4087 1256
rect 4134 1204 4162 1256
rect 4059 1146 4162 1204
rect 4059 1094 4087 1146
rect 4134 1094 4162 1146
rect 4059 1036 4162 1094
rect 4059 984 4087 1036
rect 4134 984 4162 1036
rect 4059 926 4162 984
rect 4059 874 4087 926
rect 4134 874 4162 926
rect 4059 816 4162 874
rect 4059 764 4087 816
rect 4134 764 4162 816
rect 4059 706 4162 764
rect 4059 654 4087 706
rect 4134 654 4162 706
rect 4059 596 4162 654
rect 4059 544 4087 596
rect 4134 544 4162 596
rect 4059 486 4162 544
rect 4059 434 4087 486
rect 4134 434 4162 486
rect 4059 376 4162 434
rect 4059 324 4087 376
rect 4134 324 4162 376
rect 4059 266 4162 324
rect 3941 227 4013 240
rect 3941 181 3954 227
rect 4000 181 4013 227
rect 3941 168 4013 181
rect 4059 214 4087 266
rect 4134 214 4162 266
rect 4234 240 4280 2332
rect 5839 2271 5917 2283
rect 5839 2217 5851 2271
rect 5905 2217 5917 2271
rect 5839 2205 5917 2217
rect 5174 2144 5252 2156
rect 5174 2090 5186 2144
rect 5240 2090 5252 2144
rect 5174 2078 5252 2090
rect 4883 2017 4961 2029
rect 4883 1963 4895 2017
rect 4949 1963 4961 2017
rect 4883 1951 4961 1963
rect 4615 1880 4693 1892
rect 4615 1826 4627 1880
rect 4681 1826 4693 1880
rect 4615 1814 4693 1826
rect 4418 1311 4464 1322
rect 4464 1265 4556 1311
rect 4631 1290 4677 1814
rect 4899 1442 4945 1951
rect 5190 1442 5236 2078
rect 5442 1880 5520 1892
rect 5442 1826 5454 1880
rect 5508 1826 5520 1880
rect 5442 1814 5520 1826
rect 4886 1429 4958 1442
rect 4886 1383 4899 1429
rect 4945 1383 4958 1429
rect 5177 1429 5249 1442
rect 4886 1370 4958 1383
rect 5016 1366 5119 1392
rect 5177 1383 5190 1429
rect 5236 1383 5249 1429
rect 5177 1370 5249 1383
rect 4750 1311 4796 1322
rect 5016 1315 5042 1366
rect 5093 1315 5119 1366
rect 5016 1311 5119 1315
rect 5339 1311 5385 1322
rect 4418 1254 4464 1265
rect 4418 1143 4464 1154
rect 4326 1097 4418 1143
rect 4326 807 4372 1097
rect 4418 1086 4464 1097
rect 4510 1015 4556 1265
rect 4618 1277 4690 1290
rect 4618 1231 4631 1277
rect 4677 1231 4690 1277
rect 4796 1265 5339 1311
rect 5458 1290 5504 1814
rect 5671 1311 5717 1322
rect 4750 1254 4796 1265
rect 5016 1256 5119 1265
rect 4618 1218 4690 1231
rect 5016 1205 5042 1256
rect 5093 1205 5119 1256
rect 5339 1254 5385 1265
rect 5445 1277 5517 1290
rect 5445 1231 5458 1277
rect 5504 1231 5517 1277
rect 5445 1218 5517 1231
rect 5579 1265 5671 1311
rect 4750 1143 4796 1154
rect 4658 1097 4750 1143
rect 4658 1015 4704 1097
rect 4750 1086 4796 1097
rect 5016 1146 5119 1205
rect 5016 1095 5042 1146
rect 5093 1095 5119 1146
rect 4418 975 4464 986
rect 4510 975 4704 1015
rect 5016 1036 5119 1095
rect 5339 1143 5385 1154
rect 5385 1097 5477 1143
rect 5339 1086 5385 1097
rect 4464 969 4704 975
rect 4464 929 4556 969
rect 4418 918 4464 929
rect 4418 807 4464 818
rect 4658 807 4704 969
rect 4750 975 4796 986
rect 5016 985 5042 1036
rect 5093 985 5119 1036
rect 5431 1015 5477 1097
rect 5579 1015 5625 1265
rect 5671 1254 5717 1265
rect 5671 1143 5717 1154
rect 5717 1097 5809 1143
rect 5671 1086 5717 1097
rect 5016 975 5119 985
rect 5339 975 5385 986
rect 4796 929 5339 975
rect 4750 918 4796 929
rect 5016 926 5119 929
rect 5016 875 5042 926
rect 5093 875 5119 926
rect 5339 918 5385 929
rect 5431 975 5625 1015
rect 5671 975 5717 986
rect 5431 969 5671 975
rect 4750 807 4796 818
rect 4326 761 4418 807
rect 4464 761 4556 807
rect 4418 750 4464 761
rect 4418 639 4464 650
rect 4326 593 4418 639
rect 4326 303 4372 593
rect 4418 582 4464 593
rect 4418 471 4464 482
rect 4510 471 4556 761
rect 4464 425 4556 471
rect 4658 761 4750 807
rect 4418 414 4464 425
rect 4418 303 4464 314
rect 4658 303 4704 761
rect 4750 750 4796 761
rect 5016 816 5119 875
rect 5016 765 5042 816
rect 5093 765 5119 816
rect 5016 706 5119 765
rect 5339 807 5385 818
rect 5431 807 5477 969
rect 5579 929 5671 969
rect 5671 918 5717 929
rect 5671 807 5717 818
rect 5763 807 5809 1097
rect 5385 761 5477 807
rect 5339 750 5385 761
rect 5016 655 5042 706
rect 5093 655 5119 706
rect 4750 639 4796 650
rect 4796 593 4915 639
rect 4750 582 4796 593
rect 4856 568 4915 593
rect 5016 596 5119 655
rect 5339 639 5385 650
rect 4856 555 4928 568
rect 5016 555 5042 596
rect 4856 509 4869 555
rect 4915 545 5042 555
rect 5093 555 5119 596
rect 5220 593 5339 639
rect 5220 568 5279 593
rect 5339 582 5385 593
rect 5207 555 5279 568
rect 5093 545 5220 555
rect 4915 509 5220 545
rect 5266 509 5279 555
rect 4856 496 4928 509
rect 4750 471 4796 482
rect 4856 471 4915 496
rect 4796 425 4915 471
rect 5016 486 5119 509
rect 5207 496 5279 509
rect 5016 435 5042 486
rect 5093 435 5119 486
rect 4750 414 4796 425
rect 5016 376 5119 435
rect 5220 471 5279 496
rect 5339 471 5385 482
rect 5220 425 5339 471
rect 5339 414 5385 425
rect 5016 325 5042 376
rect 5093 325 5119 376
rect 4750 303 4796 314
rect 4326 257 4418 303
rect 4464 257 4556 303
rect 4418 246 4464 257
rect 4059 156 4162 214
rect 4208 227 4280 240
rect 4208 181 4221 227
rect 4267 181 4280 227
rect 4208 168 4280 181
rect 3757 135 3803 146
rect 3803 89 3895 135
rect 3757 78 3803 89
rect 3757 -33 3803 -22
rect 3425 -90 3471 -79
rect 3547 -72 3619 -59
rect 3102 -174 3205 -115
rect 3547 -118 3560 -72
rect 3606 -118 3619 -72
rect 3665 -79 3757 -33
rect 3757 -90 3803 -79
rect 3547 -129 3619 -118
rect 2504 -201 2550 -190
rect 2836 -201 2882 -190
rect 2220 -226 2504 -201
rect 2146 -247 2504 -226
rect 2146 -284 2248 -247
rect 2504 -258 2550 -247
rect 2742 -247 2836 -201
rect 2146 -336 2173 -284
rect 2220 -336 2248 -284
rect 2146 -394 2248 -336
rect 2504 -369 2550 -358
rect 2742 -369 2788 -247
rect 2836 -258 2882 -247
rect 3102 -225 3128 -174
rect 3179 -225 3205 -174
rect 3102 -284 3205 -225
rect 3425 -201 3471 -190
rect 3757 -201 3803 -190
rect 3849 -201 3895 89
rect 4059 104 4087 156
rect 4134 104 4162 156
rect 4418 135 4464 146
rect 4059 46 4162 104
rect 4059 -6 4087 46
rect 4134 -6 4162 46
rect 4059 -64 4162 -6
rect 4059 -116 4087 -64
rect 4134 -116 4162 -64
rect 4059 -174 4162 -116
rect 4059 -201 4087 -174
rect 3471 -247 3565 -201
rect 3425 -258 3471 -247
rect 3102 -335 3128 -284
rect 3179 -335 3205 -284
rect 2146 -446 2173 -394
rect 2220 -446 2248 -394
rect 2502 -415 2504 -369
rect 2550 -415 2788 -369
rect 2836 -369 2882 -358
rect 3102 -369 3205 -335
rect 3425 -369 3471 -358
rect 2882 -394 3425 -369
rect 2882 -415 3128 -394
rect 2504 -426 2550 -415
rect 2146 -488 2248 -446
rect 1779 -555 1893 -526
rect 2172 -687 2221 -488
rect 2158 -699 2236 -687
rect 2158 -753 2170 -699
rect 2224 -753 2236 -699
rect 2158 -765 2236 -753
rect 2609 -950 2655 -415
rect 2836 -426 2882 -415
rect 3102 -445 3128 -415
rect 3179 -415 3425 -394
rect 3519 -369 3565 -247
rect 3803 -226 4087 -201
rect 4134 -201 4162 -174
rect 4326 89 4418 135
rect 4326 -201 4372 89
rect 4418 78 4464 89
rect 4418 -33 4464 -22
rect 4510 -33 4556 257
rect 4658 257 4750 303
rect 4658 143 4704 257
rect 4750 246 4796 257
rect 5016 266 5119 325
rect 5016 215 5042 266
rect 5093 215 5119 266
rect 5339 303 5385 314
rect 5431 303 5477 761
rect 5579 761 5671 807
rect 5717 761 5809 807
rect 5579 471 5625 761
rect 5671 750 5717 761
rect 5671 639 5717 650
rect 5717 593 5809 639
rect 5671 582 5717 593
rect 5671 471 5717 482
rect 5579 425 5671 471
rect 5671 414 5717 425
rect 5671 303 5717 314
rect 5763 303 5809 593
rect 5385 257 5477 303
rect 5339 246 5385 257
rect 5016 156 5119 215
rect 4464 -79 4556 -33
rect 4615 97 4704 143
rect 4750 135 4796 146
rect 4615 -59 4661 97
rect 4796 89 4915 135
rect 4750 78 4796 89
rect 4856 64 4915 89
rect 5016 105 5042 156
rect 5093 105 5119 156
rect 5339 135 5385 146
rect 4856 51 4928 64
rect 5016 51 5119 105
rect 5220 89 5339 135
rect 5431 143 5477 257
rect 5579 257 5671 303
rect 5717 257 5809 303
rect 5431 97 5520 143
rect 5220 64 5279 89
rect 5339 78 5385 89
rect 5207 51 5279 64
rect 4856 5 4869 51
rect 4915 46 5220 51
rect 4915 5 5042 46
rect 4856 -8 4928 5
rect 5016 -5 5042 5
rect 5093 5 5220 46
rect 5266 5 5279 51
rect 5093 -5 5119 5
rect 4750 -33 4796 -22
rect 4856 -33 4915 -8
rect 4602 -72 4674 -59
rect 4418 -90 4464 -79
rect 4602 -118 4615 -72
rect 4661 -118 4674 -72
rect 4796 -79 4915 -33
rect 5016 -64 5119 -5
rect 5207 -8 5279 5
rect 4750 -90 4796 -79
rect 4602 -129 4674 -118
rect 5016 -115 5042 -64
rect 5093 -115 5119 -64
rect 5220 -33 5279 -8
rect 5339 -33 5385 -22
rect 5220 -79 5339 -33
rect 5474 -59 5520 97
rect 5579 -33 5625 257
rect 5671 246 5717 257
rect 5855 240 5901 2205
rect 5973 1366 6076 1393
rect 5973 1314 6001 1366
rect 6048 1314 6076 1366
rect 5973 1256 6076 1314
rect 5973 1204 6001 1256
rect 6048 1204 6076 1256
rect 5973 1146 6076 1204
rect 5973 1094 6001 1146
rect 6048 1094 6076 1146
rect 5973 1036 6076 1094
rect 5973 984 6001 1036
rect 6048 984 6076 1036
rect 5973 926 6076 984
rect 5973 874 6001 926
rect 6048 874 6076 926
rect 5973 816 6076 874
rect 5973 764 6001 816
rect 6048 764 6076 816
rect 5973 706 6076 764
rect 5973 654 6001 706
rect 6048 654 6076 706
rect 5973 596 6076 654
rect 5973 544 6001 596
rect 6048 544 6076 596
rect 5973 486 6076 544
rect 5973 434 6001 486
rect 6048 434 6076 486
rect 5973 376 6076 434
rect 5973 324 6001 376
rect 6048 324 6076 376
rect 5973 266 6076 324
rect 5855 227 5927 240
rect 5855 181 5868 227
rect 5914 181 5927 227
rect 5855 168 5927 181
rect 5973 214 6001 266
rect 6048 214 6076 266
rect 6148 240 6194 2332
rect 6797 2144 6875 2156
rect 6797 2090 6809 2144
rect 6863 2090 6875 2144
rect 6797 2078 6875 2090
rect 6529 1880 6607 1892
rect 6529 1826 6541 1880
rect 6595 1826 6607 1880
rect 6529 1814 6607 1826
rect 6332 1311 6378 1322
rect 6378 1265 6470 1311
rect 6545 1290 6591 1814
rect 6813 1442 6859 2078
rect 6800 1429 6872 1442
rect 6800 1383 6813 1429
rect 6859 1383 6872 1429
rect 6800 1370 6872 1383
rect 6930 1366 7032 1392
rect 6664 1311 6710 1322
rect 6930 1315 6956 1366
rect 7007 1315 7032 1366
rect 6930 1311 7032 1315
rect 6332 1254 6378 1265
rect 6332 1143 6378 1154
rect 6240 1097 6332 1143
rect 6240 807 6286 1097
rect 6332 1086 6378 1097
rect 6424 1015 6470 1265
rect 6532 1277 6604 1290
rect 6532 1231 6545 1277
rect 6591 1231 6604 1277
rect 6710 1265 7032 1311
rect 6664 1254 6710 1265
rect 6930 1256 7032 1265
rect 6532 1218 6604 1231
rect 6930 1205 6956 1256
rect 7007 1205 7032 1256
rect 6664 1143 6710 1154
rect 6572 1097 6664 1143
rect 6572 1015 6618 1097
rect 6664 1086 6710 1097
rect 6930 1146 7032 1205
rect 6930 1095 6956 1146
rect 7007 1095 7032 1146
rect 6332 975 6378 986
rect 6424 975 6618 1015
rect 6930 1036 7032 1095
rect 6378 969 6618 975
rect 6378 929 6470 969
rect 6332 918 6378 929
rect 6332 807 6378 818
rect 6572 807 6618 969
rect 6664 975 6710 986
rect 6930 985 6956 1036
rect 7007 985 7032 1036
rect 6930 975 7032 985
rect 6710 929 7032 975
rect 6664 918 6710 929
rect 6930 926 7032 929
rect 6930 875 6956 926
rect 7007 875 7032 926
rect 6664 807 6710 818
rect 6240 761 6332 807
rect 6378 761 6470 807
rect 6332 750 6378 761
rect 6332 639 6378 650
rect 6240 593 6332 639
rect 6240 303 6286 593
rect 6332 582 6378 593
rect 6332 471 6378 482
rect 6424 471 6470 761
rect 6378 425 6470 471
rect 6572 761 6664 807
rect 6332 414 6378 425
rect 6332 303 6378 314
rect 6572 303 6618 761
rect 6664 750 6710 761
rect 6930 816 7032 875
rect 6930 765 6956 816
rect 7007 765 7032 816
rect 6930 706 7032 765
rect 6930 655 6956 706
rect 7007 655 7032 706
rect 6664 639 6710 650
rect 6710 593 6829 639
rect 6664 582 6710 593
rect 6770 568 6829 593
rect 6930 596 7032 655
rect 6770 555 6842 568
rect 6930 555 6956 596
rect 6770 509 6783 555
rect 6829 545 6956 555
rect 7007 545 7032 596
rect 6829 509 7032 545
rect 6770 496 6842 509
rect 6664 471 6710 482
rect 6770 471 6829 496
rect 6710 425 6829 471
rect 6930 486 7032 509
rect 6930 435 6956 486
rect 7007 435 7032 486
rect 6664 414 6710 425
rect 6930 376 7032 435
rect 6930 325 6956 376
rect 7007 325 7032 376
rect 6664 303 6710 314
rect 6240 257 6332 303
rect 6378 257 6470 303
rect 6332 246 6378 257
rect 5973 156 6076 214
rect 6122 227 6194 240
rect 6122 181 6135 227
rect 6181 181 6194 227
rect 6122 168 6194 181
rect 5671 135 5717 146
rect 5717 89 5809 135
rect 5671 78 5717 89
rect 5671 -33 5717 -22
rect 5339 -90 5385 -79
rect 5461 -72 5533 -59
rect 5016 -174 5119 -115
rect 5461 -118 5474 -72
rect 5520 -118 5533 -72
rect 5579 -79 5671 -33
rect 5671 -90 5717 -79
rect 5461 -129 5533 -118
rect 4418 -201 4464 -190
rect 4750 -201 4796 -190
rect 4134 -226 4418 -201
rect 3803 -247 4418 -226
rect 3757 -258 3803 -247
rect 4059 -284 4162 -247
rect 4418 -258 4464 -247
rect 4656 -247 4750 -201
rect 4059 -336 4087 -284
rect 4134 -336 4162 -284
rect 3757 -369 3803 -358
rect 3519 -415 3757 -369
rect 3803 -415 3805 -369
rect 4059 -394 4162 -336
rect 4418 -369 4464 -358
rect 4656 -369 4702 -247
rect 4750 -258 4796 -247
rect 5016 -225 5042 -174
rect 5093 -225 5119 -174
rect 5016 -284 5119 -225
rect 5339 -201 5385 -190
rect 5671 -201 5717 -190
rect 5763 -201 5809 89
rect 5973 104 6001 156
rect 6048 104 6076 156
rect 6332 135 6378 146
rect 5973 46 6076 104
rect 5973 -6 6001 46
rect 6048 -6 6076 46
rect 5973 -64 6076 -6
rect 5973 -116 6001 -64
rect 6048 -116 6076 -64
rect 5973 -174 6076 -116
rect 5973 -201 6001 -174
rect 5385 -247 5479 -201
rect 5339 -258 5385 -247
rect 5016 -335 5042 -284
rect 5093 -335 5119 -284
rect 3179 -445 3205 -415
rect 3425 -426 3471 -415
rect 3102 -489 3205 -445
rect 3129 -827 3179 -489
rect 3115 -839 3193 -827
rect 3115 -893 3127 -839
rect 3181 -893 3193 -839
rect 3115 -905 3193 -893
rect 3652 -950 3698 -415
rect 3757 -426 3803 -415
rect 4059 -446 4087 -394
rect 4134 -446 4162 -394
rect 4416 -415 4418 -369
rect 4464 -415 4702 -369
rect 4750 -369 4796 -358
rect 5016 -369 5119 -335
rect 5339 -369 5385 -358
rect 4796 -394 5339 -369
rect 4796 -415 5042 -394
rect 4418 -426 4464 -415
rect 4059 -488 4162 -446
rect 4085 -687 4135 -488
rect 4071 -699 4149 -687
rect 4071 -753 4083 -699
rect 4137 -753 4149 -699
rect 4071 -765 4149 -753
rect 4523 -950 4569 -415
rect 4750 -426 4796 -415
rect 5016 -445 5042 -415
rect 5093 -415 5339 -394
rect 5433 -369 5479 -247
rect 5717 -226 6001 -201
rect 6048 -201 6076 -174
rect 6240 89 6332 135
rect 6240 -201 6286 89
rect 6332 78 6378 89
rect 6332 -33 6378 -22
rect 6424 -33 6470 257
rect 6572 257 6664 303
rect 6572 143 6618 257
rect 6664 246 6710 257
rect 6930 266 7032 325
rect 6930 215 6956 266
rect 7007 215 7032 266
rect 6930 156 7032 215
rect 6378 -79 6470 -33
rect 6529 97 6618 143
rect 6664 135 6710 146
rect 6529 -59 6575 97
rect 6710 89 6829 135
rect 6664 78 6710 89
rect 6770 64 6829 89
rect 6930 105 6956 156
rect 7007 105 7032 156
rect 6770 51 6842 64
rect 6930 51 7032 105
rect 6770 5 6783 51
rect 6829 46 7032 51
rect 6829 5 6956 46
rect 6770 -8 6842 5
rect 6930 -5 6956 5
rect 7007 -5 7032 46
rect 6664 -33 6710 -22
rect 6770 -33 6829 -8
rect 6516 -72 6588 -59
rect 6332 -90 6378 -79
rect 6516 -118 6529 -72
rect 6575 -118 6588 -72
rect 6710 -79 6829 -33
rect 6930 -64 7032 -5
rect 6664 -90 6710 -79
rect 6516 -129 6588 -118
rect 6930 -115 6956 -64
rect 7007 -115 7032 -64
rect 6930 -174 7032 -115
rect 6332 -201 6378 -190
rect 6664 -201 6710 -190
rect 6048 -226 6332 -201
rect 5717 -247 6332 -226
rect 5671 -258 5717 -247
rect 5973 -284 6076 -247
rect 6332 -258 6378 -247
rect 6570 -247 6664 -201
rect 5973 -336 6001 -284
rect 6048 -336 6076 -284
rect 5671 -369 5717 -358
rect 5433 -415 5671 -369
rect 5717 -415 5719 -369
rect 5973 -394 6076 -336
rect 6332 -369 6378 -358
rect 6570 -369 6616 -247
rect 6664 -258 6710 -247
rect 6930 -225 6956 -174
rect 7007 -225 7032 -174
rect 6930 -284 7032 -225
rect 6930 -335 6956 -284
rect 7007 -335 7032 -284
rect 5093 -445 5119 -415
rect 5339 -426 5385 -415
rect 5016 -489 5119 -445
rect 5041 -827 5094 -489
rect 5029 -839 5107 -827
rect 5029 -893 5041 -839
rect 5095 -893 5107 -839
rect 5029 -905 5107 -893
rect 5566 -950 5612 -415
rect 5671 -426 5717 -415
rect 5973 -446 6001 -394
rect 6048 -446 6076 -394
rect 6330 -415 6332 -369
rect 6378 -415 6616 -369
rect 6664 -369 6710 -358
rect 6930 -369 7032 -335
rect 6710 -394 7032 -369
rect 6710 -415 6956 -394
rect 6332 -426 6378 -415
rect 5973 -488 6076 -446
rect 6000 -687 6051 -488
rect 5987 -699 6065 -687
rect 5987 -753 5999 -699
rect 6053 -753 6065 -699
rect 5987 -765 6065 -753
rect 6437 -950 6483 -415
rect 6664 -426 6710 -415
rect 6930 -445 6956 -415
rect 7007 -445 7032 -394
rect 6930 -489 7032 -445
rect 6955 -827 7009 -489
rect 6951 -839 7029 -827
rect 6951 -893 6963 -839
rect 7017 -893 7029 -839
rect 6951 -905 7029 -893
<< via1 >>
rect -595 2344 -541 2398
rect 2316 2344 2370 2398
rect 4230 2344 4284 2398
rect 6142 2344 6196 2398
rect 681 2217 735 2271
rect 1640 2217 1694 2271
rect -499 2089 -445 2143
rect 556 1952 610 2006
rect -405 1826 -351 1880
rect 324 1701 378 1755
rect -405 907 -351 961
rect 54 907 108 961
rect 315 831 369 885
rect 557 875 611 929
rect -499 150 -445 204
rect 50 150 104 204
rect 319 101 373 155
rect 1057 1963 1111 2017
rect 774 1701 828 1755
rect 774 577 828 631
rect 1029 577 1083 631
rect 622 100 676 154
rect -595 -599 -541 -545
rect 50 -600 104 -546
rect -313 -753 -259 -699
rect 447 -893 501 -839
rect 3937 2217 3991 2271
rect 2981 2090 3035 2144
rect 2713 1701 2767 1755
rect 3272 1963 3326 2017
rect 3540 1826 3594 1880
rect 5851 2217 5905 2271
rect 5186 2090 5240 2144
rect 4895 1963 4949 2017
rect 4627 1826 4681 1880
rect 5454 1826 5508 1880
rect 2170 -753 2224 -699
rect 6809 2090 6863 2144
rect 6541 1826 6595 1880
rect 3127 -893 3181 -839
rect 4083 -753 4137 -699
rect 5041 -893 5095 -839
rect 5999 -753 6053 -699
rect 6963 -893 7017 -839
<< metal2 >>
rect -607 2399 -529 2410
rect 2304 2399 2382 2410
rect 4218 2399 4296 2410
rect 6130 2399 6208 2410
rect -647 2398 7057 2399
rect -647 2344 -595 2398
rect -541 2344 2316 2398
rect 2370 2344 4230 2398
rect 4284 2344 6142 2398
rect 6196 2344 7057 2398
rect -647 2343 7057 2344
rect -607 2332 -529 2343
rect 2304 2332 2382 2343
rect 4218 2332 4296 2343
rect 6130 2332 6208 2343
rect 669 2272 747 2283
rect 1628 2272 1706 2283
rect 3925 2272 4003 2283
rect 5839 2272 5917 2283
rect -647 2271 7057 2272
rect -647 2217 681 2271
rect 735 2217 1640 2271
rect 1694 2217 3937 2271
rect 3991 2217 5851 2271
rect 5905 2217 7057 2271
rect -647 2216 7057 2217
rect 669 2205 747 2216
rect 1628 2205 1706 2216
rect 3925 2205 4003 2216
rect 5839 2205 5917 2216
rect -511 2145 -433 2155
rect 2969 2145 3047 2156
rect 5174 2145 5252 2156
rect 6797 2145 6875 2156
rect -647 2144 7057 2145
rect -647 2143 2981 2144
rect -647 2089 -499 2143
rect -445 2090 2981 2143
rect 3035 2090 5186 2144
rect 5240 2090 6809 2144
rect 6863 2090 7057 2144
rect -445 2089 7057 2090
rect -511 2077 -433 2089
rect 2969 2078 3047 2089
rect 5174 2078 5252 2089
rect 6797 2078 6875 2089
rect 1045 2018 1123 2029
rect 3260 2018 3338 2029
rect 4883 2018 4961 2029
rect -647 2017 7057 2018
rect -647 2006 1057 2017
rect -647 1962 556 2006
rect 544 1952 556 1962
rect 610 1963 1057 2006
rect 1111 1963 3272 2017
rect 3326 1963 4895 2017
rect 4949 1963 7057 2017
rect 610 1962 7057 1963
rect 610 1952 622 1962
rect 544 1940 622 1952
rect 1045 1951 1123 1962
rect 3260 1951 3338 1962
rect 4883 1951 4961 1962
rect -417 1881 -339 1892
rect 3528 1881 3606 1892
rect 4615 1881 4693 1892
rect 5442 1881 5520 1892
rect 6529 1881 6607 1892
rect -647 1880 7057 1881
rect -647 1826 -405 1880
rect -351 1826 3540 1880
rect 3594 1826 4627 1880
rect 4681 1826 5454 1880
rect 5508 1826 6541 1880
rect 6595 1826 7057 1880
rect -647 1825 7057 1826
rect -417 1814 -339 1825
rect 3528 1814 3606 1825
rect 4615 1814 4693 1825
rect 5442 1814 5520 1825
rect 6529 1814 6607 1825
rect 312 1756 390 1767
rect 762 1756 840 1767
rect 2701 1756 2779 1767
rect -647 1755 7057 1756
rect -647 1701 324 1755
rect 378 1701 774 1755
rect 828 1701 2713 1755
rect 2767 1701 7057 1755
rect -647 1700 7057 1701
rect 312 1689 390 1700
rect 762 1689 840 1700
rect 2701 1689 2779 1700
rect -417 962 -339 973
rect 42 962 120 973
rect -417 961 120 962
rect -417 907 -405 961
rect -351 907 54 961
rect 108 907 120 961
rect -417 906 120 907
rect -417 895 -339 906
rect 42 895 120 906
rect 545 929 623 941
rect 303 885 381 897
rect 545 885 557 929
rect 303 831 315 885
rect 369 875 557 885
rect 611 875 623 929
rect 369 831 623 875
rect 303 829 623 831
rect 303 819 381 829
rect 762 632 840 643
rect 1017 632 1095 643
rect 762 631 1095 632
rect 762 577 774 631
rect 828 577 1029 631
rect 1083 577 1095 631
rect 762 576 1095 577
rect 762 565 840 576
rect 1017 565 1095 576
rect -511 205 -433 216
rect 38 205 116 216
rect -511 204 116 205
rect -511 150 -499 204
rect -445 150 50 204
rect 104 150 116 204
rect -511 149 116 150
rect -511 138 -433 149
rect 38 138 116 149
rect 310 155 375 167
rect 610 155 688 166
rect 310 101 319 155
rect 373 154 688 155
rect 373 101 622 154
rect 310 100 622 101
rect 676 100 688 154
rect 310 99 688 100
rect 310 89 375 99
rect 610 88 688 99
rect -607 -545 -529 -533
rect 38 -545 116 -534
rect -607 -599 -595 -545
rect -541 -546 116 -545
rect -541 -599 50 -546
rect -607 -600 50 -599
rect 104 -600 116 -546
rect -607 -601 116 -600
rect -607 -611 -529 -601
rect 38 -612 116 -601
rect -325 -691 -247 -687
rect 2158 -691 2236 -687
rect 4071 -691 4149 -687
rect 5987 -691 6065 -687
rect -647 -699 7055 -691
rect -647 -753 -313 -699
rect -259 -753 2170 -699
rect 2224 -753 4083 -699
rect 4137 -753 5999 -699
rect 6053 -753 7055 -699
rect -647 -761 7055 -753
rect -325 -765 -247 -761
rect 2158 -765 2236 -761
rect 4071 -765 4149 -761
rect 5987 -765 6065 -761
rect 435 -831 513 -827
rect 3115 -831 3193 -827
rect 5029 -831 5107 -827
rect 6951 -831 7029 -827
rect -647 -839 7055 -831
rect -647 -893 447 -839
rect 501 -893 3127 -839
rect 3181 -893 5041 -839
rect 5095 -893 6963 -839
rect 7017 -893 7055 -839
rect -647 -901 7055 -893
rect 435 -905 513 -901
rect 3115 -905 3193 -901
rect 5029 -905 5107 -901
rect 6951 -905 7029 -901
<< labels >>
flabel metal2 7015 1730 7015 1730 0 FreeSans 480 90 0 0 A
port 1 nsew
flabel metal2 7014 1992 7014 1992 0 FreeSans 480 90 0 0 B
port 3 nsew
flabel metal2 7017 2249 7017 2249 0 FreeSans 480 90 0 0 C
port 5 nsew
flabel metal2 7040 -871 7040 -871 0 FreeSans 480 90 0 0 VDD
port 7 nsew
flabel metal2 6885 -728 6885 -728 0 FreeSans 480 90 0 0 VSS
port 11 nsew
flabel metal1 6462 -926 6462 -926 0 FreeSans 400 90 0 0 S1
port 13 nsew
flabel metal1 5590 -926 5590 -926 0 FreeSans 400 90 0 0 S2
port 15 nsew
flabel metal1 4547 -927 4547 -927 0 FreeSans 400 90 0 0 S3
port 17 nsew
flabel metal1 3677 -927 3677 -927 0 FreeSans 400 90 0 0 S4
port 19 nsew
flabel metal1 2633 -926 2633 -926 0 FreeSans 400 90 0 0 S5
port 21 nsew
flabel metal1 1296 -925 1296 -925 0 FreeSans 400 90 0 0 S6
port 23 nsew
flabel metal1 1495 587 1495 587 0 FreeSans 800 90 0 0 AND_1.A
flabel metal1 1067 556 1067 556 0 FreeSans 800 90 0 0 AND_1.B
flabel metal1 1297 -520 1297 -520 0 FreeSans 320 90 0 0 AND_1.OUT
flabel nsubdiffcont 900 159 900 159 0 FreeSans 320 90 0 0 AND_1.VDD
flabel metal1 1833 123 1833 123 0 FreeSans 320 90 0 0 AND_1.VSS
flabel metal1 350 1615 350 1615 0 FreeSans 480 90 0 0 INVERTER_magic_0.IN
flabel metal1 81 1052 81 1052 0 FreeSans 480 90 0 0 INVERTER_magic_0.OUT
flabel nsubdiffcont 475 1319 475 1319 0 FreeSans 480 90 0 0 INVERTER_magic_0.VDD
flabel psubdiffcont -283 1319 -283 1319 0 FreeSans 480 90 0 0 INVERTER_magic_0.VSS
flabel via1 346 104 346 104 0 FreeSans 480 90 0 0 INVERTER_magic_1.IN
flabel metal1 77 -459 77 -459 0 FreeSans 480 90 0 0 INVERTER_magic_1.OUT
flabel nsubdiffcont 471 -192 471 -192 0 FreeSans 480 90 0 0 INVERTER_magic_1.VDD
flabel psubdiffcont -287 -192 -287 -192 0 FreeSans 480 90 0 0 INVERTER_magic_1.VSS
flabel via1 346 859 346 859 0 FreeSans 480 90 0 0 INVERTER_magic_2.IN
flabel metal1 77 296 77 296 0 FreeSans 480 90 0 0 INVERTER_magic_2.OUT
flabel nsubdiffcont 471 563 471 563 0 FreeSans 480 90 0 0 INVERTER_magic_2.VDD
flabel psubdiffcont -287 563 -287 563 0 FreeSans 480 90 0 0 INVERTER_magic_2.VSS
flabel metal1 1086 1660 1086 1660 0 FreeSans 320 90 0 0 OR_magic_1.A
flabel metal1 1663 1657 1663 1657 0 FreeSans 320 90 0 0 OR_magic_1.B
flabel metal1 1316 768 1316 768 0 FreeSans 320 90 0 0 OR_magic_1.OUT
flabel nsubdiffcont 916 1155 916 1155 0 FreeSans 480 90 0 0 OR_magic_1.VDD
flabel psubdiffcont 2043 1155 2043 1155 0 FreeSans 480 90 0 0 OR_magic_1.VSS
flabel metal1 3009 1504 3009 1504 0 FreeSans 480 90 0 0 AND_3_magic_5.B
flabel metal1 2628 -431 2628 -431 0 FreeSans 480 90 0 0 AND_3_magic_5.OUT
flabel nsubdiffcont 3155 459 3155 459 0 FreeSans 480 90 0 0 AND_3_magic_5.VDD
flabel metal1 2342 1502 2342 1502 0 FreeSans 480 90 0 0 AND_3_magic_5.C
flabel psubdiffcont 2200 461 2200 461 0 FreeSans 480 90 0 0 AND_3_magic_5.VSS
flabel metal1 2743 1501 2743 1501 0 FreeSans 480 90 0 0 AND_3_magic_5.A
flabel metal1 3298 1504 3298 1504 0 FreeSans 480 90 0 0 AND_3_magic_2.B
flabel metal1 3679 -431 3679 -431 0 FreeSans 480 90 0 0 AND_3_magic_2.OUT
flabel nsubdiffcont 3152 459 3152 459 0 FreeSans 480 90 0 0 AND_3_magic_2.VDD
flabel metal1 3965 1502 3965 1502 0 FreeSans 480 90 0 0 AND_3_magic_2.C
flabel psubdiffcont 4107 461 4107 461 0 FreeSans 480 90 0 0 AND_3_magic_2.VSS
flabel metal1 3564 1501 3564 1501 0 FreeSans 480 90 0 0 AND_3_magic_2.A
flabel metal1 4923 1504 4923 1504 0 FreeSans 480 90 0 0 AND_3_magic_3.B
flabel metal1 4542 -431 4542 -431 0 FreeSans 480 90 0 0 AND_3_magic_3.OUT
flabel nsubdiffcont 5069 459 5069 459 0 FreeSans 480 90 0 0 AND_3_magic_3.VDD
flabel metal1 4256 1502 4256 1502 0 FreeSans 480 90 0 0 AND_3_magic_3.C
flabel psubdiffcont 4114 461 4114 461 0 FreeSans 480 90 0 0 AND_3_magic_3.VSS
flabel metal1 4657 1501 4657 1501 0 FreeSans 480 90 0 0 AND_3_magic_3.A
flabel metal1 5212 1504 5212 1504 0 FreeSans 480 90 0 0 AND_3_magic_0.B
flabel metal1 5593 -431 5593 -431 0 FreeSans 480 90 0 0 AND_3_magic_0.OUT
flabel nsubdiffcont 5066 459 5066 459 0 FreeSans 480 90 0 0 AND_3_magic_0.VDD
flabel metal1 5879 1502 5879 1502 0 FreeSans 480 90 0 0 AND_3_magic_0.C
flabel psubdiffcont 6021 461 6021 461 0 FreeSans 480 90 0 0 AND_3_magic_0.VSS
flabel metal1 5478 1501 5478 1501 0 FreeSans 480 90 0 0 AND_3_magic_0.A
flabel metal1 6837 1504 6837 1504 0 FreeSans 480 90 0 0 AND_3_magic_1.B
flabel metal1 6456 -431 6456 -431 0 FreeSans 480 90 0 0 AND_3_magic_1.OUT
flabel nsubdiffcont 6983 459 6983 459 0 FreeSans 480 90 0 0 AND_3_magic_1.VDD
flabel metal1 6170 1502 6170 1502 0 FreeSans 480 90 0 0 AND_3_magic_1.C
flabel psubdiffcont 6028 461 6028 461 0 FreeSans 480 90 0 0 AND_3_magic_1.VSS
flabel metal1 6571 1501 6571 1501 0 FreeSans 480 90 0 0 AND_3_magic_1.A
<< end >>
