magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -9237 -2107 9237 2107
<< psubdiff >>
rect -7237 85 7237 107
rect -7237 39 -7215 85
rect -7169 39 -7091 85
rect -7045 39 -6967 85
rect -6921 39 -6843 85
rect -6797 39 -6719 85
rect -6673 39 -6595 85
rect -6549 39 -6471 85
rect -6425 39 -6347 85
rect -6301 39 -6223 85
rect -6177 39 -6099 85
rect -6053 39 -5975 85
rect -5929 39 -5851 85
rect -5805 39 -5727 85
rect -5681 39 -5603 85
rect -5557 39 -5479 85
rect -5433 39 -5355 85
rect -5309 39 -5231 85
rect -5185 39 -5107 85
rect -5061 39 -4983 85
rect -4937 39 -4859 85
rect -4813 39 -4735 85
rect -4689 39 -4611 85
rect -4565 39 -4487 85
rect -4441 39 -4363 85
rect -4317 39 -4239 85
rect -4193 39 -4115 85
rect -4069 39 -3991 85
rect -3945 39 -3867 85
rect -3821 39 -3743 85
rect -3697 39 -3619 85
rect -3573 39 -3495 85
rect -3449 39 -3371 85
rect -3325 39 -3247 85
rect -3201 39 -3123 85
rect -3077 39 -2999 85
rect -2953 39 -2875 85
rect -2829 39 -2751 85
rect -2705 39 -2627 85
rect -2581 39 -2503 85
rect -2457 39 -2379 85
rect -2333 39 -2255 85
rect -2209 39 -2131 85
rect -2085 39 -2007 85
rect -1961 39 -1883 85
rect -1837 39 -1759 85
rect -1713 39 -1635 85
rect -1589 39 -1511 85
rect -1465 39 -1387 85
rect -1341 39 -1263 85
rect -1217 39 -1139 85
rect -1093 39 -1015 85
rect -969 39 -891 85
rect -845 39 -767 85
rect -721 39 -643 85
rect -597 39 -519 85
rect -473 39 -395 85
rect -349 39 -271 85
rect -225 39 -147 85
rect -101 39 -23 85
rect 23 39 101 85
rect 147 39 225 85
rect 271 39 349 85
rect 395 39 473 85
rect 519 39 597 85
rect 643 39 721 85
rect 767 39 845 85
rect 891 39 969 85
rect 1015 39 1093 85
rect 1139 39 1217 85
rect 1263 39 1341 85
rect 1387 39 1465 85
rect 1511 39 1589 85
rect 1635 39 1713 85
rect 1759 39 1837 85
rect 1883 39 1961 85
rect 2007 39 2085 85
rect 2131 39 2209 85
rect 2255 39 2333 85
rect 2379 39 2457 85
rect 2503 39 2581 85
rect 2627 39 2705 85
rect 2751 39 2829 85
rect 2875 39 2953 85
rect 2999 39 3077 85
rect 3123 39 3201 85
rect 3247 39 3325 85
rect 3371 39 3449 85
rect 3495 39 3573 85
rect 3619 39 3697 85
rect 3743 39 3821 85
rect 3867 39 3945 85
rect 3991 39 4069 85
rect 4115 39 4193 85
rect 4239 39 4317 85
rect 4363 39 4441 85
rect 4487 39 4565 85
rect 4611 39 4689 85
rect 4735 39 4813 85
rect 4859 39 4937 85
rect 4983 39 5061 85
rect 5107 39 5185 85
rect 5231 39 5309 85
rect 5355 39 5433 85
rect 5479 39 5557 85
rect 5603 39 5681 85
rect 5727 39 5805 85
rect 5851 39 5929 85
rect 5975 39 6053 85
rect 6099 39 6177 85
rect 6223 39 6301 85
rect 6347 39 6425 85
rect 6471 39 6549 85
rect 6595 39 6673 85
rect 6719 39 6797 85
rect 6843 39 6921 85
rect 6967 39 7045 85
rect 7091 39 7169 85
rect 7215 39 7237 85
rect -7237 -39 7237 39
rect -7237 -85 -7215 -39
rect -7169 -85 -7091 -39
rect -7045 -85 -6967 -39
rect -6921 -85 -6843 -39
rect -6797 -85 -6719 -39
rect -6673 -85 -6595 -39
rect -6549 -85 -6471 -39
rect -6425 -85 -6347 -39
rect -6301 -85 -6223 -39
rect -6177 -85 -6099 -39
rect -6053 -85 -5975 -39
rect -5929 -85 -5851 -39
rect -5805 -85 -5727 -39
rect -5681 -85 -5603 -39
rect -5557 -85 -5479 -39
rect -5433 -85 -5355 -39
rect -5309 -85 -5231 -39
rect -5185 -85 -5107 -39
rect -5061 -85 -4983 -39
rect -4937 -85 -4859 -39
rect -4813 -85 -4735 -39
rect -4689 -85 -4611 -39
rect -4565 -85 -4487 -39
rect -4441 -85 -4363 -39
rect -4317 -85 -4239 -39
rect -4193 -85 -4115 -39
rect -4069 -85 -3991 -39
rect -3945 -85 -3867 -39
rect -3821 -85 -3743 -39
rect -3697 -85 -3619 -39
rect -3573 -85 -3495 -39
rect -3449 -85 -3371 -39
rect -3325 -85 -3247 -39
rect -3201 -85 -3123 -39
rect -3077 -85 -2999 -39
rect -2953 -85 -2875 -39
rect -2829 -85 -2751 -39
rect -2705 -85 -2627 -39
rect -2581 -85 -2503 -39
rect -2457 -85 -2379 -39
rect -2333 -85 -2255 -39
rect -2209 -85 -2131 -39
rect -2085 -85 -2007 -39
rect -1961 -85 -1883 -39
rect -1837 -85 -1759 -39
rect -1713 -85 -1635 -39
rect -1589 -85 -1511 -39
rect -1465 -85 -1387 -39
rect -1341 -85 -1263 -39
rect -1217 -85 -1139 -39
rect -1093 -85 -1015 -39
rect -969 -85 -891 -39
rect -845 -85 -767 -39
rect -721 -85 -643 -39
rect -597 -85 -519 -39
rect -473 -85 -395 -39
rect -349 -85 -271 -39
rect -225 -85 -147 -39
rect -101 -85 -23 -39
rect 23 -85 101 -39
rect 147 -85 225 -39
rect 271 -85 349 -39
rect 395 -85 473 -39
rect 519 -85 597 -39
rect 643 -85 721 -39
rect 767 -85 845 -39
rect 891 -85 969 -39
rect 1015 -85 1093 -39
rect 1139 -85 1217 -39
rect 1263 -85 1341 -39
rect 1387 -85 1465 -39
rect 1511 -85 1589 -39
rect 1635 -85 1713 -39
rect 1759 -85 1837 -39
rect 1883 -85 1961 -39
rect 2007 -85 2085 -39
rect 2131 -85 2209 -39
rect 2255 -85 2333 -39
rect 2379 -85 2457 -39
rect 2503 -85 2581 -39
rect 2627 -85 2705 -39
rect 2751 -85 2829 -39
rect 2875 -85 2953 -39
rect 2999 -85 3077 -39
rect 3123 -85 3201 -39
rect 3247 -85 3325 -39
rect 3371 -85 3449 -39
rect 3495 -85 3573 -39
rect 3619 -85 3697 -39
rect 3743 -85 3821 -39
rect 3867 -85 3945 -39
rect 3991 -85 4069 -39
rect 4115 -85 4193 -39
rect 4239 -85 4317 -39
rect 4363 -85 4441 -39
rect 4487 -85 4565 -39
rect 4611 -85 4689 -39
rect 4735 -85 4813 -39
rect 4859 -85 4937 -39
rect 4983 -85 5061 -39
rect 5107 -85 5185 -39
rect 5231 -85 5309 -39
rect 5355 -85 5433 -39
rect 5479 -85 5557 -39
rect 5603 -85 5681 -39
rect 5727 -85 5805 -39
rect 5851 -85 5929 -39
rect 5975 -85 6053 -39
rect 6099 -85 6177 -39
rect 6223 -85 6301 -39
rect 6347 -85 6425 -39
rect 6471 -85 6549 -39
rect 6595 -85 6673 -39
rect 6719 -85 6797 -39
rect 6843 -85 6921 -39
rect 6967 -85 7045 -39
rect 7091 -85 7169 -39
rect 7215 -85 7237 -39
rect -7237 -107 7237 -85
<< psubdiffcont >>
rect -7215 39 -7169 85
rect -7091 39 -7045 85
rect -6967 39 -6921 85
rect -6843 39 -6797 85
rect -6719 39 -6673 85
rect -6595 39 -6549 85
rect -6471 39 -6425 85
rect -6347 39 -6301 85
rect -6223 39 -6177 85
rect -6099 39 -6053 85
rect -5975 39 -5929 85
rect -5851 39 -5805 85
rect -5727 39 -5681 85
rect -5603 39 -5557 85
rect -5479 39 -5433 85
rect -5355 39 -5309 85
rect -5231 39 -5185 85
rect -5107 39 -5061 85
rect -4983 39 -4937 85
rect -4859 39 -4813 85
rect -4735 39 -4689 85
rect -4611 39 -4565 85
rect -4487 39 -4441 85
rect -4363 39 -4317 85
rect -4239 39 -4193 85
rect -4115 39 -4069 85
rect -3991 39 -3945 85
rect -3867 39 -3821 85
rect -3743 39 -3697 85
rect -3619 39 -3573 85
rect -3495 39 -3449 85
rect -3371 39 -3325 85
rect -3247 39 -3201 85
rect -3123 39 -3077 85
rect -2999 39 -2953 85
rect -2875 39 -2829 85
rect -2751 39 -2705 85
rect -2627 39 -2581 85
rect -2503 39 -2457 85
rect -2379 39 -2333 85
rect -2255 39 -2209 85
rect -2131 39 -2085 85
rect -2007 39 -1961 85
rect -1883 39 -1837 85
rect -1759 39 -1713 85
rect -1635 39 -1589 85
rect -1511 39 -1465 85
rect -1387 39 -1341 85
rect -1263 39 -1217 85
rect -1139 39 -1093 85
rect -1015 39 -969 85
rect -891 39 -845 85
rect -767 39 -721 85
rect -643 39 -597 85
rect -519 39 -473 85
rect -395 39 -349 85
rect -271 39 -225 85
rect -147 39 -101 85
rect -23 39 23 85
rect 101 39 147 85
rect 225 39 271 85
rect 349 39 395 85
rect 473 39 519 85
rect 597 39 643 85
rect 721 39 767 85
rect 845 39 891 85
rect 969 39 1015 85
rect 1093 39 1139 85
rect 1217 39 1263 85
rect 1341 39 1387 85
rect 1465 39 1511 85
rect 1589 39 1635 85
rect 1713 39 1759 85
rect 1837 39 1883 85
rect 1961 39 2007 85
rect 2085 39 2131 85
rect 2209 39 2255 85
rect 2333 39 2379 85
rect 2457 39 2503 85
rect 2581 39 2627 85
rect 2705 39 2751 85
rect 2829 39 2875 85
rect 2953 39 2999 85
rect 3077 39 3123 85
rect 3201 39 3247 85
rect 3325 39 3371 85
rect 3449 39 3495 85
rect 3573 39 3619 85
rect 3697 39 3743 85
rect 3821 39 3867 85
rect 3945 39 3991 85
rect 4069 39 4115 85
rect 4193 39 4239 85
rect 4317 39 4363 85
rect 4441 39 4487 85
rect 4565 39 4611 85
rect 4689 39 4735 85
rect 4813 39 4859 85
rect 4937 39 4983 85
rect 5061 39 5107 85
rect 5185 39 5231 85
rect 5309 39 5355 85
rect 5433 39 5479 85
rect 5557 39 5603 85
rect 5681 39 5727 85
rect 5805 39 5851 85
rect 5929 39 5975 85
rect 6053 39 6099 85
rect 6177 39 6223 85
rect 6301 39 6347 85
rect 6425 39 6471 85
rect 6549 39 6595 85
rect 6673 39 6719 85
rect 6797 39 6843 85
rect 6921 39 6967 85
rect 7045 39 7091 85
rect 7169 39 7215 85
rect -7215 -85 -7169 -39
rect -7091 -85 -7045 -39
rect -6967 -85 -6921 -39
rect -6843 -85 -6797 -39
rect -6719 -85 -6673 -39
rect -6595 -85 -6549 -39
rect -6471 -85 -6425 -39
rect -6347 -85 -6301 -39
rect -6223 -85 -6177 -39
rect -6099 -85 -6053 -39
rect -5975 -85 -5929 -39
rect -5851 -85 -5805 -39
rect -5727 -85 -5681 -39
rect -5603 -85 -5557 -39
rect -5479 -85 -5433 -39
rect -5355 -85 -5309 -39
rect -5231 -85 -5185 -39
rect -5107 -85 -5061 -39
rect -4983 -85 -4937 -39
rect -4859 -85 -4813 -39
rect -4735 -85 -4689 -39
rect -4611 -85 -4565 -39
rect -4487 -85 -4441 -39
rect -4363 -85 -4317 -39
rect -4239 -85 -4193 -39
rect -4115 -85 -4069 -39
rect -3991 -85 -3945 -39
rect -3867 -85 -3821 -39
rect -3743 -85 -3697 -39
rect -3619 -85 -3573 -39
rect -3495 -85 -3449 -39
rect -3371 -85 -3325 -39
rect -3247 -85 -3201 -39
rect -3123 -85 -3077 -39
rect -2999 -85 -2953 -39
rect -2875 -85 -2829 -39
rect -2751 -85 -2705 -39
rect -2627 -85 -2581 -39
rect -2503 -85 -2457 -39
rect -2379 -85 -2333 -39
rect -2255 -85 -2209 -39
rect -2131 -85 -2085 -39
rect -2007 -85 -1961 -39
rect -1883 -85 -1837 -39
rect -1759 -85 -1713 -39
rect -1635 -85 -1589 -39
rect -1511 -85 -1465 -39
rect -1387 -85 -1341 -39
rect -1263 -85 -1217 -39
rect -1139 -85 -1093 -39
rect -1015 -85 -969 -39
rect -891 -85 -845 -39
rect -767 -85 -721 -39
rect -643 -85 -597 -39
rect -519 -85 -473 -39
rect -395 -85 -349 -39
rect -271 -85 -225 -39
rect -147 -85 -101 -39
rect -23 -85 23 -39
rect 101 -85 147 -39
rect 225 -85 271 -39
rect 349 -85 395 -39
rect 473 -85 519 -39
rect 597 -85 643 -39
rect 721 -85 767 -39
rect 845 -85 891 -39
rect 969 -85 1015 -39
rect 1093 -85 1139 -39
rect 1217 -85 1263 -39
rect 1341 -85 1387 -39
rect 1465 -85 1511 -39
rect 1589 -85 1635 -39
rect 1713 -85 1759 -39
rect 1837 -85 1883 -39
rect 1961 -85 2007 -39
rect 2085 -85 2131 -39
rect 2209 -85 2255 -39
rect 2333 -85 2379 -39
rect 2457 -85 2503 -39
rect 2581 -85 2627 -39
rect 2705 -85 2751 -39
rect 2829 -85 2875 -39
rect 2953 -85 2999 -39
rect 3077 -85 3123 -39
rect 3201 -85 3247 -39
rect 3325 -85 3371 -39
rect 3449 -85 3495 -39
rect 3573 -85 3619 -39
rect 3697 -85 3743 -39
rect 3821 -85 3867 -39
rect 3945 -85 3991 -39
rect 4069 -85 4115 -39
rect 4193 -85 4239 -39
rect 4317 -85 4363 -39
rect 4441 -85 4487 -39
rect 4565 -85 4611 -39
rect 4689 -85 4735 -39
rect 4813 -85 4859 -39
rect 4937 -85 4983 -39
rect 5061 -85 5107 -39
rect 5185 -85 5231 -39
rect 5309 -85 5355 -39
rect 5433 -85 5479 -39
rect 5557 -85 5603 -39
rect 5681 -85 5727 -39
rect 5805 -85 5851 -39
rect 5929 -85 5975 -39
rect 6053 -85 6099 -39
rect 6177 -85 6223 -39
rect 6301 -85 6347 -39
rect 6425 -85 6471 -39
rect 6549 -85 6595 -39
rect 6673 -85 6719 -39
rect 6797 -85 6843 -39
rect 6921 -85 6967 -39
rect 7045 -85 7091 -39
rect 7169 -85 7215 -39
<< metal1 >>
rect -7226 85 7226 96
rect -7226 39 -7215 85
rect -7169 39 -7091 85
rect -7045 39 -6967 85
rect -6921 39 -6843 85
rect -6797 39 -6719 85
rect -6673 39 -6595 85
rect -6549 39 -6471 85
rect -6425 39 -6347 85
rect -6301 39 -6223 85
rect -6177 39 -6099 85
rect -6053 39 -5975 85
rect -5929 39 -5851 85
rect -5805 39 -5727 85
rect -5681 39 -5603 85
rect -5557 39 -5479 85
rect -5433 39 -5355 85
rect -5309 39 -5231 85
rect -5185 39 -5107 85
rect -5061 39 -4983 85
rect -4937 39 -4859 85
rect -4813 39 -4735 85
rect -4689 39 -4611 85
rect -4565 39 -4487 85
rect -4441 39 -4363 85
rect -4317 39 -4239 85
rect -4193 39 -4115 85
rect -4069 39 -3991 85
rect -3945 39 -3867 85
rect -3821 39 -3743 85
rect -3697 39 -3619 85
rect -3573 39 -3495 85
rect -3449 39 -3371 85
rect -3325 39 -3247 85
rect -3201 39 -3123 85
rect -3077 39 -2999 85
rect -2953 39 -2875 85
rect -2829 39 -2751 85
rect -2705 39 -2627 85
rect -2581 39 -2503 85
rect -2457 39 -2379 85
rect -2333 39 -2255 85
rect -2209 39 -2131 85
rect -2085 39 -2007 85
rect -1961 39 -1883 85
rect -1837 39 -1759 85
rect -1713 39 -1635 85
rect -1589 39 -1511 85
rect -1465 39 -1387 85
rect -1341 39 -1263 85
rect -1217 39 -1139 85
rect -1093 39 -1015 85
rect -969 39 -891 85
rect -845 39 -767 85
rect -721 39 -643 85
rect -597 39 -519 85
rect -473 39 -395 85
rect -349 39 -271 85
rect -225 39 -147 85
rect -101 39 -23 85
rect 23 39 101 85
rect 147 39 225 85
rect 271 39 349 85
rect 395 39 473 85
rect 519 39 597 85
rect 643 39 721 85
rect 767 39 845 85
rect 891 39 969 85
rect 1015 39 1093 85
rect 1139 39 1217 85
rect 1263 39 1341 85
rect 1387 39 1465 85
rect 1511 39 1589 85
rect 1635 39 1713 85
rect 1759 39 1837 85
rect 1883 39 1961 85
rect 2007 39 2085 85
rect 2131 39 2209 85
rect 2255 39 2333 85
rect 2379 39 2457 85
rect 2503 39 2581 85
rect 2627 39 2705 85
rect 2751 39 2829 85
rect 2875 39 2953 85
rect 2999 39 3077 85
rect 3123 39 3201 85
rect 3247 39 3325 85
rect 3371 39 3449 85
rect 3495 39 3573 85
rect 3619 39 3697 85
rect 3743 39 3821 85
rect 3867 39 3945 85
rect 3991 39 4069 85
rect 4115 39 4193 85
rect 4239 39 4317 85
rect 4363 39 4441 85
rect 4487 39 4565 85
rect 4611 39 4689 85
rect 4735 39 4813 85
rect 4859 39 4937 85
rect 4983 39 5061 85
rect 5107 39 5185 85
rect 5231 39 5309 85
rect 5355 39 5433 85
rect 5479 39 5557 85
rect 5603 39 5681 85
rect 5727 39 5805 85
rect 5851 39 5929 85
rect 5975 39 6053 85
rect 6099 39 6177 85
rect 6223 39 6301 85
rect 6347 39 6425 85
rect 6471 39 6549 85
rect 6595 39 6673 85
rect 6719 39 6797 85
rect 6843 39 6921 85
rect 6967 39 7045 85
rect 7091 39 7169 85
rect 7215 39 7226 85
rect -7226 -39 7226 39
rect -7226 -85 -7215 -39
rect -7169 -85 -7091 -39
rect -7045 -85 -6967 -39
rect -6921 -85 -6843 -39
rect -6797 -85 -6719 -39
rect -6673 -85 -6595 -39
rect -6549 -85 -6471 -39
rect -6425 -85 -6347 -39
rect -6301 -85 -6223 -39
rect -6177 -85 -6099 -39
rect -6053 -85 -5975 -39
rect -5929 -85 -5851 -39
rect -5805 -85 -5727 -39
rect -5681 -85 -5603 -39
rect -5557 -85 -5479 -39
rect -5433 -85 -5355 -39
rect -5309 -85 -5231 -39
rect -5185 -85 -5107 -39
rect -5061 -85 -4983 -39
rect -4937 -85 -4859 -39
rect -4813 -85 -4735 -39
rect -4689 -85 -4611 -39
rect -4565 -85 -4487 -39
rect -4441 -85 -4363 -39
rect -4317 -85 -4239 -39
rect -4193 -85 -4115 -39
rect -4069 -85 -3991 -39
rect -3945 -85 -3867 -39
rect -3821 -85 -3743 -39
rect -3697 -85 -3619 -39
rect -3573 -85 -3495 -39
rect -3449 -85 -3371 -39
rect -3325 -85 -3247 -39
rect -3201 -85 -3123 -39
rect -3077 -85 -2999 -39
rect -2953 -85 -2875 -39
rect -2829 -85 -2751 -39
rect -2705 -85 -2627 -39
rect -2581 -85 -2503 -39
rect -2457 -85 -2379 -39
rect -2333 -85 -2255 -39
rect -2209 -85 -2131 -39
rect -2085 -85 -2007 -39
rect -1961 -85 -1883 -39
rect -1837 -85 -1759 -39
rect -1713 -85 -1635 -39
rect -1589 -85 -1511 -39
rect -1465 -85 -1387 -39
rect -1341 -85 -1263 -39
rect -1217 -85 -1139 -39
rect -1093 -85 -1015 -39
rect -969 -85 -891 -39
rect -845 -85 -767 -39
rect -721 -85 -643 -39
rect -597 -85 -519 -39
rect -473 -85 -395 -39
rect -349 -85 -271 -39
rect -225 -85 -147 -39
rect -101 -85 -23 -39
rect 23 -85 101 -39
rect 147 -85 225 -39
rect 271 -85 349 -39
rect 395 -85 473 -39
rect 519 -85 597 -39
rect 643 -85 721 -39
rect 767 -85 845 -39
rect 891 -85 969 -39
rect 1015 -85 1093 -39
rect 1139 -85 1217 -39
rect 1263 -85 1341 -39
rect 1387 -85 1465 -39
rect 1511 -85 1589 -39
rect 1635 -85 1713 -39
rect 1759 -85 1837 -39
rect 1883 -85 1961 -39
rect 2007 -85 2085 -39
rect 2131 -85 2209 -39
rect 2255 -85 2333 -39
rect 2379 -85 2457 -39
rect 2503 -85 2581 -39
rect 2627 -85 2705 -39
rect 2751 -85 2829 -39
rect 2875 -85 2953 -39
rect 2999 -85 3077 -39
rect 3123 -85 3201 -39
rect 3247 -85 3325 -39
rect 3371 -85 3449 -39
rect 3495 -85 3573 -39
rect 3619 -85 3697 -39
rect 3743 -85 3821 -39
rect 3867 -85 3945 -39
rect 3991 -85 4069 -39
rect 4115 -85 4193 -39
rect 4239 -85 4317 -39
rect 4363 -85 4441 -39
rect 4487 -85 4565 -39
rect 4611 -85 4689 -39
rect 4735 -85 4813 -39
rect 4859 -85 4937 -39
rect 4983 -85 5061 -39
rect 5107 -85 5185 -39
rect 5231 -85 5309 -39
rect 5355 -85 5433 -39
rect 5479 -85 5557 -39
rect 5603 -85 5681 -39
rect 5727 -85 5805 -39
rect 5851 -85 5929 -39
rect 5975 -85 6053 -39
rect 6099 -85 6177 -39
rect 6223 -85 6301 -39
rect 6347 -85 6425 -39
rect 6471 -85 6549 -39
rect 6595 -85 6673 -39
rect 6719 -85 6797 -39
rect 6843 -85 6921 -39
rect 6967 -85 7045 -39
rect 7091 -85 7169 -39
rect 7215 -85 7226 -39
rect -7226 -96 7226 -85
<< end >>
