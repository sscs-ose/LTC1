magic
tech gf180mcuC
magscale 1 10
timestamp 1699423221
<< nwell >>
rect -2844 -1287 2844 1287
<< nsubdiff >>
rect -2820 1191 2820 1263
rect -2820 -1191 -2748 1191
rect 2748 -1191 2820 1191
rect -2820 -1263 2820 -1191
<< polysilicon >>
rect -2660 1090 -2290 1103
rect -2660 1044 -2647 1090
rect -2303 1044 -2290 1090
rect -2660 1000 -2290 1044
rect -2660 -1044 -2290 -1000
rect -2660 -1090 -2647 -1044
rect -2303 -1090 -2290 -1044
rect -2660 -1103 -2290 -1090
rect -2210 1090 -1840 1103
rect -2210 1044 -2197 1090
rect -1853 1044 -1840 1090
rect -2210 1000 -1840 1044
rect -2210 -1044 -1840 -1000
rect -2210 -1090 -2197 -1044
rect -1853 -1090 -1840 -1044
rect -2210 -1103 -1840 -1090
rect -1760 1090 -1390 1103
rect -1760 1044 -1747 1090
rect -1403 1044 -1390 1090
rect -1760 1000 -1390 1044
rect -1760 -1044 -1390 -1000
rect -1760 -1090 -1747 -1044
rect -1403 -1090 -1390 -1044
rect -1760 -1103 -1390 -1090
rect -1310 1090 -940 1103
rect -1310 1044 -1297 1090
rect -953 1044 -940 1090
rect -1310 1000 -940 1044
rect -1310 -1044 -940 -1000
rect -1310 -1090 -1297 -1044
rect -953 -1090 -940 -1044
rect -1310 -1103 -940 -1090
rect -860 1090 -490 1103
rect -860 1044 -847 1090
rect -503 1044 -490 1090
rect -860 1000 -490 1044
rect -860 -1044 -490 -1000
rect -860 -1090 -847 -1044
rect -503 -1090 -490 -1044
rect -860 -1103 -490 -1090
rect -410 1090 -40 1103
rect -410 1044 -397 1090
rect -53 1044 -40 1090
rect -410 1000 -40 1044
rect -410 -1044 -40 -1000
rect -410 -1090 -397 -1044
rect -53 -1090 -40 -1044
rect -410 -1103 -40 -1090
rect 40 1090 410 1103
rect 40 1044 53 1090
rect 397 1044 410 1090
rect 40 1000 410 1044
rect 40 -1044 410 -1000
rect 40 -1090 53 -1044
rect 397 -1090 410 -1044
rect 40 -1103 410 -1090
rect 490 1090 860 1103
rect 490 1044 503 1090
rect 847 1044 860 1090
rect 490 1000 860 1044
rect 490 -1044 860 -1000
rect 490 -1090 503 -1044
rect 847 -1090 860 -1044
rect 490 -1103 860 -1090
rect 940 1090 1310 1103
rect 940 1044 953 1090
rect 1297 1044 1310 1090
rect 940 1000 1310 1044
rect 940 -1044 1310 -1000
rect 940 -1090 953 -1044
rect 1297 -1090 1310 -1044
rect 940 -1103 1310 -1090
rect 1390 1090 1760 1103
rect 1390 1044 1403 1090
rect 1747 1044 1760 1090
rect 1390 1000 1760 1044
rect 1390 -1044 1760 -1000
rect 1390 -1090 1403 -1044
rect 1747 -1090 1760 -1044
rect 1390 -1103 1760 -1090
rect 1840 1090 2210 1103
rect 1840 1044 1853 1090
rect 2197 1044 2210 1090
rect 1840 1000 2210 1044
rect 1840 -1044 2210 -1000
rect 1840 -1090 1853 -1044
rect 2197 -1090 2210 -1044
rect 1840 -1103 2210 -1090
rect 2290 1090 2660 1103
rect 2290 1044 2303 1090
rect 2647 1044 2660 1090
rect 2290 1000 2660 1044
rect 2290 -1044 2660 -1000
rect 2290 -1090 2303 -1044
rect 2647 -1090 2660 -1044
rect 2290 -1103 2660 -1090
<< polycontact >>
rect -2647 1044 -2303 1090
rect -2647 -1090 -2303 -1044
rect -2197 1044 -1853 1090
rect -2197 -1090 -1853 -1044
rect -1747 1044 -1403 1090
rect -1747 -1090 -1403 -1044
rect -1297 1044 -953 1090
rect -1297 -1090 -953 -1044
rect -847 1044 -503 1090
rect -847 -1090 -503 -1044
rect -397 1044 -53 1090
rect -397 -1090 -53 -1044
rect 53 1044 397 1090
rect 53 -1090 397 -1044
rect 503 1044 847 1090
rect 503 -1090 847 -1044
rect 953 1044 1297 1090
rect 953 -1090 1297 -1044
rect 1403 1044 1747 1090
rect 1403 -1090 1747 -1044
rect 1853 1044 2197 1090
rect 1853 -1090 2197 -1044
rect 2303 1044 2647 1090
rect 2303 -1090 2647 -1044
<< ppolyres >>
rect -2660 -1000 -2290 1000
rect -2210 -1000 -1840 1000
rect -1760 -1000 -1390 1000
rect -1310 -1000 -940 1000
rect -860 -1000 -490 1000
rect -410 -1000 -40 1000
rect 40 -1000 410 1000
rect 490 -1000 860 1000
rect 940 -1000 1310 1000
rect 1390 -1000 1760 1000
rect 1840 -1000 2210 1000
rect 2290 -1000 2660 1000
<< metal1 >>
rect -2658 1044 -2647 1090
rect -2303 1044 -2292 1090
rect -2208 1044 -2197 1090
rect -1853 1044 -1842 1090
rect -1758 1044 -1747 1090
rect -1403 1044 -1392 1090
rect -1308 1044 -1297 1090
rect -953 1044 -942 1090
rect -858 1044 -847 1090
rect -503 1044 -492 1090
rect -408 1044 -397 1090
rect -53 1044 -42 1090
rect 42 1044 53 1090
rect 397 1044 408 1090
rect 492 1044 503 1090
rect 847 1044 858 1090
rect 942 1044 953 1090
rect 1297 1044 1308 1090
rect 1392 1044 1403 1090
rect 1747 1044 1758 1090
rect 1842 1044 1853 1090
rect 2197 1044 2208 1090
rect 2292 1044 2303 1090
rect 2647 1044 2658 1090
rect -2658 -1090 -2647 -1044
rect -2303 -1090 -2292 -1044
rect -2208 -1090 -2197 -1044
rect -1853 -1090 -1842 -1044
rect -1758 -1090 -1747 -1044
rect -1403 -1090 -1392 -1044
rect -1308 -1090 -1297 -1044
rect -953 -1090 -942 -1044
rect -858 -1090 -847 -1044
rect -503 -1090 -492 -1044
rect -408 -1090 -397 -1044
rect -53 -1090 -42 -1044
rect 42 -1090 53 -1044
rect 397 -1090 408 -1044
rect 492 -1090 503 -1044
rect 847 -1090 858 -1044
rect 942 -1090 953 -1044
rect 1297 -1090 1308 -1044
rect 1392 -1090 1403 -1044
rect 1747 -1090 1758 -1044
rect 1842 -1090 1853 -1044
rect 2197 -1090 2208 -1044
rect 2292 -1090 2303 -1044
rect 2647 -1090 2658 -1044
<< properties >>
string FIXED_BBOX -2784 -1227 2784 1227
string gencell ppolyf_u
string library gf180mcu
string parameters w 1.85 l 9.996 m 1 nx 12 wmin 0.80 lmin 1.00 rho 315 val 1.768k dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
