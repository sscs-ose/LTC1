* NGSPICE file created from GF_INV1_flat.ext - technology: gf180mcuC

.subckt GF_INV1_flat VDD IN OUT VSS
X0 OUT IN.t0 VDD.t1 VDD.t0 pfet_03v3 ad=0.165p pd=1.64u as=0.165p ps=1.64u w=0.35u l=0.35u
X1 OUT IN.t1 VSS.t1 VSS.t0 nfet_03v3 ad=0.308p pd=2.28u as=0.308p ps=2.28u w=0.7u l=0.35u
R0 IN.n0 IN.t1 17.2487
R1 IN.n0 IN.t0 12.2493
R2 IN IN.n0 4.18257
R3 VDD.n0 VDD.t0 337.829
R4 VDD.n0 VDD.t1 8.28
R5 VDD VDD.n0 0.0094267
R6 OUT OUT.n0 8.33362
R7 OUT OUT.n1 5.76679
R8 VSS.n56 VSS.n55 348.781
R9 VSS.n6 VSS.n5 261.839
R10 VSS.n59 VSS.t0 245.732
R11 VSS.n43 VSS.n42 235.399
R12 VSS VSS.t1 5.6909
R13 VSS.n4 VSS.n3 2.6005
R14 VSS.n2 VSS.n1 2.6005
R15 VSS.n1 VSS.n0 2.6005
R16 VSS.n36 VSS.n35 2.6005
R17 VSS.n35 VSS.n34 2.6005
R18 VSS.n39 VSS.n38 2.6005
R19 VSS.n38 VSS.n37 2.6005
R20 VSS.n41 VSS.n40 2.6005
R21 VSS.n51 VSS.n50 2.6005
R22 VSS.n50 VSS.n49 2.6005
R23 VSS.n54 VSS.n53 2.6005
R24 VSS.n53 VSS.n52 2.6005
R25 VSS.n58 VSS.n57 2.6005
R26 VSS.n57 VSS.n56 2.6005
R27 VSS.n61 VSS.n60 2.6005
R28 VSS.n60 VSS.n59 2.6005
R29 VSS.n48 VSS.n47 2.6005
R30 VSS.n47 VSS.n46 2.6005
R31 VSS.n63 VSS.n62 2.6005
R32 VSS.n45 VSS.n44 2.6005
R33 VSS.n11 VSS.n10 2.6005
R34 VSS.n10 VSS.n9 2.6005
R35 VSS.n23 VSS.n22 2.6005
R36 VSS.n22 VSS.n21 2.6005
R37 VSS.n20 VSS.n19 2.6005
R38 VSS.n19 VSS.n18 2.6005
R39 VSS.n17 VSS.n16 2.6005
R40 VSS.n16 VSS.n15 2.6005
R41 VSS.n14 VSS.n13 2.6005
R42 VSS.n13 VSS.n12 2.6005
R43 VSS.n26 VSS.n25 2.6005
R44 VSS.n8 VSS.n7 2.6005
R45 VSS.n28 VSS.n27 2.6005
R46 VSS.n31 VSS.n30 2.6005
R47 VSS.n33 VSS.n32 2.6005
R48 VSS.n70 VSS.n69 2.6005
R49 VSS.n66 VSS.n65 2.6005
R50 VSS.n69 VSS.n68 1.77751
R51 VSS.n65 VSS.n64 1.55416
R52 VSS.n7 VSS.n6 1.53965
R53 VSS.n30 VSS.n29 1.53464
R54 VSS.n25 VSS.n24 1.18756
R55 VSS.n68 VSS.n67 0.412744
R56 VSS.n44 VSS.n43 0.387192
R57 VSS.n11 VSS.n8 0.159389
R58 VSS.n63 VSS.n61 0.155256
R59 VSS.n14 VSS.n11 0.1505
R60 VSS.n17 VSS.n14 0.1505
R61 VSS.n20 VSS.n17 0.1505
R62 VSS.n23 VSS.n20 0.1505
R63 VSS.n26 VSS.n23 0.1505
R64 VSS.n48 VSS.n45 0.148671
R65 VSS.n51 VSS.n48 0.148671
R66 VSS.n54 VSS.n51 0.148671
R67 VSS.n58 VSS.n54 0.148671
R68 VSS.n61 VSS.n58 0.148671
R69 VSS.n4 VSS.n2 0.144731
R70 VSS.n39 VSS.n36 0.144731
R71 VSS.n41 VSS.n39 0.144731
R72 VSS.n31 VSS.n28 0.144731
R73 VSS.n33 VSS.n31 0.144731
R74 VSS.n70 VSS.n66 0.144731
R75 VSS VSS.n71 0.117309
R76 VSS.n71 VSS.n33 0.112423
R77 VSS.n66 VSS.n63 0.0996745
R78 VSS.n8 VSS.n4 0.0974231
R79 VSS.n45 VSS.n41 0.0869259
R80 VSS.n28 VSS.n26 0.084688
R81 VSS.n71 VSS.n70 0.0328077
C0 VDD IN 0.217f
C1 VDD OUT 0.0775f
C2 OUT IN 0.0708f
.ends

