magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -2241 -1019 2241 1019
<< metal1 >>
rect -1241 13 1241 19
rect -1241 -13 -1235 13
rect 1235 -13 1241 13
rect -1241 -19 1241 -13
<< via1 >>
rect -1235 -13 1235 13
<< metal2 >>
rect -1241 13 1241 19
rect -1241 -13 -1235 13
rect 1235 -13 1241 13
rect -1241 -19 1241 -13
<< end >>
