magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1484 -1174 1484 1174
<< metal1 >>
rect -484 168 484 174
rect -484 142 -478 168
rect -452 142 -416 168
rect -390 142 -354 168
rect -328 142 -292 168
rect -266 142 -230 168
rect -204 142 -168 168
rect -142 142 -106 168
rect -80 142 -44 168
rect -18 142 18 168
rect 44 142 80 168
rect 106 142 142 168
rect 168 142 204 168
rect 230 142 266 168
rect 292 142 328 168
rect 354 142 390 168
rect 416 142 452 168
rect 478 142 484 168
rect -484 106 484 142
rect -484 80 -478 106
rect -452 80 -416 106
rect -390 80 -354 106
rect -328 80 -292 106
rect -266 80 -230 106
rect -204 80 -168 106
rect -142 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 142 106
rect 168 80 204 106
rect 230 80 266 106
rect 292 80 328 106
rect 354 80 390 106
rect 416 80 452 106
rect 478 80 484 106
rect -484 44 484 80
rect -484 18 -478 44
rect -452 18 -416 44
rect -390 18 -354 44
rect -328 18 -292 44
rect -266 18 -230 44
rect -204 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 204 44
rect 230 18 266 44
rect 292 18 328 44
rect 354 18 390 44
rect 416 18 452 44
rect 478 18 484 44
rect -484 -18 484 18
rect -484 -44 -478 -18
rect -452 -44 -416 -18
rect -390 -44 -354 -18
rect -328 -44 -292 -18
rect -266 -44 -230 -18
rect -204 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 204 -18
rect 230 -44 266 -18
rect 292 -44 328 -18
rect 354 -44 390 -18
rect 416 -44 452 -18
rect 478 -44 484 -18
rect -484 -80 484 -44
rect -484 -106 -478 -80
rect -452 -106 -416 -80
rect -390 -106 -354 -80
rect -328 -106 -292 -80
rect -266 -106 -230 -80
rect -204 -106 -168 -80
rect -142 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 142 -80
rect 168 -106 204 -80
rect 230 -106 266 -80
rect 292 -106 328 -80
rect 354 -106 390 -80
rect 416 -106 452 -80
rect 478 -106 484 -80
rect -484 -142 484 -106
rect -484 -168 -478 -142
rect -452 -168 -416 -142
rect -390 -168 -354 -142
rect -328 -168 -292 -142
rect -266 -168 -230 -142
rect -204 -168 -168 -142
rect -142 -168 -106 -142
rect -80 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 80 -142
rect 106 -168 142 -142
rect 168 -168 204 -142
rect 230 -168 266 -142
rect 292 -168 328 -142
rect 354 -168 390 -142
rect 416 -168 452 -142
rect 478 -168 484 -142
rect -484 -174 484 -168
<< via1 >>
rect -478 142 -452 168
rect -416 142 -390 168
rect -354 142 -328 168
rect -292 142 -266 168
rect -230 142 -204 168
rect -168 142 -142 168
rect -106 142 -80 168
rect -44 142 -18 168
rect 18 142 44 168
rect 80 142 106 168
rect 142 142 168 168
rect 204 142 230 168
rect 266 142 292 168
rect 328 142 354 168
rect 390 142 416 168
rect 452 142 478 168
rect -478 80 -452 106
rect -416 80 -390 106
rect -354 80 -328 106
rect -292 80 -266 106
rect -230 80 -204 106
rect -168 80 -142 106
rect -106 80 -80 106
rect -44 80 -18 106
rect 18 80 44 106
rect 80 80 106 106
rect 142 80 168 106
rect 204 80 230 106
rect 266 80 292 106
rect 328 80 354 106
rect 390 80 416 106
rect 452 80 478 106
rect -478 18 -452 44
rect -416 18 -390 44
rect -354 18 -328 44
rect -292 18 -266 44
rect -230 18 -204 44
rect -168 18 -142 44
rect -106 18 -80 44
rect -44 18 -18 44
rect 18 18 44 44
rect 80 18 106 44
rect 142 18 168 44
rect 204 18 230 44
rect 266 18 292 44
rect 328 18 354 44
rect 390 18 416 44
rect 452 18 478 44
rect -478 -44 -452 -18
rect -416 -44 -390 -18
rect -354 -44 -328 -18
rect -292 -44 -266 -18
rect -230 -44 -204 -18
rect -168 -44 -142 -18
rect -106 -44 -80 -18
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect 80 -44 106 -18
rect 142 -44 168 -18
rect 204 -44 230 -18
rect 266 -44 292 -18
rect 328 -44 354 -18
rect 390 -44 416 -18
rect 452 -44 478 -18
rect -478 -106 -452 -80
rect -416 -106 -390 -80
rect -354 -106 -328 -80
rect -292 -106 -266 -80
rect -230 -106 -204 -80
rect -168 -106 -142 -80
rect -106 -106 -80 -80
rect -44 -106 -18 -80
rect 18 -106 44 -80
rect 80 -106 106 -80
rect 142 -106 168 -80
rect 204 -106 230 -80
rect 266 -106 292 -80
rect 328 -106 354 -80
rect 390 -106 416 -80
rect 452 -106 478 -80
rect -478 -168 -452 -142
rect -416 -168 -390 -142
rect -354 -168 -328 -142
rect -292 -168 -266 -142
rect -230 -168 -204 -142
rect -168 -168 -142 -142
rect -106 -168 -80 -142
rect -44 -168 -18 -142
rect 18 -168 44 -142
rect 80 -168 106 -142
rect 142 -168 168 -142
rect 204 -168 230 -142
rect 266 -168 292 -142
rect 328 -168 354 -142
rect 390 -168 416 -142
rect 452 -168 478 -142
<< metal2 >>
rect -484 168 484 174
rect -484 142 -478 168
rect -452 142 -416 168
rect -390 142 -354 168
rect -328 142 -292 168
rect -266 142 -230 168
rect -204 142 -168 168
rect -142 142 -106 168
rect -80 142 -44 168
rect -18 142 18 168
rect 44 142 80 168
rect 106 142 142 168
rect 168 142 204 168
rect 230 142 266 168
rect 292 142 328 168
rect 354 142 390 168
rect 416 142 452 168
rect 478 142 484 168
rect -484 106 484 142
rect -484 80 -478 106
rect -452 80 -416 106
rect -390 80 -354 106
rect -328 80 -292 106
rect -266 80 -230 106
rect -204 80 -168 106
rect -142 80 -106 106
rect -80 80 -44 106
rect -18 80 18 106
rect 44 80 80 106
rect 106 80 142 106
rect 168 80 204 106
rect 230 80 266 106
rect 292 80 328 106
rect 354 80 390 106
rect 416 80 452 106
rect 478 80 484 106
rect -484 44 484 80
rect -484 18 -478 44
rect -452 18 -416 44
rect -390 18 -354 44
rect -328 18 -292 44
rect -266 18 -230 44
rect -204 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 204 44
rect 230 18 266 44
rect 292 18 328 44
rect 354 18 390 44
rect 416 18 452 44
rect 478 18 484 44
rect -484 -18 484 18
rect -484 -44 -478 -18
rect -452 -44 -416 -18
rect -390 -44 -354 -18
rect -328 -44 -292 -18
rect -266 -44 -230 -18
rect -204 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 204 -18
rect 230 -44 266 -18
rect 292 -44 328 -18
rect 354 -44 390 -18
rect 416 -44 452 -18
rect 478 -44 484 -18
rect -484 -80 484 -44
rect -484 -106 -478 -80
rect -452 -106 -416 -80
rect -390 -106 -354 -80
rect -328 -106 -292 -80
rect -266 -106 -230 -80
rect -204 -106 -168 -80
rect -142 -106 -106 -80
rect -80 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 80 -80
rect 106 -106 142 -80
rect 168 -106 204 -80
rect 230 -106 266 -80
rect 292 -106 328 -80
rect 354 -106 390 -80
rect 416 -106 452 -80
rect 478 -106 484 -80
rect -484 -142 484 -106
rect -484 -168 -478 -142
rect -452 -168 -416 -142
rect -390 -168 -354 -142
rect -328 -168 -292 -142
rect -266 -168 -230 -142
rect -204 -168 -168 -142
rect -142 -168 -106 -142
rect -80 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 80 -142
rect 106 -168 142 -142
rect 168 -168 204 -142
rect 230 -168 266 -142
rect 292 -168 328 -142
rect 354 -168 390 -142
rect 416 -168 452 -142
rect 478 -168 484 -142
rect -484 -174 484 -168
<< end >>
