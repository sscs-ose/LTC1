magic
tech gf180mcuC
magscale 1 10
timestamp 1714558796
<< nwell >>
rect -127 -1195 709 -667
rect 580 -2292 1412 -1764
rect -140 -3533 670 -3005
rect 2752 -3533 3687 -3005
rect 331 -4630 1216 -4102
rect 3578 -4630 4405 -4102
rect 1 -5855 856 -5327
rect 3262 -5854 4444 -5326
rect 975 -6578 1130 -6424
rect 3966 -6951 4761 -6423
<< metal1 >>
rect 1635 742 3048 768
rect 1635 690 2959 742
rect 3011 690 3048 742
rect 1635 622 3048 690
rect 7760 732 8311 756
rect 7760 680 8227 732
rect 8280 680 8311 732
rect 7760 645 8311 680
rect 1635 588 2590 622
rect -638 191 745 217
rect 2597 196 2801 210
rect -638 119 1710 191
rect 2597 180 2730 196
rect 2522 134 2730 180
rect 2791 134 2801 196
rect 2522 122 2801 134
rect -638 113 745 119
rect -638 -1158 -534 113
rect 2650 -144 3238 -31
rect 7750 -51 10195 -20
rect 7750 -105 10105 -51
rect 10160 -105 10195 -51
rect 7750 -141 10195 -105
rect 2650 -153 2763 -144
rect 1685 -327 2763 -153
rect 7566 -212 9450 -196
rect 7566 -264 9383 -212
rect 9436 -264 9450 -212
rect 7566 -274 9450 -264
rect 7566 -275 9446 -274
rect -439 -352 2763 -327
rect -439 -405 -415 -352
rect -362 -398 2763 -352
rect 6437 -368 6555 -366
rect 6437 -391 7349 -368
rect -362 -405 2746 -398
rect -439 -417 2746 -405
rect -439 -433 2634 -417
rect 2931 -445 4467 -422
rect 2931 -497 2959 -445
rect 3011 -449 4467 -445
rect 3011 -497 4385 -449
rect 2931 -501 4385 -497
rect 4437 -501 4467 -449
rect 6437 -446 6475 -391
rect 6530 -409 7349 -391
rect 6530 -446 7261 -409
rect 6437 -461 7261 -446
rect 7315 -461 7349 -409
rect 6437 -484 7349 -461
rect 6591 -485 7349 -484
rect 2931 -522 4467 -501
rect 5479 -561 7779 -542
rect 5479 -598 7707 -561
rect 3183 -614 7707 -598
rect 7760 -614 7779 -561
rect 3183 -620 7779 -614
rect 54 -832 414 -654
rect 3183 -673 3199 -620
rect 3252 -632 7779 -620
rect 3252 -673 5569 -632
rect 3183 -688 5569 -673
rect 2706 -944 5389 -918
rect 2706 -996 5311 -944
rect 5364 -996 5389 -944
rect 2706 -1018 5389 -996
rect -638 -1262 -218 -1158
rect -638 -3479 -534 -1262
rect 845 -1271 951 -1216
rect 2780 -1295 6822 -1212
rect 7859 -1231 7943 -1219
rect 2780 -1398 2965 -1295
rect 7603 -1297 7694 -1236
rect 7859 -1287 7874 -1231
rect 7931 -1287 7943 -1231
rect 9955 -1282 10327 -1234
rect 7603 -1324 7652 -1297
rect 7859 -1300 7943 -1287
rect 9939 -1680 10195 -1662
rect 9939 -1734 10109 -1680
rect 10164 -1734 10195 -1680
rect 9939 -1761 10195 -1734
rect 728 -1919 1033 -1764
rect 5188 -1984 6380 -1947
rect 5188 -2036 6295 -1984
rect 6348 -2036 6380 -1984
rect 5188 -2064 6380 -2036
rect 7556 -2285 7642 -2284
rect 838 -2368 945 -2313
rect 1549 -2368 1669 -2313
rect 7556 -2342 7569 -2285
rect 7626 -2342 7642 -2285
rect 8673 -2342 8685 -2284
rect 8743 -2342 8839 -2284
rect 5568 -2555 5665 -2554
rect 5451 -2570 5665 -2555
rect 5451 -2623 5592 -2570
rect 5644 -2623 5665 -2570
rect 5451 -2631 5665 -2623
rect 5568 -2641 5665 -2631
rect -439 -2769 53 -2744
rect -439 -2821 -412 -2769
rect -360 -2821 53 -2769
rect -439 -2850 53 -2821
rect 142 -3064 263 -3004
rect 84 -3170 263 -3064
rect 3101 -3114 3203 -3064
rect 3101 -3121 3270 -3114
rect 3146 -3171 3270 -3121
rect -638 -3583 -199 -3479
rect -638 -5834 -534 -3583
rect 820 -3609 914 -3554
rect 3824 -3609 3933 -3554
rect -338 -3764 -233 -3763
rect -439 -3792 -232 -3764
rect -439 -3844 -415 -3792
rect -363 -3844 -232 -3792
rect -439 -3870 -232 -3844
rect 855 -4111 1006 -4102
rect 743 -4257 1006 -4111
rect 3721 -4257 3986 -4102
rect 807 -4706 921 -4651
rect 1504 -4676 1635 -4625
rect 1525 -4706 1635 -4676
rect 3835 -4706 3938 -4651
rect 4548 -4706 4662 -4651
rect 76 -5153 5788 -5044
rect 153 -5492 536 -5291
rect 3110 -5318 6050 -5291
rect 3110 -5338 6555 -5318
rect 3110 -5390 6447 -5338
rect 6499 -5390 6555 -5338
rect 3110 -5436 6555 -5390
rect 3110 -5491 6050 -5436
rect -638 -5938 -221 -5834
rect 933 -5931 1038 -5876
rect 4171 -5930 4285 -5875
rect 6276 -5980 9197 -5929
rect 6276 -6032 9101 -5980
rect 9158 -6032 9197 -5980
rect 6276 -6066 9197 -6032
rect -165 -6083 -16 -6081
rect -439 -6113 -16 -6083
rect -439 -6166 -422 -6113
rect -368 -6166 -16 -6113
rect -439 -6189 -16 -6166
rect 975 -6578 1130 -6424
rect 4077 -6578 4464 -6423
rect 983 -6579 1028 -6578
rect -196 -6790 17 -6787
rect -200 -6870 20 -6790
rect -200 -6930 -190 -6870
rect -130 -6930 20 -6870
rect -200 -6970 20 -6930
rect -196 -7090 11 -6970
rect 933 -7028 1049 -6973
rect 1633 -7028 1770 -6973
rect 4183 -7027 4294 -6972
rect 4905 -7027 5018 -6972
<< via1 >>
rect 2959 690 3011 742
rect 8227 680 8280 732
rect 2730 134 2791 196
rect 10105 -105 10160 -51
rect 9383 -264 9436 -212
rect -415 -405 -362 -352
rect 2959 -497 3011 -445
rect 4385 -501 4437 -449
rect 6475 -446 6530 -391
rect 7261 -461 7315 -409
rect 7707 -614 7760 -561
rect 3199 -673 3252 -620
rect 8228 -767 8281 -715
rect 5311 -996 5364 -944
rect 7874 -1287 7931 -1231
rect 10109 -1734 10164 -1680
rect 6295 -2036 6348 -1984
rect 7569 -2342 7626 -2285
rect 8685 -2342 8743 -2284
rect 5592 -2623 5644 -2570
rect -412 -2821 -360 -2769
rect -415 -3844 -363 -3792
rect 6447 -5390 6499 -5338
rect 9101 -6032 9158 -5980
rect -422 -6166 -368 -6113
rect -190 -6930 -130 -6870
<< metal2 >>
rect 2931 742 3045 768
rect 2931 690 2959 742
rect 3011 690 3045 742
rect 2597 196 2801 210
rect 2597 134 2730 196
rect 2791 134 2801 196
rect 2597 122 2801 134
rect -439 -352 -333 -327
rect -439 -405 -415 -352
rect -362 -405 -333 -352
rect -439 -2769 -333 -405
rect 2931 -445 3045 690
rect 8200 732 8311 756
rect 8200 680 8227 732
rect 8280 680 8311 732
rect 2931 -497 2959 -445
rect 3011 -497 3045 -445
rect 2931 -522 3045 -497
rect 3183 -620 3273 -199
rect 4349 -449 4466 -196
rect 4349 -501 4385 -449
rect 4437 -501 4466 -449
rect 4349 -522 4466 -501
rect 3183 -673 3199 -620
rect 3252 -673 3273 -620
rect 3183 -688 3273 -673
rect 5283 -944 5400 -189
rect 5283 -996 5311 -944
rect 5364 -996 5400 -944
rect 5283 -1020 5400 -996
rect 6263 -1984 6380 -193
rect 6263 -2036 6295 -1984
rect 6348 -2036 6380 -1984
rect 6263 -2064 6380 -2036
rect 6438 -391 6555 -367
rect 6438 -446 6475 -391
rect 6530 -446 6555 -391
rect 5534 -2554 5664 -2553
rect 5534 -2567 5665 -2554
rect 5534 -2623 5588 -2567
rect 5644 -2623 5665 -2567
rect 5534 -2631 5665 -2623
rect 5568 -2641 5665 -2631
rect -439 -2821 -412 -2769
rect -360 -2821 -333 -2769
rect -439 -3792 -333 -2821
rect -439 -3844 -415 -3792
rect -363 -3844 -333 -3792
rect -439 -6113 -333 -3844
rect 6438 -5338 6555 -446
rect 7232 -409 7349 -193
rect 7232 -461 7261 -409
rect 7315 -461 7349 -409
rect 7232 -484 7349 -461
rect 7689 -561 7779 -542
rect 7689 -614 7707 -561
rect 7760 -614 7779 -561
rect 7689 -893 7779 -614
rect 8200 -715 8311 680
rect 10074 -51 10195 -20
rect 10074 -105 10105 -51
rect 10160 -105 10195 -51
rect 8200 -767 8228 -715
rect 8281 -767 8311 -715
rect 8200 -798 8311 -767
rect 9371 -212 9450 -196
rect 9371 -264 9383 -212
rect 9436 -264 9450 -212
rect 9371 -274 9450 -264
rect 7003 -952 7779 -893
rect 7005 -1129 7063 -952
rect 9371 -996 9446 -274
rect 9371 -1127 9462 -996
rect 9247 -1185 9462 -1127
rect 9247 -1186 9430 -1185
rect 7859 -1231 7943 -1219
rect 7859 -1287 7874 -1231
rect 7931 -1287 7943 -1231
rect 7859 -1300 7943 -1287
rect 10074 -1680 10195 -105
rect 10074 -1734 10109 -1680
rect 10164 -1734 10195 -1680
rect 10074 -1758 10195 -1734
rect 7556 -2285 7639 -2273
rect 7556 -2342 7569 -2285
rect 7626 -2342 7639 -2285
rect 7556 -2355 7639 -2342
rect 8672 -2284 8767 -2271
rect 8672 -2342 8685 -2284
rect 8743 -2342 8767 -2284
rect 8672 -2355 8767 -2342
rect 6438 -5390 6447 -5338
rect 6499 -5390 6555 -5338
rect 6438 -5436 6555 -5390
rect 9060 -2955 9197 -2940
rect 9060 -3011 9090 -2955
rect 9146 -3011 9197 -2955
rect 9060 -5980 9197 -3011
rect 9060 -6032 9101 -5980
rect 9158 -6032 9197 -5980
rect 9060 -6066 9197 -6032
rect -439 -6166 -422 -6113
rect -368 -6166 -333 -6113
rect -439 -6189 -333 -6166
rect -196 -6790 17 -6787
rect -200 -6870 20 -6790
rect -200 -6930 -190 -6870
rect -130 -6930 20 -6870
rect -200 -6970 20 -6930
<< via2 >>
rect 2731 135 2787 193
rect 5588 -2570 5644 -2567
rect 5588 -2623 5592 -2570
rect 5592 -2623 5644 -2570
rect 1219 -4603 1275 -4547
rect 7874 -1287 7931 -1231
rect 7569 -2342 7626 -2285
rect 8685 -2342 8743 -2284
rect 9090 -3011 9146 -2955
rect -190 -6930 -130 -6870
<< metal3 >>
rect 2719 203 2801 210
rect 2719 193 3118 203
rect 2719 135 2731 193
rect 2787 135 3118 193
rect 2719 123 3118 135
rect 2720 122 3118 123
rect -193 -4534 -111 -2207
rect 3037 -2272 3118 122
rect 7859 -1231 9156 -1219
rect 7859 -1287 7874 -1231
rect 7931 -1287 9156 -1231
rect 7859 -1300 9156 -1287
rect 7507 -2272 7602 -2271
rect 3037 -2273 7602 -2272
rect 3037 -2285 7639 -2273
rect 3037 -2342 7569 -2285
rect 7626 -2342 7639 -2285
rect 3037 -2353 7639 -2342
rect 7507 -2354 7639 -2353
rect 7556 -2355 7639 -2354
rect 8654 -2284 8789 -2272
rect 8654 -2342 8685 -2284
rect 8743 -2342 8789 -2284
rect 8654 -2359 8789 -2342
rect 8654 -2553 8741 -2359
rect 5558 -2567 8741 -2553
rect 5558 -2623 5588 -2567
rect 5644 -2623 8741 -2567
rect 5558 -2640 8741 -2623
rect 9075 -2955 9156 -1300
rect 9075 -3011 9090 -2955
rect 9146 -3011 9156 -2955
rect 9075 -3023 9156 -3011
rect -193 -4547 1292 -4534
rect -193 -4603 1219 -4547
rect 1275 -4603 1292 -4547
rect -193 -4615 1292 -4603
rect -193 -4616 1271 -4615
rect -193 -6787 -111 -4616
rect -196 -6790 17 -6787
rect -200 -6850 20 -6790
rect -200 -6870 92 -6850
rect -200 -6930 -190 -6870
rect -130 -6930 92 -6870
rect -200 -6932 92 -6930
rect -200 -6970 20 -6932
use Buffer_delayed_mag  Buffer_delayed_mag_0
timestamp 1714534647
transform 1 0 1756 0 1 -9
box -218 -175 878 669
use CLK_div_2_mag  CLK_div_2_mag_0
timestamp 1714558667
transform 1 0 -169 0 1 -2895
box -206 12 3133 2241
use CLK_div_3_mag  CLK_div_3_mag_0
timestamp 1714558796
transform 1 0 -263 0 1 -5153
box -40 -1 6461 3249
use CLK_div_4_mag  CLK_div_4_mag_0
timestamp 1714558667
transform 1 0 -274 0 1 -7543
box -44 -35 6589 2252
use dec_2x4_ibr_mag  dec_2x4_ibr_mag_0
timestamp 1714558529
transform 1 0 3556 0 1 -285
box -396 -5 4275 1071
use mux_4x1  mux_4x1_0
timestamp 1714480907
transform 1 0 7809 0 1 -2792
box -1194 5 2229 2107
<< labels >>
flabel metal1 4085 -626 4085 -626 0 FreeSans 1600 0 0 0 OPA0
port 0 nsew
flabel metal1 8502 -237 8502 -237 0 FreeSans 1600 0 0 0 OPA1
port 1 nsew
flabel metal1 10312 -1261 10312 -1261 0 FreeSans 1600 0 0 0 Vdiv
port 2 nsew
flabel metal1 7951 711 7951 711 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel metal1 7924 -95 7924 -95 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal1 -584 174 -584 174 0 FreeSans 1600 0 0 0 CLK
port 5 nsew
flabel metal1 -108 -7055 -108 -7055 0 FreeSans 1600 0 0 0 RST
port 6 nsew
<< end >>
