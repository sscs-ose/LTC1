magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1073 -1316 1073 1316
<< metal1 >>
rect -73 310 73 316
rect -73 284 -67 310
rect -41 284 -13 310
rect 13 284 41 310
rect 67 284 73 310
rect -73 256 73 284
rect -73 230 -67 256
rect -41 230 -13 256
rect 13 230 41 256
rect 67 230 73 256
rect -73 202 73 230
rect -73 176 -67 202
rect -41 176 -13 202
rect 13 176 41 202
rect 67 176 73 202
rect -73 148 73 176
rect -73 122 -67 148
rect -41 122 -13 148
rect 13 122 41 148
rect 67 122 73 148
rect -73 94 73 122
rect -73 68 -67 94
rect -41 68 -13 94
rect 13 68 41 94
rect 67 68 73 94
rect -73 40 73 68
rect -73 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 73 40
rect -73 -14 73 14
rect -73 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 73 -14
rect -73 -68 73 -40
rect -73 -94 -67 -68
rect -41 -94 -13 -68
rect 13 -94 41 -68
rect 67 -94 73 -68
rect -73 -122 73 -94
rect -73 -148 -67 -122
rect -41 -148 -13 -122
rect 13 -148 41 -122
rect 67 -148 73 -122
rect -73 -176 73 -148
rect -73 -202 -67 -176
rect -41 -202 -13 -176
rect 13 -202 41 -176
rect 67 -202 73 -176
rect -73 -230 73 -202
rect -73 -256 -67 -230
rect -41 -256 -13 -230
rect 13 -256 41 -230
rect 67 -256 73 -230
rect -73 -284 73 -256
rect -73 -310 -67 -284
rect -41 -310 -13 -284
rect 13 -310 41 -284
rect 67 -310 73 -284
rect -73 -316 73 -310
<< via1 >>
rect -67 284 -41 310
rect -13 284 13 310
rect 41 284 67 310
rect -67 230 -41 256
rect -13 230 13 256
rect 41 230 67 256
rect -67 176 -41 202
rect -13 176 13 202
rect 41 176 67 202
rect -67 122 -41 148
rect -13 122 13 148
rect 41 122 67 148
rect -67 68 -41 94
rect -13 68 13 94
rect 41 68 67 94
rect -67 14 -41 40
rect -13 14 13 40
rect 41 14 67 40
rect -67 -40 -41 -14
rect -13 -40 13 -14
rect 41 -40 67 -14
rect -67 -94 -41 -68
rect -13 -94 13 -68
rect 41 -94 67 -68
rect -67 -148 -41 -122
rect -13 -148 13 -122
rect 41 -148 67 -122
rect -67 -202 -41 -176
rect -13 -202 13 -176
rect 41 -202 67 -176
rect -67 -256 -41 -230
rect -13 -256 13 -230
rect 41 -256 67 -230
rect -67 -310 -41 -284
rect -13 -310 13 -284
rect 41 -310 67 -284
<< metal2 >>
rect -73 310 73 316
rect -73 284 -67 310
rect -41 284 -13 310
rect 13 284 41 310
rect 67 284 73 310
rect -73 256 73 284
rect -73 230 -67 256
rect -41 230 -13 256
rect 13 230 41 256
rect 67 230 73 256
rect -73 202 73 230
rect -73 176 -67 202
rect -41 176 -13 202
rect 13 176 41 202
rect 67 176 73 202
rect -73 148 73 176
rect -73 122 -67 148
rect -41 122 -13 148
rect 13 122 41 148
rect 67 122 73 148
rect -73 94 73 122
rect -73 68 -67 94
rect -41 68 -13 94
rect 13 68 41 94
rect 67 68 73 94
rect -73 40 73 68
rect -73 14 -67 40
rect -41 14 -13 40
rect 13 14 41 40
rect 67 14 73 40
rect -73 -14 73 14
rect -73 -40 -67 -14
rect -41 -40 -13 -14
rect 13 -40 41 -14
rect 67 -40 73 -14
rect -73 -68 73 -40
rect -73 -94 -67 -68
rect -41 -94 -13 -68
rect 13 -94 41 -68
rect 67 -94 73 -68
rect -73 -122 73 -94
rect -73 -148 -67 -122
rect -41 -148 -13 -122
rect 13 -148 41 -122
rect 67 -148 73 -122
rect -73 -176 73 -148
rect -73 -202 -67 -176
rect -41 -202 -13 -176
rect 13 -202 41 -176
rect 67 -202 73 -176
rect -73 -230 73 -202
rect -73 -256 -67 -230
rect -41 -256 -13 -230
rect 13 -256 41 -230
rect 67 -256 73 -230
rect -73 -284 73 -256
rect -73 -310 -67 -284
rect -41 -310 -13 -284
rect 13 -310 41 -284
rect 67 -310 73 -284
rect -73 -316 73 -310
<< end >>
