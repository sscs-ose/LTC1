magic
tech gf180mcuC
magscale 1 10
timestamp 1693459011
<< nwell >>
rect -744 -386 744 386
<< nsubdiff >>
rect -720 290 720 362
rect -720 -290 -648 290
rect 648 -290 720 290
rect -720 -362 720 -290
<< polysilicon >>
rect -560 189 -400 202
rect -560 143 -547 189
rect -413 143 -400 189
rect -560 100 -400 143
rect -560 -143 -400 -100
rect -560 -189 -547 -143
rect -413 -189 -400 -143
rect -560 -202 -400 -189
rect -320 189 -160 202
rect -320 143 -307 189
rect -173 143 -160 189
rect -320 100 -160 143
rect -320 -143 -160 -100
rect -320 -189 -307 -143
rect -173 -189 -160 -143
rect -320 -202 -160 -189
rect -80 189 80 202
rect -80 143 -67 189
rect 67 143 80 189
rect -80 100 80 143
rect -80 -143 80 -100
rect -80 -189 -67 -143
rect 67 -189 80 -143
rect -80 -202 80 -189
rect 160 189 320 202
rect 160 143 173 189
rect 307 143 320 189
rect 160 100 320 143
rect 160 -143 320 -100
rect 160 -189 173 -143
rect 307 -189 320 -143
rect 160 -202 320 -189
rect 400 189 560 202
rect 400 143 413 189
rect 547 143 560 189
rect 400 100 560 143
rect 400 -143 560 -100
rect 400 -189 413 -143
rect 547 -189 560 -143
rect 400 -202 560 -189
<< polycontact >>
rect -547 143 -413 189
rect -547 -189 -413 -143
rect -307 143 -173 189
rect -307 -189 -173 -143
rect -67 143 67 189
rect -67 -189 67 -143
rect 173 143 307 189
rect 173 -189 307 -143
rect 413 143 547 189
rect 413 -189 547 -143
<< ppolyres >>
rect -560 -100 -400 100
rect -320 -100 -160 100
rect -80 -100 80 100
rect 160 -100 320 100
rect 400 -100 560 100
<< metal1 >>
rect -558 143 -547 189
rect -413 143 -402 189
rect -318 143 -307 189
rect -173 143 -162 189
rect -78 143 -67 189
rect 67 143 78 189
rect 162 143 173 189
rect 307 143 318 189
rect 402 143 413 189
rect 547 143 558 189
rect -558 -189 -547 -143
rect -413 -189 -402 -143
rect -318 -189 -307 -143
rect -173 -189 -162 -143
rect -78 -189 -67 -143
rect 67 -189 78 -143
rect 162 -189 173 -143
rect 307 -189 318 -143
rect 402 -189 413 -143
rect 547 -189 558 -143
<< properties >>
string FIXED_BBOX -684 -326 684 326
string gencell ppolyf_u
string library gf180mcu
string parameters w 0.8 l 1.0 m 1 nx 5 wmin 0.80 lmin 1.00 rho 315 val 431.506 dummy 0 dw 0.07 term 0.0 sterm 0.0 caplen 0.4 snake 0 glc 0 grc 0 gtc 0 gbc 0 roverlap 0 endcov 100 full_metal 0
<< end >>
