* NGSPICE file created from nmos_3p3_GGGST2_flat_flat.ext - technology: gf180mcuC

.subckt nmos_3p3_GGGST2_flat_flat A B OUT VDD VSS
X0 VDD B.t1 a_168_68.t0 VDD.t0 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 VSS B.t2 a_24_68.t0 VSS.t0 nfet_03v3 ad=0.13p pd=1.02u as=0.13p ps=1.02u w=0.5u l=0.28u
X2 OUT a_168_68.t4 VDD.t4 VDD.t3 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X3 OUT a_168_68.t5 VSS.t6 VSS.t5 nfet_03v3 ad=0.22p pd=1.88u as=0.22p ps=1.88u w=0.5u l=0.28u
R0 A.n0 A.t2 33.763
R1 A.n1 A.n0 17.2076
R2 A.n1 A.t1 15.8587
R3 A.n0 A.t0 13.9487
R4 A A.n1 4.06507
R5 a_168_68.n0 a_168_68.t5 65.7005
R6 a_168_68.n0 a_168_68.t4 18.6271
R7 a_168_68.n3 a_168_68.n0 4.45833
R8 a_168_68.n3 a_168_68.n2 3.9018
R9 a_168_68.n2 a_168_68.t3 3.2765
R10 a_168_68.n2 a_168_68.n1 3.2765
R11 a_168_68.n5 a_168_68.n3 2.89789
R12 a_168_68.t0 a_168_68.n5 1.8205
R13 a_168_68.n5 a_168_68.n4 1.8205
R14 a_24_68.n3 a_24_68.n0 7.42041
R15 a_24_68.t2 a_24_68.n3 7.42041
R16 a_24_68.n2 a_24_68.t0 3.2765
R17 a_24_68.n2 a_24_68.n1 3.2765
R18 a_24_68.n3 a_24_68.n2 3.1505
R19 VSS.t0 VSS.n26 389.159
R20 VSS.n23 VSS.t8 241.91
R21 VSS.n27 VSS.t0 105.178
R22 VSS.n17 VSS.t7 94.6607
R23 VSS.n3 VSS.t5 42.0717
R24 VSS.n14 VSS.t3 42.0717
R25 VSS.n16 VSS.n15 9.13939
R26 VSS.n28 VSS.n16 9.13939
R27 VSS.n6 VSS.t6 7.04085
R28 VSS VSS.n16 5.2005
R29 VSS VSS.n16 5.2005
R30 VSS.n2 VSS.n1 3.76485
R31 VSS.n1 VSS.t4 3.2765
R32 VSS.n1 VSS.n0 3.2765
R33 VSS.n4 VSS.n3 2.6005
R34 VSS.n9 VSS.n8 2.6005
R35 VSS.n8 VSS.n7 2.6005
R36 VSS.n12 VSS.n11 2.6005
R37 VSS.n11 VSS.n10 2.6005
R38 VSS.n15 VSS.n13 2.6005
R39 VSS.n15 VSS.n14 2.6005
R40 VSS.n26 VSS.n16 2.6005
R41 VSS.n29 VSS.n28 2.6005
R42 VSS.n28 VSS.n27 2.6005
R43 VSS.n25 VSS.n24 2.6005
R44 VSS.n24 VSS.n23 2.6005
R45 VSS.n22 VSS.n21 2.6005
R46 VSS.n21 VSS.n20 2.6005
R47 VSS.n18 VSS.n17 2.6005
R48 VSS.n5 VSS.n4 1.64943
R49 VSS.n19 VSS.n18 1.64943
R50 VSS.n22 VSS.n19 0.559135
R51 VSS.n6 VSS.n5 0.541457
R52 VSS.n12 VSS.n9 0.0760357
R53 VSS.n13 VSS.n12 0.0760357
R54 VSS VSS.n29 0.0760357
R55 VSS.n29 VSS.n25 0.0760357
R56 VSS.n25 VSS.n22 0.0760357
R57 VSS.n13 VSS.n2 0.0712143
R58 VSS.n9 VSS.n6 0.0181786
R59 VSS VSS.n2 0.00532143
R60 VDD.t0 VDD.n5 179.732
R61 VDD.n3 VDD.t3 58.0931
R62 VDD.n8 VDD.t5 56.5038
R63 VDD.n6 VDD.n4 8.2255
R64 VDD.n12 VDD.n6 8.2255
R65 VDD VDD.n6 6.3005
R66 VDD VDD.n6 6.3005
R67 VDD.n7 VDD.t6 4.7492
R68 VDD.n5 VDD.n4 3.1505
R69 VDD.n6 VDD.t0 3.1505
R70 VDD.n13 VDD.n12 3.1505
R71 VDD.n12 VDD.n11 3.1505
R72 VDD.n10 VDD.n9 3.1505
R73 VDD.n2 VDD.n1 2.9292
R74 VDD.n4 VDD.n3 1.87106
R75 VDD.n1 VDD.t4 1.8205
R76 VDD.n1 VDD.n0 1.8205
R77 VDD.n3 VDD.n2 0.578642
R78 VDD.n9 VDD.n8 0.134373
R79 VDD VDD.n13 0.0760357
R80 VDD.n13 VDD.n10 0.0760357
R81 VDD VDD.n2 0.0647857
R82 VDD.n10 VDD.n7 0.0422857
R83 B B.n0 56.3872
R84 B.t2 B.t1 55.0112
R85 B.n0 B.t0 29.9826
R86 B.n0 B.t2 9.1255
R87 OUT.n2 OUT.n0 7.06041
R88 OUT.n2 OUT.n1 5.10528
R89 OUT OUT.n2 0.0533261
C0 OUT B 6.21e-19
C1 OUT A 2.75e-19
C2 A B 0.0624f
C3 OUT VDD 0.149f
C4 B VDD 0.106f
C5 A VDD 0.149f
.ends

