magic
tech gf180mcuC
magscale 1 10
timestamp 1695206022
<< nwell >>
rect 513 3697 734 3781
rect 287 3666 734 3697
rect 287 3660 732 3666
rect 287 3631 800 3660
rect 287 3510 1159 3631
rect 355 3496 1159 3510
rect 355 3473 800 3496
rect 1715 3243 2123 3344
rect 284 3124 350 3185
rect 146 1886 222 1938
rect 1462 1845 1555 1917
rect 10650 1013 10883 1075
rect 11442 1018 11748 1085
rect 10648 902 10967 1013
rect 11442 909 11754 1018
<< psubdiff >>
rect 1182 2200 1666 2384
<< polysilicon >>
rect 284 3124 350 3185
<< metal1 >>
rect 1867 5242 1955 5260
rect 1867 5188 1879 5242
rect 1939 5188 1955 5242
rect 1867 5175 1955 5188
rect 2317 5250 3447 5475
rect 3595 5386 3676 5401
rect 3595 5333 3611 5386
rect 3664 5333 3676 5386
rect 3595 5310 3676 5333
rect 2317 5249 3712 5250
rect 3782 5249 15023 5476
rect 2317 5140 15023 5249
rect 2322 5139 15022 5140
rect 88 5082 225 5104
rect 88 4995 118 5082
rect 203 5070 225 5082
rect 2127 5073 2221 5091
rect 2127 5070 2148 5073
rect 203 4995 2148 5070
rect 88 4991 2148 4995
rect 88 4971 225 4991
rect 2127 4986 2148 4991
rect 2210 4986 2221 5073
rect 2127 4970 2221 4986
rect 1970 4921 2036 4923
rect 2363 4921 2472 5139
rect 2617 5034 2671 5139
rect 3166 5046 3217 5050
rect 2780 5034 2826 5045
rect 2940 5034 2986 5045
rect 3099 5034 3217 5046
rect 2617 4928 2620 5034
rect 2666 4928 2671 5034
rect 3099 4928 3100 5034
rect 3146 4928 3217 5034
rect 2617 4922 2671 4928
rect 280 4867 369 4875
rect 1713 4867 1797 4875
rect 280 4862 1797 4867
rect 280 4798 292 4862
rect 353 4858 1797 4862
rect 353 4798 1723 4858
rect 280 4793 1723 4798
rect 280 4785 369 4793
rect 1713 4782 1723 4793
rect 1784 4782 1797 4858
rect 1713 4767 1797 4782
rect 1970 4869 2472 4921
rect 2620 4917 2666 4922
rect 2780 4917 2826 4928
rect 2940 4917 2986 4928
rect 3099 4916 3217 4928
rect 3341 5034 3395 5139
rect 3890 5046 3941 5050
rect 3504 5034 3550 5045
rect 3664 5034 3710 5045
rect 3823 5034 3941 5046
rect 3341 4928 3344 5034
rect 3390 4928 3395 5034
rect 3823 4928 3824 5034
rect 3870 4928 3941 5034
rect 3341 4922 3395 4928
rect 3344 4917 3390 4922
rect 3504 4917 3550 4928
rect 3664 4917 3710 4928
rect 3823 4916 3941 4928
rect 4065 4990 4119 5139
rect 4065 4928 4068 4990
rect 4114 4928 4119 4990
rect 4065 4922 4119 4928
rect 4217 4990 4286 5001
rect 4388 4991 4434 5001
rect 4217 4928 4228 4990
rect 4274 4928 4286 4990
rect 4068 4917 4114 4922
rect 325 4693 1663 4694
rect 1970 4693 2050 4869
rect 2135 4811 2218 4820
rect 2135 4737 2144 4811
rect 2206 4737 2218 4811
rect 2135 4725 2218 4737
rect 325 4687 2050 4693
rect -827 4544 2050 4687
rect -827 2417 -630 4544
rect 325 4393 2050 4544
rect -403 4239 -315 4248
rect -403 4227 -306 4239
rect -403 4171 -377 4227
rect -318 4171 -306 4227
rect -403 4156 -306 4171
rect -124 4222 -54 4234
rect -124 4167 -114 4222
rect -58 4167 -54 4222
rect -566 4082 -483 4087
rect -572 4078 -483 4082
rect -572 4014 -552 4078
rect -498 4014 -483 4078
rect -572 3998 -483 4014
rect -827 2404 -629 2417
rect -827 2331 -732 2404
rect -653 2331 -629 2404
rect -827 2321 -629 2331
rect -572 1940 -486 3998
rect -403 3088 -314 4156
rect -124 4155 -54 4167
rect 839 4215 922 4226
rect 839 4163 856 4215
rect 912 4163 922 4215
rect 2150 4196 2208 4725
rect 839 4147 922 4163
rect 1016 4150 1098 4155
rect 1016 4098 1034 4150
rect 1086 4098 1098 4150
rect 1598 4138 2208 4196
rect 2363 4162 2472 4869
rect 2646 4805 2727 4817
rect 3166 4812 3217 4916
rect 3166 4806 3320 4812
rect 2563 4803 2727 4805
rect 2563 4800 2664 4803
rect 2563 4746 2576 4800
rect 2630 4753 2664 4800
rect 2713 4753 2727 4803
rect 2630 4746 2727 4753
rect 2563 4738 2727 4746
rect 2646 4737 2727 4738
rect 2774 4793 3320 4806
rect 3370 4803 3451 4817
rect 3890 4812 3941 4916
rect 4217 4915 4286 4928
rect 4382 4990 4437 4991
rect 4382 4928 4388 4990
rect 4434 4928 4437 4990
rect 3890 4806 4048 4812
rect 3370 4793 3388 4803
rect 2774 4757 3388 4793
rect 2620 4600 2666 4604
rect 2774 4601 2826 4757
rect 2872 4710 2952 4711
rect 2872 4708 2971 4710
rect 2872 4705 2884 4708
rect 2872 4657 2883 4705
rect 2872 4656 2884 4657
rect 2936 4656 2971 4708
rect 2872 4653 2971 4656
rect 3019 4705 3120 4711
rect 3019 4657 3030 4705
rect 3019 4653 3031 4657
rect 3083 4654 3120 4705
rect 3083 4653 3095 4654
rect 3166 4606 3217 4757
rect 3274 4753 3388 4757
rect 3437 4753 3451 4803
rect 3274 4746 3451 4753
rect 3370 4737 3451 4746
rect 3498 4793 4048 4806
rect 4094 4803 4175 4817
rect 4382 4812 4437 4928
rect 4629 4990 4683 5139
rect 4629 4928 4632 4990
rect 4678 4928 4683 4990
rect 4629 4922 4683 4928
rect 4781 4990 4850 5001
rect 4952 4991 4998 5001
rect 4781 4928 4792 4990
rect 4838 4928 4850 4990
rect 4632 4917 4678 4922
rect 4781 4915 4850 4928
rect 4946 4990 5001 4991
rect 4946 4928 4952 4990
rect 4998 4928 5001 4990
rect 4382 4806 4605 4812
rect 4094 4793 4112 4803
rect 3498 4757 4112 4793
rect 2615 4593 2672 4600
rect 2615 4459 2620 4593
rect 2666 4459 2672 4593
rect 2769 4593 2836 4601
rect 2940 4598 2986 4604
rect 2769 4526 2780 4593
rect 2826 4526 2836 4593
rect 2937 4593 2994 4598
rect 2937 4459 2940 4593
rect 2986 4459 2994 4593
rect 2615 4363 2672 4459
rect 2780 4448 2826 4459
rect 2937 4363 2994 4459
rect 3098 4593 3217 4606
rect 3344 4600 3390 4604
rect 3498 4601 3550 4757
rect 3743 4705 3844 4711
rect 3743 4657 3754 4705
rect 3743 4653 3755 4657
rect 3807 4654 3844 4705
rect 3807 4653 3819 4654
rect 3890 4606 3941 4757
rect 4002 4753 4112 4757
rect 4161 4753 4175 4803
rect 4002 4746 4175 4753
rect 4094 4737 4175 4746
rect 4222 4793 4605 4806
rect 4658 4803 4739 4817
rect 4946 4812 5001 4928
rect 4658 4793 4676 4803
rect 4222 4757 4676 4793
rect 3098 4459 3100 4593
rect 3146 4459 3217 4593
rect 3098 4441 3217 4459
rect 3339 4593 3396 4600
rect 3339 4459 3344 4593
rect 3390 4459 3396 4593
rect 3339 4363 3396 4459
rect 3493 4593 3560 4601
rect 3664 4598 3710 4604
rect 3493 4510 3504 4593
rect 3493 4458 3497 4510
rect 3550 4459 3560 4593
rect 3549 4458 3560 4459
rect 3493 4446 3560 4458
rect 3661 4593 3718 4598
rect 3661 4459 3664 4593
rect 3710 4459 3718 4593
rect 3661 4363 3718 4459
rect 3822 4593 3941 4606
rect 4068 4600 4114 4604
rect 4222 4601 4274 4757
rect 4549 4753 4676 4757
rect 4725 4753 4739 4803
rect 4549 4746 4739 4753
rect 4658 4737 4739 4746
rect 4786 4811 5116 4812
rect 4786 4759 4800 4811
rect 4852 4759 5045 4811
rect 5100 4759 5116 4811
rect 4786 4757 5116 4759
rect 4342 4710 4422 4711
rect 4342 4705 4496 4710
rect 4342 4657 4357 4705
rect 4342 4653 4358 4657
rect 4410 4653 4496 4705
rect 3822 4459 3824 4593
rect 3870 4459 3941 4593
rect 3822 4441 3941 4459
rect 4063 4593 4120 4600
rect 4063 4459 4068 4593
rect 4114 4459 4120 4593
rect 4217 4593 4284 4601
rect 4388 4598 4434 4604
rect 4632 4600 4678 4604
rect 4786 4601 4838 4757
rect 4906 4710 4986 4711
rect 4906 4657 4921 4710
rect 4973 4658 5060 4710
rect 4969 4657 5060 4658
rect 4906 4653 5060 4657
rect 4217 4526 4228 4593
rect 4274 4526 4284 4593
rect 4385 4593 4442 4598
rect 4385 4459 4388 4593
rect 4434 4459 4442 4593
rect 4063 4363 4120 4459
rect 4228 4448 4274 4459
rect 4385 4363 4442 4459
rect 4627 4593 4684 4600
rect 4627 4459 4632 4593
rect 4678 4459 4684 4593
rect 4781 4593 4848 4601
rect 4952 4598 4998 4604
rect 4781 4526 4792 4593
rect 4838 4526 4848 4593
rect 4949 4593 5006 4598
rect 4949 4459 4952 4593
rect 4998 4459 5006 4593
rect 4627 4363 4684 4459
rect 4792 4448 4838 4459
rect 4949 4363 5006 4459
rect 5149 4547 5259 4563
rect 5149 4464 5169 4547
rect 5241 4464 5259 4547
rect 5149 4453 5259 4464
rect 2519 4343 5094 4363
rect 2519 4297 2668 4343
rect 2895 4297 3392 4343
rect 3619 4297 4116 4343
rect 4343 4297 4680 4343
rect 4907 4297 5094 4343
rect 2519 4254 5094 4297
rect 2519 4208 5095 4254
rect 1016 4093 1098 4098
rect 2363 4018 4934 4162
rect 2363 3976 2527 4018
rect 2123 3942 2527 3976
rect 2123 3896 2174 3942
rect 2464 3896 2527 3942
rect 2123 3870 2527 3896
rect 2623 3937 2677 4018
rect 3172 3949 3223 3953
rect 2786 3937 2832 3948
rect 2946 3937 2992 3948
rect 3105 3937 3223 3949
rect 2207 3787 2274 3870
rect 2623 3831 2626 3937
rect 2672 3831 2677 3937
rect 3105 3831 3106 3937
rect 3152 3831 3223 3937
rect 2623 3825 2677 3831
rect 2626 3820 2672 3825
rect 2786 3820 2832 3831
rect 2946 3820 2992 3831
rect 3105 3819 3223 3831
rect 3347 3893 3401 4018
rect 3347 3831 3350 3893
rect 3396 3831 3401 3893
rect 3347 3825 3401 3831
rect 3499 3893 3568 3904
rect 3670 3894 3716 3904
rect 3499 3831 3510 3893
rect 3556 3831 3568 3893
rect 3350 3820 3396 3825
rect 2207 3741 2218 3787
rect 2264 3741 2275 3787
rect 2375 3741 2386 3787
rect 2432 3741 2443 3787
rect 1868 3663 2334 3673
rect 287 3631 1020 3637
rect 287 3621 1159 3631
rect 112 3496 1159 3621
rect 1868 3609 1879 3663
rect 1939 3660 2334 3663
rect 1939 3659 2272 3660
rect 1939 3609 2270 3659
rect 1868 3607 2270 3609
rect 2328 3614 2334 3660
rect 2322 3607 2334 3614
rect 1868 3601 2334 3607
rect 2380 3670 2443 3741
rect 2597 3720 2683 3721
rect 2597 3718 2733 3720
rect 2380 3612 2527 3670
rect 2597 3666 2610 3718
rect 2673 3706 2733 3718
rect 3172 3715 3223 3819
rect 3499 3818 3568 3831
rect 3664 3893 3719 3894
rect 3664 3831 3670 3893
rect 3716 3831 3719 3893
rect 3172 3709 3329 3715
rect 2597 3656 2670 3666
rect 2719 3656 2733 3706
rect 2597 3647 2733 3656
rect 2652 3640 2733 3647
rect 2780 3696 3329 3709
rect 3376 3706 3457 3720
rect 3664 3715 3719 3831
rect 3911 3893 3965 4018
rect 3911 3831 3914 3893
rect 3960 3831 3965 3893
rect 3911 3825 3965 3831
rect 4063 3893 4132 3904
rect 4234 3894 4280 3904
rect 4063 3831 4074 3893
rect 4120 3831 4132 3893
rect 3914 3820 3960 3825
rect 4063 3818 4132 3831
rect 4228 3893 4283 3894
rect 4228 3831 4234 3893
rect 4280 3831 4283 3893
rect 3664 3709 3787 3715
rect 3376 3696 3394 3706
rect 2780 3660 3394 3696
rect 112 3478 1020 3496
rect 132 3476 1020 3478
rect 132 3475 1018 3476
rect 310 3473 800 3475
rect 1274 3334 1353 3531
rect 2209 3496 2272 3509
rect 2209 3362 2222 3496
rect 2268 3362 2272 3496
rect 1715 3276 2123 3344
rect 2209 3276 2272 3362
rect 2380 3496 2443 3612
rect 2626 3503 2672 3507
rect 2780 3504 2832 3660
rect 2878 3613 2958 3614
rect 2878 3608 2977 3613
rect 2878 3560 2889 3608
rect 2878 3556 2890 3560
rect 2942 3556 2977 3608
rect 3025 3608 3048 3614
rect 3025 3560 3036 3608
rect 3100 3562 3126 3614
rect 3084 3560 3126 3562
rect 3025 3556 3126 3560
rect 3172 3509 3223 3660
rect 3283 3656 3394 3660
rect 3443 3656 3457 3706
rect 3283 3649 3457 3656
rect 3376 3640 3457 3649
rect 3504 3663 3787 3709
rect 3839 3696 3894 3715
rect 3940 3706 4021 3720
rect 4228 3715 4283 3831
rect 4475 3893 4529 4018
rect 4475 3831 4478 3893
rect 4524 3831 4529 3893
rect 4475 3825 4529 3831
rect 4627 3893 4696 3904
rect 4798 3894 4844 3904
rect 4627 3831 4638 3893
rect 4684 3831 4696 3893
rect 4478 3820 4524 3825
rect 4627 3818 4696 3831
rect 4792 3893 4847 3894
rect 4792 3831 4798 3893
rect 4844 3831 4847 3893
rect 4792 3724 4847 3831
rect 4792 3723 4962 3724
rect 4228 3709 4453 3715
rect 3940 3696 3958 3706
rect 3839 3663 3958 3696
rect 3504 3660 3958 3663
rect 2380 3479 2382 3496
rect 2428 3479 2443 3496
rect 2380 3427 2381 3479
rect 2433 3427 2443 3479
rect 2380 3362 2382 3427
rect 2428 3362 2443 3427
rect 2380 3351 2443 3362
rect 2621 3496 2678 3503
rect 2621 3362 2626 3496
rect 2672 3362 2678 3496
rect 2775 3496 2842 3504
rect 2946 3501 2992 3507
rect 2775 3429 2786 3496
rect 2832 3429 2842 3496
rect 2943 3496 3000 3501
rect 2943 3362 2946 3496
rect 2992 3362 3000 3496
rect 1715 3266 2527 3276
rect 2621 3266 2678 3362
rect 2786 3351 2832 3362
rect 2943 3266 3000 3362
rect 3104 3496 3223 3509
rect 3350 3503 3396 3507
rect 3504 3504 3556 3660
rect 3832 3656 3958 3660
rect 4007 3656 4021 3706
rect 3832 3649 4021 3656
rect 3940 3640 4021 3649
rect 4068 3696 4453 3709
rect 4504 3706 4585 3720
rect 4792 3709 4858 3723
rect 4504 3696 4522 3706
rect 4068 3660 4522 3696
rect 3624 3613 3704 3614
rect 3624 3608 3778 3613
rect 3624 3560 3639 3608
rect 3624 3556 3640 3560
rect 3692 3556 3778 3608
rect 3104 3362 3106 3496
rect 3152 3362 3223 3496
rect 3104 3344 3223 3362
rect 3345 3496 3402 3503
rect 3345 3362 3350 3496
rect 3396 3362 3402 3496
rect 3499 3496 3566 3504
rect 3670 3501 3716 3507
rect 3914 3503 3960 3507
rect 4068 3504 4120 3660
rect 4397 3656 4522 3660
rect 4571 3656 4585 3706
rect 4397 3649 4585 3656
rect 4504 3640 4585 3649
rect 4632 3671 4858 3709
rect 4910 3671 4962 3723
rect 4632 3660 4962 3671
rect 4188 3613 4268 3614
rect 4188 3608 4342 3613
rect 4188 3560 4203 3608
rect 4188 3556 4204 3560
rect 4256 3556 4342 3608
rect 3499 3429 3510 3496
rect 3556 3429 3566 3496
rect 3667 3496 3724 3501
rect 3667 3362 3670 3496
rect 3716 3362 3724 3496
rect 3345 3266 3402 3362
rect 3510 3351 3556 3362
rect 3667 3266 3724 3362
rect 3909 3496 3966 3503
rect 3909 3362 3914 3496
rect 3960 3362 3966 3496
rect 4063 3496 4130 3504
rect 4234 3501 4280 3507
rect 4478 3503 4524 3507
rect 4632 3504 4684 3660
rect 4752 3613 4832 3614
rect 4752 3611 4906 3613
rect 4752 3559 4764 3611
rect 4816 3559 4906 3611
rect 4752 3556 4906 3559
rect 4063 3429 4074 3496
rect 4120 3429 4130 3496
rect 4231 3496 4288 3501
rect 4231 3362 4234 3496
rect 4280 3362 4288 3496
rect 3909 3266 3966 3362
rect 4074 3351 4120 3362
rect 4231 3266 4288 3362
rect 4473 3496 4530 3503
rect 4473 3362 4478 3496
rect 4524 3362 4530 3496
rect 4627 3496 4694 3504
rect 4798 3501 4844 3507
rect 4627 3429 4638 3496
rect 4684 3429 4694 3496
rect 4795 3496 4852 3501
rect 4795 3362 4798 3496
rect 4844 3362 4852 3496
rect 4473 3266 4530 3362
rect 4638 3351 4684 3362
rect 4795 3266 4852 3362
rect 5008 3266 5094 4208
rect 5149 3675 5204 4453
rect 5454 4164 5607 5139
rect 5752 5036 5806 5139
rect 6301 5048 6352 5052
rect 5915 5036 5961 5047
rect 6075 5036 6121 5047
rect 6234 5036 6352 5048
rect 5752 4930 5755 5036
rect 5801 4930 5806 5036
rect 6234 4930 6235 5036
rect 6281 4930 6352 5036
rect 5752 4924 5806 4930
rect 5755 4919 5801 4924
rect 5915 4919 5961 4930
rect 6075 4919 6121 4930
rect 6234 4918 6352 4930
rect 6476 5036 6530 5139
rect 7025 5048 7076 5052
rect 6639 5036 6685 5047
rect 6799 5036 6845 5047
rect 6958 5036 7076 5048
rect 6476 4930 6479 5036
rect 6525 4930 6530 5036
rect 6958 4930 6959 5036
rect 7005 4930 7076 5036
rect 6476 4924 6530 4930
rect 6479 4919 6525 4924
rect 6639 4919 6685 4930
rect 6799 4919 6845 4930
rect 6958 4918 7076 4930
rect 7200 4992 7254 5139
rect 7200 4930 7203 4992
rect 7249 4930 7254 4992
rect 7200 4924 7254 4930
rect 7352 4992 7421 5003
rect 7523 4993 7569 5003
rect 7352 4930 7363 4992
rect 7409 4930 7421 4992
rect 7203 4919 7249 4924
rect 5781 4807 5862 4819
rect 6301 4814 6352 4918
rect 6301 4808 6455 4814
rect 5698 4805 5862 4807
rect 5698 4802 5799 4805
rect 5698 4748 5711 4802
rect 5765 4755 5799 4802
rect 5848 4755 5862 4805
rect 5765 4748 5862 4755
rect 5698 4740 5862 4748
rect 5781 4739 5862 4740
rect 5909 4795 6455 4808
rect 6505 4805 6586 4819
rect 7025 4814 7076 4918
rect 7352 4917 7421 4930
rect 7517 4992 7572 4993
rect 7517 4930 7523 4992
rect 7569 4930 7572 4992
rect 7025 4808 7183 4814
rect 6505 4795 6523 4805
rect 5909 4759 6523 4795
rect 5755 4602 5801 4606
rect 5909 4603 5961 4759
rect 6007 4712 6087 4713
rect 6007 4710 6106 4712
rect 6007 4707 6019 4710
rect 6007 4659 6018 4707
rect 6007 4658 6019 4659
rect 6071 4658 6106 4710
rect 6007 4655 6106 4658
rect 6154 4707 6255 4713
rect 6154 4659 6165 4707
rect 6154 4655 6166 4659
rect 6218 4656 6255 4707
rect 6218 4655 6230 4656
rect 6301 4608 6352 4759
rect 6409 4755 6523 4759
rect 6572 4755 6586 4805
rect 6409 4748 6586 4755
rect 6505 4739 6586 4748
rect 6633 4795 7183 4808
rect 7229 4805 7310 4819
rect 7517 4814 7572 4930
rect 7764 4992 7818 5139
rect 7764 4930 7767 4992
rect 7813 4930 7818 4992
rect 7764 4924 7818 4930
rect 7916 4992 7985 5003
rect 8087 4993 8133 5003
rect 7916 4930 7927 4992
rect 7973 4930 7985 4992
rect 7767 4919 7813 4924
rect 7916 4917 7985 4930
rect 8081 4992 8136 4993
rect 8081 4930 8087 4992
rect 8133 4930 8136 4992
rect 7517 4808 7740 4814
rect 7229 4795 7247 4805
rect 6633 4759 7247 4795
rect 5750 4595 5807 4602
rect 5750 4461 5755 4595
rect 5801 4461 5807 4595
rect 5904 4595 5971 4603
rect 6075 4600 6121 4606
rect 5904 4528 5915 4595
rect 5961 4528 5971 4595
rect 6072 4595 6129 4600
rect 6072 4461 6075 4595
rect 6121 4461 6129 4595
rect 5750 4365 5807 4461
rect 5915 4450 5961 4461
rect 6072 4365 6129 4461
rect 6233 4595 6352 4608
rect 6479 4602 6525 4606
rect 6633 4603 6685 4759
rect 6878 4707 6979 4713
rect 6878 4659 6889 4707
rect 6878 4655 6890 4659
rect 6942 4656 6979 4707
rect 6942 4655 6954 4656
rect 7025 4608 7076 4759
rect 7137 4755 7247 4759
rect 7296 4755 7310 4805
rect 7137 4748 7310 4755
rect 7229 4739 7310 4748
rect 7357 4795 7740 4808
rect 7793 4805 7874 4819
rect 8081 4814 8136 4930
rect 7793 4795 7811 4805
rect 7357 4759 7811 4795
rect 6233 4461 6235 4595
rect 6281 4461 6352 4595
rect 6233 4443 6352 4461
rect 6474 4595 6531 4602
rect 6474 4461 6479 4595
rect 6525 4461 6531 4595
rect 6474 4365 6531 4461
rect 6628 4595 6695 4603
rect 6799 4600 6845 4606
rect 6628 4512 6639 4595
rect 6628 4460 6632 4512
rect 6685 4461 6695 4595
rect 6684 4460 6695 4461
rect 6628 4448 6695 4460
rect 6796 4595 6853 4600
rect 6796 4461 6799 4595
rect 6845 4461 6853 4595
rect 6796 4365 6853 4461
rect 6957 4595 7076 4608
rect 7203 4602 7249 4606
rect 7357 4603 7409 4759
rect 7684 4755 7811 4759
rect 7860 4755 7874 4805
rect 7684 4748 7874 4755
rect 7793 4739 7874 4748
rect 7921 4813 8251 4814
rect 7921 4761 7935 4813
rect 7987 4761 8251 4813
rect 7921 4759 8251 4761
rect 7477 4712 7557 4713
rect 7477 4707 7631 4712
rect 7477 4659 7492 4707
rect 7477 4655 7493 4659
rect 7545 4655 7631 4707
rect 6957 4461 6959 4595
rect 7005 4461 7076 4595
rect 6957 4443 7076 4461
rect 7198 4595 7255 4602
rect 7198 4461 7203 4595
rect 7249 4461 7255 4595
rect 7352 4595 7419 4603
rect 7523 4600 7569 4606
rect 7767 4602 7813 4606
rect 7921 4603 7973 4759
rect 8041 4712 8121 4713
rect 8041 4659 8056 4712
rect 8108 4660 8195 4712
rect 8104 4659 8195 4660
rect 8041 4655 8195 4659
rect 7352 4528 7363 4595
rect 7409 4528 7419 4595
rect 7520 4595 7577 4600
rect 7520 4461 7523 4595
rect 7569 4461 7577 4595
rect 7198 4365 7255 4461
rect 7363 4450 7409 4461
rect 7520 4365 7577 4461
rect 7762 4595 7819 4602
rect 7762 4461 7767 4595
rect 7813 4461 7819 4595
rect 7916 4595 7983 4603
rect 8087 4600 8133 4606
rect 7916 4528 7927 4595
rect 7973 4528 7983 4595
rect 8084 4595 8141 4600
rect 8084 4461 8087 4595
rect 8133 4461 8141 4595
rect 7762 4365 7819 4461
rect 7927 4450 7973 4461
rect 8084 4365 8141 4461
rect 5654 4345 8229 4365
rect 5654 4299 5803 4345
rect 6030 4299 6527 4345
rect 6754 4299 7251 4345
rect 7478 4299 7815 4345
rect 8042 4299 8229 4345
rect 5654 4256 8229 4299
rect 5654 4210 8230 4256
rect 5454 4160 8069 4164
rect 5454 4019 8092 4160
rect 5454 3978 5662 4019
rect 5258 3944 5662 3978
rect 5258 3898 5309 3944
rect 5599 3898 5662 3944
rect 5258 3872 5662 3898
rect 5758 3939 5812 4019
rect 6307 3951 6358 3955
rect 5921 3939 5967 3950
rect 6081 3939 6127 3950
rect 6240 3939 6358 3951
rect 5342 3789 5409 3872
rect 5758 3833 5761 3939
rect 5807 3833 5812 3939
rect 6240 3833 6241 3939
rect 6287 3833 6358 3939
rect 5758 3827 5812 3833
rect 5761 3822 5807 3827
rect 5921 3822 5967 3833
rect 6081 3822 6127 3833
rect 6240 3821 6358 3833
rect 6482 3895 6536 4019
rect 6482 3833 6485 3895
rect 6531 3833 6536 3895
rect 6482 3827 6536 3833
rect 6634 3895 6703 3906
rect 6805 3896 6851 3906
rect 6634 3833 6645 3895
rect 6691 3833 6703 3895
rect 6485 3822 6531 3827
rect 5342 3743 5353 3789
rect 5399 3743 5410 3789
rect 5510 3743 5521 3789
rect 5567 3743 5578 3789
rect 5149 3662 5469 3675
rect 5149 3661 5407 3662
rect 5149 3609 5405 3661
rect 5463 3616 5469 3662
rect 5457 3609 5469 3616
rect 5149 3603 5469 3609
rect 5515 3672 5578 3743
rect 5732 3722 5818 3723
rect 5732 3720 5868 3722
rect 5515 3614 5662 3672
rect 5732 3668 5745 3720
rect 5808 3708 5868 3720
rect 6307 3717 6358 3821
rect 6634 3820 6703 3833
rect 6799 3895 6854 3896
rect 6799 3833 6805 3895
rect 6851 3833 6854 3895
rect 6307 3711 6464 3717
rect 5732 3658 5805 3668
rect 5854 3658 5868 3708
rect 5732 3649 5868 3658
rect 5787 3642 5868 3649
rect 5915 3698 6464 3711
rect 6511 3708 6592 3722
rect 6799 3717 6854 3833
rect 7046 3895 7100 4019
rect 7046 3833 7049 3895
rect 7095 3833 7100 3895
rect 7046 3827 7100 3833
rect 7198 3895 7267 3906
rect 7369 3896 7415 3906
rect 7198 3833 7209 3895
rect 7255 3833 7267 3895
rect 7049 3822 7095 3827
rect 7198 3820 7267 3833
rect 7363 3895 7418 3896
rect 7363 3833 7369 3895
rect 7415 3833 7418 3895
rect 6799 3711 6922 3717
rect 6511 3698 6529 3708
rect 5915 3662 6529 3698
rect 5149 3602 5204 3603
rect 5344 3498 5407 3511
rect 5344 3364 5357 3498
rect 5403 3364 5407 3498
rect 5344 3278 5407 3364
rect 5515 3498 5578 3614
rect 5761 3505 5807 3509
rect 5915 3506 5967 3662
rect 6013 3615 6093 3616
rect 6013 3610 6112 3615
rect 6013 3562 6024 3610
rect 6013 3558 6025 3562
rect 6077 3558 6112 3610
rect 6160 3610 6183 3616
rect 6160 3562 6171 3610
rect 6235 3564 6261 3616
rect 6219 3562 6261 3564
rect 6160 3558 6261 3562
rect 6307 3511 6358 3662
rect 6418 3658 6529 3662
rect 6578 3658 6592 3708
rect 6418 3651 6592 3658
rect 6511 3642 6592 3651
rect 6639 3665 6922 3711
rect 6974 3698 7029 3717
rect 7075 3708 7156 3722
rect 7363 3717 7418 3833
rect 7610 3895 7664 4019
rect 7610 3833 7613 3895
rect 7659 3833 7664 3895
rect 7610 3827 7664 3833
rect 7762 3895 7831 3906
rect 7933 3896 7979 3906
rect 7762 3833 7773 3895
rect 7819 3833 7831 3895
rect 7613 3822 7659 3827
rect 7762 3820 7831 3833
rect 7927 3895 7982 3896
rect 7927 3833 7933 3895
rect 7979 3833 7982 3895
rect 7927 3726 7982 3833
rect 7927 3725 8097 3726
rect 7363 3711 7588 3717
rect 7075 3698 7093 3708
rect 6974 3665 7093 3698
rect 6639 3662 7093 3665
rect 5515 3481 5517 3498
rect 5563 3481 5578 3498
rect 5515 3429 5516 3481
rect 5568 3429 5578 3481
rect 5515 3364 5517 3429
rect 5563 3364 5578 3429
rect 5515 3353 5578 3364
rect 5756 3498 5813 3505
rect 5756 3364 5761 3498
rect 5807 3364 5813 3498
rect 5910 3498 5977 3506
rect 6081 3503 6127 3509
rect 5910 3431 5921 3498
rect 5967 3431 5977 3498
rect 6078 3498 6135 3503
rect 6078 3364 6081 3498
rect 6127 3364 6135 3498
rect 1715 3263 5094 3266
rect 1715 3243 2176 3263
rect 2123 3207 2176 3243
rect 2470 3254 5094 3263
rect 5258 3268 5662 3278
rect 5756 3268 5813 3364
rect 5921 3353 5967 3364
rect 6078 3268 6135 3364
rect 6239 3498 6358 3511
rect 6485 3505 6531 3509
rect 6639 3506 6691 3662
rect 6967 3658 7093 3662
rect 7142 3658 7156 3708
rect 6967 3651 7156 3658
rect 7075 3642 7156 3651
rect 7203 3698 7588 3711
rect 7639 3708 7720 3722
rect 7927 3711 7993 3725
rect 7639 3698 7657 3708
rect 7203 3662 7657 3698
rect 6759 3615 6839 3616
rect 6759 3610 6913 3615
rect 6759 3562 6774 3610
rect 6759 3558 6775 3562
rect 6827 3558 6913 3610
rect 6239 3364 6241 3498
rect 6287 3364 6358 3498
rect 6239 3346 6358 3364
rect 6480 3498 6537 3505
rect 6480 3364 6485 3498
rect 6531 3364 6537 3498
rect 6634 3498 6701 3506
rect 6805 3503 6851 3509
rect 7049 3505 7095 3509
rect 7203 3506 7255 3662
rect 7532 3658 7657 3662
rect 7706 3658 7720 3708
rect 7532 3651 7720 3658
rect 7639 3642 7720 3651
rect 7767 3673 7993 3711
rect 8045 3673 8097 3725
rect 7767 3662 8097 3673
rect 7323 3615 7403 3616
rect 7323 3610 7477 3615
rect 7323 3562 7338 3610
rect 7323 3558 7339 3562
rect 7391 3558 7477 3610
rect 6634 3431 6645 3498
rect 6691 3431 6701 3498
rect 6802 3498 6859 3503
rect 6802 3364 6805 3498
rect 6851 3364 6859 3498
rect 6480 3268 6537 3364
rect 6645 3353 6691 3364
rect 6802 3268 6859 3364
rect 7044 3498 7101 3505
rect 7044 3364 7049 3498
rect 7095 3364 7101 3498
rect 7198 3498 7265 3506
rect 7369 3503 7415 3509
rect 7613 3505 7659 3509
rect 7767 3506 7819 3662
rect 7887 3615 7967 3616
rect 7887 3613 8041 3615
rect 7887 3561 7899 3613
rect 7951 3561 8041 3613
rect 7887 3558 8041 3561
rect 7198 3431 7209 3498
rect 7255 3431 7265 3498
rect 7366 3498 7423 3503
rect 7366 3364 7369 3498
rect 7415 3364 7423 3498
rect 7044 3268 7101 3364
rect 7209 3353 7255 3364
rect 7366 3268 7423 3364
rect 7608 3498 7665 3505
rect 7608 3364 7613 3498
rect 7659 3364 7665 3498
rect 7762 3498 7829 3506
rect 7933 3503 7979 3509
rect 7762 3431 7773 3498
rect 7819 3431 7829 3498
rect 7930 3498 7987 3503
rect 7930 3364 7933 3498
rect 7979 3364 7987 3498
rect 7608 3268 7665 3364
rect 7773 3353 7819 3364
rect 7930 3268 7987 3364
rect 8143 3268 8229 4210
rect 8596 4162 8721 5139
rect 8866 5034 8920 5139
rect 9415 5046 9466 5050
rect 9029 5034 9075 5045
rect 9189 5034 9235 5045
rect 9348 5034 9466 5046
rect 8866 4928 8869 5034
rect 8915 4928 8920 5034
rect 9348 4928 9349 5034
rect 9395 4928 9466 5034
rect 8866 4922 8920 4928
rect 8869 4917 8915 4922
rect 9029 4917 9075 4928
rect 9189 4917 9235 4928
rect 9348 4916 9466 4928
rect 9590 5034 9644 5139
rect 10139 5046 10190 5050
rect 9753 5034 9799 5045
rect 9913 5034 9959 5045
rect 10072 5034 10190 5046
rect 9590 4928 9593 5034
rect 9639 4928 9644 5034
rect 10072 4928 10073 5034
rect 10119 4928 10190 5034
rect 9590 4922 9644 4928
rect 9593 4917 9639 4922
rect 9753 4917 9799 4928
rect 9913 4917 9959 4928
rect 10072 4916 10190 4928
rect 10314 4990 10368 5139
rect 10314 4928 10317 4990
rect 10363 4928 10368 4990
rect 10314 4922 10368 4928
rect 10466 4990 10535 5001
rect 10637 4991 10683 5001
rect 10466 4928 10477 4990
rect 10523 4928 10535 4990
rect 10317 4917 10363 4922
rect 8895 4805 8976 4817
rect 9415 4812 9466 4916
rect 9415 4806 9569 4812
rect 8812 4803 8976 4805
rect 8812 4800 8913 4803
rect 8812 4746 8825 4800
rect 8879 4753 8913 4800
rect 8962 4753 8976 4803
rect 8879 4746 8976 4753
rect 8812 4738 8976 4746
rect 8895 4737 8976 4738
rect 9023 4793 9569 4806
rect 9619 4803 9700 4817
rect 10139 4812 10190 4916
rect 10466 4915 10535 4928
rect 10631 4990 10686 4991
rect 10631 4928 10637 4990
rect 10683 4928 10686 4990
rect 10139 4806 10297 4812
rect 9619 4793 9637 4803
rect 9023 4757 9637 4793
rect 8869 4600 8915 4604
rect 9023 4601 9075 4757
rect 9121 4710 9201 4711
rect 9121 4708 9220 4710
rect 9121 4705 9133 4708
rect 9121 4657 9132 4705
rect 9121 4656 9133 4657
rect 9185 4656 9220 4708
rect 9121 4653 9220 4656
rect 9268 4705 9369 4711
rect 9268 4657 9279 4705
rect 9268 4653 9280 4657
rect 9332 4654 9369 4705
rect 9332 4653 9344 4654
rect 9415 4606 9466 4757
rect 9523 4753 9637 4757
rect 9686 4753 9700 4803
rect 9523 4746 9700 4753
rect 9619 4737 9700 4746
rect 9747 4793 10297 4806
rect 10343 4803 10424 4817
rect 10631 4812 10686 4928
rect 10878 4990 10932 5139
rect 10878 4928 10881 4990
rect 10927 4928 10932 4990
rect 10878 4922 10932 4928
rect 11030 4990 11099 5001
rect 11201 4991 11247 5001
rect 11030 4928 11041 4990
rect 11087 4928 11099 4990
rect 10881 4917 10927 4922
rect 11030 4915 11099 4928
rect 11195 4990 11250 4991
rect 11195 4928 11201 4990
rect 11247 4928 11250 4990
rect 10631 4806 10854 4812
rect 10343 4793 10361 4803
rect 9747 4757 10361 4793
rect 8864 4593 8921 4600
rect 8864 4459 8869 4593
rect 8915 4459 8921 4593
rect 9018 4593 9085 4601
rect 9189 4598 9235 4604
rect 9018 4526 9029 4593
rect 9075 4526 9085 4593
rect 9186 4593 9243 4598
rect 9186 4459 9189 4593
rect 9235 4459 9243 4593
rect 8864 4363 8921 4459
rect 9029 4448 9075 4459
rect 9186 4363 9243 4459
rect 9347 4593 9466 4606
rect 9593 4600 9639 4604
rect 9747 4601 9799 4757
rect 9992 4705 10093 4711
rect 9992 4657 10003 4705
rect 9992 4653 10004 4657
rect 10056 4654 10093 4705
rect 10056 4653 10068 4654
rect 10139 4606 10190 4757
rect 10251 4753 10361 4757
rect 10410 4753 10424 4803
rect 10251 4746 10424 4753
rect 10343 4737 10424 4746
rect 10471 4793 10854 4806
rect 10907 4803 10988 4817
rect 11195 4812 11250 4928
rect 11584 4812 11663 4823
rect 10907 4793 10925 4803
rect 10471 4757 10925 4793
rect 9347 4459 9349 4593
rect 9395 4459 9466 4593
rect 9347 4441 9466 4459
rect 9588 4593 9645 4600
rect 9588 4459 9593 4593
rect 9639 4459 9645 4593
rect 9588 4363 9645 4459
rect 9742 4593 9809 4601
rect 9913 4598 9959 4604
rect 9742 4510 9753 4593
rect 9742 4458 9746 4510
rect 9799 4459 9809 4593
rect 9798 4458 9809 4459
rect 9742 4446 9809 4458
rect 9910 4593 9967 4598
rect 9910 4459 9913 4593
rect 9959 4459 9967 4593
rect 9910 4363 9967 4459
rect 10071 4593 10190 4606
rect 10317 4600 10363 4604
rect 10471 4601 10523 4757
rect 10798 4753 10925 4757
rect 10974 4753 10988 4803
rect 10798 4746 10988 4753
rect 10907 4737 10988 4746
rect 11035 4811 11663 4812
rect 11035 4759 11049 4811
rect 11101 4810 11663 4811
rect 11101 4759 11594 4810
rect 11035 4757 11594 4759
rect 11651 4757 11663 4810
rect 10591 4710 10671 4711
rect 10591 4705 10745 4710
rect 10591 4657 10606 4705
rect 10591 4653 10607 4657
rect 10659 4653 10745 4705
rect 10071 4459 10073 4593
rect 10119 4459 10190 4593
rect 10071 4441 10190 4459
rect 10312 4593 10369 4600
rect 10312 4459 10317 4593
rect 10363 4459 10369 4593
rect 10466 4593 10533 4601
rect 10637 4598 10683 4604
rect 10881 4600 10927 4604
rect 11035 4601 11087 4757
rect 11584 4745 11663 4757
rect 11155 4710 11235 4711
rect 11155 4657 11170 4710
rect 11222 4658 11309 4710
rect 11218 4657 11309 4658
rect 11155 4653 11309 4657
rect 10466 4526 10477 4593
rect 10523 4526 10533 4593
rect 10634 4593 10691 4598
rect 10634 4459 10637 4593
rect 10683 4459 10691 4593
rect 10312 4363 10369 4459
rect 10477 4448 10523 4459
rect 10634 4363 10691 4459
rect 10876 4593 10933 4600
rect 10876 4459 10881 4593
rect 10927 4459 10933 4593
rect 11030 4593 11097 4601
rect 11201 4598 11247 4604
rect 11030 4526 11041 4593
rect 11087 4526 11097 4593
rect 11198 4593 11255 4598
rect 11198 4459 11201 4593
rect 11247 4459 11255 4593
rect 10876 4363 10933 4459
rect 11041 4448 11087 4459
rect 11198 4363 11255 4459
rect 11372 4544 11479 4563
rect 11372 4480 11395 4544
rect 11456 4480 11479 4544
rect 11372 4454 11479 4480
rect 8768 4343 11343 4363
rect 8768 4297 8917 4343
rect 9144 4297 9641 4343
rect 9868 4297 10365 4343
rect 10592 4297 10929 4343
rect 11156 4297 11343 4343
rect 8768 4254 11343 4297
rect 8768 4208 11344 4254
rect 8596 4160 11183 4162
rect 8596 4019 11186 4160
rect 8596 3976 8776 4019
rect 8372 3942 8776 3976
rect 8372 3896 8423 3942
rect 8713 3896 8776 3942
rect 8372 3870 8776 3896
rect 8872 3937 8926 4019
rect 9421 3949 9472 3953
rect 9035 3937 9081 3948
rect 9195 3937 9241 3948
rect 9354 3937 9472 3949
rect 8456 3787 8523 3870
rect 8872 3831 8875 3937
rect 8921 3831 8926 3937
rect 9354 3831 9355 3937
rect 9401 3831 9472 3937
rect 8872 3825 8926 3831
rect 8875 3820 8921 3825
rect 9035 3820 9081 3831
rect 9195 3820 9241 3831
rect 9354 3819 9472 3831
rect 9596 3893 9650 4019
rect 9596 3831 9599 3893
rect 9645 3831 9650 3893
rect 9596 3825 9650 3831
rect 9748 3893 9817 3904
rect 9919 3894 9965 3904
rect 9748 3831 9759 3893
rect 9805 3831 9817 3893
rect 9599 3820 9645 3825
rect 8456 3741 8467 3787
rect 8513 3741 8524 3787
rect 8624 3741 8635 3787
rect 8681 3741 8692 3787
rect 8278 3665 8583 3673
rect 8278 3612 8289 3665
rect 8343 3660 8583 3665
rect 8343 3659 8521 3660
rect 8343 3612 8519 3659
rect 8278 3607 8519 3612
rect 8577 3614 8583 3660
rect 8571 3607 8583 3614
rect 8278 3601 8583 3607
rect 8629 3670 8692 3741
rect 8846 3720 8932 3721
rect 8846 3718 8982 3720
rect 8629 3612 8776 3670
rect 8846 3666 8859 3718
rect 8922 3706 8982 3718
rect 9421 3715 9472 3819
rect 9748 3818 9817 3831
rect 9913 3893 9968 3894
rect 9913 3831 9919 3893
rect 9965 3831 9968 3893
rect 9421 3709 9578 3715
rect 8846 3656 8919 3666
rect 8968 3656 8982 3706
rect 8846 3647 8982 3656
rect 8901 3640 8982 3647
rect 9029 3696 9578 3709
rect 9625 3706 9706 3720
rect 9913 3715 9968 3831
rect 10160 3893 10214 4019
rect 10160 3831 10163 3893
rect 10209 3831 10214 3893
rect 10160 3825 10214 3831
rect 10312 3893 10381 3904
rect 10483 3894 10529 3904
rect 10312 3831 10323 3893
rect 10369 3831 10381 3893
rect 10163 3820 10209 3825
rect 10312 3818 10381 3831
rect 10477 3893 10532 3894
rect 10477 3831 10483 3893
rect 10529 3831 10532 3893
rect 9913 3709 10036 3715
rect 9625 3696 9643 3706
rect 9029 3660 9643 3696
rect 8458 3496 8521 3509
rect 8458 3362 8471 3496
rect 8517 3362 8521 3496
rect 8458 3276 8521 3362
rect 8629 3496 8692 3612
rect 8875 3503 8921 3507
rect 9029 3504 9081 3660
rect 9127 3613 9207 3614
rect 9127 3608 9226 3613
rect 9127 3560 9138 3608
rect 9127 3556 9139 3560
rect 9191 3556 9226 3608
rect 9274 3608 9297 3614
rect 9274 3560 9285 3608
rect 9349 3562 9375 3614
rect 9333 3560 9375 3562
rect 9274 3556 9375 3560
rect 9421 3509 9472 3660
rect 9532 3656 9643 3660
rect 9692 3656 9706 3706
rect 9532 3649 9706 3656
rect 9625 3640 9706 3649
rect 9753 3663 10036 3709
rect 10088 3696 10143 3715
rect 10189 3706 10270 3720
rect 10477 3715 10532 3831
rect 10724 3893 10778 4019
rect 10724 3831 10727 3893
rect 10773 3831 10778 3893
rect 10724 3825 10778 3831
rect 10876 3893 10945 3904
rect 11047 3894 11093 3904
rect 10876 3831 10887 3893
rect 10933 3831 10945 3893
rect 10727 3820 10773 3825
rect 10876 3818 10945 3831
rect 11041 3893 11096 3894
rect 11041 3831 11047 3893
rect 11093 3831 11096 3893
rect 11041 3724 11096 3831
rect 11041 3723 11211 3724
rect 10477 3709 10702 3715
rect 10189 3696 10207 3706
rect 10088 3663 10207 3696
rect 9753 3660 10207 3663
rect 8629 3479 8631 3496
rect 8677 3479 8692 3496
rect 8629 3427 8630 3479
rect 8682 3427 8692 3479
rect 8629 3362 8631 3427
rect 8677 3362 8692 3427
rect 8629 3351 8692 3362
rect 8870 3496 8927 3503
rect 8870 3362 8875 3496
rect 8921 3362 8927 3496
rect 9024 3496 9091 3504
rect 9195 3501 9241 3507
rect 9024 3429 9035 3496
rect 9081 3429 9091 3496
rect 9192 3496 9249 3501
rect 9192 3362 9195 3496
rect 9241 3362 9249 3496
rect 5258 3265 8229 3268
rect 5258 3254 5311 3265
rect 2470 3246 5311 3254
rect 2470 3207 2674 3246
rect 2123 3200 2674 3207
rect 2901 3200 3398 3246
rect 3625 3200 3962 3246
rect 4189 3200 4526 3246
rect 4753 3209 5311 3246
rect 5605 3256 8229 3265
rect 8372 3266 8776 3276
rect 8870 3266 8927 3362
rect 9035 3351 9081 3362
rect 9192 3266 9249 3362
rect 9353 3496 9472 3509
rect 9599 3503 9645 3507
rect 9753 3504 9805 3660
rect 10081 3656 10207 3660
rect 10256 3656 10270 3706
rect 10081 3649 10270 3656
rect 10189 3640 10270 3649
rect 10317 3696 10702 3709
rect 10753 3706 10834 3720
rect 11041 3709 11107 3723
rect 10753 3696 10771 3706
rect 10317 3660 10771 3696
rect 9873 3613 9953 3614
rect 9873 3608 10027 3613
rect 9873 3560 9888 3608
rect 9873 3556 9889 3560
rect 9941 3556 10027 3608
rect 9353 3362 9355 3496
rect 9401 3362 9472 3496
rect 9353 3344 9472 3362
rect 9594 3496 9651 3503
rect 9594 3362 9599 3496
rect 9645 3362 9651 3496
rect 9748 3496 9815 3504
rect 9919 3501 9965 3507
rect 10163 3503 10209 3507
rect 10317 3504 10369 3660
rect 10646 3656 10771 3660
rect 10820 3656 10834 3706
rect 10646 3649 10834 3656
rect 10753 3640 10834 3649
rect 10881 3671 11107 3709
rect 11159 3671 11211 3723
rect 10881 3660 11211 3671
rect 10437 3613 10517 3614
rect 10437 3608 10591 3613
rect 10437 3560 10452 3608
rect 10437 3556 10453 3560
rect 10505 3556 10591 3608
rect 9748 3429 9759 3496
rect 9805 3429 9815 3496
rect 9916 3496 9973 3501
rect 9916 3362 9919 3496
rect 9965 3362 9973 3496
rect 9594 3266 9651 3362
rect 9759 3351 9805 3362
rect 9916 3266 9973 3362
rect 10158 3496 10215 3503
rect 10158 3362 10163 3496
rect 10209 3362 10215 3496
rect 10312 3496 10379 3504
rect 10483 3501 10529 3507
rect 10727 3503 10773 3507
rect 10881 3504 10933 3660
rect 11001 3613 11081 3614
rect 11001 3611 11155 3613
rect 11001 3559 11013 3611
rect 11065 3559 11155 3611
rect 11001 3556 11155 3559
rect 10312 3429 10323 3496
rect 10369 3429 10379 3496
rect 10480 3496 10537 3501
rect 10480 3362 10483 3496
rect 10529 3362 10537 3496
rect 10158 3266 10215 3362
rect 10323 3351 10369 3362
rect 10480 3266 10537 3362
rect 10722 3496 10779 3503
rect 10722 3362 10727 3496
rect 10773 3362 10779 3496
rect 10876 3496 10943 3504
rect 11047 3501 11093 3507
rect 10876 3429 10887 3496
rect 10933 3429 10943 3496
rect 11044 3496 11101 3501
rect 11044 3362 11047 3496
rect 11093 3362 11101 3496
rect 10722 3266 10779 3362
rect 10887 3351 10933 3362
rect 11044 3266 11101 3362
rect 11257 3271 11343 4208
rect 11404 3677 11476 4454
rect 11771 4166 11880 5139
rect 12025 5038 12079 5139
rect 12574 5050 12625 5054
rect 12188 5038 12234 5049
rect 12348 5038 12394 5049
rect 12507 5038 12625 5050
rect 12025 4932 12028 5038
rect 12074 4932 12079 5038
rect 12507 4932 12508 5038
rect 12554 4932 12625 5038
rect 12025 4926 12079 4932
rect 12028 4921 12074 4926
rect 12188 4921 12234 4932
rect 12348 4921 12394 4932
rect 12507 4920 12625 4932
rect 12749 5038 12803 5139
rect 13298 5050 13349 5054
rect 12912 5038 12958 5049
rect 13072 5038 13118 5049
rect 13231 5038 13349 5050
rect 12749 4932 12752 5038
rect 12798 4932 12803 5038
rect 13231 4932 13232 5038
rect 13278 4932 13349 5038
rect 12749 4926 12803 4932
rect 12752 4921 12798 4926
rect 12912 4921 12958 4932
rect 13072 4921 13118 4932
rect 13231 4920 13349 4932
rect 13473 4994 13527 5139
rect 13473 4932 13476 4994
rect 13522 4932 13527 4994
rect 13473 4926 13527 4932
rect 13625 4994 13694 5005
rect 13796 4995 13842 5005
rect 13625 4932 13636 4994
rect 13682 4932 13694 4994
rect 13476 4921 13522 4926
rect 12054 4809 12135 4821
rect 12574 4816 12625 4920
rect 12574 4810 12728 4816
rect 11971 4807 12135 4809
rect 11971 4804 12072 4807
rect 11971 4750 11984 4804
rect 12038 4757 12072 4804
rect 12121 4757 12135 4807
rect 12038 4750 12135 4757
rect 11971 4742 12135 4750
rect 12054 4741 12135 4742
rect 12182 4797 12728 4810
rect 12778 4807 12859 4821
rect 13298 4816 13349 4920
rect 13625 4919 13694 4932
rect 13790 4994 13845 4995
rect 13790 4932 13796 4994
rect 13842 4932 13845 4994
rect 13298 4810 13456 4816
rect 12778 4797 12796 4807
rect 12182 4761 12796 4797
rect 12028 4604 12074 4608
rect 12182 4605 12234 4761
rect 12280 4714 12360 4715
rect 12280 4712 12379 4714
rect 12280 4709 12292 4712
rect 12280 4661 12291 4709
rect 12280 4660 12292 4661
rect 12344 4660 12379 4712
rect 12280 4657 12379 4660
rect 12427 4709 12528 4715
rect 12427 4661 12438 4709
rect 12427 4657 12439 4661
rect 12491 4658 12528 4709
rect 12491 4657 12503 4658
rect 12574 4610 12625 4761
rect 12682 4757 12796 4761
rect 12845 4757 12859 4807
rect 12682 4750 12859 4757
rect 12778 4741 12859 4750
rect 12906 4797 13456 4810
rect 13502 4807 13583 4821
rect 13790 4816 13845 4932
rect 14037 4994 14091 5139
rect 14037 4932 14040 4994
rect 14086 4932 14091 4994
rect 14037 4926 14091 4932
rect 14189 4994 14258 5005
rect 14360 4995 14406 5005
rect 14189 4932 14200 4994
rect 14246 4932 14258 4994
rect 14040 4921 14086 4926
rect 14189 4919 14258 4932
rect 14354 4994 14409 4995
rect 14354 4932 14360 4994
rect 14406 4932 14409 4994
rect 13790 4810 14013 4816
rect 13502 4797 13520 4807
rect 12906 4761 13520 4797
rect 12023 4597 12080 4604
rect 12023 4463 12028 4597
rect 12074 4463 12080 4597
rect 12177 4597 12244 4605
rect 12348 4602 12394 4608
rect 12177 4530 12188 4597
rect 12234 4530 12244 4597
rect 12345 4597 12402 4602
rect 12345 4463 12348 4597
rect 12394 4463 12402 4597
rect 12023 4367 12080 4463
rect 12188 4452 12234 4463
rect 12345 4367 12402 4463
rect 12506 4597 12625 4610
rect 12752 4604 12798 4608
rect 12906 4605 12958 4761
rect 13151 4709 13252 4715
rect 13151 4661 13162 4709
rect 13151 4657 13163 4661
rect 13215 4658 13252 4709
rect 13215 4657 13227 4658
rect 13298 4610 13349 4761
rect 13410 4757 13520 4761
rect 13569 4757 13583 4807
rect 13410 4750 13583 4757
rect 13502 4741 13583 4750
rect 13630 4797 14013 4810
rect 14066 4807 14147 4821
rect 14354 4816 14409 4932
rect 14066 4797 14084 4807
rect 13630 4761 14084 4797
rect 12506 4463 12508 4597
rect 12554 4463 12625 4597
rect 12506 4445 12625 4463
rect 12747 4597 12804 4604
rect 12747 4463 12752 4597
rect 12798 4463 12804 4597
rect 12747 4367 12804 4463
rect 12901 4597 12968 4605
rect 13072 4602 13118 4608
rect 12901 4514 12912 4597
rect 12901 4462 12905 4514
rect 12958 4463 12968 4597
rect 12957 4462 12968 4463
rect 12901 4450 12968 4462
rect 13069 4597 13126 4602
rect 13069 4463 13072 4597
rect 13118 4463 13126 4597
rect 13069 4367 13126 4463
rect 13230 4597 13349 4610
rect 13476 4604 13522 4608
rect 13630 4605 13682 4761
rect 13957 4757 14084 4761
rect 14133 4757 14147 4807
rect 13957 4750 14147 4757
rect 14066 4741 14147 4750
rect 14194 4815 14524 4816
rect 14194 4763 14208 4815
rect 14260 4763 14524 4815
rect 14194 4761 14524 4763
rect 13750 4714 13830 4715
rect 13750 4709 13904 4714
rect 13750 4661 13765 4709
rect 13750 4657 13766 4661
rect 13818 4657 13904 4709
rect 13230 4463 13232 4597
rect 13278 4463 13349 4597
rect 13230 4445 13349 4463
rect 13471 4597 13528 4604
rect 13471 4463 13476 4597
rect 13522 4463 13528 4597
rect 13625 4597 13692 4605
rect 13796 4602 13842 4608
rect 14040 4604 14086 4608
rect 14194 4605 14246 4761
rect 14314 4714 14394 4715
rect 14314 4661 14329 4714
rect 14381 4662 14468 4714
rect 14377 4661 14468 4662
rect 14314 4657 14468 4661
rect 13625 4530 13636 4597
rect 13682 4530 13692 4597
rect 13793 4597 13850 4602
rect 13793 4463 13796 4597
rect 13842 4463 13850 4597
rect 13471 4367 13528 4463
rect 13636 4452 13682 4463
rect 13793 4367 13850 4463
rect 14035 4597 14092 4604
rect 14035 4463 14040 4597
rect 14086 4463 14092 4597
rect 14189 4597 14256 4605
rect 14360 4602 14406 4608
rect 14189 4530 14200 4597
rect 14246 4530 14256 4597
rect 14357 4597 14414 4602
rect 14357 4463 14360 4597
rect 14406 4463 14414 4597
rect 14035 4367 14092 4463
rect 14200 4452 14246 4463
rect 14357 4367 14414 4463
rect 11927 4347 14536 4367
rect 11927 4301 12076 4347
rect 12303 4301 12800 4347
rect 13027 4301 13524 4347
rect 13751 4301 14088 4347
rect 14315 4301 14536 4347
rect 11927 4212 14536 4301
rect 11771 4160 14342 4166
rect 11771 4019 14343 4160
rect 11771 3980 11935 4019
rect 11531 3946 11935 3980
rect 11531 3900 11582 3946
rect 11872 3900 11935 3946
rect 11531 3874 11935 3900
rect 12031 3941 12085 4019
rect 12580 3953 12631 3957
rect 12194 3941 12240 3952
rect 12354 3941 12400 3952
rect 12513 3941 12631 3953
rect 11615 3791 11682 3874
rect 12031 3835 12034 3941
rect 12080 3835 12085 3941
rect 12513 3835 12514 3941
rect 12560 3835 12631 3941
rect 12031 3829 12085 3835
rect 12034 3824 12080 3829
rect 12194 3824 12240 3835
rect 12354 3824 12400 3835
rect 12513 3823 12631 3835
rect 12755 3897 12809 4019
rect 12755 3835 12758 3897
rect 12804 3835 12809 3897
rect 12755 3829 12809 3835
rect 12907 3897 12976 3908
rect 13078 3898 13124 3908
rect 12907 3835 12918 3897
rect 12964 3835 12976 3897
rect 12758 3824 12804 3829
rect 11615 3745 11626 3791
rect 11672 3745 11683 3791
rect 11783 3745 11794 3791
rect 11840 3745 11851 3791
rect 11404 3664 11742 3677
rect 11404 3663 11680 3664
rect 11404 3611 11678 3663
rect 11736 3618 11742 3664
rect 11730 3611 11742 3618
rect 11404 3605 11742 3611
rect 11788 3674 11851 3745
rect 12005 3724 12091 3725
rect 12005 3722 12141 3724
rect 11788 3616 11935 3674
rect 12005 3670 12018 3722
rect 12081 3710 12141 3722
rect 12580 3719 12631 3823
rect 12907 3822 12976 3835
rect 13072 3897 13127 3898
rect 13072 3835 13078 3897
rect 13124 3835 13127 3897
rect 12580 3713 12737 3719
rect 12005 3660 12078 3670
rect 12127 3660 12141 3710
rect 12005 3651 12141 3660
rect 12060 3644 12141 3651
rect 12188 3700 12737 3713
rect 12784 3710 12865 3724
rect 13072 3719 13127 3835
rect 13319 3897 13373 4019
rect 13319 3835 13322 3897
rect 13368 3835 13373 3897
rect 13319 3829 13373 3835
rect 13471 3897 13540 3908
rect 13642 3898 13688 3908
rect 13471 3835 13482 3897
rect 13528 3835 13540 3897
rect 13322 3824 13368 3829
rect 13471 3822 13540 3835
rect 13636 3897 13691 3898
rect 13636 3835 13642 3897
rect 13688 3835 13691 3897
rect 13072 3713 13195 3719
rect 12784 3700 12802 3710
rect 12188 3664 12802 3700
rect 11617 3500 11680 3513
rect 11617 3366 11630 3500
rect 11676 3366 11680 3500
rect 11617 3280 11680 3366
rect 11788 3500 11851 3616
rect 12034 3507 12080 3511
rect 12188 3508 12240 3664
rect 12286 3617 12366 3618
rect 12286 3612 12385 3617
rect 12286 3564 12297 3612
rect 12286 3560 12298 3564
rect 12350 3560 12385 3612
rect 12433 3612 12456 3618
rect 12433 3564 12444 3612
rect 12508 3566 12534 3618
rect 12492 3564 12534 3566
rect 12433 3560 12534 3564
rect 12580 3513 12631 3664
rect 12691 3660 12802 3664
rect 12851 3660 12865 3710
rect 12691 3653 12865 3660
rect 12784 3644 12865 3653
rect 12912 3667 13195 3713
rect 13247 3700 13302 3719
rect 13348 3710 13429 3724
rect 13636 3719 13691 3835
rect 13883 3897 13937 4019
rect 13883 3835 13886 3897
rect 13932 3835 13937 3897
rect 13883 3829 13937 3835
rect 14035 3897 14104 3908
rect 14206 3898 14252 3908
rect 14035 3835 14046 3897
rect 14092 3835 14104 3897
rect 13886 3824 13932 3829
rect 14035 3822 14104 3835
rect 14200 3897 14255 3898
rect 14200 3835 14206 3897
rect 14252 3835 14255 3897
rect 14200 3728 14255 3835
rect 14200 3727 14370 3728
rect 13636 3713 13861 3719
rect 13348 3700 13366 3710
rect 13247 3667 13366 3700
rect 12912 3664 13366 3667
rect 11788 3483 11790 3500
rect 11836 3483 11851 3500
rect 11788 3431 11789 3483
rect 11841 3431 11851 3483
rect 11788 3366 11790 3431
rect 11836 3366 11851 3431
rect 11788 3355 11851 3366
rect 12029 3500 12086 3507
rect 12029 3366 12034 3500
rect 12080 3366 12086 3500
rect 12183 3500 12250 3508
rect 12354 3505 12400 3511
rect 12183 3433 12194 3500
rect 12240 3433 12250 3500
rect 12351 3500 12408 3505
rect 12351 3366 12354 3500
rect 12400 3366 12408 3500
rect 11257 3270 11408 3271
rect 11531 3270 11935 3280
rect 12029 3270 12086 3366
rect 12194 3355 12240 3366
rect 12351 3270 12408 3366
rect 12512 3500 12631 3513
rect 12758 3507 12804 3511
rect 12912 3508 12964 3664
rect 13240 3660 13366 3664
rect 13415 3660 13429 3710
rect 13240 3653 13429 3660
rect 13348 3644 13429 3653
rect 13476 3700 13861 3713
rect 13912 3710 13993 3724
rect 14200 3713 14266 3727
rect 13912 3700 13930 3710
rect 13476 3664 13930 3700
rect 13032 3617 13112 3618
rect 13032 3612 13186 3617
rect 13032 3564 13047 3612
rect 13032 3560 13048 3564
rect 13100 3560 13186 3612
rect 12512 3366 12514 3500
rect 12560 3366 12631 3500
rect 12512 3348 12631 3366
rect 12753 3500 12810 3507
rect 12753 3366 12758 3500
rect 12804 3366 12810 3500
rect 12907 3500 12974 3508
rect 13078 3505 13124 3511
rect 13322 3507 13368 3511
rect 13476 3508 13528 3664
rect 13805 3660 13930 3664
rect 13979 3660 13993 3710
rect 13805 3653 13993 3660
rect 13912 3644 13993 3653
rect 14040 3675 14266 3713
rect 14318 3675 14370 3727
rect 14040 3664 14370 3675
rect 13596 3617 13676 3618
rect 13596 3612 13750 3617
rect 13596 3564 13611 3612
rect 13596 3560 13612 3564
rect 13664 3560 13750 3612
rect 12907 3433 12918 3500
rect 12964 3433 12974 3500
rect 13075 3500 13132 3505
rect 13075 3366 13078 3500
rect 13124 3366 13132 3500
rect 12753 3270 12810 3366
rect 12918 3355 12964 3366
rect 13075 3270 13132 3366
rect 13317 3500 13374 3507
rect 13317 3366 13322 3500
rect 13368 3366 13374 3500
rect 13471 3500 13538 3508
rect 13642 3505 13688 3511
rect 13886 3507 13932 3511
rect 14040 3508 14092 3664
rect 14160 3617 14240 3618
rect 14160 3615 14314 3617
rect 14160 3563 14172 3615
rect 14224 3563 14314 3615
rect 14160 3560 14314 3563
rect 13471 3433 13482 3500
rect 13528 3433 13538 3500
rect 13639 3500 13696 3505
rect 13639 3366 13642 3500
rect 13688 3366 13696 3500
rect 13317 3270 13374 3366
rect 13482 3355 13528 3366
rect 13639 3270 13696 3366
rect 13881 3500 13938 3507
rect 13881 3366 13886 3500
rect 13932 3366 13938 3500
rect 14035 3500 14102 3508
rect 14206 3505 14252 3511
rect 14035 3433 14046 3500
rect 14092 3433 14102 3500
rect 14203 3500 14260 3505
rect 14203 3366 14206 3500
rect 14252 3366 14260 3500
rect 13881 3270 13938 3366
rect 14046 3355 14092 3366
rect 14203 3270 14260 3366
rect 14416 3270 14536 4212
rect 11257 3267 14536 3270
rect 11257 3266 11584 3267
rect 8372 3263 11584 3266
rect 8372 3256 8425 3263
rect 5605 3248 8425 3256
rect 5605 3209 5809 3248
rect 4753 3202 5809 3209
rect 6036 3202 6533 3248
rect 6760 3202 7097 3248
rect 7324 3202 7661 3248
rect 7888 3207 8425 3248
rect 8719 3246 11584 3263
rect 8719 3207 8923 3246
rect 7888 3202 8923 3207
rect 4753 3201 8923 3202
rect 4753 3200 5970 3201
rect 101 3180 201 3184
rect 101 3127 136 3180
rect 189 3127 201 3180
rect 2123 3170 5970 3200
rect 101 3123 201 3127
rect 2525 3117 5970 3170
rect 6033 3200 8923 3201
rect 9150 3200 9647 3246
rect 9874 3200 10211 3246
rect 10438 3200 10775 3246
rect 11002 3211 11584 3246
rect 11878 3250 14536 3267
rect 11878 3211 12082 3250
rect 11002 3204 12082 3211
rect 12309 3204 12806 3250
rect 13033 3204 13370 3250
rect 13597 3204 13934 3250
rect 14161 3204 14536 3250
rect 11002 3200 14536 3204
rect 6033 3117 14536 3200
rect 873 3088 1020 3102
rect 2525 3089 14536 3117
rect -403 3041 -131 3088
rect -403 2579 -314 3041
rect 440 3002 620 3077
rect 873 3019 900 3088
rect 1003 3019 1020 3088
rect 11268 3038 11374 3040
rect 873 3005 1020 3019
rect 2915 3023 11374 3038
rect 2915 2944 2929 3023
rect 3008 3021 11374 3023
rect 3008 2944 11284 3021
rect 2915 2930 11284 2944
rect 11352 2930 11374 3021
rect 2915 2927 11374 2930
rect 11268 2912 11374 2927
rect 1528 2889 1655 2893
rect 1528 2836 1543 2889
rect 1622 2836 1655 2889
rect 1528 2832 1655 2836
rect 2105 2848 5347 2869
rect 516 2684 621 2806
rect 1211 2786 1321 2798
rect 1211 2781 1234 2786
rect -403 2512 -372 2579
rect -319 2512 -314 2579
rect 196 2575 621 2684
rect 1091 2735 1234 2781
rect -403 2024 -314 2512
rect 296 2475 395 2575
rect 1091 2515 1137 2735
rect 1211 2727 1234 2735
rect 1297 2727 1321 2786
rect 2105 2780 5238 2848
rect 5316 2780 5347 2848
rect 2105 2754 5347 2780
rect 5471 2854 14428 2866
rect 5471 2850 14343 2854
rect 5471 2770 5488 2850
rect 5557 2836 14343 2850
rect 5557 2784 7614 2836
rect 7669 2790 14343 2836
rect 14411 2790 14428 2854
rect 7669 2784 14428 2790
rect 5557 2770 14428 2784
rect 5471 2751 14428 2770
rect 1211 2715 1321 2727
rect 11464 2687 11582 2702
rect 8687 2681 11582 2687
rect 8687 2673 11484 2681
rect 2194 2661 2316 2669
rect 8429 2661 8550 2662
rect 2193 2647 8550 2661
rect 2193 2552 2214 2647
rect 2283 2627 8550 2647
rect 2283 2571 8457 2627
rect 8525 2571 8550 2627
rect 8687 2615 8702 2673
rect 8769 2615 11484 2673
rect 8687 2586 11484 2615
rect 11567 2586 11582 2681
rect 2283 2552 8550 2571
rect 11464 2570 11582 2586
rect 2193 2540 8550 2552
rect 2194 2527 2316 2540
rect 8422 2537 8550 2540
rect 1008 2465 1137 2515
rect -265 2409 -156 2427
rect -265 2336 -253 2409
rect -174 2336 -156 2409
rect -265 2318 -156 2336
rect -403 1977 -138 2024
rect 747 1998 875 2007
rect 653 1990 875 1998
rect -572 1928 -485 1940
rect -572 1874 -551 1928
rect -497 1874 -485 1928
rect -572 1868 -485 1874
rect -565 1863 -485 1868
rect -403 1640 -314 1977
rect 118 1938 243 1942
rect 653 1940 776 1990
rect 118 1886 146 1938
rect 222 1886 243 1938
rect 747 1919 776 1940
rect 856 1919 875 1990
rect 747 1893 875 1919
rect 1008 1981 1054 2465
rect 2459 2458 5100 2469
rect 2457 2449 5100 2458
rect 1182 2383 1666 2384
rect 1155 2288 2114 2383
rect 2457 2381 2469 2449
rect 2526 2448 5100 2449
rect 2526 2387 5034 2448
rect 5087 2387 5100 2448
rect 2526 2381 5100 2387
rect 2457 2373 5100 2381
rect 2459 2366 5100 2373
rect 5760 2440 11223 2469
rect 5760 2435 11150 2440
rect 5760 2376 5782 2435
rect 5855 2434 11150 2435
rect 5855 2376 8455 2434
rect 5760 2372 8455 2376
rect 8509 2372 11150 2434
rect 5760 2366 11150 2372
rect 5763 2364 11150 2366
rect 11211 2364 11223 2440
rect 5763 2363 11223 2364
rect 5763 2359 5877 2363
rect 11139 2353 11223 2363
rect 1155 2275 2680 2288
rect 3693 2275 8780 2302
rect 1155 2222 1159 2275
rect 1214 2222 2680 2275
rect 3687 2274 8780 2275
rect 1155 2195 2680 2222
rect 2065 2169 2680 2195
rect 3686 2269 8780 2274
rect 3686 2259 8708 2269
rect 3686 2190 3701 2259
rect 3768 2217 8708 2259
rect 8766 2217 8780 2269
rect 3768 2201 8780 2217
rect 10530 2287 10750 2291
rect 14636 2287 15022 5139
rect 10530 2280 15022 2287
rect 10530 2217 10552 2280
rect 10604 2217 10664 2280
rect 10716 2217 15022 2280
rect 3768 2190 3789 2201
rect 3686 2181 3789 2190
rect 10530 2155 15022 2217
rect 5027 2150 5112 2153
rect 8113 2150 8194 2151
rect 3841 2140 8196 2150
rect 3841 2134 5043 2140
rect 3841 2069 3858 2134
rect 3917 2070 5043 2134
rect 5099 2139 8196 2140
rect 5099 2070 8131 2139
rect 3917 2069 8131 2070
rect 3841 2067 8131 2069
rect 8187 2067 8196 2139
rect 10530 2103 10590 2155
rect 10679 2103 15022 2155
rect 10530 2100 15022 2103
rect 10532 2069 15022 2100
rect 3841 2047 8196 2067
rect 2161 1993 2283 2015
rect 1008 1935 1343 1981
rect 2161 1958 2189 1993
rect 118 1883 243 1886
rect -403 1630 -309 1640
rect -403 1629 -368 1630
rect -403 1556 -370 1629
rect -315 1556 -309 1630
rect -403 1548 -309 1556
rect -383 1544 -309 1548
rect 1008 1486 1054 1935
rect 1462 1908 1555 1917
rect 1462 1853 1476 1908
rect 1537 1853 1555 1908
rect 2031 1900 2189 1958
rect 2161 1898 2189 1900
rect 2258 1898 2283 1993
rect 2456 1986 2758 1994
rect 2456 1934 2467 1986
rect 2526 1934 2758 1986
rect 3689 1961 3771 1969
rect 2456 1916 2758 1934
rect 3529 1960 3771 1961
rect 2161 1873 2283 1898
rect 2929 1912 3012 1918
rect 1462 1845 1555 1853
rect 2929 1860 2943 1912
rect 3001 1860 3012 1912
rect 3529 1908 3697 1960
rect 3759 1908 3771 1960
rect 3529 1903 3771 1908
rect 3689 1896 3771 1903
rect 4005 1960 4119 1964
rect 5763 1960 5877 1966
rect 4005 1952 5877 1960
rect 4005 1886 4018 1952
rect 4103 1950 5877 1952
rect 4103 1888 5782 1950
rect 5862 1888 5877 1950
rect 4103 1886 5877 1888
rect 4005 1878 5877 1886
rect 4005 1871 4119 1878
rect 5763 1872 5877 1878
rect 2929 1846 3012 1860
rect 1462 1844 1554 1845
rect 6096 1841 8801 1989
rect 10802 1961 10870 1964
rect 9016 1952 10870 1961
rect 9016 1900 9024 1952
rect 9082 1951 10870 1952
rect 9082 1900 10807 1951
rect 9016 1899 10807 1900
rect 10865 1899 10870 1951
rect 9016 1892 10870 1899
rect 9016 1887 9096 1892
rect 10802 1886 10870 1892
rect 4219 1799 5576 1811
rect 11464 1807 11640 1876
rect 4219 1741 4230 1799
rect 4286 1795 5576 1799
rect 4286 1741 5479 1795
rect 4219 1731 5479 1741
rect 4220 1729 5479 1731
rect 5454 1726 5479 1729
rect 5561 1726 5576 1795
rect 9066 1775 10671 1785
rect 5454 1709 5576 1726
rect 9058 1689 10671 1775
rect 5018 1652 5101 1664
rect 5018 1583 5026 1652
rect 5088 1649 5101 1652
rect 5088 1583 6192 1649
rect 7008 1588 7166 1646
rect 9058 1628 10596 1689
rect 10657 1628 10671 1689
rect 9058 1610 10671 1628
rect 9066 1609 10671 1610
rect 10755 1740 11010 1803
rect 9090 1605 10669 1609
rect 5018 1577 6192 1583
rect 5018 1565 5101 1577
rect 7108 1493 7166 1588
rect 1005 1485 1080 1486
rect 1004 1478 1080 1485
rect -259 1345 -160 1454
rect 1004 1412 1013 1478
rect 1065 1412 1080 1478
rect 1004 1401 1080 1412
rect 7108 1446 7375 1493
rect 7927 1457 8052 1512
rect 8990 1464 9098 1480
rect 7108 1370 7166 1446
rect 7103 1359 7185 1370
rect -260 1328 6112 1345
rect -260 1244 5972 1328
rect 6035 1244 6112 1328
rect 7103 1306 7117 1359
rect 7169 1306 7185 1359
rect 7103 1293 7185 1306
rect -260 1146 6112 1244
rect -260 1117 7071 1146
rect 7997 1129 8052 1457
rect 8990 1412 9018 1464
rect 9080 1412 9098 1464
rect 10755 1414 10818 1740
rect 8990 1401 9098 1412
rect 9159 1339 9364 1411
rect 10562 1351 10818 1414
rect 11571 1411 11640 1807
rect 11714 1699 11773 2069
rect 11714 1655 11765 1699
rect 11571 1339 11790 1411
rect 12060 1350 12227 1408
rect 9159 1146 9231 1339
rect 9148 1134 9232 1146
rect -274 1063 7071 1117
rect 7993 1117 8065 1129
rect 7993 1063 8005 1117
rect 8058 1063 8065 1117
rect -274 977 7247 1063
rect 7993 1051 8065 1063
rect 9148 1066 9161 1134
rect 9221 1066 9232 1134
rect 9148 1046 9232 1066
rect 10916 1018 11443 1139
rect 10916 1013 11754 1018
rect 10648 977 11754 1013
rect -274 838 12117 977
rect 6985 763 12117 838
<< via1 >>
rect 1879 5188 1939 5242
rect 3611 5333 3664 5386
rect 118 4995 203 5082
rect 2148 4986 2210 5073
rect 292 4798 353 4862
rect 1723 4782 1784 4858
rect 2144 4737 2206 4811
rect -377 4171 -318 4227
rect -114 4167 -58 4222
rect -552 4014 -498 4078
rect -732 2331 -653 2404
rect 856 4163 912 4215
rect 140 4071 192 4123
rect 582 4099 634 4151
rect 1034 4098 1086 4150
rect 2576 4746 2630 4800
rect 2884 4656 2936 4708
rect 3031 4653 3083 4705
rect 3611 4655 3666 4707
rect 3755 4653 3807 4705
rect 3497 4458 3549 4510
rect 4800 4759 4852 4811
rect 5045 4759 5100 4811
rect 4358 4653 4410 4705
rect 4921 4658 4973 4710
rect 5169 4464 5241 4547
rect 1879 3609 1939 3663
rect 2270 3607 2322 3659
rect 2610 3666 2673 3718
rect 2890 3556 2942 3608
rect 3048 3562 3100 3614
rect 3787 3663 3839 3715
rect 2381 3427 2433 3479
rect 3640 3556 3692 3608
rect 4858 3671 4910 3723
rect 4204 3556 4256 3608
rect 4764 3559 4816 3611
rect 5711 4748 5765 4802
rect 6019 4658 6071 4710
rect 6166 4655 6218 4707
rect 6753 4657 6807 4711
rect 6890 4655 6942 4707
rect 6632 4460 6684 4512
rect 7935 4761 7987 4813
rect 7493 4655 7545 4707
rect 8056 4660 8108 4712
rect 5405 3609 5457 3661
rect 5745 3668 5808 3720
rect 6025 3558 6077 3610
rect 6183 3564 6235 3616
rect 6922 3665 6974 3717
rect 5516 3429 5568 3481
rect 6775 3558 6827 3610
rect 7993 3673 8045 3725
rect 7339 3558 7391 3610
rect 7899 3561 7951 3613
rect 8825 4746 8879 4800
rect 9133 4656 9185 4708
rect 9280 4653 9332 4705
rect 9866 4655 9920 4708
rect 10004 4653 10056 4705
rect 9746 4458 9798 4510
rect 11049 4759 11101 4811
rect 11594 4757 11651 4810
rect 10607 4653 10659 4705
rect 11170 4658 11222 4710
rect 11395 4480 11456 4544
rect 8289 3612 8343 3665
rect 8519 3607 8571 3659
rect 8859 3666 8922 3718
rect 9139 3556 9191 3608
rect 9297 3562 9349 3614
rect 10036 3663 10088 3715
rect 8630 3427 8682 3479
rect 9889 3556 9941 3608
rect 11107 3671 11159 3723
rect 10453 3556 10505 3608
rect 11013 3559 11065 3611
rect 11984 4750 12038 4804
rect 12292 4660 12344 4712
rect 12439 4657 12491 4709
rect 13018 4661 13079 4713
rect 13163 4657 13215 4709
rect 12905 4462 12957 4514
rect 14208 4763 14260 4815
rect 13766 4657 13818 4709
rect 14329 4662 14381 4714
rect 11678 3611 11730 3663
rect 12018 3670 12081 3722
rect 12298 3560 12350 3612
rect 12456 3566 12508 3618
rect 13195 3667 13247 3719
rect 11789 3431 11841 3483
rect 13048 3560 13100 3612
rect 14266 3675 14318 3727
rect 13612 3560 13664 3612
rect 14172 3563 14224 3615
rect 136 3127 189 3180
rect 271 3127 335 3179
rect 5970 3117 6033 3201
rect 900 3019 1003 3088
rect 2929 2944 3008 3023
rect 11284 2930 11352 3021
rect 1543 2836 1622 2889
rect -372 2512 -319 2579
rect 1234 2727 1297 2786
rect 5238 2780 5316 2848
rect 5488 2770 5557 2850
rect 7614 2784 7669 2836
rect 14343 2790 14411 2854
rect 2214 2552 2283 2647
rect 8457 2571 8525 2627
rect 8702 2615 8769 2673
rect 11484 2586 11567 2681
rect -253 2336 -174 2409
rect 649 2223 704 2276
rect -551 1874 -497 1928
rect 146 1886 222 1938
rect 776 1919 856 1990
rect 2469 2381 2526 2449
rect 5034 2387 5087 2448
rect 5782 2376 5855 2435
rect 8455 2372 8509 2434
rect 11150 2364 11211 2440
rect 1159 2222 1214 2275
rect 3701 2190 3768 2259
rect 8708 2217 8766 2269
rect 10552 2217 10604 2280
rect 10664 2217 10716 2280
rect 3858 2069 3917 2134
rect 5043 2070 5099 2140
rect 8131 2067 8187 2139
rect 10590 2103 10679 2155
rect -368 1629 -315 1630
rect -370 1556 -315 1629
rect 1476 1853 1537 1908
rect 2189 1898 2258 1993
rect 2467 1934 2526 1986
rect 2943 1860 3001 1912
rect 3697 1908 3759 1960
rect 4018 1886 4103 1952
rect 5782 1888 5862 1950
rect 9024 1900 9082 1952
rect 10807 1899 10865 1951
rect 4230 1741 4286 1799
rect 5479 1726 5561 1795
rect 5026 1583 5088 1652
rect 10596 1628 10657 1689
rect 1013 1412 1065 1478
rect 8256 1457 8309 1509
rect 5972 1244 6035 1328
rect 7117 1306 7169 1359
rect 7613 1354 7668 1406
rect 7762 1356 7832 1408
rect 9018 1412 9080 1464
rect 11175 1739 11229 1791
rect 11323 1738 11376 1790
rect 8501 1357 8560 1410
rect 8005 1063 8058 1117
rect 9161 1066 9221 1134
<< metal2 >>
rect 3595 5394 3676 5401
rect 3595 5327 3606 5394
rect 3667 5327 3676 5394
rect 3595 5305 3676 5327
rect 1868 5242 1955 5259
rect 1868 5188 1879 5242
rect 1939 5188 1955 5242
rect 88 5082 225 5104
rect 88 4995 118 5082
rect 203 4995 225 5082
rect 88 4971 225 4995
rect -387 4227 -306 4239
rect -387 4171 -377 4227
rect -318 4225 -306 4227
rect -124 4225 -54 4234
rect -318 4222 -54 4225
rect -318 4171 -114 4222
rect -387 4169 -114 4171
rect -387 4156 -306 4169
rect -124 4167 -114 4169
rect -58 4167 -54 4222
rect -124 4155 -54 4167
rect 133 4135 194 4971
rect 280 4862 369 4875
rect 280 4798 292 4862
rect 353 4798 369 4862
rect 280 4785 369 4798
rect 1713 4858 1797 4875
rect 127 4123 196 4135
rect -566 4078 -483 4087
rect -566 4014 -552 4078
rect -498 4071 -483 4078
rect 127 4071 140 4123
rect 192 4071 196 4123
rect -498 4014 195 4071
rect -566 4010 195 4014
rect -566 3998 -483 4010
rect 285 3191 365 4785
rect 1713 4782 1723 4858
rect 1784 4782 1797 4858
rect 1713 4767 1797 4782
rect 1024 4352 1095 4370
rect 579 4281 1095 4352
rect 579 4155 650 4281
rect 570 4151 650 4155
rect 570 4099 582 4151
rect 634 4099 650 4151
rect 839 4215 922 4224
rect 839 4163 856 4215
rect 912 4163 922 4215
rect 839 4147 922 4163
rect 1024 4155 1095 4281
rect 570 4092 650 4099
rect 100 3180 201 3182
rect 100 3127 136 3180
rect 189 3127 201 3180
rect 100 3123 201 3127
rect 257 3179 365 3191
rect 257 3127 271 3179
rect 335 3127 365 3179
rect 100 2786 171 3123
rect 257 3115 365 3127
rect 843 3102 922 4147
rect 1019 4150 1099 4155
rect 1019 4098 1034 4150
rect 1086 4098 1099 4150
rect 1019 4092 1099 4098
rect 1019 4091 1092 4092
rect 843 3088 1020 3102
rect 843 3019 900 3088
rect 1003 3019 1020 3088
rect 843 3005 1020 3019
rect 1528 2889 1655 2894
rect 1528 2836 1543 2889
rect 1622 2836 1655 2889
rect 1528 2832 1655 2836
rect 1211 2786 1321 2798
rect 100 2727 1234 2786
rect 1297 2727 1321 2786
rect 100 2715 1321 2727
rect -386 2584 -314 2594
rect 1535 2584 1616 2832
rect -386 2579 1616 2584
rect -386 2512 -372 2579
rect -319 2512 1616 2579
rect -386 2503 1616 2512
rect -386 2500 -314 2503
rect -750 2407 -629 2417
rect -265 2409 -156 2427
rect -265 2407 -253 2409
rect -750 2404 -253 2407
rect -750 2331 -732 2404
rect -653 2336 -253 2404
rect -174 2336 -156 2409
rect -653 2331 -156 2336
rect -750 2326 -156 2331
rect -750 2321 -629 2326
rect -265 2318 -156 2326
rect 618 2276 1223 2285
rect 618 2223 649 2276
rect 704 2275 1223 2276
rect 704 2223 1159 2275
rect 618 2222 1159 2223
rect 1214 2222 1223 2275
rect 618 2208 1223 2222
rect 747 1990 875 2007
rect -565 1935 -485 1940
rect 116 1938 241 1943
rect 116 1935 146 1938
rect -565 1928 146 1935
rect -565 1874 -551 1928
rect -497 1886 146 1928
rect 222 1935 241 1938
rect 222 1886 242 1935
rect 747 1919 776 1990
rect 856 1919 875 1990
rect 747 1916 875 1919
rect 1462 1916 1555 1917
rect 747 1908 1558 1916
rect 747 1893 1476 1908
rect -497 1874 242 1886
rect -565 1868 242 1874
rect -565 1863 -485 1868
rect 760 1853 1476 1893
rect 1537 1853 1558 1908
rect 760 1842 1558 1853
rect 1719 1774 1792 4767
rect 1868 3663 1955 5188
rect 2127 5073 2221 5091
rect 2127 4986 2148 5073
rect 2210 5049 2221 5073
rect 2210 4991 4976 5049
rect 2210 4986 2221 4991
rect 2127 4970 2221 4986
rect 2135 4811 2218 4820
rect 2135 4737 2144 4811
rect 2206 4810 2218 4811
rect 2206 4805 2624 4810
rect 2206 4800 2642 4805
rect 2206 4746 2576 4800
rect 2630 4746 2642 4800
rect 2206 4738 2642 4746
rect 2206 4737 2629 4738
rect 2135 4730 2629 4737
rect 2135 4725 2218 4730
rect 2244 4545 2342 4563
rect 2244 4471 2260 4545
rect 2325 4471 2342 4545
rect 2244 4453 2342 4471
rect 1868 3609 1879 3663
rect 1939 3609 1955 3663
rect 1868 3601 1955 3609
rect 2268 3659 2325 4453
rect 2268 3607 2270 3659
rect 2322 3607 2325 3659
rect 2571 3721 2629 4730
rect 2879 4708 2938 4720
rect 2879 4656 2884 4708
rect 2936 4656 2938 4708
rect 2879 4641 2938 4656
rect 3018 4708 3075 4991
rect 3177 4878 4854 4934
rect 3018 4705 3118 4708
rect 3018 4653 3031 4705
rect 3083 4653 3118 4705
rect 3019 4650 3118 4653
rect 2571 3718 2685 3721
rect 2571 3666 2610 3718
rect 2673 3666 2685 3718
rect 2571 3658 2685 3666
rect 2602 3657 2685 3658
rect 2879 3611 2935 4641
rect 3177 3617 3233 4878
rect 4798 4811 4854 4878
rect 4798 4771 4800 4811
rect 4734 4759 4800 4771
rect 4852 4759 4854 4811
rect 3595 4722 3686 4731
rect 3595 4649 3604 4722
rect 3678 4649 3686 4722
rect 4734 4715 4854 4759
rect 4192 4708 4346 4709
rect 3743 4705 3842 4708
rect 3743 4653 3755 4705
rect 3807 4653 3842 4705
rect 3743 4650 3842 4653
rect 3595 4634 3686 4649
rect 3036 3614 3233 3617
rect 2268 3595 2325 3607
rect 2878 3608 2954 3611
rect 2878 3595 2890 3608
rect 2268 3556 2890 3595
rect 2942 3556 2954 3608
rect 3036 3562 3048 3614
rect 3100 3562 3233 3614
rect 3036 3561 3233 3562
rect 3493 4510 3551 4522
rect 3493 4458 3497 4510
rect 3549 4458 3551 4510
rect 3493 3610 3551 4458
rect 3786 3717 3842 4650
rect 3785 3715 3842 3717
rect 3785 3663 3787 3715
rect 3839 3663 3842 3715
rect 3785 3659 3842 3663
rect 3786 3651 3842 3659
rect 4192 4705 4445 4708
rect 4192 4653 4358 4705
rect 4410 4653 4445 4705
rect 4192 4650 4445 4653
rect 4192 3611 4248 4650
rect 4734 3613 4790 4715
rect 4918 4710 4976 4991
rect 6153 4993 8111 5051
rect 4918 4658 4921 4710
rect 4973 4658 4976 4710
rect 4867 4602 4976 4658
rect 5032 4811 5117 4828
rect 5032 4759 5045 4811
rect 5100 4759 5117 4811
rect 5032 4757 5117 4759
rect 5698 4802 5777 4807
rect 4867 3820 4923 4602
rect 4867 3745 4953 3820
rect 4846 3723 4953 3745
rect 4846 3671 4858 3723
rect 4910 3671 4953 3723
rect 4846 3668 4953 3671
rect 4734 3611 4829 3613
rect 3493 3608 3704 3610
rect 3036 3560 3102 3561
rect 2268 3547 2954 3556
rect 3493 3556 3640 3608
rect 3692 3556 3704 3608
rect 3493 3553 3704 3556
rect 4192 3608 4291 3611
rect 4192 3556 4204 3608
rect 4256 3556 4291 3608
rect 4734 3559 4764 3611
rect 4816 3559 4829 3611
rect 4734 3557 4829 3559
rect 4192 3553 4291 3556
rect 2268 3545 2942 3547
rect 2268 3538 2934 3545
rect 4192 3482 4248 3553
rect 2369 3479 4248 3482
rect 2369 3427 2381 3479
rect 2433 3427 4248 3479
rect 2369 3426 4248 3427
rect 4897 3549 4953 3668
rect 2379 3425 2435 3426
rect 4897 3263 4954 3549
rect 2905 3023 3030 3057
rect 2905 2944 2929 3023
rect 3008 2944 3030 3023
rect 2905 2927 3030 2944
rect 2194 2647 2316 2669
rect 2194 2552 2214 2647
rect 2283 2552 2316 2647
rect 2194 2527 2316 2552
rect 2197 2015 2255 2527
rect 2457 2449 2537 2458
rect 2457 2381 2469 2449
rect 2526 2381 2537 2449
rect 2457 2373 2537 2381
rect 2161 1993 2283 2015
rect 2457 1994 2536 2373
rect 2161 1898 2189 1993
rect 2258 1898 2283 1993
rect 2456 1986 2539 1994
rect 2456 1934 2467 1986
rect 2526 1934 2539 1986
rect 2456 1916 2539 1934
rect 2929 1921 3007 2927
rect 3686 2259 3789 2274
rect 3686 2190 3701 2259
rect 3768 2190 3789 2259
rect 3686 2181 3789 2190
rect 3691 1969 3767 2181
rect 3846 2141 3938 2149
rect 3845 2134 3938 2141
rect 3845 2069 3858 2134
rect 3917 2069 3938 2134
rect 3845 2052 3938 2069
rect 3689 1960 3771 1969
rect 2161 1873 2283 1898
rect 2929 1912 3012 1921
rect 2929 1860 2943 1912
rect 3001 1860 3012 1912
rect 3689 1908 3697 1960
rect 3759 1908 3771 1960
rect 3689 1896 3771 1908
rect 2929 1846 3012 1860
rect 3845 1774 3918 2052
rect 4005 1952 4119 1964
rect 4005 1886 4018 1952
rect 4103 1886 4119 1952
rect 4005 1871 4119 1886
rect 1719 1701 3918 1774
rect -383 1638 -309 1640
rect 4007 1638 4100 1871
rect 4219 1799 4295 1811
rect 4219 1741 4230 1799
rect 4286 1741 4295 1799
rect 4219 1731 4295 1741
rect -383 1630 4100 1638
rect -383 1629 -368 1630
rect -383 1556 -370 1629
rect -315 1556 4100 1630
rect -383 1545 4100 1556
rect -383 1544 -309 1545
rect 4220 1486 4293 1731
rect 1005 1485 4293 1486
rect 1004 1478 4293 1485
rect 1004 1412 1013 1478
rect 1065 1413 4293 1478
rect 1065 1412 1080 1413
rect 1004 1401 1080 1412
rect 4830 960 4954 3263
rect 5032 2457 5094 4757
rect 5698 4748 5711 4802
rect 5765 4748 5777 4802
rect 5698 4740 5777 4748
rect 5152 4556 5262 4563
rect 5152 4462 5162 4556
rect 5251 4462 5262 4556
rect 5152 4453 5262 4462
rect 5706 4213 5764 4740
rect 5249 4155 5764 4213
rect 5249 2931 5307 4155
rect 5706 3723 5764 4155
rect 6014 4710 6073 4722
rect 6014 4658 6019 4710
rect 6071 4658 6073 4710
rect 6014 4643 6073 4658
rect 6153 4710 6210 4993
rect 6312 4880 7989 4936
rect 6153 4707 6253 4710
rect 6153 4655 6166 4707
rect 6218 4655 6253 4707
rect 6154 4652 6253 4655
rect 5706 3720 5820 3723
rect 5403 3661 5460 3674
rect 5403 3609 5405 3661
rect 5457 3609 5460 3661
rect 5706 3668 5745 3720
rect 5808 3668 5820 3720
rect 5706 3660 5820 3668
rect 5737 3659 5820 3660
rect 6014 3613 6070 4643
rect 6312 3619 6368 4880
rect 7933 4813 7989 4880
rect 7933 4773 7935 4813
rect 7869 4761 7935 4773
rect 7987 4761 7989 4813
rect 6715 4720 6812 4733
rect 6715 4649 6729 4720
rect 6800 4711 6812 4720
rect 7869 4717 7989 4761
rect 6807 4657 6812 4711
rect 7327 4710 7481 4711
rect 6800 4649 6812 4657
rect 6878 4707 6977 4710
rect 6878 4655 6890 4707
rect 6942 4655 6977 4707
rect 6878 4652 6977 4655
rect 6715 4634 6812 4649
rect 6171 3616 6368 3619
rect 5403 3597 5460 3609
rect 6013 3610 6089 3613
rect 6013 3597 6025 3610
rect 5403 3558 6025 3597
rect 6077 3558 6089 3610
rect 6171 3564 6183 3616
rect 6235 3564 6368 3616
rect 6171 3563 6368 3564
rect 6628 4512 6686 4524
rect 6628 4460 6632 4512
rect 6684 4460 6686 4512
rect 6628 3612 6686 4460
rect 6921 3719 6977 4652
rect 6920 3717 6977 3719
rect 6920 3665 6922 3717
rect 6974 3665 6977 3717
rect 6920 3661 6977 3665
rect 6921 3653 6977 3661
rect 7327 4707 7580 4710
rect 7327 4655 7493 4707
rect 7545 4655 7580 4707
rect 7327 4652 7580 4655
rect 7327 3613 7383 4652
rect 7869 3615 7925 4717
rect 8053 4712 8111 4993
rect 9267 4991 11225 5049
rect 8812 4800 8891 4805
rect 8812 4746 8825 4800
rect 8879 4746 8891 4800
rect 8812 4738 8891 4746
rect 8053 4660 8056 4712
rect 8108 4660 8111 4712
rect 8002 4604 8111 4660
rect 8002 3814 8058 4604
rect 8258 4547 8375 4563
rect 8258 4472 8268 4547
rect 8350 4472 8375 4547
rect 8258 4455 8375 4472
rect 8002 3758 8183 3814
rect 8002 3747 8058 3758
rect 7981 3725 8058 3747
rect 7981 3673 7993 3725
rect 8045 3673 8058 3725
rect 7981 3670 8058 3673
rect 7869 3613 7964 3615
rect 6628 3610 6839 3612
rect 6171 3562 6237 3563
rect 5403 3549 6089 3558
rect 6628 3558 6775 3610
rect 6827 3558 6839 3610
rect 6628 3555 6839 3558
rect 7327 3610 7426 3613
rect 7327 3558 7339 3610
rect 7391 3558 7426 3610
rect 7869 3561 7899 3613
rect 7951 3561 7964 3613
rect 7869 3559 7964 3561
rect 7327 3555 7426 3558
rect 5403 3547 6077 3549
rect 5403 3540 6069 3547
rect 7327 3484 7383 3555
rect 5504 3481 7383 3484
rect 5504 3429 5516 3481
rect 5568 3429 7383 3481
rect 5504 3428 7383 3429
rect 5514 3427 5570 3428
rect 5956 3201 6101 3204
rect 5956 3117 5970 3201
rect 6033 3117 6101 3201
rect 5956 3113 6101 3117
rect 5249 2869 5306 2931
rect 5204 2848 5347 2869
rect 5204 2780 5238 2848
rect 5316 2780 5347 2848
rect 5204 2754 5347 2780
rect 5471 2850 5574 2866
rect 5471 2770 5488 2850
rect 5557 2770 5574 2850
rect 5471 2751 5574 2770
rect 5027 2448 5095 2457
rect 5027 2387 5034 2448
rect 5087 2387 5095 2448
rect 5027 2373 5095 2387
rect 5027 2148 5112 2153
rect 5019 2140 5124 2148
rect 5019 2070 5043 2140
rect 5099 2070 5124 2140
rect 5019 1664 5124 2070
rect 5475 1811 5568 2751
rect 5763 2435 5877 2453
rect 5763 2376 5782 2435
rect 5855 2376 5877 2435
rect 5763 2359 5877 2376
rect 5774 1966 5864 2359
rect 5763 1950 5877 1966
rect 5763 1888 5782 1950
rect 5862 1888 5877 1950
rect 5763 1872 5877 1888
rect 5454 1795 5576 1811
rect 5454 1726 5479 1795
rect 5561 1726 5576 1795
rect 5454 1709 5576 1726
rect 5018 1652 5124 1664
rect 5018 1583 5026 1652
rect 5088 1583 5124 1652
rect 5018 1569 5124 1583
rect 5018 1565 5101 1569
rect 5960 1328 6101 3113
rect 7604 2836 7682 2861
rect 7604 2784 7614 2836
rect 7669 2784 7682 2836
rect 7604 1421 7682 2784
rect 8127 2151 8183 3758
rect 8278 3677 8337 4455
rect 8438 4290 8529 4298
rect 8438 4223 8450 4290
rect 8516 4283 8529 4290
rect 8820 4283 8878 4738
rect 8516 4225 8878 4283
rect 8516 4223 8529 4225
rect 8438 4217 8529 4223
rect 8820 3721 8878 4225
rect 9128 4708 9187 4720
rect 9128 4656 9133 4708
rect 9185 4656 9187 4708
rect 9128 4641 9187 4656
rect 9267 4708 9324 4991
rect 9426 4878 11103 4934
rect 9267 4705 9367 4708
rect 9267 4653 9280 4705
rect 9332 4653 9367 4705
rect 9268 4650 9367 4653
rect 8820 3718 8934 3721
rect 8278 3665 8352 3677
rect 8278 3612 8289 3665
rect 8343 3612 8352 3665
rect 8278 3599 8352 3612
rect 8517 3659 8574 3672
rect 8517 3607 8519 3659
rect 8571 3607 8574 3659
rect 8820 3666 8859 3718
rect 8922 3666 8934 3718
rect 8820 3658 8934 3666
rect 8851 3657 8934 3658
rect 9128 3611 9184 4641
rect 9426 3617 9482 4878
rect 11047 4811 11103 4878
rect 11047 4771 11049 4811
rect 10983 4759 11049 4771
rect 11101 4759 11103 4811
rect 9828 4718 9925 4731
rect 9828 4646 9841 4718
rect 9911 4708 9925 4718
rect 10983 4715 11103 4759
rect 10441 4708 10595 4709
rect 9920 4655 9925 4708
rect 9911 4646 9925 4655
rect 9992 4705 10091 4708
rect 9992 4653 10004 4705
rect 10056 4653 10091 4705
rect 9992 4650 10091 4653
rect 9828 4634 9925 4646
rect 9285 3614 9482 3617
rect 8113 2139 8194 2151
rect 8113 2067 8131 2139
rect 8187 2067 8194 2139
rect 8113 2053 8194 2067
rect 8278 1979 8337 3599
rect 8517 3595 8574 3607
rect 9127 3608 9203 3611
rect 9127 3595 9139 3608
rect 8517 3556 9139 3595
rect 9191 3556 9203 3608
rect 9285 3562 9297 3614
rect 9349 3562 9482 3614
rect 9285 3561 9482 3562
rect 9742 4510 9800 4522
rect 9742 4458 9746 4510
rect 9798 4458 9800 4510
rect 9742 3610 9800 4458
rect 10035 3717 10091 4650
rect 10034 3715 10091 3717
rect 10034 3663 10036 3715
rect 10088 3663 10091 3715
rect 10034 3659 10091 3663
rect 10035 3651 10091 3659
rect 10441 4705 10694 4708
rect 10441 4653 10607 4705
rect 10659 4653 10694 4705
rect 10441 4650 10694 4653
rect 10441 3611 10497 4650
rect 10983 3613 11039 4715
rect 11167 4710 11225 4991
rect 12426 4995 14384 5053
rect 11584 4818 11663 4823
rect 11583 4810 11663 4818
rect 11583 4757 11594 4810
rect 11651 4757 11663 4810
rect 11583 4751 11663 4757
rect 11584 4745 11663 4751
rect 11971 4804 12050 4809
rect 11971 4750 11984 4804
rect 12038 4750 12050 4804
rect 11167 4658 11170 4710
rect 11222 4658 11225 4710
rect 11116 4602 11225 4658
rect 11116 3798 11172 4602
rect 11372 4551 11479 4563
rect 11372 4472 11389 4551
rect 11465 4472 11479 4551
rect 11372 4454 11479 4472
rect 11589 4225 11658 4745
rect 11971 4742 12050 4750
rect 11282 4156 11658 4225
rect 11116 3745 11211 3798
rect 11095 3723 11211 3745
rect 11095 3671 11107 3723
rect 11159 3671 11211 3723
rect 11095 3668 11211 3671
rect 10983 3611 11078 3613
rect 9742 3608 9953 3610
rect 9285 3560 9351 3561
rect 8517 3547 9203 3556
rect 9742 3556 9889 3608
rect 9941 3556 9953 3608
rect 9742 3553 9953 3556
rect 10441 3608 10540 3611
rect 10441 3556 10453 3608
rect 10505 3556 10540 3608
rect 10983 3559 11013 3611
rect 11065 3559 11078 3611
rect 10983 3557 11078 3559
rect 10441 3553 10540 3556
rect 8517 3545 9191 3547
rect 8517 3538 9183 3545
rect 10441 3482 10497 3553
rect 8618 3479 8682 3482
rect 8618 3427 8630 3479
rect 8618 3426 8682 3427
rect 10491 3426 10497 3482
rect 8626 3404 8682 3426
rect 8687 2673 8781 2684
rect 8429 2639 8550 2662
rect 8429 2602 8447 2639
rect 8398 2555 8447 2602
rect 8537 2555 8550 2639
rect 8687 2615 8702 2673
rect 8769 2615 8781 2673
rect 8687 2600 8781 2615
rect 8398 2541 8550 2555
rect 8443 2434 8515 2448
rect 8443 2372 8455 2434
rect 8509 2372 8515 2434
rect 8443 2363 8515 2372
rect 7788 1920 8339 1979
rect 7600 1406 7683 1421
rect 7788 1420 7847 1920
rect 8445 1830 8512 2363
rect 8693 2288 8780 2600
rect 11154 2475 11211 3668
rect 11282 3040 11351 4156
rect 11475 4065 11565 4066
rect 11979 4065 12037 4742
rect 11475 4007 12037 4065
rect 11268 3021 11374 3040
rect 11268 2930 11284 3021
rect 11352 2930 11374 3021
rect 11268 2912 11374 2930
rect 11475 2702 11565 4007
rect 11979 3725 12037 4007
rect 12287 4712 12346 4724
rect 12287 4660 12292 4712
rect 12344 4660 12346 4712
rect 12287 4645 12346 4660
rect 12426 4712 12483 4995
rect 12585 4882 14262 4938
rect 12426 4709 12526 4712
rect 12426 4657 12439 4709
rect 12491 4657 12526 4709
rect 12427 4654 12526 4657
rect 11979 3722 12093 3725
rect 11676 3663 11733 3676
rect 11676 3611 11678 3663
rect 11730 3611 11733 3663
rect 11979 3670 12018 3722
rect 12081 3670 12093 3722
rect 11979 3662 12093 3670
rect 12010 3661 12093 3662
rect 12287 3615 12343 4645
rect 12585 3621 12641 4882
rect 14206 4815 14262 4882
rect 14206 4775 14208 4815
rect 14142 4763 14208 4775
rect 14260 4763 14262 4815
rect 12997 4722 13094 4731
rect 12997 4652 13007 4722
rect 13083 4652 13094 4722
rect 14142 4719 14262 4763
rect 13600 4712 13754 4713
rect 13151 4709 13250 4712
rect 13151 4657 13163 4709
rect 13215 4707 13250 4709
rect 13600 4709 13853 4712
rect 13215 4657 13264 4707
rect 13151 4654 13264 4657
rect 12997 4634 13094 4652
rect 12444 3618 12641 3621
rect 11676 3599 11733 3611
rect 12286 3612 12362 3615
rect 12286 3599 12298 3612
rect 11676 3560 12298 3599
rect 12350 3560 12362 3612
rect 12444 3566 12456 3618
rect 12508 3566 12641 3618
rect 12444 3565 12641 3566
rect 12901 4514 12959 4526
rect 12901 4462 12905 4514
rect 12957 4462 12959 4514
rect 12901 3614 12959 4462
rect 13188 3719 13264 4654
rect 13188 3667 13195 3719
rect 13247 3667 13264 3719
rect 13188 3663 13264 3667
rect 13600 4657 13766 4709
rect 13818 4657 13853 4709
rect 13600 4654 13853 4657
rect 13194 3655 13250 3663
rect 13600 3615 13656 4654
rect 14142 3617 14198 4719
rect 14326 4714 14384 4995
rect 14326 4665 14329 4714
rect 14280 4662 14329 4665
rect 14381 4662 14384 4714
rect 14275 4606 14384 4662
rect 14275 3749 14364 4606
rect 14254 3737 14364 3749
rect 14254 3727 14411 3737
rect 14254 3675 14266 3727
rect 14318 3675 14411 3727
rect 14254 3672 14411 3675
rect 14142 3615 14237 3617
rect 12901 3612 13112 3614
rect 12444 3564 12510 3565
rect 11676 3551 12362 3560
rect 12901 3560 13048 3612
rect 13100 3560 13112 3612
rect 12901 3557 13112 3560
rect 13600 3612 13699 3615
rect 13600 3560 13612 3612
rect 13664 3560 13699 3612
rect 14142 3563 14172 3615
rect 14224 3563 14237 3615
rect 14142 3561 14237 3563
rect 13600 3557 13699 3560
rect 11676 3549 12350 3551
rect 11676 3542 12342 3549
rect 13600 3486 13656 3557
rect 11777 3483 13656 3486
rect 11777 3431 11789 3483
rect 11841 3431 13656 3483
rect 11777 3430 13656 3431
rect 11787 3429 11843 3430
rect 14327 2866 14411 3672
rect 14327 2854 14421 2866
rect 14327 2791 14343 2854
rect 14330 2790 14343 2791
rect 14411 2790 14421 2854
rect 14330 2780 14421 2790
rect 11464 2681 11582 2702
rect 11464 2586 11484 2681
rect 11567 2586 11582 2681
rect 11464 2570 11582 2586
rect 11154 2455 11212 2475
rect 11139 2440 11223 2455
rect 11139 2364 11150 2440
rect 11211 2364 11223 2440
rect 11139 2353 11223 2364
rect 8692 2269 8780 2288
rect 8692 2217 8708 2269
rect 8766 2217 8780 2269
rect 8692 2204 8780 2217
rect 10530 2280 10750 2291
rect 10530 2217 10552 2280
rect 10604 2217 10664 2280
rect 10716 2217 10750 2280
rect 10530 2155 10750 2217
rect 10530 2103 10590 2155
rect 10679 2103 10750 2155
rect 10530 2100 10750 2103
rect 9016 1952 9096 1961
rect 9016 1900 9024 1952
rect 9082 1900 9096 1952
rect 9016 1887 9096 1900
rect 8213 1763 8512 1830
rect 8213 1525 8280 1763
rect 8213 1509 8319 1525
rect 8213 1457 8256 1509
rect 8309 1457 8319 1509
rect 9027 1480 9093 1887
rect 10548 1689 10673 2100
rect 10802 1952 10870 1964
rect 11162 1952 11223 1962
rect 10802 1951 11223 1952
rect 10802 1899 10807 1951
rect 10865 1899 11223 1951
rect 10802 1891 11223 1899
rect 10802 1886 10870 1891
rect 11162 1801 11223 1891
rect 11162 1791 11240 1801
rect 11162 1739 11175 1791
rect 11229 1739 11240 1791
rect 11162 1728 11240 1739
rect 11305 1790 11383 1802
rect 11305 1738 11323 1790
rect 11376 1738 11383 1790
rect 11305 1729 11383 1738
rect 10548 1628 10596 1689
rect 10657 1628 10673 1689
rect 10548 1605 10673 1628
rect 10581 1604 10673 1605
rect 8213 1439 8319 1457
rect 8990 1477 9098 1480
rect 8990 1464 9099 1477
rect 5960 1244 5972 1328
rect 6035 1244 6101 1328
rect 7103 1359 7185 1370
rect 7103 1306 7117 1359
rect 7169 1306 7185 1359
rect 7600 1354 7613 1406
rect 7668 1354 7683 1406
rect 7600 1346 7683 1354
rect 7745 1408 7847 1420
rect 7745 1356 7762 1408
rect 7832 1356 7847 1408
rect 7745 1345 7847 1356
rect 8487 1410 8581 1414
rect 8487 1357 8501 1410
rect 8560 1357 8581 1410
rect 8990 1412 9018 1464
rect 9080 1412 9099 1464
rect 8990 1401 9098 1412
rect 8487 1348 8581 1357
rect 7103 1293 7185 1306
rect 5960 1233 6101 1244
rect 7108 1273 7185 1293
rect 8502 1273 8562 1348
rect 5960 1227 6042 1233
rect 7108 1213 8562 1273
rect 9148 1134 9232 1146
rect 7993 1124 8065 1129
rect 9148 1124 9161 1134
rect 7993 1117 9161 1124
rect 7993 1063 8005 1117
rect 8058 1066 9161 1117
rect 9221 1066 9232 1134
rect 8058 1063 9232 1066
rect 7993 1054 9232 1063
rect 7993 1051 8065 1054
rect 9148 1046 9232 1054
rect 4831 903 4954 960
rect 11323 903 11380 1729
rect 4831 786 11380 903
<< via2 >>
rect 3606 5386 3667 5394
rect 3606 5333 3611 5386
rect 3611 5333 3664 5386
rect 3664 5333 3667 5386
rect 3606 5327 3667 5333
rect 2260 4471 2325 4545
rect 3604 4707 3678 4722
rect 3604 4655 3611 4707
rect 3611 4655 3666 4707
rect 3666 4655 3678 4707
rect 3604 4649 3678 4655
rect 5162 4547 5251 4556
rect 5162 4464 5169 4547
rect 5169 4464 5241 4547
rect 5241 4464 5251 4547
rect 5162 4462 5251 4464
rect 6729 4711 6800 4720
rect 6729 4657 6753 4711
rect 6753 4657 6800 4711
rect 6729 4649 6800 4657
rect 8268 4472 8350 4547
rect 8450 4223 8516 4290
rect 9841 4708 9911 4718
rect 9841 4655 9866 4708
rect 9866 4655 9911 4708
rect 9841 4646 9911 4655
rect 11389 4544 11465 4551
rect 11389 4480 11395 4544
rect 11395 4480 11456 4544
rect 11456 4480 11465 4544
rect 11389 4472 11465 4480
rect 8447 2627 8537 2639
rect 8447 2571 8457 2627
rect 8457 2571 8525 2627
rect 8525 2571 8537 2627
rect 8447 2555 8537 2571
rect 13007 4713 13083 4722
rect 13007 4661 13018 4713
rect 13018 4661 13079 4713
rect 13079 4661 13083 4713
rect 13007 4652 13083 4661
<< metal3 >>
rect 3595 5394 3676 5401
rect 3595 5327 3606 5394
rect 3667 5327 3676 5394
rect 3595 4782 3676 5327
rect 3595 4722 13107 4782
rect 3595 4649 3604 4722
rect 3678 4720 13007 4722
rect 3678 4649 6729 4720
rect 6800 4718 13007 4720
rect 6800 4649 9841 4718
rect 3595 4646 9841 4649
rect 9911 4652 13007 4718
rect 13083 4652 13107 4722
rect 9911 4646 13107 4652
rect 3595 4634 13107 4646
rect 2244 4556 11480 4563
rect 2244 4545 5162 4556
rect 2244 4471 2260 4545
rect 2325 4471 5162 4545
rect 2244 4462 5162 4471
rect 5251 4551 11480 4556
rect 5251 4547 11389 4551
rect 5251 4472 8268 4547
rect 8350 4472 11389 4547
rect 11465 4472 11480 4551
rect 5251 4462 11480 4472
rect 2244 4391 11480 4462
rect 8438 4290 8531 4302
rect 8438 4286 8450 4290
rect 8398 4223 8450 4286
rect 8516 4223 8531 4290
rect 8398 4209 8531 4223
rect 8398 2665 8509 4209
rect 8398 2639 8550 2665
rect 8398 2555 8447 2639
rect 8537 2555 8550 2639
rect 8398 2541 8550 2555
use and2_mag  and2_mag_0
timestamp 1695127730
transform 1 0 -188 0 -1 4489
box -70 -188 1009 863
use and2_mag  and2_mag_1
timestamp 1695127730
transform 1 0 1217 0 1 2472
box -70 -188 1009 863
use and2_mag  and2_mag_2
timestamp 1695127730
transform 1 0 -195 0 -1 2302
box -70 -188 1009 863
use and2_mag  and2_mag_3
timestamp 1695127730
transform 1 0 8176 0 -1 1774
box -70 -188 1009 863
use Buffer_delayed_mag  Buffer_delayed_mag_0
timestamp 1694693600
transform 1 0 6232 0 -1 1777
box -218 -175 878 631
use Buffer_delayed_mag  Buffer_delayed_mag_1
timestamp 1694693600
transform 1 0 9835 0 -1 1535
box -218 -175 878 631
use GF_INV_MAG  GF_INV_MAG_0
timestamp 1695119997
transform 1 0 734 0 1 2875
box -118 -175 286 631
use GF_INV_MAG  GF_INV_MAG_1
timestamp 1695119997
transform 1 0 9435 0 -1 1537
box -118 -175 286 631
use GF_INV_MAG  GF_INV_MAG_2
timestamp 1695119997
transform 1 0 11832 0 -1 1539
box -118 -175 286 631
use JK_FF_mag  JK_FF_mag_0
timestamp 1695127730
transform 1 0 2513 0 -1 5259
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_1
timestamp 1695127730
transform 1 0 5648 0 -1 5261
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_2
timestamp 1695127730
transform 1 0 8762 0 -1 5259
box -390 0 2603 2148
use JK_FF_mag  JK_FF_mag_3
timestamp 1695127730
transform 1 0 11921 0 -1 5263
box -390 0 2603 2148
use nand3_mag  nand3_mag_0
timestamp 1694691991
transform 1 0 -188 0 1 2763
box -70 -188 671 863
use nand3_mag  nand3_mag_1
timestamp 1694691991
transform 1 0 7311 0 -1 1771
box -70 -188 671 863
use nor_3_mag  nor_3_mag_0
timestamp 1695119997
transform 1 0 10521 0 -1 2682
box 329 440 1054 1778
use or_2  or_2_0
timestamp 1694669839
transform 1 0 1154 0 1 2104
box 0 0 1 1
use or_2  or_2_1
timestamp 1694669839
transform 1 0 1468 0 1 3710
box 0 0 1 1
use or_2_mag  or_2_mag_0
timestamp 1695127730
transform 1 0 379 0 -1 5033
box 330 510 1401 1521
use or_2_mag  or_2_mag_1
timestamp 1695127730
transform 1 0 817 0 -1 2795
box 330 510 1401 1521
use or_2_mag  or_2_mag_3
timestamp 1695127730
transform 1 0 2289 0 -1 2798
box 330 510 1401 1521
<< labels >>
flabel metal1 3090 1030 3090 1030 0 FreeSans 640 0 0 0 VDD
port 0 nsew
flabel metal1 4600 5390 4600 5390 0 FreeSans 640 0 0 0 VSS
port 1 nsew
flabel via2 3640 5360 3640 5360 0 FreeSans 640 0 0 0 RST
port 2 nsew
flabel via1 1910 5220 1910 5220 0 FreeSans 640 0 0 0 CLK
port 3 nsew
flabel metal1 12200 1380 12200 1380 0 FreeSans 640 0 0 0 Vdiv11
port 4 nsew
flabel metal2 4940 3710 4940 3710 0 FreeSans 640 0 0 0 Q3
port 5 nsew
flabel metal1 8080 3710 8080 3710 0 FreeSans 640 0 0 0 Q2
port 6 nsew
flabel metal2 11190 3710 11190 3710 0 FreeSans 640 0 0 0 Q1
port 7 nsew
flabel metal2 14350 3720 14350 3720 0 FreeSans 640 0 0 0 Q0
port 8 nsew
<< end >>
