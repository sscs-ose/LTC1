magic
tech gf180mcuC
magscale 1 10
timestamp 1699956126
<< pwell >>
rect -162 -168 162 168
<< nmos >>
rect -50 -100 50 100
<< ndiff >>
rect -138 87 -50 100
rect -138 -87 -125 87
rect -79 -87 -50 87
rect -138 -100 -50 -87
rect 50 87 138 100
rect 50 -87 79 87
rect 125 -87 138 87
rect 50 -100 138 -87
<< ndiffc >>
rect -125 -87 -79 87
rect 79 -87 125 87
<< polysilicon >>
rect -50 100 50 144
rect -50 -144 50 -100
<< metal1 >>
rect -125 87 -79 98
rect -125 -98 -79 -87
rect 79 87 125 98
rect 79 -98 125 -87
<< properties >>
string gencell nfet_03v3
string library gf180mcu
string parameters w 1 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.28 wmin 0.22 full_metal 0 compatible {nfet_03v3 nfet_06v0 nfet_06v0_nvt}
<< end >>
