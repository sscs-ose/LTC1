* NGSPICE file created from Transmission_Gate_Layout_flat.ext - technology: gf180mcuC

.subckt Transmission_Gate_Layout_flat VSS VDD CLK VIN VOUT
X0 VOUT CLK.t0 VIN.t33 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X1 VIN CLK.t1 VOUT.t32 VSS.t10 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X2 VIN a_n120_68.t6 VOUT.t46 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 VIN CLK.t2 VOUT.t31 VSS.t10 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X4 VOUT CLK.t3 VIN.t32 VSS.t9 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X5 VOUT a_n120_68.t7 VIN.t47 VDD.t10 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X6 VOUT a_n120_68.t8 VIN.t8 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X7 VIN a_n120_68.t9 VOUT.t9 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X8 VOUT a_n120_68.t10 VIN.t35 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X9 VIN a_n120_68.t11 VOUT.t36 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X10 VIN a_n120_68.t12 VOUT.t44 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X11 VIN a_n120_68.t13 VOUT.t45 VDD.t5 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X12 VIN CLK.t4 VOUT.t29 VSS.t8 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X13 VOUT CLK.t5 VIN.t31 VSS.t4 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X14 VIN CLK.t6 VOUT.t27 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X15 VOUT a_n120_68.t14 VIN.t6 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X16 VIN a_n120_68.t15 VOUT.t7 VDD.t5 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X17 VOUT CLK.t8 VIN.t30 VSS.t4 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X18 VIN CLK.t9 VOUT.t25 VSS.t10 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X19 VOUT CLK.t10 VIN.t29 VSS.t9 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X20 VOUT CLK.t11 VIN.t28 VSS.t9 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X21 VIN a_n120_68.t16 VOUT.t34 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X22 VOUT a_n120_68.t17 VIN.t37 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X23 VOUT a_n120_68.t18 VIN.t38 VDD.t10 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X24 VOUT a_n120_68.t19 VIN.t42 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X25 VIN CLK.t13 VOUT.t22 VSS.t8 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X26 VOUT CLK.t14 VIN.t27 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X27 VIN a_n120_68.t20 VOUT.t43 VDD.t11 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X28 VIN a_n120_68.t21 VOUT.t4 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X29 VIN CLK.t15 VOUT.t20 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X30 VOUT a_n120_68.t22 VIN.t5 VDD.t10 pfet_03v3 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.28u
X31 VOUT a_n120_68.t23 VIN.t2 VDD.t9 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X32 VIN a_n120_68.t24 VOUT.t3 VDD.t8 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X33 VIN CLK.t16 VOUT.t19 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X34 VIN CLK.t17 VOUT.t18 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X35 VIN CLK.t18 VOUT.t17 VSS.t8 nfet_03v3 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.28u
X36 VIN a_n120_68.t25 VOUT.t41 VDD.t7 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X37 VOUT a_n120_68.t26 VIN.t0 VDD.t6 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X38 VOUT CLK.t20 VIN.t26 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X39 VOUT CLK.t21 VIN.t25 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X40 VIN a_n120_68.t27 VOUT.t1 VDD.t5 pfet_03v3 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.28u
X41 VOUT a_n120_68.t28 VIN.t39 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X42 VIN CLK.t23 VOUT.t14 VSS.t6 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X43 VOUT CLK.t24 VIN.t24 VSS.t5 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X44 VOUT a_n120_68.t29 VIN.t40 VDD.t4 pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X45 VOUT CLK.t26 VIN.t23 VSS.t4 nfet_03v3 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.28u
X46 VOUT CLK.t27 VIN.t22 VSS.t3 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
X47 VIN CLK.t29 VOUT.t10 VSS.t0 nfet_03v3 ad=0.325p pd=1.77u as=0.325p ps=1.77u w=1.25u l=0.28u
R0 CLK.t25 CLK.t12 82.9076
R1 CLK.t22 CLK.t25 82.9076
R2 CLK.t19 CLK.n6 56.4451
R3 CLK.t13 CLK.t4 50.3184
R4 CLK.t18 CLK.t13 50.3184
R5 CLK.t0 CLK.t20 50.3184
R6 CLK.t27 CLK.t0 50.3184
R7 CLK.t23 CLK.t15 50.3184
R8 CLK.t6 CLK.t23 50.3184
R9 CLK.t10 CLK.t3 50.3184
R10 CLK.t11 CLK.t10 50.3184
R11 CLK.t29 CLK.t16 50.3184
R12 CLK.t17 CLK.t29 50.3184
R13 CLK.t21 CLK.t14 50.3184
R14 CLK.t24 CLK.t21 50.3184
R15 CLK.t9 CLK.t2 50.3184
R16 CLK.t1 CLK.t9 50.3184
R17 CLK.t5 CLK.t26 50.3184
R18 CLK.t8 CLK.t5 50.3184
R19 CLK.t7 CLK.t19 50.3184
R20 CLK.t28 CLK.t7 50.3184
R21 CLK.n7 CLK.t22 49.7969
R22 CLK.n0 CLK.t18 39.7594
R23 CLK.n7 CLK.t28 31.1559
R24 CLK.n1 CLK.n0 20.8576
R25 CLK.n2 CLK.n1 20.8576
R26 CLK.n3 CLK.n2 20.8576
R27 CLK.n4 CLK.n3 20.8576
R28 CLK.n5 CLK.n4 20.8576
R29 CLK.n6 CLK.n5 20.8576
R30 CLK.n0 CLK.t27 18.9023
R31 CLK.n1 CLK.t6 18.9023
R32 CLK.n2 CLK.t11 18.9023
R33 CLK.n3 CLK.t17 18.9023
R34 CLK.n4 CLK.t24 18.9023
R35 CLK.n5 CLK.t1 18.9023
R36 CLK.n6 CLK.t8 18.9023
R37 CLK.n8 CLK.n7 17.8594
R38 CLK CLK.n8 8.0005
R39 CLK CLK.n8 8.0005
R40 VIN.n42 VIN.n40 5.21612
R41 VIN.n48 VIN.t23 4.4609
R42 VIN.n47 VIN.t31 4.4609
R43 VIN.n46 VIN.t30 4.4609
R44 VIN.n44 VIN.n43 4.4609
R45 VIN.n42 VIN.n41 4.4609
R46 VIN.n22 VIN.n21 3.90572
R47 VIN.n36 VIN.n33 3.90572
R48 VIN.n30 VIN.n29 3.90572
R49 VIN.n12 VIN.n9 3.84485
R50 VIN.n4 VIN.n1 3.84485
R51 VIN.n62 VIN.n61 3.84485
R52 VIN.n66 VIN.n65 3.3285
R53 VIN.n68 VIN.n67 3.3285
R54 VIN.n70 VIN.n69 3.3285
R55 VIN.n55 VIN.t47 3.3285
R56 VIN.n54 VIN.t5 3.3285
R57 VIN.n53 VIN.t38 3.3285
R58 VIN.n22 VIN.n19 3.1505
R59 VIN.n23 VIN.n17 3.1505
R60 VIN.n36 VIN.n35 3.1505
R61 VIN.n39 VIN.n38 3.1505
R62 VIN.n30 VIN.n27 3.1505
R63 VIN.n31 VIN.n25 3.1505
R64 VIN.n64 VIN.n55 2.72398
R65 VIN.n12 VIN.n11 2.6005
R66 VIN.n15 VIN.n14 2.6005
R67 VIN.n4 VIN.n3 2.6005
R68 VIN.n7 VIN.n6 2.6005
R69 VIN.n62 VIN.n59 2.6005
R70 VIN.n63 VIN.n57 2.6005
R71 VIN.n46 VIN.n45 2.47941
R72 VIN.n17 VIN.t32 1.3109
R73 VIN.n17 VIN.n16 1.3109
R74 VIN.n19 VIN.t29 1.3109
R75 VIN.n19 VIN.n18 1.3109
R76 VIN.n21 VIN.t28 1.3109
R77 VIN.n21 VIN.n20 1.3109
R78 VIN.n38 VIN.t22 1.3109
R79 VIN.n38 VIN.n37 1.3109
R80 VIN.n35 VIN.t33 1.3109
R81 VIN.n35 VIN.n34 1.3109
R82 VIN.n33 VIN.t26 1.3109
R83 VIN.n33 VIN.n32 1.3109
R84 VIN.n25 VIN.t27 1.3109
R85 VIN.n25 VIN.n24 1.3109
R86 VIN.n27 VIN.t25 1.3109
R87 VIN.n27 VIN.n26 1.3109
R88 VIN.n29 VIN.t24 1.3109
R89 VIN.n29 VIN.n28 1.3109
R90 VIN.n15 VIN.n12 1.24485
R91 VIN.n7 VIN.n4 1.24485
R92 VIN.n55 VIN.n54 1.24485
R93 VIN.n54 VIN.n53 1.24485
R94 VIN.n63 VIN.n62 1.24485
R95 VIN.n68 VIN.n66 1.24485
R96 VIN.n70 VIN.n68 1.24485
R97 VIN.n53 VIN.n52 1.2018
R98 VIN.n66 VIN.n64 1.2018
R99 VIN VIN.n70 1.05507
R100 VIN.n45 VIN.n44 0.957239
R101 VIN.n49 VIN.n48 0.957239
R102 VIN.n23 VIN.n22 0.755717
R103 VIN.n39 VIN.n36 0.755717
R104 VIN.n44 VIN.n42 0.755717
R105 VIN.n48 VIN.n47 0.755717
R106 VIN.n47 VIN.n46 0.755717
R107 VIN.n31 VIN.n30 0.755717
R108 VIN.n57 VIN.t8 0.7285
R109 VIN.n57 VIN.n56 0.7285
R110 VIN.n59 VIN.t2 0.7285
R111 VIN.n59 VIN.n58 0.7285
R112 VIN.n61 VIN.t42 0.7285
R113 VIN.n61 VIN.n60 0.7285
R114 VIN.n14 VIN.t39 0.7285
R115 VIN.n14 VIN.n13 0.7285
R116 VIN.n11 VIN.t40 0.7285
R117 VIN.n11 VIN.n10 0.7285
R118 VIN.n9 VIN.t37 0.7285
R119 VIN.n9 VIN.n8 0.7285
R120 VIN.n6 VIN.t35 0.7285
R121 VIN.n6 VIN.n5 0.7285
R122 VIN.n3 VIN.t6 0.7285
R123 VIN.n3 VIN.n2 0.7285
R124 VIN.n1 VIN.t0 0.7285
R125 VIN.n1 VIN.n0 0.7285
R126 VIN.n50 VIN.n49 0.626587
R127 VIN.n52 VIN.n51 0.626587
R128 VIN.n51 VIN.n15 0.575717
R129 VIN.n52 VIN.n7 0.575717
R130 VIN.n64 VIN.n63 0.575717
R131 VIN.n50 VIN.n23 0.331152
R132 VIN.n45 VIN.n39 0.331152
R133 VIN.n49 VIN.n31 0.331152
R134 VIN.n51 VIN.n50 0.239196
R135 VOUT.n44 VOUT.n41 3.90572
R136 VOUT.n52 VOUT.n49 3.90572
R137 VOUT.n67 VOUT.n66 3.90572
R138 VOUT.n22 VOUT.n21 3.84485
R139 VOUT.n14 VOUT.n13 3.84485
R140 VOUT.n4 VOUT.n1 3.84485
R141 VOUT.n44 VOUT.n43 3.1505
R142 VOUT.n47 VOUT.n46 3.1505
R143 VOUT.n52 VOUT.n51 3.1505
R144 VOUT.n55 VOUT.n54 3.1505
R145 VOUT.n57 VOUT.n39 3.1505
R146 VOUT.n58 VOUT.n37 3.1505
R147 VOUT.n59 VOUT.n35 3.1505
R148 VOUT.n67 VOUT.n64 3.1505
R149 VOUT.n68 VOUT.n62 3.1505
R150 VOUT.n22 VOUT.n19 2.6005
R151 VOUT.n23 VOUT.n17 2.6005
R152 VOUT.n14 VOUT.n11 2.6005
R153 VOUT.n15 VOUT.n9 2.6005
R154 VOUT.n33 VOUT.n32 2.6005
R155 VOUT.n30 VOUT.n29 2.6005
R156 VOUT.n27 VOUT.n26 2.6005
R157 VOUT.n4 VOUT.n3 2.6005
R158 VOUT.n7 VOUT.n6 2.6005
R159 VOUT.n62 VOUT.t29 1.3109
R160 VOUT.n62 VOUT.n61 1.3109
R161 VOUT.n64 VOUT.t22 1.3109
R162 VOUT.n64 VOUT.n63 1.3109
R163 VOUT.n66 VOUT.t17 1.3109
R164 VOUT.n66 VOUT.n65 1.3109
R165 VOUT.n35 VOUT.t20 1.3109
R166 VOUT.n35 VOUT.n34 1.3109
R167 VOUT.n37 VOUT.t14 1.3109
R168 VOUT.n37 VOUT.n36 1.3109
R169 VOUT.n39 VOUT.t27 1.3109
R170 VOUT.n39 VOUT.n38 1.3109
R171 VOUT.n46 VOUT.t18 1.3109
R172 VOUT.n46 VOUT.n45 1.3109
R173 VOUT.n43 VOUT.t10 1.3109
R174 VOUT.n43 VOUT.n42 1.3109
R175 VOUT.n41 VOUT.t19 1.3109
R176 VOUT.n41 VOUT.n40 1.3109
R177 VOUT.n54 VOUT.t32 1.3109
R178 VOUT.n54 VOUT.n53 1.3109
R179 VOUT.n51 VOUT.t25 1.3109
R180 VOUT.n51 VOUT.n50 1.3109
R181 VOUT.n49 VOUT.t31 1.3109
R182 VOUT.n49 VOUT.n48 1.3109
R183 VOUT.n23 VOUT.n22 1.24485
R184 VOUT.n15 VOUT.n14 1.24485
R185 VOUT.n30 VOUT.n27 1.24485
R186 VOUT.n33 VOUT.n30 1.24485
R187 VOUT.n7 VOUT.n4 1.24485
R188 VOUT.n24 VOUT.n23 1.2018
R189 VOUT.n27 VOUT.n24 1.2018
R190 VOUT.n56 VOUT.n55 0.957239
R191 VOUT.n57 VOUT.n56 0.957239
R192 VOUT.n70 VOUT.n7 0.947457
R193 VOUT.n60 VOUT.n33 0.904413
R194 VOUT.n47 VOUT.n44 0.755717
R195 VOUT.n55 VOUT.n52 0.755717
R196 VOUT.n59 VOUT.n58 0.755717
R197 VOUT.n58 VOUT.n57 0.755717
R198 VOUT.n68 VOUT.n67 0.755717
R199 VOUT.n6 VOUT.t45 0.7285
R200 VOUT.n6 VOUT.n5 0.7285
R201 VOUT.n3 VOUT.t7 0.7285
R202 VOUT.n3 VOUT.n2 0.7285
R203 VOUT.n1 VOUT.t1 0.7285
R204 VOUT.n1 VOUT.n0 0.7285
R205 VOUT.n26 VOUT.t36 0.7285
R206 VOUT.n26 VOUT.n25 0.7285
R207 VOUT.n29 VOUT.t3 0.7285
R208 VOUT.n29 VOUT.n28 0.7285
R209 VOUT.n32 VOUT.t4 0.7285
R210 VOUT.n32 VOUT.n31 0.7285
R211 VOUT.n17 VOUT.t46 0.7285
R212 VOUT.n17 VOUT.n16 0.7285
R213 VOUT.n19 VOUT.t43 0.7285
R214 VOUT.n19 VOUT.n18 0.7285
R215 VOUT.n21 VOUT.t34 0.7285
R216 VOUT.n21 VOUT.n20 0.7285
R217 VOUT.n9 VOUT.t41 0.7285
R218 VOUT.n9 VOUT.n8 0.7285
R219 VOUT.n11 VOUT.t44 0.7285
R220 VOUT.n11 VOUT.n10 0.7285
R221 VOUT.n13 VOUT.t9 0.7285
R222 VOUT.n13 VOUT.n12 0.7285
R223 VOUT.n69 VOUT.n60 0.581587
R224 VOUT.n24 VOUT.n15 0.575717
R225 VOUT VOUT.n70 0.479848
R226 VOUT.n69 VOUT.n68 0.376152
R227 VOUT.n56 VOUT.n47 0.331152
R228 VOUT.n60 VOUT.n59 0.331152
R229 VOUT.n70 VOUT.n69 0.00245652
R230 VSS.n42 VSS.t5 95.3395
R231 VSS.n6 VSS.t6 82.6276
R232 VSS.n3 VSS.t3 57.2039
R233 VSS.n39 VSS.t10 44.492
R234 VSS.n18 VSS.t0 36.0174
R235 VSS.n12 VSS.t9 23.3056
R236 VSS.n33 VSS.t4 14.831
R237 VSS.n2 VSS.t8 6.09629
R238 VSS.n21 VSS.t2 5.21612
R239 VSS.n24 VSS.t1 4.5767
R240 VSS.n21 VSS.t11 4.4609
R241 VSS.n22 VSS.t7 4.4609
R242 VSS.n1 VSS.n0 2.6005
R243 VSS.n5 VSS.n4 2.6005
R244 VSS.n4 VSS.n3 2.6005
R245 VSS.n8 VSS.n7 2.6005
R246 VSS.n7 VSS.n6 2.6005
R247 VSS.n11 VSS.n10 2.6005
R248 VSS.n10 VSS.n9 2.6005
R249 VSS.n14 VSS.n13 2.6005
R250 VSS.n13 VSS.n12 2.6005
R251 VSS.n17 VSS.n16 2.6005
R252 VSS.n16 VSS.n15 2.6005
R253 VSS.n20 VSS.n19 2.6005
R254 VSS.n19 VSS.n18 2.6005
R255 VSS.n47 VSS.n46 2.6005
R256 VSS.n46 VSS.n45 2.6005
R257 VSS.n44 VSS.n43 2.6005
R258 VSS.n43 VSS.n42 2.6005
R259 VSS.n41 VSS.n40 2.6005
R260 VSS.n40 VSS.n39 2.6005
R261 VSS.n38 VSS.n37 2.6005
R262 VSS.n37 VSS.n36 2.6005
R263 VSS.n35 VSS.n34 2.6005
R264 VSS.n34 VSS.n33 2.6005
R265 VSS.n32 VSS.n31 2.6005
R266 VSS.n31 VSS.n30 2.6005
R267 VSS.n29 VSS.n28 2.6005
R268 VSS.n28 VSS.n27 2.6005
R269 VSS.n26 VSS.n25 2.6005
R270 VSS.n2 VSS.n1 1.71016
R271 VSS.n22 VSS.n21 0.755717
R272 VSS.n23 VSS.n22 0.691152
R273 VSS.n5 VSS.n2 0.482242
R274 VSS.n25 VSS.n24 0.11254
R275 VSS.n8 VSS.n5 0.0760357
R276 VSS.n11 VSS.n8 0.0760357
R277 VSS.n14 VSS.n11 0.0760357
R278 VSS.n17 VSS.n14 0.0760357
R279 VSS.n20 VSS.n17 0.0760357
R280 VSS.n47 VSS.n44 0.0760357
R281 VSS.n44 VSS.n41 0.0760357
R282 VSS.n41 VSS.n38 0.0760357
R283 VSS.n38 VSS.n35 0.0760357
R284 VSS.n35 VSS.n32 0.0760357
R285 VSS.n32 VSS.n29 0.0760357
R286 VSS.n29 VSS.n26 0.0760357
R287 VSS.n26 VSS.n23 0.0639821
R288 VSS VSS.n47 0.0422857
R289 VSS VSS.n20 0.03425
R290 a_n120_68.t20 a_n120_68.t16 82.9076
R291 a_n120_68.t6 a_n120_68.t20 82.9076
R292 a_n120_68.t14 a_n120_68.t10 82.9076
R293 a_n120_68.t26 a_n120_68.t14 82.9076
R294 a_n120_68.t12 a_n120_68.t9 82.9076
R295 a_n120_68.t25 a_n120_68.t12 82.9076
R296 a_n120_68.t29 a_n120_68.t28 82.9076
R297 a_n120_68.t17 a_n120_68.t29 82.9076
R298 a_n120_68.t24 a_n120_68.t21 82.9076
R299 a_n120_68.t11 a_n120_68.t24 82.9076
R300 a_n120_68.t23 a_n120_68.t19 82.9076
R301 a_n120_68.t8 a_n120_68.t23 82.9076
R302 a_n120_68.t15 a_n120_68.t13 82.9076
R303 a_n120_68.t27 a_n120_68.t15 82.9076
R304 a_n120_68.t22 a_n120_68.t7 82.9076
R305 a_n120_68.t18 a_n120_68.t22 82.9076
R306 a_n120_68.n11 a_n120_68.t18 74.3934
R307 a_n120_68.n5 a_n120_68.t27 56.0541
R308 a_n120_68.t7 a_n120_68.n10 56.0541
R309 a_n120_68.n10 a_n120_68.t6 35.1969
R310 a_n120_68.n9 a_n120_68.t26 35.1969
R311 a_n120_68.n8 a_n120_68.t25 35.1969
R312 a_n120_68.n7 a_n120_68.t17 35.1969
R313 a_n120_68.n6 a_n120_68.t11 35.1969
R314 a_n120_68.n5 a_n120_68.t8 35.1969
R315 a_n120_68.n6 a_n120_68.n5 20.8576
R316 a_n120_68.n7 a_n120_68.n6 20.8576
R317 a_n120_68.n8 a_n120_68.n7 20.8576
R318 a_n120_68.n9 a_n120_68.n8 20.8576
R319 a_n120_68.n10 a_n120_68.n9 20.8576
R320 a_n120_68.n15 a_n120_68.n14 5.21612
R321 a_n120_68.n2 a_n120_68.n0 4.57285
R322 a_n120_68.n13 a_n120_68.n12 4.4609
R323 a_n120_68.n16 a_n120_68.n15 4.4609
R324 a_n120_68.n2 a_n120_68.n1 3.3285
R325 a_n120_68.n4 a_n120_68.n3 3.3285
R326 a_n120_68.n4 a_n120_68.n2 1.24485
R327 a_n120_68.n15 a_n120_68.n13 0.755717
R328 a_n120_68.n11 a_n120_68.n4 0.750969
R329 a_n120_68.n13 a_n120_68.n11 0.510317
R330 VDD.n47 VDD.t6 40.9622
R331 VDD.n0 VDD.t5 20.4814
R332 VDD.n31 VDD.t0 20.4814
R333 VDD.n40 VDD.t10 17.8099
R334 VDD.n15 VDD.t4 16.029
R335 VDD.n18 VDD.t7 13.3576
R336 VDD.n43 VDD.t11 11.5766
R337 VDD.n3 VDD.t9 8.90522
R338 VDD.n24 VDD.n23 8.2255
R339 VDD.n48 VDD.n24 8.2255
R340 VDD VDD.n24 6.3005
R341 VDD VDD.n24 6.3005
R342 VDD.n25 VDD.t2 4.57285
R343 VDD.n9 VDD.t8 3.56239
R344 VDD.n26 VDD.t3 3.3285
R345 VDD.n25 VDD.t1 3.3285
R346 VDD.n1 VDD.n0 3.1505
R347 VDD.n5 VDD.n4 3.1505
R348 VDD.n4 VDD.n3 3.1505
R349 VDD.n8 VDD.n7 3.1505
R350 VDD.n7 VDD.n6 3.1505
R351 VDD.n11 VDD.n10 3.1505
R352 VDD.n10 VDD.n9 3.1505
R353 VDD.n14 VDD.n13 3.1505
R354 VDD.n13 VDD.n12 3.1505
R355 VDD.n17 VDD.n16 3.1505
R356 VDD.n16 VDD.n15 3.1505
R357 VDD.n20 VDD.n19 3.1505
R358 VDD.n19 VDD.n18 3.1505
R359 VDD.n23 VDD.n21 3.1505
R360 VDD.n23 VDD.n22 3.1505
R361 VDD.n46 VDD.n24 3.1505
R362 VDD.n49 VDD.n48 3.1505
R363 VDD.n48 VDD.n47 3.1505
R364 VDD.n45 VDD.n44 3.1505
R365 VDD.n44 VDD.n43 3.1505
R366 VDD.n42 VDD.n41 3.1505
R367 VDD.n41 VDD.n40 3.1505
R368 VDD.n39 VDD.n38 3.1505
R369 VDD.n38 VDD.n37 3.1505
R370 VDD.n36 VDD.n35 3.1505
R371 VDD.n35 VDD.n34 3.1505
R372 VDD.n33 VDD.n32 3.1505
R373 VDD.n32 VDD.n31 3.1505
R374 VDD.n30 VDD.n29 3.1505
R375 VDD.n2 VDD.n1 1.89487
R376 VDD.n26 VDD.n25 1.24485
R377 VDD.n27 VDD.n26 0.935717
R378 VDD.t6 VDD.n46 0.890972
R379 VDD.n5 VDD.n2 0.616836
R380 VDD.n29 VDD.n28 0.460561
R381 VDD.n8 VDD.n5 0.0760357
R382 VDD.n11 VDD.n8 0.0760357
R383 VDD.n14 VDD.n11 0.0760357
R384 VDD.n17 VDD.n14 0.0760357
R385 VDD.n20 VDD.n17 0.0760357
R386 VDD.n21 VDD.n20 0.0760357
R387 VDD VDD.n21 0.0760357
R388 VDD VDD.n49 0.0760357
R389 VDD.n49 VDD.n45 0.0760357
R390 VDD.n45 VDD.n42 0.0760357
R391 VDD.n42 VDD.n39 0.0760357
R392 VDD.n39 VDD.n36 0.0760357
R393 VDD.n36 VDD.n33 0.0760357
R394 VDD.n33 VDD.n30 0.0760357
R395 VDD.n30 VDD.n27 0.0262143
C0 CLK VOUT 0.319f
C1 VIN VDD 1.63f
C2 VIN VOUT 11.5f
C3 CLK VIN 0.334f
C4 VOUT VDD 0.171f
C5 CLK VDD 0.343f
.ends

