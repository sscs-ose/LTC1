magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -3099 -2045 3099 2045
<< psubdiff >>
rect -1099 23 1099 45
rect -1099 -23 -1077 23
rect -1031 -23 -953 23
rect -907 -23 -829 23
rect -783 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 783 23
rect 829 -23 907 23
rect 953 -23 1031 23
rect 1077 -23 1099 23
rect -1099 -45 1099 -23
<< psubdiffcont >>
rect -1077 -23 -1031 23
rect -953 -23 -907 23
rect -829 -23 -783 23
rect -705 -23 -659 23
rect -581 -23 -535 23
rect -457 -23 -411 23
rect -333 -23 -287 23
rect -209 -23 -163 23
rect -85 -23 -39 23
rect 39 -23 85 23
rect 163 -23 209 23
rect 287 -23 333 23
rect 411 -23 457 23
rect 535 -23 581 23
rect 659 -23 705 23
rect 783 -23 829 23
rect 907 -23 953 23
rect 1031 -23 1077 23
<< metal1 >>
rect -1088 23 1088 34
rect -1088 -23 -1077 23
rect -1031 -23 -953 23
rect -907 -23 -829 23
rect -783 -23 -705 23
rect -659 -23 -581 23
rect -535 -23 -457 23
rect -411 -23 -333 23
rect -287 -23 -209 23
rect -163 -23 -85 23
rect -39 -23 39 23
rect 85 -23 163 23
rect 209 -23 287 23
rect 333 -23 411 23
rect 457 -23 535 23
rect 581 -23 659 23
rect 705 -23 783 23
rect 829 -23 907 23
rect 953 -23 1031 23
rect 1077 -23 1088 23
rect -1088 -34 1088 -23
<< end >>
