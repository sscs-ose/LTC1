magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -14993 -2097 14993 2097
<< psubdiff >>
rect -12993 75 12993 97
rect -12993 29 -12971 75
rect -12925 29 -12867 75
rect -12821 29 -12763 75
rect -12717 29 -12659 75
rect -12613 29 -12555 75
rect -12509 29 -12451 75
rect -12405 29 -12347 75
rect -12301 29 -12243 75
rect -12197 29 -12139 75
rect -12093 29 -12035 75
rect -11989 29 -11931 75
rect -11885 29 -11827 75
rect -11781 29 -11723 75
rect -11677 29 -11619 75
rect -11573 29 -11515 75
rect -11469 29 -11411 75
rect -11365 29 -11307 75
rect -11261 29 -11203 75
rect -11157 29 -11099 75
rect -11053 29 -10995 75
rect -10949 29 -10891 75
rect -10845 29 -10787 75
rect -10741 29 -10683 75
rect -10637 29 -10579 75
rect -10533 29 -10475 75
rect -10429 29 -10371 75
rect -10325 29 -10267 75
rect -10221 29 -10163 75
rect -10117 29 -10059 75
rect -10013 29 -9955 75
rect -9909 29 -9851 75
rect -9805 29 -9747 75
rect -9701 29 -9643 75
rect -9597 29 -9539 75
rect -9493 29 -9435 75
rect -9389 29 -9331 75
rect -9285 29 -9227 75
rect -9181 29 -9123 75
rect -9077 29 -9019 75
rect -8973 29 -8915 75
rect -8869 29 -8811 75
rect -8765 29 -8707 75
rect -8661 29 -8603 75
rect -8557 29 -8499 75
rect -8453 29 -8395 75
rect -8349 29 -8291 75
rect -8245 29 -8187 75
rect -8141 29 -8083 75
rect -8037 29 -7979 75
rect -7933 29 -7875 75
rect -7829 29 -7771 75
rect -7725 29 -7667 75
rect -7621 29 -7563 75
rect -7517 29 -7459 75
rect -7413 29 -7355 75
rect -7309 29 -7251 75
rect -7205 29 -7147 75
rect -7101 29 -7043 75
rect -6997 29 -6939 75
rect -6893 29 -6835 75
rect -6789 29 -6731 75
rect -6685 29 -6627 75
rect -6581 29 -6523 75
rect -6477 29 -6419 75
rect -6373 29 -6315 75
rect -6269 29 -6211 75
rect -6165 29 -6107 75
rect -6061 29 -6003 75
rect -5957 29 -5899 75
rect -5853 29 -5795 75
rect -5749 29 -5691 75
rect -5645 29 -5587 75
rect -5541 29 -5483 75
rect -5437 29 -5379 75
rect -5333 29 -5275 75
rect -5229 29 -5171 75
rect -5125 29 -5067 75
rect -5021 29 -4963 75
rect -4917 29 -4859 75
rect -4813 29 -4755 75
rect -4709 29 -4651 75
rect -4605 29 -4547 75
rect -4501 29 -4443 75
rect -4397 29 -4339 75
rect -4293 29 -4235 75
rect -4189 29 -4131 75
rect -4085 29 -4027 75
rect -3981 29 -3923 75
rect -3877 29 -3819 75
rect -3773 29 -3715 75
rect -3669 29 -3611 75
rect -3565 29 -3507 75
rect -3461 29 -3403 75
rect -3357 29 -3299 75
rect -3253 29 -3195 75
rect -3149 29 -3091 75
rect -3045 29 -2987 75
rect -2941 29 -2883 75
rect -2837 29 -2779 75
rect -2733 29 -2675 75
rect -2629 29 -2571 75
rect -2525 29 -2467 75
rect -2421 29 -2363 75
rect -2317 29 -2259 75
rect -2213 29 -2155 75
rect -2109 29 -2051 75
rect -2005 29 -1947 75
rect -1901 29 -1843 75
rect -1797 29 -1739 75
rect -1693 29 -1635 75
rect -1589 29 -1531 75
rect -1485 29 -1427 75
rect -1381 29 -1323 75
rect -1277 29 -1219 75
rect -1173 29 -1115 75
rect -1069 29 -1011 75
rect -965 29 -907 75
rect -861 29 -803 75
rect -757 29 -699 75
rect -653 29 -595 75
rect -549 29 -491 75
rect -445 29 -387 75
rect -341 29 -283 75
rect -237 29 -179 75
rect -133 29 -75 75
rect -29 29 29 75
rect 75 29 133 75
rect 179 29 237 75
rect 283 29 341 75
rect 387 29 445 75
rect 491 29 549 75
rect 595 29 653 75
rect 699 29 757 75
rect 803 29 861 75
rect 907 29 965 75
rect 1011 29 1069 75
rect 1115 29 1173 75
rect 1219 29 1277 75
rect 1323 29 1381 75
rect 1427 29 1485 75
rect 1531 29 1589 75
rect 1635 29 1693 75
rect 1739 29 1797 75
rect 1843 29 1901 75
rect 1947 29 2005 75
rect 2051 29 2109 75
rect 2155 29 2213 75
rect 2259 29 2317 75
rect 2363 29 2421 75
rect 2467 29 2525 75
rect 2571 29 2629 75
rect 2675 29 2733 75
rect 2779 29 2837 75
rect 2883 29 2941 75
rect 2987 29 3045 75
rect 3091 29 3149 75
rect 3195 29 3253 75
rect 3299 29 3357 75
rect 3403 29 3461 75
rect 3507 29 3565 75
rect 3611 29 3669 75
rect 3715 29 3773 75
rect 3819 29 3877 75
rect 3923 29 3981 75
rect 4027 29 4085 75
rect 4131 29 4189 75
rect 4235 29 4293 75
rect 4339 29 4397 75
rect 4443 29 4501 75
rect 4547 29 4605 75
rect 4651 29 4709 75
rect 4755 29 4813 75
rect 4859 29 4917 75
rect 4963 29 5021 75
rect 5067 29 5125 75
rect 5171 29 5229 75
rect 5275 29 5333 75
rect 5379 29 5437 75
rect 5483 29 5541 75
rect 5587 29 5645 75
rect 5691 29 5749 75
rect 5795 29 5853 75
rect 5899 29 5957 75
rect 6003 29 6061 75
rect 6107 29 6165 75
rect 6211 29 6269 75
rect 6315 29 6373 75
rect 6419 29 6477 75
rect 6523 29 6581 75
rect 6627 29 6685 75
rect 6731 29 6789 75
rect 6835 29 6893 75
rect 6939 29 6997 75
rect 7043 29 7101 75
rect 7147 29 7205 75
rect 7251 29 7309 75
rect 7355 29 7413 75
rect 7459 29 7517 75
rect 7563 29 7621 75
rect 7667 29 7725 75
rect 7771 29 7829 75
rect 7875 29 7933 75
rect 7979 29 8037 75
rect 8083 29 8141 75
rect 8187 29 8245 75
rect 8291 29 8349 75
rect 8395 29 8453 75
rect 8499 29 8557 75
rect 8603 29 8661 75
rect 8707 29 8765 75
rect 8811 29 8869 75
rect 8915 29 8973 75
rect 9019 29 9077 75
rect 9123 29 9181 75
rect 9227 29 9285 75
rect 9331 29 9389 75
rect 9435 29 9493 75
rect 9539 29 9597 75
rect 9643 29 9701 75
rect 9747 29 9805 75
rect 9851 29 9909 75
rect 9955 29 10013 75
rect 10059 29 10117 75
rect 10163 29 10221 75
rect 10267 29 10325 75
rect 10371 29 10429 75
rect 10475 29 10533 75
rect 10579 29 10637 75
rect 10683 29 10741 75
rect 10787 29 10845 75
rect 10891 29 10949 75
rect 10995 29 11053 75
rect 11099 29 11157 75
rect 11203 29 11261 75
rect 11307 29 11365 75
rect 11411 29 11469 75
rect 11515 29 11573 75
rect 11619 29 11677 75
rect 11723 29 11781 75
rect 11827 29 11885 75
rect 11931 29 11989 75
rect 12035 29 12093 75
rect 12139 29 12197 75
rect 12243 29 12301 75
rect 12347 29 12405 75
rect 12451 29 12509 75
rect 12555 29 12613 75
rect 12659 29 12717 75
rect 12763 29 12821 75
rect 12867 29 12925 75
rect 12971 29 12993 75
rect -12993 -29 12993 29
rect -12993 -75 -12971 -29
rect -12925 -75 -12867 -29
rect -12821 -75 -12763 -29
rect -12717 -75 -12659 -29
rect -12613 -75 -12555 -29
rect -12509 -75 -12451 -29
rect -12405 -75 -12347 -29
rect -12301 -75 -12243 -29
rect -12197 -75 -12139 -29
rect -12093 -75 -12035 -29
rect -11989 -75 -11931 -29
rect -11885 -75 -11827 -29
rect -11781 -75 -11723 -29
rect -11677 -75 -11619 -29
rect -11573 -75 -11515 -29
rect -11469 -75 -11411 -29
rect -11365 -75 -11307 -29
rect -11261 -75 -11203 -29
rect -11157 -75 -11099 -29
rect -11053 -75 -10995 -29
rect -10949 -75 -10891 -29
rect -10845 -75 -10787 -29
rect -10741 -75 -10683 -29
rect -10637 -75 -10579 -29
rect -10533 -75 -10475 -29
rect -10429 -75 -10371 -29
rect -10325 -75 -10267 -29
rect -10221 -75 -10163 -29
rect -10117 -75 -10059 -29
rect -10013 -75 -9955 -29
rect -9909 -75 -9851 -29
rect -9805 -75 -9747 -29
rect -9701 -75 -9643 -29
rect -9597 -75 -9539 -29
rect -9493 -75 -9435 -29
rect -9389 -75 -9331 -29
rect -9285 -75 -9227 -29
rect -9181 -75 -9123 -29
rect -9077 -75 -9019 -29
rect -8973 -75 -8915 -29
rect -8869 -75 -8811 -29
rect -8765 -75 -8707 -29
rect -8661 -75 -8603 -29
rect -8557 -75 -8499 -29
rect -8453 -75 -8395 -29
rect -8349 -75 -8291 -29
rect -8245 -75 -8187 -29
rect -8141 -75 -8083 -29
rect -8037 -75 -7979 -29
rect -7933 -75 -7875 -29
rect -7829 -75 -7771 -29
rect -7725 -75 -7667 -29
rect -7621 -75 -7563 -29
rect -7517 -75 -7459 -29
rect -7413 -75 -7355 -29
rect -7309 -75 -7251 -29
rect -7205 -75 -7147 -29
rect -7101 -75 -7043 -29
rect -6997 -75 -6939 -29
rect -6893 -75 -6835 -29
rect -6789 -75 -6731 -29
rect -6685 -75 -6627 -29
rect -6581 -75 -6523 -29
rect -6477 -75 -6419 -29
rect -6373 -75 -6315 -29
rect -6269 -75 -6211 -29
rect -6165 -75 -6107 -29
rect -6061 -75 -6003 -29
rect -5957 -75 -5899 -29
rect -5853 -75 -5795 -29
rect -5749 -75 -5691 -29
rect -5645 -75 -5587 -29
rect -5541 -75 -5483 -29
rect -5437 -75 -5379 -29
rect -5333 -75 -5275 -29
rect -5229 -75 -5171 -29
rect -5125 -75 -5067 -29
rect -5021 -75 -4963 -29
rect -4917 -75 -4859 -29
rect -4813 -75 -4755 -29
rect -4709 -75 -4651 -29
rect -4605 -75 -4547 -29
rect -4501 -75 -4443 -29
rect -4397 -75 -4339 -29
rect -4293 -75 -4235 -29
rect -4189 -75 -4131 -29
rect -4085 -75 -4027 -29
rect -3981 -75 -3923 -29
rect -3877 -75 -3819 -29
rect -3773 -75 -3715 -29
rect -3669 -75 -3611 -29
rect -3565 -75 -3507 -29
rect -3461 -75 -3403 -29
rect -3357 -75 -3299 -29
rect -3253 -75 -3195 -29
rect -3149 -75 -3091 -29
rect -3045 -75 -2987 -29
rect -2941 -75 -2883 -29
rect -2837 -75 -2779 -29
rect -2733 -75 -2675 -29
rect -2629 -75 -2571 -29
rect -2525 -75 -2467 -29
rect -2421 -75 -2363 -29
rect -2317 -75 -2259 -29
rect -2213 -75 -2155 -29
rect -2109 -75 -2051 -29
rect -2005 -75 -1947 -29
rect -1901 -75 -1843 -29
rect -1797 -75 -1739 -29
rect -1693 -75 -1635 -29
rect -1589 -75 -1531 -29
rect -1485 -75 -1427 -29
rect -1381 -75 -1323 -29
rect -1277 -75 -1219 -29
rect -1173 -75 -1115 -29
rect -1069 -75 -1011 -29
rect -965 -75 -907 -29
rect -861 -75 -803 -29
rect -757 -75 -699 -29
rect -653 -75 -595 -29
rect -549 -75 -491 -29
rect -445 -75 -387 -29
rect -341 -75 -283 -29
rect -237 -75 -179 -29
rect -133 -75 -75 -29
rect -29 -75 29 -29
rect 75 -75 133 -29
rect 179 -75 237 -29
rect 283 -75 341 -29
rect 387 -75 445 -29
rect 491 -75 549 -29
rect 595 -75 653 -29
rect 699 -75 757 -29
rect 803 -75 861 -29
rect 907 -75 965 -29
rect 1011 -75 1069 -29
rect 1115 -75 1173 -29
rect 1219 -75 1277 -29
rect 1323 -75 1381 -29
rect 1427 -75 1485 -29
rect 1531 -75 1589 -29
rect 1635 -75 1693 -29
rect 1739 -75 1797 -29
rect 1843 -75 1901 -29
rect 1947 -75 2005 -29
rect 2051 -75 2109 -29
rect 2155 -75 2213 -29
rect 2259 -75 2317 -29
rect 2363 -75 2421 -29
rect 2467 -75 2525 -29
rect 2571 -75 2629 -29
rect 2675 -75 2733 -29
rect 2779 -75 2837 -29
rect 2883 -75 2941 -29
rect 2987 -75 3045 -29
rect 3091 -75 3149 -29
rect 3195 -75 3253 -29
rect 3299 -75 3357 -29
rect 3403 -75 3461 -29
rect 3507 -75 3565 -29
rect 3611 -75 3669 -29
rect 3715 -75 3773 -29
rect 3819 -75 3877 -29
rect 3923 -75 3981 -29
rect 4027 -75 4085 -29
rect 4131 -75 4189 -29
rect 4235 -75 4293 -29
rect 4339 -75 4397 -29
rect 4443 -75 4501 -29
rect 4547 -75 4605 -29
rect 4651 -75 4709 -29
rect 4755 -75 4813 -29
rect 4859 -75 4917 -29
rect 4963 -75 5021 -29
rect 5067 -75 5125 -29
rect 5171 -75 5229 -29
rect 5275 -75 5333 -29
rect 5379 -75 5437 -29
rect 5483 -75 5541 -29
rect 5587 -75 5645 -29
rect 5691 -75 5749 -29
rect 5795 -75 5853 -29
rect 5899 -75 5957 -29
rect 6003 -75 6061 -29
rect 6107 -75 6165 -29
rect 6211 -75 6269 -29
rect 6315 -75 6373 -29
rect 6419 -75 6477 -29
rect 6523 -75 6581 -29
rect 6627 -75 6685 -29
rect 6731 -75 6789 -29
rect 6835 -75 6893 -29
rect 6939 -75 6997 -29
rect 7043 -75 7101 -29
rect 7147 -75 7205 -29
rect 7251 -75 7309 -29
rect 7355 -75 7413 -29
rect 7459 -75 7517 -29
rect 7563 -75 7621 -29
rect 7667 -75 7725 -29
rect 7771 -75 7829 -29
rect 7875 -75 7933 -29
rect 7979 -75 8037 -29
rect 8083 -75 8141 -29
rect 8187 -75 8245 -29
rect 8291 -75 8349 -29
rect 8395 -75 8453 -29
rect 8499 -75 8557 -29
rect 8603 -75 8661 -29
rect 8707 -75 8765 -29
rect 8811 -75 8869 -29
rect 8915 -75 8973 -29
rect 9019 -75 9077 -29
rect 9123 -75 9181 -29
rect 9227 -75 9285 -29
rect 9331 -75 9389 -29
rect 9435 -75 9493 -29
rect 9539 -75 9597 -29
rect 9643 -75 9701 -29
rect 9747 -75 9805 -29
rect 9851 -75 9909 -29
rect 9955 -75 10013 -29
rect 10059 -75 10117 -29
rect 10163 -75 10221 -29
rect 10267 -75 10325 -29
rect 10371 -75 10429 -29
rect 10475 -75 10533 -29
rect 10579 -75 10637 -29
rect 10683 -75 10741 -29
rect 10787 -75 10845 -29
rect 10891 -75 10949 -29
rect 10995 -75 11053 -29
rect 11099 -75 11157 -29
rect 11203 -75 11261 -29
rect 11307 -75 11365 -29
rect 11411 -75 11469 -29
rect 11515 -75 11573 -29
rect 11619 -75 11677 -29
rect 11723 -75 11781 -29
rect 11827 -75 11885 -29
rect 11931 -75 11989 -29
rect 12035 -75 12093 -29
rect 12139 -75 12197 -29
rect 12243 -75 12301 -29
rect 12347 -75 12405 -29
rect 12451 -75 12509 -29
rect 12555 -75 12613 -29
rect 12659 -75 12717 -29
rect 12763 -75 12821 -29
rect 12867 -75 12925 -29
rect 12971 -75 12993 -29
rect -12993 -97 12993 -75
<< psubdiffcont >>
rect -12971 29 -12925 75
rect -12867 29 -12821 75
rect -12763 29 -12717 75
rect -12659 29 -12613 75
rect -12555 29 -12509 75
rect -12451 29 -12405 75
rect -12347 29 -12301 75
rect -12243 29 -12197 75
rect -12139 29 -12093 75
rect -12035 29 -11989 75
rect -11931 29 -11885 75
rect -11827 29 -11781 75
rect -11723 29 -11677 75
rect -11619 29 -11573 75
rect -11515 29 -11469 75
rect -11411 29 -11365 75
rect -11307 29 -11261 75
rect -11203 29 -11157 75
rect -11099 29 -11053 75
rect -10995 29 -10949 75
rect -10891 29 -10845 75
rect -10787 29 -10741 75
rect -10683 29 -10637 75
rect -10579 29 -10533 75
rect -10475 29 -10429 75
rect -10371 29 -10325 75
rect -10267 29 -10221 75
rect -10163 29 -10117 75
rect -10059 29 -10013 75
rect -9955 29 -9909 75
rect -9851 29 -9805 75
rect -9747 29 -9701 75
rect -9643 29 -9597 75
rect -9539 29 -9493 75
rect -9435 29 -9389 75
rect -9331 29 -9285 75
rect -9227 29 -9181 75
rect -9123 29 -9077 75
rect -9019 29 -8973 75
rect -8915 29 -8869 75
rect -8811 29 -8765 75
rect -8707 29 -8661 75
rect -8603 29 -8557 75
rect -8499 29 -8453 75
rect -8395 29 -8349 75
rect -8291 29 -8245 75
rect -8187 29 -8141 75
rect -8083 29 -8037 75
rect -7979 29 -7933 75
rect -7875 29 -7829 75
rect -7771 29 -7725 75
rect -7667 29 -7621 75
rect -7563 29 -7517 75
rect -7459 29 -7413 75
rect -7355 29 -7309 75
rect -7251 29 -7205 75
rect -7147 29 -7101 75
rect -7043 29 -6997 75
rect -6939 29 -6893 75
rect -6835 29 -6789 75
rect -6731 29 -6685 75
rect -6627 29 -6581 75
rect -6523 29 -6477 75
rect -6419 29 -6373 75
rect -6315 29 -6269 75
rect -6211 29 -6165 75
rect -6107 29 -6061 75
rect -6003 29 -5957 75
rect -5899 29 -5853 75
rect -5795 29 -5749 75
rect -5691 29 -5645 75
rect -5587 29 -5541 75
rect -5483 29 -5437 75
rect -5379 29 -5333 75
rect -5275 29 -5229 75
rect -5171 29 -5125 75
rect -5067 29 -5021 75
rect -4963 29 -4917 75
rect -4859 29 -4813 75
rect -4755 29 -4709 75
rect -4651 29 -4605 75
rect -4547 29 -4501 75
rect -4443 29 -4397 75
rect -4339 29 -4293 75
rect -4235 29 -4189 75
rect -4131 29 -4085 75
rect -4027 29 -3981 75
rect -3923 29 -3877 75
rect -3819 29 -3773 75
rect -3715 29 -3669 75
rect -3611 29 -3565 75
rect -3507 29 -3461 75
rect -3403 29 -3357 75
rect -3299 29 -3253 75
rect -3195 29 -3149 75
rect -3091 29 -3045 75
rect -2987 29 -2941 75
rect -2883 29 -2837 75
rect -2779 29 -2733 75
rect -2675 29 -2629 75
rect -2571 29 -2525 75
rect -2467 29 -2421 75
rect -2363 29 -2317 75
rect -2259 29 -2213 75
rect -2155 29 -2109 75
rect -2051 29 -2005 75
rect -1947 29 -1901 75
rect -1843 29 -1797 75
rect -1739 29 -1693 75
rect -1635 29 -1589 75
rect -1531 29 -1485 75
rect -1427 29 -1381 75
rect -1323 29 -1277 75
rect -1219 29 -1173 75
rect -1115 29 -1069 75
rect -1011 29 -965 75
rect -907 29 -861 75
rect -803 29 -757 75
rect -699 29 -653 75
rect -595 29 -549 75
rect -491 29 -445 75
rect -387 29 -341 75
rect -283 29 -237 75
rect -179 29 -133 75
rect -75 29 -29 75
rect 29 29 75 75
rect 133 29 179 75
rect 237 29 283 75
rect 341 29 387 75
rect 445 29 491 75
rect 549 29 595 75
rect 653 29 699 75
rect 757 29 803 75
rect 861 29 907 75
rect 965 29 1011 75
rect 1069 29 1115 75
rect 1173 29 1219 75
rect 1277 29 1323 75
rect 1381 29 1427 75
rect 1485 29 1531 75
rect 1589 29 1635 75
rect 1693 29 1739 75
rect 1797 29 1843 75
rect 1901 29 1947 75
rect 2005 29 2051 75
rect 2109 29 2155 75
rect 2213 29 2259 75
rect 2317 29 2363 75
rect 2421 29 2467 75
rect 2525 29 2571 75
rect 2629 29 2675 75
rect 2733 29 2779 75
rect 2837 29 2883 75
rect 2941 29 2987 75
rect 3045 29 3091 75
rect 3149 29 3195 75
rect 3253 29 3299 75
rect 3357 29 3403 75
rect 3461 29 3507 75
rect 3565 29 3611 75
rect 3669 29 3715 75
rect 3773 29 3819 75
rect 3877 29 3923 75
rect 3981 29 4027 75
rect 4085 29 4131 75
rect 4189 29 4235 75
rect 4293 29 4339 75
rect 4397 29 4443 75
rect 4501 29 4547 75
rect 4605 29 4651 75
rect 4709 29 4755 75
rect 4813 29 4859 75
rect 4917 29 4963 75
rect 5021 29 5067 75
rect 5125 29 5171 75
rect 5229 29 5275 75
rect 5333 29 5379 75
rect 5437 29 5483 75
rect 5541 29 5587 75
rect 5645 29 5691 75
rect 5749 29 5795 75
rect 5853 29 5899 75
rect 5957 29 6003 75
rect 6061 29 6107 75
rect 6165 29 6211 75
rect 6269 29 6315 75
rect 6373 29 6419 75
rect 6477 29 6523 75
rect 6581 29 6627 75
rect 6685 29 6731 75
rect 6789 29 6835 75
rect 6893 29 6939 75
rect 6997 29 7043 75
rect 7101 29 7147 75
rect 7205 29 7251 75
rect 7309 29 7355 75
rect 7413 29 7459 75
rect 7517 29 7563 75
rect 7621 29 7667 75
rect 7725 29 7771 75
rect 7829 29 7875 75
rect 7933 29 7979 75
rect 8037 29 8083 75
rect 8141 29 8187 75
rect 8245 29 8291 75
rect 8349 29 8395 75
rect 8453 29 8499 75
rect 8557 29 8603 75
rect 8661 29 8707 75
rect 8765 29 8811 75
rect 8869 29 8915 75
rect 8973 29 9019 75
rect 9077 29 9123 75
rect 9181 29 9227 75
rect 9285 29 9331 75
rect 9389 29 9435 75
rect 9493 29 9539 75
rect 9597 29 9643 75
rect 9701 29 9747 75
rect 9805 29 9851 75
rect 9909 29 9955 75
rect 10013 29 10059 75
rect 10117 29 10163 75
rect 10221 29 10267 75
rect 10325 29 10371 75
rect 10429 29 10475 75
rect 10533 29 10579 75
rect 10637 29 10683 75
rect 10741 29 10787 75
rect 10845 29 10891 75
rect 10949 29 10995 75
rect 11053 29 11099 75
rect 11157 29 11203 75
rect 11261 29 11307 75
rect 11365 29 11411 75
rect 11469 29 11515 75
rect 11573 29 11619 75
rect 11677 29 11723 75
rect 11781 29 11827 75
rect 11885 29 11931 75
rect 11989 29 12035 75
rect 12093 29 12139 75
rect 12197 29 12243 75
rect 12301 29 12347 75
rect 12405 29 12451 75
rect 12509 29 12555 75
rect 12613 29 12659 75
rect 12717 29 12763 75
rect 12821 29 12867 75
rect 12925 29 12971 75
rect -12971 -75 -12925 -29
rect -12867 -75 -12821 -29
rect -12763 -75 -12717 -29
rect -12659 -75 -12613 -29
rect -12555 -75 -12509 -29
rect -12451 -75 -12405 -29
rect -12347 -75 -12301 -29
rect -12243 -75 -12197 -29
rect -12139 -75 -12093 -29
rect -12035 -75 -11989 -29
rect -11931 -75 -11885 -29
rect -11827 -75 -11781 -29
rect -11723 -75 -11677 -29
rect -11619 -75 -11573 -29
rect -11515 -75 -11469 -29
rect -11411 -75 -11365 -29
rect -11307 -75 -11261 -29
rect -11203 -75 -11157 -29
rect -11099 -75 -11053 -29
rect -10995 -75 -10949 -29
rect -10891 -75 -10845 -29
rect -10787 -75 -10741 -29
rect -10683 -75 -10637 -29
rect -10579 -75 -10533 -29
rect -10475 -75 -10429 -29
rect -10371 -75 -10325 -29
rect -10267 -75 -10221 -29
rect -10163 -75 -10117 -29
rect -10059 -75 -10013 -29
rect -9955 -75 -9909 -29
rect -9851 -75 -9805 -29
rect -9747 -75 -9701 -29
rect -9643 -75 -9597 -29
rect -9539 -75 -9493 -29
rect -9435 -75 -9389 -29
rect -9331 -75 -9285 -29
rect -9227 -75 -9181 -29
rect -9123 -75 -9077 -29
rect -9019 -75 -8973 -29
rect -8915 -75 -8869 -29
rect -8811 -75 -8765 -29
rect -8707 -75 -8661 -29
rect -8603 -75 -8557 -29
rect -8499 -75 -8453 -29
rect -8395 -75 -8349 -29
rect -8291 -75 -8245 -29
rect -8187 -75 -8141 -29
rect -8083 -75 -8037 -29
rect -7979 -75 -7933 -29
rect -7875 -75 -7829 -29
rect -7771 -75 -7725 -29
rect -7667 -75 -7621 -29
rect -7563 -75 -7517 -29
rect -7459 -75 -7413 -29
rect -7355 -75 -7309 -29
rect -7251 -75 -7205 -29
rect -7147 -75 -7101 -29
rect -7043 -75 -6997 -29
rect -6939 -75 -6893 -29
rect -6835 -75 -6789 -29
rect -6731 -75 -6685 -29
rect -6627 -75 -6581 -29
rect -6523 -75 -6477 -29
rect -6419 -75 -6373 -29
rect -6315 -75 -6269 -29
rect -6211 -75 -6165 -29
rect -6107 -75 -6061 -29
rect -6003 -75 -5957 -29
rect -5899 -75 -5853 -29
rect -5795 -75 -5749 -29
rect -5691 -75 -5645 -29
rect -5587 -75 -5541 -29
rect -5483 -75 -5437 -29
rect -5379 -75 -5333 -29
rect -5275 -75 -5229 -29
rect -5171 -75 -5125 -29
rect -5067 -75 -5021 -29
rect -4963 -75 -4917 -29
rect -4859 -75 -4813 -29
rect -4755 -75 -4709 -29
rect -4651 -75 -4605 -29
rect -4547 -75 -4501 -29
rect -4443 -75 -4397 -29
rect -4339 -75 -4293 -29
rect -4235 -75 -4189 -29
rect -4131 -75 -4085 -29
rect -4027 -75 -3981 -29
rect -3923 -75 -3877 -29
rect -3819 -75 -3773 -29
rect -3715 -75 -3669 -29
rect -3611 -75 -3565 -29
rect -3507 -75 -3461 -29
rect -3403 -75 -3357 -29
rect -3299 -75 -3253 -29
rect -3195 -75 -3149 -29
rect -3091 -75 -3045 -29
rect -2987 -75 -2941 -29
rect -2883 -75 -2837 -29
rect -2779 -75 -2733 -29
rect -2675 -75 -2629 -29
rect -2571 -75 -2525 -29
rect -2467 -75 -2421 -29
rect -2363 -75 -2317 -29
rect -2259 -75 -2213 -29
rect -2155 -75 -2109 -29
rect -2051 -75 -2005 -29
rect -1947 -75 -1901 -29
rect -1843 -75 -1797 -29
rect -1739 -75 -1693 -29
rect -1635 -75 -1589 -29
rect -1531 -75 -1485 -29
rect -1427 -75 -1381 -29
rect -1323 -75 -1277 -29
rect -1219 -75 -1173 -29
rect -1115 -75 -1069 -29
rect -1011 -75 -965 -29
rect -907 -75 -861 -29
rect -803 -75 -757 -29
rect -699 -75 -653 -29
rect -595 -75 -549 -29
rect -491 -75 -445 -29
rect -387 -75 -341 -29
rect -283 -75 -237 -29
rect -179 -75 -133 -29
rect -75 -75 -29 -29
rect 29 -75 75 -29
rect 133 -75 179 -29
rect 237 -75 283 -29
rect 341 -75 387 -29
rect 445 -75 491 -29
rect 549 -75 595 -29
rect 653 -75 699 -29
rect 757 -75 803 -29
rect 861 -75 907 -29
rect 965 -75 1011 -29
rect 1069 -75 1115 -29
rect 1173 -75 1219 -29
rect 1277 -75 1323 -29
rect 1381 -75 1427 -29
rect 1485 -75 1531 -29
rect 1589 -75 1635 -29
rect 1693 -75 1739 -29
rect 1797 -75 1843 -29
rect 1901 -75 1947 -29
rect 2005 -75 2051 -29
rect 2109 -75 2155 -29
rect 2213 -75 2259 -29
rect 2317 -75 2363 -29
rect 2421 -75 2467 -29
rect 2525 -75 2571 -29
rect 2629 -75 2675 -29
rect 2733 -75 2779 -29
rect 2837 -75 2883 -29
rect 2941 -75 2987 -29
rect 3045 -75 3091 -29
rect 3149 -75 3195 -29
rect 3253 -75 3299 -29
rect 3357 -75 3403 -29
rect 3461 -75 3507 -29
rect 3565 -75 3611 -29
rect 3669 -75 3715 -29
rect 3773 -75 3819 -29
rect 3877 -75 3923 -29
rect 3981 -75 4027 -29
rect 4085 -75 4131 -29
rect 4189 -75 4235 -29
rect 4293 -75 4339 -29
rect 4397 -75 4443 -29
rect 4501 -75 4547 -29
rect 4605 -75 4651 -29
rect 4709 -75 4755 -29
rect 4813 -75 4859 -29
rect 4917 -75 4963 -29
rect 5021 -75 5067 -29
rect 5125 -75 5171 -29
rect 5229 -75 5275 -29
rect 5333 -75 5379 -29
rect 5437 -75 5483 -29
rect 5541 -75 5587 -29
rect 5645 -75 5691 -29
rect 5749 -75 5795 -29
rect 5853 -75 5899 -29
rect 5957 -75 6003 -29
rect 6061 -75 6107 -29
rect 6165 -75 6211 -29
rect 6269 -75 6315 -29
rect 6373 -75 6419 -29
rect 6477 -75 6523 -29
rect 6581 -75 6627 -29
rect 6685 -75 6731 -29
rect 6789 -75 6835 -29
rect 6893 -75 6939 -29
rect 6997 -75 7043 -29
rect 7101 -75 7147 -29
rect 7205 -75 7251 -29
rect 7309 -75 7355 -29
rect 7413 -75 7459 -29
rect 7517 -75 7563 -29
rect 7621 -75 7667 -29
rect 7725 -75 7771 -29
rect 7829 -75 7875 -29
rect 7933 -75 7979 -29
rect 8037 -75 8083 -29
rect 8141 -75 8187 -29
rect 8245 -75 8291 -29
rect 8349 -75 8395 -29
rect 8453 -75 8499 -29
rect 8557 -75 8603 -29
rect 8661 -75 8707 -29
rect 8765 -75 8811 -29
rect 8869 -75 8915 -29
rect 8973 -75 9019 -29
rect 9077 -75 9123 -29
rect 9181 -75 9227 -29
rect 9285 -75 9331 -29
rect 9389 -75 9435 -29
rect 9493 -75 9539 -29
rect 9597 -75 9643 -29
rect 9701 -75 9747 -29
rect 9805 -75 9851 -29
rect 9909 -75 9955 -29
rect 10013 -75 10059 -29
rect 10117 -75 10163 -29
rect 10221 -75 10267 -29
rect 10325 -75 10371 -29
rect 10429 -75 10475 -29
rect 10533 -75 10579 -29
rect 10637 -75 10683 -29
rect 10741 -75 10787 -29
rect 10845 -75 10891 -29
rect 10949 -75 10995 -29
rect 11053 -75 11099 -29
rect 11157 -75 11203 -29
rect 11261 -75 11307 -29
rect 11365 -75 11411 -29
rect 11469 -75 11515 -29
rect 11573 -75 11619 -29
rect 11677 -75 11723 -29
rect 11781 -75 11827 -29
rect 11885 -75 11931 -29
rect 11989 -75 12035 -29
rect 12093 -75 12139 -29
rect 12197 -75 12243 -29
rect 12301 -75 12347 -29
rect 12405 -75 12451 -29
rect 12509 -75 12555 -29
rect 12613 -75 12659 -29
rect 12717 -75 12763 -29
rect 12821 -75 12867 -29
rect 12925 -75 12971 -29
<< metal1 >>
rect -12982 75 12982 86
rect -12982 29 -12971 75
rect -12925 29 -12867 75
rect -12821 29 -12763 75
rect -12717 29 -12659 75
rect -12613 29 -12555 75
rect -12509 29 -12451 75
rect -12405 29 -12347 75
rect -12301 29 -12243 75
rect -12197 29 -12139 75
rect -12093 29 -12035 75
rect -11989 29 -11931 75
rect -11885 29 -11827 75
rect -11781 29 -11723 75
rect -11677 29 -11619 75
rect -11573 29 -11515 75
rect -11469 29 -11411 75
rect -11365 29 -11307 75
rect -11261 29 -11203 75
rect -11157 29 -11099 75
rect -11053 29 -10995 75
rect -10949 29 -10891 75
rect -10845 29 -10787 75
rect -10741 29 -10683 75
rect -10637 29 -10579 75
rect -10533 29 -10475 75
rect -10429 29 -10371 75
rect -10325 29 -10267 75
rect -10221 29 -10163 75
rect -10117 29 -10059 75
rect -10013 29 -9955 75
rect -9909 29 -9851 75
rect -9805 29 -9747 75
rect -9701 29 -9643 75
rect -9597 29 -9539 75
rect -9493 29 -9435 75
rect -9389 29 -9331 75
rect -9285 29 -9227 75
rect -9181 29 -9123 75
rect -9077 29 -9019 75
rect -8973 29 -8915 75
rect -8869 29 -8811 75
rect -8765 29 -8707 75
rect -8661 29 -8603 75
rect -8557 29 -8499 75
rect -8453 29 -8395 75
rect -8349 29 -8291 75
rect -8245 29 -8187 75
rect -8141 29 -8083 75
rect -8037 29 -7979 75
rect -7933 29 -7875 75
rect -7829 29 -7771 75
rect -7725 29 -7667 75
rect -7621 29 -7563 75
rect -7517 29 -7459 75
rect -7413 29 -7355 75
rect -7309 29 -7251 75
rect -7205 29 -7147 75
rect -7101 29 -7043 75
rect -6997 29 -6939 75
rect -6893 29 -6835 75
rect -6789 29 -6731 75
rect -6685 29 -6627 75
rect -6581 29 -6523 75
rect -6477 29 -6419 75
rect -6373 29 -6315 75
rect -6269 29 -6211 75
rect -6165 29 -6107 75
rect -6061 29 -6003 75
rect -5957 29 -5899 75
rect -5853 29 -5795 75
rect -5749 29 -5691 75
rect -5645 29 -5587 75
rect -5541 29 -5483 75
rect -5437 29 -5379 75
rect -5333 29 -5275 75
rect -5229 29 -5171 75
rect -5125 29 -5067 75
rect -5021 29 -4963 75
rect -4917 29 -4859 75
rect -4813 29 -4755 75
rect -4709 29 -4651 75
rect -4605 29 -4547 75
rect -4501 29 -4443 75
rect -4397 29 -4339 75
rect -4293 29 -4235 75
rect -4189 29 -4131 75
rect -4085 29 -4027 75
rect -3981 29 -3923 75
rect -3877 29 -3819 75
rect -3773 29 -3715 75
rect -3669 29 -3611 75
rect -3565 29 -3507 75
rect -3461 29 -3403 75
rect -3357 29 -3299 75
rect -3253 29 -3195 75
rect -3149 29 -3091 75
rect -3045 29 -2987 75
rect -2941 29 -2883 75
rect -2837 29 -2779 75
rect -2733 29 -2675 75
rect -2629 29 -2571 75
rect -2525 29 -2467 75
rect -2421 29 -2363 75
rect -2317 29 -2259 75
rect -2213 29 -2155 75
rect -2109 29 -2051 75
rect -2005 29 -1947 75
rect -1901 29 -1843 75
rect -1797 29 -1739 75
rect -1693 29 -1635 75
rect -1589 29 -1531 75
rect -1485 29 -1427 75
rect -1381 29 -1323 75
rect -1277 29 -1219 75
rect -1173 29 -1115 75
rect -1069 29 -1011 75
rect -965 29 -907 75
rect -861 29 -803 75
rect -757 29 -699 75
rect -653 29 -595 75
rect -549 29 -491 75
rect -445 29 -387 75
rect -341 29 -283 75
rect -237 29 -179 75
rect -133 29 -75 75
rect -29 29 29 75
rect 75 29 133 75
rect 179 29 237 75
rect 283 29 341 75
rect 387 29 445 75
rect 491 29 549 75
rect 595 29 653 75
rect 699 29 757 75
rect 803 29 861 75
rect 907 29 965 75
rect 1011 29 1069 75
rect 1115 29 1173 75
rect 1219 29 1277 75
rect 1323 29 1381 75
rect 1427 29 1485 75
rect 1531 29 1589 75
rect 1635 29 1693 75
rect 1739 29 1797 75
rect 1843 29 1901 75
rect 1947 29 2005 75
rect 2051 29 2109 75
rect 2155 29 2213 75
rect 2259 29 2317 75
rect 2363 29 2421 75
rect 2467 29 2525 75
rect 2571 29 2629 75
rect 2675 29 2733 75
rect 2779 29 2837 75
rect 2883 29 2941 75
rect 2987 29 3045 75
rect 3091 29 3149 75
rect 3195 29 3253 75
rect 3299 29 3357 75
rect 3403 29 3461 75
rect 3507 29 3565 75
rect 3611 29 3669 75
rect 3715 29 3773 75
rect 3819 29 3877 75
rect 3923 29 3981 75
rect 4027 29 4085 75
rect 4131 29 4189 75
rect 4235 29 4293 75
rect 4339 29 4397 75
rect 4443 29 4501 75
rect 4547 29 4605 75
rect 4651 29 4709 75
rect 4755 29 4813 75
rect 4859 29 4917 75
rect 4963 29 5021 75
rect 5067 29 5125 75
rect 5171 29 5229 75
rect 5275 29 5333 75
rect 5379 29 5437 75
rect 5483 29 5541 75
rect 5587 29 5645 75
rect 5691 29 5749 75
rect 5795 29 5853 75
rect 5899 29 5957 75
rect 6003 29 6061 75
rect 6107 29 6165 75
rect 6211 29 6269 75
rect 6315 29 6373 75
rect 6419 29 6477 75
rect 6523 29 6581 75
rect 6627 29 6685 75
rect 6731 29 6789 75
rect 6835 29 6893 75
rect 6939 29 6997 75
rect 7043 29 7101 75
rect 7147 29 7205 75
rect 7251 29 7309 75
rect 7355 29 7413 75
rect 7459 29 7517 75
rect 7563 29 7621 75
rect 7667 29 7725 75
rect 7771 29 7829 75
rect 7875 29 7933 75
rect 7979 29 8037 75
rect 8083 29 8141 75
rect 8187 29 8245 75
rect 8291 29 8349 75
rect 8395 29 8453 75
rect 8499 29 8557 75
rect 8603 29 8661 75
rect 8707 29 8765 75
rect 8811 29 8869 75
rect 8915 29 8973 75
rect 9019 29 9077 75
rect 9123 29 9181 75
rect 9227 29 9285 75
rect 9331 29 9389 75
rect 9435 29 9493 75
rect 9539 29 9597 75
rect 9643 29 9701 75
rect 9747 29 9805 75
rect 9851 29 9909 75
rect 9955 29 10013 75
rect 10059 29 10117 75
rect 10163 29 10221 75
rect 10267 29 10325 75
rect 10371 29 10429 75
rect 10475 29 10533 75
rect 10579 29 10637 75
rect 10683 29 10741 75
rect 10787 29 10845 75
rect 10891 29 10949 75
rect 10995 29 11053 75
rect 11099 29 11157 75
rect 11203 29 11261 75
rect 11307 29 11365 75
rect 11411 29 11469 75
rect 11515 29 11573 75
rect 11619 29 11677 75
rect 11723 29 11781 75
rect 11827 29 11885 75
rect 11931 29 11989 75
rect 12035 29 12093 75
rect 12139 29 12197 75
rect 12243 29 12301 75
rect 12347 29 12405 75
rect 12451 29 12509 75
rect 12555 29 12613 75
rect 12659 29 12717 75
rect 12763 29 12821 75
rect 12867 29 12925 75
rect 12971 29 12982 75
rect -12982 -29 12982 29
rect -12982 -75 -12971 -29
rect -12925 -75 -12867 -29
rect -12821 -75 -12763 -29
rect -12717 -75 -12659 -29
rect -12613 -75 -12555 -29
rect -12509 -75 -12451 -29
rect -12405 -75 -12347 -29
rect -12301 -75 -12243 -29
rect -12197 -75 -12139 -29
rect -12093 -75 -12035 -29
rect -11989 -75 -11931 -29
rect -11885 -75 -11827 -29
rect -11781 -75 -11723 -29
rect -11677 -75 -11619 -29
rect -11573 -75 -11515 -29
rect -11469 -75 -11411 -29
rect -11365 -75 -11307 -29
rect -11261 -75 -11203 -29
rect -11157 -75 -11099 -29
rect -11053 -75 -10995 -29
rect -10949 -75 -10891 -29
rect -10845 -75 -10787 -29
rect -10741 -75 -10683 -29
rect -10637 -75 -10579 -29
rect -10533 -75 -10475 -29
rect -10429 -75 -10371 -29
rect -10325 -75 -10267 -29
rect -10221 -75 -10163 -29
rect -10117 -75 -10059 -29
rect -10013 -75 -9955 -29
rect -9909 -75 -9851 -29
rect -9805 -75 -9747 -29
rect -9701 -75 -9643 -29
rect -9597 -75 -9539 -29
rect -9493 -75 -9435 -29
rect -9389 -75 -9331 -29
rect -9285 -75 -9227 -29
rect -9181 -75 -9123 -29
rect -9077 -75 -9019 -29
rect -8973 -75 -8915 -29
rect -8869 -75 -8811 -29
rect -8765 -75 -8707 -29
rect -8661 -75 -8603 -29
rect -8557 -75 -8499 -29
rect -8453 -75 -8395 -29
rect -8349 -75 -8291 -29
rect -8245 -75 -8187 -29
rect -8141 -75 -8083 -29
rect -8037 -75 -7979 -29
rect -7933 -75 -7875 -29
rect -7829 -75 -7771 -29
rect -7725 -75 -7667 -29
rect -7621 -75 -7563 -29
rect -7517 -75 -7459 -29
rect -7413 -75 -7355 -29
rect -7309 -75 -7251 -29
rect -7205 -75 -7147 -29
rect -7101 -75 -7043 -29
rect -6997 -75 -6939 -29
rect -6893 -75 -6835 -29
rect -6789 -75 -6731 -29
rect -6685 -75 -6627 -29
rect -6581 -75 -6523 -29
rect -6477 -75 -6419 -29
rect -6373 -75 -6315 -29
rect -6269 -75 -6211 -29
rect -6165 -75 -6107 -29
rect -6061 -75 -6003 -29
rect -5957 -75 -5899 -29
rect -5853 -75 -5795 -29
rect -5749 -75 -5691 -29
rect -5645 -75 -5587 -29
rect -5541 -75 -5483 -29
rect -5437 -75 -5379 -29
rect -5333 -75 -5275 -29
rect -5229 -75 -5171 -29
rect -5125 -75 -5067 -29
rect -5021 -75 -4963 -29
rect -4917 -75 -4859 -29
rect -4813 -75 -4755 -29
rect -4709 -75 -4651 -29
rect -4605 -75 -4547 -29
rect -4501 -75 -4443 -29
rect -4397 -75 -4339 -29
rect -4293 -75 -4235 -29
rect -4189 -75 -4131 -29
rect -4085 -75 -4027 -29
rect -3981 -75 -3923 -29
rect -3877 -75 -3819 -29
rect -3773 -75 -3715 -29
rect -3669 -75 -3611 -29
rect -3565 -75 -3507 -29
rect -3461 -75 -3403 -29
rect -3357 -75 -3299 -29
rect -3253 -75 -3195 -29
rect -3149 -75 -3091 -29
rect -3045 -75 -2987 -29
rect -2941 -75 -2883 -29
rect -2837 -75 -2779 -29
rect -2733 -75 -2675 -29
rect -2629 -75 -2571 -29
rect -2525 -75 -2467 -29
rect -2421 -75 -2363 -29
rect -2317 -75 -2259 -29
rect -2213 -75 -2155 -29
rect -2109 -75 -2051 -29
rect -2005 -75 -1947 -29
rect -1901 -75 -1843 -29
rect -1797 -75 -1739 -29
rect -1693 -75 -1635 -29
rect -1589 -75 -1531 -29
rect -1485 -75 -1427 -29
rect -1381 -75 -1323 -29
rect -1277 -75 -1219 -29
rect -1173 -75 -1115 -29
rect -1069 -75 -1011 -29
rect -965 -75 -907 -29
rect -861 -75 -803 -29
rect -757 -75 -699 -29
rect -653 -75 -595 -29
rect -549 -75 -491 -29
rect -445 -75 -387 -29
rect -341 -75 -283 -29
rect -237 -75 -179 -29
rect -133 -75 -75 -29
rect -29 -75 29 -29
rect 75 -75 133 -29
rect 179 -75 237 -29
rect 283 -75 341 -29
rect 387 -75 445 -29
rect 491 -75 549 -29
rect 595 -75 653 -29
rect 699 -75 757 -29
rect 803 -75 861 -29
rect 907 -75 965 -29
rect 1011 -75 1069 -29
rect 1115 -75 1173 -29
rect 1219 -75 1277 -29
rect 1323 -75 1381 -29
rect 1427 -75 1485 -29
rect 1531 -75 1589 -29
rect 1635 -75 1693 -29
rect 1739 -75 1797 -29
rect 1843 -75 1901 -29
rect 1947 -75 2005 -29
rect 2051 -75 2109 -29
rect 2155 -75 2213 -29
rect 2259 -75 2317 -29
rect 2363 -75 2421 -29
rect 2467 -75 2525 -29
rect 2571 -75 2629 -29
rect 2675 -75 2733 -29
rect 2779 -75 2837 -29
rect 2883 -75 2941 -29
rect 2987 -75 3045 -29
rect 3091 -75 3149 -29
rect 3195 -75 3253 -29
rect 3299 -75 3357 -29
rect 3403 -75 3461 -29
rect 3507 -75 3565 -29
rect 3611 -75 3669 -29
rect 3715 -75 3773 -29
rect 3819 -75 3877 -29
rect 3923 -75 3981 -29
rect 4027 -75 4085 -29
rect 4131 -75 4189 -29
rect 4235 -75 4293 -29
rect 4339 -75 4397 -29
rect 4443 -75 4501 -29
rect 4547 -75 4605 -29
rect 4651 -75 4709 -29
rect 4755 -75 4813 -29
rect 4859 -75 4917 -29
rect 4963 -75 5021 -29
rect 5067 -75 5125 -29
rect 5171 -75 5229 -29
rect 5275 -75 5333 -29
rect 5379 -75 5437 -29
rect 5483 -75 5541 -29
rect 5587 -75 5645 -29
rect 5691 -75 5749 -29
rect 5795 -75 5853 -29
rect 5899 -75 5957 -29
rect 6003 -75 6061 -29
rect 6107 -75 6165 -29
rect 6211 -75 6269 -29
rect 6315 -75 6373 -29
rect 6419 -75 6477 -29
rect 6523 -75 6581 -29
rect 6627 -75 6685 -29
rect 6731 -75 6789 -29
rect 6835 -75 6893 -29
rect 6939 -75 6997 -29
rect 7043 -75 7101 -29
rect 7147 -75 7205 -29
rect 7251 -75 7309 -29
rect 7355 -75 7413 -29
rect 7459 -75 7517 -29
rect 7563 -75 7621 -29
rect 7667 -75 7725 -29
rect 7771 -75 7829 -29
rect 7875 -75 7933 -29
rect 7979 -75 8037 -29
rect 8083 -75 8141 -29
rect 8187 -75 8245 -29
rect 8291 -75 8349 -29
rect 8395 -75 8453 -29
rect 8499 -75 8557 -29
rect 8603 -75 8661 -29
rect 8707 -75 8765 -29
rect 8811 -75 8869 -29
rect 8915 -75 8973 -29
rect 9019 -75 9077 -29
rect 9123 -75 9181 -29
rect 9227 -75 9285 -29
rect 9331 -75 9389 -29
rect 9435 -75 9493 -29
rect 9539 -75 9597 -29
rect 9643 -75 9701 -29
rect 9747 -75 9805 -29
rect 9851 -75 9909 -29
rect 9955 -75 10013 -29
rect 10059 -75 10117 -29
rect 10163 -75 10221 -29
rect 10267 -75 10325 -29
rect 10371 -75 10429 -29
rect 10475 -75 10533 -29
rect 10579 -75 10637 -29
rect 10683 -75 10741 -29
rect 10787 -75 10845 -29
rect 10891 -75 10949 -29
rect 10995 -75 11053 -29
rect 11099 -75 11157 -29
rect 11203 -75 11261 -29
rect 11307 -75 11365 -29
rect 11411 -75 11469 -29
rect 11515 -75 11573 -29
rect 11619 -75 11677 -29
rect 11723 -75 11781 -29
rect 11827 -75 11885 -29
rect 11931 -75 11989 -29
rect 12035 -75 12093 -29
rect 12139 -75 12197 -29
rect 12243 -75 12301 -29
rect 12347 -75 12405 -29
rect 12451 -75 12509 -29
rect 12555 -75 12613 -29
rect 12659 -75 12717 -29
rect 12763 -75 12821 -29
rect 12867 -75 12925 -29
rect 12971 -75 12982 -29
rect -12982 -86 12982 -75
<< end >>
