magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -906 33210 16833 58443
<< metal2 >>
rect 8733 41714 9612 52826
rect 13707 49592 13910 50992
rect 10638 47992 10996 49392
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_0
timestamp 1713338890
transform 1 0 14795 0 1 35896
box -38 -686 38 686
use M2_M1_CDNS_6903358316533  M2_M1_CDNS_6903358316533_1
timestamp 1713338890
transform 1 0 14795 0 1 50296
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_0
timestamp 1713338890
transform 1 0 14795 0 1 35896
box -38 -686 38 686
use M3_M2_CDNS_6903358316534  M3_M2_CDNS_6903358316534_1
timestamp 1713338890
transform 1 0 14795 0 1 50296
box -38 -686 38 686
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_0
timestamp 1713338890
transform 1 0 6892 0 1 35896
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_1
timestamp 1713338890
transform 1 0 8086 0 1 37496
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_2
timestamp 1713338890
transform 1 0 13376 0 1 35896
box -534 -658 534 658
use M3_M2_CDNS_69033583165370  M3_M2_CDNS_69033583165370_3
timestamp 1713338890
transform 1 0 13376 0 1 50290
box -534 -658 534 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_0
timestamp 1713338890
transform 1 0 9647 0 1 35896
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_1
timestamp 1713338890
transform 1 0 11575 0 1 37496
box -906 -658 906 658
use M3_M2_CDNS_69033583165373  M3_M2_CDNS_69033583165373_2
timestamp 1713338890
transform 1 0 11575 0 1 48698
box -906 -658 906 658
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_0
timestamp 1713338890
transform 1 0 2555 0 1 38371
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_1
timestamp 1713338890
transform 1 0 2927 0 1 37999
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_2
timestamp 1713338890
transform 1 0 2803 0 1 38123
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_3
timestamp 1713338890
transform 1 0 2679 0 1 38247
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_4
timestamp 1713338890
transform 1 0 3299 0 1 37627
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_5
timestamp 1713338890
transform 1 0 3795 0 1 37131
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_6
timestamp 1713338890
transform 1 0 3671 0 1 37255
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_7
timestamp 1713338890
transform 1 0 3547 0 1 37379
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_8
timestamp 1713338890
transform 1 0 3423 0 1 37503
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_9
timestamp 1713338890
transform 1 0 3919 0 1 37007
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_10
timestamp 1713338890
transform 1 0 4043 0 1 36883
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_11
timestamp 1713338890
transform 1 0 4167 0 1 36759
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_12
timestamp 1713338890
transform 1 0 3051 0 1 37875
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_13
timestamp 1713338890
transform 1 0 3175 0 1 37751
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_14
timestamp 1713338890
transform 1 0 4498 0 1 38690
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_15
timestamp 1713338890
transform 1 0 4746 0 1 38442
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_16
timestamp 1713338890
transform 1 0 4622 0 1 38566
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_17
timestamp 1713338890
transform 1 0 5490 0 1 37698
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_18
timestamp 1713338890
transform 1 0 5242 0 1 37946
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_19
timestamp 1713338890
transform 1 0 5366 0 1 37822
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_20
timestamp 1713338890
transform 1 0 5118 0 1 38070
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_21
timestamp 1713338890
transform 1 0 4994 0 1 38194
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_22
timestamp 1713338890
transform 1 0 4870 0 1 38318
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_23
timestamp 1713338890
transform 1 0 1132 0 1 42056
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_24
timestamp 1713338890
transform 1 0 2000 0 1 41188
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_25
timestamp 1713338890
transform 1 0 1876 0 1 41312
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_26
timestamp 1713338890
transform 1 0 1752 0 1 41436
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_27
timestamp 1713338890
transform 1 0 1628 0 1 41560
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_28
timestamp 1713338890
transform 1 0 1504 0 1 41684
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_29
timestamp 1713338890
transform 1 0 1380 0 1 41808
box -38 -844 38 844
use M3_M2_CDNS_69033583165374  M3_M2_CDNS_69033583165374_30
timestamp 1713338890
transform 1 0 1256 0 1 41932
box -38 -844 38 844
use M3_M2_CDNS_69033583165375  M3_M2_CDNS_69033583165375_0
timestamp 1713338890
transform 1 0 6110 0 1 37492
box -38 -658 38 658
use M3_M2_CDNS_69033583165375  M3_M2_CDNS_69033583165375_1
timestamp 1713338890
transform 1 0 5986 0 1 37493
box -38 -658 38 658
use M3_M2_CDNS_69033583165375  M3_M2_CDNS_69033583165375_2
timestamp 1713338890
transform 1 0 5862 0 1 37514
box -38 -658 38 658
use M3_M2_CDNS_69033583165376  M3_M2_CDNS_69033583165376_0
timestamp 1713338890
transform 1 0 5614 0 1 37630
box -38 -782 38 782
use M3_M2_CDNS_69033583165377  M3_M2_CDNS_69033583165377_0
timestamp 1713338890
transform 1 0 5738 0 1 37563
box -38 -720 38 720
use M3_M2_CDNS_69033583165385  M3_M2_CDNS_69033583165385_0
timestamp 1713338890
transform 1 0 9150 0 1 52151
box -348 -596 348 596
use M3_M2_CDNS_69033583165386  M3_M2_CDNS_69033583165386_0
timestamp 1713338890
transform 1 0 8050 0 1 50990
box -410 -472 410 472
use M3_M2_CDNS_69033583165387  M3_M2_CDNS_69033583165387_0
timestamp 1713338890
transform 1 0 8050 0 1 54607
box -410 -1836 410 1836
use M3_M2_CDNS_69033583165388  M3_M2_CDNS_69033583165388_0
timestamp 1713338890
transform 1 0 6592 0 1 54844
box -410 -1588 410 1588
<< end >>
