magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1445 -1019 1445 1019
<< metal2 >>
rect -445 14 445 19
rect -445 -14 -440 14
rect -412 -14 -369 14
rect -341 -14 -298 14
rect -270 -14 -227 14
rect -199 -14 -156 14
rect -128 -14 -85 14
rect -57 -14 -14 14
rect 14 -14 57 14
rect 85 -14 128 14
rect 156 -14 199 14
rect 227 -14 270 14
rect 298 -14 341 14
rect 369 -14 412 14
rect 440 -14 445 14
rect -445 -19 445 -14
<< via2 >>
rect -440 -14 -412 14
rect -369 -14 -341 14
rect -298 -14 -270 14
rect -227 -14 -199 14
rect -156 -14 -128 14
rect -85 -14 -57 14
rect -14 -14 14 14
rect 57 -14 85 14
rect 128 -14 156 14
rect 199 -14 227 14
rect 270 -14 298 14
rect 341 -14 369 14
rect 412 -14 440 14
<< metal3 >>
rect -445 14 445 19
rect -445 -14 -440 14
rect -412 -14 -369 14
rect -341 -14 -298 14
rect -270 -14 -227 14
rect -199 -14 -156 14
rect -128 -14 -85 14
rect -57 -14 -14 14
rect 14 -14 57 14
rect 85 -14 128 14
rect 156 -14 199 14
rect 227 -14 270 14
rect 298 -14 341 14
rect 369 -14 412 14
rect 440 -14 445 14
rect -445 -19 445 -14
<< end >>
