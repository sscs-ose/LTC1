** sch_path: /home/shahid/GF180Projects/mux/Xschem/2x1_mux.sch
**.subckt 2x1_mux VDD VSS Sel OUT I0 I1
*.iopin VDD
*.iopin VSS
*.ipin Sel
*.opin OUT
*.ipin I0
*.ipin I1
x1 net2 VSS VDD OUT net3 NAND
x2 Sel VSS VDD net3 I1 NAND
x3 I0 VSS VDD net2 net1 NAND
x4 VSS Sel net1 VDD inv_my
**.ends

* expanding   symbol:  NAND.sym # of pins=5
** sym_path: /home/shahid/GF180Projects/mux/Xschem/NAND.sym
** sch_path: /home/shahid/GF180Projects/mux/Xschem/NAND.sch
.subckt NAND IN1 VSS VDD OUT IN2
*.ipin IN2
*.ipin IN1
*.iopin VSS
*.iopin VDD
*.opin OUT
XM3 net1 IN2 VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM4 OUT IN1 net1 VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM5 OUT IN1 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN2 VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  inv_my.sym # of pins=4
** sym_path: /home/shahid/GF180Projects/mux/Xschem/inv_my.sym
** sch_path: /home/shahid/GF180Projects/mux/Xschem/inv_my.sch
.subckt inv_my VSS IN OUT VDD
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
XM1 OUT IN VSS VSS nfet_03v3 L=0.28u W=0.22u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pfet_03v3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.end
