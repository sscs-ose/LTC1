magic
tech gf180mcuC
magscale 1 10
timestamp 1697622990
<< nwell >>
rect 8578 11491 8995 11493
rect 8561 11488 8995 11491
<< metal1 >>
rect 18808 63061 19203 63067
rect -3079 62802 -2804 62816
rect -3079 62742 -3054 62802
rect -2994 62800 -2804 62802
rect -2994 62742 -2890 62800
rect -3079 62740 -2890 62742
rect -2830 62740 -2804 62800
rect -3079 62688 -2804 62740
rect -3079 62677 -2888 62688
rect -3390 62675 -2888 62677
rect -3390 62615 -3054 62675
rect -2994 62628 -2888 62675
rect -2828 62628 -2804 62688
rect -2994 62615 -2804 62628
rect -3390 62549 -2804 62615
rect -3079 62548 -2804 62549
rect -3079 62537 -2883 62548
rect -3079 62477 -3054 62537
rect -2994 62488 -2883 62537
rect -2823 62488 -2804 62548
rect -2994 62477 -2804 62488
rect -3079 62466 -2804 62477
rect -1982 62677 19203 63061
rect -4059 61402 -3689 61414
rect -4411 61374 -3689 61402
rect -4411 61361 -3847 61374
rect -4411 61301 -4013 61361
rect -3953 61314 -3847 61361
rect -3787 61314 -3689 61374
rect -3953 61301 -3689 61314
rect -4411 61237 -3689 61301
rect -4059 61234 -3689 61237
rect -4059 61223 -3842 61234
rect -4059 61163 -4013 61223
rect -3953 61174 -3842 61223
rect -3782 61174 -3689 61234
rect -3953 61163 -3689 61174
rect -4059 61136 -3689 61163
rect -2698 52730 -2423 52744
rect -2698 52670 -2673 52730
rect -2613 52728 -2423 52730
rect -2613 52670 -2509 52728
rect -2698 52668 -2509 52670
rect -2449 52668 -2423 52728
rect -2698 52639 -2423 52668
rect -3477 52616 -2423 52639
rect -3477 52603 -2507 52616
rect -3477 52543 -2673 52603
rect -2613 52556 -2507 52603
rect -2447 52556 -2423 52616
rect -2613 52543 -2423 52556
rect -3477 52491 -2423 52543
rect -2698 52476 -2423 52491
rect -2698 52465 -2502 52476
rect -2698 52405 -2673 52465
rect -2613 52416 -2502 52465
rect -2442 52416 -2423 52476
rect -2613 52405 -2423 52416
rect -2698 52394 -2423 52405
rect -3907 52246 -3537 52258
rect -4131 52218 -3537 52246
rect -4131 52205 -3695 52218
rect -4131 52145 -3861 52205
rect -3801 52158 -3695 52205
rect -3635 52158 -3537 52218
rect -3801 52145 -3537 52158
rect -4131 52081 -3537 52145
rect -3907 52078 -3537 52081
rect -3907 52067 -3690 52078
rect -3907 52007 -3861 52067
rect -3801 52018 -3690 52067
rect -3630 52018 -3537 52078
rect -3801 52007 -3537 52018
rect -3907 51980 -3537 52007
rect -2388 44204 -2113 44218
rect -2388 44144 -2363 44204
rect -2303 44202 -2113 44204
rect -2303 44144 -2199 44202
rect -2388 44142 -2199 44144
rect -2139 44142 -2113 44202
rect -2388 44090 -2113 44142
rect -2388 44077 -2197 44090
rect -2388 44073 -2363 44077
rect -3246 44017 -2363 44073
rect -2303 44030 -2197 44077
rect -2137 44030 -2113 44090
rect -2303 44017 -2113 44030
rect -3246 43950 -2113 44017
rect -3246 43939 -2192 43950
rect -3246 43925 -2363 43939
rect -2388 43879 -2363 43925
rect -2303 43890 -2192 43939
rect -2132 43890 -2113 43950
rect -2303 43879 -2113 43890
rect -2388 43868 -2113 43879
rect -2381 43663 -2106 43677
rect -2381 43603 -2356 43663
rect -2296 43661 -2106 43663
rect -2296 43603 -2192 43661
rect -2381 43601 -2192 43603
rect -2132 43601 -2106 43661
rect -2381 43549 -2106 43601
rect -2381 43547 -2190 43549
rect -3246 43536 -2190 43547
rect -3246 43476 -2356 43536
rect -2296 43489 -2190 43536
rect -2130 43489 -2106 43549
rect -2296 43476 -2106 43489
rect -3246 43409 -2106 43476
rect -3246 43399 -2185 43409
rect -2381 43398 -2185 43399
rect -2381 43338 -2356 43398
rect -2296 43349 -2185 43398
rect -2125 43349 -2106 43409
rect -2296 43338 -2106 43349
rect -2381 43327 -2106 43338
rect -2489 36770 -2214 36784
rect -2489 36710 -2464 36770
rect -2404 36768 -2214 36770
rect -2404 36710 -2300 36768
rect -2489 36708 -2300 36710
rect -2240 36708 -2214 36768
rect -2489 36680 -2214 36708
rect -3157 36656 -2214 36680
rect -3157 36643 -2298 36656
rect -3157 36583 -2464 36643
rect -2404 36596 -2298 36643
rect -2238 36596 -2214 36656
rect -2404 36583 -2214 36596
rect -3157 36532 -2214 36583
rect -2489 36516 -2214 36532
rect -2489 36505 -2293 36516
rect -2489 36445 -2464 36505
rect -2404 36456 -2293 36505
rect -2233 36456 -2214 36516
rect -2404 36445 -2214 36456
rect -2489 36434 -2214 36445
rect -3588 25044 -3261 25051
rect -3588 24984 -3575 25044
rect -3515 24984 -3455 25044
rect -3395 24984 -3335 25044
rect -3275 24984 -3261 25044
rect -3588 24965 -3261 24984
rect -3896 24924 -3261 24965
rect -3896 24864 -3575 24924
rect -3515 24864 -3455 24924
rect -3395 24864 -3335 24924
rect -3275 24864 -3261 24924
rect -3896 24824 -3261 24864
rect -3588 24804 -3261 24824
rect -3588 24744 -3575 24804
rect -3515 24744 -3455 24804
rect -3395 24744 -3335 24804
rect -3275 24744 -3261 24804
rect -3588 24732 -3261 24744
rect -1982 24212 -1598 62677
rect -734 55462 -180 55520
rect 4523 55463 5059 55511
rect 2762 54729 2988 54776
rect 8386 54369 8903 54424
rect -1113 48238 -1066 48601
rect 7285 41464 7336 42465
rect 7526 40566 7997 40618
rect 61 39776 236 39866
rect 4351 39720 4955 39766
rect 2010 28029 2740 28118
rect 2010 28021 2605 28029
rect 2010 27961 2039 28021
rect 2099 28018 2415 28021
rect 2099 27961 2218 28018
rect 2010 27958 2218 27961
rect 2278 27961 2415 28018
rect 2475 27969 2605 28021
rect 2665 27969 2740 28029
rect 2475 27961 2740 27969
rect 2278 27958 2740 27961
rect 2010 27894 2740 27958
rect 2010 27834 2042 27894
rect 2102 27886 2605 27894
rect 2102 27883 2407 27886
rect 2102 27834 2218 27883
rect 2010 27823 2218 27834
rect 2278 27826 2407 27883
rect 2467 27834 2605 27886
rect 2665 27834 2740 27894
rect 2467 27826 2740 27834
rect 2278 27823 2740 27826
rect 2010 27720 2740 27823
rect 5020 26011 5999 26363
rect -1982 24059 -1230 24212
rect -1982 23938 -1598 24059
rect -1383 23938 -1230 24059
rect -1982 23785 -806 23938
rect -1982 22452 -1598 23785
rect 5647 23168 5999 26011
rect 2715 22816 11131 23168
rect 18808 22570 19203 62677
rect 18790 22452 19220 22570
rect -1982 22068 19220 22452
rect 18790 21990 19220 22068
rect 9800 17600 10310 17660
rect 9800 17540 9832 17600
rect 9892 17540 9960 17600
rect 10020 17597 10310 17600
rect 10020 17540 10111 17597
rect 9800 17537 10111 17540
rect 10171 17537 10310 17597
rect 9800 17482 10310 17537
rect 7638 17441 10310 17482
rect 7638 17381 9830 17441
rect 9890 17439 10177 17441
rect 9890 17381 10001 17439
rect 7638 17379 10001 17381
rect 10061 17381 10177 17439
rect 10237 17381 10310 17441
rect 10061 17379 10310 17381
rect 7638 17338 10310 17379
rect 7638 16685 7782 17338
rect 9800 17278 10310 17338
rect 9800 17262 10193 17278
rect 9800 17257 10044 17262
rect 9800 17197 9842 17257
rect 9902 17202 10044 17257
rect 10104 17218 10193 17262
rect 10253 17218 10310 17278
rect 10104 17202 10310 17218
rect 9902 17197 10310 17202
rect 9800 17160 10310 17197
rect 13355 17337 25065 18084
rect 4098 16541 7782 16685
rect 9750 16937 10260 16990
rect 9750 16930 10050 16937
rect 9750 16927 9919 16930
rect 9750 16867 9791 16927
rect 9851 16870 9919 16927
rect 9979 16877 10050 16930
rect 10110 16877 10260 16937
rect 9979 16870 10260 16877
rect 9851 16867 10260 16870
rect 9750 16753 10260 16867
rect 9750 16748 10103 16753
rect 9750 16730 9955 16748
rect 9750 16670 9786 16730
rect 9846 16688 9955 16730
rect 10015 16693 10103 16748
rect 10163 16693 10260 16753
rect 10015 16688 10260 16693
rect 9846 16670 10260 16688
rect 9750 16620 10260 16670
rect 9750 16610 10137 16620
rect 9750 16579 9960 16610
rect 9750 16519 9763 16579
rect 9823 16550 9960 16579
rect 10020 16560 10137 16610
rect 10197 16560 10260 16620
rect 10020 16550 10260 16560
rect 9823 16519 10260 16550
rect 9750 16490 10260 16519
rect 1520 15970 1593 16058
rect 1320 15880 1398 15964
rect 1740 15510 1998 15563
rect 1863 15507 1996 15510
rect 9778 15355 9980 16490
rect 1530 15295 2126 15296
rect 1530 15240 2128 15295
rect 1532 15239 2128 15240
rect 3928 15153 9980 15355
rect 11733 14403 11992 14405
rect 2167 13969 7519 14172
rect 5930 11533 6133 13969
rect 6482 11515 6685 13969
rect 7316 11533 7519 13969
rect 9781 13966 11992 14403
rect 9781 11862 10218 13966
rect 11532 13843 11992 13966
rect 13355 13958 14102 17337
rect 22731 16830 23374 16880
rect 22731 16802 22811 16830
rect 22672 16770 22811 16802
rect 22871 16770 22931 16830
rect 22991 16770 23051 16830
rect 23111 16770 23171 16830
rect 23231 16770 23291 16830
rect 23351 16770 23374 16830
rect 22672 16710 23374 16770
rect 22672 16650 22811 16710
rect 22871 16650 22931 16710
rect 22991 16650 23051 16710
rect 23111 16650 23171 16710
rect 23231 16650 23291 16710
rect 23351 16650 23374 16710
rect 22672 16626 23374 16650
rect 22731 16591 23374 16626
rect 22735 16435 23393 16495
rect 22735 16430 22818 16435
rect 22669 16375 22818 16430
rect 22878 16375 22938 16435
rect 22998 16375 23058 16435
rect 23118 16375 23178 16435
rect 23238 16375 23298 16435
rect 23358 16375 23393 16435
rect 22669 16315 23393 16375
rect 22669 16255 22818 16315
rect 22878 16255 22938 16315
rect 22998 16255 23058 16315
rect 23118 16255 23178 16315
rect 23238 16255 23298 16315
rect 23358 16255 23393 16315
rect 22669 16232 23393 16255
rect 22735 16213 23393 16232
rect 22738 16210 23393 16213
rect 24318 16043 25065 17337
rect 55673 16043 56135 16047
rect 24318 15847 67173 16043
rect 67680 15847 88740 15857
rect 24318 15482 88740 15847
rect 24318 15472 68127 15482
rect 24318 15296 67173 15472
rect 22079 15270 22652 15272
rect 21918 15254 22652 15270
rect 21918 15194 22090 15254
rect 22150 15194 22210 15254
rect 22270 15194 22330 15254
rect 22390 15194 22450 15254
rect 22510 15194 22570 15254
rect 22630 15194 22652 15254
rect 21918 15134 22652 15194
rect 21918 15074 22090 15134
rect 22150 15074 22210 15134
rect 22270 15074 22330 15134
rect 22390 15074 22450 15134
rect 22510 15074 22570 15134
rect 22630 15074 22652 15134
rect 21918 15051 22652 15074
rect 21918 15049 22491 15051
rect 55490 14890 56420 15296
rect 22045 14662 22661 14694
rect 21999 14636 22694 14662
rect 21999 14576 22059 14636
rect 22119 14576 22179 14636
rect 22239 14576 22299 14636
rect 22359 14576 22419 14636
rect 22479 14576 22539 14636
rect 22599 14576 22694 14636
rect 21999 14516 22694 14576
rect 21999 14470 22059 14516
rect 17927 14293 18154 14470
rect 22045 14456 22059 14470
rect 22119 14456 22179 14516
rect 22239 14456 22299 14516
rect 22359 14456 22419 14516
rect 22479 14456 22539 14516
rect 22599 14470 22694 14516
rect 22599 14456 22661 14470
rect 22045 14427 22661 14456
rect 17890 14268 18200 14293
rect 17890 14216 17931 14268
rect 17983 14216 18035 14268
rect 18087 14216 18139 14268
rect 18191 14216 18200 14268
rect 17890 14164 18200 14216
rect 19228 14168 19380 14254
rect 17890 14112 17931 14164
rect 17983 14112 18035 14164
rect 18087 14112 18139 14164
rect 18191 14112 18200 14164
rect 17890 14060 18200 14112
rect 17890 14008 17931 14060
rect 17983 14008 18035 14060
rect 18087 14008 18139 14060
rect 18191 14008 18200 14060
rect 10844 13451 11116 13516
rect 10844 13397 10855 13451
rect 10913 13397 10993 13451
rect 11051 13397 11116 13451
rect 10844 13324 11116 13397
rect 10844 13270 10858 13324
rect 10916 13322 11116 13324
rect 10916 13270 10997 13322
rect 10844 13268 10997 13270
rect 11055 13268 11116 13322
rect 10844 13252 11116 13268
rect 10844 13212 11222 13252
rect 12351 13241 12512 13253
rect 10844 13180 11335 13212
rect 12222 13195 12512 13241
rect 12351 13184 12512 13195
rect 10844 13171 10997 13180
rect 10844 13117 10857 13171
rect 10915 13126 10997 13171
rect 11055 13140 11335 13180
rect 11055 13126 11222 13140
rect 10915 13117 11222 13126
rect 10844 13100 11222 13117
rect 11365 12710 11683 12801
rect 11365 12650 11397 12710
rect 11457 12707 11683 12710
rect 11457 12650 11581 12707
rect 11365 12647 11581 12650
rect 11641 12647 11683 12707
rect 11365 12582 11683 12647
rect 11365 12522 11394 12582
rect 11454 12574 11683 12582
rect 11454 12522 11579 12574
rect 11365 12514 11579 12522
rect 11639 12514 11683 12574
rect 11365 12437 11683 12514
rect 12387 12469 12512 13184
rect 11365 12377 11395 12437
rect 11455 12377 11572 12437
rect 11632 12377 11683 12437
rect 11365 12334 11683 12377
rect 12257 12416 12529 12469
rect 12257 12362 12268 12416
rect 12326 12362 12406 12416
rect 12464 12362 12529 12416
rect 12257 12289 12529 12362
rect 12257 12235 12271 12289
rect 12329 12287 12529 12289
rect 12329 12235 12410 12287
rect 12257 12233 12410 12235
rect 12468 12233 12529 12287
rect 12257 12217 12529 12233
rect 12257 12145 12533 12217
rect 12257 12136 12410 12145
rect 12257 12082 12270 12136
rect 12328 12091 12410 12136
rect 12468 12091 12533 12145
rect 12328 12082 12533 12091
rect 12257 12065 12533 12082
rect 8578 11669 8995 11731
rect 8578 11666 8872 11669
rect 8578 11665 8727 11666
rect 8578 11605 8605 11665
rect 8665 11606 8727 11665
rect 8787 11609 8872 11666
rect 8932 11609 8995 11669
rect 8787 11606 8995 11609
rect 8665 11605 8995 11606
rect 8578 11554 8995 11605
rect 9781 11564 12433 11862
rect 8578 11553 8742 11554
rect 8578 11493 8611 11553
rect 8671 11494 8742 11553
rect 8802 11494 8881 11554
rect 8941 11494 8995 11554
rect 8671 11493 8995 11494
rect 8578 11491 8995 11493
rect 9959 11492 12433 11564
rect 8561 11488 8995 11491
rect 1646 10690 2266 10779
rect 2407 10345 2529 10437
rect -63 7610 319 10120
rect 11236 9994 11632 10070
rect 11236 9983 11517 9994
rect 11236 9923 11340 9983
rect 11400 9934 11517 9983
rect 11577 9934 11632 9994
rect 11400 9923 11632 9934
rect 11236 9862 11632 9923
rect 11236 9852 11410 9862
rect 11236 9792 11274 9852
rect 11334 9802 11410 9852
rect 11470 9857 11632 9862
rect 11470 9802 11557 9857
rect 11334 9797 11557 9802
rect 11617 9797 11632 9857
rect 11334 9792 11632 9797
rect 11236 9772 11632 9792
rect 4086 9217 5247 9311
rect 12063 8509 12433 11492
rect 11423 7986 11671 8029
rect 11423 7926 11436 7986
rect 11496 7926 11570 7986
rect 11630 7926 11671 7986
rect 11423 7894 11671 7926
rect 12747 7909 13129 7920
rect 11423 7874 11740 7894
rect 11423 7872 11837 7874
rect 11423 7812 11431 7872
rect 11491 7860 11837 7872
rect 11491 7812 11560 7860
rect 11423 7800 11560 7812
rect 11620 7802 11837 7860
rect 12692 7851 13129 7909
rect 11620 7800 11740 7802
rect 11423 7782 11740 7800
rect 12747 7798 13129 7851
rect 11423 7781 11671 7782
rect 5268 7610 6063 7709
rect -63 7568 6063 7610
rect -63 7564 5727 7568
rect -63 7548 5588 7564
rect -63 7488 5391 7548
rect 5451 7504 5588 7548
rect 5648 7508 5727 7564
rect 5787 7564 6063 7568
rect 5787 7508 5871 7564
rect 5648 7504 5871 7508
rect 5931 7504 6063 7564
rect 5451 7488 6063 7504
rect -63 7444 6063 7488
rect -63 7430 5850 7444
rect -63 7423 5676 7430
rect -63 7418 5503 7423
rect -63 7358 5354 7418
rect 5414 7363 5503 7418
rect 5563 7370 5676 7423
rect 5736 7384 5850 7430
rect 5910 7384 6063 7444
rect 5736 7370 6063 7384
rect 5563 7363 6063 7370
rect 5414 7358 6063 7363
rect -63 7315 6063 7358
rect 10683 7569 11112 7726
rect 10683 7355 11727 7569
rect 10753 7354 11727 7355
rect -63 7310 5939 7315
rect -63 7306 5637 7310
rect -63 7298 5474 7306
rect -63 7238 5323 7298
rect 5383 7246 5474 7298
rect 5534 7250 5637 7306
rect 5697 7250 5798 7310
rect 5858 7255 5939 7310
rect 5999 7255 6063 7315
rect 13007 7311 13129 7798
rect 5858 7250 6063 7255
rect 5534 7246 6063 7250
rect 5383 7238 6063 7246
rect -63 7228 6063 7238
rect 5268 7226 6063 7228
rect 12940 7309 13192 7311
rect 12940 7249 12962 7309
rect 13022 7249 13098 7309
rect 13158 7249 13192 7309
rect 12940 7196 13192 7249
rect 8560 7077 9108 7137
rect 12940 7136 12957 7196
rect 13017 7189 13192 7196
rect 13017 7136 13093 7189
rect 12940 7129 13093 7136
rect 13153 7129 13192 7189
rect 12940 7111 13192 7129
rect 8560 7072 8949 7077
rect 8560 7012 8594 7072
rect 8654 7012 8737 7072
rect 8797 7017 8949 7072
rect 9009 7017 9108 7077
rect 8797 7012 9108 7017
rect 8560 6960 9108 7012
rect 8560 6900 8594 6960
rect 8654 6900 8742 6960
rect 8802 6900 8980 6960
rect 9040 6900 9108 6960
rect 8560 6879 9108 6900
rect 12397 5486 12483 5488
rect 12397 5407 12791 5486
rect 12397 5396 12675 5407
rect 12397 5336 12498 5396
rect 12558 5347 12675 5396
rect 12735 5347 12791 5407
rect 12558 5336 12791 5347
rect 12397 5275 12791 5336
rect 12397 5265 12568 5275
rect 12397 5205 12432 5265
rect 12492 5215 12568 5265
rect 12628 5270 12791 5275
rect 12628 5215 12715 5270
rect 12492 5210 12715 5215
rect 12775 5210 12791 5270
rect 12492 5205 12791 5210
rect 12397 5185 12791 5205
rect 5586 4579 6428 4675
rect 4778 -986 5148 -932
rect 4778 -1046 4824 -986
rect 4884 -988 5148 -986
rect 4884 -1046 4988 -988
rect 4778 -1048 4988 -1046
rect 5048 -1048 5148 -988
rect 4778 -1072 5148 -1048
rect 4422 -1100 5148 -1072
rect 4422 -1113 4990 -1100
rect 4422 -1173 4824 -1113
rect 4884 -1160 4990 -1113
rect 5050 -1160 5148 -1100
rect 4884 -1173 5148 -1160
rect 4422 -1237 5148 -1173
rect 4778 -1240 5148 -1237
rect 4778 -1251 4995 -1240
rect 4778 -1311 4824 -1251
rect 4884 -1300 4995 -1251
rect 5055 -1300 5148 -1240
rect 4884 -1311 5148 -1300
rect 4778 -1338 5148 -1311
rect 4844 -1524 5214 -1512
rect 4488 -1552 5214 -1524
rect 4488 -1565 5056 -1552
rect 4488 -1625 4890 -1565
rect 4950 -1612 5056 -1565
rect 5116 -1612 5214 -1552
rect 4950 -1625 5214 -1612
rect 4488 -1689 5214 -1625
rect 4844 -1692 5214 -1689
rect 4844 -1703 5061 -1692
rect 4844 -1763 4890 -1703
rect 4950 -1752 5061 -1703
rect 5121 -1752 5214 -1692
rect 4950 -1763 5214 -1752
rect 4844 -1790 5214 -1763
rect 4506 -2249 4874 -2240
rect 4506 -2309 4792 -2249
rect 4852 -2309 4874 -2249
rect 4506 -2330 4874 -2309
rect 4377 -2352 4874 -2330
rect 4377 -2412 4543 -2352
rect 4603 -2412 4683 -2352
rect 4743 -2412 4874 -2352
rect 4377 -2441 4874 -2412
rect 4506 -2473 4874 -2441
rect 4506 -2533 4545 -2473
rect 4605 -2476 4874 -2473
rect 4605 -2533 4691 -2476
rect 4506 -2536 4691 -2533
rect 4751 -2481 4874 -2476
rect 4751 -2536 4811 -2481
rect 4506 -2541 4811 -2536
rect 4871 -2541 4874 -2481
rect 4506 -2563 4874 -2541
rect 5001 -2620 5371 -2608
rect 4645 -2648 5371 -2620
rect 4645 -2661 5213 -2648
rect 4645 -2721 5047 -2661
rect 5107 -2708 5213 -2661
rect 5273 -2708 5371 -2648
rect 5107 -2721 5371 -2708
rect 4645 -2785 5371 -2721
rect 5001 -2788 5371 -2785
rect 5001 -2799 5218 -2788
rect 5001 -2859 5047 -2799
rect 5107 -2848 5218 -2799
rect 5278 -2848 5371 -2788
rect 5107 -2859 5371 -2848
rect 5001 -2886 5371 -2859
rect 4905 -3038 5275 -3026
rect 4549 -3066 5275 -3038
rect 4549 -3079 5117 -3066
rect 4549 -3139 4951 -3079
rect 5011 -3126 5117 -3079
rect 5177 -3126 5275 -3066
rect 5011 -3139 5275 -3126
rect 4549 -3203 5275 -3139
rect 4905 -3206 5275 -3203
rect 4905 -3217 5122 -3206
rect 4905 -3277 4951 -3217
rect 5011 -3266 5122 -3217
rect 5182 -3266 5275 -3206
rect 5011 -3277 5275 -3266
rect 4905 -3304 5275 -3277
rect 4882 -3452 5252 -3440
rect 4526 -3480 5252 -3452
rect 4526 -3493 5094 -3480
rect 4526 -3553 4928 -3493
rect 4988 -3540 5094 -3493
rect 5154 -3540 5252 -3480
rect 4988 -3553 5252 -3540
rect 4526 -3617 5252 -3553
rect 4882 -3620 5252 -3617
rect 4882 -3631 5099 -3620
rect 4882 -3691 4928 -3631
rect 4988 -3680 5099 -3631
rect 5159 -3680 5252 -3620
rect 4988 -3691 5252 -3680
rect 4882 -3718 5252 -3691
rect 4928 -3931 5298 -3919
rect 4572 -3959 5298 -3931
rect 4572 -3972 5140 -3959
rect 4572 -4032 4974 -3972
rect 5034 -4019 5140 -3972
rect 5200 -4019 5298 -3959
rect 5034 -4032 5298 -4019
rect 4572 -4096 5298 -4032
rect 4928 -4099 5298 -4096
rect 4928 -4110 5145 -4099
rect 4928 -4170 4974 -4110
rect 5034 -4159 5145 -4110
rect 5205 -4159 5298 -4099
rect 5034 -4170 5298 -4159
rect 4928 -4197 5298 -4170
rect 5033 -4474 5403 -4462
rect 4677 -4502 5403 -4474
rect 4677 -4515 5245 -4502
rect 4677 -4575 5079 -4515
rect 5139 -4562 5245 -4515
rect 5305 -4562 5403 -4502
rect 5139 -4575 5403 -4562
rect 4677 -4639 5403 -4575
rect 5033 -4642 5403 -4639
rect 5033 -4653 5250 -4642
rect 5033 -4713 5079 -4653
rect 5139 -4702 5250 -4653
rect 5310 -4702 5403 -4642
rect 5139 -4713 5403 -4702
rect 5033 -4740 5403 -4713
rect 5638 -5420 5862 -5418
rect 8579 -5420 9022 3070
rect 9531 -5420 9974 3070
rect 10350 -5420 10793 3070
rect 13382 -3641 14075 13958
rect 17890 13943 18200 14008
rect 17890 13891 17919 13943
rect 17971 13891 18023 13943
rect 18075 13891 18127 13943
rect 18179 13891 18200 13943
rect 17890 13839 18200 13891
rect 17890 13787 17919 13839
rect 17971 13787 18023 13839
rect 18075 13787 18127 13839
rect 18179 13787 18200 13839
rect 17890 13738 18200 13787
rect 19198 14114 19410 14168
rect 20406 14143 20600 14210
rect 28009 14162 45862 14382
rect 20393 14129 20705 14143
rect 19198 14062 19222 14114
rect 19274 14062 19326 14114
rect 19378 14062 19410 14114
rect 19198 14010 19410 14062
rect 19198 13958 19222 14010
rect 19274 13958 19326 14010
rect 19378 13958 19410 14010
rect 19198 13906 19410 13958
rect 19198 13854 19222 13906
rect 19274 13854 19326 13906
rect 19378 13854 19410 13906
rect 19198 13802 19410 13854
rect 20370 14091 20705 14129
rect 20370 14039 20393 14091
rect 20445 14039 20497 14091
rect 20549 14039 20601 14091
rect 20653 14039 20705 14091
rect 22087 14087 23144 14135
rect 20370 13987 20705 14039
rect 20370 13935 20393 13987
rect 20445 13935 20497 13987
rect 20549 13935 20601 13987
rect 20653 13935 20705 13987
rect 20370 13883 20705 13935
rect 21918 13926 22114 14087
rect 22275 14086 22915 14087
rect 22275 13927 22497 14086
rect 22656 13927 22915 14086
rect 22275 13926 22915 13927
rect 23076 13926 23144 14087
rect 22087 13904 23144 13926
rect 28009 14102 37931 14162
rect 37991 14102 38051 14162
rect 38111 14102 38171 14162
rect 38231 14102 38291 14162
rect 38351 14102 38411 14162
rect 38471 14102 45862 14162
rect 28009 14042 45862 14102
rect 28009 13982 37931 14042
rect 37991 13982 38051 14042
rect 38111 13982 38171 14042
rect 38231 13982 38291 14042
rect 38351 13982 38411 14042
rect 38471 13982 45862 14042
rect 28009 13917 45862 13982
rect 20370 13831 20393 13883
rect 20445 13831 20497 13883
rect 20549 13831 20601 13883
rect 20653 13831 20705 13883
rect 20370 13811 20705 13831
rect 19198 13750 19222 13802
rect 19274 13750 19326 13802
rect 19378 13750 19410 13802
rect 19198 13738 19410 13750
rect 21938 13658 22849 13700
rect 21833 13522 21964 13658
rect 22100 13657 22678 13658
rect 22100 13523 22388 13657
rect 22522 13523 22678 13657
rect 22100 13522 22678 13523
rect 22814 13522 22849 13658
rect 21938 13497 22849 13522
rect 21781 13264 22530 13292
rect 21781 13162 21813 13264
rect 21915 13263 22385 13264
rect 21915 13163 22053 13263
rect 22153 13163 22385 13263
rect 21915 13162 22385 13163
rect 22487 13162 22530 13264
rect 21781 13142 22530 13162
rect 28009 13000 28474 13917
rect 29826 13329 30426 13389
rect 29802 13269 29826 13323
rect 29886 13269 29946 13329
rect 30006 13269 30066 13329
rect 30126 13269 30186 13329
rect 30246 13269 30306 13329
rect 30366 13323 30426 13329
rect 30366 13269 31638 13323
rect 29802 13209 31638 13269
rect 29802 13149 29826 13209
rect 29886 13149 29946 13209
rect 30006 13149 30066 13209
rect 30126 13149 30186 13209
rect 30246 13149 30306 13209
rect 30366 13149 31638 13209
rect 29802 13134 31638 13149
rect 28009 12882 28470 13000
rect 22767 12489 24077 12615
rect 25831 12525 28470 12882
rect 22767 12487 23800 12489
rect 22767 12486 23246 12487
rect 22823 12412 22947 12486
rect 23122 12412 23246 12486
rect 23406 12412 23530 12487
rect 23676 12412 23800 12487
rect 23953 12412 24077 12489
rect 25830 12503 28470 12525
rect 25830 12433 26744 12503
rect 24624 12412 24967 12413
rect 25540 12412 25770 12413
rect 25830 12412 26545 12433
rect 16702 12108 17532 12110
rect 16702 11903 18051 12108
rect 22793 11960 26545 12412
rect 16702 11653 17532 11903
rect 16702 11448 18065 11653
rect 26224 11549 26277 11586
rect 16702 11170 17532 11448
rect 22449 11211 22560 11220
rect 19654 11192 19738 11204
rect 16702 10965 18065 11170
rect 19654 11132 19666 11192
rect 19726 11132 19738 11192
rect 19654 11121 19738 11132
rect 19895 11197 19979 11209
rect 19895 11137 19907 11197
rect 19967 11137 19979 11197
rect 20134 11199 20218 11211
rect 20134 11139 20146 11199
rect 19895 11126 19979 11137
rect 20206 11128 20218 11199
rect 20361 11199 20445 11211
rect 20361 11139 20373 11199
rect 20433 11139 20445 11199
rect 20361 11128 20445 11139
rect 22449 11171 22956 11211
rect 22449 11111 22477 11171
rect 22537 11111 22956 11171
rect 22449 11110 22956 11111
rect 22449 11027 22560 11110
rect 22449 10967 22472 11027
rect 22532 10967 22560 11027
rect 16702 10715 17532 10965
rect 22449 10942 22560 10967
rect 16702 10510 18070 10715
rect 16702 9691 17532 10510
rect 20845 10390 21011 10561
rect 21224 10390 21390 10578
rect 21511 10390 21677 10561
rect 20845 10386 21677 10390
rect 21966 10388 22132 10574
rect 21966 10386 23117 10388
rect 20845 10224 23117 10386
rect 21511 10222 23117 10224
rect 31449 10181 31638 13134
rect 31886 11708 32351 13917
rect 44097 13154 44562 13917
rect 44130 13150 44562 13154
rect 45397 13145 45862 13917
rect 64769 13781 65603 13916
rect 64769 13718 64920 13781
rect 47691 13711 64920 13718
rect 64990 13777 65603 13781
rect 64990 13711 65179 13777
rect 47691 13707 65179 13711
rect 65249 13712 65603 13777
rect 65249 13707 65420 13712
rect 47691 13642 65420 13707
rect 65490 13642 65603 13712
rect 47691 13630 65603 13642
rect 47691 13560 64924 13630
rect 64994 13600 65603 13630
rect 64994 13560 65191 13600
rect 47691 13530 65191 13560
rect 65261 13559 65603 13600
rect 65261 13530 65415 13559
rect 47691 13489 65415 13530
rect 65485 13489 65603 13559
rect 47691 13463 65603 13489
rect 47691 13461 65181 13463
rect 47691 13391 64923 13461
rect 64993 13393 65181 13461
rect 65251 13416 65603 13463
rect 65251 13393 65413 13416
rect 64993 13391 65413 13393
rect 47691 13346 65413 13391
rect 65483 13346 65603 13416
rect 47691 13286 65603 13346
rect 47691 13216 64973 13286
rect 65043 13281 65603 13286
rect 65043 13216 65175 13281
rect 47691 13211 65175 13216
rect 65245 13269 65603 13281
rect 65245 13211 65338 13269
rect 47691 13199 65338 13211
rect 65408 13199 65603 13269
rect 47691 13149 65603 13199
rect 41677 12670 41885 12734
rect 41677 12547 41720 12670
rect 41843 12547 41885 12670
rect 41677 12421 41885 12547
rect 41677 12296 41719 12421
rect 41844 12296 41885 12421
rect 41677 12214 41885 12296
rect 41677 12196 42058 12214
rect 41677 12073 41720 12196
rect 41843 12073 42058 12196
rect 41677 12061 42058 12073
rect 37793 10788 38571 10840
rect 37793 10728 37873 10788
rect 37933 10728 37993 10788
rect 38053 10728 38113 10788
rect 38173 10728 38233 10788
rect 38293 10728 38353 10788
rect 38413 10728 38571 10788
rect 37793 10668 38571 10728
rect 37793 10608 37873 10668
rect 37933 10608 37993 10668
rect 38053 10608 38113 10668
rect 38173 10608 38233 10668
rect 38293 10608 38353 10668
rect 38413 10608 38571 10668
rect 37793 10547 38571 10608
rect 19888 9897 22600 10122
rect 31449 10073 32313 10181
rect 31449 9975 31638 10073
rect 28770 9909 28848 9964
rect 29009 9914 29087 9964
rect 29248 9916 29326 9964
rect 29474 9916 29552 9964
rect 16702 9264 17980 9691
rect 22373 9505 22600 9897
rect 28768 9897 28852 9909
rect 28768 9837 28780 9897
rect 28840 9837 28852 9897
rect 28768 9826 28852 9837
rect 29009 9902 29093 9914
rect 29009 9842 29021 9902
rect 29081 9842 29093 9902
rect 29009 9831 29093 9842
rect 29248 9904 29332 9916
rect 29248 9844 29260 9904
rect 29320 9844 29332 9904
rect 29248 9833 29332 9844
rect 29474 9904 29559 9916
rect 29474 9844 29487 9904
rect 29547 9844 29559 9904
rect 29474 9833 29559 9844
rect 28770 9794 28848 9826
rect 29009 9794 29087 9831
rect 29248 9794 29326 9833
rect 29474 9794 29552 9833
rect 22373 9472 22743 9505
rect 22373 9390 22985 9472
rect 22373 9358 22743 9390
rect 16702 8606 17532 9264
rect 19614 9158 19692 9209
rect 19853 9163 19931 9209
rect 20318 9165 20396 9209
rect 19612 9146 19696 9158
rect 19612 9086 19624 9146
rect 19684 9086 19696 9146
rect 19612 9075 19696 9086
rect 19853 9151 19937 9163
rect 20318 9153 20403 9165
rect 19853 9091 19865 9151
rect 19925 9091 19937 9151
rect 19853 9080 19937 9091
rect 20092 9093 20104 9153
rect 20164 9093 20176 9153
rect 20092 9082 20176 9093
rect 20318 9093 20331 9153
rect 20391 9093 20403 9153
rect 20318 9082 20403 9093
rect 19614 9039 19692 9075
rect 19853 9039 19931 9080
rect 20092 9039 20170 9082
rect 20318 9039 20396 9082
rect 26167 8889 26249 8932
rect 16702 8179 18037 8606
rect 27648 8585 27807 9468
rect 27901 8593 28060 9476
rect 28305 8593 28464 9476
rect 28660 8589 28819 9472
rect 30473 8717 30883 9048
rect 26351 8450 26523 8578
rect 16702 4973 17532 8179
rect 22865 7922 22989 8384
rect 23323 7922 23447 8384
rect 24418 7922 24542 8396
rect 25281 7922 25405 8393
rect 25975 7922 26099 8413
rect 26224 8326 26523 8450
rect 26343 8324 26523 8326
rect 26351 7922 26523 8324
rect 22840 7885 26523 7922
rect 22840 7883 23415 7885
rect 22840 7878 23176 7883
rect 22840 7818 22935 7878
rect 22995 7823 23176 7878
rect 23236 7825 23415 7883
rect 23475 7825 23642 7885
rect 23702 7825 26523 7885
rect 23236 7823 26523 7825
rect 22995 7818 26523 7823
rect 22840 7798 26523 7818
rect 26351 7706 26523 7798
rect 18490 7270 18630 7520
rect 28714 6915 28792 6970
rect 28953 6920 29031 6970
rect 29192 6922 29270 6970
rect 29418 6922 29496 6970
rect 28712 6903 28796 6915
rect 22095 6822 22546 6850
rect 28712 6843 28724 6903
rect 28784 6843 28796 6903
rect 28712 6832 28796 6843
rect 28953 6908 29037 6920
rect 28953 6848 28965 6908
rect 29025 6848 29037 6908
rect 28953 6837 29037 6848
rect 29192 6910 29276 6922
rect 29192 6850 29204 6910
rect 29264 6850 29276 6910
rect 29192 6839 29276 6850
rect 29418 6910 29503 6922
rect 29418 6850 29431 6910
rect 29491 6850 29503 6910
rect 29418 6839 29503 6850
rect 17937 6751 18038 6809
rect 22095 6791 22102 6822
rect 17937 6711 19507 6751
rect 17937 6674 19508 6711
rect 21988 6705 22102 6791
rect 22219 6821 22546 6822
rect 22219 6706 22399 6821
rect 22514 6706 22546 6821
rect 28714 6800 28792 6832
rect 28953 6800 29031 6837
rect 29192 6800 29270 6839
rect 29418 6800 29496 6839
rect 22219 6705 22546 6706
rect 22085 6683 22546 6705
rect 17937 6646 18068 6674
rect 17938 6614 18068 6646
rect 18128 6614 18188 6674
rect 18248 6614 18308 6674
rect 18368 6614 18428 6674
rect 18488 6614 18548 6674
rect 18608 6614 18668 6674
rect 18728 6614 18788 6674
rect 18848 6614 18908 6674
rect 18968 6614 19028 6674
rect 19088 6614 19148 6674
rect 19208 6614 19268 6674
rect 19328 6614 19388 6674
rect 19448 6614 19508 6674
rect 17938 6585 19508 6614
rect 26889 5053 27137 6444
rect 27452 5078 27700 6469
rect 27937 5086 28185 6477
rect 28962 6257 29078 6331
rect 31485 6257 31602 9975
rect 32011 9884 32303 9911
rect 32011 9822 32070 9884
rect 32132 9822 32303 9884
rect 32011 9792 32303 9822
rect 28962 6141 31602 6257
rect 33295 9275 33729 9309
rect 36032 9299 36466 10247
rect 36737 9299 37171 10223
rect 36032 9275 37171 9299
rect 33295 8865 37171 9275
rect 33295 8841 36466 8865
rect 32225 5373 32329 5795
rect 33295 5113 33729 8841
rect 47691 8256 48260 13149
rect 64769 13020 65603 13149
rect 55240 9830 56170 9840
rect 47615 8242 48260 8256
rect 47615 8241 47935 8242
rect 47615 8163 47780 8241
rect 47858 8163 47935 8241
rect 47615 8162 47935 8163
rect 48015 8162 48260 8242
rect 47615 8150 48260 8162
rect 47690 7940 48260 8150
rect 50084 9609 57840 9830
rect 50084 7719 50305 9609
rect 53921 9320 54794 9377
rect 53921 9256 54010 9320
rect 54070 9316 54130 9320
rect 54190 9319 54250 9320
rect 54070 9256 54129 9316
rect 54190 9260 54246 9319
rect 54310 9260 54370 9320
rect 54430 9319 54490 9320
rect 54430 9260 54487 9319
rect 54550 9260 54794 9320
rect 54189 9259 54246 9260
rect 54306 9259 54487 9260
rect 54547 9259 54794 9260
rect 54189 9256 54794 9259
rect 53921 9206 54794 9256
rect 53921 9202 54371 9206
rect 53921 9200 54251 9202
rect 54311 9200 54371 9202
rect 54431 9200 54794 9206
rect 53921 9140 54010 9200
rect 54070 9140 54128 9200
rect 54190 9140 54250 9200
rect 54311 9142 54370 9200
rect 54431 9199 54490 9200
rect 54431 9146 54489 9199
rect 54310 9140 54370 9142
rect 54430 9140 54489 9146
rect 54550 9140 54794 9200
rect 53921 9139 54489 9140
rect 54549 9139 54794 9140
rect 53921 9088 54794 9139
rect 50084 7338 50292 7719
rect 43227 7112 43321 7123
rect 46153 7119 46241 7191
rect 46418 7119 46522 7199
rect 46706 7119 46809 7195
rect 46908 7119 47009 7188
rect 48084 7130 50292 7338
rect 57619 7531 57840 9609
rect 61491 9327 62361 9385
rect 61491 9263 61580 9327
rect 61640 9323 61700 9327
rect 61760 9326 61820 9327
rect 61640 9263 61699 9323
rect 61760 9267 61816 9326
rect 61880 9267 61940 9327
rect 62000 9326 62060 9327
rect 62000 9267 62057 9326
rect 62120 9267 62361 9327
rect 61759 9266 61816 9267
rect 61876 9266 62057 9267
rect 62117 9266 62361 9267
rect 61759 9263 62361 9266
rect 61491 9213 62361 9263
rect 61491 9209 61941 9213
rect 61491 9207 61821 9209
rect 61881 9207 61941 9209
rect 62001 9207 62361 9213
rect 61491 9147 61580 9207
rect 61640 9147 61698 9207
rect 61760 9147 61820 9207
rect 61881 9149 61940 9207
rect 62001 9206 62060 9207
rect 62001 9153 62059 9206
rect 61880 9147 61940 9149
rect 62000 9147 62059 9153
rect 62120 9147 62361 9207
rect 61491 9146 62059 9147
rect 62119 9146 62361 9147
rect 61491 9099 62361 9146
rect 58049 7531 58270 8320
rect 66783 7933 67158 15296
rect 57619 7310 58270 7531
rect 43227 7111 43449 7112
rect 43820 7111 43992 7112
rect 43227 6941 43278 7111
rect 43448 6941 43821 7111
rect 43991 7110 44714 7111
rect 43991 6942 44532 7110
rect 44700 6942 44714 7110
rect 46136 7091 47059 7119
rect 46136 7086 46925 7091
rect 46136 7008 46183 7086
rect 46259 7083 46925 7086
rect 46259 7081 46709 7083
rect 46259 7008 46429 7081
rect 46136 7003 46429 7008
rect 46505 7005 46709 7081
rect 46785 7013 46925 7083
rect 47001 7013 47059 7091
rect 46785 7005 47059 7013
rect 46505 7003 47059 7005
rect 46136 6961 47059 7003
rect 43991 6941 44714 6942
rect 43227 6940 43449 6941
rect 43820 6940 43992 6941
rect 43227 6919 43321 6940
rect 38263 6633 39669 6671
rect 38263 6430 39317 6633
rect 38287 6427 39317 6430
rect 39523 6427 39913 6633
rect 38287 6418 39669 6427
rect 38287 6414 38493 6418
rect 43759 6087 44718 6127
rect 43759 6009 43813 6087
rect 43889 6074 44718 6087
rect 43889 6009 44062 6074
rect 43759 5996 44062 6009
rect 44138 6073 44718 6074
rect 44138 6069 44518 6073
rect 44138 5996 44296 6069
rect 43759 5991 44296 5996
rect 44372 5995 44518 6069
rect 44594 5995 44718 6073
rect 44372 5991 44718 5995
rect 43759 5971 44718 5991
rect 16702 4546 24378 4973
rect 40140 4953 42232 5122
rect 16702 3267 17532 4546
rect 21250 3267 21677 4546
rect 30400 4524 30604 4659
rect 27094 4444 27485 4463
rect 27094 4443 27342 4444
rect 27094 4315 27111 4443
rect 27239 4315 27342 4443
rect 27094 4314 27342 4315
rect 27472 4314 27485 4444
rect 27094 4248 27485 4314
rect 30400 4399 30434 4524
rect 30559 4399 30604 4524
rect 30400 4263 30604 4399
rect 27094 4118 27107 4248
rect 27237 4247 27485 4248
rect 27237 4119 27343 4247
rect 27471 4119 27485 4247
rect 30300 4262 30604 4263
rect 30300 4139 30435 4262
rect 30558 4139 30604 4262
rect 42800 4230 42910 4490
rect 43290 4210 43400 4470
rect 30300 4138 30604 4139
rect 30400 4129 30604 4138
rect 27237 4118 27485 4119
rect 27094 4108 27485 4118
rect 27110 3940 27240 4108
rect 16702 2840 24359 3267
rect 16702 1379 17532 2840
rect 21227 1379 21654 2840
rect 44729 2789 45104 4670
rect 48084 2343 48292 7130
rect 50084 6664 50292 7130
rect 56251 6721 56621 6792
rect 58049 6680 58270 7310
rect 66784 6887 67156 7933
rect 64336 6799 67156 6887
rect 64234 6728 67156 6799
rect 64336 6639 67156 6728
rect 66784 6577 67156 6639
rect 49311 5107 64328 5157
rect 48076 2220 48292 2343
rect 48596 4954 64328 5107
rect 48596 4904 49514 4954
rect 48596 1659 48799 4904
rect 49311 4006 49514 4904
rect 49799 4761 50002 4954
rect 51438 4912 51796 4954
rect 51593 4761 51796 4912
rect 49799 4558 51796 4761
rect 53695 4666 54568 4724
rect 53695 4602 53784 4666
rect 53844 4662 53904 4666
rect 53964 4665 54024 4666
rect 53844 4602 53903 4662
rect 53964 4606 54020 4665
rect 54084 4606 54144 4666
rect 54204 4665 54264 4666
rect 54204 4606 54261 4665
rect 54324 4606 54568 4666
rect 53963 4605 54020 4606
rect 54080 4605 54261 4606
rect 54321 4605 54568 4606
rect 53963 4602 54568 4605
rect 49799 4006 50002 4558
rect 53695 4552 54568 4602
rect 53695 4548 54145 4552
rect 53695 4546 54025 4548
rect 54085 4546 54145 4548
rect 54205 4546 54568 4552
rect 53695 4486 53784 4546
rect 53844 4486 53902 4546
rect 53964 4486 54024 4546
rect 54085 4488 54144 4546
rect 54205 4545 54264 4546
rect 54205 4492 54263 4545
rect 54084 4486 54144 4488
rect 54204 4486 54263 4492
rect 54324 4486 54568 4546
rect 53695 4485 54263 4486
rect 54323 4485 54568 4486
rect 53695 4412 54568 4485
rect 53695 4319 54344 4412
rect 53701 4315 54344 4319
rect 53701 4314 54194 4315
rect 49311 3803 50002 4006
rect 49311 1659 49514 3803
rect 50335 2374 50478 3627
rect 47450 1456 49514 1659
rect 50081 2231 50478 2374
rect 16702 952 24382 1379
rect 47945 1007 48083 1256
rect 50081 1007 50224 2231
rect 50335 1992 50478 2231
rect 56403 2041 56855 2118
rect 16702 -1185 17532 952
rect 19771 -1203 20198 952
rect 47943 864 50224 1007
rect 50715 -448 51181 505
rect 52024 -448 52490 458
rect 53443 -448 53909 458
rect 54484 -448 54950 458
rect 74047 -448 74513 -207
rect 47429 -914 74513 -448
rect 88322 -822 88697 15482
rect 98848 4721 99160 4739
rect 98848 4666 98886 4721
rect 98945 4715 99160 4721
rect 98945 4666 99061 4715
rect 98848 4660 99061 4666
rect 99120 4660 99160 4715
rect 98848 4566 99482 4660
rect 98848 4562 99062 4566
rect 98848 4507 98884 4562
rect 98943 4511 99062 4562
rect 99121 4511 99482 4566
rect 98943 4507 99482 4511
rect 98848 4440 99482 4507
rect 98848 4397 99160 4440
rect 98848 4342 98887 4397
rect 98946 4392 99160 4397
rect 98946 4342 99075 4392
rect 98848 4337 99075 4342
rect 99134 4337 99160 4392
rect 91327 4259 92059 4316
rect 98848 4305 99160 4337
rect 91327 4195 91416 4259
rect 91476 4255 91536 4259
rect 91596 4258 91656 4259
rect 91476 4195 91535 4255
rect 91596 4199 91652 4258
rect 91716 4199 91776 4259
rect 91836 4258 91896 4259
rect 91836 4199 91893 4258
rect 91956 4199 92059 4259
rect 91595 4198 91652 4199
rect 91712 4198 91893 4199
rect 91953 4198 92059 4199
rect 91595 4195 92059 4198
rect 91327 4145 92059 4195
rect 91327 4141 91777 4145
rect 91327 4139 91657 4141
rect 91717 4139 91777 4141
rect 91837 4139 92059 4145
rect 91327 4079 91416 4139
rect 91476 4079 91534 4139
rect 91596 4079 91656 4139
rect 91717 4081 91776 4139
rect 91837 4138 91896 4139
rect 91837 4085 91895 4138
rect 91716 4079 91776 4081
rect 91836 4079 91895 4085
rect 91956 4079 92059 4139
rect 91327 4078 91895 4079
rect 91955 4078 92059 4079
rect 91327 4051 92059 4078
rect 95080 2670 95620 2970
rect 95080 2610 95232 2670
rect 95292 2610 95352 2670
rect 95412 2610 95472 2670
rect 95532 2610 95620 2670
rect 95080 2550 95620 2610
rect 95080 2490 95232 2550
rect 95292 2490 95352 2550
rect 95412 2490 95472 2550
rect 95532 2490 95620 2550
rect 95080 2430 95620 2490
rect 95080 2370 95232 2430
rect 95292 2370 95352 2430
rect 95412 2370 95472 2430
rect 95532 2370 95620 2430
rect 95080 2270 95620 2370
rect 90062 -69 90216 161
rect 90062 -223 91541 -69
rect 90062 -240 90357 -223
rect 89933 -298 90357 -240
rect 89933 -310 90127 -298
rect 89933 -370 90003 -310
rect 90063 -358 90127 -310
rect 90187 -358 90357 -298
rect 90063 -370 90357 -358
rect 89933 -410 90357 -370
rect 91387 -410 91541 -223
rect 93502 -410 93656 120
rect 89933 -427 93656 -410
rect 89933 -487 90021 -427
rect 90081 -439 93656 -427
rect 90081 -487 90145 -439
rect 89933 -499 90145 -487
rect 90205 -499 93656 -439
rect 89933 -564 93656 -499
rect 89933 -570 90316 -564
rect 50307 -915 50773 -914
rect 52557 -915 53023 -914
rect 55367 -915 55833 -914
rect 18080 -1503 18860 -1470
rect 18080 -1510 18665 -1503
rect 18080 -1515 18415 -1510
rect 18080 -1628 18108 -1515
rect 18235 -1623 18415 -1515
rect 18542 -1616 18665 -1510
rect 18792 -1616 18860 -1503
rect 18542 -1623 18860 -1616
rect 18235 -1628 18860 -1623
rect 18080 -1660 18860 -1628
rect 58411 -2964 58526 -2610
rect 58344 -3011 58612 -2964
rect 58344 -3036 58526 -3011
rect 58344 -3095 58356 -3036
rect 58411 -3070 58526 -3036
rect 58581 -3070 58612 -3011
rect 58411 -3095 58612 -3070
rect 58344 -3209 58612 -3095
rect 58344 -3210 58521 -3209
rect 58344 -3269 58355 -3210
rect 58410 -3268 58521 -3210
rect 58576 -3268 58612 -3209
rect 58410 -3269 58612 -3268
rect 58344 -3325 58612 -3269
rect 20040 -3641 20542 -3449
rect 13382 -3920 20542 -3641
rect 13382 -4128 14075 -3920
rect 60197 -5340 60663 -914
rect 64717 -5340 65183 -914
rect 66293 -5340 66759 -914
rect 68159 -3639 68520 -3628
rect 68159 -3694 68215 -3639
rect 68274 -3640 68520 -3639
rect 68274 -3694 68389 -3640
rect 68159 -3695 68389 -3694
rect 68448 -3695 68520 -3640
rect 68159 -3805 69109 -3695
rect 68159 -3860 68216 -3805
rect 68275 -3810 69109 -3805
rect 68275 -3860 68414 -3810
rect 68159 -3865 68414 -3860
rect 68473 -3865 68520 -3810
rect 68159 -3896 68520 -3865
rect 70747 -5340 71213 -914
rect 73441 -5340 73907 -914
rect 87273 -1197 88697 -822
rect 98561 -760 98873 -742
rect 98561 -815 98599 -760
rect 98658 -766 98873 -760
rect 98658 -815 98774 -766
rect 98561 -821 98774 -815
rect 98833 -821 98873 -766
rect 98561 -900 98873 -821
rect 98561 -915 99246 -900
rect 98561 -919 98775 -915
rect 98561 -974 98597 -919
rect 98656 -970 98775 -919
rect 98834 -970 99246 -915
rect 98656 -974 99246 -970
rect 98561 -1057 99246 -974
rect 98561 -1084 98873 -1057
rect 98561 -1139 98600 -1084
rect 98659 -1089 98873 -1084
rect 98659 -1139 98788 -1089
rect 98561 -1144 98788 -1139
rect 98847 -1144 98873 -1089
rect 98561 -1181 98873 -1144
rect 87273 -4550 87648 -1197
rect 98576 -1964 98937 -1953
rect 98576 -2019 98632 -1964
rect 98691 -1965 98937 -1964
rect 98691 -2019 98806 -1965
rect 98576 -2020 98806 -2019
rect 98865 -2020 98937 -1965
rect 98576 -2130 99239 -2020
rect 98576 -2185 98633 -2130
rect 98692 -2135 99239 -2130
rect 98692 -2185 98831 -2135
rect 98576 -2190 98831 -2185
rect 98890 -2190 98937 -2135
rect 98576 -2221 98937 -2190
rect 98546 -2861 98907 -2850
rect 98546 -2916 98602 -2861
rect 98661 -2862 98907 -2861
rect 98661 -2916 98776 -2862
rect 98546 -2917 98776 -2916
rect 98835 -2917 98907 -2862
rect 98546 -3027 99209 -2917
rect 98546 -3082 98603 -3027
rect 98662 -3032 99209 -3027
rect 98662 -3082 98801 -3032
rect 98546 -3087 98801 -3082
rect 98860 -3087 98907 -3032
rect 98546 -3118 98907 -3087
rect 98538 -3344 98899 -3333
rect 98538 -3399 98594 -3344
rect 98653 -3345 98899 -3344
rect 98653 -3399 98768 -3345
rect 98538 -3400 98768 -3399
rect 98827 -3400 98899 -3345
rect 98538 -3510 99201 -3400
rect 98538 -3565 98595 -3510
rect 98654 -3515 99201 -3510
rect 98654 -3565 98793 -3515
rect 98538 -3570 98793 -3565
rect 98852 -3570 98899 -3515
rect 98538 -3601 98899 -3570
rect 98576 -3896 98937 -3885
rect 98576 -3951 98632 -3896
rect 98691 -3897 98937 -3896
rect 98691 -3951 98806 -3897
rect 98576 -3952 98806 -3951
rect 98865 -3952 98937 -3897
rect 98576 -4062 99239 -3952
rect 98576 -4117 98633 -4062
rect 98692 -4067 99239 -4062
rect 98692 -4117 98831 -4067
rect 98576 -4122 98831 -4117
rect 98890 -4122 98937 -4067
rect 98576 -4153 98937 -4122
rect 87090 -4720 87760 -4550
rect 87090 -4780 87132 -4720
rect 87192 -4780 87252 -4720
rect 87312 -4780 87372 -4720
rect 87432 -4780 87760 -4720
rect 87090 -4840 87760 -4780
rect 87090 -4900 87132 -4840
rect 87192 -4900 87252 -4840
rect 87312 -4900 87372 -4840
rect 87432 -4900 87760 -4840
rect 87090 -4960 87760 -4900
rect 87090 -5020 87132 -4960
rect 87192 -5020 87252 -4960
rect 87312 -5020 87372 -4960
rect 87432 -5020 87760 -4960
rect 87090 -5090 87760 -5020
rect 5638 -5640 46550 -5420
rect 5638 -26120 5862 -5640
rect 46330 -7116 46550 -5640
rect 56830 -5580 97660 -5340
rect 56830 -7113 57070 -5580
rect 46330 -7305 49145 -7116
rect 6386 -8123 6433 -7467
rect 13089 -7874 13136 -7507
rect 28743 -7995 28833 -7665
rect 13833 -10333 13879 -9997
rect 13098 -12624 13146 -12186
rect 28843 -12493 28889 -11707
rect 25725 -14613 27275 -14562
rect 14185 -16057 14240 -15620
rect 27991 -15636 28043 -14884
rect 28905 -18073 28951 -17807
rect 42594 -18574 45406 -18222
rect 46330 -26120 46550 -7305
rect 54749 -7361 57070 -7113
rect 54726 -8904 56321 -8804
rect 48724 -9293 48793 -9131
rect 48405 -9337 48793 -9293
rect 48405 -9397 48442 -9337
rect 48502 -9349 48793 -9337
rect 48502 -9397 48581 -9349
rect 48405 -9409 48581 -9397
rect 48641 -9409 48793 -9349
rect 48405 -9453 48793 -9409
rect 48405 -9513 48436 -9453
rect 48496 -9474 48793 -9453
rect 48496 -9513 48584 -9474
rect 48405 -9534 48584 -9513
rect 48644 -9534 48793 -9474
rect 48405 -9567 48793 -9534
rect 48405 -9627 48439 -9567
rect 48499 -9590 48793 -9567
rect 48499 -9627 48584 -9590
rect 48405 -9650 48584 -9627
rect 48644 -9650 48793 -9590
rect 48405 -9663 48793 -9650
rect 48724 -10104 48793 -9663
rect 52279 -11322 53565 -11166
rect 52279 -11364 53571 -11322
rect 52279 -11367 53315 -11364
rect 52279 -11375 53073 -11367
rect 52279 -11377 52804 -11375
rect 52279 -11390 52549 -11377
rect 52279 -11450 52344 -11390
rect 52404 -11437 52549 -11390
rect 52609 -11435 52804 -11377
rect 52864 -11427 53073 -11375
rect 53133 -11424 53315 -11367
rect 53375 -11424 53571 -11364
rect 53133 -11427 53571 -11424
rect 52864 -11435 53571 -11427
rect 52609 -11437 53571 -11435
rect 52404 -11450 53571 -11437
rect 52279 -11546 53571 -11450
rect 52279 -11547 53402 -11546
rect 52279 -11559 53243 -11547
rect 52279 -11562 53030 -11559
rect 52279 -11572 52785 -11562
rect 52279 -11580 52552 -11572
rect 52279 -11640 52346 -11580
rect 52406 -11632 52552 -11580
rect 52612 -11622 52785 -11572
rect 52845 -11619 53030 -11562
rect 53090 -11607 53243 -11559
rect 53303 -11606 53402 -11547
rect 53462 -11606 53571 -11546
rect 53303 -11607 53571 -11606
rect 53090 -11619 53571 -11607
rect 52845 -11622 53571 -11619
rect 52612 -11632 53571 -11622
rect 52406 -11640 53571 -11632
rect 52279 -11732 53571 -11640
rect 52279 -11740 53351 -11732
rect 52279 -11750 53153 -11740
rect 52279 -11753 52914 -11750
rect 52279 -11755 52703 -11753
rect 52279 -11756 52505 -11755
rect 52279 -11816 52337 -11756
rect 52397 -11815 52505 -11756
rect 52565 -11813 52703 -11755
rect 52763 -11810 52914 -11753
rect 52974 -11800 53153 -11750
rect 53213 -11792 53351 -11740
rect 53411 -11792 53571 -11732
rect 53213 -11800 53571 -11792
rect 52974 -11810 53571 -11800
rect 52763 -11813 53571 -11810
rect 52565 -11815 53571 -11813
rect 52397 -11816 53571 -11815
rect 52279 -11848 53571 -11816
rect 48991 -14110 49554 -14074
rect 56118 -14110 56321 -8904
rect 48991 -14140 56322 -14110
rect 48789 -14152 56322 -14140
rect 48789 -14212 49195 -14152
rect 49255 -14212 49315 -14152
rect 49375 -14212 49435 -14152
rect 49495 -14212 56322 -14152
rect 48789 -14272 56322 -14212
rect 48789 -14332 49195 -14272
rect 49255 -14332 49315 -14272
rect 49375 -14332 49435 -14272
rect 49495 -14315 56322 -14272
rect 49495 -14332 49554 -14315
rect 48789 -14335 49554 -14332
rect 48991 -14450 49554 -14335
rect 5638 -26332 46550 -26120
rect 5780 -26340 46550 -26332
rect 56830 -26120 57070 -7361
rect 57536 -8443 57583 -7347
rect 64239 -8183 64286 -7477
rect 79893 -8205 79983 -7375
rect 64983 -10117 65030 -10037
rect 64983 -10164 65333 -10117
rect 64983 -10343 65030 -10164
rect 64248 -12534 64296 -11606
rect 79993 -12443 80039 -11737
rect 77165 -14593 77995 -14542
rect 65335 -15997 65390 -15493
rect 65336 -16516 65388 -15997
rect 79141 -16316 79193 -14894
rect 79617 -17833 80103 -17787
rect 80055 -18003 80101 -17833
rect 93784 -18554 96726 -18202
rect 97420 -26120 97660 -5580
rect 98574 -7470 98910 -7460
rect 98574 -7530 98602 -7470
rect 98662 -7530 98722 -7470
rect 98782 -7530 98842 -7470
rect 98902 -7530 98910 -7470
rect 98574 -7590 99250 -7530
rect 98574 -7650 98602 -7590
rect 98662 -7650 98722 -7590
rect 98782 -7650 98842 -7590
rect 98902 -7650 99250 -7590
rect 98574 -7690 99250 -7650
rect 98574 -7710 98910 -7690
rect 98574 -7770 98602 -7710
rect 98662 -7770 98722 -7710
rect 98782 -7770 98842 -7710
rect 98902 -7770 98910 -7710
rect 98574 -7800 98910 -7770
rect 56830 -26360 97660 -26120
<< via1 >>
rect -3054 62742 -2994 62802
rect -2890 62740 -2830 62800
rect -3054 62615 -2994 62675
rect -2888 62628 -2828 62688
rect -3054 62477 -2994 62537
rect -2883 62488 -2823 62548
rect -4013 61301 -3953 61361
rect -3847 61314 -3787 61374
rect -4013 61163 -3953 61223
rect -3842 61174 -3782 61234
rect -2673 52670 -2613 52730
rect -2509 52668 -2449 52728
rect -2673 52543 -2613 52603
rect -2507 52556 -2447 52616
rect -2673 52405 -2613 52465
rect -2502 52416 -2442 52476
rect -3861 52145 -3801 52205
rect -3695 52158 -3635 52218
rect -3861 52007 -3801 52067
rect -3690 52018 -3630 52078
rect -2363 44144 -2303 44204
rect -2199 44142 -2139 44202
rect -2363 44017 -2303 44077
rect -2197 44030 -2137 44090
rect -2363 43879 -2303 43939
rect -2192 43890 -2132 43950
rect -2356 43603 -2296 43663
rect -2192 43601 -2132 43661
rect -2356 43476 -2296 43536
rect -2190 43489 -2130 43549
rect -2356 43338 -2296 43398
rect -2185 43349 -2125 43409
rect -2464 36710 -2404 36770
rect -2300 36708 -2240 36768
rect -2464 36583 -2404 36643
rect -2298 36596 -2238 36656
rect -2464 36445 -2404 36505
rect -2293 36456 -2233 36516
rect -3575 24984 -3515 25044
rect -3455 24984 -3395 25044
rect -3335 24984 -3275 25044
rect -3575 24864 -3515 24924
rect -3455 24864 -3395 24924
rect -3335 24864 -3275 24924
rect -3575 24744 -3515 24804
rect -3455 24744 -3395 24804
rect -3335 24744 -3275 24804
rect 2039 27961 2099 28021
rect 2218 27958 2278 28018
rect 2415 27961 2475 28021
rect 2605 27969 2665 28029
rect 2042 27834 2102 27894
rect 2218 27823 2278 27883
rect 2407 27826 2467 27886
rect 2605 27834 2665 27894
rect 9832 17540 9892 17600
rect 9960 17540 10020 17600
rect 10111 17537 10171 17597
rect 9830 17381 9890 17441
rect 10001 17379 10061 17439
rect 10177 17381 10237 17441
rect 9842 17197 9902 17257
rect 10044 17202 10104 17262
rect 10193 17218 10253 17278
rect 9791 16867 9851 16927
rect 9919 16870 9979 16930
rect 10050 16877 10110 16937
rect 9786 16670 9846 16730
rect 9955 16688 10015 16748
rect 10103 16693 10163 16753
rect 9763 16519 9823 16579
rect 9960 16550 10020 16610
rect 10137 16560 10197 16620
rect 22811 16770 22871 16830
rect 22931 16770 22991 16830
rect 23051 16770 23111 16830
rect 23171 16770 23231 16830
rect 23291 16770 23351 16830
rect 22811 16650 22871 16710
rect 22931 16650 22991 16710
rect 23051 16650 23111 16710
rect 23171 16650 23231 16710
rect 23291 16650 23351 16710
rect 22818 16375 22878 16435
rect 22938 16375 22998 16435
rect 23058 16375 23118 16435
rect 23178 16375 23238 16435
rect 23298 16375 23358 16435
rect 22818 16255 22878 16315
rect 22938 16255 22998 16315
rect 23058 16255 23118 16315
rect 23178 16255 23238 16315
rect 23298 16255 23358 16315
rect 22090 15194 22150 15254
rect 22210 15194 22270 15254
rect 22330 15194 22390 15254
rect 22450 15194 22510 15254
rect 22570 15194 22630 15254
rect 22090 15074 22150 15134
rect 22210 15074 22270 15134
rect 22330 15074 22390 15134
rect 22450 15074 22510 15134
rect 22570 15074 22630 15134
rect 22059 14576 22119 14636
rect 22179 14576 22239 14636
rect 22299 14576 22359 14636
rect 22419 14576 22479 14636
rect 22539 14576 22599 14636
rect 22059 14456 22119 14516
rect 22179 14456 22239 14516
rect 22299 14456 22359 14516
rect 22419 14456 22479 14516
rect 22539 14456 22599 14516
rect 17931 14216 17983 14268
rect 18035 14216 18087 14268
rect 18139 14216 18191 14268
rect 17931 14112 17983 14164
rect 18035 14112 18087 14164
rect 18139 14112 18191 14164
rect 17931 14008 17983 14060
rect 18035 14008 18087 14060
rect 18139 14008 18191 14060
rect 10855 13397 10913 13451
rect 10993 13397 11051 13451
rect 10858 13270 10916 13324
rect 10997 13268 11055 13322
rect 10857 13117 10915 13171
rect 10997 13126 11055 13180
rect 11397 12650 11457 12710
rect 11581 12647 11641 12707
rect 11394 12522 11454 12582
rect 11579 12514 11639 12574
rect 11395 12377 11455 12437
rect 11572 12377 11632 12437
rect 12268 12362 12326 12416
rect 12406 12362 12464 12416
rect 12271 12235 12329 12289
rect 12410 12233 12468 12287
rect 12270 12082 12328 12136
rect 12410 12091 12468 12145
rect 8605 11605 8665 11665
rect 8727 11606 8787 11666
rect 8872 11609 8932 11669
rect 8611 11493 8671 11553
rect 8742 11494 8802 11554
rect 8881 11494 8941 11554
rect 11340 9923 11400 9983
rect 11517 9934 11577 9994
rect 11274 9792 11334 9852
rect 11410 9802 11470 9862
rect 11557 9797 11617 9857
rect 11436 7926 11496 7986
rect 11570 7926 11630 7986
rect 11431 7812 11491 7872
rect 11560 7800 11620 7860
rect 5391 7488 5451 7548
rect 5588 7504 5648 7564
rect 5727 7508 5787 7568
rect 5871 7504 5931 7564
rect 5354 7358 5414 7418
rect 5503 7363 5563 7423
rect 5676 7370 5736 7430
rect 5850 7384 5910 7444
rect 5323 7238 5383 7298
rect 5474 7246 5534 7306
rect 5637 7250 5697 7310
rect 5798 7250 5858 7310
rect 5939 7255 5999 7315
rect 12962 7249 13022 7309
rect 13098 7249 13158 7309
rect 12957 7136 13017 7196
rect 13093 7129 13153 7189
rect 8594 7012 8654 7072
rect 8737 7012 8797 7072
rect 8949 7017 9009 7077
rect 8594 6900 8654 6960
rect 8742 6900 8802 6960
rect 8980 6900 9040 6960
rect 12498 5336 12558 5396
rect 12675 5347 12735 5407
rect 12432 5205 12492 5265
rect 12568 5215 12628 5275
rect 12715 5210 12775 5270
rect 4824 -1046 4884 -986
rect 4988 -1048 5048 -988
rect 4824 -1173 4884 -1113
rect 4990 -1160 5050 -1100
rect 4824 -1311 4884 -1251
rect 4995 -1300 5055 -1240
rect 4890 -1625 4950 -1565
rect 5056 -1612 5116 -1552
rect 4890 -1763 4950 -1703
rect 5061 -1752 5121 -1692
rect 4792 -2309 4852 -2249
rect 4543 -2412 4603 -2352
rect 4683 -2412 4743 -2352
rect 4545 -2533 4605 -2473
rect 4691 -2536 4751 -2476
rect 4811 -2541 4871 -2481
rect 5047 -2721 5107 -2661
rect 5213 -2708 5273 -2648
rect 5047 -2859 5107 -2799
rect 5218 -2848 5278 -2788
rect 4951 -3139 5011 -3079
rect 5117 -3126 5177 -3066
rect 4951 -3277 5011 -3217
rect 5122 -3266 5182 -3206
rect 4928 -3553 4988 -3493
rect 5094 -3540 5154 -3480
rect 4928 -3691 4988 -3631
rect 5099 -3680 5159 -3620
rect 4974 -4032 5034 -3972
rect 5140 -4019 5200 -3959
rect 4974 -4170 5034 -4110
rect 5145 -4159 5205 -4099
rect 5079 -4575 5139 -4515
rect 5245 -4562 5305 -4502
rect 5079 -4713 5139 -4653
rect 5250 -4702 5310 -4642
rect 17919 13891 17971 13943
rect 18023 13891 18075 13943
rect 18127 13891 18179 13943
rect 17919 13787 17971 13839
rect 18023 13787 18075 13839
rect 18127 13787 18179 13839
rect 19222 14062 19274 14114
rect 19326 14062 19378 14114
rect 19222 13958 19274 14010
rect 19326 13958 19378 14010
rect 19222 13854 19274 13906
rect 19326 13854 19378 13906
rect 20393 14039 20445 14091
rect 20497 14039 20549 14091
rect 20601 14039 20653 14091
rect 20393 13935 20445 13987
rect 20497 13935 20549 13987
rect 20601 13935 20653 13987
rect 22114 13926 22275 14087
rect 22497 13927 22656 14086
rect 22915 13926 23076 14087
rect 37931 14102 37991 14162
rect 38051 14102 38111 14162
rect 38171 14102 38231 14162
rect 38291 14102 38351 14162
rect 38411 14102 38471 14162
rect 37931 13982 37991 14042
rect 38051 13982 38111 14042
rect 38171 13982 38231 14042
rect 38291 13982 38351 14042
rect 38411 13982 38471 14042
rect 20393 13831 20445 13883
rect 20497 13831 20549 13883
rect 20601 13831 20653 13883
rect 19222 13750 19274 13802
rect 19326 13750 19378 13802
rect 21964 13522 22100 13658
rect 22388 13523 22522 13657
rect 22678 13522 22814 13658
rect 21813 13162 21915 13264
rect 22053 13163 22153 13263
rect 22385 13162 22487 13264
rect 29826 13269 29886 13329
rect 29946 13269 30006 13329
rect 30066 13269 30126 13329
rect 30186 13269 30246 13329
rect 30306 13269 30366 13329
rect 29826 13149 29886 13209
rect 29946 13149 30006 13209
rect 30066 13149 30126 13209
rect 30186 13149 30246 13209
rect 30306 13149 30366 13209
rect 19666 11132 19726 11192
rect 19907 11137 19967 11197
rect 20146 11139 20206 11199
rect 20373 11139 20433 11199
rect 22477 11111 22537 11171
rect 22472 10967 22532 11027
rect 64920 13711 64990 13781
rect 65179 13707 65249 13777
rect 65420 13642 65490 13712
rect 64924 13560 64994 13630
rect 65191 13530 65261 13600
rect 65415 13489 65485 13559
rect 64923 13391 64993 13461
rect 65181 13393 65251 13463
rect 65413 13346 65483 13416
rect 64973 13216 65043 13286
rect 65175 13211 65245 13281
rect 65338 13199 65408 13269
rect 41720 12547 41843 12670
rect 41719 12296 41844 12421
rect 41720 12073 41843 12196
rect 37873 10728 37933 10788
rect 37993 10728 38053 10788
rect 38113 10728 38173 10788
rect 38233 10728 38293 10788
rect 38353 10728 38413 10788
rect 37873 10608 37933 10668
rect 37993 10608 38053 10668
rect 38113 10608 38173 10668
rect 38233 10608 38293 10668
rect 38353 10608 38413 10668
rect 28780 9837 28840 9897
rect 29021 9842 29081 9902
rect 29260 9844 29320 9904
rect 29487 9844 29547 9904
rect 19624 9086 19684 9146
rect 19865 9091 19925 9151
rect 20104 9093 20164 9153
rect 20331 9093 20391 9153
rect 22935 7818 22995 7878
rect 23176 7823 23236 7883
rect 23415 7825 23475 7885
rect 23642 7825 23702 7885
rect 28724 6843 28784 6903
rect 28965 6848 29025 6908
rect 29204 6850 29264 6910
rect 29431 6850 29491 6910
rect 22102 6705 22219 6822
rect 22399 6706 22514 6821
rect 18068 6614 18128 6674
rect 18188 6614 18248 6674
rect 18308 6614 18368 6674
rect 18428 6614 18488 6674
rect 18548 6614 18608 6674
rect 18668 6614 18728 6674
rect 18788 6614 18848 6674
rect 18908 6614 18968 6674
rect 19028 6614 19088 6674
rect 19148 6614 19208 6674
rect 19268 6614 19328 6674
rect 19388 6614 19448 6674
rect 32070 9822 32132 9884
rect 47780 8163 47858 8241
rect 47935 8162 48015 8242
rect 54010 9256 54070 9320
rect 54130 9316 54190 9320
rect 54250 9319 54310 9320
rect 54129 9260 54190 9316
rect 54246 9260 54310 9319
rect 54370 9260 54430 9320
rect 54490 9319 54550 9320
rect 54487 9260 54550 9319
rect 54129 9256 54189 9260
rect 54246 9259 54306 9260
rect 54487 9259 54547 9260
rect 54251 9200 54311 9202
rect 54371 9200 54431 9206
rect 54010 9140 54070 9200
rect 54128 9140 54190 9200
rect 54250 9142 54311 9200
rect 54370 9146 54431 9200
rect 54490 9199 54550 9200
rect 54250 9140 54310 9142
rect 54370 9140 54430 9146
rect 54489 9140 54550 9199
rect 54489 9139 54549 9140
rect 61580 9263 61640 9327
rect 61700 9323 61760 9327
rect 61820 9326 61880 9327
rect 61699 9267 61760 9323
rect 61816 9267 61880 9326
rect 61940 9267 62000 9327
rect 62060 9326 62120 9327
rect 62057 9267 62120 9326
rect 61699 9263 61759 9267
rect 61816 9266 61876 9267
rect 62057 9266 62117 9267
rect 61821 9207 61881 9209
rect 61941 9207 62001 9213
rect 61580 9147 61640 9207
rect 61698 9147 61760 9207
rect 61820 9149 61881 9207
rect 61940 9153 62001 9207
rect 62060 9206 62120 9207
rect 61820 9147 61880 9149
rect 61940 9147 62000 9153
rect 62059 9147 62120 9206
rect 62059 9146 62119 9147
rect 43278 6941 43448 7111
rect 43821 6941 43991 7111
rect 44532 6942 44700 7110
rect 46183 7008 46259 7086
rect 46429 7003 46505 7081
rect 46709 7005 46785 7083
rect 46925 7013 47001 7091
rect 39317 6427 39523 6633
rect 43813 6009 43889 6087
rect 44062 5996 44138 6074
rect 44296 5991 44372 6069
rect 44518 5995 44594 6073
rect 27111 4315 27239 4443
rect 27342 4314 27472 4444
rect 30434 4399 30559 4524
rect 27107 4118 27237 4248
rect 27343 4119 27471 4247
rect 30435 4139 30558 4262
rect 53784 4602 53844 4666
rect 53904 4662 53964 4666
rect 54024 4665 54084 4666
rect 53903 4606 53964 4662
rect 54020 4606 54084 4665
rect 54144 4606 54204 4666
rect 54264 4665 54324 4666
rect 54261 4606 54324 4665
rect 53903 4602 53963 4606
rect 54020 4605 54080 4606
rect 54261 4605 54321 4606
rect 54025 4546 54085 4548
rect 54145 4546 54205 4552
rect 53784 4486 53844 4546
rect 53902 4486 53964 4546
rect 54024 4488 54085 4546
rect 54144 4492 54205 4546
rect 54264 4545 54324 4546
rect 54024 4486 54084 4488
rect 54144 4486 54204 4492
rect 54263 4486 54324 4545
rect 54263 4485 54323 4486
rect 98886 4666 98945 4721
rect 99061 4660 99120 4715
rect 98884 4507 98943 4562
rect 99062 4511 99121 4566
rect 98887 4342 98946 4397
rect 99075 4337 99134 4392
rect 91416 4195 91476 4259
rect 91536 4255 91596 4259
rect 91656 4258 91716 4259
rect 91535 4199 91596 4255
rect 91652 4199 91716 4258
rect 91776 4199 91836 4259
rect 91896 4258 91956 4259
rect 91893 4199 91956 4258
rect 91535 4195 91595 4199
rect 91652 4198 91712 4199
rect 91893 4198 91953 4199
rect 91657 4139 91717 4141
rect 91777 4139 91837 4145
rect 91416 4079 91476 4139
rect 91534 4079 91596 4139
rect 91656 4081 91717 4139
rect 91776 4085 91837 4139
rect 91896 4138 91956 4139
rect 91656 4079 91716 4081
rect 91776 4079 91836 4085
rect 91895 4079 91956 4138
rect 91895 4078 91955 4079
rect 95232 2610 95292 2670
rect 95352 2610 95412 2670
rect 95472 2610 95532 2670
rect 95232 2490 95292 2550
rect 95352 2490 95412 2550
rect 95472 2490 95532 2550
rect 95232 2370 95292 2430
rect 95352 2370 95412 2430
rect 95472 2370 95532 2430
rect 90003 -370 90063 -310
rect 90127 -358 90187 -298
rect 90021 -487 90081 -427
rect 90145 -499 90205 -439
rect 18108 -1628 18235 -1515
rect 18415 -1623 18542 -1510
rect 18665 -1616 18792 -1503
rect 58356 -3095 58411 -3036
rect 58526 -3070 58581 -3011
rect 58355 -3269 58410 -3210
rect 58521 -3268 58576 -3209
rect 68215 -3694 68274 -3639
rect 68389 -3695 68448 -3640
rect 68216 -3860 68275 -3805
rect 68414 -3865 68473 -3810
rect 98599 -815 98658 -760
rect 98774 -821 98833 -766
rect 98597 -974 98656 -919
rect 98775 -970 98834 -915
rect 98600 -1139 98659 -1084
rect 98788 -1144 98847 -1089
rect 98632 -2019 98691 -1964
rect 98806 -2020 98865 -1965
rect 98633 -2185 98692 -2130
rect 98831 -2190 98890 -2135
rect 98602 -2916 98661 -2861
rect 98776 -2917 98835 -2862
rect 98603 -3082 98662 -3027
rect 98801 -3087 98860 -3032
rect 98594 -3399 98653 -3344
rect 98768 -3400 98827 -3345
rect 98595 -3565 98654 -3510
rect 98793 -3570 98852 -3515
rect 98632 -3951 98691 -3896
rect 98806 -3952 98865 -3897
rect 98633 -4117 98692 -4062
rect 98831 -4122 98890 -4067
rect 87132 -4780 87192 -4720
rect 87252 -4780 87312 -4720
rect 87372 -4780 87432 -4720
rect 87132 -4900 87192 -4840
rect 87252 -4900 87312 -4840
rect 87372 -4900 87432 -4840
rect 87132 -5020 87192 -4960
rect 87252 -5020 87312 -4960
rect 87372 -5020 87432 -4960
rect 48442 -9397 48502 -9337
rect 48581 -9409 48641 -9349
rect 48436 -9513 48496 -9453
rect 48584 -9534 48644 -9474
rect 48439 -9627 48499 -9567
rect 48584 -9650 48644 -9590
rect 52344 -11450 52404 -11390
rect 52549 -11437 52609 -11377
rect 52804 -11435 52864 -11375
rect 53073 -11427 53133 -11367
rect 53315 -11424 53375 -11364
rect 52346 -11640 52406 -11580
rect 52552 -11632 52612 -11572
rect 52785 -11622 52845 -11562
rect 53030 -11619 53090 -11559
rect 53243 -11607 53303 -11547
rect 53402 -11606 53462 -11546
rect 52337 -11816 52397 -11756
rect 52505 -11815 52565 -11755
rect 52703 -11813 52763 -11753
rect 52914 -11810 52974 -11750
rect 53153 -11800 53213 -11740
rect 53351 -11792 53411 -11732
rect 49195 -14212 49255 -14152
rect 49315 -14212 49375 -14152
rect 49435 -14212 49495 -14152
rect 49195 -14332 49255 -14272
rect 49315 -14332 49375 -14272
rect 49435 -14332 49495 -14272
rect 98602 -7530 98662 -7470
rect 98722 -7530 98782 -7470
rect 98842 -7530 98902 -7470
rect 98602 -7650 98662 -7590
rect 98722 -7650 98782 -7590
rect 98842 -7650 98902 -7590
rect 98602 -7770 98662 -7710
rect 98722 -7770 98782 -7710
rect 98842 -7770 98902 -7710
<< metal2 >>
rect -3079 62802 -2804 62816
rect -3079 62742 -3054 62802
rect -2994 62800 -2804 62802
rect -2994 62742 -2890 62800
rect -3079 62740 -2890 62742
rect -2830 62740 -2804 62800
rect -3079 62688 -2804 62740
rect -3079 62675 -2888 62688
rect -3079 62615 -3054 62675
rect -2994 62628 -2888 62675
rect -2828 62628 -2804 62688
rect -2994 62615 -2804 62628
rect -3079 62548 -2804 62615
rect -3079 62537 -2883 62548
rect -3079 62477 -3054 62537
rect -2994 62488 -2883 62537
rect -2823 62488 -2804 62548
rect -2994 62477 -2804 62488
rect -3079 62466 -2804 62477
rect -4059 61374 -3689 61414
rect -4059 61361 -3847 61374
rect -4059 61301 -4013 61361
rect -3953 61314 -3847 61361
rect -3787 61314 -3689 61374
rect -3953 61301 -3689 61314
rect -4059 61234 -3689 61301
rect -4059 61223 -3842 61234
rect -4059 61163 -4013 61223
rect -3953 61174 -3842 61223
rect -3782 61174 -3689 61234
rect -3953 61163 -3689 61174
rect -4059 61136 -3689 61163
rect -2698 52730 -2423 52744
rect -2698 52670 -2673 52730
rect -2613 52728 -2423 52730
rect -2613 52670 -2509 52728
rect -2698 52668 -2509 52670
rect -2449 52668 -2423 52728
rect -2698 52616 -2423 52668
rect -2698 52603 -2507 52616
rect -2698 52543 -2673 52603
rect -2613 52556 -2507 52603
rect -2447 52556 -2423 52616
rect -2613 52543 -2423 52556
rect -2698 52476 -2423 52543
rect -2698 52465 -2502 52476
rect -2698 52405 -2673 52465
rect -2613 52416 -2502 52465
rect -2442 52416 -2423 52476
rect -2613 52405 -2423 52416
rect -2698 52394 -2423 52405
rect -3907 52218 -3537 52258
rect -3907 52205 -3695 52218
rect -3907 52145 -3861 52205
rect -3801 52158 -3695 52205
rect -3635 52158 -3537 52218
rect -3801 52145 -3537 52158
rect -3907 52078 -3537 52145
rect -3907 52067 -3690 52078
rect -3907 52007 -3861 52067
rect -3801 52018 -3690 52067
rect -3630 52018 -3537 52078
rect -3801 52007 -3537 52018
rect -3907 51980 -3537 52007
rect -2388 44204 -2113 44218
rect -2388 44144 -2363 44204
rect -2303 44202 -2113 44204
rect -2303 44144 -2199 44202
rect -2388 44142 -2199 44144
rect -2139 44142 -2113 44202
rect -2388 44090 -2113 44142
rect -2388 44077 -2197 44090
rect -2388 44017 -2363 44077
rect -2303 44030 -2197 44077
rect -2137 44030 -2113 44090
rect -2303 44017 -2113 44030
rect -2388 43950 -2113 44017
rect -2388 43939 -2192 43950
rect -2388 43879 -2363 43939
rect -2303 43890 -2192 43939
rect -2132 43890 -2113 43950
rect -2303 43879 -2113 43890
rect -2388 43868 -2113 43879
rect -2381 43663 -2106 43677
rect -2381 43603 -2356 43663
rect -2296 43661 -2106 43663
rect -2296 43603 -2192 43661
rect -2381 43601 -2192 43603
rect -2132 43601 -2106 43661
rect -2381 43549 -2106 43601
rect -2381 43536 -2190 43549
rect -2381 43476 -2356 43536
rect -2296 43489 -2190 43536
rect -2130 43489 -2106 43549
rect -2296 43476 -2106 43489
rect -2381 43409 -2106 43476
rect -2381 43398 -2185 43409
rect -2381 43338 -2356 43398
rect -2296 43349 -2185 43398
rect -2125 43349 -2106 43409
rect -2296 43338 -2106 43349
rect -2381 43327 -2106 43338
rect -2489 36770 -2214 36784
rect -2489 36710 -2464 36770
rect -2404 36768 -2214 36770
rect -2404 36710 -2300 36768
rect -2489 36708 -2300 36710
rect -2240 36708 -2214 36768
rect -2489 36656 -2214 36708
rect -2489 36643 -2298 36656
rect -2489 36583 -2464 36643
rect -2404 36596 -2298 36643
rect -2238 36596 -2214 36656
rect -2404 36583 -2214 36596
rect -2489 36516 -2214 36583
rect -2489 36505 -2293 36516
rect -2489 36445 -2464 36505
rect -2404 36456 -2293 36505
rect -2233 36456 -2214 36516
rect -2404 36445 -2214 36456
rect -2489 36434 -2214 36445
rect 2010 28029 2740 28118
rect 2010 28021 2605 28029
rect 2010 27961 2039 28021
rect 2099 28018 2415 28021
rect 2099 27961 2218 28018
rect 2010 27958 2218 27961
rect 2278 27961 2415 28018
rect 2475 27969 2605 28021
rect 2665 27969 2740 28029
rect 2475 27961 2740 27969
rect 2278 27958 2740 27961
rect 2010 27894 2740 27958
rect 2010 27834 2042 27894
rect 2102 27886 2605 27894
rect 2102 27883 2407 27886
rect 2102 27834 2218 27883
rect 2010 27823 2218 27834
rect 2278 27826 2407 27883
rect 2467 27834 2605 27886
rect 2665 27834 2740 27894
rect 2467 27826 2740 27834
rect 2278 27823 2740 27826
rect 2010 27720 2740 27823
rect -3588 25044 -3261 25051
rect -3592 24984 -3575 25044
rect -3515 24984 -3455 25044
rect -3395 24984 -3335 25044
rect -3275 25043 -3165 25044
rect -3275 24984 -1026 25043
rect -3592 24951 -1026 24984
rect -3592 24924 -464 24951
rect -3592 24864 -3575 24924
rect -3515 24864 -3455 24924
rect -3395 24864 -3335 24924
rect -3275 24864 -464 24924
rect -3592 24840 -464 24864
rect -3592 24804 -1026 24840
rect -3592 24744 -3575 24804
rect -3515 24744 -3455 24804
rect -3395 24744 -3335 24804
rect -3275 24748 -1026 24804
rect -3275 24744 -3165 24748
rect -3592 24732 -3165 24744
rect -1775 20749 -1405 23311
rect 8582 21782 9071 21859
rect 8582 21762 8972 21782
rect 8582 21696 8757 21762
rect 8829 21716 8972 21762
rect 9044 21716 9071 21782
rect 8829 21696 9071 21716
rect 8582 21609 9071 21696
rect 8582 21599 8908 21609
rect 8582 21533 8646 21599
rect 8718 21543 8908 21599
rect 8980 21543 9071 21609
rect 8718 21533 9071 21543
rect 8582 21358 9071 21533
rect 8582 21348 8884 21358
rect 8582 21282 8664 21348
rect 8736 21292 8884 21348
rect 8956 21292 9071 21358
rect 8736 21282 9071 21292
rect 8582 21236 9071 21282
rect -265 20749 1066 20974
rect -1794 20716 1066 20749
rect -1794 20696 369 20716
rect -1794 20630 154 20696
rect 226 20650 369 20696
rect 441 20650 1066 20716
rect 226 20630 1066 20650
rect -1794 20543 1066 20630
rect -1794 20533 305 20543
rect -1794 20467 43 20533
rect 115 20477 305 20533
rect 377 20477 1066 20543
rect 115 20467 1066 20477
rect -1794 20340 1066 20467
rect -265 20292 1066 20340
rect -265 20282 281 20292
rect -265 20216 61 20282
rect 133 20226 281 20282
rect 353 20226 1066 20292
rect 133 20216 1066 20226
rect -265 19888 1066 20216
rect 2458 16522 2515 16888
rect -198 15447 -142 15448
rect -298 15391 -132 15447
rect -198 15252 -142 15391
rect 2503 15111 2561 15299
rect 1122 14386 1678 14442
rect 2080 14352 2136 14528
rect 919 13812 975 14048
rect 1943 11782 1999 12188
rect 8582 11731 8987 21236
rect 41677 20265 44259 20474
rect 9800 17600 10310 17660
rect 9800 17540 9832 17600
rect 9892 17540 9960 17600
rect 10020 17597 10310 17600
rect 10020 17540 10111 17597
rect 9800 17537 10111 17540
rect 10171 17537 10310 17597
rect 9800 17470 10310 17537
rect 9800 17441 21600 17470
rect 9800 17381 9830 17441
rect 9890 17439 10177 17441
rect 9890 17381 10001 17439
rect 9800 17379 10001 17381
rect 10061 17381 10177 17439
rect 10237 17381 21600 17441
rect 10061 17379 21600 17381
rect 9800 17278 21600 17379
rect 9800 17262 10193 17278
rect 9800 17257 10044 17262
rect 9800 17197 9842 17257
rect 9902 17202 10044 17257
rect 10104 17218 10193 17262
rect 10253 17250 21600 17278
rect 10253 17218 10310 17250
rect 10104 17202 10310 17218
rect 9902 17197 10310 17202
rect 9800 17160 10310 17197
rect 9750 16937 10260 16990
rect 9750 16930 10050 16937
rect 9750 16927 9919 16930
rect 9750 16867 9791 16927
rect 9851 16870 9919 16927
rect 9979 16877 10050 16930
rect 10110 16914 10260 16937
rect 10110 16877 20684 16914
rect 9979 16870 20684 16877
rect 9851 16867 20684 16870
rect 9750 16753 20684 16867
rect 9750 16748 10103 16753
rect 9750 16730 9955 16748
rect 9750 16670 9786 16730
rect 9846 16688 9955 16730
rect 10015 16693 10103 16748
rect 10163 16693 20684 16753
rect 10015 16688 20684 16693
rect 9846 16670 20684 16688
rect 9750 16646 20684 16670
rect 9750 16620 10260 16646
rect 9750 16610 10137 16620
rect 9750 16579 9960 16610
rect 9750 16519 9763 16579
rect 9823 16550 9960 16579
rect 10020 16560 10137 16610
rect 10197 16560 10260 16620
rect 10020 16550 10260 16560
rect 9823 16519 10260 16550
rect 9750 16490 10260 16519
rect 12240 16138 19962 16431
rect 12240 14461 12533 16138
rect 19669 15309 19962 16138
rect 20416 15743 20684 16646
rect 21380 16095 21600 17250
rect 22731 16830 23374 16880
rect 22731 16770 22811 16830
rect 22871 16770 22931 16830
rect 22991 16770 23051 16830
rect 23111 16770 23171 16830
rect 23231 16770 23291 16830
rect 23351 16799 23374 16830
rect 23351 16770 37528 16799
rect 22731 16710 37528 16770
rect 22731 16650 22811 16710
rect 22871 16650 22931 16710
rect 22991 16650 23051 16710
rect 23111 16650 23171 16710
rect 23231 16650 23291 16710
rect 23351 16650 37528 16710
rect 22731 16594 37528 16650
rect 22731 16591 23374 16594
rect 22735 16494 23393 16495
rect 22735 16435 36567 16494
rect 22735 16375 22818 16435
rect 22878 16375 22938 16435
rect 22998 16375 23058 16435
rect 23118 16375 23178 16435
rect 23238 16375 23298 16435
rect 23358 16375 36567 16435
rect 22735 16315 36567 16375
rect 22735 16255 22818 16315
rect 22878 16255 22938 16315
rect 22998 16255 23058 16315
rect 23118 16255 23178 16315
rect 23238 16255 23298 16315
rect 23358 16289 36567 16315
rect 23358 16255 23393 16289
rect 22735 16213 23393 16255
rect 22738 16210 23393 16213
rect 21380 16087 24210 16095
rect 21380 15884 35629 16087
rect 21380 15875 24210 15884
rect 20416 15712 24234 15743
rect 20416 15506 33629 15712
rect 20416 15475 24234 15506
rect 19669 15286 23314 15309
rect 19669 15254 31910 15286
rect 19669 15194 22090 15254
rect 22150 15194 22210 15254
rect 22270 15194 22330 15254
rect 22390 15194 22450 15254
rect 22510 15194 22570 15254
rect 22630 15194 31910 15254
rect 19669 15134 31910 15194
rect 10823 14168 12533 14461
rect 12941 14846 19271 15094
rect 19669 15074 22090 15134
rect 22150 15074 22210 15134
rect 22270 15074 22330 15134
rect 22390 15074 22450 15134
rect 22510 15074 22570 15134
rect 22630 15074 31910 15134
rect 19669 15039 31910 15074
rect 19669 15016 23314 15039
rect 10823 13451 11116 14168
rect 10823 13397 10855 13451
rect 10913 13397 10993 13451
rect 11051 13397 11116 13451
rect 10823 13324 11116 13397
rect 10823 13270 10858 13324
rect 10916 13322 11116 13324
rect 10916 13270 10997 13322
rect 10823 13268 10997 13270
rect 11055 13268 11116 13322
rect 10823 13180 11116 13268
rect 10823 13171 10997 13180
rect 10823 13117 10857 13171
rect 10915 13126 10997 13171
rect 11055 13126 11116 13180
rect 10915 13117 11116 13126
rect 10823 13099 11116 13117
rect 11365 12710 11683 12801
rect 11365 12650 11397 12710
rect 11457 12707 11683 12710
rect 11457 12650 11581 12707
rect 11365 12647 11581 12650
rect 11641 12647 11683 12707
rect 11365 12582 11683 12647
rect 11365 12522 11394 12582
rect 11454 12574 11683 12582
rect 11454 12522 11579 12574
rect 11365 12514 11579 12522
rect 11639 12514 11683 12574
rect 11365 12437 11683 12514
rect 11365 12377 11395 12437
rect 11455 12377 11572 12437
rect 11632 12377 11683 12437
rect 11365 12334 11683 12377
rect 12236 12459 12529 12469
rect 12236 12416 12533 12459
rect 12236 12362 12268 12416
rect 12326 12362 12406 12416
rect 12464 12362 12533 12416
rect 12236 12289 12533 12362
rect 12236 12235 12271 12289
rect 12329 12287 12533 12289
rect 12329 12235 12410 12287
rect 12236 12233 12410 12235
rect 12468 12233 12533 12287
rect 12236 12145 12533 12233
rect 12236 12136 12410 12145
rect 12236 12082 12270 12136
rect 12328 12091 12410 12136
rect 12468 12091 12533 12145
rect 12328 12082 12533 12091
rect 12236 12064 12533 12082
rect 8578 11669 8995 11731
rect 8578 11666 8871 11669
rect 8578 11665 8725 11666
rect 8578 11605 8605 11665
rect 8665 11606 8725 11665
rect 8787 11609 8871 11666
rect 8932 11609 8995 11669
rect 8787 11606 8995 11609
rect 8665 11605 8995 11606
rect 8578 11554 8995 11605
rect 8578 11494 8610 11554
rect 8670 11553 8741 11554
rect 8671 11494 8741 11553
rect 8802 11494 8881 11554
rect 8941 11494 8995 11554
rect 8578 11493 8611 11494
rect 8671 11493 8995 11494
rect 8578 11488 8995 11493
rect 11239 10062 11632 10070
rect 12240 10062 12533 12064
rect 11238 10056 12533 10062
rect 11236 9994 12533 10056
rect 11236 9983 11517 9994
rect 11236 9923 11340 9983
rect 11400 9934 11517 9983
rect 11577 9934 12533 9994
rect 11400 9923 12533 9934
rect 11236 9862 12533 9923
rect 11236 9852 11410 9862
rect 11236 9792 11274 9852
rect 11334 9802 11410 9852
rect 11470 9857 12533 9862
rect 11470 9802 11557 9857
rect 11334 9797 11557 9802
rect 11617 9797 12533 9857
rect 11334 9792 12533 9797
rect 11236 9772 12533 9792
rect 11238 9769 12533 9772
rect 12941 8826 13189 14846
rect 19023 14678 19271 14846
rect 22059 14694 22659 14696
rect 22045 14678 22661 14694
rect 19023 14636 30057 14678
rect 19023 14576 22059 14636
rect 22119 14576 22179 14636
rect 22239 14576 22299 14636
rect 22359 14576 22419 14636
rect 22479 14576 22539 14636
rect 22599 14576 30057 14636
rect 19023 14516 30057 14576
rect 19023 14456 22059 14516
rect 22119 14456 22179 14516
rect 22239 14456 22299 14516
rect 22359 14456 22419 14516
rect 22479 14456 22539 14516
rect 22599 14456 30057 14516
rect 19023 14430 30057 14456
rect 22045 14427 22661 14430
rect 17357 14268 18262 14318
rect 17357 14216 17931 14268
rect 17983 14216 18035 14268
rect 18087 14216 18139 14268
rect 18191 14216 18262 14268
rect 17357 14185 18262 14216
rect 17357 14165 17787 14185
rect 17357 14099 17572 14165
rect 17644 14119 17787 14165
rect 17859 14164 18262 14185
rect 17859 14119 17931 14164
rect 17644 14112 17931 14119
rect 17983 14112 18035 14164
rect 18087 14117 18139 14164
rect 18120 14112 18139 14117
rect 18191 14112 18262 14164
rect 17644 14099 18048 14112
rect 17357 14060 18048 14099
rect 18120 14060 18262 14112
rect 17357 14012 17931 14060
rect 17357 14002 17723 14012
rect 17357 13936 17461 14002
rect 17533 13946 17723 14002
rect 17795 14008 17931 14012
rect 17983 14008 18035 14060
rect 18120 14051 18139 14060
rect 18087 14008 18139 14051
rect 18191 14008 18262 14060
rect 17795 13950 18262 14008
rect 17795 13946 17912 13950
rect 17533 13936 17912 13946
rect 17984 13943 18262 13950
rect 17357 13884 17912 13936
rect 17984 13891 18023 13943
rect 18075 13891 18127 13943
rect 18179 13891 18262 13943
rect 17984 13884 18262 13891
rect 17357 13839 18262 13884
rect 17357 13787 17919 13839
rect 17971 13787 18023 13839
rect 18075 13787 18127 13839
rect 18179 13787 18262 13839
rect 17357 13761 18262 13787
rect 17357 13751 17699 13761
rect 17357 13685 17479 13751
rect 17551 13695 17699 13751
rect 17771 13700 18262 13761
rect 19198 14114 19410 14168
rect 19198 14062 19222 14114
rect 19274 14062 19326 14114
rect 19378 14062 19410 14114
rect 19198 14010 19410 14062
rect 19198 13958 19222 14010
rect 19274 13958 19326 14010
rect 19378 13958 19410 14010
rect 19198 13906 19410 13958
rect 19198 13854 19222 13906
rect 19274 13854 19326 13906
rect 19378 13854 19410 13906
rect 19198 13802 19410 13854
rect 19198 13750 19222 13802
rect 19274 13750 19326 13802
rect 19378 13750 19410 13802
rect 20130 14145 20656 14238
rect 20130 14109 20725 14145
rect 20130 14099 20472 14109
rect 20130 14033 20252 14099
rect 20324 14091 20472 14099
rect 20544 14091 20725 14109
rect 20324 14039 20393 14091
rect 20445 14043 20472 14091
rect 20445 14039 20497 14043
rect 20549 14039 20601 14091
rect 20653 14039 20725 14091
rect 20324 14033 20725 14039
rect 20130 13987 20725 14033
rect 20130 13935 20393 13987
rect 20445 13935 20497 13987
rect 20549 13935 20601 13987
rect 20653 13935 20725 13987
rect 20130 13910 20725 13935
rect 20130 13844 20243 13910
rect 20315 13904 20725 13910
rect 22087 14087 23144 14135
rect 22087 13926 22114 14087
rect 22275 14086 22915 14087
rect 22275 13927 22497 14086
rect 22656 13927 22915 14086
rect 22275 13926 22915 13927
rect 23076 13926 28904 14087
rect 22087 13904 23144 13926
rect 20315 13883 20470 13904
rect 20542 13883 20725 13904
rect 20315 13844 20393 13883
rect 20130 13831 20393 13844
rect 20445 13838 20470 13883
rect 20445 13831 20497 13838
rect 20549 13831 20601 13883
rect 20653 13831 20725 13883
rect 20130 13787 20725 13831
rect 19198 13738 19410 13750
rect 17771 13695 17916 13700
rect 17551 13685 17916 13695
rect 17357 13634 17916 13685
rect 17988 13634 18262 13700
rect 17357 13556 18262 13634
rect 11423 8578 13189 8826
rect 13467 13461 13922 13516
rect 17357 13490 17697 13556
rect 17769 13490 18262 13556
rect 17357 13461 18262 13490
rect 13467 13285 18262 13461
rect 13467 13116 18226 13285
rect 11423 7986 11671 8578
rect 11423 7926 11436 7986
rect 11496 7926 11570 7986
rect 11630 7926 11671 7986
rect 11423 7872 11671 7926
rect 11423 7812 11431 7872
rect 11491 7860 11671 7872
rect 11491 7812 11560 7860
rect 11423 7800 11560 7812
rect 11620 7800 11671 7860
rect 11423 7781 11671 7800
rect 5268 7568 6063 7709
rect 5268 7564 5727 7568
rect 5268 7548 5588 7564
rect 5268 7488 5391 7548
rect 5451 7504 5588 7548
rect 5648 7508 5727 7564
rect 5787 7564 6063 7568
rect 5787 7508 5871 7564
rect 5648 7504 5871 7508
rect 5931 7504 6063 7564
rect 5451 7488 6063 7504
rect 5268 7444 6063 7488
rect 5268 7430 5850 7444
rect 5268 7423 5676 7430
rect 5268 7418 5503 7423
rect 5268 7358 5354 7418
rect 5414 7363 5503 7418
rect 5563 7370 5676 7423
rect 5736 7384 5850 7430
rect 5910 7384 6063 7444
rect 5736 7370 6063 7384
rect 5563 7363 6063 7370
rect 5414 7358 6063 7363
rect 5268 7315 6063 7358
rect 5268 7310 5939 7315
rect 5268 7306 5637 7310
rect 5268 7298 5474 7306
rect 5268 7238 5323 7298
rect 5383 7246 5474 7298
rect 5534 7250 5637 7306
rect 5697 7250 5798 7310
rect 5858 7255 5939 7310
rect 5999 7255 6063 7315
rect 5858 7250 6063 7255
rect 5534 7246 6063 7250
rect 5383 7238 6063 7246
rect 5268 7226 6063 7238
rect 12940 7309 13192 7311
rect 12940 7249 12962 7309
rect 13022 7249 13098 7309
rect 13158 7249 13192 7309
rect 12940 7196 13192 7249
rect 8560 7077 9108 7137
rect 12940 7136 12957 7196
rect 13017 7189 13192 7196
rect 13017 7136 13093 7189
rect 12940 7129 13093 7136
rect 13153 7129 13192 7189
rect 12940 7111 13192 7129
rect 8560 7072 8949 7077
rect 8560 7070 8594 7072
rect 8654 7070 8737 7072
rect 8560 7010 8588 7070
rect 8654 7012 8729 7070
rect 8797 7017 8949 7072
rect 9009 7017 9108 7077
rect 8797 7012 9108 7017
rect 8648 7010 8729 7012
rect 8789 7010 9108 7012
rect 8560 6960 9108 7010
rect 8560 6900 8594 6960
rect 8654 6955 8742 6960
rect 8802 6955 8980 6960
rect 8654 6900 8735 6955
rect 8802 6900 8975 6955
rect 9040 6900 9108 6960
rect 8560 6895 8735 6900
rect 8795 6895 8975 6900
rect 9035 6895 9108 6900
rect 8560 6879 9108 6895
rect 12397 5486 12483 5488
rect 12397 5469 12848 5486
rect 12382 5466 12848 5469
rect 12941 5466 13189 7111
rect 12382 5407 13189 5466
rect 12382 5396 12675 5407
rect 12382 5336 12498 5396
rect 12558 5347 12675 5396
rect 12735 5347 13189 5407
rect 12558 5336 13189 5347
rect 12382 5275 13189 5336
rect 12382 5265 12568 5275
rect 12382 5205 12432 5265
rect 12492 5215 12568 5265
rect 12628 5270 13189 5275
rect 12628 5215 12715 5270
rect 12492 5210 12715 5215
rect 12775 5218 13189 5270
rect 12775 5210 12848 5218
rect 12492 5205 12848 5210
rect 12382 5176 12848 5205
rect 4778 -986 5148 -932
rect 4778 -1046 4824 -986
rect 4884 -988 5148 -986
rect 4884 -1046 4988 -988
rect 4778 -1048 4988 -1046
rect 5048 -1048 5148 -988
rect 4778 -1100 5148 -1048
rect 4778 -1113 4990 -1100
rect 4778 -1173 4824 -1113
rect 4884 -1160 4990 -1113
rect 5050 -1160 5148 -1100
rect 4884 -1173 5148 -1160
rect 4778 -1240 5148 -1173
rect 4778 -1251 4995 -1240
rect 4778 -1311 4824 -1251
rect 4884 -1300 4995 -1251
rect 5055 -1300 5148 -1240
rect 4884 -1311 5148 -1300
rect 4778 -1338 5148 -1311
rect 4844 -1552 5214 -1512
rect 4844 -1565 5056 -1552
rect 4844 -1625 4890 -1565
rect 4950 -1612 5056 -1565
rect 5116 -1612 5214 -1552
rect 4950 -1625 5214 -1612
rect 4844 -1692 5214 -1625
rect 4844 -1703 5061 -1692
rect 4844 -1763 4890 -1703
rect 4950 -1752 5061 -1703
rect 5121 -1752 5214 -1692
rect 4950 -1763 5214 -1752
rect 4844 -1790 5214 -1763
rect 4506 -2249 4874 -2240
rect 4506 -2309 4792 -2249
rect 4852 -2255 4874 -2249
rect 4852 -2309 11467 -2255
rect 4506 -2352 11467 -2309
rect 4506 -2412 4543 -2352
rect 4603 -2412 4683 -2352
rect 4743 -2412 11467 -2352
rect 4506 -2455 11467 -2412
rect 4506 -2473 4874 -2455
rect 4506 -2533 4545 -2473
rect 4605 -2476 4874 -2473
rect 4605 -2533 4691 -2476
rect 4506 -2536 4691 -2533
rect 4751 -2481 4874 -2476
rect 4751 -2536 4811 -2481
rect 4506 -2541 4811 -2536
rect 4871 -2541 4874 -2481
rect 4506 -2563 4874 -2541
rect 5001 -2648 5371 -2608
rect 5001 -2661 5213 -2648
rect 5001 -2721 5047 -2661
rect 5107 -2708 5213 -2661
rect 5273 -2708 5371 -2648
rect 5107 -2721 5371 -2708
rect 5001 -2788 5371 -2721
rect 5001 -2799 5218 -2788
rect 5001 -2859 5047 -2799
rect 5107 -2848 5218 -2799
rect 5278 -2848 5371 -2788
rect 5107 -2859 5371 -2848
rect 5001 -2886 5371 -2859
rect 4905 -3066 5275 -3026
rect 4905 -3079 5117 -3066
rect 4905 -3139 4951 -3079
rect 5011 -3126 5117 -3079
rect 5177 -3126 5275 -3066
rect 5011 -3139 5275 -3126
rect 4905 -3206 5275 -3139
rect 4905 -3217 5122 -3206
rect 4905 -3277 4951 -3217
rect 5011 -3266 5122 -3217
rect 5182 -3266 5275 -3206
rect 5011 -3277 5275 -3266
rect 4905 -3304 5275 -3277
rect 4882 -3480 5252 -3440
rect 4882 -3493 5094 -3480
rect 4882 -3553 4928 -3493
rect 4988 -3540 5094 -3493
rect 5154 -3540 5252 -3480
rect 4988 -3553 5252 -3540
rect 4882 -3620 5252 -3553
rect 4882 -3631 5099 -3620
rect 4882 -3691 4928 -3631
rect 4988 -3680 5099 -3631
rect 5159 -3680 5252 -3620
rect 4988 -3691 5252 -3680
rect 4882 -3718 5252 -3691
rect 11285 -3874 11467 -2455
rect 13467 -3380 13922 13116
rect 17908 12969 18198 13116
rect 19228 12977 19380 13738
rect 20406 12980 20725 13787
rect 21938 13658 22849 13700
rect 25430 13658 26138 13671
rect 21938 13522 21964 13658
rect 22100 13657 22678 13658
rect 22100 13523 22388 13657
rect 22522 13523 22678 13657
rect 22100 13522 22678 13523
rect 22814 13642 26138 13658
rect 22814 13538 25496 13642
rect 25600 13538 25684 13642
rect 25788 13538 25879 13642
rect 25983 13538 26138 13642
rect 22814 13522 26138 13538
rect 21938 13497 22849 13522
rect 25430 13504 26138 13522
rect 25430 13503 26015 13504
rect 21799 13290 22548 13292
rect 21799 13264 25263 13290
rect 21799 13162 21813 13264
rect 21915 13263 22385 13264
rect 21915 13163 22053 13263
rect 22153 13163 22385 13263
rect 21915 13162 22385 13163
rect 22487 13162 25263 13264
rect 21799 13142 25263 13162
rect 22003 13130 25263 13142
rect 17908 12820 18711 12969
rect 19228 12825 19543 12977
rect 19391 12008 19543 12825
rect 20406 12807 22149 12980
rect 21976 12098 22149 12807
rect 25103 12633 25263 13130
rect 25103 12473 28368 12633
rect 21863 11925 22149 12098
rect 27026 11727 27558 11886
rect 28208 11854 28368 12473
rect 28743 12234 28904 13926
rect 29809 13377 30057 14430
rect 29808 13329 30422 13377
rect 29808 13269 29826 13329
rect 29886 13269 29946 13329
rect 30006 13269 30066 13329
rect 30126 13269 30186 13329
rect 30246 13269 30306 13329
rect 30366 13269 30422 13329
rect 29808 13209 30422 13269
rect 29808 13149 29826 13209
rect 29886 13149 29946 13209
rect 30006 13149 30066 13209
rect 30126 13149 30186 13209
rect 30246 13149 30306 13209
rect 30366 13149 30422 13209
rect 29808 13140 30422 13149
rect 28743 12073 30776 12234
rect 30615 11894 30776 12073
rect 27026 11650 27185 11727
rect 28208 11694 30139 11854
rect 30615 11733 30983 11894
rect 26304 11491 27236 11650
rect 19654 11192 19738 11204
rect 19654 11132 19666 11192
rect 19726 11132 19738 11192
rect 19654 11121 19738 11132
rect 19895 11197 19979 11209
rect 19895 11137 19907 11197
rect 19967 11137 19979 11197
rect 19895 11126 19979 11137
rect 20120 11199 20230 11220
rect 20120 11139 20146 11199
rect 20206 11139 20230 11199
rect 20120 11110 20230 11139
rect 20361 11199 20445 11211
rect 20361 11139 20373 11199
rect 20433 11139 20445 11199
rect 20361 11128 20445 11139
rect 22449 11208 22560 11220
rect 22449 11171 22574 11208
rect 21983 11113 22080 11125
rect 22449 11113 22477 11171
rect 21983 11111 22477 11113
rect 22537 11111 22574 11171
rect 21983 11072 22574 11111
rect 21983 11027 22575 11072
rect 21983 10967 22472 11027
rect 22532 10967 22575 11027
rect 21983 10919 22575 10967
rect 21984 10918 22575 10919
rect 27077 11032 27236 11491
rect 27077 10873 27324 11032
rect 29660 10913 29767 11694
rect 30822 10849 30983 11733
rect 31663 9951 31910 15039
rect 33423 12307 33629 15506
rect 33149 12101 33629 12307
rect 33423 11895 33629 12101
rect 28768 9897 28852 9909
rect 28768 9837 28780 9897
rect 28840 9837 28852 9897
rect 28768 9826 28852 9837
rect 29009 9902 29093 9914
rect 29009 9842 29021 9902
rect 29081 9842 29093 9902
rect 29009 9831 29093 9842
rect 29248 9904 29332 9916
rect 29248 9844 29260 9904
rect 29320 9844 29332 9904
rect 29248 9833 29332 9844
rect 29475 9904 29559 9916
rect 29475 9844 29487 9904
rect 29547 9844 29559 9904
rect 29475 9833 29559 9844
rect 30909 9884 32327 9951
rect 35426 9902 35629 15884
rect 36362 11499 36567 16289
rect 37323 12528 37528 16594
rect 41677 15783 41886 20265
rect 37851 14162 38494 14212
rect 37851 14102 37931 14162
rect 37991 14102 38051 14162
rect 38111 14102 38171 14162
rect 38231 14102 38291 14162
rect 38351 14102 38411 14162
rect 38471 14102 38494 14162
rect 37851 14042 38494 14102
rect 37851 13982 37931 14042
rect 37991 13982 38051 14042
rect 38111 13982 38171 14042
rect 38231 13982 38291 14042
rect 38351 13982 38411 14042
rect 38471 13982 38494 14042
rect 37851 13923 38494 13982
rect 37852 10840 37971 13923
rect 38108 10840 38227 13923
rect 38374 10840 38493 13923
rect 41677 12670 41885 15783
rect 64769 13781 65603 13916
rect 64769 13711 64920 13781
rect 64990 13777 65603 13781
rect 64990 13711 65179 13777
rect 64769 13707 65179 13711
rect 65249 13759 65603 13777
rect 65249 13712 71106 13759
rect 65249 13707 65420 13712
rect 64769 13642 65420 13707
rect 65490 13642 71106 13712
rect 64769 13630 71106 13642
rect 64769 13560 64924 13630
rect 64994 13600 71106 13630
rect 64994 13560 65191 13600
rect 64769 13530 65191 13560
rect 65261 13559 71106 13600
rect 65261 13530 65415 13559
rect 64769 13489 65415 13530
rect 65485 13489 71106 13559
rect 64769 13463 71106 13489
rect 64769 13461 65181 13463
rect 64769 13391 64923 13461
rect 64993 13393 65181 13461
rect 65251 13416 71106 13463
rect 65251 13393 65413 13416
rect 64993 13391 65413 13393
rect 64769 13346 65413 13391
rect 65483 13346 71106 13416
rect 64769 13318 71106 13346
rect 64769 13286 65603 13318
rect 64769 13216 64973 13286
rect 65043 13281 65603 13286
rect 65043 13216 65175 13281
rect 64769 13211 65175 13216
rect 65245 13269 65603 13281
rect 65245 13211 65338 13269
rect 64769 13199 65338 13211
rect 65408 13199 65603 13269
rect 64769 13020 65603 13199
rect 39735 12603 41562 12604
rect 39735 12349 41564 12603
rect 37793 10788 38571 10840
rect 37793 10728 37873 10788
rect 37933 10728 37993 10788
rect 38053 10728 38113 10788
rect 38173 10728 38233 10788
rect 38293 10728 38353 10788
rect 38413 10728 38571 10788
rect 37793 10668 38571 10728
rect 37793 10608 37873 10668
rect 37933 10608 37993 10668
rect 38053 10608 38113 10668
rect 38173 10608 38233 10668
rect 38293 10608 38353 10668
rect 38413 10608 38571 10668
rect 37793 10547 38571 10608
rect 38124 10314 38319 10344
rect 30909 9822 32070 9884
rect 32132 9822 32327 9884
rect 30909 9794 32327 9822
rect 34743 9821 35629 9902
rect 31663 9749 31910 9794
rect 32011 9792 32327 9794
rect 32170 9693 32327 9792
rect 35426 9791 35629 9821
rect 38116 9812 38319 10314
rect 35450 9784 35605 9791
rect 35021 9697 35271 9715
rect 34756 9668 35271 9697
rect 34756 9620 35439 9668
rect 34858 9581 35439 9620
rect 38116 9581 38311 9812
rect 34858 9492 38311 9581
rect 29769 9190 31596 9392
rect 35150 9389 38311 9492
rect 35367 9386 38311 9389
rect 41307 9609 41564 12349
rect 41677 12547 41720 12670
rect 41843 12547 41885 12670
rect 41677 12421 41885 12547
rect 41677 12296 41719 12421
rect 41844 12296 41885 12421
rect 41677 12214 41885 12296
rect 41677 12196 42058 12214
rect 41677 12073 41720 12196
rect 41843 12073 42058 12196
rect 41677 12061 42058 12073
rect 19612 9146 19696 9158
rect 19612 9086 19624 9146
rect 19684 9086 19696 9146
rect 19612 9075 19696 9086
rect 19853 9151 19937 9163
rect 19853 9091 19865 9151
rect 19925 9091 19937 9151
rect 19853 9080 19937 9091
rect 20060 9153 20200 9180
rect 20060 9093 20104 9153
rect 20164 9093 20200 9153
rect 20060 9070 20200 9093
rect 20319 9153 20403 9165
rect 20319 9093 20331 9153
rect 20391 9093 20403 9153
rect 20319 9082 20403 9093
rect 26250 8881 27154 9033
rect 29769 8898 29971 9190
rect 30473 9034 30883 9048
rect 30473 9021 30665 9034
rect 30473 8961 30533 9021
rect 30593 8974 30665 9021
rect 30725 9033 30883 9034
rect 30725 8974 30790 9033
rect 30593 8973 30790 8974
rect 30850 8973 30883 9033
rect 30593 8961 30883 8973
rect 30473 8924 30883 8961
rect 30473 8908 30663 8924
rect 21824 8205 22125 8362
rect 19342 7505 19505 8018
rect 21968 7600 22125 8205
rect 27002 8017 27154 8881
rect 29614 8696 30098 8898
rect 30473 8848 30530 8908
rect 30590 8864 30663 8908
rect 30723 8864 30790 8924
rect 30850 8864 30883 8924
rect 30590 8848 30883 8864
rect 30473 8797 30883 8848
rect 30473 8795 30652 8797
rect 30473 8735 30527 8795
rect 30587 8737 30652 8795
rect 30712 8737 30790 8797
rect 30850 8737 30883 8797
rect 30587 8735 30883 8737
rect 30473 8717 30883 8735
rect 22923 7878 23007 7890
rect 22923 7818 22935 7878
rect 22995 7818 23007 7878
rect 22923 7807 23007 7818
rect 23164 7883 23248 7895
rect 23164 7823 23176 7883
rect 23236 7823 23248 7883
rect 23164 7812 23248 7823
rect 23403 7885 23487 7897
rect 23403 7825 23415 7885
rect 23475 7825 23487 7885
rect 23403 7814 23487 7825
rect 23630 7885 23714 7897
rect 23630 7825 23642 7885
rect 23702 7825 23714 7885
rect 27002 7865 27262 8017
rect 23630 7814 23714 7825
rect 19076 7342 19505 7505
rect 21969 7489 22125 7600
rect 21177 7488 22125 7489
rect 19076 6748 19239 7342
rect 20972 7320 22125 7488
rect 17938 6711 19507 6748
rect 17938 6674 19508 6711
rect 17938 6614 18068 6674
rect 18128 6614 18188 6674
rect 18248 6614 18308 6674
rect 18368 6614 18428 6674
rect 18488 6614 18548 6674
rect 18608 6614 18668 6674
rect 18728 6614 18788 6674
rect 18848 6614 18908 6674
rect 18968 6614 19028 6674
rect 19088 6614 19148 6674
rect 19208 6614 19268 6674
rect 19328 6614 19388 6674
rect 19448 6614 19508 6674
rect 17938 6585 19508 6614
rect 20972 6253 21508 7320
rect 22095 6822 26596 6907
rect 28712 6903 28796 6915
rect 28712 6843 28724 6903
rect 28784 6843 28796 6903
rect 28712 6832 28796 6843
rect 28953 6908 29037 6920
rect 28953 6848 28965 6908
rect 29025 6848 29037 6908
rect 28953 6837 29037 6848
rect 29192 6910 29276 6922
rect 29192 6850 29204 6910
rect 29264 6850 29276 6910
rect 29192 6839 29276 6850
rect 29419 6910 29503 6922
rect 29419 6850 29431 6910
rect 29491 6850 29503 6910
rect 29419 6839 29503 6850
rect 22095 6791 22102 6822
rect 22083 6707 22102 6791
rect 22085 6705 22102 6707
rect 22219 6821 26596 6822
rect 22219 6706 22399 6821
rect 22514 6706 26596 6821
rect 22219 6705 26596 6706
rect 22085 6683 22546 6705
rect 20972 5718 22844 6253
rect 18271 -745 18995 -726
rect 18271 -858 18296 -745
rect 18423 -858 18995 -745
rect 18271 -887 18995 -858
rect 18271 -906 18760 -887
rect 18271 -1019 18501 -906
rect 18628 -1000 18760 -906
rect 18887 -1000 18995 -887
rect 18628 -1019 18995 -1000
rect 18271 -1063 18995 -1019
rect 18080 -1502 18860 -1470
rect 18080 -1503 18671 -1502
rect 18080 -1510 18665 -1503
rect 18080 -1515 18415 -1510
rect 18542 -1515 18665 -1510
rect 18080 -1628 18108 -1515
rect 18235 -1623 18415 -1515
rect 18544 -1616 18665 -1515
rect 18798 -1615 18860 -1502
rect 18792 -1616 18860 -1615
rect 18235 -1628 18417 -1623
rect 18544 -1628 18860 -1616
rect 18080 -1660 18860 -1628
rect 22309 -2588 22844 5718
rect 26394 5828 26596 6705
rect 31394 5828 31596 9190
rect 38043 7647 38298 9386
rect 41307 9354 48122 9609
rect 47867 8256 48122 9354
rect 53921 9320 54794 9377
rect 53921 9256 54010 9320
rect 54070 9316 54130 9320
rect 54190 9319 54250 9320
rect 54070 9256 54129 9316
rect 54190 9260 54246 9319
rect 54189 9259 54246 9260
rect 54310 9260 54370 9320
rect 54430 9319 54490 9320
rect 54430 9260 54487 9319
rect 54306 9259 54487 9260
rect 54550 9260 54794 9320
rect 54547 9259 54794 9260
rect 54189 9256 54794 9259
rect 53921 9206 54794 9256
rect 53921 9202 54371 9206
rect 53921 9200 54251 9202
rect 53921 9140 54010 9200
rect 54070 9140 54128 9200
rect 54190 9140 54250 9200
rect 54311 9200 54371 9202
rect 54311 9142 54370 9200
rect 54431 9200 54794 9206
rect 54431 9199 54490 9200
rect 54431 9146 54489 9199
rect 54310 9140 54370 9142
rect 54430 9140 54489 9146
rect 53921 9139 54489 9140
rect 54550 9140 54794 9200
rect 54549 9139 54794 9140
rect 53921 9088 54794 9139
rect 61491 9327 62361 9385
rect 61491 9263 61580 9327
rect 61640 9323 61700 9327
rect 61760 9326 61820 9327
rect 61640 9263 61699 9323
rect 61760 9267 61816 9326
rect 61759 9266 61816 9267
rect 61880 9267 61940 9327
rect 62000 9326 62060 9327
rect 62000 9267 62057 9326
rect 61876 9266 62057 9267
rect 62120 9267 62361 9327
rect 62117 9266 62361 9267
rect 61759 9263 62361 9266
rect 61491 9213 62361 9263
rect 61491 9209 61941 9213
rect 61491 9207 61821 9209
rect 61491 9147 61580 9207
rect 61640 9147 61698 9207
rect 61760 9147 61820 9207
rect 61881 9207 61941 9209
rect 61881 9149 61940 9207
rect 62001 9207 62361 9213
rect 62001 9206 62060 9207
rect 62001 9153 62059 9206
rect 61880 9147 61940 9149
rect 62000 9147 62059 9153
rect 61491 9146 62059 9147
rect 62120 9147 62361 9207
rect 62119 9146 62361 9147
rect 61491 9099 62361 9146
rect 47615 8252 48122 8256
rect 47615 8242 48258 8252
rect 47615 8241 47935 8242
rect 47615 8163 47780 8241
rect 47858 8163 47935 8241
rect 47615 8162 47935 8163
rect 48015 8162 48258 8242
rect 47615 8150 48258 8162
rect 47690 8137 48258 8150
rect 47690 7940 48260 8137
rect 47852 7647 48122 7648
rect 38043 7392 48122 7647
rect 44110 7124 44460 7130
rect 43227 7111 44715 7124
rect 43227 6941 43278 7111
rect 43448 6941 43821 7111
rect 43991 6941 44531 7111
rect 44701 6941 44715 7111
rect 46136 7091 47059 7119
rect 46136 7086 46925 7091
rect 46136 7008 46183 7086
rect 46259 7083 46925 7086
rect 46259 7081 46709 7083
rect 46259 7008 46429 7081
rect 46136 7003 46429 7008
rect 46505 7005 46709 7081
rect 46785 7013 46925 7083
rect 47001 7013 47059 7091
rect 47852 7063 48122 7392
rect 46785 7005 47059 7013
rect 46505 7003 47059 7005
rect 46136 6961 47059 7003
rect 43227 6919 44715 6941
rect 44110 6850 44480 6919
rect 44110 6810 44460 6850
rect 38263 6633 39669 6671
rect 38263 6430 38287 6633
rect 38493 6427 39317 6633
rect 39523 6427 39669 6633
rect 38287 6418 39669 6427
rect 38287 6414 38493 6418
rect 43759 6087 44718 6127
rect 43759 6009 43813 6087
rect 43889 6074 44718 6087
rect 43889 6009 44062 6074
rect 43759 5996 44062 6009
rect 44138 6073 44718 6074
rect 44138 6069 44518 6073
rect 44138 5996 44296 6069
rect 43759 5991 44296 5996
rect 44372 5995 44518 6069
rect 44594 5995 44718 6073
rect 44372 5991 44718 5995
rect 43759 5971 44718 5991
rect 26394 5626 31596 5828
rect 30400 4524 30604 4659
rect 47853 4548 48122 7063
rect 98848 4724 99160 4739
rect 27094 4444 27485 4463
rect 27094 4314 27110 4444
rect 27240 4314 27342 4444
rect 27472 4314 27485 4444
rect 27094 4248 27485 4314
rect 27094 4118 27107 4248
rect 27237 4118 27342 4248
rect 27472 4118 27485 4248
rect 30400 4399 30434 4524
rect 30559 4399 30604 4524
rect 30400 4263 30604 4399
rect 45792 4279 48122 4548
rect 53695 4666 54568 4724
rect 53695 4602 53784 4666
rect 53844 4662 53904 4666
rect 53964 4665 54024 4666
rect 53844 4602 53903 4662
rect 53964 4606 54020 4665
rect 53963 4605 54020 4606
rect 54084 4606 54144 4666
rect 54204 4665 54264 4666
rect 54204 4606 54261 4665
rect 54080 4605 54261 4606
rect 54324 4606 54568 4666
rect 54321 4605 54568 4606
rect 53963 4602 54568 4605
rect 53695 4552 54568 4602
rect 53695 4548 54145 4552
rect 53695 4546 54025 4548
rect 53695 4486 53784 4546
rect 53844 4486 53902 4546
rect 53964 4486 54024 4546
rect 54085 4546 54145 4548
rect 54085 4488 54144 4546
rect 54205 4546 54568 4552
rect 54205 4545 54264 4546
rect 54205 4492 54263 4545
rect 54084 4486 54144 4488
rect 54204 4486 54263 4492
rect 53695 4485 54263 4486
rect 54324 4486 54568 4546
rect 54323 4485 54568 4486
rect 53695 4412 54568 4485
rect 98848 4666 98886 4724
rect 98948 4718 99160 4724
rect 98948 4666 99061 4718
rect 98848 4660 99061 4666
rect 99123 4660 99160 4718
rect 98848 4569 99160 4660
rect 98848 4565 99062 4569
rect 98848 4507 98884 4565
rect 98946 4511 99062 4565
rect 99124 4511 99160 4569
rect 98946 4507 99160 4511
rect 53695 4319 54344 4412
rect 53701 4315 54344 4319
rect 98848 4400 99160 4507
rect 98848 4342 98887 4400
rect 98949 4395 99160 4400
rect 98949 4342 99075 4395
rect 98848 4337 99075 4342
rect 99137 4337 99160 4395
rect 53701 4314 54194 4315
rect 30400 4138 30434 4263
rect 30559 4138 30604 4263
rect 30400 4129 30604 4138
rect 91327 4259 92059 4316
rect 98848 4305 99160 4337
rect 91327 4195 91416 4259
rect 91476 4255 91536 4259
rect 91596 4258 91656 4259
rect 91476 4195 91535 4255
rect 91596 4199 91652 4258
rect 91595 4198 91652 4199
rect 91716 4199 91776 4259
rect 91836 4258 91896 4259
rect 91836 4199 91893 4258
rect 91712 4198 91893 4199
rect 91956 4199 92059 4259
rect 91953 4198 92059 4199
rect 91595 4195 92059 4198
rect 91327 4145 92059 4195
rect 91327 4141 91777 4145
rect 91327 4139 91657 4141
rect 27094 4108 27485 4118
rect 91327 4079 91416 4139
rect 91476 4079 91534 4139
rect 91596 4079 91656 4139
rect 91717 4139 91777 4141
rect 91717 4081 91776 4139
rect 91837 4139 92059 4145
rect 91837 4138 91896 4139
rect 91837 4085 91895 4138
rect 91716 4079 91776 4081
rect 91836 4079 91895 4085
rect 91327 4078 91895 4079
rect 91956 4079 92059 4139
rect 91955 4078 92059 4079
rect 91327 4051 92059 4078
rect 95080 2785 95620 2970
rect 95080 2670 96818 2785
rect 95080 2610 95232 2670
rect 95292 2610 95352 2670
rect 95412 2610 95472 2670
rect 95532 2610 96818 2670
rect 95080 2550 96818 2610
rect 95080 2490 95232 2550
rect 95292 2490 95352 2550
rect 95412 2490 95472 2550
rect 95532 2490 96818 2550
rect 95080 2430 96818 2490
rect 95080 2370 95232 2430
rect 95292 2370 95352 2430
rect 95412 2370 95472 2430
rect 95532 2390 96818 2430
rect 95532 2370 95620 2390
rect 95080 2270 95620 2370
rect 94369 368 94922 651
rect 89933 -298 90316 -240
rect 89933 -310 90127 -298
rect 89933 -317 90003 -310
rect 86599 -370 90003 -317
rect 90063 -358 90127 -310
rect 90187 -358 90316 -298
rect 90063 -370 90316 -358
rect 86599 -427 90316 -370
rect 86599 -487 90021 -427
rect 90081 -439 90316 -427
rect 90081 -487 90145 -439
rect 86599 -499 90145 -487
rect 90205 -499 90316 -439
rect 86599 -523 90316 -499
rect 89933 -570 90316 -523
rect 22309 -3123 47333 -2588
rect 58344 -3008 58612 -2964
rect 58344 -3033 58523 -3008
rect 58344 -3095 58353 -3033
rect 58411 -3070 58523 -3033
rect 58581 -3070 58612 -3008
rect 58411 -3095 58612 -3070
rect 13467 -3705 17126 -3380
rect 17805 -3874 17987 -3316
rect 4928 -3959 5298 -3919
rect 4928 -3972 5140 -3959
rect 4928 -4032 4974 -3972
rect 5034 -4019 5140 -3972
rect 5200 -4019 5298 -3959
rect 5034 -4032 5298 -4019
rect 4928 -4099 5298 -4032
rect 11285 -4056 17987 -3874
rect 11296 -4081 17960 -4056
rect 4928 -4110 5145 -4099
rect 4928 -4170 4974 -4110
rect 5034 -4159 5145 -4110
rect 5205 -4159 5298 -4099
rect 5034 -4170 5298 -4159
rect 4928 -4197 5298 -4170
rect 5033 -4502 5403 -4462
rect 5033 -4515 5245 -4502
rect 5033 -4575 5079 -4515
rect 5139 -4562 5245 -4515
rect 5305 -4562 5403 -4502
rect 5139 -4575 5403 -4562
rect 5033 -4642 5403 -4575
rect 5033 -4653 5250 -4642
rect 5033 -4713 5079 -4653
rect 5139 -4702 5250 -4653
rect 5310 -4702 5403 -4642
rect 5139 -4713 5403 -4702
rect 5033 -4740 5403 -4713
rect 46962 -5017 47332 -3123
rect 58344 -3206 58612 -3095
rect 58344 -3207 58518 -3206
rect 58344 -3269 58352 -3207
rect 58410 -3268 58518 -3207
rect 58576 -3268 58612 -3206
rect 58410 -3269 58612 -3268
rect 58344 -3325 58612 -3269
rect 68159 -3636 68520 -3628
rect 68159 -3694 68215 -3636
rect 68277 -3637 68520 -3636
rect 68277 -3694 68389 -3637
rect 68159 -3695 68389 -3694
rect 68451 -3695 68520 -3637
rect 68159 -3802 68520 -3695
rect 68159 -3860 68216 -3802
rect 68278 -3807 68520 -3802
rect 68278 -3860 68414 -3807
rect 68159 -3865 68414 -3860
rect 68476 -3865 68520 -3807
rect 68159 -3896 68520 -3865
rect 87090 -4720 87760 -4550
rect 87090 -4780 87130 -4720
rect 87192 -4780 87250 -4720
rect 87312 -4780 87370 -4720
rect 87432 -4780 87760 -4720
rect 87090 -4840 87760 -4780
rect 87090 -4900 87130 -4840
rect 87192 -4900 87250 -4840
rect 87312 -4900 87370 -4840
rect 87432 -4900 87760 -4840
rect 87090 -4960 87760 -4900
rect 45298 -5387 48300 -5017
rect 87090 -5020 87132 -4960
rect 87192 -5020 87250 -4960
rect 87312 -5020 87370 -4960
rect 87432 -5020 87760 -4960
rect 87090 -5090 87760 -5020
rect 47930 -9293 48300 -5387
rect 94639 -7468 94922 368
rect 96448 -5325 96818 2390
rect 98561 -757 98873 -742
rect 98561 -815 98599 -757
rect 98661 -763 98873 -757
rect 98661 -815 98774 -763
rect 98561 -821 98774 -815
rect 98836 -821 98873 -763
rect 98561 -912 98873 -821
rect 98561 -916 98775 -912
rect 98561 -974 98597 -916
rect 98659 -970 98775 -916
rect 98837 -970 98873 -912
rect 98659 -974 98873 -970
rect 98561 -1081 98873 -974
rect 98561 -1139 98600 -1081
rect 98662 -1086 98873 -1081
rect 98662 -1139 98788 -1086
rect 98561 -1144 98788 -1139
rect 98850 -1144 98873 -1086
rect 98561 -1181 98873 -1144
rect 98576 -1961 98937 -1953
rect 98576 -2019 98632 -1961
rect 98694 -1962 98937 -1961
rect 98694 -2019 98806 -1962
rect 98576 -2020 98806 -2019
rect 98868 -2020 98937 -1962
rect 98576 -2127 98937 -2020
rect 98576 -2185 98633 -2127
rect 98695 -2132 98937 -2127
rect 98695 -2185 98831 -2132
rect 98576 -2190 98831 -2185
rect 98893 -2190 98937 -2132
rect 98576 -2221 98937 -2190
rect 98546 -2858 98907 -2850
rect 98546 -2916 98602 -2858
rect 98664 -2859 98907 -2858
rect 98664 -2916 98776 -2859
rect 98546 -2917 98776 -2916
rect 98838 -2917 98907 -2859
rect 98546 -3024 98907 -2917
rect 98546 -3082 98603 -3024
rect 98665 -3029 98907 -3024
rect 98665 -3082 98801 -3029
rect 98546 -3087 98801 -3082
rect 98863 -3087 98907 -3029
rect 98546 -3118 98907 -3087
rect 98538 -3341 98899 -3333
rect 98538 -3399 98594 -3341
rect 98656 -3342 98899 -3341
rect 98656 -3399 98768 -3342
rect 98538 -3400 98768 -3399
rect 98830 -3400 98899 -3342
rect 98538 -3507 98899 -3400
rect 98538 -3565 98595 -3507
rect 98657 -3512 98899 -3507
rect 98657 -3565 98793 -3512
rect 98538 -3570 98793 -3565
rect 98855 -3570 98899 -3512
rect 98538 -3601 98899 -3570
rect 98576 -3893 98937 -3885
rect 98576 -3951 98632 -3893
rect 98694 -3894 98937 -3893
rect 98694 -3951 98806 -3894
rect 98576 -3952 98806 -3951
rect 98868 -3952 98937 -3894
rect 98576 -4059 98937 -3952
rect 98576 -4117 98633 -4059
rect 98695 -4064 98937 -4059
rect 98695 -4117 98831 -4064
rect 98576 -4122 98831 -4117
rect 98893 -4122 98937 -4064
rect 98576 -4153 98937 -4122
rect 98574 -7468 98910 -7460
rect 94639 -7470 98910 -7468
rect 94639 -7530 98602 -7470
rect 98662 -7530 98722 -7470
rect 98782 -7530 98842 -7470
rect 98902 -7530 98910 -7470
rect 94639 -7590 98910 -7530
rect 94639 -7650 98602 -7590
rect 98662 -7650 98722 -7590
rect 98782 -7650 98842 -7590
rect 98902 -7650 98910 -7590
rect 94639 -7710 98910 -7650
rect 94639 -7751 98602 -7710
rect 98574 -7770 98602 -7751
rect 98662 -7770 98722 -7710
rect 98782 -7770 98842 -7710
rect 98902 -7770 98910 -7710
rect 98574 -7800 98910 -7770
rect 47930 -9337 48775 -9293
rect 47930 -9397 48442 -9337
rect 48502 -9349 48775 -9337
rect 48502 -9397 48581 -9349
rect 47930 -9409 48581 -9397
rect 48641 -9409 48775 -9349
rect 47930 -9453 48775 -9409
rect 47930 -9513 48436 -9453
rect 48496 -9474 48775 -9453
rect 48496 -9513 48584 -9474
rect 47930 -9534 48584 -9513
rect 48644 -9534 48775 -9474
rect 47930 -9567 48775 -9534
rect 47930 -9627 48439 -9567
rect 48499 -9590 48775 -9567
rect 48499 -9627 48584 -9590
rect 47930 -9650 48584 -9627
rect 48644 -9650 48775 -9590
rect 47930 -9663 48775 -9650
rect 52279 -11322 53565 -11166
rect 52279 -11364 53571 -11322
rect 52279 -11367 53315 -11364
rect 52279 -11375 53073 -11367
rect 52279 -11377 52804 -11375
rect 52279 -11390 52549 -11377
rect 52279 -11450 52344 -11390
rect 52404 -11437 52549 -11390
rect 52609 -11435 52804 -11377
rect 52864 -11427 53073 -11375
rect 53133 -11424 53315 -11367
rect 53375 -11424 53571 -11364
rect 53133 -11427 53571 -11424
rect 52864 -11435 53571 -11427
rect 52609 -11437 53571 -11435
rect 52404 -11450 53571 -11437
rect 52279 -11546 53571 -11450
rect 52279 -11547 53402 -11546
rect 52279 -11559 53243 -11547
rect 52279 -11562 53030 -11559
rect 52279 -11572 52785 -11562
rect 52279 -11580 52552 -11572
rect 52279 -11640 52346 -11580
rect 52406 -11632 52552 -11580
rect 52612 -11622 52785 -11572
rect 52845 -11619 53030 -11562
rect 53090 -11607 53243 -11559
rect 53303 -11606 53402 -11547
rect 53462 -11606 53571 -11546
rect 53303 -11607 53571 -11606
rect 53090 -11619 53571 -11607
rect 52845 -11622 53571 -11619
rect 52612 -11632 53571 -11622
rect 52406 -11640 53571 -11632
rect 52279 -11732 53571 -11640
rect 52279 -11740 53351 -11732
rect 52279 -11750 53153 -11740
rect 52279 -11753 52914 -11750
rect 52279 -11755 52703 -11753
rect 52279 -11756 52505 -11755
rect 52279 -11816 52337 -11756
rect 52397 -11815 52505 -11756
rect 52565 -11813 52703 -11755
rect 52763 -11810 52914 -11753
rect 52974 -11800 53153 -11750
rect 53213 -11792 53351 -11740
rect 53411 -11792 53571 -11732
rect 53213 -11800 53571 -11792
rect 52974 -11810 53571 -11800
rect 52763 -11813 53571 -11810
rect 52565 -11815 53571 -11813
rect 52397 -11816 53571 -11815
rect 52279 -11848 53571 -11816
rect 48991 -14152 49554 -14074
rect 48991 -14212 49195 -14152
rect 49255 -14212 49315 -14152
rect 49375 -14212 49435 -14152
rect 49495 -14212 49554 -14152
rect 48991 -14272 49554 -14212
rect 48991 -14332 49195 -14272
rect 49255 -14332 49315 -14272
rect 49375 -14332 49435 -14272
rect 49495 -14332 49554 -14272
rect 48991 -14450 49554 -14332
<< via2 >>
rect -3054 62742 -2994 62802
rect -2890 62740 -2830 62800
rect -3054 62615 -2994 62675
rect -2888 62628 -2828 62688
rect -3054 62477 -2994 62537
rect -2883 62488 -2823 62548
rect -4013 61301 -3953 61361
rect -3847 61314 -3787 61374
rect -4013 61163 -3953 61223
rect -3842 61174 -3782 61234
rect -2673 52670 -2613 52730
rect -2509 52668 -2449 52728
rect -2673 52543 -2613 52603
rect -2507 52556 -2447 52616
rect -2673 52405 -2613 52465
rect -2502 52416 -2442 52476
rect -3861 52145 -3801 52205
rect -3695 52158 -3635 52218
rect -3861 52007 -3801 52067
rect -3690 52018 -3630 52078
rect -2363 44144 -2303 44204
rect -2199 44142 -2139 44202
rect -2363 44017 -2303 44077
rect -2197 44030 -2137 44090
rect -2363 43879 -2303 43939
rect -2192 43890 -2132 43950
rect -2356 43603 -2296 43663
rect -2192 43601 -2132 43661
rect -2356 43476 -2296 43536
rect -2190 43489 -2130 43549
rect -2356 43338 -2296 43398
rect -2185 43349 -2125 43409
rect -2464 36710 -2404 36770
rect -2300 36708 -2240 36768
rect -2464 36583 -2404 36643
rect -2298 36596 -2238 36656
rect -2464 36445 -2404 36505
rect -2293 36456 -2233 36516
rect 2039 27961 2099 28021
rect 2218 27958 2278 28018
rect 2415 27961 2475 28021
rect 2605 27969 2665 28029
rect 2042 27834 2102 27894
rect 2218 27823 2278 27883
rect 2407 27826 2467 27886
rect 2605 27834 2665 27894
rect 8757 21696 8829 21762
rect 8972 21716 9044 21782
rect 8646 21533 8718 21599
rect 8908 21543 8980 21609
rect 8664 21282 8736 21348
rect 8884 21292 8956 21358
rect 154 20630 226 20696
rect 369 20650 441 20716
rect 43 20467 115 20533
rect 305 20477 377 20543
rect 61 20216 133 20282
rect 281 20226 353 20292
rect 11397 12650 11457 12710
rect 11581 12647 11641 12707
rect 11394 12522 11454 12582
rect 11579 12514 11639 12574
rect 11395 12377 11455 12437
rect 11572 12377 11632 12437
rect 8605 11605 8665 11665
rect 8725 11606 8727 11666
rect 8727 11606 8785 11666
rect 8871 11609 8872 11669
rect 8872 11609 8931 11669
rect 8610 11553 8670 11554
rect 8610 11494 8611 11553
rect 8611 11494 8670 11553
rect 8741 11494 8742 11554
rect 8742 11494 8801 11554
rect 8881 11494 8941 11554
rect 17572 14099 17644 14165
rect 17787 14119 17859 14185
rect 18048 14112 18087 14117
rect 18087 14112 18120 14117
rect 18048 14060 18120 14112
rect 17461 13936 17533 14002
rect 17723 13946 17795 14012
rect 18048 14051 18087 14060
rect 18087 14051 18120 14060
rect 17912 13943 17984 13950
rect 17912 13891 17919 13943
rect 17919 13891 17971 13943
rect 17971 13891 17984 13943
rect 17912 13884 17984 13891
rect 17479 13685 17551 13751
rect 17699 13695 17771 13761
rect 20252 14033 20324 14099
rect 20472 14091 20544 14109
rect 20472 14043 20497 14091
rect 20497 14043 20544 14091
rect 20243 13844 20315 13910
rect 20470 13883 20542 13904
rect 20470 13838 20497 13883
rect 20497 13838 20542 13883
rect 17916 13634 17988 13700
rect 17697 13490 17769 13556
rect 5391 7488 5451 7548
rect 5588 7504 5648 7564
rect 5727 7508 5787 7568
rect 5871 7504 5931 7564
rect 5354 7358 5414 7418
rect 5503 7363 5563 7423
rect 5676 7370 5736 7430
rect 5850 7384 5910 7444
rect 5323 7238 5383 7298
rect 5474 7246 5534 7306
rect 5637 7250 5697 7310
rect 5798 7250 5858 7310
rect 5939 7255 5999 7315
rect 8588 7012 8594 7070
rect 8594 7012 8648 7070
rect 8729 7012 8737 7070
rect 8737 7012 8789 7070
rect 8949 7017 9009 7077
rect 8588 7010 8648 7012
rect 8729 7010 8789 7012
rect 8594 6900 8654 6960
rect 8735 6900 8742 6955
rect 8742 6900 8795 6955
rect 8975 6900 8980 6955
rect 8980 6900 9035 6955
rect 8735 6895 8795 6900
rect 8975 6895 9035 6900
rect 4824 -1046 4884 -986
rect 4988 -1048 5048 -988
rect 4824 -1173 4884 -1113
rect 4990 -1160 5050 -1100
rect 4824 -1311 4884 -1251
rect 4995 -1300 5055 -1240
rect 4890 -1625 4950 -1565
rect 5056 -1612 5116 -1552
rect 4890 -1763 4950 -1703
rect 5061 -1752 5121 -1692
rect 5047 -2721 5107 -2661
rect 5213 -2708 5273 -2648
rect 5047 -2859 5107 -2799
rect 5218 -2848 5278 -2788
rect 4951 -3139 5011 -3079
rect 5117 -3126 5177 -3066
rect 4951 -3277 5011 -3217
rect 5122 -3266 5182 -3206
rect 4928 -3553 4988 -3493
rect 5094 -3540 5154 -3480
rect 4928 -3691 4988 -3631
rect 5099 -3680 5159 -3620
rect 25496 13538 25600 13642
rect 25684 13538 25788 13642
rect 25879 13538 25983 13642
rect 19666 11132 19726 11192
rect 19907 11137 19967 11197
rect 20146 11139 20206 11199
rect 20373 11139 20433 11199
rect 28780 9837 28840 9897
rect 29021 9842 29081 9902
rect 29260 9844 29320 9904
rect 29487 9844 29547 9904
rect 19624 9086 19684 9146
rect 19865 9091 19925 9151
rect 20104 9093 20164 9153
rect 20331 9093 20391 9153
rect 30533 8961 30593 9021
rect 30665 8974 30725 9034
rect 30790 8973 30850 9033
rect 30530 8848 30590 8908
rect 30663 8864 30723 8924
rect 30790 8864 30850 8924
rect 30527 8735 30587 8795
rect 30652 8737 30712 8797
rect 30790 8737 30850 8797
rect 22935 7818 22995 7878
rect 23176 7823 23236 7883
rect 23415 7825 23475 7885
rect 23642 7825 23702 7885
rect 28724 6843 28784 6903
rect 28965 6848 29025 6908
rect 29204 6850 29264 6910
rect 29431 6850 29491 6910
rect 18296 -858 18423 -745
rect 18501 -1019 18628 -906
rect 18760 -1000 18887 -887
rect 18671 -1503 18798 -1502
rect 18108 -1628 18235 -1515
rect 18417 -1623 18542 -1515
rect 18542 -1623 18544 -1515
rect 18671 -1615 18792 -1503
rect 18792 -1615 18798 -1503
rect 18417 -1628 18544 -1623
rect 54010 9256 54070 9316
rect 54129 9256 54189 9316
rect 54246 9259 54306 9319
rect 54370 9260 54430 9320
rect 54487 9259 54547 9319
rect 54010 9140 54070 9200
rect 54128 9140 54188 9200
rect 54251 9142 54311 9202
rect 54371 9146 54431 9206
rect 54489 9139 54549 9199
rect 61580 9263 61640 9323
rect 61699 9263 61759 9323
rect 61816 9266 61876 9326
rect 61940 9267 62000 9327
rect 62057 9266 62117 9326
rect 61580 9147 61640 9207
rect 61698 9147 61758 9207
rect 61821 9149 61881 9209
rect 61941 9153 62001 9213
rect 62059 9146 62119 9206
rect 43278 6941 43448 7111
rect 43821 6941 43991 7111
rect 44531 7110 44701 7111
rect 44531 6942 44532 7110
rect 44532 6942 44700 7110
rect 44700 6942 44701 7110
rect 44531 6941 44701 6942
rect 46183 7008 46259 7086
rect 46429 7003 46505 7081
rect 46709 7005 46785 7083
rect 46925 7013 47001 7091
rect 38287 6427 38493 6633
rect 43813 6009 43889 6087
rect 44062 5996 44138 6074
rect 44296 5991 44372 6069
rect 44518 5995 44594 6073
rect 27110 4443 27240 4444
rect 27110 4315 27111 4443
rect 27111 4315 27239 4443
rect 27239 4315 27240 4443
rect 27110 4314 27240 4315
rect 27342 4314 27472 4444
rect 27107 4118 27237 4248
rect 27342 4247 27472 4248
rect 27342 4119 27343 4247
rect 27343 4119 27471 4247
rect 27471 4119 27472 4247
rect 27342 4118 27472 4119
rect 30434 4399 30559 4524
rect 53784 4602 53844 4662
rect 53903 4602 53963 4662
rect 54020 4605 54080 4665
rect 54144 4606 54204 4666
rect 54261 4605 54321 4665
rect 53784 4486 53844 4546
rect 53902 4486 53962 4546
rect 54025 4488 54085 4548
rect 54145 4492 54205 4552
rect 54263 4485 54323 4545
rect 98886 4721 98948 4724
rect 98886 4666 98945 4721
rect 98945 4666 98948 4721
rect 99061 4715 99123 4718
rect 99061 4660 99120 4715
rect 99120 4660 99123 4715
rect 99062 4566 99124 4569
rect 98884 4562 98946 4565
rect 98884 4507 98943 4562
rect 98943 4507 98946 4562
rect 99062 4511 99121 4566
rect 99121 4511 99124 4566
rect 98887 4397 98949 4400
rect 98887 4342 98946 4397
rect 98946 4342 98949 4397
rect 99075 4392 99137 4395
rect 99075 4337 99134 4392
rect 99134 4337 99137 4392
rect 30434 4262 30559 4263
rect 30434 4139 30435 4262
rect 30435 4139 30558 4262
rect 30558 4139 30559 4262
rect 30434 4138 30559 4139
rect 91416 4195 91476 4255
rect 91535 4195 91595 4255
rect 91652 4198 91712 4258
rect 91776 4199 91836 4259
rect 91893 4198 91953 4258
rect 91416 4079 91476 4139
rect 91534 4079 91594 4139
rect 91657 4081 91717 4141
rect 91777 4085 91837 4145
rect 91895 4078 91955 4138
rect 58523 -3011 58581 -3008
rect 58353 -3036 58411 -3033
rect 58353 -3095 58356 -3036
rect 58356 -3095 58411 -3036
rect 58523 -3070 58526 -3011
rect 58526 -3070 58581 -3011
rect 4974 -4032 5034 -3972
rect 5140 -4019 5200 -3959
rect 4974 -4170 5034 -4110
rect 5145 -4159 5205 -4099
rect 5079 -4575 5139 -4515
rect 5245 -4562 5305 -4502
rect 5079 -4713 5139 -4653
rect 5250 -4702 5310 -4642
rect 58352 -3210 58410 -3207
rect 58352 -3269 58355 -3210
rect 58355 -3269 58410 -3210
rect 58518 -3209 58576 -3206
rect 58518 -3268 58521 -3209
rect 58521 -3268 58576 -3209
rect 68215 -3639 68277 -3636
rect 68215 -3694 68274 -3639
rect 68274 -3694 68277 -3639
rect 68389 -3640 68451 -3637
rect 68389 -3695 68448 -3640
rect 68448 -3695 68451 -3640
rect 68216 -3805 68278 -3802
rect 68216 -3860 68275 -3805
rect 68275 -3860 68278 -3805
rect 68414 -3810 68476 -3807
rect 68414 -3865 68473 -3810
rect 68473 -3865 68476 -3810
rect 87130 -4780 87132 -4720
rect 87132 -4780 87190 -4720
rect 87250 -4780 87252 -4720
rect 87252 -4780 87310 -4720
rect 87370 -4780 87372 -4720
rect 87372 -4780 87430 -4720
rect 87130 -4900 87132 -4840
rect 87132 -4900 87190 -4840
rect 87250 -4900 87252 -4840
rect 87252 -4900 87310 -4840
rect 87370 -4900 87372 -4840
rect 87372 -4900 87430 -4840
rect 87132 -5020 87192 -4960
rect 87250 -5020 87252 -4960
rect 87252 -5020 87310 -4960
rect 87370 -5020 87372 -4960
rect 87372 -5020 87430 -4960
rect 98599 -760 98661 -757
rect 98599 -815 98658 -760
rect 98658 -815 98661 -760
rect 98774 -766 98836 -763
rect 98774 -821 98833 -766
rect 98833 -821 98836 -766
rect 98775 -915 98837 -912
rect 98597 -919 98659 -916
rect 98597 -974 98656 -919
rect 98656 -974 98659 -919
rect 98775 -970 98834 -915
rect 98834 -970 98837 -915
rect 98600 -1084 98662 -1081
rect 98600 -1139 98659 -1084
rect 98659 -1139 98662 -1084
rect 98788 -1089 98850 -1086
rect 98788 -1144 98847 -1089
rect 98847 -1144 98850 -1089
rect 98632 -1964 98694 -1961
rect 98632 -2019 98691 -1964
rect 98691 -2019 98694 -1964
rect 98806 -1965 98868 -1962
rect 98806 -2020 98865 -1965
rect 98865 -2020 98868 -1965
rect 98633 -2130 98695 -2127
rect 98633 -2185 98692 -2130
rect 98692 -2185 98695 -2130
rect 98831 -2135 98893 -2132
rect 98831 -2190 98890 -2135
rect 98890 -2190 98893 -2135
rect 98602 -2861 98664 -2858
rect 98602 -2916 98661 -2861
rect 98661 -2916 98664 -2861
rect 98776 -2862 98838 -2859
rect 98776 -2917 98835 -2862
rect 98835 -2917 98838 -2862
rect 98603 -3027 98665 -3024
rect 98603 -3082 98662 -3027
rect 98662 -3082 98665 -3027
rect 98801 -3032 98863 -3029
rect 98801 -3087 98860 -3032
rect 98860 -3087 98863 -3032
rect 98594 -3344 98656 -3341
rect 98594 -3399 98653 -3344
rect 98653 -3399 98656 -3344
rect 98768 -3345 98830 -3342
rect 98768 -3400 98827 -3345
rect 98827 -3400 98830 -3345
rect 98595 -3510 98657 -3507
rect 98595 -3565 98654 -3510
rect 98654 -3565 98657 -3510
rect 98793 -3515 98855 -3512
rect 98793 -3570 98852 -3515
rect 98852 -3570 98855 -3515
rect 98632 -3896 98694 -3893
rect 98632 -3951 98691 -3896
rect 98691 -3951 98694 -3896
rect 98806 -3897 98868 -3894
rect 98806 -3952 98865 -3897
rect 98865 -3952 98868 -3897
rect 98633 -4062 98695 -4059
rect 98633 -4117 98692 -4062
rect 98692 -4117 98695 -4062
rect 98831 -4067 98893 -4064
rect 98831 -4122 98890 -4067
rect 98890 -4122 98893 -4067
rect 52344 -11450 52404 -11390
rect 52549 -11437 52609 -11377
rect 52804 -11435 52864 -11375
rect 53073 -11427 53133 -11367
rect 53315 -11424 53375 -11364
rect 52346 -11640 52406 -11580
rect 52552 -11632 52612 -11572
rect 52785 -11622 52845 -11562
rect 53030 -11619 53090 -11559
rect 53243 -11607 53303 -11547
rect 53402 -11606 53462 -11546
rect 52337 -11816 52397 -11756
rect 52505 -11815 52565 -11755
rect 52703 -11813 52763 -11753
rect 52914 -11810 52974 -11750
rect 53153 -11800 53213 -11740
rect 53351 -11792 53411 -11732
<< metal3 >>
rect -3079 62802 -2804 62816
rect -3079 62742 -3054 62802
rect -2994 62800 -2804 62802
rect -2994 62742 -2890 62800
rect -3079 62740 -2890 62742
rect -2830 62740 -2804 62800
rect -3079 62739 -2804 62740
rect -3089 62688 7594 62739
rect -3089 62675 -2888 62688
rect -3089 62615 -3054 62675
rect -2994 62628 -2888 62675
rect -2828 62628 7594 62688
rect -2994 62615 7594 62628
rect -3089 62548 7594 62615
rect -3089 62537 -2883 62548
rect -3089 62487 -3054 62537
rect -3079 62477 -3054 62487
rect -2994 62488 -2883 62537
rect -2823 62488 7594 62548
rect -2994 62487 7594 62488
rect -2994 62477 -2804 62487
rect -3079 62466 -2804 62477
rect -4059 61382 -3685 61414
rect -4059 61374 -2311 61382
rect -4059 61361 -3847 61374
rect -4059 61301 -4013 61361
rect -3953 61314 -3847 61361
rect -3787 61314 -2311 61374
rect -3953 61301 -2311 61314
rect -4059 61234 -2311 61301
rect -4059 61223 -3842 61234
rect -4059 61163 -4013 61223
rect -3953 61174 -3842 61223
rect -3782 61174 -2311 61234
rect -3953 61163 -2311 61174
rect -4059 61157 -2311 61163
rect -4059 61153 -3685 61157
rect -4059 61136 -3689 61153
rect -2118 60500 -1893 60774
rect -2698 52730 -2423 52744
rect -2698 52670 -2673 52730
rect -2613 52728 -2423 52730
rect -2613 52670 -2509 52728
rect -2698 52668 -2509 52670
rect -2449 52668 -2423 52728
rect -2698 52616 -2423 52668
rect -2698 52603 -2507 52616
rect -2698 52543 -2673 52603
rect -2613 52556 -2507 52603
rect -2447 52575 -2423 52616
rect -2447 52556 861 52575
rect -2613 52543 861 52556
rect -2698 52476 861 52543
rect -2698 52465 -2502 52476
rect -2698 52405 -2673 52465
rect -2613 52416 -2502 52465
rect -2442 52416 861 52476
rect -2613 52405 861 52416
rect -2698 52399 861 52405
rect -2698 52394 -2423 52399
rect -3907 52218 -3536 52258
rect -3907 52205 -3695 52218
rect -3907 52145 -3861 52205
rect -3801 52158 -3695 52205
rect -3635 52195 -3536 52218
rect -3635 52158 1088 52195
rect -3801 52145 1088 52158
rect -3907 52078 1088 52145
rect -3907 52067 -3690 52078
rect -3907 52007 -3861 52067
rect -3801 52018 -3690 52067
rect -3630 52018 1088 52078
rect -3801 52007 1088 52018
rect -3907 51994 1088 52007
rect -3907 51980 -3537 51994
rect -2076 51992 -1875 51994
rect -2076 50862 -1875 51119
rect -2388 44204 -2113 44218
rect -2388 44144 -2363 44204
rect -2303 44202 -2113 44204
rect -2303 44144 -2199 44202
rect -2388 44142 -2199 44144
rect -2139 44142 -2113 44202
rect -2388 44090 -2113 44142
rect -2388 44077 -2197 44090
rect -2388 44017 -2363 44077
rect -2303 44030 -2197 44077
rect -2137 44030 -2113 44090
rect -2303 44017 -2113 44030
rect -2388 43950 -2113 44017
rect -2388 43939 -2192 43950
rect -2388 43879 -2363 43939
rect -2303 43890 -2192 43939
rect -2132 43933 -2113 43950
rect 1490 43933 1578 44198
rect -2132 43890 1578 43933
rect -2303 43879 1578 43890
rect -2388 43868 1578 43879
rect -2336 43845 1578 43868
rect -2336 43798 -2269 43845
rect 1490 43798 1578 43845
rect -2381 43663 -2106 43677
rect -2381 43603 -2356 43663
rect -2296 43661 -2106 43663
rect -2296 43603 -2192 43661
rect -2381 43601 -2192 43603
rect -2132 43601 -2106 43661
rect -2381 43549 -2106 43601
rect -2381 43536 -2190 43549
rect -2381 43476 -2356 43536
rect -2296 43489 -2190 43536
rect -2130 43489 -2106 43549
rect -2296 43476 -2106 43489
rect -2381 43409 -2106 43476
rect -2381 43398 -2185 43409
rect -2381 43338 -2356 43398
rect -2296 43349 -2185 43398
rect -2125 43349 -2106 43409
rect -2296 43338 -2106 43349
rect -2381 43327 -2106 43338
rect -2489 36770 -2214 36784
rect -2489 36710 -2464 36770
rect -2404 36768 -2214 36770
rect -2404 36710 -2300 36768
rect -2489 36708 -2300 36710
rect -2240 36708 -2214 36768
rect -2489 36656 -2214 36708
rect -2489 36643 -2298 36656
rect -2489 36583 -2464 36643
rect -2404 36596 -2298 36643
rect -2238 36596 -2214 36656
rect -2404 36583 -2214 36596
rect -2489 36516 -2214 36583
rect -2489 36505 -2293 36516
rect -2489 36445 -2464 36505
rect -2404 36456 -2293 36505
rect -2233 36456 -2214 36516
rect -2404 36445 -2214 36456
rect -2489 36434 -2214 36445
rect 6888 32662 7411 33451
rect -4689 32139 7411 32662
rect -4689 18858 -4166 32139
rect 2010 28029 2740 28118
rect 2010 28021 2605 28029
rect 2010 27961 2039 28021
rect 2099 28018 2415 28021
rect 2099 27961 2218 28018
rect 2010 27958 2218 27961
rect 2278 27961 2415 28018
rect 2475 27969 2605 28021
rect 2665 27969 2740 28029
rect 2475 27961 2740 27969
rect 2278 27958 2740 27961
rect 2010 27894 2740 27958
rect 2010 27834 2042 27894
rect 2102 27886 2605 27894
rect 2102 27883 2407 27886
rect 2102 27834 2218 27883
rect 2010 27823 2218 27834
rect 2278 27826 2407 27883
rect 2467 27834 2605 27886
rect 2665 27834 2740 27894
rect 2467 27826 2740 27834
rect 2278 27823 2740 27826
rect 2010 27720 2740 27823
rect 2011 21918 2709 27720
rect 2011 21782 22718 21918
rect 2011 21762 8972 21782
rect 2011 21696 8757 21762
rect 8829 21716 8972 21762
rect 9044 21716 22718 21782
rect 8829 21696 22718 21716
rect 2011 21609 22718 21696
rect 2011 21599 8908 21609
rect 2011 21533 8646 21599
rect 8718 21543 8908 21599
rect 8980 21543 22718 21609
rect 8718 21533 22718 21543
rect 2011 21358 22718 21533
rect 2011 21348 8884 21358
rect 2011 21282 8664 21348
rect 8736 21292 8884 21348
rect 8956 21292 22718 21358
rect 8736 21282 22718 21292
rect 2011 21220 22718 21282
rect -265 20781 1066 20974
rect -265 20716 20745 20781
rect -265 20696 369 20716
rect -265 20630 154 20696
rect 226 20650 369 20696
rect 441 20650 20745 20716
rect 226 20630 20745 20650
rect -265 20543 20745 20630
rect -265 20533 305 20543
rect -265 20467 43 20533
rect 115 20477 305 20533
rect 377 20477 20745 20543
rect 115 20467 20745 20477
rect -265 20292 20745 20467
rect -265 20282 281 20292
rect -265 20216 61 20282
rect 133 20226 281 20282
rect 353 20226 20745 20292
rect 133 20216 20745 20226
rect -265 20107 20745 20216
rect -265 19888 1066 20107
rect -4689 18335 17883 18858
rect 17360 14316 17883 18335
rect 17360 14185 18261 14316
rect 17360 14165 17787 14185
rect 17360 14099 17572 14165
rect 17644 14119 17787 14165
rect 17859 14119 18261 14185
rect 17644 14117 18261 14119
rect 17644 14099 18048 14117
rect 17360 14051 18048 14099
rect 18120 14051 18261 14117
rect 17360 14012 18261 14051
rect 17360 14002 17723 14012
rect 17360 13936 17461 14002
rect 17533 13946 17723 14002
rect 17795 13950 18261 14012
rect 17795 13946 17912 13950
rect 17533 13936 17912 13946
rect 17360 13884 17912 13936
rect 17984 13884 18261 13950
rect 17360 13761 18261 13884
rect 17360 13751 17699 13761
rect 17360 13685 17479 13751
rect 17551 13695 17699 13751
rect 17771 13700 18261 13761
rect 20071 14109 20745 20107
rect 22020 17766 22718 21220
rect 22020 17741 49711 17766
rect 22020 17109 91956 17741
rect 22020 17094 55075 17109
rect 22020 17068 49711 17094
rect 20071 14099 20472 14109
rect 20071 14033 20252 14099
rect 20324 14043 20472 14099
rect 20544 14043 20745 14109
rect 20324 14033 20745 14043
rect 20071 13910 20745 14033
rect 20071 13844 20243 13910
rect 20315 13904 20745 13910
rect 20315 13844 20470 13904
rect 20071 13838 20470 13844
rect 20542 13838 20745 13904
rect 20071 13708 20745 13838
rect 17771 13695 17916 13700
rect 17551 13685 17916 13695
rect 17360 13634 17916 13685
rect 17988 13634 18261 13700
rect 26035 13671 26139 13672
rect 25430 13657 26202 13671
rect 17360 13556 18261 13634
rect 17360 13490 17697 13556
rect 17769 13490 18261 13556
rect 17360 13289 18261 13490
rect 25426 13642 26202 13657
rect 25426 13538 25496 13642
rect 25600 13538 25684 13642
rect 25788 13538 25879 13642
rect 25983 13538 26202 13642
rect 25426 13428 26202 13538
rect 11365 12714 11683 12801
rect 5394 12710 11683 12714
rect 5394 12650 11397 12710
rect 11457 12707 11683 12710
rect 11457 12650 11581 12707
rect 5394 12647 11581 12650
rect 11641 12647 11683 12707
rect 5394 12582 11683 12647
rect 5394 12522 11394 12582
rect 11454 12574 11683 12582
rect 11454 12522 11579 12574
rect 5394 12514 11579 12522
rect 11639 12514 11683 12574
rect 5394 12473 11683 12514
rect 5394 12470 5595 12473
rect 5394 12390 5422 12470
rect 5502 12393 5595 12470
rect 5675 12437 11683 12473
rect 5675 12393 11395 12437
rect 5502 12390 11395 12393
rect 5394 12377 11395 12390
rect 11455 12377 11572 12437
rect 11632 12377 11683 12437
rect 5394 12363 11683 12377
rect 5394 12279 5745 12363
rect 11365 12334 11683 12363
rect 5394 12199 5421 12279
rect 5501 12277 5745 12279
rect 5501 12199 5582 12277
rect 5394 12197 5582 12199
rect 5662 12197 5745 12277
rect 5394 12132 5745 12197
rect 8578 11669 8996 11732
rect 8578 11666 8871 11669
rect 8578 11665 8725 11666
rect 8578 11605 8605 11665
rect 8665 11606 8725 11665
rect 8785 11609 8871 11666
rect 8931 11609 8996 11669
rect 8785 11606 8996 11609
rect 8665 11605 8996 11606
rect 8578 11554 8996 11605
rect 8578 11494 8610 11554
rect 8670 11494 8741 11554
rect 8801 11494 8881 11554
rect 8941 11494 8996 11554
rect 8578 11488 8996 11494
rect 5268 7568 6063 7709
rect 5268 7564 5727 7568
rect 5268 7548 5588 7564
rect 5268 7488 5391 7548
rect 5451 7504 5588 7548
rect 5648 7508 5727 7564
rect 5787 7564 6063 7568
rect 5787 7508 5871 7564
rect 5648 7504 5871 7508
rect 5931 7504 6063 7564
rect 5451 7488 6063 7504
rect 5268 7444 6063 7488
rect 5268 7430 5850 7444
rect 5268 7423 5676 7430
rect 5268 7418 5503 7423
rect 5268 7358 5354 7418
rect 5414 7363 5503 7418
rect 5563 7370 5676 7423
rect 5736 7384 5850 7430
rect 5910 7384 6063 7444
rect 5736 7370 6063 7384
rect 5563 7363 6063 7370
rect 5414 7358 6063 7363
rect 5268 7315 6063 7358
rect 5268 7310 5939 7315
rect 5268 7306 5637 7310
rect 5268 7298 5474 7306
rect 5268 7238 5323 7298
rect 5383 7246 5474 7298
rect 5534 7250 5637 7306
rect 5697 7250 5798 7310
rect 5858 7255 5939 7310
rect 5999 7255 6063 7315
rect 5858 7250 6063 7255
rect 5534 7246 6063 7250
rect 5383 7238 6063 7246
rect 5268 7226 6063 7238
rect 8648 7137 8897 11488
rect 19634 11244 19861 11247
rect 19622 11199 20513 11244
rect 19622 11197 20146 11199
rect 19622 11192 19907 11197
rect 19622 11132 19666 11192
rect 19726 11137 19907 11192
rect 19967 11139 20146 11197
rect 20206 11139 20373 11199
rect 20433 11139 20513 11199
rect 19967 11137 20513 11139
rect 19726 11132 20513 11137
rect 19622 11090 20513 11132
rect 19634 9198 19861 11090
rect 20286 9198 20513 11090
rect 19580 9187 19979 9198
rect 20206 9187 20513 9198
rect 19580 9153 20513 9187
rect 19580 9151 20104 9153
rect 19580 9146 19865 9151
rect 19580 9086 19624 9146
rect 19684 9091 19865 9146
rect 19925 9093 20104 9151
rect 20164 9093 20331 9153
rect 20391 9093 20513 9153
rect 19925 9091 20513 9093
rect 19684 9086 20513 9091
rect 19580 9044 20513 9086
rect 20286 8003 20513 9044
rect 25973 9080 26202 13428
rect 28727 10002 32041 10065
rect 28718 9904 32041 10002
rect 28718 9902 29260 9904
rect 28718 9897 29021 9902
rect 28718 9837 28780 9897
rect 28840 9842 29021 9897
rect 29081 9844 29260 9902
rect 29320 9844 29487 9904
rect 29547 9844 32041 9904
rect 29081 9842 32041 9844
rect 28840 9837 32041 9842
rect 28718 9814 32041 9837
rect 28718 9777 29681 9814
rect 30509 9080 30918 9085
rect 25973 9034 30918 9080
rect 25973 9021 30665 9034
rect 25973 8961 30533 9021
rect 30593 8974 30665 9021
rect 30725 9033 30918 9034
rect 30725 8974 30790 9033
rect 30593 8973 30790 8974
rect 30850 8973 30918 9033
rect 30593 8961 30918 8973
rect 25973 8924 30918 8961
rect 25973 8908 30663 8924
rect 25973 8851 30530 8908
rect 30355 8848 30530 8851
rect 30590 8864 30663 8908
rect 30723 8864 30790 8924
rect 30850 8864 30918 8924
rect 30590 8848 30918 8864
rect 30355 8797 30918 8848
rect 30355 8795 30652 8797
rect 30355 8735 30527 8795
rect 30587 8737 30652 8795
rect 30712 8737 30790 8797
rect 30850 8737 30918 8797
rect 30587 8735 30918 8737
rect 30355 8672 30918 8735
rect 20286 7955 20641 8003
rect 20286 7885 26699 7955
rect 20286 7883 23415 7885
rect 20286 7878 23176 7883
rect 20286 7818 22935 7878
rect 22995 7823 23176 7878
rect 23236 7825 23415 7883
rect 23475 7825 23642 7885
rect 23702 7825 26699 7885
rect 23236 7823 26699 7825
rect 22995 7818 26699 7823
rect 20286 7728 26699 7818
rect 8560 7077 9108 7137
rect 8560 7070 8949 7077
rect 8560 7010 8588 7070
rect 8648 7010 8729 7070
rect 8789 7017 8949 7070
rect 9009 7017 9108 7077
rect 8789 7010 9108 7017
rect 8560 6960 9108 7010
rect 8560 6900 8594 6960
rect 8654 6955 9108 6960
rect 8654 6900 8735 6955
rect 8560 6895 8735 6900
rect 8795 6895 8975 6955
rect 9035 6895 9108 6955
rect 8560 6879 9108 6895
rect 20318 352 20641 7728
rect 26472 6980 26699 7728
rect 31790 6980 32041 9814
rect 49039 9313 49671 17068
rect 53921 9320 54794 9377
rect 53921 9319 54370 9320
rect 53921 9316 54246 9319
rect 53921 9313 54010 9316
rect 49039 9256 54010 9313
rect 54070 9256 54129 9316
rect 54189 9259 54246 9316
rect 54306 9260 54370 9319
rect 54430 9319 54794 9320
rect 54430 9260 54487 9319
rect 54306 9259 54487 9260
rect 54547 9313 54794 9319
rect 61491 9327 62361 9385
rect 61491 9326 61940 9327
rect 61491 9323 61816 9326
rect 61491 9313 61580 9323
rect 54547 9263 61580 9313
rect 61640 9263 61699 9323
rect 61759 9266 61816 9323
rect 61876 9267 61940 9326
rect 62000 9326 62361 9327
rect 62000 9267 62057 9326
rect 61876 9266 62057 9267
rect 62117 9313 62361 9326
rect 62117 9266 62375 9313
rect 61759 9263 62375 9266
rect 54547 9259 62375 9263
rect 54189 9256 62375 9259
rect 49039 9213 62375 9256
rect 49039 9209 61941 9213
rect 49039 9207 61821 9209
rect 49039 9206 61580 9207
rect 49039 9202 54371 9206
rect 49039 9200 54251 9202
rect 49039 9140 54010 9200
rect 54070 9140 54128 9200
rect 54188 9142 54251 9200
rect 54311 9146 54371 9202
rect 54431 9199 61580 9206
rect 54431 9146 54489 9199
rect 54311 9142 54489 9146
rect 54188 9140 54489 9142
rect 49039 9139 54489 9140
rect 54549 9147 61580 9199
rect 61640 9147 61698 9207
rect 61758 9149 61821 9207
rect 61881 9153 61941 9209
rect 62001 9206 62375 9213
rect 62001 9153 62059 9206
rect 61881 9149 62059 9153
rect 61758 9147 62059 9149
rect 54549 9146 62059 9147
rect 62119 9146 62375 9206
rect 54549 9139 62375 9146
rect 49039 9087 62375 9139
rect 26472 6910 32041 6980
rect 26472 6908 29204 6910
rect 26472 6903 28965 6908
rect 26472 6843 28724 6903
rect 28784 6848 28965 6903
rect 29025 6850 29204 6908
rect 29264 6850 29431 6910
rect 29491 6850 32041 6910
rect 29025 6848 32041 6850
rect 28784 6843 32041 6848
rect 26472 6753 32041 6843
rect 27167 4463 27415 6753
rect 31790 6741 32041 6753
rect 32327 7125 32533 7128
rect 32327 7124 43272 7125
rect 44110 7124 44460 7130
rect 32327 7111 44715 7124
rect 32327 6941 43278 7111
rect 43448 6941 43821 7111
rect 43991 6941 44531 7111
rect 44701 6941 44715 7111
rect 46136 7091 47059 7119
rect 46136 7086 46925 7091
rect 46136 7008 46183 7086
rect 46259 7083 46925 7086
rect 46259 7081 46709 7083
rect 46259 7008 46429 7081
rect 46136 7003 46429 7008
rect 46505 7005 46709 7081
rect 46785 7013 46925 7083
rect 47001 7013 47059 7091
rect 46785 7005 47059 7013
rect 46505 7003 47059 7005
rect 46136 6961 47059 7003
rect 32327 6919 44715 6941
rect 30400 5978 30606 5983
rect 32327 5978 32533 6919
rect 38287 6633 38493 6919
rect 44110 6850 44480 6919
rect 44110 6810 44460 6850
rect 38287 6414 38493 6427
rect 46593 6163 46752 6961
rect 47454 6163 47743 6195
rect 46512 6130 47745 6163
rect 30400 5772 32533 5978
rect 43759 6087 47745 6130
rect 43759 6009 43813 6087
rect 43889 6074 47745 6087
rect 43889 6009 44062 6074
rect 43759 5996 44062 6009
rect 44138 6073 47745 6074
rect 44138 6069 44518 6073
rect 44138 5996 44296 6069
rect 43759 5991 44296 5996
rect 44372 5995 44518 6069
rect 44594 5995 47745 6073
rect 44372 5991 47745 5995
rect 43759 5971 47745 5991
rect 46512 5937 47745 5971
rect 30400 4524 30606 5772
rect 27094 4444 27485 4463
rect 27094 4314 27110 4444
rect 27240 4314 27342 4444
rect 27472 4314 27485 4444
rect 27094 4248 27485 4314
rect 27094 4118 27107 4248
rect 27237 4118 27342 4248
rect 27472 4118 27485 4248
rect 30400 4399 30434 4524
rect 30559 4399 30606 4524
rect 30400 4263 30606 4399
rect 30400 4138 30434 4263
rect 30559 4138 30606 4263
rect 30400 4129 30606 4138
rect 27094 4108 27485 4118
rect 47454 3849 47743 5937
rect 49039 4545 49671 9087
rect 91324 4952 91956 17109
rect 91324 4724 99215 4952
rect 53695 4666 54568 4724
rect 53695 4665 54144 4666
rect 53695 4662 54020 4665
rect 53695 4602 53784 4662
rect 53844 4602 53903 4662
rect 53963 4605 54020 4662
rect 54080 4606 54144 4665
rect 54204 4665 54568 4666
rect 54204 4606 54261 4665
rect 54080 4605 54261 4606
rect 54321 4605 54568 4665
rect 53963 4602 54568 4605
rect 53695 4552 54568 4602
rect 53695 4548 54145 4552
rect 53695 4546 54025 4548
rect 53695 4545 53784 4546
rect 49039 4486 53784 4545
rect 53844 4486 53902 4546
rect 53962 4488 54025 4546
rect 54085 4492 54145 4548
rect 54205 4545 54568 4552
rect 91324 4666 98886 4724
rect 98948 4718 99215 4724
rect 98948 4666 99061 4718
rect 91324 4660 99061 4666
rect 99123 4660 99215 4718
rect 91324 4569 99215 4660
rect 91324 4565 99062 4569
rect 54205 4492 54263 4545
rect 54085 4488 54263 4492
rect 53962 4486 54263 4488
rect 49039 4485 54263 4486
rect 54323 4485 57420 4545
rect 49039 4319 57420 4485
rect 49039 4304 49671 4319
rect 49161 4303 49588 4304
rect 49161 3849 49588 3854
rect 47454 3560 49588 3849
rect 17589 29 20641 352
rect 4778 -986 5148 -932
rect 4778 -1046 4824 -986
rect 4884 -988 5148 -986
rect 4884 -1046 4988 -988
rect 4778 -1048 4988 -1046
rect 5048 -1004 5148 -988
rect 5048 -1048 15958 -1004
rect 4778 -1100 15958 -1048
rect 4778 -1113 4990 -1100
rect 4778 -1173 4824 -1113
rect 4884 -1160 4990 -1113
rect 5050 -1160 15958 -1100
rect 4884 -1173 15958 -1160
rect 4778 -1240 15958 -1173
rect 4778 -1251 4995 -1240
rect 4778 -1311 4824 -1251
rect 4884 -1300 4995 -1251
rect 5055 -1300 15958 -1240
rect 4884 -1311 15958 -1300
rect 4778 -1321 15958 -1311
rect 4778 -1338 5148 -1321
rect 4844 -1552 14921 -1512
rect 4844 -1565 5056 -1552
rect 4844 -1625 4890 -1565
rect 4950 -1612 5056 -1565
rect 5116 -1612 14921 -1552
rect 4950 -1625 14921 -1612
rect 4844 -1692 14921 -1625
rect 4844 -1703 5061 -1692
rect 4844 -1763 4890 -1703
rect 4950 -1752 5061 -1703
rect 5121 -1752 14921 -1692
rect 4950 -1756 14921 -1752
rect 4950 -1763 5222 -1756
rect 4844 -1773 5222 -1763
rect 4844 -1790 5214 -1773
rect 14677 -2260 14921 -1756
rect 15641 -1813 15958 -1321
rect 17649 -1459 17851 29
rect 18284 -745 21310 -725
rect 18284 -858 18296 -745
rect 18423 -858 21310 -745
rect 18284 -887 21310 -858
rect 18284 -906 18760 -887
rect 18284 -1019 18501 -906
rect 18628 -1000 18760 -906
rect 18887 -1000 21310 -887
rect 18628 -1019 21310 -1000
rect 18284 -1061 21310 -1019
rect 20974 -1269 21310 -1061
rect 17649 -1502 18861 -1459
rect 17649 -1515 18671 -1502
rect 17649 -1628 18108 -1515
rect 18235 -1628 18417 -1515
rect 18544 -1615 18671 -1515
rect 18798 -1615 18861 -1502
rect 20974 -1605 26713 -1269
rect 18544 -1628 18861 -1615
rect 17649 -1661 18861 -1628
rect 15641 -2130 25855 -1813
rect 24985 -2260 25196 -2248
rect 14677 -2504 25212 -2260
rect 5001 -2623 5379 -2608
rect 4971 -2648 24848 -2623
rect 4971 -2661 5213 -2648
rect 4971 -2721 5047 -2661
rect 5107 -2708 5213 -2661
rect 5273 -2708 24848 -2648
rect 5107 -2721 24848 -2708
rect 4971 -2774 24848 -2721
rect 5001 -2788 5379 -2774
rect 5001 -2799 5218 -2788
rect 5001 -2859 5047 -2799
rect 5107 -2848 5218 -2799
rect 5278 -2848 5379 -2788
rect 5107 -2859 5379 -2848
rect 5001 -2869 5379 -2859
rect 5001 -2886 5371 -2869
rect 4975 -3026 16639 -2983
rect 4905 -3066 16639 -3026
rect 4905 -3079 5117 -3066
rect 4905 -3139 4951 -3079
rect 5011 -3126 5117 -3079
rect 5177 -3126 16639 -3066
rect 5011 -3139 16639 -3126
rect 4905 -3206 16639 -3139
rect 4905 -3217 5122 -3206
rect 4905 -3277 4951 -3217
rect 5011 -3266 5122 -3217
rect 5182 -3232 16639 -3206
rect 5182 -3266 5283 -3232
rect 5011 -3277 5283 -3266
rect 4905 -3287 5283 -3277
rect 4905 -3304 5275 -3287
rect 4882 -3462 5260 -3440
rect 4882 -3480 16212 -3462
rect 4882 -3493 5094 -3480
rect 4882 -3553 4928 -3493
rect 4988 -3540 5094 -3493
rect 5154 -3540 16212 -3480
rect 4988 -3553 16212 -3540
rect 4882 -3620 16212 -3553
rect 4882 -3631 5099 -3620
rect 4882 -3691 4928 -3631
rect 4988 -3680 5099 -3631
rect 5159 -3643 16212 -3620
rect 5159 -3680 5260 -3643
rect 4988 -3691 5260 -3680
rect 4882 -3701 5260 -3691
rect 4882 -3718 5252 -3701
rect 5001 -3919 7452 -3878
rect 4928 -3959 7452 -3919
rect 4928 -3972 5140 -3959
rect 4928 -4032 4974 -3972
rect 5034 -4019 5140 -3972
rect 5200 -4019 7452 -3959
rect 5034 -4032 7452 -4019
rect 4928 -4099 7452 -4032
rect 4928 -4110 5145 -4099
rect 4928 -4170 4974 -4110
rect 5034 -4159 5145 -4110
rect 5205 -4103 7452 -4099
rect 5205 -4159 5306 -4103
rect 5034 -4170 5306 -4159
rect 4928 -4180 5306 -4170
rect 4928 -4197 5298 -4180
rect 7227 -4372 7452 -4103
rect 5070 -4462 6102 -4418
rect 5033 -4502 6102 -4462
rect 5033 -4515 5245 -4502
rect 5033 -4575 5079 -4515
rect 5139 -4562 5245 -4515
rect 5305 -4562 6102 -4502
rect 5139 -4575 6102 -4562
rect 5033 -4630 6102 -4575
rect 5033 -4642 5411 -4630
rect 5033 -4653 5250 -4642
rect 5033 -4713 5079 -4653
rect 5139 -4702 5250 -4653
rect 5310 -4702 5411 -4642
rect 5139 -4713 5411 -4702
rect 5033 -4723 5411 -4713
rect 5033 -4740 5403 -4723
rect 16031 -5048 16212 -3643
rect 16390 -5174 16639 -3232
rect 24697 -5269 24848 -2774
rect 24985 -5303 25196 -2504
rect 25538 -3786 25855 -2130
rect 26377 -2241 26713 -1605
rect 49161 -1981 49588 3560
rect 57127 213 57420 4319
rect 91324 4507 98884 4565
rect 98946 4511 99062 4565
rect 99124 4511 99215 4569
rect 98946 4507 99215 4511
rect 91324 4400 99215 4507
rect 91324 4342 98887 4400
rect 98949 4395 99215 4400
rect 98949 4342 99075 4395
rect 91324 4337 99075 4342
rect 99137 4337 99215 4395
rect 91324 4320 99215 4337
rect 91324 4259 92059 4320
rect 98838 4305 99160 4320
rect 91324 4258 91776 4259
rect 91324 4255 91652 4258
rect 91324 4195 91416 4255
rect 91476 4195 91535 4255
rect 91595 4198 91652 4255
rect 91712 4199 91776 4258
rect 91836 4258 92059 4259
rect 91836 4199 91893 4258
rect 91712 4198 91893 4199
rect 91953 4198 92059 4258
rect 91595 4195 92059 4198
rect 91324 4145 92059 4195
rect 91324 4141 91777 4145
rect 91324 4139 91657 4141
rect 91324 4079 91416 4139
rect 91476 4079 91534 4139
rect 91594 4081 91657 4139
rect 91717 4085 91777 4141
rect 91837 4138 92059 4145
rect 91837 4085 91895 4138
rect 91717 4081 91895 4085
rect 91594 4079 91895 4081
rect 91324 4078 91895 4079
rect 91955 4078 92059 4138
rect 91324 4051 92059 4078
rect 91324 4026 91956 4051
rect 55465 -151 57420 213
rect 26377 -2577 36376 -2241
rect 49161 -2408 51945 -1981
rect 25538 -4103 32240 -3786
rect 31923 -5255 32240 -4103
rect 36040 -6541 36376 -2577
rect 51518 -4201 51945 -2408
rect 51284 -4233 52067 -4201
rect 51284 -4260 51573 -4233
rect 51284 -4341 51332 -4260
rect 51413 -4314 51573 -4260
rect 51654 -4264 52067 -4233
rect 51654 -4314 51848 -4264
rect 51413 -4341 51848 -4314
rect 51284 -4345 51848 -4341
rect 51929 -4345 52067 -4264
rect 51284 -4383 52067 -4345
rect 51284 -4402 51559 -4383
rect 51284 -4483 51316 -4402
rect 51397 -4464 51559 -4402
rect 51640 -4414 52067 -4383
rect 51640 -4464 51821 -4414
rect 51397 -4483 51821 -4464
rect 51284 -4495 51821 -4483
rect 51902 -4495 52067 -4414
rect 51284 -4560 52067 -4495
rect 51284 -4564 51547 -4560
rect 51284 -4645 51301 -4564
rect 51382 -4641 51547 -4564
rect 51628 -4564 52067 -4560
rect 51628 -4641 51855 -4564
rect 51382 -4645 51855 -4641
rect 51936 -4645 52067 -4564
rect 51284 -4719 52067 -4645
rect 36093 -14454 36324 -6662
rect 52279 -11322 53565 -11166
rect 52279 -11364 53571 -11322
rect 52279 -11367 53315 -11364
rect 52279 -11375 53073 -11367
rect 52279 -11377 52804 -11375
rect 52279 -11390 52549 -11377
rect 52279 -11450 52344 -11390
rect 52404 -11437 52549 -11390
rect 52609 -11435 52804 -11377
rect 52864 -11427 53073 -11375
rect 53133 -11424 53315 -11367
rect 53375 -11424 53571 -11364
rect 53133 -11427 53571 -11424
rect 52864 -11435 53571 -11427
rect 52609 -11437 53571 -11435
rect 52404 -11450 53571 -11437
rect 52279 -11479 53571 -11450
rect 55465 -11479 55829 -151
rect 98561 -757 98873 -742
rect 56983 -815 98599 -757
rect 98661 -763 98873 -757
rect 98661 -815 98774 -763
rect 56983 -821 98774 -815
rect 98836 -821 98873 -763
rect 56983 -912 98873 -821
rect 56983 -916 98775 -912
rect 56983 -974 98597 -916
rect 98659 -970 98775 -916
rect 98837 -970 98873 -912
rect 98659 -974 98873 -970
rect 56983 -1081 98873 -974
rect 56983 -1139 98600 -1081
rect 98662 -1086 98873 -1081
rect 98662 -1139 98788 -1086
rect 56983 -1144 98788 -1139
rect 98850 -1144 98873 -1086
rect 56983 -1181 98873 -1144
rect 56983 -1186 98866 -1181
rect 56983 -5243 57309 -1186
rect 67147 -1961 98964 -1936
rect 67147 -2019 98632 -1961
rect 98694 -1962 98964 -1961
rect 98694 -2019 98806 -1962
rect 67147 -2020 98806 -2019
rect 98868 -2020 98964 -1962
rect 67147 -2127 98964 -2020
rect 67147 -2185 98633 -2127
rect 98695 -2132 98964 -2127
rect 98695 -2185 98831 -2132
rect 67147 -2190 98831 -2185
rect 98893 -2190 98964 -2132
rect 67147 -2230 98964 -2190
rect 58351 -2964 58627 -2793
rect 58344 -3008 58627 -2964
rect 58344 -3033 58523 -3008
rect 58344 -3095 58353 -3033
rect 58411 -3070 58523 -3033
rect 58581 -3070 58627 -3008
rect 58411 -3095 58627 -3070
rect 58344 -3206 58627 -3095
rect 58344 -3207 58518 -3206
rect 58344 -3269 58352 -3207
rect 58410 -3268 58518 -3207
rect 58576 -3268 58627 -3206
rect 58410 -3269 58627 -3268
rect 58344 -3325 58627 -3269
rect 58351 -3328 58627 -3325
rect 58377 -5154 58602 -3328
rect 67147 -4968 67396 -2230
rect 98546 -2858 98907 -2850
rect 98546 -2905 98602 -2858
rect 75818 -2916 98602 -2905
rect 98664 -2859 98907 -2858
rect 98664 -2916 98776 -2859
rect 75818 -2917 98776 -2916
rect 98838 -2917 98907 -2859
rect 75818 -3024 98907 -2917
rect 75818 -3082 98603 -3024
rect 98665 -3029 98907 -3024
rect 98665 -3082 98801 -3029
rect 75818 -3087 98801 -3082
rect 98863 -3087 98907 -3029
rect 75818 -3114 98907 -3087
rect 68159 -3635 68520 -3628
rect 68156 -3636 68691 -3635
rect 68156 -3661 68215 -3636
rect 68107 -3683 68215 -3661
rect 67579 -3694 68215 -3683
rect 68277 -3637 68691 -3636
rect 68277 -3694 68389 -3637
rect 67579 -3695 68389 -3694
rect 68451 -3695 68691 -3637
rect 67579 -3802 68691 -3695
rect 67579 -3854 68216 -3802
rect 67579 -5030 67750 -3854
rect 68107 -3860 68216 -3854
rect 68278 -3807 68691 -3802
rect 68278 -3860 68414 -3807
rect 68107 -3865 68414 -3860
rect 68476 -3865 68691 -3807
rect 68107 -3886 68691 -3865
rect 68156 -3911 68691 -3886
rect 57040 -5346 57252 -5243
rect 68640 -5267 69133 -5096
rect 75848 -5104 75996 -3114
rect 98546 -3118 98907 -3114
rect 76086 -3341 98994 -3305
rect 76086 -3399 98594 -3341
rect 98656 -3342 98994 -3341
rect 98656 -3399 98768 -3342
rect 76086 -3400 98768 -3399
rect 98830 -3400 98994 -3342
rect 76086 -3507 98994 -3400
rect 76086 -3565 98595 -3507
rect 98657 -3512 98994 -3507
rect 98657 -3565 98793 -3512
rect 76086 -3570 98793 -3565
rect 98855 -3570 98994 -3512
rect 76086 -3614 98994 -3570
rect 75883 -5179 75961 -5104
rect 76158 -5181 76323 -3614
rect 98576 -3892 98937 -3885
rect 83093 -3893 99108 -3892
rect 83093 -3951 98632 -3893
rect 98694 -3894 99108 -3893
rect 98694 -3951 98806 -3894
rect 83093 -3952 98806 -3951
rect 98868 -3952 99108 -3894
rect 83093 -4059 99108 -3952
rect 83093 -4117 98633 -4059
rect 98695 -4064 99108 -4059
rect 98695 -4117 98831 -4064
rect 83093 -4122 98831 -4117
rect 98893 -4122 99108 -4064
rect 83093 -4168 99108 -4122
rect 83093 -5156 83369 -4168
rect 87090 -4720 87760 -4550
rect 87090 -4780 87130 -4720
rect 87190 -4780 87250 -4720
rect 87310 -4780 87370 -4720
rect 87430 -4780 87760 -4720
rect 87090 -4840 87760 -4780
rect 87090 -4900 87130 -4840
rect 87190 -4900 87250 -4840
rect 87310 -4900 87370 -4840
rect 87430 -4900 87760 -4840
rect 87090 -4960 87760 -4900
rect 87090 -5020 87132 -4960
rect 87192 -5020 87250 -4960
rect 87310 -5020 87370 -4960
rect 87430 -5020 87760 -4960
rect 87090 -5090 87760 -5020
rect 52279 -11546 55829 -11479
rect 52279 -11547 53402 -11546
rect 52279 -11559 53243 -11547
rect 52279 -11562 53030 -11559
rect 52279 -11572 52785 -11562
rect 52279 -11580 52552 -11572
rect 52279 -11640 52346 -11580
rect 52406 -11632 52552 -11580
rect 52612 -11622 52785 -11572
rect 52845 -11619 53030 -11562
rect 53090 -11607 53243 -11559
rect 53303 -11606 53402 -11547
rect 53462 -11606 55829 -11546
rect 53303 -11607 55829 -11606
rect 53090 -11619 55829 -11607
rect 52845 -11622 55829 -11619
rect 52612 -11632 55829 -11622
rect 52406 -11640 55829 -11632
rect 52279 -11732 55829 -11640
rect 52279 -11740 53351 -11732
rect 52279 -11750 53153 -11740
rect 52279 -11753 52914 -11750
rect 52279 -11755 52703 -11753
rect 52279 -11756 52505 -11755
rect 52279 -11816 52337 -11756
rect 52397 -11815 52505 -11756
rect 52565 -11813 52703 -11755
rect 52763 -11810 52914 -11753
rect 52974 -11800 53153 -11750
rect 53213 -11792 53351 -11740
rect 53411 -11792 55829 -11732
rect 53213 -11800 55829 -11792
rect 52974 -11810 55829 -11800
rect 52763 -11813 55829 -11810
rect 52565 -11815 55829 -11813
rect 52397 -11816 55829 -11815
rect 52279 -11843 55829 -11816
rect 52279 -11848 53571 -11843
rect 87243 -14434 87474 -5992
rect 34855 -14685 36324 -14454
rect 78405 -14665 87474 -14434
<< via3 >>
rect 5422 12390 5502 12470
rect 5595 12393 5675 12473
rect 5421 12199 5501 12279
rect 5582 12197 5662 12277
rect 5391 7488 5451 7548
rect 5588 7504 5648 7564
rect 5727 7508 5787 7568
rect 5871 7504 5931 7564
rect 5354 7358 5414 7418
rect 5503 7363 5563 7423
rect 5676 7370 5736 7430
rect 5850 7384 5910 7444
rect 5323 7238 5383 7298
rect 5474 7246 5534 7306
rect 5637 7250 5697 7310
rect 5798 7250 5858 7310
rect 5939 7255 5999 7315
rect 51332 -4341 51413 -4260
rect 51573 -4314 51654 -4233
rect 51848 -4345 51929 -4264
rect 51316 -4483 51397 -4402
rect 51559 -4464 51640 -4383
rect 51821 -4495 51902 -4414
rect 51301 -4645 51382 -4564
rect 51547 -4641 51628 -4560
rect 51855 -4645 51936 -4564
<< metal4 >>
rect -7940 41508 -7091 41515
rect -7940 41159 -2689 41508
rect -7940 40575 -2522 41159
rect -7940 -27439 -7091 40575
rect 5385 12473 5993 29177
rect 27663 28397 28023 28607
rect 27811 28389 28023 28397
rect 5385 12470 5595 12473
rect 5385 12390 5422 12470
rect 5502 12393 5595 12470
rect 5675 12393 5993 12473
rect 5502 12390 5993 12393
rect 5385 12279 5993 12390
rect 5385 12199 5421 12279
rect 5501 12277 5993 12279
rect 5501 12199 5582 12277
rect 5385 12197 5582 12199
rect 5662 12197 5993 12277
rect 5385 7709 5993 12197
rect 5268 7568 6063 7709
rect 5268 7564 5727 7568
rect 5268 7548 5588 7564
rect 5268 7488 5391 7548
rect 5451 7504 5588 7548
rect 5648 7508 5727 7564
rect 5787 7564 6063 7568
rect 5787 7508 5871 7564
rect 5648 7504 5871 7508
rect 5931 7504 6063 7564
rect 5451 7488 6063 7504
rect 5268 7444 6063 7488
rect 5268 7430 5850 7444
rect 5268 7423 5676 7430
rect 5268 7418 5503 7423
rect 5268 7358 5354 7418
rect 5414 7363 5503 7418
rect 5563 7370 5676 7423
rect 5736 7384 5850 7430
rect 5910 7384 6063 7444
rect 5736 7370 6063 7384
rect 5563 7363 6063 7370
rect 5414 7358 6063 7363
rect 5268 7315 6063 7358
rect 5268 7310 5939 7315
rect 5268 7306 5637 7310
rect 5268 7298 5474 7306
rect 5268 7238 5323 7298
rect 5383 7246 5474 7298
rect 5534 7250 5637 7306
rect 5697 7250 5798 7310
rect 5858 7255 5939 7310
rect 5999 7255 6063 7315
rect 5858 7250 6063 7255
rect 5534 7246 6063 7250
rect 5383 7238 6063 7246
rect 5268 7226 6063 7238
rect 5385 -5287 5993 7226
rect 51271 -4204 52095 -4173
rect 27683 -4233 64047 -4204
rect 27683 -4260 51573 -4233
rect 27683 -4341 51332 -4260
rect 51413 -4314 51573 -4260
rect 51654 -4264 64047 -4233
rect 51654 -4314 51848 -4264
rect 51413 -4341 51848 -4314
rect 27683 -4345 51848 -4341
rect 51929 -4345 64047 -4264
rect 27683 -4383 64047 -4345
rect 27683 -4402 51559 -4383
rect 27683 -4483 51316 -4402
rect 51397 -4464 51559 -4402
rect 51640 -4414 64047 -4383
rect 51640 -4464 51821 -4414
rect 51397 -4483 51821 -4464
rect 27683 -4495 51821 -4483
rect 51902 -4495 64047 -4414
rect 27683 -4560 64047 -4495
rect 27683 -4564 51547 -4560
rect 27683 -4645 51301 -4564
rect 51382 -4641 51547 -4564
rect 51628 -4564 64047 -4560
rect 51628 -4641 51855 -4564
rect 51382 -4645 51855 -4641
rect 51936 -4645 64047 -4564
rect 27683 -4719 64047 -4645
rect 5385 -5895 8343 -5287
rect 39445 -6852 59430 -6272
rect 11279 -27389 12128 -26499
rect 21483 -27389 22332 -26499
rect 11279 -27439 22332 -27389
rect -7940 -27686 22332 -27439
rect 28864 -27686 29713 -26251
rect 62449 -27498 66334 -26649
rect 62449 -27686 63298 -27498
rect -7940 -28288 63298 -27686
rect 21483 -28535 63298 -28288
rect 65485 -27544 66334 -27498
rect 72203 -27544 73052 -26649
rect 65485 -27594 73052 -27544
rect 80015 -27594 80864 -26550
rect 65485 -28393 80864 -27594
rect 72203 -28443 80864 -28393
<< metal5 >>
rect 27811 28210 28023 28746
rect 95916 21264 96692 22542
rect 95916 20488 98134 21264
rect 97352 20450 98134 20488
rect 97352 118 98128 20450
rect 87362 -658 98128 118
use 7b_divider_magic  7b_divider_magic_0 ~/GF180Projects/Layout/Magic/VCO1/divider
timestamp 1697518002
transform 1 0 57381 0 1 -16876
box -441 -10214 40218 12749
use 7b_divider_magic  7b_divider_magic_1
timestamp 1697518002
transform 0 -1 9619 -1 0 62378
box -441 -10214 40218 12749
use 7b_divider_magic  7b_divider_magic_2
timestamp 1697518002
transform 1 0 6231 0 1 -16896
box -441 -10214 40218 12749
use A_MUX  A_MUX_0 ~/GF180Projects/Layout/Magic/VCO1/A_MUx
timestamp 1697518002
transform 1 0 42495 0 1 4782
box -285 -452 3979 2227
use A_MUX  A_MUX_1
timestamp 1697518002
transform 1 0 18282 0 -1 12510
box -285 -452 3979 2227
use A_MUX  A_MUX_2
timestamp 1697518002
transform 1 0 18240 0 1 7818
box -285 -452 3979 2227
use A_MUX  A_MUX_3
timestamp 1697518002
transform -1 0 30924 0 -1 11425
box -285 -452 3979 2227
use A_MUX  A_MUX_4
timestamp 1697518002
transform -1 0 30867 0 -1 8419
box -285 -452 3979 2227
use A_MUX  A_MUX_5
timestamp 1697518002
transform 1 0 16712 0 1 -3124
box -285 -452 3979 2227
use A_MUX  A_MUX_6
timestamp 1697518002
transform 1 0 36417 0 -1 12138
box -285 -452 3979 2227
use cap_11p  cap_11p_0 ~/GF180Projects/Layout/Magic/ATIF/CP
timestamp 1697518002
transform 1 0 94240 0 1 13088
box -26450 -13708 -6739 632
use cap_240p  cap_240p_0 ~/GF180Projects/Layout/Magic/ATIF/CP
timestamp 1697518021
transform 1 0 89483 0 -1 28277
box -68140 -68970 6839 8429
use CP_1  CP_1_0 ~/GF180Projects/Layout/Magic/ATIF/CP
timestamp 1697518002
transform 1 0 33105 0 1 10459
box -1133 -1188 2101 1774
use Current_Mirror_Top  Current_Mirror_Top_0 ~/GF180Projects/Layout/Magic/VCO1/Current_mirror_Top
timestamp 1697518002
transform -1 0 2228 0 1 10249
box -1992 -209 4486 7070
use INV_2  INV_2_0 ~/GF180Projects/Layout/Magic/VCO1/INV_2
timestamp 1697518002
transform 1 0 11673 0 1 7901
box 21 -485 1081 648
use INV_2  INV_2_1
timestamp 1697518002
transform 1 0 11228 0 1 13239
box 21 -485 1081 648
use PFD_T2  PFD_T2_0 ~/GF180Projects/Layout/Magic/ATIF/PFD_2
timestamp 1697518002
transform 1 0 22661 0 1 8437
box -28 -113 4062 3793
use RES_74k  RES_74k_1 ~/GF180Projects/Layout/Magic/ATIF/Res/RES_p
timestamp 1697518002
transform -1 0 51462 0 -1 12102
box 3672 -1094 9598 4966
use Tappered_Buffer  Tappered_Buffer_0 ~/GF180Projects/Layout/Magic/VCO1/Tappered_Buffer
timestamp 1697518002
transform 1 0 50570 0 1 3553
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_1
timestamp 1697518002
transform 1 0 50390 0 1 8230
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_2
timestamp 1697518002
transform 1 0 58351 0 1 8237
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_4
timestamp 1697518002
transform -1 0 94996 0 1 3197
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_5
timestamp 1697518002
transform 1 0 48878 0 -1 -10328
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_6
timestamp 1697518002
transform -1 0 4941 0 1 26954
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_7
timestamp 1697518002
transform -1 0 11108 0 1 10738
box -161 -3147 5956 876
use Tappered_Buffer  Tappered_Buffer_8
timestamp 1697518002
transform -1 0 12287 0 1 6101
box -161 -3147 5956 876
use VCO_DFF_C  VCO_DFF_C_0 ~/GF180Projects/Layout/Magic/VCO1/VCO_DFF_C
timestamp 1697518002
transform 1 0 24282 0 1 -1600
box 0 -27 23932 7170
<< labels >>
flabel metal1 22036 6756 22036 6756 0 FreeSans 1600 0 0 0 S3
port 19 nsew
flabel metal1 21995 13993 21995 13993 0 FreeSans 1600 0 0 0 UP_INPUT
port 25 nsew
flabel metal1 18022 14399 18022 14399 0 FreeSans 1600 0 0 0 F_IN
port 29 nsew
flabel metal1 32279 5743 32279 5743 0 FreeSans 1600 0 0 0 VCTRL2
port 39 nsew
flabel metal1 33470 8331 33470 8331 0 FreeSans 1600 0 0 0 VSS
port 40 nsew
flabel metal1 30024 14122 30024 14122 0 FreeSans 1600 0 0 0 VDD
port 41 nsew
flabel metal1 42870 4240 42870 4240 0 FreeSans 1600 0 0 0 VCTRL_IN
port 42 nsew
flabel metal1 43370 4280 43370 4280 0 FreeSans 1600 0 0 0 S4
port 43 nsew
flabel metal1 21788 13207 21788 13207 0 FreeSans 1600 0 0 0 S2
port 20 nsew
flabel metal1 21858 13590 21858 13590 0 FreeSans 1600 0 0 0 DN_INPUT
port 26 nsew
flabel metal1 19290 14218 19290 14218 0 FreeSans 1600 0 0 0 S1
port 23 nsew
flabel metal1 17988 6714 17988 6714 0 FreeSans 1600 0 0 0 S6
port 24 nsew
flabel metal1 26249 11574 26249 11574 0 FreeSans 1600 0 0 0 UP1
port 44 nsew
flabel metal1 26214 8908 26214 8908 0 FreeSans 1600 0 0 0 DN1
port 45 nsew
flabel metal1 22703 16344 22703 16344 0 FreeSans 1600 0 0 0 LF_OFFCHIP
port 49 nsew
flabel metal1 22694 16690 22694 16690 0 FreeSans 1600 0 0 0 S5
port 50 nsew
flabel metal1 56568 6749 56568 6749 0 FreeSans 1600 0 0 0 OUTB
port 51 nsew
flabel metal1 56817 2078 56817 2078 0 FreeSans 1600 0 0 0 OUT
port 52 nsew
flabel metal1 99070 -7610 99070 -7610 0 FreeSans 1600 0 0 0 OUT1
port 53 nsew
flabel metal1 99167 -991 99167 -991 0 FreeSans 1600 0 0 0 D16
port 54 nsew
flabel metal1 99137 -2090 99137 -2090 0 FreeSans 1600 0 0 0 D13
port 55 nsew
flabel metal1 99090 -2966 99090 -2966 0 FreeSans 1600 0 0 0 D12
port 56 nsew
flabel metal1 99146 -3471 99146 -3471 0 FreeSans 1600 0 0 0 D14
port 57 nsew
flabel metal1 99171 -4022 99171 -4022 0 FreeSans 1600 0 0 0 D15
port 58 nsew
flabel metal1 4423 -2365 4423 -2365 0 FreeSans 1600 0 0 0 S7
port 59 nsew
flabel metal1 4793 -4573 4793 -4573 0 FreeSans 1600 0 0 0 D4
port 60 nsew
flabel metal1 4742 -4063 4742 -4063 0 FreeSans 1600 0 0 0 D6
port 61 nsew
flabel metal1 4675 -3537 4675 -3537 0 FreeSans 1600 0 0 0 D1
port 62 nsew
flabel metal1 4723 -3078 4723 -3078 0 FreeSans 1600 0 0 0 D5
port 63 nsew
flabel metal1 4752 -2715 4752 -2715 0 FreeSans 1600 0 0 0 D0
port 64 nsew
flabel metal1 4646 -1595 4646 -1595 0 FreeSans 1600 0 0 0 D2
port 65 nsew
flabel metal1 4579 -1155 4579 -1155 0 FreeSans 1600 0 0 0 D3
port 66 nsew
flabel metal1 -3298 62608 -3298 62608 0 FreeSans 1600 0 0 0 D11
port 67 nsew
flabel metal1 -3395 52547 -3395 52547 0 FreeSans 1600 0 0 0 D8
port 68 nsew
flabel metal1 -3154 44010 -3154 44010 0 FreeSans 1600 0 0 0 D7
port 69 nsew
flabel metal1 -3184 43467 -3184 43467 0 FreeSans 1600 0 0 0 D9
port 70 nsew
flabel metal1 -3049 36634 -3049 36634 0 FreeSans 1600 0 0 0 D10
port 71 nsew
flabel metal1 -3814 24857 -3814 24857 0 FreeSans 1600 0 0 0 PRE_SCALAR
port 72 nsew
flabel metal1 4188 9245 4188 9245 0 FreeSans 1600 0 0 0 UP_OUT
port 73 nsew
flabel metal1 5730 4634 5730 4634 0 FreeSans 1600 0 0 0 DN_OUT
port 74 nsew
flabel metal2 21999 15127 21999 15127 0 FreeSans 1600 0 0 0 UP
port 75 nsew
flabel metal2 22016 14545 22016 14545 0 FreeSans 1600 0 0 0 DN
port 76 nsew
flabel metal1 99365 4556 99365 4556 0 FreeSans 1600 0 0 0 VDD_TEST
port 77 nsew
flabel metal1 39830 6510 39830 6510 0 FreeSans 1600 0 0 0 VCTRL_OBV
port 78 nsew
flabel metal1 18550 7330 18550 7330 0 FreeSans 1600 0 0 0 DIV_OUT2
port 79 nsew
flabel metal1 13110 -7700 13110 -7700 0 FreeSans 1600 0 0 0 Q02
port 80 nsew
flabel metal1 13860 -10180 13860 -10180 0 FreeSans 1600 0 0 0 Q07
port 81 nsew
flabel metal1 28770 -7800 28770 -7800 0 FreeSans 1600 0 0 0 Q01
port 82 nsew
flabel metal1 14210 -15910 14210 -15910 0 FreeSans 1600 0 0 0 Q05
port 83 nsew
flabel metal1 13110 -12310 13110 -12310 0 FreeSans 1600 0 0 0 Q06
port 84 nsew
flabel metal1 28860 -12250 28860 -12250 0 FreeSans 1600 0 0 0 Q03
port 85 nsew
flabel metal1 28010 -15010 28010 -15010 0 FreeSans 1600 0 0 0 Q04
port 86 nsew
flabel metal1 28920 -18000 28920 -18000 0 FreeSans 1600 0 0 0 P02
port 87 nsew
flabel metal1 6410 -8020 6410 -8020 0 FreeSans 1600 0 0 0 LD0
port 88 nsew
flabel metal1 43780 -18390 43780 -18390 0 FreeSans 1600 0 0 0 OUT01
port 89 nsew
flabel metal1 95190 -18410 95190 -18410 0 FreeSans 3200 0 0 0 OUT11
port 91 nsew
flabel metal1 57550 -8180 57550 -8180 0 FreeSans 3200 0 0 0 LD1
port 93 nsew
flabel metal1 64250 -7650 64250 -7650 0 FreeSans 3200 0 0 0 Q12
port 94 nsew
flabel metal1 79910 -7950 79910 -7950 0 FreeSans 3200 0 0 0 Q11
port 95 nsew
flabel metal1 64260 -11900 64260 -11900 0 FreeSans 3200 0 0 0 Q16
port 96 nsew
flabel metal1 80010 -12090 80010 -12090 0 FreeSans 3200 0 0 0 Q13
port 97 nsew
flabel metal1 65360 -15960 65360 -15960 0 FreeSans 3200 0 0 0 Q15
port 98 nsew
flabel metal1 79160 -15880 79160 -15880 0 FreeSans 3200 0 0 0 Q14
port 99 nsew
flabel metal1 65000 -10230 65000 -10230 0 FreeSans 3200 0 0 0 Q17
port 100 nsew
flabel metal1 80070 -17980 80070 -17980 0 FreeSans 3200 0 0 0 P12
port 101 nsew
flabel metal1 58470 -2667 58470 -2667 0 FreeSans 3200 0 0 0 D17G
port 102 nsew
flabel metal1 69038 -3769 69038 -3769 0 FreeSans 3200 0 0 0 D16G
port 103 nsew
flabel metal1 -4324 61270 -4324 61270 0 FreeSans 3200 0 0 0 D27G
port 104 nsew
flabel metal1 -4077 52130 -4077 52130 0 FreeSans 3200 0 0 0 D26G
port 105 nsew
flabel metal1 8667 22935 8667 22935 0 FreeSans 3200 0 0 0 OUT21
port 106 nsew
flabel metal1 4687 55482 4687 55482 0 FreeSans 3200 0 0 0 Q26
port 108 nsew
flabel metal1 2862 54749 2862 54749 0 FreeSans 3200 0 0 0 Q27
port 109 nsew
flabel metal1 8628 54398 8628 54398 0 FreeSans 3200 0 0 0 Q25
port 110 nsew
flabel metal1 -561 55487 -561 55487 0 FreeSans 3200 0 0 0 Q22
port 111 nsew
flabel metal1 -1095 48432 -1095 48432 0 FreeSans 3200 0 0 0 LD2
port 112 nsew
flabel metal1 137 39812 137 39812 0 FreeSans 3200 0 0 0 Q21
port 114 nsew
flabel metal1 4469 39744 4469 39744 0 FreeSans 3200 0 0 0 Q23
port 115 nsew
flabel metal1 7673 40583 7673 40583 0 FreeSans 3200 0 0 0 Q24
port 116 nsew
flabel metal1 48873 -14249 48873 -14249 0 FreeSans 1600 0 0 0 DIV_OUT
port 117 nsew
flabel metal1 2488 10382 2488 10382 0 FreeSans 1600 0 0 0 ITAIL
port 118 nsew
flabel metal1 5143 15231 5143 15231 0 FreeSans 1600 0 0 0 ITAIL_SINK
port 120 nsew
flabel metal1 53770 15520 53770 15520 0 FreeSans 1600 0 0 0 A1
port 121 nsew
flabel metal1 5149 16633 5149 16633 0 FreeSans 1600 0 0 0 ITAIL_SRC
port 119 nsew
flabel metal2 2480 16670 2480 16670 0 FreeSans 1600 0 0 0 A0
port 122 nsew
flabel metal2 2530 15190 2530 15190 0 FreeSans 1600 0 0 0 A3
port 123 nsew
flabel metal1 1916 15531 1916 15531 0 FreeSans 480 180 0 0 G_sink_up
port 4 nsew
flabel metal1 1919 15268 1919 15268 0 FreeSans 480 180 0 0 G_sink_dn
port 5 nsew
flabel metal1 1382 15902 1382 15902 0 FreeSans 480 180 0 0 G_source_dn
port 2 nsew
flabel metal1 1578 15993 1578 15993 0 FreeSans 480 180 0 0 G_source_up
port 1 nsew
flabel metal2 2100 14450 2100 14450 0 FreeSans 1600 0 0 0 G1_2
port 124 nsew
flabel metal2 1230 14410 1230 14410 0 FreeSans 1600 0 0 0 SD0_1
port 125 nsew
flabel metal2 1970 11950 1970 11950 0 FreeSans 1600 0 0 0 SD2_1
port 126 nsew
flabel metal1 1720 10740 1720 10740 0 FreeSans 1600 0 0 0 G2_1
port 127 nsew
flabel metal2 940 13900 940 13900 0 FreeSans 1600 0 0 0 G1_1
port 128 nsew
flabel metal2 -170 15280 -170 15280 0 FreeSans 1600 0 0 0 SD01
port 129 nsew
<< end >>
