* NGSPICE file created from TG_magic_flat.ext - technology: gf180mcuC

.subckt TG_magic_flat B VDD VSS CLK A
X0 B CLK.t0 A.t6 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 B a_267_n568.t6 A.t33 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 B a_267_n568.t7 A.t34 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 A a_267_n568.t8 B.t35 VDD.t6 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X4 A a_267_n568.t9 B.t13 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 B a_267_n568.t10 A.t14 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X6 B CLK.t1 A.t5 VSS.t8 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X7 B a_267_n568.t11 A.t15 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X8 A a_267_n568.t12 B.t18 VDD.t5 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 A CLK.t2 B.t10 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X10 B a_267_n568.t13 A.t19 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X11 B a_267_n568.t14 A.t20 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X12 B CLK.t3 A.t4 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X13 A a_267_n568.t15 B.t21 VDD.t5 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X14 A a_267_n568.t16 B.t22 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X15 A CLK.t5 B.t8 VSS.t6 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X16 B a_267_n568.t17 A.t23 VDD.t8 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X17 B a_267_n568.t18 A.t30 VDD.t10 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X18 B CLK.t6 A.t3 VSS.t5 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X19 A a_267_n568.t19 B.t31 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X20 B a_267_n568.t20 A.t32 VDD.t8 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X21 A CLK.t9 B.t6 VSS.t2 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X22 B a_267_n568.t21 A.t24 VDD.t8 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X23 B CLK.t11 A.t2 VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X24 A a_267_n568.t22 B.t25 VDD.t6 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X25 A CLK.t12 B.t4 VSS.t0 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X26 A a_267_n568.t23 B.t16 VDD.t5 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X27 B a_267_n568.t24 A.t17 VDD.t9 pfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X28 B a_267_n568.t25 A.t28 VDD.t8 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X29 A a_267_n568.t26 B.t29 VDD.t6 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X30 A CLK.t14 B.t3 VSS.t2 nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X31 A a_267_n568.t27 B.t26 VDD.t7 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X32 B CLK.t16 A.t1 VSS.t1 nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X33 A a_267_n568.t28 B.t27 VDD.t6 pfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X34 A CLK.t17 B.t1 VSS.t0 nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X35 A a_267_n568.t29 B.t0 VDD.t5 pfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
R0 CLK.t8 CLK.t16 83.8201
R1 CLK.n6 CLK.t10 52.6648
R2 CLK.t7 CLK.t13 43.8005
R3 CLK.t15 CLK.t7 43.8005
R4 CLK.t10 CLK.t15 43.8005
R5 CLK.t4 CLK.t8 43.8005
R6 CLK.n6 CLK.t4 23.2041
R7 CLK CLK.n6 21.9984
R8 CLK.n0 CLK.t12 21.9005
R9 CLK.n0 CLK.t17 21.9005
R10 CLK.n1 CLK.t0 21.9005
R11 CLK.n1 CLK.t1 21.9005
R12 CLK.n2 CLK.t2 21.9005
R13 CLK.n2 CLK.t5 21.9005
R14 CLK.n3 CLK.t3 21.9005
R15 CLK.n3 CLK.t6 21.9005
R16 CLK.n4 CLK.t9 21.9005
R17 CLK.n4 CLK.t14 21.9005
R18 CLK.n5 CLK.t11 21.9005
R19 CLK.t16 CLK.n5 21.9005
R20 CLK.n1 CLK.n0 15.8172
R21 CLK.n2 CLK.n1 15.8172
R22 CLK.n3 CLK.n2 15.8172
R23 CLK.n4 CLK.n3 15.8172
R24 CLK.n5 CLK.n4 15.8172
R25 A.n47 A.n45 5.44589
R26 A A.n52 5.33254
R27 A.n26 A.n25 5.07789
R28 A.n51 A.t2 4.7885
R29 A.n50 A.t1 4.7885
R30 A.n47 A.n46 4.7885
R31 A.n31 A.t33 4.4205
R32 A.n32 A.t17 4.4205
R33 A.n33 A.t15 4.4205
R34 A.n34 A.t34 4.4205
R35 A.n28 A.n22 4.4205
R36 A.n27 A.n23 4.4205
R37 A.n26 A.n24 4.4205
R38 A.n44 A.n41 3.80789
R39 A.n39 A.n36 3.80789
R40 A.n8 A.n7 3.25789
R41 A.n19 A.n18 3.25789
R42 A.n44 A.n43 3.1505
R43 A.n39 A.n38 3.1505
R44 A.n8 A.n5 2.6005
R45 A.n9 A.n3 2.6005
R46 A.n10 A.n1 2.6005
R47 A.n19 A.n16 2.6005
R48 A.n20 A.n14 2.6005
R49 A.n21 A.n12 2.6005
R50 A.n1 A.t24 1.8205
R51 A.n1 A.n0 1.8205
R52 A.n3 A.t23 1.8205
R53 A.n3 A.n2 1.8205
R54 A.n5 A.t28 1.8205
R55 A.n5 A.n4 1.8205
R56 A.n7 A.t32 1.8205
R57 A.n7 A.n6 1.8205
R58 A.n12 A.t20 1.8205
R59 A.n12 A.n11 1.8205
R60 A.n14 A.t14 1.8205
R61 A.n14 A.n13 1.8205
R62 A.n16 A.t30 1.8205
R63 A.n16 A.n15 1.8205
R64 A.n18 A.t19 1.8205
R65 A.n18 A.n17 1.8205
R66 A.n43 A.t5 1.6385
R67 A.n43 A.n42 1.6385
R68 A.n41 A.t6 1.6385
R69 A.n41 A.n40 1.6385
R70 A.n38 A.t3 1.6385
R71 A.n38 A.n37 1.6385
R72 A.n36 A.t4 1.6385
R73 A.n36 A.n35 1.6385
R74 A.n48 A.n47 0.884196
R75 A.n50 A.n49 0.884196
R76 A.n29 A.n28 0.882239
R77 A.n31 A.n30 0.882239
R78 A.n52 A.n51 0.8105
R79 A.n10 A.n9 0.657891
R80 A.n9 A.n8 0.657891
R81 A.n21 A.n20 0.657891
R82 A.n20 A.n19 0.657891
R83 A.n28 A.n27 0.657891
R84 A.n27 A.n26 0.657891
R85 A.n32 A.n31 0.657891
R86 A.n33 A.n32 0.657891
R87 A.n34 A.n33 0.657891
R88 A.n51 A.n50 0.657891
R89 A.n49 A.n48 0.6005
R90 A.n30 A.n29 0.6005
R91 A.n48 A.n44 0.284196
R92 A.n49 A.n39 0.284196
R93 A.n30 A.n10 0.282239
R94 A.n29 A.n21 0.282239
R95 A.n52 A.n34 0.237239
R96 B.n39 B.n38 3.80789
R97 B.n49 B.n48 3.80789
R98 B.n44 B.n43 3.80789
R99 B.n4 B.n1 3.25789
R100 B.n15 B.n12 3.25789
R101 B.n27 B.n24 3.25789
R102 B.n39 B.n36 3.1505
R103 B.n49 B.n46 3.1505
R104 B.n44 B.n41 3.1505
R105 B.n34 B.n22 3.05463
R106 B.n7 B.n6 2.6005
R107 B.n4 B.n3 2.6005
R108 B.n10 B.n9 2.6005
R109 B.n15 B.n14 2.6005
R110 B.n18 B.n17 2.6005
R111 B.n21 B.n20 2.6005
R112 B.n27 B.n26 2.6005
R113 B.n30 B.n29 2.6005
R114 B.n33 B.n32 2.6005
R115 B.n32 B.t25 1.8205
R116 B.n32 B.n31 1.8205
R117 B.n29 B.t27 1.8205
R118 B.n29 B.n28 1.8205
R119 B.n26 B.t29 1.8205
R120 B.n26 B.n25 1.8205
R121 B.n24 B.t35 1.8205
R122 B.n24 B.n23 1.8205
R123 B.n9 B.t18 1.8205
R124 B.n9 B.n8 1.8205
R125 B.n1 B.t0 1.8205
R126 B.n1 B.n0 1.8205
R127 B.n3 B.t16 1.8205
R128 B.n3 B.n2 1.8205
R129 B.n6 B.t21 1.8205
R130 B.n6 B.n5 1.8205
R131 B.n20 B.t26 1.8205
R132 B.n20 B.n19 1.8205
R133 B.n17 B.t13 1.8205
R134 B.n17 B.n16 1.8205
R135 B.n14 B.t22 1.8205
R136 B.n14 B.n13 1.8205
R137 B.n12 B.t31 1.8205
R138 B.n12 B.n11 1.8205
R139 B.n36 B.t4 1.6385
R140 B.n36 B.n35 1.6385
R141 B.n38 B.t1 1.6385
R142 B.n38 B.n37 1.6385
R143 B.n46 B.t6 1.6385
R144 B.n46 B.n45 1.6385
R145 B.n48 B.t3 1.6385
R146 B.n48 B.n47 1.6385
R147 B.n41 B.t10 1.6385
R148 B.n41 B.n40 1.6385
R149 B.n43 B.t8 1.6385
R150 B.n43 B.n42 1.6385
R151 B.n50 B.n49 0.896962
R152 B.n22 B.n10 0.86137
R153 B.n7 B.n4 0.657891
R154 B.n18 B.n15 0.657891
R155 B.n21 B.n18 0.657891
R156 B.n30 B.n27 0.657891
R157 B.n33 B.n30 0.657891
R158 B.n10 B.n7 0.655976
R159 B.n51 B.n50 0.613266
R160 B B.n52 0.468109
R161 B.n52 B.n51 0.432891
R162 B.n22 B.n21 0.323909
R163 B.n51 B.n39 0.284196
R164 B.n50 B.n44 0.284196
R165 B.n34 B.n33 0.272457
R166 B.n52 B.n34 0.0591957
R167 VSS.n2 VSS.t5 292.235
R168 VSS.n7 VSS.t3 185.615
R169 VSS.n1 VSS.t0 184.615
R170 VSS.n2 VSS.t6 180.065
R171 VSS.n12 VSS.t2 112.171
R172 VSS.n15 VSS.t1 67.8933
R173 VSS.n16 VSS.n14 13.1409
R174 VSS.n6 VSS.t7 5.44589
R175 VSS.n6 VSS.t4 4.7885
R176 VSS.n8 VSS.n7 2.6005
R177 VSS.n0 VSS.t8 2.6005
R178 VSS.n4 VSS.n3 2.6005
R179 VSS.n3 VSS.n2 2.6005
R180 VSS.n13 VSS.n5 2.6005
R181 VSS.n13 VSS.n12 2.6005
R182 VSS.n17 VSS.n16 2.6005
R183 VSS.n16 VSS.n15 2.6005
R184 VSS.n11 VSS.n10 2.6005
R185 VSS.n10 VSS.n9 2.6005
R186 VSS.n1 VSS.n0 1.86933
R187 VSS.n4 VSS.n1 0.489014
R188 VSS.n8 VSS.n6 0.477419
R189 VSS.n14 VSS.n13 0.430325
R190 VSS.n5 VSS.n4 0.11481
R191 VSS.n17 VSS.n11 0.11481
R192 VSS.n11 VSS.n8 0.11481
R193 VSS VSS.n17 0.11119
R194 VSS VSS.n5 0.00412069
R195 a_267_n568.t24 a_267_n568.t6 43.8005
R196 a_267_n568.t11 a_267_n568.t24 43.8005
R197 a_267_n568.t26 a_267_n568.t8 43.8005
R198 a_267_n568.t28 a_267_n568.t26 43.8005
R199 a_267_n568.t22 a_267_n568.t28 43.8005
R200 a_267_n568.t10 a_267_n568.t14 43.8005
R201 a_267_n568.t18 a_267_n568.t10 43.8005
R202 a_267_n568.t13 a_267_n568.t18 43.8005
R203 a_267_n568.t16 a_267_n568.t19 43.8005
R204 a_267_n568.t9 a_267_n568.t16 43.8005
R205 a_267_n568.t27 a_267_n568.t9 43.8005
R206 a_267_n568.t17 a_267_n568.t21 43.8005
R207 a_267_n568.t25 a_267_n568.t17 43.8005
R208 a_267_n568.t20 a_267_n568.t25 43.8005
R209 a_267_n568.t23 a_267_n568.t29 43.8005
R210 a_267_n568.t15 a_267_n568.t23 43.8005
R211 a_267_n568.t12 a_267_n568.t15 43.8005
R212 a_267_n568.n5 a_267_n568.t22 40.7345
R213 a_267_n568.t7 a_267_n568.n8 40.7345
R214 a_267_n568.n10 a_267_n568.n9 28.094
R215 a_267_n568.n5 a_267_n568.t13 25.5505
R216 a_267_n568.n6 a_267_n568.t27 25.5505
R217 a_267_n568.n7 a_267_n568.t20 25.5505
R218 a_267_n568.n8 a_267_n568.t12 25.5505
R219 a_267_n568.n9 a_267_n568.t11 21.9005
R220 a_267_n568.n9 a_267_n568.t7 21.9005
R221 a_267_n568.n6 a_267_n568.n5 15.1845
R222 a_267_n568.n7 a_267_n568.n6 15.1845
R223 a_267_n568.n8 a_267_n568.n7 15.1845
R224 a_267_n568.n14 a_267_n568.n13 5.44589
R225 a_267_n568.n2 a_267_n568.n0 5.07789
R226 a_267_n568.n15 a_267_n568.n14 4.7885
R227 a_267_n568.n12 a_267_n568.n11 4.4205
R228 a_267_n568.n2 a_267_n568.n1 4.4205
R229 a_267_n568.n4 a_267_n568.n3 4.4205
R230 a_267_n568.n14 a_267_n568.n12 1.1392
R231 a_267_n568.n4 a_267_n568.n2 0.657891
R232 a_267_n568.n10 a_267_n568.n4 0.286152
R233 a_267_n568.n12 a_267_n568.n10 0.282239
R234 VDD.n14 VDD.t8 59.8916
R235 VDD.n1 VDD.t6 42.1945
R236 VDD.n6 VDD.t0 40.6581
R237 VDD.n14 VDD.t7 36.9031
R238 VDD.n17 VDD.t5 22.989
R239 VDD.n11 VDD.t9 13.9146
R240 VDD.n16 VDD.n15 12.1031
R241 VDD.n3 VDD.t3 5.07789
R242 VDD.n5 VDD.t2 4.4205
R243 VDD.n4 VDD.t4 4.4205
R244 VDD.n3 VDD.t1 4.4205
R245 VDD.n0 VDD.t10 3.1505
R246 VDD.n15 VDD.n2 3.1505
R247 VDD.n15 VDD.n14 3.1505
R248 VDD.n19 VDD.n18 3.1505
R249 VDD.n18 VDD.n17 3.1505
R250 VDD.n13 VDD.n12 3.1505
R251 VDD.n12 VDD.n11 3.1505
R252 VDD.n10 VDD.n9 3.1505
R253 VDD.n9 VDD.n8 3.1505
R254 VDD.n7 VDD.n6 3.1505
R255 VDD.n1 VDD.n0 2.06641
R256 VDD.n2 VDD.n1 0.667563
R257 VDD.n5 VDD.n4 0.657891
R258 VDD.n4 VDD.n3 0.657891
R259 VDD.n7 VDD.n5 0.481332
R260 VDD.n19 VDD.n13 0.11481
R261 VDD.n13 VDD.n10 0.11481
R262 VDD.n10 VDD.n7 0.11481
R263 VDD VDD.n2 0.113776
R264 VDD.n18 VDD.n16 0.111026
R265 VDD VDD.n19 0.00153448
C0 VDD B 0.175f
C1 A CLK 0.256f
C2 VDD CLK 0.384f
C3 B CLK 0.155f
C4 VDD A 1.43f
C5 B A 4.86f
.ends

