magic
tech gf180mcuC
magscale 1 10
timestamp 1691518522
<< nwell >>
rect 37 220 1644 1873
<< pwell >>
rect 99 -636 379 36
rect 502 -636 1582 36
<< nmos >>
rect 211 -232 267 -32
rect 614 -232 670 -32
rect 774 -232 830 -32
rect 934 -232 990 -32
rect 1094 -232 1150 -32
rect 1254 -232 1310 -32
rect 1414 -232 1470 -32
rect 211 -568 267 -368
rect 614 -568 670 -368
rect 774 -568 830 -368
rect 934 -568 990 -368
rect 1094 -568 1150 -368
rect 1254 -568 1310 -368
rect 1414 -568 1470 -368
<< pmos >>
rect 211 1358 267 1558
rect 614 1358 670 1558
rect 774 1358 830 1558
rect 934 1358 990 1558
rect 1094 1358 1150 1558
rect 1254 1358 1310 1558
rect 1414 1358 1470 1558
rect 211 1022 267 1222
rect 614 1022 670 1222
rect 774 1022 830 1222
rect 934 1022 990 1222
rect 1094 1022 1150 1222
rect 1254 1022 1310 1222
rect 1414 1022 1470 1222
rect 211 686 267 886
rect 614 686 670 886
rect 774 686 830 886
rect 934 686 990 886
rect 1094 686 1150 886
rect 1254 686 1310 886
rect 1414 686 1470 886
rect 211 350 267 550
rect 614 350 670 550
rect 774 350 830 550
rect 934 350 990 550
rect 1094 350 1150 550
rect 1254 350 1310 550
rect 1414 350 1470 550
<< ndiff >>
rect 123 -45 211 -32
rect 123 -219 136 -45
rect 182 -219 211 -45
rect 123 -232 211 -219
rect 267 -45 355 -32
rect 267 -219 296 -45
rect 342 -219 355 -45
rect 267 -232 355 -219
rect 526 -45 614 -32
rect 526 -219 539 -45
rect 585 -219 614 -45
rect 526 -232 614 -219
rect 670 -45 774 -32
rect 670 -219 699 -45
rect 745 -219 774 -45
rect 670 -232 774 -219
rect 830 -45 934 -32
rect 830 -219 859 -45
rect 905 -219 934 -45
rect 830 -232 934 -219
rect 990 -45 1094 -32
rect 990 -219 1019 -45
rect 1065 -219 1094 -45
rect 990 -232 1094 -219
rect 1150 -45 1254 -32
rect 1150 -219 1179 -45
rect 1225 -219 1254 -45
rect 1150 -232 1254 -219
rect 1310 -45 1414 -32
rect 1310 -219 1339 -45
rect 1385 -219 1414 -45
rect 1310 -232 1414 -219
rect 1470 -45 1558 -32
rect 1470 -219 1499 -45
rect 1545 -219 1558 -45
rect 1470 -232 1558 -219
rect 123 -381 211 -368
rect 123 -555 136 -381
rect 182 -555 211 -381
rect 123 -568 211 -555
rect 267 -381 355 -368
rect 267 -555 296 -381
rect 342 -555 355 -381
rect 267 -568 355 -555
rect 526 -381 614 -368
rect 526 -555 539 -381
rect 585 -555 614 -381
rect 526 -568 614 -555
rect 670 -381 774 -368
rect 670 -555 699 -381
rect 745 -555 774 -381
rect 670 -568 774 -555
rect 830 -381 934 -368
rect 830 -555 859 -381
rect 905 -555 934 -381
rect 830 -568 934 -555
rect 990 -381 1094 -368
rect 990 -555 1019 -381
rect 1065 -555 1094 -381
rect 990 -568 1094 -555
rect 1150 -381 1254 -368
rect 1150 -555 1179 -381
rect 1225 -555 1254 -381
rect 1150 -568 1254 -555
rect 1310 -381 1414 -368
rect 1310 -555 1339 -381
rect 1385 -555 1414 -381
rect 1310 -568 1414 -555
rect 1470 -381 1558 -368
rect 1470 -555 1499 -381
rect 1545 -555 1558 -381
rect 1470 -568 1558 -555
<< pdiff >>
rect 123 1545 211 1558
rect 123 1371 136 1545
rect 182 1371 211 1545
rect 123 1358 211 1371
rect 267 1545 355 1558
rect 267 1371 296 1545
rect 342 1371 355 1545
rect 267 1358 355 1371
rect 526 1545 614 1558
rect 526 1371 539 1545
rect 585 1371 614 1545
rect 526 1358 614 1371
rect 670 1545 774 1558
rect 670 1371 699 1545
rect 745 1371 774 1545
rect 670 1358 774 1371
rect 830 1545 934 1558
rect 830 1371 859 1545
rect 905 1371 934 1545
rect 830 1358 934 1371
rect 990 1545 1094 1558
rect 990 1371 1019 1545
rect 1065 1371 1094 1545
rect 990 1358 1094 1371
rect 1150 1545 1254 1558
rect 1150 1371 1179 1545
rect 1225 1371 1254 1545
rect 1150 1358 1254 1371
rect 1310 1545 1414 1558
rect 1310 1371 1339 1545
rect 1385 1371 1414 1545
rect 1310 1358 1414 1371
rect 1470 1545 1558 1558
rect 1470 1371 1499 1545
rect 1545 1371 1558 1545
rect 1470 1358 1558 1371
rect 123 1209 211 1222
rect 123 1035 136 1209
rect 182 1035 211 1209
rect 123 1022 211 1035
rect 267 1209 355 1222
rect 267 1035 296 1209
rect 342 1035 355 1209
rect 267 1022 355 1035
rect 526 1209 614 1222
rect 526 1035 539 1209
rect 585 1035 614 1209
rect 526 1022 614 1035
rect 670 1209 774 1222
rect 670 1035 699 1209
rect 745 1035 774 1209
rect 670 1022 774 1035
rect 830 1209 934 1222
rect 830 1035 859 1209
rect 905 1035 934 1209
rect 830 1022 934 1035
rect 990 1209 1094 1222
rect 990 1035 1019 1209
rect 1065 1035 1094 1209
rect 990 1022 1094 1035
rect 1150 1209 1254 1222
rect 1150 1035 1179 1209
rect 1225 1035 1254 1209
rect 1150 1022 1254 1035
rect 1310 1209 1414 1222
rect 1310 1035 1339 1209
rect 1385 1035 1414 1209
rect 1310 1022 1414 1035
rect 1470 1209 1558 1222
rect 1470 1035 1499 1209
rect 1545 1035 1558 1209
rect 1470 1022 1558 1035
rect 123 873 211 886
rect 123 699 136 873
rect 182 699 211 873
rect 123 686 211 699
rect 267 873 355 886
rect 267 699 296 873
rect 342 699 355 873
rect 267 686 355 699
rect 526 873 614 886
rect 526 699 539 873
rect 585 699 614 873
rect 526 686 614 699
rect 670 873 774 886
rect 670 699 699 873
rect 745 699 774 873
rect 670 686 774 699
rect 830 873 934 886
rect 830 699 859 873
rect 905 699 934 873
rect 830 686 934 699
rect 990 873 1094 886
rect 990 699 1019 873
rect 1065 699 1094 873
rect 990 686 1094 699
rect 1150 873 1254 886
rect 1150 699 1179 873
rect 1225 699 1254 873
rect 1150 686 1254 699
rect 1310 873 1414 886
rect 1310 699 1339 873
rect 1385 699 1414 873
rect 1310 686 1414 699
rect 1470 873 1558 886
rect 1470 699 1499 873
rect 1545 699 1558 873
rect 1470 686 1558 699
rect 123 537 211 550
rect 123 363 136 537
rect 182 363 211 537
rect 123 350 211 363
rect 267 537 355 550
rect 267 363 296 537
rect 342 363 355 537
rect 267 350 355 363
rect 526 537 614 550
rect 526 363 539 537
rect 585 363 614 537
rect 526 350 614 363
rect 670 537 774 550
rect 670 363 699 537
rect 745 363 774 537
rect 670 350 774 363
rect 830 537 934 550
rect 830 363 859 537
rect 905 363 934 537
rect 830 350 934 363
rect 990 537 1094 550
rect 990 363 1019 537
rect 1065 363 1094 537
rect 990 350 1094 363
rect 1150 537 1254 550
rect 1150 363 1179 537
rect 1225 363 1254 537
rect 1150 350 1254 363
rect 1310 537 1414 550
rect 1310 363 1339 537
rect 1385 363 1414 537
rect 1310 350 1414 363
rect 1470 537 1558 550
rect 1470 363 1499 537
rect 1545 363 1558 537
rect 1470 350 1558 363
<< ndiffc >>
rect 136 -219 182 -45
rect 296 -219 342 -45
rect 539 -219 585 -45
rect 699 -219 745 -45
rect 859 -219 905 -45
rect 1019 -219 1065 -45
rect 1179 -219 1225 -45
rect 1339 -219 1385 -45
rect 1499 -219 1545 -45
rect 136 -555 182 -381
rect 296 -555 342 -381
rect 539 -555 585 -381
rect 699 -555 745 -381
rect 859 -555 905 -381
rect 1019 -555 1065 -381
rect 1179 -555 1225 -381
rect 1339 -555 1385 -381
rect 1499 -555 1545 -381
<< pdiffc >>
rect 136 1371 182 1545
rect 296 1371 342 1545
rect 539 1371 585 1545
rect 699 1371 745 1545
rect 859 1371 905 1545
rect 1019 1371 1065 1545
rect 1179 1371 1225 1545
rect 1339 1371 1385 1545
rect 1499 1371 1545 1545
rect 136 1035 182 1209
rect 296 1035 342 1209
rect 539 1035 585 1209
rect 699 1035 745 1209
rect 859 1035 905 1209
rect 1019 1035 1065 1209
rect 1179 1035 1225 1209
rect 1339 1035 1385 1209
rect 1499 1035 1545 1209
rect 136 699 182 873
rect 296 699 342 873
rect 539 699 585 873
rect 699 699 745 873
rect 859 699 905 873
rect 1019 699 1065 873
rect 1179 699 1225 873
rect 1339 699 1385 873
rect 1499 699 1545 873
rect 136 363 182 537
rect 296 363 342 537
rect 539 363 585 537
rect 699 363 745 537
rect 859 363 905 537
rect 1019 363 1065 537
rect 1179 363 1225 537
rect 1339 363 1385 537
rect 1499 363 1545 537
<< psubdiff >>
rect 67 -767 1614 -737
rect 67 -821 97 -767
rect 258 -821 318 -767
rect 479 -821 539 -767
rect 700 -821 760 -767
rect 921 -821 981 -767
rect 1142 -821 1202 -767
rect 1363 -821 1423 -767
rect 1584 -821 1614 -767
rect 67 -851 1614 -821
<< nsubdiff >>
rect 67 1813 1614 1843
rect 67 1759 97 1813
rect 258 1759 318 1813
rect 479 1759 539 1813
rect 700 1759 760 1813
rect 921 1759 981 1813
rect 1142 1759 1202 1813
rect 1363 1759 1423 1813
rect 1584 1759 1614 1813
rect 67 1729 1614 1759
<< psubdiffcont >>
rect 97 -821 258 -767
rect 318 -821 479 -767
rect 539 -821 700 -767
rect 760 -821 921 -767
rect 981 -821 1142 -767
rect 1202 -821 1363 -767
rect 1423 -821 1584 -767
<< nsubdiffcont >>
rect 97 1759 258 1813
rect 318 1759 479 1813
rect 539 1759 700 1813
rect 760 1759 921 1813
rect 981 1759 1142 1813
rect 1202 1759 1363 1813
rect 1423 1759 1584 1813
<< polysilicon >>
rect 211 1558 267 1602
rect 614 1558 670 1602
rect 774 1558 830 1602
rect 934 1558 990 1602
rect 1094 1558 1150 1602
rect 1254 1558 1310 1602
rect 1414 1558 1470 1602
rect 211 1222 267 1358
rect 614 1222 670 1358
rect 774 1222 830 1358
rect 934 1222 990 1358
rect 1094 1222 1150 1358
rect 1254 1222 1310 1358
rect 1414 1222 1470 1358
rect 211 886 267 1022
rect 614 886 670 1022
rect 774 886 830 1022
rect 934 886 990 1022
rect 1094 886 1150 1022
rect 1254 886 1310 1022
rect 1414 886 1470 1022
rect 211 550 267 686
rect 406 642 481 654
rect 614 642 670 686
rect 406 641 670 642
rect 406 595 421 641
rect 467 595 670 641
rect 406 594 670 595
rect 406 580 481 594
rect 614 550 670 594
rect 774 550 830 686
rect 934 550 990 686
rect 1094 550 1150 686
rect 1254 550 1310 686
rect 1414 550 1470 686
rect 42 70 118 82
rect 211 70 267 350
rect 614 279 670 350
rect 774 279 830 350
rect 934 279 990 350
rect 1094 279 1150 350
rect 1254 279 1310 350
rect 1414 279 1470 350
rect 614 229 1471 279
rect 42 68 267 70
rect 42 22 56 68
rect 104 22 267 68
rect 42 9 118 22
rect 211 -32 267 22
rect 614 -32 670 12
rect 774 -32 830 12
rect 934 -32 990 12
rect 1094 -32 1150 12
rect 1254 -32 1310 12
rect 1414 -32 1470 12
rect 211 -368 267 -232
rect 614 -276 670 -232
rect 774 -276 830 -232
rect 934 -276 990 -232
rect 1094 -276 1150 -232
rect 1254 -276 1310 -232
rect 1414 -276 1470 -232
rect 614 -324 1470 -276
rect 614 -368 670 -324
rect 774 -368 830 -324
rect 934 -368 990 -324
rect 1094 -368 1150 -324
rect 1254 -368 1310 -324
rect 1414 -368 1470 -324
rect 211 -588 267 -568
rect 614 -588 670 -568
rect 211 -644 670 -588
rect 774 -612 830 -568
rect 934 -612 990 -568
rect 1094 -612 1150 -568
rect 1254 -612 1310 -568
rect 1414 -612 1470 -568
<< polycontact >>
rect 421 595 467 641
rect 56 22 104 68
<< metal1 >>
rect 37 1813 1644 1873
rect 37 1759 97 1813
rect 258 1759 318 1813
rect 479 1759 539 1813
rect 700 1759 760 1813
rect 921 1759 981 1813
rect 1142 1759 1202 1813
rect 1363 1759 1423 1813
rect 1584 1759 1644 1813
rect 37 1699 1644 1759
rect 136 1545 182 1699
rect 539 1602 1545 1650
rect 136 1209 182 1371
rect 136 873 182 1035
rect 136 537 182 699
rect 136 352 182 363
rect 296 1545 342 1556
rect 296 1209 342 1371
rect 296 873 342 1035
rect 296 640 342 699
rect 539 1545 585 1602
rect 539 1209 585 1371
rect 539 873 585 1035
rect 406 641 481 654
rect 406 640 421 641
rect 296 595 421 640
rect 467 595 481 641
rect 296 594 481 595
rect 296 537 342 594
rect 406 580 481 594
rect 13 334 90 347
rect 13 312 24 334
rect -43 278 24 312
rect 80 278 90 334
rect -43 259 90 278
rect -43 258 13 259
rect 42 69 118 82
rect -43 68 118 69
rect -43 22 56 68
rect 104 22 118 68
rect -43 20 118 22
rect 42 9 118 20
rect 136 -45 182 -34
rect 136 -381 182 -219
rect 136 -707 182 -555
rect 296 -45 342 363
rect 539 537 585 699
rect 699 1545 745 1556
rect 699 1209 745 1371
rect 699 873 745 1035
rect 699 565 745 699
rect 698 537 745 565
rect 698 519 699 537
rect 405 333 482 345
rect 405 279 419 333
rect 473 329 482 333
rect 539 329 585 363
rect 473 282 585 329
rect 473 279 482 282
rect 405 267 482 279
rect 296 -381 342 -219
rect 296 -566 342 -555
rect 539 -45 585 282
rect 699 306 745 363
rect 859 1545 905 1602
rect 859 1209 905 1371
rect 859 873 905 1035
rect 859 537 905 699
rect 1019 1545 1065 1556
rect 1019 1209 1065 1371
rect 1019 873 1065 1035
rect 1019 537 1065 699
rect 859 352 905 363
rect 1018 306 1065 363
rect 1179 1545 1225 1602
rect 1179 1209 1225 1371
rect 1179 873 1225 1035
rect 1179 537 1225 699
rect 1339 1545 1385 1556
rect 1339 1209 1385 1371
rect 1339 873 1385 1035
rect 1339 537 1385 699
rect 1179 352 1225 363
rect 1338 306 1385 363
rect 1499 1545 1545 1602
rect 1499 1209 1545 1371
rect 1499 873 1545 1035
rect 1499 537 1545 699
rect 1499 352 1545 363
rect 699 304 1385 306
rect 699 260 1724 304
rect 1339 258 1724 260
rect 1339 60 1385 258
rect 539 -381 585 -219
rect 539 -613 585 -555
rect 699 13 1385 60
rect 699 -45 745 13
rect 699 -381 745 -219
rect 699 -566 745 -555
rect 859 -45 905 -34
rect 859 -381 905 -219
rect 859 -613 905 -555
rect 1019 -45 1065 13
rect 1019 -381 1065 -219
rect 1019 -566 1065 -555
rect 1179 -45 1225 -34
rect 1179 -381 1225 -219
rect 1179 -613 1225 -555
rect 1339 -45 1385 13
rect 1339 -381 1385 -219
rect 1339 -566 1385 -555
rect 1499 -45 1545 -34
rect 1499 -381 1545 -219
rect 1499 -613 1545 -555
rect 539 -661 1545 -613
rect 37 -767 1644 -707
rect 37 -821 97 -767
rect 258 -821 318 -767
rect 479 -821 539 -767
rect 700 -821 760 -767
rect 921 -821 981 -767
rect 1142 -821 1202 -767
rect 1363 -821 1423 -767
rect 1584 -821 1644 -767
rect 37 -881 1644 -821
<< via1 >>
rect 24 278 80 334
rect 419 279 473 333
<< metal2 >>
rect 13 334 90 347
rect 405 334 482 345
rect 13 278 24 334
rect 80 333 482 334
rect 80 279 419 333
rect 473 279 482 333
rect 80 278 482 279
rect 13 259 90 278
rect 405 267 482 278
<< labels >>
flabel metal1 1624 282 1624 282 0 FreeSans 800 0 0 0 B
port 12 nsew
flabel nsubdiffcont 842 1781 842 1781 0 FreeSans 800 0 0 0 VDD
port 13 nsew
flabel psubdiffcont 833 -798 833 -798 0 FreeSans 800 0 0 0 VSS
port 14 nsew
flabel metal1 38 42 38 42 0 FreeSans 800 0 0 0 CLK
port 15 nsew
flabel metal1 10 287 10 287 0 FreeSans 800 0 0 0 A
port 17 nsew
<< end >>
