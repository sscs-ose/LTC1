magic
tech gf180mcuD
magscale 1 5
timestamp 1713338890
<< checkpaint >>
rect -1329 -1019 1329 1019
<< metal1 >>
rect -329 13 329 19
rect -329 -13 -323 13
rect -297 -13 -261 13
rect -235 -13 -199 13
rect -173 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 173 13
rect 199 -13 235 13
rect 261 -13 297 13
rect 323 -13 329 13
rect -329 -19 329 -13
<< via1 >>
rect -323 -13 -297 13
rect -261 -13 -235 13
rect -199 -13 -173 13
rect -137 -13 -111 13
rect -75 -13 -49 13
rect -13 -13 13 13
rect 49 -13 75 13
rect 111 -13 137 13
rect 173 -13 199 13
rect 235 -13 261 13
rect 297 -13 323 13
<< metal2 >>
rect -329 13 329 19
rect -329 -13 -323 13
rect -297 -13 -261 13
rect -235 -13 -199 13
rect -173 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 173 13
rect 199 -13 235 13
rect 261 -13 297 13
rect 323 -13 329 13
rect -329 -19 329 -13
<< end >>
