** sch_path: /home/shahid/GF180Projects/Layout/Xschem/VCO/PLL_TOP_FINAL/TB_TOP_MUX_F8_sch.sch
**.subckt TB_TOP_MUX_F8_sch
V1 VSS GND 0
V3 VCTRL2 VSS 3.3
V4 VCTRL_IN VSS 0.6
V6 F_IN VSS pulse(0 3.3 0 100p 100p 50n 100n)
I4 VDD ITAIL 100u
V8 S1 VSS 0
V9 S2 VSS 0
V10 S3 VSS 0
V11 S4 VSS 0
V12 S6 VSS 0
V13 DN_INPUT VSS pulse(0 3.3 10n 100p 100p 500n 1000n)
V14 UP_INPUT VSS pulse(0 3.3 0 100p 100p 500n 1000n)
V15 VDD_TEST VSS 3.3
C1 LF_OFFCHIP VSS 11.27p m=1
R1 LF_OFFCHIP net1 74k m=1
C2 net1 VSS 239p m=1
V16 S5 VSS 0
V17 D0 VSS 0
V18 D1 VSS 3.3
V19 D2 VSS 0
V20 D3 VSS 0
V21 D4 VSS 0
V22 D5 VSS 3.3
V23 D6 VSS 3.3
V29 D12 VSS 0
V30 D13 VSS 0
V31 D14 VSS 0
V32 D15 VSS 3.3
V2 S7 VSS 0
V5 VDD VSS pwl(0 0 0.05US 0 0.050001US 3.3)
V7 D7 VSS 0
V34 D8 VSS 0
V35 D9 VSS 0
V36 D10 VSS 3.3
V24 DIV_OUT2 VSS pulse(0 3.3 700n 100p 100p 500n 1000n)
x1 VDD_TEST D12 D0 UP_INPUT D13 D1 DN_INPUT VSS D14 D2 PRE_SCALAR UP_OUT D15 D3 F_IN DN_OUT GND D4 ITAIL DIV_OUT D5 S1 S6 D6
+ VCTRL_IN D7 VCTRL2 S2 D8 S3 OUT D9 OUTB S4 LF_OFFCHIP D10 S5 S7 VSS OUT1 DIV_OUT2 GND GND GND GND VDD pex_PLL_TOP_MUX_8
**** begin user architecture code


*.include pex_A_MUX.spice
*.include pex_VCO_DFF_C.spice
*.include Tappered-Buffer_1_pex.spice
*.include pex_PFD_T2.spice
*.include pex_CP.spice
*.include Res_74k_pex.spice
*.include pex_cap_11p.spice
*.include pex_cap_240p.spice
.include pex_PLL_TOP_MUX_8.spice
*.include pex_7b_divider_magic.spice
*.include pex_PLL_TOP_MUX_2.spice
*.include Tappered-Buffer_1_pex.spice
*.option RSHUNT=1e18
**.option ABSTOL=1e-12
**.option VNTOL=1e-12
**.option CHGTOL=1e-14
**.option RELTOL=1e-5
.option gmin=1e-15
**.option trtol=1
**.OPTION ITL4=500
.control
save all
save x1.vco_dff_c_0.vctrl.t19
+ x1.pre_scalar.n0
+ pre_scalar
+ x1.vss.t6260
+ x1.vdd.n7823
+ x1.vctrl_in.t6
+ x1.vctrl2.t62
+ x1.vco_dff_c_0.vco_c_0.outb.t53
+ x1.vco_dff_c_0.vco_c_0.inv_2_5.in.n34
+ x1.vco_dff_c_0.vco_c_0.inv_2_3.out.n2
+ x1.vco_dff_c_0.vco_c_0.inv_2_2.in.n30
+ x1.vco_dff_c_0.vco_c_0.inv_2_0.in.n51
+ x1.vco_dff_c_0.outb.t31
+ x1.vco_dff_c_0.out.t10
+ x1.up_out.t60
+ x1.up_input.n12
+ x1.up1.n10
+ x1.up.n28
+ x1.dn
+ x1.a_mux_6.in1.n194
+ x1.a_mux_5.in1.t163
+ x1.a_mux_2.out.n14
+ x1.a_mux_1.out
+ x1.a_mux_6.out
+ x1.7b_divider_magic_2.p2_gen_magic_0.dff_magic_0.tg_magic_3.out
+ x1.7b_divider_magic_2.p2_gen_magic_0.dff_magic_0.tg_magic_3.clk
+ x1.7b_divider_magic_2.p2_gen_magic_0.dff_magic_0.tg_magic_2.in.n10
+ x1.7b_divider_magic_2.p2.t16
+ x1.7b_divider_magic_2.out1.t8
+ x1.7b_divider_magic_2.divide_by_2_1.tg_magic_3.out
+ x1.7b_divider_magic_2.divide_by_2_1.tg_magic_3.clk
+ x1.7b_divider_magic_1.p2_gen_magic_0.dff_magic_0.tg_magic_1.in.n19
+ x1.7b_divider_magic_1.ld
+ x1.7b_divider_magic_1.divide_by_2_1.tg_magic_2.in.n14
+ x1.7b_divider_magic_1.divide_by_2_0.tg_magic_3.out
+ x1.7b_divider_magic_1.divide_by_2_0.tg_magic_3.in
+ x1.7b_divider_magic_0.out1
+ x1.7b_divider_magic_0.ld.n38
+ x1.vctrl_obv
+ x1.a_mux_6.out.n27
+ out1
+ out
+ outb
+ net1
+ lf_offchip
+ itail1
+ itail
+ f_in
+ dn_out
+ up_out
+ dn_input
+ div_out
*set ngbehavior=hsa
*set ng_nomodcheck
tran 500n 130u
write TB_TOP_MUX_F7_sch.raw
.endc



.include /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice moscap_typical
.lib /home/shahid/OSPDKs/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical

**** end user architecture code
**.ends
.GLOBAL GND
.end
