magic
tech gf180mcuC
magscale 1 10
timestamp 1695285543
<< nwell >>
rect -2839 5952 -2275 6462
rect -2076 5952 -1512 6462
rect -1265 5952 -701 6462
rect -2839 4981 -2275 5491
rect -2076 4981 -1512 5491
rect -1265 4981 -701 5491
rect -2839 4006 -2275 4516
rect -2076 4005 -1512 4515
rect -1265 4005 -701 4515
<< pwell >>
rect -2548 5924 -2488 5925
rect -1785 5924 -1725 5925
rect -974 5924 -914 5925
rect -2548 5880 -2485 5924
rect -1785 5880 -1722 5924
rect -974 5880 -911 5924
rect -2777 5644 -2337 5880
rect -2014 5644 -1574 5880
rect -1203 5644 -763 5880
rect -2548 4953 -2488 4954
rect -1785 4953 -1725 4954
rect -974 4953 -914 4954
rect -2548 4909 -2485 4953
rect -1785 4909 -1722 4953
rect -974 4909 -911 4953
rect -2777 4673 -2337 4909
rect -2014 4673 -1574 4909
rect -1203 4673 -763 4909
rect -2548 3978 -2488 3979
rect -446 3978 4332 7401
rect -2548 3934 -2485 3978
rect -1785 3977 -1725 3978
rect -974 3977 -914 3978
rect -2777 3698 -2337 3934
rect -1785 3933 -1722 3977
rect -974 3933 -911 3977
rect -446 3967 3704 3978
rect -2014 3697 -1574 3933
rect -1203 3697 -763 3933
rect -446 3898 3732 3967
rect 3783 3963 4332 3978
rect 3798 3898 4332 3963
rect -446 3633 4332 3898
rect -2839 2762 3809 3138
rect -2839 2271 3809 2647
<< nmos >>
rect 317 6838 417 6958
rect 521 6838 621 6958
rect 725 6838 825 6958
rect 929 6838 1029 6958
rect 1133 6838 1233 6958
rect 1337 6838 1437 6958
rect 1541 6838 1641 6958
rect 1745 6838 1845 6958
rect 1949 6838 2049 6958
rect 2153 6838 2253 6958
rect 2357 6838 2457 6958
rect 2561 6838 2661 6958
rect 2765 6838 2865 6958
rect 2969 6838 3069 6958
rect 3173 6838 3273 6958
rect 3377 6838 3477 6958
rect 317 6433 417 6553
rect 521 6433 621 6553
rect 725 6433 825 6553
rect 929 6433 1029 6553
rect 1133 6433 1233 6553
rect 1337 6433 1437 6553
rect 1541 6433 1641 6553
rect 1745 6433 1845 6553
rect 1949 6433 2049 6553
rect 2153 6433 2253 6553
rect 2357 6433 2457 6553
rect 2561 6433 2661 6553
rect 2765 6433 2865 6553
rect 2969 6433 3069 6553
rect 3173 6433 3273 6553
rect 3377 6433 3477 6553
rect 317 6041 417 6161
rect 521 6041 621 6161
rect 725 6041 825 6161
rect 929 6041 1029 6161
rect 1133 6041 1233 6161
rect 1337 6041 1437 6161
rect 1541 6041 1641 6161
rect 1745 6041 1845 6161
rect 1949 6041 2049 6161
rect 2153 6041 2253 6161
rect 2357 6041 2457 6161
rect 2561 6041 2661 6161
rect 2765 6041 2865 6161
rect 2969 6041 3069 6161
rect 3173 6041 3273 6161
rect 3377 6041 3477 6161
rect -2665 5712 -2609 5812
rect -2505 5712 -2449 5812
rect -1902 5712 -1846 5812
rect -1742 5712 -1686 5812
rect -1091 5712 -1035 5812
rect -931 5712 -875 5812
rect 317 5636 417 5756
rect 521 5636 621 5756
rect 725 5636 825 5756
rect 929 5636 1029 5756
rect 1133 5636 1233 5756
rect 1337 5636 1437 5756
rect 1541 5636 1641 5756
rect 1745 5636 1845 5756
rect 1949 5636 2049 5756
rect 2153 5636 2253 5756
rect 2357 5636 2457 5756
rect 2561 5636 2661 5756
rect 2765 5636 2865 5756
rect 2969 5636 3069 5756
rect 3173 5636 3273 5756
rect 3377 5636 3477 5756
rect 317 5244 417 5364
rect 521 5244 621 5364
rect 725 5244 825 5364
rect 929 5244 1029 5364
rect 1133 5244 1233 5364
rect 1337 5244 1437 5364
rect 1541 5244 1641 5364
rect 1745 5244 1845 5364
rect 1949 5244 2049 5364
rect 2153 5244 2253 5364
rect 2357 5244 2457 5364
rect 2561 5244 2661 5364
rect 2765 5244 2865 5364
rect 2969 5244 3069 5364
rect 3173 5244 3273 5364
rect 3377 5244 3477 5364
rect -2665 4741 -2609 4841
rect -2505 4741 -2449 4841
rect -1902 4741 -1846 4841
rect -1742 4741 -1686 4841
rect -1091 4741 -1035 4841
rect -931 4741 -875 4841
rect 317 4839 417 4959
rect 521 4839 621 4959
rect 725 4839 825 4959
rect 929 4839 1029 4959
rect 1133 4839 1233 4959
rect 1337 4839 1437 4959
rect 1541 4839 1641 4959
rect 1745 4839 1845 4959
rect 1949 4839 2049 4959
rect 2153 4839 2253 4959
rect 2357 4839 2457 4959
rect 2561 4839 2661 4959
rect 2765 4839 2865 4959
rect 2969 4839 3069 4959
rect 3173 4839 3273 4959
rect 3377 4839 3477 4959
rect 317 4447 417 4567
rect 521 4447 621 4567
rect 725 4447 825 4567
rect 929 4447 1029 4567
rect 1133 4447 1233 4567
rect 1337 4447 1437 4567
rect 1541 4447 1641 4567
rect 1745 4447 1845 4567
rect 1949 4447 2049 4567
rect 2153 4447 2253 4567
rect 2357 4447 2457 4567
rect 2561 4447 2661 4567
rect 2765 4447 2865 4567
rect 2969 4447 3069 4567
rect 3173 4447 3273 4567
rect 3377 4447 3477 4567
rect -2665 3766 -2609 3866
rect -2505 3766 -2449 3866
rect 317 4042 417 4162
rect 521 4042 621 4162
rect 725 4042 825 4162
rect 929 4042 1029 4162
rect 1133 4042 1233 4162
rect 1337 4042 1437 4162
rect 1541 4042 1641 4162
rect 1745 4042 1845 4162
rect 1949 4042 2049 4162
rect 2153 4042 2253 4162
rect 2357 4042 2457 4162
rect 2561 4042 2661 4162
rect 2765 4042 2865 4162
rect 2969 4042 3069 4162
rect 3173 4042 3273 4162
rect 3377 4042 3477 4162
rect -1902 3765 -1846 3865
rect -1742 3765 -1686 3865
rect -1091 3765 -1035 3865
rect -931 3765 -875 3865
rect -2727 2830 -2627 3070
rect -2523 2830 -2423 3070
rect -2319 2830 -2219 3070
rect -2115 2830 -2015 3070
rect -1911 2830 -1811 3070
rect -1707 2830 -1607 3070
rect -1503 2830 -1403 3070
rect -1299 2830 -1199 3070
rect -1095 2830 -995 3070
rect -891 2830 -791 3070
rect -687 2830 -587 3070
rect -483 2830 -383 3070
rect -279 2830 -179 3070
rect -75 2830 25 3070
rect 129 2830 229 3070
rect 333 2830 433 3070
rect 537 2830 637 3070
rect 741 2830 841 3070
rect 945 2830 1045 3070
rect 1149 2830 1249 3070
rect 1353 2830 1453 3070
rect 1557 2830 1657 3070
rect 1761 2830 1861 3070
rect 1965 2830 2065 3070
rect 2169 2830 2269 3070
rect 2373 2830 2473 3070
rect 2577 2830 2677 3070
rect 2781 2830 2881 3070
rect 2985 2830 3085 3070
rect 3189 2830 3289 3070
rect 3393 2830 3493 3070
rect 3597 2830 3697 3070
rect -2727 2339 -2627 2579
rect -2523 2339 -2423 2579
rect -2319 2339 -2219 2579
rect -2115 2339 -2015 2579
rect -1911 2339 -1811 2579
rect -1707 2339 -1607 2579
rect -1503 2339 -1403 2579
rect -1299 2339 -1199 2579
rect -1095 2339 -995 2579
rect -891 2339 -791 2579
rect -687 2339 -587 2579
rect -483 2339 -383 2579
rect -279 2339 -179 2579
rect -75 2339 25 2579
rect 129 2339 229 2579
rect 333 2339 433 2579
rect 537 2339 637 2579
rect 741 2339 841 2579
rect 945 2339 1045 2579
rect 1149 2339 1249 2579
rect 1353 2339 1453 2579
rect 1557 2339 1657 2579
rect 1761 2339 1861 2579
rect 1965 2339 2065 2579
rect 2169 2339 2269 2579
rect 2373 2339 2473 2579
rect 2577 2339 2677 2579
rect 2781 2339 2881 2579
rect 2985 2339 3085 2579
rect 3189 2339 3289 2579
rect 3393 2339 3493 2579
rect 3597 2339 3697 2579
<< pmos >>
rect -2665 6082 -2609 6182
rect -2505 6082 -2449 6182
rect -1902 6082 -1846 6182
rect -1742 6082 -1686 6182
rect -1091 6082 -1035 6182
rect -931 6082 -875 6182
rect -2665 5111 -2609 5211
rect -2505 5111 -2449 5211
rect -1902 5111 -1846 5211
rect -1742 5111 -1686 5211
rect -1091 5111 -1035 5211
rect -931 5111 -875 5211
rect -2665 4136 -2609 4236
rect -2505 4136 -2449 4236
rect -1902 4135 -1846 4235
rect -1742 4135 -1686 4235
rect -1091 4135 -1035 4235
rect -931 4135 -875 4235
<< ndiff >>
rect 229 6945 317 6958
rect 229 6851 242 6945
rect 288 6851 317 6945
rect 229 6838 317 6851
rect 417 6945 521 6958
rect 417 6851 446 6945
rect 492 6851 521 6945
rect 417 6838 521 6851
rect 621 6945 725 6958
rect 621 6851 650 6945
rect 696 6851 725 6945
rect 621 6838 725 6851
rect 825 6945 929 6958
rect 825 6851 854 6945
rect 900 6851 929 6945
rect 825 6838 929 6851
rect 1029 6945 1133 6958
rect 1029 6851 1058 6945
rect 1104 6851 1133 6945
rect 1029 6838 1133 6851
rect 1233 6945 1337 6958
rect 1233 6851 1262 6945
rect 1308 6851 1337 6945
rect 1233 6838 1337 6851
rect 1437 6945 1541 6958
rect 1437 6851 1466 6945
rect 1512 6851 1541 6945
rect 1437 6838 1541 6851
rect 1641 6945 1745 6958
rect 1641 6851 1670 6945
rect 1716 6851 1745 6945
rect 1641 6838 1745 6851
rect 1845 6945 1949 6958
rect 1845 6851 1874 6945
rect 1920 6851 1949 6945
rect 1845 6838 1949 6851
rect 2049 6945 2153 6958
rect 2049 6851 2078 6945
rect 2124 6851 2153 6945
rect 2049 6838 2153 6851
rect 2253 6945 2357 6958
rect 2253 6851 2282 6945
rect 2328 6851 2357 6945
rect 2253 6838 2357 6851
rect 2457 6945 2561 6958
rect 2457 6851 2486 6945
rect 2532 6851 2561 6945
rect 2457 6838 2561 6851
rect 2661 6945 2765 6958
rect 2661 6851 2690 6945
rect 2736 6851 2765 6945
rect 2661 6838 2765 6851
rect 2865 6945 2969 6958
rect 2865 6851 2894 6945
rect 2940 6851 2969 6945
rect 2865 6838 2969 6851
rect 3069 6945 3173 6958
rect 3069 6851 3098 6945
rect 3144 6851 3173 6945
rect 3069 6838 3173 6851
rect 3273 6945 3377 6958
rect 3273 6851 3302 6945
rect 3348 6851 3377 6945
rect 3273 6838 3377 6851
rect 3477 6945 3565 6958
rect 3477 6851 3506 6945
rect 3552 6851 3565 6945
rect 3477 6838 3565 6851
rect 229 6540 317 6553
rect 229 6446 242 6540
rect 288 6446 317 6540
rect 229 6433 317 6446
rect 417 6540 521 6553
rect 417 6446 446 6540
rect 492 6446 521 6540
rect 417 6433 521 6446
rect 621 6540 725 6553
rect 621 6446 650 6540
rect 696 6446 725 6540
rect 621 6433 725 6446
rect 825 6540 929 6553
rect 825 6446 854 6540
rect 900 6446 929 6540
rect 825 6433 929 6446
rect 1029 6540 1133 6553
rect 1029 6446 1058 6540
rect 1104 6446 1133 6540
rect 1029 6433 1133 6446
rect 1233 6540 1337 6553
rect 1233 6446 1262 6540
rect 1308 6446 1337 6540
rect 1233 6433 1337 6446
rect 1437 6540 1541 6553
rect 1437 6446 1466 6540
rect 1512 6446 1541 6540
rect 1437 6433 1541 6446
rect 1641 6540 1745 6553
rect 1641 6446 1670 6540
rect 1716 6446 1745 6540
rect 1641 6433 1745 6446
rect 1845 6540 1949 6553
rect 1845 6446 1874 6540
rect 1920 6446 1949 6540
rect 1845 6433 1949 6446
rect 2049 6540 2153 6553
rect 2049 6446 2078 6540
rect 2124 6446 2153 6540
rect 2049 6433 2153 6446
rect 2253 6540 2357 6553
rect 2253 6446 2282 6540
rect 2328 6446 2357 6540
rect 2253 6433 2357 6446
rect 2457 6540 2561 6553
rect 2457 6446 2486 6540
rect 2532 6446 2561 6540
rect 2457 6433 2561 6446
rect 2661 6540 2765 6553
rect 2661 6446 2690 6540
rect 2736 6446 2765 6540
rect 2661 6433 2765 6446
rect 2865 6540 2969 6553
rect 2865 6446 2894 6540
rect 2940 6446 2969 6540
rect 2865 6433 2969 6446
rect 3069 6540 3173 6553
rect 3069 6446 3098 6540
rect 3144 6446 3173 6540
rect 3069 6433 3173 6446
rect 3273 6540 3377 6553
rect 3273 6446 3302 6540
rect 3348 6446 3377 6540
rect 3273 6433 3377 6446
rect 3477 6540 3565 6553
rect 3477 6446 3506 6540
rect 3552 6446 3565 6540
rect 3477 6433 3565 6446
rect 229 6148 317 6161
rect 229 6054 242 6148
rect 288 6054 317 6148
rect 229 6041 317 6054
rect 417 6148 521 6161
rect 417 6054 446 6148
rect 492 6054 521 6148
rect 417 6041 521 6054
rect 621 6148 725 6161
rect 621 6054 650 6148
rect 696 6054 725 6148
rect 621 6041 725 6054
rect 825 6148 929 6161
rect 825 6054 854 6148
rect 900 6054 929 6148
rect 825 6041 929 6054
rect 1029 6148 1133 6161
rect 1029 6054 1058 6148
rect 1104 6054 1133 6148
rect 1029 6041 1133 6054
rect 1233 6148 1337 6161
rect 1233 6054 1262 6148
rect 1308 6054 1337 6148
rect 1233 6041 1337 6054
rect 1437 6148 1541 6161
rect 1437 6054 1466 6148
rect 1512 6054 1541 6148
rect 1437 6041 1541 6054
rect 1641 6148 1745 6161
rect 1641 6054 1670 6148
rect 1716 6054 1745 6148
rect 1641 6041 1745 6054
rect 1845 6148 1949 6161
rect 1845 6054 1874 6148
rect 1920 6054 1949 6148
rect 1845 6041 1949 6054
rect 2049 6148 2153 6161
rect 2049 6054 2078 6148
rect 2124 6054 2153 6148
rect 2049 6041 2153 6054
rect 2253 6148 2357 6161
rect 2253 6054 2282 6148
rect 2328 6054 2357 6148
rect 2253 6041 2357 6054
rect 2457 6148 2561 6161
rect 2457 6054 2486 6148
rect 2532 6054 2561 6148
rect 2457 6041 2561 6054
rect 2661 6148 2765 6161
rect 2661 6054 2690 6148
rect 2736 6054 2765 6148
rect 2661 6041 2765 6054
rect 2865 6148 2969 6161
rect 2865 6054 2894 6148
rect 2940 6054 2969 6148
rect 2865 6041 2969 6054
rect 3069 6148 3173 6161
rect 3069 6054 3098 6148
rect 3144 6054 3173 6148
rect 3069 6041 3173 6054
rect 3273 6148 3377 6161
rect 3273 6054 3302 6148
rect 3348 6054 3377 6148
rect 3273 6041 3377 6054
rect 3477 6148 3565 6161
rect 3477 6054 3506 6148
rect 3552 6054 3565 6148
rect 3477 6041 3565 6054
rect -2753 5799 -2665 5812
rect -2753 5725 -2740 5799
rect -2694 5725 -2665 5799
rect -2753 5712 -2665 5725
rect -2609 5799 -2505 5812
rect -2609 5725 -2580 5799
rect -2534 5725 -2505 5799
rect -2609 5712 -2505 5725
rect -2449 5799 -2361 5812
rect -2449 5725 -2420 5799
rect -2374 5725 -2361 5799
rect -2449 5712 -2361 5725
rect -1990 5799 -1902 5812
rect -1990 5725 -1977 5799
rect -1931 5725 -1902 5799
rect -1990 5712 -1902 5725
rect -1846 5799 -1742 5812
rect -1846 5725 -1817 5799
rect -1771 5725 -1742 5799
rect -1846 5712 -1742 5725
rect -1686 5799 -1598 5812
rect -1686 5725 -1657 5799
rect -1611 5725 -1598 5799
rect -1686 5712 -1598 5725
rect -1179 5799 -1091 5812
rect -1179 5725 -1166 5799
rect -1120 5725 -1091 5799
rect -1179 5712 -1091 5725
rect -1035 5799 -931 5812
rect -1035 5725 -1006 5799
rect -960 5725 -931 5799
rect -1035 5712 -931 5725
rect -875 5799 -787 5812
rect -875 5725 -846 5799
rect -800 5725 -787 5799
rect -875 5712 -787 5725
rect 229 5743 317 5756
rect 229 5649 242 5743
rect 288 5649 317 5743
rect 229 5636 317 5649
rect 417 5743 521 5756
rect 417 5649 446 5743
rect 492 5649 521 5743
rect 417 5636 521 5649
rect 621 5743 725 5756
rect 621 5649 650 5743
rect 696 5649 725 5743
rect 621 5636 725 5649
rect 825 5743 929 5756
rect 825 5649 854 5743
rect 900 5649 929 5743
rect 825 5636 929 5649
rect 1029 5743 1133 5756
rect 1029 5649 1058 5743
rect 1104 5649 1133 5743
rect 1029 5636 1133 5649
rect 1233 5743 1337 5756
rect 1233 5649 1262 5743
rect 1308 5649 1337 5743
rect 1233 5636 1337 5649
rect 1437 5743 1541 5756
rect 1437 5649 1466 5743
rect 1512 5649 1541 5743
rect 1437 5636 1541 5649
rect 1641 5743 1745 5756
rect 1641 5649 1670 5743
rect 1716 5649 1745 5743
rect 1641 5636 1745 5649
rect 1845 5743 1949 5756
rect 1845 5649 1874 5743
rect 1920 5649 1949 5743
rect 1845 5636 1949 5649
rect 2049 5743 2153 5756
rect 2049 5649 2078 5743
rect 2124 5649 2153 5743
rect 2049 5636 2153 5649
rect 2253 5743 2357 5756
rect 2253 5649 2282 5743
rect 2328 5649 2357 5743
rect 2253 5636 2357 5649
rect 2457 5743 2561 5756
rect 2457 5649 2486 5743
rect 2532 5649 2561 5743
rect 2457 5636 2561 5649
rect 2661 5743 2765 5756
rect 2661 5649 2690 5743
rect 2736 5649 2765 5743
rect 2661 5636 2765 5649
rect 2865 5743 2969 5756
rect 2865 5649 2894 5743
rect 2940 5649 2969 5743
rect 2865 5636 2969 5649
rect 3069 5743 3173 5756
rect 3069 5649 3098 5743
rect 3144 5649 3173 5743
rect 3069 5636 3173 5649
rect 3273 5743 3377 5756
rect 3273 5649 3302 5743
rect 3348 5649 3377 5743
rect 3273 5636 3377 5649
rect 3477 5743 3565 5756
rect 3477 5649 3506 5743
rect 3552 5649 3565 5743
rect 3477 5636 3565 5649
rect 229 5351 317 5364
rect 229 5257 242 5351
rect 288 5257 317 5351
rect 229 5244 317 5257
rect 417 5351 521 5364
rect 417 5257 446 5351
rect 492 5257 521 5351
rect 417 5244 521 5257
rect 621 5351 725 5364
rect 621 5257 650 5351
rect 696 5257 725 5351
rect 621 5244 725 5257
rect 825 5351 929 5364
rect 825 5257 854 5351
rect 900 5257 929 5351
rect 825 5244 929 5257
rect 1029 5351 1133 5364
rect 1029 5257 1058 5351
rect 1104 5257 1133 5351
rect 1029 5244 1133 5257
rect 1233 5351 1337 5364
rect 1233 5257 1262 5351
rect 1308 5257 1337 5351
rect 1233 5244 1337 5257
rect 1437 5351 1541 5364
rect 1437 5257 1466 5351
rect 1512 5257 1541 5351
rect 1437 5244 1541 5257
rect 1641 5351 1745 5364
rect 1641 5257 1670 5351
rect 1716 5257 1745 5351
rect 1641 5244 1745 5257
rect 1845 5351 1949 5364
rect 1845 5257 1874 5351
rect 1920 5257 1949 5351
rect 1845 5244 1949 5257
rect 2049 5351 2153 5364
rect 2049 5257 2078 5351
rect 2124 5257 2153 5351
rect 2049 5244 2153 5257
rect 2253 5351 2357 5364
rect 2253 5257 2282 5351
rect 2328 5257 2357 5351
rect 2253 5244 2357 5257
rect 2457 5351 2561 5364
rect 2457 5257 2486 5351
rect 2532 5257 2561 5351
rect 2457 5244 2561 5257
rect 2661 5351 2765 5364
rect 2661 5257 2690 5351
rect 2736 5257 2765 5351
rect 2661 5244 2765 5257
rect 2865 5351 2969 5364
rect 2865 5257 2894 5351
rect 2940 5257 2969 5351
rect 2865 5244 2969 5257
rect 3069 5351 3173 5364
rect 3069 5257 3098 5351
rect 3144 5257 3173 5351
rect 3069 5244 3173 5257
rect 3273 5351 3377 5364
rect 3273 5257 3302 5351
rect 3348 5257 3377 5351
rect 3273 5244 3377 5257
rect 3477 5351 3565 5364
rect 3477 5257 3506 5351
rect 3552 5257 3565 5351
rect 3477 5244 3565 5257
rect -2753 4828 -2665 4841
rect -2753 4754 -2740 4828
rect -2694 4754 -2665 4828
rect -2753 4741 -2665 4754
rect -2609 4828 -2505 4841
rect -2609 4754 -2580 4828
rect -2534 4754 -2505 4828
rect -2609 4741 -2505 4754
rect -2449 4828 -2361 4841
rect -2449 4754 -2420 4828
rect -2374 4754 -2361 4828
rect -2449 4741 -2361 4754
rect -1990 4828 -1902 4841
rect -1990 4754 -1977 4828
rect -1931 4754 -1902 4828
rect -1990 4741 -1902 4754
rect -1846 4828 -1742 4841
rect -1846 4754 -1817 4828
rect -1771 4754 -1742 4828
rect -1846 4741 -1742 4754
rect -1686 4828 -1598 4841
rect -1686 4754 -1657 4828
rect -1611 4754 -1598 4828
rect -1686 4741 -1598 4754
rect -1179 4828 -1091 4841
rect -1179 4754 -1166 4828
rect -1120 4754 -1091 4828
rect -1179 4741 -1091 4754
rect -1035 4828 -931 4841
rect -1035 4754 -1006 4828
rect -960 4754 -931 4828
rect -1035 4741 -931 4754
rect -875 4828 -787 4841
rect -875 4754 -846 4828
rect -800 4754 -787 4828
rect -875 4741 -787 4754
rect 229 4946 317 4959
rect 229 4852 242 4946
rect 288 4852 317 4946
rect 229 4839 317 4852
rect 417 4946 521 4959
rect 417 4852 446 4946
rect 492 4852 521 4946
rect 417 4839 521 4852
rect 621 4946 725 4959
rect 621 4852 650 4946
rect 696 4852 725 4946
rect 621 4839 725 4852
rect 825 4946 929 4959
rect 825 4852 854 4946
rect 900 4852 929 4946
rect 825 4839 929 4852
rect 1029 4946 1133 4959
rect 1029 4852 1058 4946
rect 1104 4852 1133 4946
rect 1029 4839 1133 4852
rect 1233 4946 1337 4959
rect 1233 4852 1262 4946
rect 1308 4852 1337 4946
rect 1233 4839 1337 4852
rect 1437 4946 1541 4959
rect 1437 4852 1466 4946
rect 1512 4852 1541 4946
rect 1437 4839 1541 4852
rect 1641 4946 1745 4959
rect 1641 4852 1670 4946
rect 1716 4852 1745 4946
rect 1641 4839 1745 4852
rect 1845 4946 1949 4959
rect 1845 4852 1874 4946
rect 1920 4852 1949 4946
rect 1845 4839 1949 4852
rect 2049 4946 2153 4959
rect 2049 4852 2078 4946
rect 2124 4852 2153 4946
rect 2049 4839 2153 4852
rect 2253 4946 2357 4959
rect 2253 4852 2282 4946
rect 2328 4852 2357 4946
rect 2253 4839 2357 4852
rect 2457 4946 2561 4959
rect 2457 4852 2486 4946
rect 2532 4852 2561 4946
rect 2457 4839 2561 4852
rect 2661 4946 2765 4959
rect 2661 4852 2690 4946
rect 2736 4852 2765 4946
rect 2661 4839 2765 4852
rect 2865 4946 2969 4959
rect 2865 4852 2894 4946
rect 2940 4852 2969 4946
rect 2865 4839 2969 4852
rect 3069 4946 3173 4959
rect 3069 4852 3098 4946
rect 3144 4852 3173 4946
rect 3069 4839 3173 4852
rect 3273 4946 3377 4959
rect 3273 4852 3302 4946
rect 3348 4852 3377 4946
rect 3273 4839 3377 4852
rect 3477 4946 3565 4959
rect 3477 4852 3506 4946
rect 3552 4852 3565 4946
rect 3477 4839 3565 4852
rect 229 4554 317 4567
rect 229 4460 242 4554
rect 288 4460 317 4554
rect 229 4447 317 4460
rect 417 4554 521 4567
rect 417 4460 446 4554
rect 492 4460 521 4554
rect 417 4447 521 4460
rect 621 4554 725 4567
rect 621 4460 650 4554
rect 696 4460 725 4554
rect 621 4447 725 4460
rect 825 4554 929 4567
rect 825 4460 854 4554
rect 900 4460 929 4554
rect 825 4447 929 4460
rect 1029 4554 1133 4567
rect 1029 4460 1058 4554
rect 1104 4460 1133 4554
rect 1029 4447 1133 4460
rect 1233 4554 1337 4567
rect 1233 4460 1262 4554
rect 1308 4460 1337 4554
rect 1233 4447 1337 4460
rect 1437 4554 1541 4567
rect 1437 4460 1466 4554
rect 1512 4460 1541 4554
rect 1437 4447 1541 4460
rect 1641 4554 1745 4567
rect 1641 4460 1670 4554
rect 1716 4460 1745 4554
rect 1641 4447 1745 4460
rect 1845 4554 1949 4567
rect 1845 4460 1874 4554
rect 1920 4460 1949 4554
rect 1845 4447 1949 4460
rect 2049 4554 2153 4567
rect 2049 4460 2078 4554
rect 2124 4460 2153 4554
rect 2049 4447 2153 4460
rect 2253 4554 2357 4567
rect 2253 4460 2282 4554
rect 2328 4460 2357 4554
rect 2253 4447 2357 4460
rect 2457 4554 2561 4567
rect 2457 4460 2486 4554
rect 2532 4460 2561 4554
rect 2457 4447 2561 4460
rect 2661 4554 2765 4567
rect 2661 4460 2690 4554
rect 2736 4460 2765 4554
rect 2661 4447 2765 4460
rect 2865 4554 2969 4567
rect 2865 4460 2894 4554
rect 2940 4460 2969 4554
rect 2865 4447 2969 4460
rect 3069 4554 3173 4567
rect 3069 4460 3098 4554
rect 3144 4460 3173 4554
rect 3069 4447 3173 4460
rect 3273 4554 3377 4567
rect 3273 4460 3302 4554
rect 3348 4460 3377 4554
rect 3273 4447 3377 4460
rect 3477 4554 3565 4567
rect 3477 4460 3506 4554
rect 3552 4460 3565 4554
rect 3477 4447 3565 4460
rect -2753 3853 -2665 3866
rect -2753 3779 -2740 3853
rect -2694 3779 -2665 3853
rect -2753 3766 -2665 3779
rect -2609 3853 -2505 3866
rect -2609 3779 -2580 3853
rect -2534 3779 -2505 3853
rect -2609 3766 -2505 3779
rect -2449 3853 -2361 3866
rect 229 4149 317 4162
rect 229 4055 242 4149
rect 288 4055 317 4149
rect 229 4042 317 4055
rect 417 4149 521 4162
rect 417 4055 446 4149
rect 492 4055 521 4149
rect 417 4042 521 4055
rect 621 4149 725 4162
rect 621 4055 650 4149
rect 696 4055 725 4149
rect 621 4042 725 4055
rect 825 4149 929 4162
rect 825 4055 854 4149
rect 900 4055 929 4149
rect 825 4042 929 4055
rect 1029 4149 1133 4162
rect 1029 4055 1058 4149
rect 1104 4055 1133 4149
rect 1029 4042 1133 4055
rect 1233 4149 1337 4162
rect 1233 4055 1262 4149
rect 1308 4055 1337 4149
rect 1233 4042 1337 4055
rect 1437 4149 1541 4162
rect 1437 4055 1466 4149
rect 1512 4055 1541 4149
rect 1437 4042 1541 4055
rect 1641 4149 1745 4162
rect 1641 4055 1670 4149
rect 1716 4055 1745 4149
rect 1641 4042 1745 4055
rect 1845 4149 1949 4162
rect 1845 4055 1874 4149
rect 1920 4055 1949 4149
rect 1845 4042 1949 4055
rect 2049 4149 2153 4162
rect 2049 4055 2078 4149
rect 2124 4055 2153 4149
rect 2049 4042 2153 4055
rect 2253 4149 2357 4162
rect 2253 4055 2282 4149
rect 2328 4055 2357 4149
rect 2253 4042 2357 4055
rect 2457 4149 2561 4162
rect 2457 4055 2486 4149
rect 2532 4055 2561 4149
rect 2457 4042 2561 4055
rect 2661 4149 2765 4162
rect 2661 4055 2690 4149
rect 2736 4055 2765 4149
rect 2661 4042 2765 4055
rect 2865 4149 2969 4162
rect 2865 4055 2894 4149
rect 2940 4055 2969 4149
rect 2865 4042 2969 4055
rect 3069 4149 3173 4162
rect 3069 4055 3098 4149
rect 3144 4055 3173 4149
rect 3069 4042 3173 4055
rect 3273 4149 3377 4162
rect 3273 4055 3302 4149
rect 3348 4055 3377 4149
rect 3273 4042 3377 4055
rect 3477 4149 3565 4162
rect 3477 4055 3506 4149
rect 3552 4055 3565 4149
rect 3477 4042 3565 4055
rect -2449 3779 -2420 3853
rect -2374 3779 -2361 3853
rect -2449 3766 -2361 3779
rect -1990 3852 -1902 3865
rect -1990 3778 -1977 3852
rect -1931 3778 -1902 3852
rect -1990 3765 -1902 3778
rect -1846 3852 -1742 3865
rect -1846 3778 -1817 3852
rect -1771 3778 -1742 3852
rect -1846 3765 -1742 3778
rect -1686 3852 -1598 3865
rect -1686 3778 -1657 3852
rect -1611 3778 -1598 3852
rect -1686 3765 -1598 3778
rect -1179 3852 -1091 3865
rect -1179 3778 -1166 3852
rect -1120 3778 -1091 3852
rect -1179 3765 -1091 3778
rect -1035 3852 -931 3865
rect -1035 3778 -1006 3852
rect -960 3778 -931 3852
rect -1035 3765 -931 3778
rect -875 3852 -787 3865
rect -875 3778 -846 3852
rect -800 3778 -787 3852
rect -875 3765 -787 3778
rect -2815 3057 -2727 3070
rect -2815 2843 -2802 3057
rect -2756 2843 -2727 3057
rect -2815 2830 -2727 2843
rect -2627 3057 -2523 3070
rect -2627 2843 -2598 3057
rect -2552 2843 -2523 3057
rect -2627 2830 -2523 2843
rect -2423 3057 -2319 3070
rect -2423 2843 -2394 3057
rect -2348 2843 -2319 3057
rect -2423 2830 -2319 2843
rect -2219 3057 -2115 3070
rect -2219 2843 -2190 3057
rect -2144 2843 -2115 3057
rect -2219 2830 -2115 2843
rect -2015 3057 -1911 3070
rect -2015 2843 -1986 3057
rect -1940 2843 -1911 3057
rect -2015 2830 -1911 2843
rect -1811 3057 -1707 3070
rect -1811 2843 -1782 3057
rect -1736 2843 -1707 3057
rect -1811 2830 -1707 2843
rect -1607 3057 -1503 3070
rect -1607 2843 -1578 3057
rect -1532 2843 -1503 3057
rect -1607 2830 -1503 2843
rect -1403 3057 -1299 3070
rect -1403 2843 -1374 3057
rect -1328 2843 -1299 3057
rect -1403 2830 -1299 2843
rect -1199 3057 -1095 3070
rect -1199 2843 -1170 3057
rect -1124 2843 -1095 3057
rect -1199 2830 -1095 2843
rect -995 3057 -891 3070
rect -995 2843 -966 3057
rect -920 2843 -891 3057
rect -995 2830 -891 2843
rect -791 3057 -687 3070
rect -791 2843 -762 3057
rect -716 2843 -687 3057
rect -791 2830 -687 2843
rect -587 3057 -483 3070
rect -587 2843 -558 3057
rect -512 2843 -483 3057
rect -587 2830 -483 2843
rect -383 3057 -279 3070
rect -383 2843 -354 3057
rect -308 2843 -279 3057
rect -383 2830 -279 2843
rect -179 3057 -75 3070
rect -179 2843 -150 3057
rect -104 2843 -75 3057
rect -179 2830 -75 2843
rect 25 3057 129 3070
rect 25 2843 54 3057
rect 100 2843 129 3057
rect 25 2830 129 2843
rect 229 3057 333 3070
rect 229 2843 258 3057
rect 304 2843 333 3057
rect 229 2830 333 2843
rect 433 3057 537 3070
rect 433 2843 462 3057
rect 508 2843 537 3057
rect 433 2830 537 2843
rect 637 3057 741 3070
rect 637 2843 666 3057
rect 712 2843 741 3057
rect 637 2830 741 2843
rect 841 3057 945 3070
rect 841 2843 870 3057
rect 916 2843 945 3057
rect 841 2830 945 2843
rect 1045 3057 1149 3070
rect 1045 2843 1074 3057
rect 1120 2843 1149 3057
rect 1045 2830 1149 2843
rect 1249 3057 1353 3070
rect 1249 2843 1278 3057
rect 1324 2843 1353 3057
rect 1249 2830 1353 2843
rect 1453 3057 1557 3070
rect 1453 2843 1482 3057
rect 1528 2843 1557 3057
rect 1453 2830 1557 2843
rect 1657 3057 1761 3070
rect 1657 2843 1686 3057
rect 1732 2843 1761 3057
rect 1657 2830 1761 2843
rect 1861 3057 1965 3070
rect 1861 2843 1890 3057
rect 1936 2843 1965 3057
rect 1861 2830 1965 2843
rect 2065 3057 2169 3070
rect 2065 2843 2094 3057
rect 2140 2843 2169 3057
rect 2065 2830 2169 2843
rect 2269 3057 2373 3070
rect 2269 2843 2298 3057
rect 2344 2843 2373 3057
rect 2269 2830 2373 2843
rect 2473 3057 2577 3070
rect 2473 2843 2502 3057
rect 2548 2843 2577 3057
rect 2473 2830 2577 2843
rect 2677 3057 2781 3070
rect 2677 2843 2706 3057
rect 2752 2843 2781 3057
rect 2677 2830 2781 2843
rect 2881 3057 2985 3070
rect 2881 2843 2910 3057
rect 2956 2843 2985 3057
rect 2881 2830 2985 2843
rect 3085 3057 3189 3070
rect 3085 2843 3114 3057
rect 3160 2843 3189 3057
rect 3085 2830 3189 2843
rect 3289 3057 3393 3070
rect 3289 2843 3318 3057
rect 3364 2843 3393 3057
rect 3289 2830 3393 2843
rect 3493 3057 3597 3070
rect 3493 2843 3522 3057
rect 3568 2843 3597 3057
rect 3493 2830 3597 2843
rect 3697 3057 3785 3070
rect 3697 2843 3726 3057
rect 3772 2843 3785 3057
rect 3697 2830 3785 2843
rect -2815 2566 -2727 2579
rect -2815 2352 -2802 2566
rect -2756 2352 -2727 2566
rect -2815 2339 -2727 2352
rect -2627 2566 -2523 2579
rect -2627 2352 -2598 2566
rect -2552 2352 -2523 2566
rect -2627 2339 -2523 2352
rect -2423 2566 -2319 2579
rect -2423 2352 -2394 2566
rect -2348 2352 -2319 2566
rect -2423 2339 -2319 2352
rect -2219 2566 -2115 2579
rect -2219 2352 -2190 2566
rect -2144 2352 -2115 2566
rect -2219 2339 -2115 2352
rect -2015 2566 -1911 2579
rect -2015 2352 -1986 2566
rect -1940 2352 -1911 2566
rect -2015 2339 -1911 2352
rect -1811 2566 -1707 2579
rect -1811 2352 -1782 2566
rect -1736 2352 -1707 2566
rect -1811 2339 -1707 2352
rect -1607 2566 -1503 2579
rect -1607 2352 -1578 2566
rect -1532 2352 -1503 2566
rect -1607 2339 -1503 2352
rect -1403 2566 -1299 2579
rect -1403 2352 -1374 2566
rect -1328 2352 -1299 2566
rect -1403 2339 -1299 2352
rect -1199 2566 -1095 2579
rect -1199 2352 -1170 2566
rect -1124 2352 -1095 2566
rect -1199 2339 -1095 2352
rect -995 2566 -891 2579
rect -995 2352 -966 2566
rect -920 2352 -891 2566
rect -995 2339 -891 2352
rect -791 2566 -687 2579
rect -791 2352 -762 2566
rect -716 2352 -687 2566
rect -791 2339 -687 2352
rect -587 2566 -483 2579
rect -587 2352 -558 2566
rect -512 2352 -483 2566
rect -587 2339 -483 2352
rect -383 2566 -279 2579
rect -383 2352 -354 2566
rect -308 2352 -279 2566
rect -383 2339 -279 2352
rect -179 2566 -75 2579
rect -179 2352 -150 2566
rect -104 2352 -75 2566
rect -179 2339 -75 2352
rect 25 2566 129 2579
rect 25 2352 54 2566
rect 100 2352 129 2566
rect 25 2339 129 2352
rect 229 2566 333 2579
rect 229 2352 258 2566
rect 304 2352 333 2566
rect 229 2339 333 2352
rect 433 2566 537 2579
rect 433 2352 462 2566
rect 508 2352 537 2566
rect 433 2339 537 2352
rect 637 2566 741 2579
rect 637 2352 666 2566
rect 712 2352 741 2566
rect 637 2339 741 2352
rect 841 2566 945 2579
rect 841 2352 870 2566
rect 916 2352 945 2566
rect 841 2339 945 2352
rect 1045 2566 1149 2579
rect 1045 2352 1074 2566
rect 1120 2352 1149 2566
rect 1045 2339 1149 2352
rect 1249 2566 1353 2579
rect 1249 2352 1278 2566
rect 1324 2352 1353 2566
rect 1249 2339 1353 2352
rect 1453 2566 1557 2579
rect 1453 2352 1482 2566
rect 1528 2352 1557 2566
rect 1453 2339 1557 2352
rect 1657 2566 1761 2579
rect 1657 2352 1686 2566
rect 1732 2352 1761 2566
rect 1657 2339 1761 2352
rect 1861 2566 1965 2579
rect 1861 2352 1890 2566
rect 1936 2352 1965 2566
rect 1861 2339 1965 2352
rect 2065 2566 2169 2579
rect 2065 2352 2094 2566
rect 2140 2352 2169 2566
rect 2065 2339 2169 2352
rect 2269 2566 2373 2579
rect 2269 2352 2298 2566
rect 2344 2352 2373 2566
rect 2269 2339 2373 2352
rect 2473 2566 2577 2579
rect 2473 2352 2502 2566
rect 2548 2352 2577 2566
rect 2473 2339 2577 2352
rect 2677 2566 2781 2579
rect 2677 2352 2706 2566
rect 2752 2352 2781 2566
rect 2677 2339 2781 2352
rect 2881 2566 2985 2579
rect 2881 2352 2910 2566
rect 2956 2352 2985 2566
rect 2881 2339 2985 2352
rect 3085 2566 3189 2579
rect 3085 2352 3114 2566
rect 3160 2352 3189 2566
rect 3085 2339 3189 2352
rect 3289 2566 3393 2579
rect 3289 2352 3318 2566
rect 3364 2352 3393 2566
rect 3289 2339 3393 2352
rect 3493 2566 3597 2579
rect 3493 2352 3522 2566
rect 3568 2352 3597 2566
rect 3493 2339 3597 2352
rect 3697 2566 3785 2579
rect 3697 2352 3726 2566
rect 3772 2352 3785 2566
rect 3697 2339 3785 2352
<< pdiff >>
rect -2753 6169 -2665 6182
rect -2753 6095 -2740 6169
rect -2694 6095 -2665 6169
rect -2753 6082 -2665 6095
rect -2609 6169 -2505 6182
rect -2609 6095 -2580 6169
rect -2534 6095 -2505 6169
rect -2609 6082 -2505 6095
rect -2449 6169 -2361 6182
rect -2449 6095 -2420 6169
rect -2374 6095 -2361 6169
rect -2449 6082 -2361 6095
rect -1990 6169 -1902 6182
rect -1990 6095 -1977 6169
rect -1931 6095 -1902 6169
rect -1990 6082 -1902 6095
rect -1846 6169 -1742 6182
rect -1846 6095 -1817 6169
rect -1771 6095 -1742 6169
rect -1846 6082 -1742 6095
rect -1686 6169 -1598 6182
rect -1686 6095 -1657 6169
rect -1611 6095 -1598 6169
rect -1686 6082 -1598 6095
rect -1179 6169 -1091 6182
rect -1179 6095 -1166 6169
rect -1120 6095 -1091 6169
rect -1179 6082 -1091 6095
rect -1035 6169 -931 6182
rect -1035 6095 -1006 6169
rect -960 6095 -931 6169
rect -1035 6082 -931 6095
rect -875 6169 -787 6182
rect -875 6095 -846 6169
rect -800 6095 -787 6169
rect -875 6082 -787 6095
rect -2753 5198 -2665 5211
rect -2753 5124 -2740 5198
rect -2694 5124 -2665 5198
rect -2753 5111 -2665 5124
rect -2609 5198 -2505 5211
rect -2609 5124 -2580 5198
rect -2534 5124 -2505 5198
rect -2609 5111 -2505 5124
rect -2449 5198 -2361 5211
rect -2449 5124 -2420 5198
rect -2374 5124 -2361 5198
rect -2449 5111 -2361 5124
rect -1990 5198 -1902 5211
rect -1990 5124 -1977 5198
rect -1931 5124 -1902 5198
rect -1990 5111 -1902 5124
rect -1846 5198 -1742 5211
rect -1846 5124 -1817 5198
rect -1771 5124 -1742 5198
rect -1846 5111 -1742 5124
rect -1686 5198 -1598 5211
rect -1686 5124 -1657 5198
rect -1611 5124 -1598 5198
rect -1686 5111 -1598 5124
rect -1179 5198 -1091 5211
rect -1179 5124 -1166 5198
rect -1120 5124 -1091 5198
rect -1179 5111 -1091 5124
rect -1035 5198 -931 5211
rect -1035 5124 -1006 5198
rect -960 5124 -931 5198
rect -1035 5111 -931 5124
rect -875 5198 -787 5211
rect -875 5124 -846 5198
rect -800 5124 -787 5198
rect -875 5111 -787 5124
rect -2753 4223 -2665 4236
rect -2753 4149 -2740 4223
rect -2694 4149 -2665 4223
rect -2753 4136 -2665 4149
rect -2609 4223 -2505 4236
rect -2609 4149 -2580 4223
rect -2534 4149 -2505 4223
rect -2609 4136 -2505 4149
rect -2449 4223 -2361 4236
rect -2449 4149 -2420 4223
rect -2374 4149 -2361 4223
rect -2449 4136 -2361 4149
rect -1990 4222 -1902 4235
rect -1990 4148 -1977 4222
rect -1931 4148 -1902 4222
rect -1990 4135 -1902 4148
rect -1846 4222 -1742 4235
rect -1846 4148 -1817 4222
rect -1771 4148 -1742 4222
rect -1846 4135 -1742 4148
rect -1686 4222 -1598 4235
rect -1686 4148 -1657 4222
rect -1611 4148 -1598 4222
rect -1686 4135 -1598 4148
rect -1179 4222 -1091 4235
rect -1179 4148 -1166 4222
rect -1120 4148 -1091 4222
rect -1179 4135 -1091 4148
rect -1035 4222 -931 4235
rect -1035 4148 -1006 4222
rect -960 4148 -931 4222
rect -1035 4135 -931 4148
rect -875 4222 -787 4235
rect -875 4148 -846 4222
rect -800 4148 -787 4222
rect -875 4135 -787 4148
<< ndiffc >>
rect 242 6851 288 6945
rect 446 6851 492 6945
rect 650 6851 696 6945
rect 854 6851 900 6945
rect 1058 6851 1104 6945
rect 1262 6851 1308 6945
rect 1466 6851 1512 6945
rect 1670 6851 1716 6945
rect 1874 6851 1920 6945
rect 2078 6851 2124 6945
rect 2282 6851 2328 6945
rect 2486 6851 2532 6945
rect 2690 6851 2736 6945
rect 2894 6851 2940 6945
rect 3098 6851 3144 6945
rect 3302 6851 3348 6945
rect 3506 6851 3552 6945
rect 242 6446 288 6540
rect 446 6446 492 6540
rect 650 6446 696 6540
rect 854 6446 900 6540
rect 1058 6446 1104 6540
rect 1262 6446 1308 6540
rect 1466 6446 1512 6540
rect 1670 6446 1716 6540
rect 1874 6446 1920 6540
rect 2078 6446 2124 6540
rect 2282 6446 2328 6540
rect 2486 6446 2532 6540
rect 2690 6446 2736 6540
rect 2894 6446 2940 6540
rect 3098 6446 3144 6540
rect 3302 6446 3348 6540
rect 3506 6446 3552 6540
rect 242 6054 288 6148
rect 446 6054 492 6148
rect 650 6054 696 6148
rect 854 6054 900 6148
rect 1058 6054 1104 6148
rect 1262 6054 1308 6148
rect 1466 6054 1512 6148
rect 1670 6054 1716 6148
rect 1874 6054 1920 6148
rect 2078 6054 2124 6148
rect 2282 6054 2328 6148
rect 2486 6054 2532 6148
rect 2690 6054 2736 6148
rect 2894 6054 2940 6148
rect 3098 6054 3144 6148
rect 3302 6054 3348 6148
rect 3506 6054 3552 6148
rect -2740 5725 -2694 5799
rect -2580 5725 -2534 5799
rect -2420 5725 -2374 5799
rect -1977 5725 -1931 5799
rect -1817 5725 -1771 5799
rect -1657 5725 -1611 5799
rect -1166 5725 -1120 5799
rect -1006 5725 -960 5799
rect -846 5725 -800 5799
rect 242 5649 288 5743
rect 446 5649 492 5743
rect 650 5649 696 5743
rect 854 5649 900 5743
rect 1058 5649 1104 5743
rect 1262 5649 1308 5743
rect 1466 5649 1512 5743
rect 1670 5649 1716 5743
rect 1874 5649 1920 5743
rect 2078 5649 2124 5743
rect 2282 5649 2328 5743
rect 2486 5649 2532 5743
rect 2690 5649 2736 5743
rect 2894 5649 2940 5743
rect 3098 5649 3144 5743
rect 3302 5649 3348 5743
rect 3506 5649 3552 5743
rect 242 5257 288 5351
rect 446 5257 492 5351
rect 650 5257 696 5351
rect 854 5257 900 5351
rect 1058 5257 1104 5351
rect 1262 5257 1308 5351
rect 1466 5257 1512 5351
rect 1670 5257 1716 5351
rect 1874 5257 1920 5351
rect 2078 5257 2124 5351
rect 2282 5257 2328 5351
rect 2486 5257 2532 5351
rect 2690 5257 2736 5351
rect 2894 5257 2940 5351
rect 3098 5257 3144 5351
rect 3302 5257 3348 5351
rect 3506 5257 3552 5351
rect -2740 4754 -2694 4828
rect -2580 4754 -2534 4828
rect -2420 4754 -2374 4828
rect -1977 4754 -1931 4828
rect -1817 4754 -1771 4828
rect -1657 4754 -1611 4828
rect -1166 4754 -1120 4828
rect -1006 4754 -960 4828
rect -846 4754 -800 4828
rect 242 4852 288 4946
rect 446 4852 492 4946
rect 650 4852 696 4946
rect 854 4852 900 4946
rect 1058 4852 1104 4946
rect 1262 4852 1308 4946
rect 1466 4852 1512 4946
rect 1670 4852 1716 4946
rect 1874 4852 1920 4946
rect 2078 4852 2124 4946
rect 2282 4852 2328 4946
rect 2486 4852 2532 4946
rect 2690 4852 2736 4946
rect 2894 4852 2940 4946
rect 3098 4852 3144 4946
rect 3302 4852 3348 4946
rect 3506 4852 3552 4946
rect 242 4460 288 4554
rect 446 4460 492 4554
rect 650 4460 696 4554
rect 854 4460 900 4554
rect 1058 4460 1104 4554
rect 1262 4460 1308 4554
rect 1466 4460 1512 4554
rect 1670 4460 1716 4554
rect 1874 4460 1920 4554
rect 2078 4460 2124 4554
rect 2282 4460 2328 4554
rect 2486 4460 2532 4554
rect 2690 4460 2736 4554
rect 2894 4460 2940 4554
rect 3098 4460 3144 4554
rect 3302 4460 3348 4554
rect 3506 4460 3552 4554
rect -2740 3779 -2694 3853
rect -2580 3779 -2534 3853
rect 242 4055 288 4149
rect 446 4055 492 4149
rect 650 4055 696 4149
rect 854 4055 900 4149
rect 1058 4055 1104 4149
rect 1262 4055 1308 4149
rect 1466 4055 1512 4149
rect 1670 4055 1716 4149
rect 1874 4055 1920 4149
rect 2078 4055 2124 4149
rect 2282 4055 2328 4149
rect 2486 4055 2532 4149
rect 2690 4055 2736 4149
rect 2894 4055 2940 4149
rect 3098 4055 3144 4149
rect 3302 4055 3348 4149
rect 3506 4055 3552 4149
rect -2420 3779 -2374 3853
rect -1977 3778 -1931 3852
rect -1817 3778 -1771 3852
rect -1657 3778 -1611 3852
rect -1166 3778 -1120 3852
rect -1006 3778 -960 3852
rect -846 3778 -800 3852
rect -2802 2843 -2756 3057
rect -2598 2843 -2552 3057
rect -2394 2843 -2348 3057
rect -2190 2843 -2144 3057
rect -1986 2843 -1940 3057
rect -1782 2843 -1736 3057
rect -1578 2843 -1532 3057
rect -1374 2843 -1328 3057
rect -1170 2843 -1124 3057
rect -966 2843 -920 3057
rect -762 2843 -716 3057
rect -558 2843 -512 3057
rect -354 2843 -308 3057
rect -150 2843 -104 3057
rect 54 2843 100 3057
rect 258 2843 304 3057
rect 462 2843 508 3057
rect 666 2843 712 3057
rect 870 2843 916 3057
rect 1074 2843 1120 3057
rect 1278 2843 1324 3057
rect 1482 2843 1528 3057
rect 1686 2843 1732 3057
rect 1890 2843 1936 3057
rect 2094 2843 2140 3057
rect 2298 2843 2344 3057
rect 2502 2843 2548 3057
rect 2706 2843 2752 3057
rect 2910 2843 2956 3057
rect 3114 2843 3160 3057
rect 3318 2843 3364 3057
rect 3522 2843 3568 3057
rect 3726 2843 3772 3057
rect -2802 2352 -2756 2566
rect -2598 2352 -2552 2566
rect -2394 2352 -2348 2566
rect -2190 2352 -2144 2566
rect -1986 2352 -1940 2566
rect -1782 2352 -1736 2566
rect -1578 2352 -1532 2566
rect -1374 2352 -1328 2566
rect -1170 2352 -1124 2566
rect -966 2352 -920 2566
rect -762 2352 -716 2566
rect -558 2352 -512 2566
rect -354 2352 -308 2566
rect -150 2352 -104 2566
rect 54 2352 100 2566
rect 258 2352 304 2566
rect 462 2352 508 2566
rect 666 2352 712 2566
rect 870 2352 916 2566
rect 1074 2352 1120 2566
rect 1278 2352 1324 2566
rect 1482 2352 1528 2566
rect 1686 2352 1732 2566
rect 1890 2352 1936 2566
rect 2094 2352 2140 2566
rect 2298 2352 2344 2566
rect 2502 2352 2548 2566
rect 2706 2352 2752 2566
rect 2910 2352 2956 2566
rect 3114 2352 3160 2566
rect 3318 2352 3364 2566
rect 3522 2352 3568 2566
rect 3726 2352 3772 2566
<< pdiffc >>
rect -2740 6095 -2694 6169
rect -2580 6095 -2534 6169
rect -2420 6095 -2374 6169
rect -1977 6095 -1931 6169
rect -1817 6095 -1771 6169
rect -1657 6095 -1611 6169
rect -1166 6095 -1120 6169
rect -1006 6095 -960 6169
rect -846 6095 -800 6169
rect -2740 5124 -2694 5198
rect -2580 5124 -2534 5198
rect -2420 5124 -2374 5198
rect -1977 5124 -1931 5198
rect -1817 5124 -1771 5198
rect -1657 5124 -1611 5198
rect -1166 5124 -1120 5198
rect -1006 5124 -960 5198
rect -846 5124 -800 5198
rect -2740 4149 -2694 4223
rect -2580 4149 -2534 4223
rect -2420 4149 -2374 4223
rect -1977 4148 -1931 4222
rect -1817 4148 -1771 4222
rect -1657 4148 -1611 4222
rect -1166 4148 -1120 4222
rect -1006 4148 -960 4222
rect -846 4148 -800 4222
<< psubdiff >>
rect -422 7360 4308 7377
rect -422 7270 -407 7360
rect -307 7270 -207 7360
rect -107 7270 -7 7360
rect 93 7270 193 7360
rect 293 7270 393 7360
rect 493 7270 593 7360
rect 693 7270 793 7360
rect 893 7270 993 7360
rect 1093 7270 1193 7360
rect 1293 7270 1393 7360
rect 1493 7270 1593 7360
rect 1693 7270 1793 7360
rect 1893 7270 1993 7360
rect 2093 7270 2193 7360
rect 2293 7270 2393 7360
rect 2493 7270 2593 7360
rect 2693 7270 2793 7360
rect 2893 7270 2993 7360
rect 3093 7270 3193 7360
rect 3293 7270 3393 7360
rect 3493 7270 3593 7360
rect 3693 7270 3793 7360
rect 3893 7270 3993 7360
rect 4093 7270 4193 7360
rect 4293 7270 4308 7360
rect -422 7257 4308 7270
rect -422 7160 -292 7257
rect -422 7070 -407 7160
rect -307 7070 -292 7160
rect 4178 7160 4308 7257
rect -422 6960 -292 7070
rect -422 6870 -407 6960
rect -307 6870 -292 6960
rect 4178 7070 4193 7160
rect 4293 7070 4308 7160
rect 4178 6960 4308 7070
rect -422 6760 -292 6870
rect 4178 6870 4193 6960
rect 4293 6870 4308 6960
rect -422 6670 -407 6760
rect -307 6670 -292 6760
rect 4178 6760 4308 6870
rect -422 6560 -292 6670
rect -422 6470 -407 6560
rect -307 6470 -292 6560
rect 4178 6670 4193 6760
rect 4293 6670 4308 6760
rect 4178 6560 4308 6670
rect -422 6360 -292 6470
rect 4178 6470 4193 6560
rect 4293 6470 4308 6560
rect -422 6270 -407 6360
rect -307 6270 -292 6360
rect 4178 6360 4308 6470
rect -422 6160 -292 6270
rect 4178 6270 4193 6360
rect 4293 6270 4308 6360
rect -422 6070 -407 6160
rect -307 6070 -292 6160
rect -422 5960 -292 6070
rect 4178 6160 4308 6270
rect 4178 6070 4193 6160
rect 4293 6070 4308 6160
rect -422 5870 -407 5960
rect -307 5870 -292 5960
rect 4178 5960 4308 6070
rect -422 5760 -292 5870
rect -422 5670 -407 5760
rect -307 5670 -292 5760
rect 4178 5870 4193 5960
rect 4293 5870 4308 5960
rect 4178 5760 4308 5870
rect -2827 5618 -2273 5634
rect -2827 5570 -2796 5618
rect -2327 5570 -2273 5618
rect -2827 5552 -2273 5570
rect -2064 5618 -1510 5634
rect -2064 5570 -2033 5618
rect -1564 5570 -1510 5618
rect -2064 5552 -1510 5570
rect -1253 5618 -699 5634
rect -1253 5570 -1222 5618
rect -753 5570 -699 5618
rect -1253 5552 -699 5570
rect -422 5560 -292 5670
rect 4178 5670 4193 5760
rect 4293 5670 4308 5760
rect -422 5470 -407 5560
rect -307 5470 -292 5560
rect 4178 5560 4308 5670
rect -422 5360 -292 5470
rect 4178 5470 4193 5560
rect 4293 5470 4308 5560
rect -422 5270 -407 5360
rect -307 5270 -292 5360
rect -422 5160 -292 5270
rect 4178 5360 4308 5470
rect 4178 5270 4193 5360
rect 4293 5270 4308 5360
rect -422 5070 -407 5160
rect -307 5070 -292 5160
rect 4178 5160 4308 5270
rect -422 4960 -292 5070
rect -422 4870 -407 4960
rect -307 4870 -292 4960
rect 4178 5070 4193 5160
rect 4293 5070 4308 5160
rect 4178 4960 4308 5070
rect -422 4760 -292 4870
rect 4178 4870 4193 4960
rect 4293 4870 4308 4960
rect -422 4670 -407 4760
rect -307 4670 -292 4760
rect 4178 4760 4308 4870
rect -2827 4647 -2273 4663
rect -2827 4599 -2796 4647
rect -2327 4599 -2273 4647
rect -2827 4581 -2273 4599
rect -2064 4647 -1510 4663
rect -2064 4599 -2033 4647
rect -1564 4599 -1510 4647
rect -2064 4581 -1510 4599
rect -1253 4647 -699 4663
rect -1253 4599 -1222 4647
rect -753 4599 -699 4647
rect -1253 4581 -699 4599
rect -422 4560 -292 4670
rect 4178 4670 4193 4760
rect 4293 4670 4308 4760
rect -422 4470 -407 4560
rect -307 4470 -292 4560
rect -422 4360 -292 4470
rect 4178 4560 4308 4670
rect 4178 4470 4193 4560
rect 4293 4470 4308 4560
rect -422 4270 -407 4360
rect -307 4270 -292 4360
rect 4178 4360 4308 4470
rect -422 4160 -292 4270
rect 4178 4270 4193 4360
rect 4293 4270 4308 4360
rect -422 4070 -407 4160
rect -307 4070 -292 4160
rect -422 3960 -292 4070
rect 4178 4160 4308 4270
rect 4178 4070 4193 4160
rect 4293 4070 4308 4160
rect -422 3870 -407 3960
rect -307 3870 -292 3960
rect 4178 3960 4308 4070
rect -422 3777 -292 3870
rect 4178 3870 4193 3960
rect 4293 3870 4308 3960
rect 4178 3777 4308 3870
rect -422 3760 4308 3777
rect -2827 3672 -2273 3688
rect -2827 3624 -2796 3672
rect -2327 3624 -2273 3672
rect -2827 3606 -2273 3624
rect -2064 3671 -1510 3687
rect -2064 3623 -2033 3671
rect -1564 3623 -1510 3671
rect -2064 3605 -1510 3623
rect -1253 3671 -699 3687
rect -1253 3623 -1222 3671
rect -753 3623 -699 3671
rect -422 3670 -407 3760
rect -307 3670 -207 3760
rect -107 3670 -7 3760
rect 93 3670 193 3760
rect 293 3670 393 3760
rect 493 3670 593 3760
rect 693 3670 793 3760
rect 893 3670 993 3760
rect 1093 3670 1193 3760
rect 1293 3670 1393 3760
rect 1493 3670 1593 3760
rect 1693 3670 1793 3760
rect 1893 3670 1993 3760
rect 2093 3670 2193 3760
rect 2293 3670 2393 3760
rect 2493 3670 2593 3760
rect 2693 3670 2793 3760
rect 2893 3670 2993 3760
rect 3093 3670 3193 3760
rect 3293 3670 3393 3760
rect 3493 3670 3593 3760
rect 3693 3670 3793 3760
rect 3893 3670 3993 3760
rect 4093 3670 4193 3760
rect 4293 3670 4308 3760
rect -422 3657 4308 3670
rect -1253 3605 -699 3623
rect -2839 3437 3876 3463
rect -2839 3306 -2791 3437
rect -2646 3306 -2491 3437
rect -2346 3306 -2191 3437
rect -2046 3306 -1891 3437
rect -1746 3306 -1591 3437
rect -1446 3306 -1291 3437
rect -1146 3306 -991 3437
rect -846 3306 -691 3437
rect -546 3306 -391 3437
rect -246 3306 -91 3437
rect 54 3306 209 3437
rect 354 3306 509 3437
rect 654 3306 809 3437
rect 954 3306 1109 3437
rect 1254 3306 1409 3437
rect 1554 3306 1709 3437
rect 1854 3306 2009 3437
rect 2154 3306 2309 3437
rect 2454 3306 2609 3437
rect 2754 3306 2909 3437
rect 3054 3306 3209 3437
rect 3354 3306 3509 3437
rect 3654 3306 3876 3437
rect -2839 3276 3876 3306
rect -2839 2128 3876 2157
rect -2839 1997 -2795 2128
rect -2650 1997 -2495 2128
rect -2350 1997 -2195 2128
rect -2050 1997 -1895 2128
rect -1750 1997 -1595 2128
rect -1450 1997 -1295 2128
rect -1150 1997 -995 2128
rect -850 1997 -695 2128
rect -550 1997 -395 2128
rect -250 1997 -95 2128
rect 50 1997 205 2128
rect 350 1997 505 2128
rect 650 1997 805 2128
rect 950 1997 1105 2128
rect 1250 1997 1405 2128
rect 1550 1997 1705 2128
rect 1850 1997 2005 2128
rect 2150 1997 2305 2128
rect 2450 1997 2605 2128
rect 2750 1997 2905 2128
rect 3050 1997 3205 2128
rect 3350 1997 3505 2128
rect 3650 1997 3876 2128
rect -2839 1970 3876 1997
<< nsubdiff >>
rect -2761 6416 -2355 6436
rect -2761 6360 -2724 6416
rect -2412 6360 -2355 6416
rect -2761 6339 -2355 6360
rect -1998 6416 -1592 6436
rect -1998 6360 -1961 6416
rect -1649 6360 -1592 6416
rect -1998 6339 -1592 6360
rect -1187 6416 -781 6436
rect -1187 6360 -1150 6416
rect -838 6360 -781 6416
rect -1187 6339 -781 6360
rect -2761 5445 -2355 5465
rect -2761 5389 -2724 5445
rect -2412 5389 -2355 5445
rect -2761 5368 -2355 5389
rect -1998 5445 -1592 5465
rect -1998 5389 -1961 5445
rect -1649 5389 -1592 5445
rect -1998 5368 -1592 5389
rect -1187 5445 -781 5465
rect -1187 5389 -1150 5445
rect -838 5389 -781 5445
rect -1187 5368 -781 5389
rect -2761 4470 -2355 4490
rect -2761 4414 -2724 4470
rect -2412 4414 -2355 4470
rect -2761 4393 -2355 4414
rect -1998 4469 -1592 4489
rect -1998 4413 -1961 4469
rect -1649 4413 -1592 4469
rect -1998 4392 -1592 4413
rect -1187 4469 -781 4489
rect -1187 4413 -1150 4469
rect -838 4413 -781 4469
rect -1187 4392 -781 4413
<< psubdiffcont >>
rect -407 7270 -307 7360
rect -207 7270 -107 7360
rect -7 7270 93 7360
rect 193 7270 293 7360
rect 393 7270 493 7360
rect 593 7270 693 7360
rect 793 7270 893 7360
rect 993 7270 1093 7360
rect 1193 7270 1293 7360
rect 1393 7270 1493 7360
rect 1593 7270 1693 7360
rect 1793 7270 1893 7360
rect 1993 7270 2093 7360
rect 2193 7270 2293 7360
rect 2393 7270 2493 7360
rect 2593 7270 2693 7360
rect 2793 7270 2893 7360
rect 2993 7270 3093 7360
rect 3193 7270 3293 7360
rect 3393 7270 3493 7360
rect 3593 7270 3693 7360
rect 3793 7270 3893 7360
rect 3993 7270 4093 7360
rect 4193 7270 4293 7360
rect -407 7070 -307 7160
rect -407 6870 -307 6960
rect 4193 7070 4293 7160
rect 4193 6870 4293 6960
rect -407 6670 -307 6760
rect -407 6470 -307 6560
rect 4193 6670 4293 6760
rect 4193 6470 4293 6560
rect -407 6270 -307 6360
rect 4193 6270 4293 6360
rect -407 6070 -307 6160
rect 4193 6070 4293 6160
rect -407 5870 -307 5960
rect -407 5670 -307 5760
rect 4193 5870 4293 5960
rect -2796 5570 -2327 5618
rect -2033 5570 -1564 5618
rect -1222 5570 -753 5618
rect 4193 5670 4293 5760
rect -407 5470 -307 5560
rect 4193 5470 4293 5560
rect -407 5270 -307 5360
rect 4193 5270 4293 5360
rect -407 5070 -307 5160
rect -407 4870 -307 4960
rect 4193 5070 4293 5160
rect 4193 4870 4293 4960
rect -407 4670 -307 4760
rect -2796 4599 -2327 4647
rect -2033 4599 -1564 4647
rect -1222 4599 -753 4647
rect 4193 4670 4293 4760
rect -407 4470 -307 4560
rect 4193 4470 4293 4560
rect -407 4270 -307 4360
rect 4193 4270 4293 4360
rect -407 4070 -307 4160
rect 4193 4070 4293 4160
rect -407 3870 -307 3960
rect 4193 3870 4293 3960
rect -2796 3624 -2327 3672
rect -2033 3623 -1564 3671
rect -1222 3623 -753 3671
rect -407 3670 -307 3760
rect -207 3670 -107 3760
rect -7 3670 93 3760
rect 193 3670 293 3760
rect 393 3670 493 3760
rect 593 3670 693 3760
rect 793 3670 893 3760
rect 993 3670 1093 3760
rect 1193 3670 1293 3760
rect 1393 3670 1493 3760
rect 1593 3670 1693 3760
rect 1793 3670 1893 3760
rect 1993 3670 2093 3760
rect 2193 3670 2293 3760
rect 2393 3670 2493 3760
rect 2593 3670 2693 3760
rect 2793 3670 2893 3760
rect 2993 3670 3093 3760
rect 3193 3670 3293 3760
rect 3393 3670 3493 3760
rect 3593 3670 3693 3760
rect 3793 3670 3893 3760
rect 3993 3670 4093 3760
rect 4193 3670 4293 3760
rect -2791 3306 -2646 3437
rect -2491 3306 -2346 3437
rect -2191 3306 -2046 3437
rect -1891 3306 -1746 3437
rect -1591 3306 -1446 3437
rect -1291 3306 -1146 3437
rect -991 3306 -846 3437
rect -691 3306 -546 3437
rect -391 3306 -246 3437
rect -91 3306 54 3437
rect 209 3306 354 3437
rect 509 3306 654 3437
rect 809 3306 954 3437
rect 1109 3306 1254 3437
rect 1409 3306 1554 3437
rect 1709 3306 1854 3437
rect 2009 3306 2154 3437
rect 2309 3306 2454 3437
rect 2609 3306 2754 3437
rect 2909 3306 3054 3437
rect 3209 3306 3354 3437
rect 3509 3306 3654 3437
rect -2795 1997 -2650 2128
rect -2495 1997 -2350 2128
rect -2195 1997 -2050 2128
rect -1895 1997 -1750 2128
rect -1595 1997 -1450 2128
rect -1295 1997 -1150 2128
rect -995 1997 -850 2128
rect -695 1997 -550 2128
rect -395 1997 -250 2128
rect -95 1997 50 2128
rect 205 1997 350 2128
rect 505 1997 650 2128
rect 805 1997 950 2128
rect 1105 1997 1250 2128
rect 1405 1997 1550 2128
rect 1705 1997 1850 2128
rect 2005 1997 2150 2128
rect 2305 1997 2450 2128
rect 2605 1997 2750 2128
rect 2905 1997 3050 2128
rect 3205 1997 3350 2128
rect 3505 1997 3650 2128
<< nsubdiffcont >>
rect -2724 6360 -2412 6416
rect -1961 6360 -1649 6416
rect -1150 6360 -838 6416
rect -2724 5389 -2412 5445
rect -1961 5389 -1649 5445
rect -1150 5389 -838 5445
rect -2724 4414 -2412 4470
rect -1961 4413 -1649 4469
rect -1150 4413 -838 4469
<< polysilicon >>
rect 317 7107 3477 7137
rect 256 7094 3477 7107
rect 256 7043 271 7094
rect 322 7060 3477 7094
rect 322 7043 417 7060
rect 256 7028 417 7043
rect 317 6958 417 7028
rect 521 6958 621 7002
rect 725 6958 825 7002
rect 929 6958 1029 7060
rect 1133 6958 1233 7060
rect 1337 6958 1437 7002
rect 1541 6958 1641 7002
rect 1745 6958 1845 7060
rect 1949 6958 2049 7060
rect 2153 6958 2253 7002
rect 2357 6958 2457 7002
rect 2561 6958 2661 7060
rect 2765 6958 2865 7060
rect 2969 6958 3069 7002
rect 3173 6958 3273 7002
rect 3377 6958 3477 7060
rect 317 6794 417 6838
rect 521 6739 621 6838
rect 725 6739 825 6838
rect 929 6794 1029 6838
rect 1133 6794 1233 6838
rect 1337 6739 1437 6838
rect 1541 6739 1641 6838
rect 1745 6794 1845 6838
rect 1949 6794 2049 6838
rect 2153 6739 2253 6838
rect 2357 6739 2457 6838
rect 2561 6794 2661 6838
rect 2765 6794 2865 6838
rect 2969 6739 3069 6838
rect 3173 6739 3273 6838
rect 3377 6794 3477 6838
rect 317 6700 3477 6739
rect 131 6686 3477 6700
rect 131 6635 145 6686
rect 196 6662 3477 6686
rect 196 6635 417 6662
rect 131 6621 417 6635
rect 317 6553 417 6621
rect 521 6553 621 6597
rect 725 6553 825 6597
rect 929 6553 1029 6662
rect 1133 6553 1233 6662
rect 1337 6553 1437 6597
rect 1541 6553 1641 6597
rect 1745 6553 1845 6662
rect 1949 6553 2049 6662
rect 2153 6553 2253 6597
rect 2357 6553 2457 6597
rect 2561 6553 2661 6662
rect 2765 6553 2865 6662
rect 2969 6553 3069 6597
rect 3173 6553 3273 6597
rect 3377 6553 3477 6662
rect 317 6389 417 6433
rect 521 6340 621 6433
rect 725 6340 825 6433
rect 929 6389 1029 6433
rect 1133 6389 1233 6433
rect 1337 6340 1437 6433
rect 1541 6340 1641 6433
rect 1745 6389 1845 6433
rect 1949 6389 2049 6433
rect 2153 6340 2253 6433
rect 2357 6340 2457 6433
rect 2561 6389 2661 6433
rect 2765 6389 2865 6433
rect 2969 6340 3069 6433
rect 3173 6340 3273 6433
rect 3377 6389 3477 6433
rect 317 6310 3477 6340
rect -2665 6182 -2609 6226
rect -2505 6182 -2449 6226
rect -1902 6182 -1846 6226
rect -1742 6182 -1686 6226
rect -1091 6182 -1035 6226
rect -931 6182 -875 6226
rect 256 6297 3477 6310
rect 256 6246 271 6297
rect 322 6263 3477 6297
rect 322 6246 417 6263
rect 256 6231 417 6246
rect 317 6161 417 6231
rect 521 6161 621 6205
rect 725 6161 825 6205
rect 929 6161 1029 6263
rect 1133 6161 1233 6263
rect 1337 6161 1437 6205
rect 1541 6161 1641 6205
rect 1745 6161 1845 6263
rect 1949 6161 2049 6263
rect 2153 6161 2253 6205
rect 2357 6161 2457 6205
rect 2561 6161 2661 6263
rect 2765 6161 2865 6263
rect 2969 6161 3069 6205
rect 3173 6161 3273 6205
rect 3377 6161 3477 6263
rect -2665 6038 -2609 6082
rect -2739 6024 -2609 6038
rect -2739 5965 -2725 6024
rect -2662 5965 -2609 6024
rect -2739 5950 -2609 5965
rect -2665 5812 -2609 5950
rect -2505 5937 -2449 6082
rect -1902 6038 -1846 6082
rect -1976 6024 -1846 6038
rect -1976 5965 -1962 6024
rect -1899 5965 -1846 6024
rect -1976 5950 -1846 5965
rect -2561 5924 -2449 5937
rect -2561 5865 -2548 5924
rect -2485 5865 -2449 5924
rect -2561 5852 -2449 5865
rect -2505 5812 -2449 5852
rect -1902 5812 -1846 5950
rect -1742 5937 -1686 6082
rect -1091 6038 -1035 6082
rect -1165 6024 -1035 6038
rect -1165 5965 -1151 6024
rect -1088 5965 -1035 6024
rect -1165 5950 -1035 5965
rect -1798 5924 -1686 5937
rect -1798 5865 -1785 5924
rect -1722 5865 -1686 5924
rect -1798 5852 -1686 5865
rect -1742 5812 -1686 5852
rect -1091 5812 -1035 5950
rect -931 5937 -875 6082
rect -987 5924 -875 5937
rect -987 5865 -974 5924
rect -911 5865 -875 5924
rect -987 5852 -875 5865
rect -931 5812 -875 5852
rect 317 5997 417 6041
rect 521 5942 621 6041
rect 725 5942 825 6041
rect 929 5997 1029 6041
rect 1133 5997 1233 6041
rect 1337 5942 1437 6041
rect 1541 5942 1641 6041
rect 1745 5997 1845 6041
rect 1949 5997 2049 6041
rect 2153 5942 2253 6041
rect 2357 5942 2457 6041
rect 2561 5997 2661 6041
rect 2765 5997 2865 6041
rect 2969 5942 3069 6041
rect 3173 5942 3273 6041
rect 3377 5997 3477 6041
rect 317 5903 3477 5942
rect 131 5889 3477 5903
rect 131 5838 145 5889
rect 196 5865 3477 5889
rect 196 5838 417 5865
rect 131 5824 417 5838
rect -2665 5668 -2609 5712
rect -2505 5668 -2449 5712
rect -1902 5668 -1846 5712
rect -1742 5668 -1686 5712
rect -1091 5668 -1035 5712
rect -931 5668 -875 5712
rect 317 5756 417 5824
rect 521 5756 621 5800
rect 725 5756 825 5800
rect 929 5756 1029 5865
rect 1133 5756 1233 5865
rect 1337 5756 1437 5800
rect 1541 5756 1641 5800
rect 1745 5756 1845 5865
rect 1949 5756 2049 5865
rect 2153 5756 2253 5800
rect 2357 5756 2457 5800
rect 2561 5756 2661 5865
rect 2765 5756 2865 5865
rect 2969 5756 3069 5800
rect 3173 5756 3273 5800
rect 3377 5756 3477 5865
rect 317 5592 417 5636
rect 521 5543 621 5636
rect 725 5543 825 5636
rect 929 5592 1029 5636
rect 1133 5592 1233 5636
rect 1337 5543 1437 5636
rect 1541 5543 1641 5636
rect 1745 5592 1845 5636
rect 1949 5592 2049 5636
rect 2153 5543 2253 5636
rect 2357 5543 2457 5636
rect 2561 5592 2661 5636
rect 2765 5592 2865 5636
rect 2969 5543 3069 5636
rect 3173 5543 3273 5636
rect 3377 5592 3477 5636
rect 317 5513 3477 5543
rect 256 5500 3477 5513
rect 256 5449 271 5500
rect 322 5466 3477 5500
rect 322 5449 417 5466
rect 256 5434 417 5449
rect 317 5364 417 5434
rect 521 5364 621 5408
rect 725 5364 825 5408
rect 929 5364 1029 5466
rect 1133 5364 1233 5466
rect 1337 5364 1437 5408
rect 1541 5364 1641 5408
rect 1745 5364 1845 5466
rect 1949 5364 2049 5466
rect 2153 5364 2253 5408
rect 2357 5364 2457 5408
rect 2561 5364 2661 5466
rect 2765 5364 2865 5466
rect 2969 5364 3069 5408
rect 3173 5364 3273 5408
rect 3377 5364 3477 5466
rect -2665 5211 -2609 5255
rect -2505 5211 -2449 5255
rect -1902 5211 -1846 5255
rect -1742 5211 -1686 5255
rect -1091 5211 -1035 5255
rect -931 5211 -875 5255
rect 317 5200 417 5244
rect -2665 5067 -2609 5111
rect -2739 5053 -2609 5067
rect -2739 4994 -2725 5053
rect -2662 4994 -2609 5053
rect -2739 4979 -2609 4994
rect -2665 4841 -2609 4979
rect -2505 4966 -2449 5111
rect -1902 5067 -1846 5111
rect -1976 5053 -1846 5067
rect -1976 4994 -1962 5053
rect -1899 4994 -1846 5053
rect -1976 4979 -1846 4994
rect -2561 4953 -2449 4966
rect -2561 4894 -2548 4953
rect -2485 4894 -2449 4953
rect -2561 4881 -2449 4894
rect -2505 4841 -2449 4881
rect -1902 4841 -1846 4979
rect -1742 4966 -1686 5111
rect -1091 5067 -1035 5111
rect -1165 5053 -1035 5067
rect -1165 4994 -1151 5053
rect -1088 4994 -1035 5053
rect -1165 4979 -1035 4994
rect -1798 4953 -1686 4966
rect -1798 4894 -1785 4953
rect -1722 4894 -1686 4953
rect -1798 4881 -1686 4894
rect -1742 4841 -1686 4881
rect -1091 4841 -1035 4979
rect -931 4966 -875 5111
rect -987 4953 -875 4966
rect -987 4894 -974 4953
rect -911 4894 -875 4953
rect -987 4881 -875 4894
rect -931 4841 -875 4881
rect 521 5145 621 5244
rect 725 5145 825 5244
rect 929 5200 1029 5244
rect 1133 5200 1233 5244
rect 1337 5145 1437 5244
rect 1541 5145 1641 5244
rect 1745 5200 1845 5244
rect 1949 5200 2049 5244
rect 2153 5145 2253 5244
rect 2357 5145 2457 5244
rect 2561 5200 2661 5244
rect 2765 5200 2865 5244
rect 2969 5145 3069 5244
rect 3173 5145 3273 5244
rect 3377 5200 3477 5244
rect 317 5106 3477 5145
rect 131 5092 3477 5106
rect 131 5041 145 5092
rect 196 5068 3477 5092
rect 196 5041 417 5068
rect 131 5027 417 5041
rect 317 4959 417 5027
rect 521 4959 621 5003
rect 725 4959 825 5003
rect 929 4959 1029 5068
rect 1133 4959 1233 5068
rect 1337 4959 1437 5003
rect 1541 4959 1641 5003
rect 1745 4959 1845 5068
rect 1949 4959 2049 5068
rect 2153 4959 2253 5003
rect 2357 4959 2457 5003
rect 2561 4959 2661 5068
rect 2765 4959 2865 5068
rect 2969 4959 3069 5003
rect 3173 4959 3273 5003
rect 3377 4959 3477 5068
rect 317 4795 417 4839
rect -2665 4697 -2609 4741
rect -2505 4697 -2449 4741
rect -1902 4697 -1846 4741
rect -1742 4697 -1686 4741
rect -1091 4697 -1035 4741
rect -931 4697 -875 4741
rect 521 4746 621 4839
rect 725 4746 825 4839
rect 929 4795 1029 4839
rect 1133 4795 1233 4839
rect 1337 4746 1437 4839
rect 1541 4746 1641 4839
rect 1745 4795 1845 4839
rect 1949 4795 2049 4839
rect 2153 4746 2253 4839
rect 2357 4746 2457 4839
rect 2561 4795 2661 4839
rect 2765 4795 2865 4839
rect 2969 4746 3069 4839
rect 3173 4746 3273 4839
rect 3377 4795 3477 4839
rect 317 4716 3477 4746
rect 256 4703 3477 4716
rect 256 4652 271 4703
rect 322 4669 3477 4703
rect 322 4652 417 4669
rect 256 4637 417 4652
rect 317 4567 417 4637
rect 521 4567 621 4611
rect 725 4567 825 4611
rect 929 4567 1029 4669
rect 1133 4567 1233 4669
rect 1337 4567 1437 4611
rect 1541 4567 1641 4611
rect 1745 4567 1845 4669
rect 1949 4567 2049 4669
rect 2153 4567 2253 4611
rect 2357 4567 2457 4611
rect 2561 4567 2661 4669
rect 2765 4567 2865 4669
rect 2969 4567 3069 4611
rect 3173 4567 3273 4611
rect 3377 4567 3477 4669
rect 317 4403 417 4447
rect -2665 4236 -2609 4280
rect -2505 4236 -2449 4280
rect -1902 4235 -1846 4279
rect -1742 4235 -1686 4279
rect -1091 4235 -1035 4279
rect -931 4235 -875 4279
rect 521 4348 621 4447
rect 725 4348 825 4447
rect 929 4403 1029 4447
rect 1133 4403 1233 4447
rect 1337 4348 1437 4447
rect 1541 4348 1641 4447
rect 1745 4403 1845 4447
rect 1949 4403 2049 4447
rect 2153 4348 2253 4447
rect 2357 4348 2457 4447
rect 2561 4403 2661 4447
rect 2765 4403 2865 4447
rect 2969 4348 3069 4447
rect 3173 4348 3273 4447
rect 3377 4403 3477 4447
rect 317 4309 3477 4348
rect -2665 4092 -2609 4136
rect -2739 4078 -2609 4092
rect -2739 4019 -2725 4078
rect -2662 4019 -2609 4078
rect -2739 4004 -2609 4019
rect -2665 3866 -2609 4004
rect -2505 3991 -2449 4136
rect 131 4295 3477 4309
rect 131 4244 145 4295
rect 196 4271 3477 4295
rect 196 4244 417 4271
rect 131 4230 417 4244
rect 317 4162 417 4230
rect 521 4162 621 4206
rect 725 4162 825 4206
rect 929 4162 1029 4271
rect 1133 4162 1233 4271
rect 1337 4162 1437 4206
rect 1541 4162 1641 4206
rect 1745 4162 1845 4271
rect 1949 4162 2049 4271
rect 2153 4162 2253 4206
rect 2357 4162 2457 4206
rect 2561 4162 2661 4271
rect 2765 4162 2865 4271
rect 2969 4162 3069 4206
rect 3173 4162 3273 4206
rect 3377 4162 3477 4271
rect -1902 4091 -1846 4135
rect -1976 4077 -1846 4091
rect -1976 4018 -1962 4077
rect -1899 4018 -1846 4077
rect -1976 4003 -1846 4018
rect -2561 3978 -2449 3991
rect -2561 3919 -2548 3978
rect -2485 3919 -2449 3978
rect -2561 3906 -2449 3919
rect -2505 3866 -2449 3906
rect -1902 3865 -1846 4003
rect -1742 3990 -1686 4135
rect -1091 4091 -1035 4135
rect -1165 4077 -1035 4091
rect -1165 4018 -1151 4077
rect -1088 4018 -1035 4077
rect -1165 4003 -1035 4018
rect -1798 3977 -1686 3990
rect -1798 3918 -1785 3977
rect -1722 3918 -1686 3977
rect -1798 3905 -1686 3918
rect -1742 3865 -1686 3905
rect -1091 3865 -1035 4003
rect -931 3990 -875 4135
rect -987 3977 -875 3990
rect -987 3918 -974 3977
rect -911 3918 -875 3977
rect -987 3905 -875 3918
rect -931 3865 -875 3905
rect 317 3998 417 4042
rect 75 3960 167 3981
rect 75 3909 95 3960
rect 146 3949 167 3960
rect 521 3949 621 4042
rect 725 3949 825 4042
rect 929 3998 1029 4042
rect 1133 3998 1233 4042
rect 1337 3949 1437 4042
rect 1541 3949 1641 4042
rect 1745 3998 1845 4042
rect 1949 3998 2049 4042
rect 2153 3949 2253 4042
rect 2357 3949 2457 4042
rect 2561 3998 2661 4042
rect 2765 3998 2865 4042
rect 2969 3949 3069 4042
rect 3173 3949 3273 4042
rect 3377 3998 3477 4042
rect 146 3909 3273 3949
rect 75 3899 3273 3909
rect 75 3889 167 3899
rect -2665 3722 -2609 3766
rect -2505 3722 -2449 3766
rect -1902 3721 -1846 3765
rect -1742 3721 -1686 3765
rect -1091 3721 -1035 3765
rect -931 3721 -875 3765
rect -3007 3255 -2921 3269
rect -3007 3251 3697 3255
rect -3007 3202 -2989 3251
rect -2941 3202 3697 3251
rect -3007 3197 3697 3202
rect -3007 3186 -2921 3197
rect -2727 3070 -2627 3197
rect -2523 3070 -2423 3114
rect -2319 3070 -2219 3114
rect -2115 3070 -2015 3197
rect -1911 3070 -1811 3197
rect -1707 3070 -1607 3114
rect -1503 3070 -1403 3114
rect -1299 3070 -1199 3197
rect -1095 3070 -995 3197
rect -891 3070 -791 3114
rect -687 3070 -587 3114
rect -483 3070 -383 3197
rect -279 3070 -179 3197
rect -75 3070 25 3114
rect 129 3070 229 3114
rect 333 3070 433 3197
rect 537 3070 637 3197
rect 741 3070 841 3114
rect 945 3070 1045 3114
rect 1149 3070 1249 3197
rect 1353 3070 1453 3197
rect 1557 3070 1657 3114
rect 1761 3070 1861 3114
rect 1965 3070 2065 3197
rect 2169 3070 2269 3197
rect 2373 3070 2473 3114
rect 2577 3070 2677 3114
rect 2781 3070 2881 3197
rect 2985 3070 3085 3197
rect 3189 3070 3289 3114
rect 3393 3070 3493 3114
rect 3597 3070 3697 3197
rect -2727 2786 -2627 2830
rect -3010 2731 -2923 2744
rect -2523 2731 -2423 2830
rect -2319 2731 -2219 2830
rect -2115 2786 -2015 2830
rect -1911 2786 -1811 2830
rect -1707 2731 -1607 2830
rect -1503 2731 -1403 2830
rect -1299 2786 -1199 2830
rect -1095 2786 -995 2830
rect -891 2731 -791 2830
rect -687 2731 -587 2830
rect -483 2786 -383 2830
rect -279 2786 -179 2830
rect -75 2731 25 2830
rect 129 2731 229 2830
rect 333 2786 433 2830
rect 537 2786 637 2830
rect 741 2731 841 2830
rect 945 2731 1045 2830
rect 1149 2786 1249 2830
rect 1353 2786 1453 2830
rect 1557 2731 1657 2830
rect 1761 2731 1861 2830
rect 1965 2786 2065 2830
rect 2169 2786 2269 2830
rect 2373 2731 2473 2830
rect 2577 2731 2677 2830
rect 2781 2786 2881 2830
rect 2985 2786 3085 2830
rect 3189 2731 3289 2830
rect 3393 2731 3493 2830
rect 3597 2786 3697 2830
rect -3010 2730 3697 2731
rect -3010 2677 -2997 2730
rect -2941 2677 3697 2730
rect -3010 2672 3697 2677
rect -3010 2663 -2923 2672
rect -2727 2579 -2627 2672
rect -2523 2579 -2423 2623
rect -2319 2579 -2219 2623
rect -2115 2579 -2015 2672
rect -1911 2579 -1811 2672
rect -1707 2579 -1607 2623
rect -1503 2579 -1403 2623
rect -1299 2579 -1199 2672
rect -1095 2579 -995 2672
rect -891 2579 -791 2623
rect -687 2579 -587 2623
rect -483 2579 -383 2672
rect -279 2579 -179 2672
rect -75 2579 25 2623
rect 129 2579 229 2623
rect 333 2579 433 2672
rect 537 2579 637 2672
rect 741 2579 841 2623
rect 945 2579 1045 2623
rect 1149 2579 1249 2672
rect 1353 2579 1453 2672
rect 1557 2579 1657 2623
rect 1761 2579 1861 2623
rect 1965 2579 2065 2672
rect 2169 2579 2269 2672
rect 2373 2579 2473 2623
rect 2577 2579 2677 2623
rect 2781 2579 2881 2672
rect 2985 2579 3085 2672
rect 3189 2579 3289 2623
rect 3393 2579 3493 2623
rect 3597 2579 3697 2672
rect -2727 2295 -2627 2339
rect -3005 2236 -2913 2252
rect -2523 2236 -2423 2339
rect -2319 2236 -2219 2339
rect -2115 2295 -2015 2339
rect -1911 2295 -1811 2339
rect -1707 2236 -1607 2339
rect -1503 2236 -1403 2339
rect -1299 2295 -1199 2339
rect -1095 2295 -995 2339
rect -891 2236 -791 2339
rect -687 2236 -587 2339
rect -483 2295 -383 2339
rect -279 2295 -179 2339
rect -75 2236 25 2339
rect 129 2236 229 2339
rect 333 2295 433 2339
rect 537 2295 637 2339
rect 741 2236 841 2339
rect 945 2236 1045 2339
rect 1149 2295 1249 2339
rect 1353 2295 1453 2339
rect 1557 2236 1657 2339
rect 1761 2236 1861 2339
rect 1965 2295 2065 2339
rect 2169 2295 2269 2339
rect 2373 2236 2473 2339
rect 2577 2236 2677 2339
rect 2781 2295 2881 2339
rect 2985 2295 3085 2339
rect 3189 2236 3289 2339
rect 3393 2236 3493 2339
rect 3597 2295 3697 2339
rect -3005 2231 3493 2236
rect -3005 2180 -2989 2231
rect -2941 2180 3493 2231
rect -3005 2177 3493 2180
rect -3005 2164 -2913 2177
<< polycontact >>
rect 271 7043 322 7094
rect 145 6635 196 6686
rect 271 6246 322 6297
rect -2725 5965 -2662 6024
rect -1962 5965 -1899 6024
rect -2548 5865 -2485 5924
rect -1151 5965 -1088 6024
rect -1785 5865 -1722 5924
rect -974 5865 -911 5924
rect 145 5838 196 5889
rect 271 5449 322 5500
rect -2725 4994 -2662 5053
rect -1962 4994 -1899 5053
rect -2548 4894 -2485 4953
rect -1151 4994 -1088 5053
rect -1785 4894 -1722 4953
rect -974 4894 -911 4953
rect 145 5041 196 5092
rect 271 4652 322 4703
rect -2725 4019 -2662 4078
rect 145 4244 196 4295
rect -1962 4018 -1899 4077
rect -2548 3919 -2485 3978
rect -1151 4018 -1088 4077
rect -1785 3918 -1722 3977
rect -974 3918 -911 3977
rect 95 3909 146 3960
rect -2989 3202 -2941 3251
rect -2997 2677 -2941 2730
rect -2989 2180 -2941 2231
<< metal1 >>
rect 3645 7677 3729 7689
rect 3645 7621 3661 7677
rect 3716 7621 3729 7677
rect 3645 7608 3729 7621
rect 3846 7674 3930 7686
rect 3846 7618 3862 7674
rect 3917 7618 3930 7674
rect 3846 7605 3930 7618
rect 3643 7543 3727 7555
rect 3643 7487 3659 7543
rect 3714 7487 3727 7543
rect 3643 7474 3727 7487
rect 3851 7538 3935 7550
rect 3851 7482 3867 7538
rect 3922 7482 3935 7538
rect 3851 7469 3935 7482
rect -422 7360 -292 7377
rect -422 7270 -407 7360
rect -307 7343 -292 7360
rect -222 7360 -92 7377
rect -222 7343 -207 7360
rect -307 7297 -207 7343
rect -307 7270 -292 7297
rect -422 7257 -292 7270
rect -222 7270 -207 7297
rect -107 7343 -92 7360
rect -22 7360 108 7377
rect -22 7343 -7 7360
rect -107 7297 -7 7343
rect -107 7270 -92 7297
rect -222 7257 -92 7270
rect -22 7270 -7 7297
rect 93 7343 108 7360
rect 178 7360 308 7377
rect 178 7343 193 7360
rect 93 7297 193 7343
rect 93 7270 108 7297
rect -22 7257 108 7270
rect 178 7270 193 7297
rect 293 7343 308 7360
rect 378 7360 508 7377
rect 378 7343 393 7360
rect 293 7297 393 7343
rect 293 7270 308 7297
rect 178 7257 308 7270
rect 378 7270 393 7297
rect 493 7343 508 7360
rect 578 7360 708 7377
rect 578 7343 593 7360
rect 493 7297 593 7343
rect 493 7270 508 7297
rect 378 7257 508 7270
rect 578 7270 593 7297
rect 693 7343 708 7360
rect 778 7360 908 7377
rect 778 7343 793 7360
rect 693 7297 793 7343
rect 693 7270 708 7297
rect 578 7257 708 7270
rect 778 7270 793 7297
rect 893 7343 908 7360
rect 978 7360 1108 7377
rect 978 7343 993 7360
rect 893 7297 993 7343
rect 893 7270 908 7297
rect 778 7257 908 7270
rect 978 7270 993 7297
rect 1093 7343 1108 7360
rect 1178 7360 1308 7377
rect 1178 7343 1193 7360
rect 1093 7297 1193 7343
rect 1093 7270 1108 7297
rect 978 7257 1108 7270
rect 1178 7270 1193 7297
rect 1293 7343 1308 7360
rect 1378 7360 1508 7377
rect 1378 7343 1393 7360
rect 1293 7297 1393 7343
rect 1293 7270 1308 7297
rect 1178 7257 1308 7270
rect 1378 7270 1393 7297
rect 1493 7343 1508 7360
rect 1578 7360 1708 7377
rect 1578 7343 1593 7360
rect 1493 7297 1593 7343
rect 1493 7270 1508 7297
rect 1378 7257 1508 7270
rect 1578 7270 1593 7297
rect 1693 7343 1708 7360
rect 1778 7360 1908 7377
rect 1778 7343 1793 7360
rect 1693 7297 1793 7343
rect 1693 7270 1708 7297
rect 1578 7257 1708 7270
rect 1778 7270 1793 7297
rect 1893 7343 1908 7360
rect 1978 7360 2108 7377
rect 1978 7343 1993 7360
rect 1893 7297 1993 7343
rect 1893 7270 1908 7297
rect 1778 7257 1908 7270
rect 1978 7270 1993 7297
rect 2093 7343 2108 7360
rect 2178 7360 2308 7377
rect 2178 7343 2193 7360
rect 2093 7297 2193 7343
rect 2093 7270 2108 7297
rect 1978 7257 2108 7270
rect 2178 7270 2193 7297
rect 2293 7343 2308 7360
rect 2378 7360 2508 7377
rect 2378 7343 2393 7360
rect 2293 7297 2393 7343
rect 2293 7270 2308 7297
rect 2178 7257 2308 7270
rect 2378 7270 2393 7297
rect 2493 7343 2508 7360
rect 2578 7360 2708 7377
rect 2578 7343 2593 7360
rect 2493 7297 2593 7343
rect 2493 7270 2508 7297
rect 2378 7257 2508 7270
rect 2578 7270 2593 7297
rect 2693 7343 2708 7360
rect 2778 7360 2908 7377
rect 2778 7343 2793 7360
rect 2693 7297 2793 7343
rect 2693 7270 2708 7297
rect 2578 7257 2708 7270
rect 2778 7270 2793 7297
rect 2893 7343 2908 7360
rect 2978 7360 3108 7377
rect 2978 7343 2993 7360
rect 2893 7297 2993 7343
rect 2893 7270 2908 7297
rect 2778 7257 2908 7270
rect 2978 7270 2993 7297
rect 3093 7343 3108 7360
rect 3178 7360 3308 7377
rect 3178 7343 3193 7360
rect 3093 7297 3193 7343
rect 3093 7270 3108 7297
rect 2978 7257 3108 7270
rect 3178 7270 3193 7297
rect 3293 7343 3308 7360
rect 3378 7360 3508 7377
rect 3378 7343 3393 7360
rect 3293 7297 3393 7343
rect 3293 7270 3308 7297
rect 3178 7257 3308 7270
rect 3378 7270 3393 7297
rect 3493 7343 3508 7360
rect 3578 7360 3708 7377
rect 3578 7343 3593 7360
rect 3493 7297 3593 7343
rect 3493 7270 3508 7297
rect 3378 7257 3508 7270
rect 3578 7270 3593 7297
rect 3693 7343 3708 7360
rect 3778 7360 3908 7377
rect 3778 7343 3793 7360
rect 3693 7297 3793 7343
rect 3693 7270 3708 7297
rect 3578 7257 3708 7270
rect 3778 7270 3793 7297
rect 3893 7343 3908 7360
rect 3978 7360 4108 7377
rect 3978 7343 3993 7360
rect 3893 7297 3993 7343
rect 3893 7270 3908 7297
rect 3778 7257 3908 7270
rect 3978 7270 3993 7297
rect 4093 7343 4108 7360
rect 4178 7360 4308 7377
rect 4178 7343 4193 7360
rect 4093 7297 4193 7343
rect 4093 7270 4108 7297
rect 3978 7257 4108 7270
rect 4178 7270 4193 7297
rect 4293 7270 4308 7360
rect 4178 7257 4308 7270
rect -393 7177 -347 7257
rect 4220 7177 4266 7257
rect -422 7160 -292 7177
rect -422 7070 -407 7160
rect -307 7070 -292 7160
rect 454 7130 3348 7170
rect 4178 7160 4308 7177
rect -422 7057 -292 7070
rect 81 7101 159 7113
rect -393 6977 -347 7057
rect 81 7047 93 7101
rect 147 7097 159 7101
rect 256 7097 335 7107
rect 147 7094 335 7097
rect 147 7051 271 7094
rect 147 7047 159 7051
rect 81 7039 159 7047
rect 256 7043 271 7051
rect 322 7043 335 7094
rect 256 7028 335 7043
rect 446 7084 3355 7130
rect -422 6960 -292 6977
rect -422 6870 -407 6960
rect -307 6870 -292 6960
rect 446 6957 492 7084
rect 641 7026 699 7028
rect 629 7019 711 7026
rect 629 6963 642 7019
rect 698 6963 711 7019
rect -422 6857 -292 6870
rect 242 6945 288 6956
rect -393 6777 -347 6857
rect 443 6945 494 6957
rect 629 6951 711 6963
rect 854 6957 900 7084
rect 443 6851 446 6945
rect 492 6851 494 6945
rect 228 6841 310 6851
rect 228 6785 240 6841
rect 296 6785 310 6841
rect 443 6839 494 6851
rect 650 6945 696 6951
rect 650 6840 696 6851
rect 851 6945 902 6957
rect 851 6851 854 6945
rect 900 6851 902 6945
rect 851 6839 902 6851
rect 1058 6945 1104 6956
rect 1058 6848 1104 6851
rect 1234 6945 1325 7084
rect 1450 7019 1532 7026
rect 1450 6963 1462 7019
rect 1518 6963 1532 7019
rect 1450 6951 1532 6963
rect 1234 6851 1262 6945
rect 1308 6851 1325 6945
rect -422 6760 -292 6777
rect 228 6776 310 6785
rect 1038 6838 1119 6848
rect 1038 6782 1051 6838
rect 1107 6782 1119 6838
rect -422 6670 -407 6760
rect -307 6670 -292 6760
rect 1038 6774 1119 6782
rect 1038 6746 1096 6774
rect -422 6657 -292 6670
rect -90 6692 -12 6704
rect 650 6700 1096 6746
rect -393 6577 -347 6657
rect -90 6638 -78 6692
rect -24 6688 -12 6692
rect 131 6688 210 6700
rect -24 6686 210 6688
rect -24 6642 145 6686
rect -24 6638 -12 6642
rect -90 6632 -12 6638
rect 131 6635 145 6642
rect 196 6635 210 6686
rect 523 6661 597 6673
rect 523 6656 533 6661
rect 131 6621 210 6635
rect 326 6610 533 6656
rect -422 6560 -292 6577
rect -422 6470 -407 6560
rect -307 6470 -292 6560
rect 326 6552 372 6610
rect 523 6605 533 6610
rect 589 6605 597 6661
rect 523 6593 597 6605
rect -3641 6446 -2275 6462
rect -2076 6446 -1512 6462
rect -1265 6446 -701 6462
rect -422 6457 -292 6470
rect 239 6540 372 6552
rect -3641 6416 -701 6446
rect -3641 6403 -2724 6416
rect -3641 6336 -3203 6403
rect -3136 6360 -2724 6403
rect -2412 6360 -1961 6416
rect -1649 6360 -1150 6416
rect -838 6360 -701 6416
rect -393 6377 -347 6457
rect 239 6446 242 6540
rect 288 6481 372 6540
rect 443 6540 494 6552
rect 288 6446 290 6481
rect 239 6434 290 6446
rect 443 6446 446 6540
rect 492 6446 494 6540
rect 443 6434 494 6446
rect 650 6540 696 6700
rect 1042 6603 1124 6611
rect 650 6435 696 6446
rect 851 6540 902 6552
rect 851 6446 854 6540
rect 900 6446 902 6540
rect 1042 6547 1057 6603
rect 1113 6547 1124 6603
rect 1042 6540 1124 6547
rect 1042 6539 1058 6540
rect 851 6434 902 6446
rect 1104 6539 1124 6540
rect 1234 6540 1325 6851
rect 1466 6945 1512 6951
rect 1466 6840 1512 6851
rect 1643 6945 1734 7084
rect 1643 6851 1670 6945
rect 1716 6851 1734 6945
rect 1445 6768 1530 6783
rect 1445 6712 1458 6768
rect 1514 6712 1530 6768
rect 1445 6702 1530 6712
rect 1058 6435 1104 6446
rect 1234 6446 1262 6540
rect 1308 6446 1325 6540
rect -3136 6336 -701 6360
rect -3641 6331 -701 6336
rect -3641 6312 -2275 6331
rect -2076 6312 -1512 6331
rect -1265 6312 -701 6331
rect -422 6360 -292 6377
rect -2743 6169 -2692 6312
rect -2743 6095 -2740 6169
rect -2694 6095 -2692 6169
rect -2743 6093 -2692 6095
rect -2580 6169 -2534 6180
rect -2740 6084 -2694 6093
rect -2580 6042 -2534 6095
rect -2420 6169 -2374 6312
rect -2420 6084 -2374 6095
rect -1980 6169 -1929 6312
rect -1980 6095 -1977 6169
rect -1931 6095 -1929 6169
rect -1980 6093 -1929 6095
rect -1817 6169 -1771 6180
rect -1977 6084 -1931 6093
rect -1817 6042 -1771 6095
rect -1657 6169 -1611 6312
rect -1657 6084 -1611 6095
rect -1169 6169 -1118 6312
rect -1169 6095 -1166 6169
rect -1120 6095 -1118 6169
rect -1169 6093 -1118 6095
rect -1006 6169 -960 6180
rect -1166 6084 -1120 6093
rect -1006 6042 -960 6095
rect -846 6169 -800 6312
rect -422 6270 -407 6360
rect -307 6270 -292 6360
rect 446 6350 492 6434
rect 854 6350 900 6434
rect 1234 6350 1325 6446
rect 1466 6540 1512 6702
rect 1466 6435 1512 6446
rect 1643 6540 1734 6851
rect 1874 6945 1920 6956
rect 1874 6848 1920 6851
rect 2058 6945 2149 7084
rect 2266 7019 2348 7026
rect 2266 6963 2278 7019
rect 2334 6963 2348 7019
rect 2266 6951 2348 6963
rect 2058 6851 2078 6945
rect 2124 6851 2149 6945
rect 1852 6838 1933 6848
rect 1852 6782 1863 6838
rect 1919 6782 1933 6838
rect 1852 6774 1933 6782
rect 1643 6446 1670 6540
rect 1716 6446 1734 6540
rect 1852 6601 1936 6614
rect 1852 6545 1866 6601
rect 1922 6545 1936 6601
rect 1852 6540 1936 6545
rect 1852 6537 1874 6540
rect 1643 6350 1734 6446
rect 1920 6537 1936 6540
rect 2058 6540 2149 6851
rect 2282 6945 2328 6951
rect 2282 6840 2328 6851
rect 2461 6945 2552 7084
rect 2894 6957 2940 7084
rect 3079 7019 3161 7026
rect 3079 6963 3092 7019
rect 3148 6963 3161 7019
rect 2461 6851 2486 6945
rect 2532 6851 2552 6945
rect 2260 6763 2345 6771
rect 2260 6707 2273 6763
rect 2329 6707 2345 6763
rect 2260 6699 2345 6707
rect 1874 6435 1920 6446
rect 2058 6446 2078 6540
rect 2124 6446 2149 6540
rect 2058 6350 2149 6446
rect 2282 6540 2328 6699
rect 2282 6435 2328 6446
rect 2461 6540 2552 6851
rect 2690 6945 2736 6956
rect 2690 6850 2736 6851
rect 2891 6945 2941 6957
rect 3079 6951 3161 6963
rect 3302 6958 3348 7084
rect 4178 7070 4193 7160
rect 4293 7070 4308 7160
rect 4178 7057 4308 7070
rect 4220 6977 4266 7057
rect 4178 6960 4308 6977
rect 2891 6851 2894 6945
rect 2940 6851 2941 6945
rect 2674 6838 2754 6850
rect 2891 6839 2941 6851
rect 3098 6945 3144 6951
rect 3098 6840 3144 6851
rect 3300 6945 3349 6958
rect 3300 6851 3302 6945
rect 3348 6851 3349 6945
rect 3300 6839 3349 6851
rect 3506 6945 3552 6956
rect 4178 6870 4193 6960
rect 4293 6870 4308 6960
rect 4178 6857 4308 6870
rect 2674 6782 2683 6838
rect 2739 6791 2754 6838
rect 3506 6792 3552 6851
rect 3824 6796 3906 6812
rect 3824 6792 3837 6796
rect 3494 6791 3837 6792
rect 2739 6782 3837 6791
rect 2674 6774 3837 6782
rect 2678 6746 3837 6774
rect 2678 6745 3552 6746
rect 2461 6446 2486 6540
rect 2532 6446 2552 6540
rect 2672 6599 2754 6609
rect 2672 6543 2685 6599
rect 2741 6543 2754 6599
rect 2672 6540 2754 6543
rect 2672 6532 2690 6540
rect 2461 6350 2552 6446
rect 2736 6532 2754 6540
rect 2891 6540 2942 6552
rect 2690 6435 2736 6446
rect 2891 6446 2894 6540
rect 2940 6446 2942 6540
rect 2891 6434 2942 6446
rect 3098 6540 3144 6745
rect 3824 6742 3837 6746
rect 3891 6742 3906 6796
rect 4220 6777 4266 6857
rect 3824 6736 3906 6742
rect 4178 6760 4308 6777
rect 4178 6670 4193 6760
rect 4293 6670 4308 6760
rect 4178 6657 4308 6670
rect 3488 6600 3571 6609
rect 3098 6435 3144 6446
rect 3299 6540 3350 6552
rect 3299 6446 3302 6540
rect 3348 6446 3350 6540
rect 3488 6546 3502 6600
rect 3556 6546 3571 6600
rect 4220 6577 4266 6657
rect 3488 6540 3571 6546
rect 3488 6535 3506 6540
rect 3299 6434 3350 6446
rect 3552 6535 3571 6540
rect 4178 6560 4308 6577
rect 4178 6470 4193 6560
rect 4293 6470 4308 6560
rect 4178 6457 4308 6470
rect 3506 6435 3552 6446
rect 2894 6350 2940 6434
rect 3302 6350 3348 6434
rect 4220 6377 4266 6457
rect 4178 6360 4308 6377
rect -422 6257 -292 6270
rect 80 6302 158 6311
rect 256 6302 335 6310
rect -393 6177 -347 6257
rect 80 6246 92 6302
rect 148 6297 335 6302
rect 148 6246 271 6297
rect 322 6246 335 6297
rect 80 6237 158 6246
rect 256 6231 335 6246
rect 446 6304 3357 6350
rect 446 6287 3355 6304
rect -846 6084 -800 6095
rect -422 6160 -292 6177
rect 446 6160 492 6287
rect 641 6229 699 6231
rect 629 6222 711 6229
rect 629 6166 642 6222
rect 698 6166 711 6222
rect -422 6070 -407 6160
rect -307 6070 -292 6160
rect -422 6057 -292 6070
rect 242 6148 288 6159
rect -2580 6038 -2471 6042
rect -1817 6038 -1708 6042
rect -1006 6038 -897 6042
rect -634 6038 -553 6052
rect -2739 6024 -2650 6038
rect -2739 5996 -2725 6024
rect -2840 5965 -2725 5996
rect -2662 5965 -2650 6024
rect -2580 5996 -2031 6038
rect -1976 6024 -1887 6038
rect -1976 5996 -1962 6024
rect -2504 5992 -1962 5996
rect -2840 5960 -2650 5965
rect -3625 5950 -2650 5960
rect -3625 5902 -2794 5950
rect -2559 5924 -2474 5935
rect -2559 5902 -2548 5924
rect -3625 5878 -2548 5902
rect -2840 5865 -2548 5878
rect -2485 5865 -2474 5924
rect -2840 5856 -2474 5865
rect -2740 5799 -2694 5810
rect -2580 5809 -2534 5810
rect -2740 5645 -2694 5725
rect -2593 5799 -2526 5809
rect -2593 5725 -2580 5799
rect -2534 5725 -2526 5799
rect -2593 5711 -2526 5725
rect -2420 5799 -2374 5992
rect -2077 5965 -1962 5992
rect -1899 5965 -1887 6024
rect -1817 6002 -1512 6038
rect -1165 6028 -1076 6038
rect -1817 5996 -1600 6002
rect -1741 5992 -1600 5996
rect -2077 5950 -1887 5965
rect -2077 5902 -2031 5950
rect -1657 5946 -1600 5992
rect -1544 5992 -1512 6002
rect -1176 6024 -1076 6028
rect -1176 6022 -1151 6024
rect -1176 5996 -1165 6022
rect -1544 5946 -1534 5992
rect -1266 5966 -1165 5996
rect -1266 5965 -1151 5966
rect -1088 5965 -1076 6024
rect -1006 6036 -488 6038
rect -1006 5996 -621 6036
rect -930 5992 -621 5996
rect -1266 5950 -1076 5965
rect -1796 5924 -1711 5935
rect -1796 5902 -1785 5924
rect -2077 5865 -1785 5902
rect -1722 5865 -1711 5924
rect -2077 5856 -1711 5865
rect -1657 5934 -1534 5946
rect -2420 5714 -2374 5725
rect -1977 5799 -1931 5810
rect -1817 5809 -1771 5810
rect -1977 5645 -1931 5725
rect -1830 5799 -1763 5809
rect -1830 5725 -1817 5799
rect -1771 5725 -1763 5799
rect -1830 5711 -1763 5725
rect -1657 5799 -1611 5934
rect -985 5924 -900 5935
rect -1315 5902 -1233 5903
rect -985 5902 -974 5924
rect -1315 5865 -974 5902
rect -911 5865 -900 5924
rect -1315 5809 -1299 5865
rect -1243 5856 -900 5865
rect -1243 5809 -1233 5856
rect -1315 5798 -1233 5809
rect -1166 5799 -1120 5810
rect -1006 5809 -960 5810
rect -1657 5714 -1611 5725
rect -1166 5645 -1120 5725
rect -1019 5799 -952 5809
rect -1019 5725 -1006 5799
rect -960 5725 -952 5799
rect -1019 5711 -952 5725
rect -846 5799 -800 5992
rect -634 5980 -621 5992
rect -565 5992 -488 6036
rect -565 5980 -553 5992
rect -634 5970 -553 5980
rect -393 5977 -347 6057
rect 443 6148 494 6160
rect 629 6154 711 6166
rect 854 6160 900 6287
rect 443 6054 446 6148
rect 492 6054 494 6148
rect 228 6044 310 6054
rect 228 5988 240 6044
rect 296 5988 310 6044
rect 443 6042 494 6054
rect 650 6148 696 6154
rect 650 6043 696 6054
rect 851 6148 902 6160
rect 851 6054 854 6148
rect 900 6054 902 6148
rect 851 6042 902 6054
rect 1058 6148 1104 6159
rect 1058 6051 1104 6054
rect 1234 6148 1325 6287
rect 1450 6222 1532 6229
rect 1450 6166 1462 6222
rect 1518 6166 1532 6222
rect 1450 6154 1532 6166
rect 1234 6054 1262 6148
rect 1308 6054 1325 6148
rect 228 5979 310 5988
rect 1038 6041 1119 6051
rect 1038 5985 1051 6041
rect 1107 5985 1119 6041
rect 1038 5977 1119 5985
rect -422 5960 -292 5977
rect -422 5870 -407 5960
rect -307 5870 -292 5960
rect 1038 5949 1096 5977
rect 650 5903 1096 5949
rect -422 5857 -292 5870
rect -93 5887 -15 5894
rect 131 5889 210 5903
rect 131 5887 145 5889
rect -393 5777 -347 5857
rect -93 5831 -79 5887
rect -23 5838 145 5887
rect 196 5838 210 5889
rect 523 5864 597 5876
rect 523 5859 533 5864
rect -23 5831 210 5838
rect -93 5822 -15 5831
rect 131 5824 210 5831
rect 326 5813 533 5859
rect -846 5714 -800 5725
rect -422 5760 -292 5777
rect -422 5670 -407 5760
rect -307 5670 -292 5760
rect 326 5755 372 5813
rect 523 5808 533 5813
rect 589 5808 597 5864
rect 523 5796 597 5808
rect -422 5657 -292 5670
rect 239 5743 372 5755
rect -3025 5629 -2939 5643
rect -2863 5638 -2247 5645
rect -2100 5638 -1484 5645
rect -1289 5638 -673 5645
rect -2863 5629 -673 5638
rect -3025 5628 -673 5629
rect -3025 5563 -3013 5628
rect -2948 5618 -673 5628
rect -2948 5570 -2796 5618
rect -2327 5571 -2033 5618
rect -2327 5570 -2247 5571
rect -2948 5563 -2247 5570
rect -3025 5562 -2247 5563
rect -3025 5556 -2939 5562
rect -2863 5547 -2247 5562
rect -2100 5570 -2033 5571
rect -1564 5571 -1222 5618
rect -1564 5570 -1484 5571
rect -2100 5547 -1484 5570
rect -1289 5570 -1222 5571
rect -753 5570 -673 5618
rect -393 5577 -347 5657
rect 239 5649 242 5743
rect 288 5684 372 5743
rect 443 5743 494 5755
rect 288 5649 290 5684
rect 239 5637 290 5649
rect 443 5649 446 5743
rect 492 5649 494 5743
rect 443 5637 494 5649
rect 650 5743 696 5903
rect 1042 5806 1124 5814
rect 650 5638 696 5649
rect 851 5743 902 5755
rect 851 5649 854 5743
rect 900 5649 902 5743
rect 1042 5750 1057 5806
rect 1113 5750 1124 5806
rect 1042 5743 1124 5750
rect 1042 5742 1058 5743
rect 851 5637 902 5649
rect 1104 5742 1124 5743
rect 1234 5743 1325 6054
rect 1466 6148 1512 6154
rect 1466 6043 1512 6054
rect 1643 6148 1734 6287
rect 1643 6054 1670 6148
rect 1716 6054 1734 6148
rect 1445 5971 1530 5986
rect 1445 5915 1458 5971
rect 1514 5915 1530 5971
rect 1445 5905 1530 5915
rect 1058 5638 1104 5649
rect 1234 5649 1262 5743
rect 1308 5649 1325 5743
rect -1289 5547 -673 5570
rect -422 5560 -292 5577
rect -3218 5472 -3108 5473
rect -2839 5472 -2275 5491
rect -2076 5472 -1512 5491
rect -1265 5472 -701 5491
rect -3218 5452 -701 5472
rect -422 5470 -407 5560
rect -307 5470 -292 5560
rect 446 5553 492 5637
rect 854 5553 900 5637
rect 1234 5553 1325 5649
rect 1466 5743 1512 5905
rect 1466 5638 1512 5649
rect 1643 5743 1734 6054
rect 1874 6148 1920 6159
rect 1874 6051 1920 6054
rect 2058 6148 2149 6287
rect 2266 6222 2348 6229
rect 2266 6166 2278 6222
rect 2334 6166 2348 6222
rect 2266 6154 2348 6166
rect 2058 6054 2078 6148
rect 2124 6054 2149 6148
rect 1852 6041 1933 6051
rect 1852 5985 1863 6041
rect 1919 5985 1933 6041
rect 1852 5977 1933 5985
rect 1643 5649 1670 5743
rect 1716 5649 1734 5743
rect 1852 5804 1936 5817
rect 1852 5748 1866 5804
rect 1922 5748 1936 5804
rect 1852 5743 1936 5748
rect 1852 5740 1874 5743
rect 1643 5553 1734 5649
rect 1920 5740 1936 5743
rect 2058 5743 2149 6054
rect 2282 6148 2328 6154
rect 2282 6043 2328 6054
rect 2461 6148 2552 6287
rect 2894 6160 2940 6287
rect 3079 6222 3161 6229
rect 3079 6166 3092 6222
rect 3148 6166 3161 6222
rect 2461 6054 2486 6148
rect 2532 6054 2552 6148
rect 2260 5966 2345 5974
rect 2260 5910 2273 5966
rect 2329 5910 2345 5966
rect 2260 5902 2345 5910
rect 1874 5638 1920 5649
rect 2058 5649 2078 5743
rect 2124 5649 2149 5743
rect 2058 5553 2149 5649
rect 2282 5743 2328 5902
rect 2282 5638 2328 5649
rect 2461 5743 2552 6054
rect 2690 6148 2736 6159
rect 2690 6053 2736 6054
rect 2891 6148 2941 6160
rect 3079 6154 3161 6166
rect 3302 6161 3348 6287
rect 4178 6270 4193 6360
rect 4293 6270 4308 6360
rect 4178 6257 4308 6270
rect 4220 6177 4266 6257
rect 2891 6054 2894 6148
rect 2940 6054 2941 6148
rect 2674 6041 2754 6053
rect 2891 6042 2941 6054
rect 3098 6148 3144 6154
rect 3098 6043 3144 6054
rect 3300 6148 3349 6161
rect 4178 6160 4308 6177
rect 3300 6054 3302 6148
rect 3348 6054 3349 6148
rect 3300 6042 3349 6054
rect 3506 6148 3552 6159
rect 4178 6070 4193 6160
rect 4293 6070 4308 6160
rect 4178 6057 4308 6070
rect 2674 5985 2683 6041
rect 2739 5994 2754 6041
rect 3506 5995 3552 6054
rect 3824 5998 3906 6009
rect 3824 5995 3836 5998
rect 3506 5994 3836 5995
rect 2739 5985 3836 5994
rect 2674 5977 3836 5985
rect 2678 5949 3836 5977
rect 2678 5948 3552 5949
rect 2461 5649 2486 5743
rect 2532 5649 2552 5743
rect 2672 5802 2754 5812
rect 2672 5746 2685 5802
rect 2741 5746 2754 5802
rect 2672 5743 2754 5746
rect 2672 5735 2690 5743
rect 2461 5553 2552 5649
rect 2736 5735 2754 5743
rect 2891 5743 2942 5755
rect 2690 5638 2736 5649
rect 2891 5649 2894 5743
rect 2940 5649 2942 5743
rect 2891 5637 2942 5649
rect 3098 5743 3144 5948
rect 3824 5942 3836 5949
rect 3892 5942 3906 5998
rect 4220 5977 4266 6057
rect 3824 5933 3906 5942
rect 4178 5960 4308 5977
rect 4178 5870 4193 5960
rect 4293 5870 4308 5960
rect 4178 5857 4308 5870
rect 3488 5803 3571 5812
rect 3098 5638 3144 5649
rect 3299 5743 3350 5755
rect 3299 5649 3302 5743
rect 3348 5649 3350 5743
rect 3488 5749 3502 5803
rect 3556 5749 3571 5803
rect 4220 5777 4266 5857
rect 3488 5743 3571 5749
rect 3488 5738 3506 5743
rect 3299 5637 3350 5649
rect 3552 5738 3571 5743
rect 4178 5760 4308 5777
rect 4178 5670 4193 5760
rect 4293 5670 4308 5760
rect 4178 5657 4308 5670
rect 3506 5638 3552 5649
rect 2894 5553 2940 5637
rect 3302 5553 3348 5637
rect 4220 5577 4266 5657
rect 4178 5560 4308 5577
rect -422 5457 -292 5470
rect 80 5506 158 5517
rect 256 5506 335 5513
rect -3218 5385 -3203 5452
rect -3136 5445 -701 5452
rect -3136 5389 -2724 5445
rect -2412 5389 -1961 5445
rect -1649 5389 -1150 5445
rect -838 5389 -701 5445
rect -3136 5385 -701 5389
rect -3218 5357 -701 5385
rect -393 5377 -347 5457
rect 80 5450 92 5506
rect 148 5500 335 5506
rect 148 5450 271 5500
rect 80 5443 158 5450
rect 256 5449 271 5450
rect 322 5449 335 5500
rect 256 5434 335 5449
rect 446 5507 3357 5553
rect 446 5490 3355 5507
rect -2839 5341 -2275 5357
rect -2076 5341 -1512 5357
rect -1265 5341 -701 5357
rect -422 5360 -292 5377
rect 446 5363 492 5490
rect 641 5432 699 5434
rect 629 5425 711 5432
rect 629 5369 642 5425
rect 698 5369 711 5425
rect -2743 5198 -2692 5341
rect -2743 5124 -2740 5198
rect -2694 5124 -2692 5198
rect -2743 5122 -2692 5124
rect -2580 5198 -2534 5209
rect -2740 5113 -2694 5122
rect -2580 5071 -2534 5124
rect -2420 5198 -2374 5341
rect -2227 5226 -2149 5236
rect -2227 5172 -2215 5226
rect -2161 5222 -2149 5226
rect -2161 5176 -2031 5222
rect -2161 5172 -2149 5176
rect -2227 5160 -2149 5172
rect -2420 5113 -2374 5124
rect -2580 5067 -2471 5071
rect -2739 5053 -2650 5067
rect -2739 5025 -2725 5053
rect -2840 5023 -2725 5025
rect -2887 4994 -2725 5023
rect -2662 4994 -2650 5053
rect -2580 5025 -2275 5067
rect -2504 5021 -2275 5025
rect -2887 4991 -2650 4994
rect -3642 4979 -2650 4991
rect -3642 4931 -2790 4979
rect -2559 4953 -2474 4964
rect -2559 4931 -2548 4953
rect -3642 4917 -2548 4931
rect -2887 4912 -2548 4917
rect -2840 4894 -2548 4912
rect -2485 4894 -2474 4953
rect -2840 4885 -2474 4894
rect -2740 4828 -2694 4839
rect -2580 4838 -2534 4839
rect -2740 4674 -2694 4754
rect -2593 4828 -2526 4838
rect -2593 4754 -2580 4828
rect -2534 4754 -2526 4828
rect -2593 4740 -2526 4754
rect -2420 4828 -2374 5021
rect -2321 4814 -2275 5021
rect -2077 5025 -2031 5176
rect -1980 5198 -1929 5341
rect -1980 5124 -1977 5198
rect -1931 5124 -1929 5198
rect -1980 5122 -1929 5124
rect -1817 5198 -1771 5209
rect -1977 5113 -1931 5122
rect -1817 5071 -1771 5124
rect -1657 5198 -1611 5341
rect -1169 5198 -1118 5341
rect -1021 5270 -943 5282
rect -1021 5216 -1009 5270
rect -955 5216 -943 5270
rect -1021 5204 -943 5216
rect -1657 5113 -1611 5124
rect -1354 5174 -1271 5189
rect -1354 5120 -1340 5174
rect -1286 5120 -1271 5174
rect -1169 5124 -1166 5198
rect -1120 5124 -1118 5198
rect -1169 5122 -1118 5124
rect -1006 5198 -959 5204
rect -960 5193 -959 5198
rect -846 5198 -800 5341
rect -422 5270 -407 5360
rect -307 5270 -292 5360
rect -422 5257 -292 5270
rect 242 5351 288 5362
rect 443 5351 494 5363
rect 629 5357 711 5369
rect 854 5363 900 5490
rect 443 5257 446 5351
rect 492 5257 494 5351
rect -1354 5105 -1271 5120
rect -1166 5113 -1120 5122
rect -1817 5067 -1708 5071
rect -1976 5053 -1887 5067
rect -1976 5025 -1962 5053
rect -2077 4994 -1962 5025
rect -1899 4994 -1887 5053
rect -1817 5038 -1512 5067
rect -1817 5025 -1593 5038
rect -1741 5021 -1593 5025
rect -2077 4979 -1887 4994
rect -1657 4984 -1593 5021
rect -1539 5021 -1512 5038
rect -1336 5025 -1290 5105
rect -1006 5071 -960 5124
rect -393 5177 -347 5257
rect 228 5247 310 5257
rect 228 5191 240 5247
rect 296 5191 310 5247
rect 443 5245 494 5257
rect 650 5351 696 5357
rect 650 5246 696 5257
rect 851 5351 902 5363
rect 851 5257 854 5351
rect 900 5257 902 5351
rect 851 5245 902 5257
rect 1058 5351 1104 5362
rect 1058 5254 1104 5257
rect 1234 5351 1325 5490
rect 1450 5425 1532 5432
rect 1450 5369 1462 5425
rect 1518 5369 1532 5425
rect 1450 5357 1532 5369
rect 1234 5257 1262 5351
rect 1308 5257 1325 5351
rect 228 5182 310 5191
rect 1038 5244 1119 5254
rect 1038 5188 1051 5244
rect 1107 5188 1119 5244
rect 1038 5180 1119 5188
rect -846 5113 -800 5124
rect -422 5160 -292 5177
rect -1006 5067 -897 5071
rect -422 5070 -407 5160
rect -307 5070 -292 5160
rect 1038 5152 1096 5180
rect 650 5106 1096 5152
rect -1165 5053 -1076 5067
rect -1165 5025 -1151 5053
rect -1539 4984 -1527 5021
rect -1657 4978 -1527 4984
rect -1336 4994 -1151 5025
rect -1088 4994 -1076 5053
rect -1006 5043 -670 5067
rect -422 5057 -292 5070
rect -94 5095 -11 5101
rect 131 5095 210 5106
rect -1006 5025 -551 5043
rect -930 5021 -551 5025
rect -1336 4979 -1076 4994
rect -1796 4953 -1711 4964
rect -2098 4931 -2028 4933
rect -1796 4931 -1785 4953
rect -2098 4920 -1785 4931
rect -2098 4864 -2088 4920
rect -2032 4894 -1785 4920
rect -1722 4894 -1711 4953
rect -2032 4885 -1711 4894
rect -1657 4931 -1611 4978
rect -985 4953 -900 4964
rect -985 4931 -974 4953
rect -1657 4894 -974 4931
rect -911 4894 -900 4953
rect -1657 4885 -900 4894
rect -2032 4864 -2028 4885
rect -2098 4852 -2028 4864
rect -1977 4828 -1931 4839
rect -1817 4838 -1771 4839
rect -2321 4805 -2218 4814
rect -2321 4755 -2284 4805
rect -2420 4743 -2374 4754
rect -2296 4751 -2284 4755
rect -2230 4751 -2218 4805
rect -2296 4742 -2218 4751
rect -1977 4674 -1931 4754
rect -1830 4828 -1763 4838
rect -1830 4754 -1817 4828
rect -1771 4754 -1763 4828
rect -1830 4740 -1763 4754
rect -1657 4828 -1611 4885
rect -1657 4743 -1611 4754
rect -1166 4828 -1120 4839
rect -1006 4838 -960 4839
rect -1166 4674 -1120 4754
rect -1019 4828 -952 4838
rect -1019 4754 -1006 4828
rect -960 4754 -952 4828
rect -1019 4740 -952 4754
rect -846 4828 -800 5021
rect -716 5015 -551 5021
rect -716 4965 -617 5015
rect -630 4961 -617 4965
rect -563 4961 -551 5015
rect -393 4977 -347 5057
rect -94 5039 -79 5095
rect -23 5092 210 5095
rect -23 5041 145 5092
rect 196 5041 210 5092
rect 523 5067 597 5079
rect 523 5062 533 5067
rect -23 5039 210 5041
rect -94 5029 -11 5039
rect 131 5027 210 5039
rect 326 5016 533 5062
rect -630 4954 -551 4961
rect -422 4960 -292 4977
rect -422 4870 -407 4960
rect -307 4870 -292 4960
rect 326 4958 372 5016
rect 523 5011 533 5016
rect 589 5011 597 5067
rect 523 4999 597 5011
rect -422 4857 -292 4870
rect 239 4946 372 4958
rect -393 4777 -347 4857
rect 239 4852 242 4946
rect 288 4887 372 4946
rect 443 4946 494 4958
rect 288 4852 290 4887
rect -245 4838 -173 4852
rect 239 4840 290 4852
rect 443 4852 446 4946
rect 492 4852 494 4946
rect 443 4840 494 4852
rect 650 4946 696 5106
rect 1042 5009 1124 5017
rect 650 4841 696 4852
rect 851 4946 902 4958
rect 851 4852 854 4946
rect 900 4852 902 4946
rect 1042 4953 1057 5009
rect 1113 4953 1124 5009
rect 1042 4946 1124 4953
rect 1042 4945 1058 4946
rect 851 4840 902 4852
rect 1104 4945 1124 4946
rect 1234 4946 1325 5257
rect 1466 5351 1512 5357
rect 1466 5246 1512 5257
rect 1643 5351 1734 5490
rect 1643 5257 1670 5351
rect 1716 5257 1734 5351
rect 1445 5174 1530 5189
rect 1445 5118 1458 5174
rect 1514 5118 1530 5174
rect 1445 5108 1530 5118
rect 1058 4841 1104 4852
rect 1234 4852 1262 4946
rect 1308 4852 1325 4946
rect -245 4782 -238 4838
rect -182 4782 128 4838
rect -846 4743 -800 4754
rect -422 4760 -292 4777
rect -245 4770 -173 4782
rect -2863 4665 -2247 4674
rect -2100 4665 -1484 4674
rect -1289 4665 -673 4674
rect -3024 4658 -2943 4665
rect -2863 4658 -673 4665
rect -3024 4657 -673 4658
rect -422 4670 -407 4760
rect -307 4670 -292 4760
rect -422 4657 -292 4670
rect 72 4721 128 4782
rect 446 4756 492 4840
rect 854 4756 900 4840
rect 1234 4756 1325 4852
rect 1466 4946 1512 5108
rect 1466 4841 1512 4852
rect 1643 4946 1734 5257
rect 1874 5351 1920 5362
rect 1874 5254 1920 5257
rect 2058 5351 2149 5490
rect 2266 5425 2348 5432
rect 2266 5369 2278 5425
rect 2334 5369 2348 5425
rect 2266 5357 2348 5369
rect 2058 5257 2078 5351
rect 2124 5257 2149 5351
rect 1852 5244 1933 5254
rect 1852 5188 1863 5244
rect 1919 5188 1933 5244
rect 1852 5180 1933 5188
rect 1643 4852 1670 4946
rect 1716 4852 1734 4946
rect 1852 5007 1936 5020
rect 1852 4951 1866 5007
rect 1922 4951 1936 5007
rect 1852 4946 1936 4951
rect 1852 4943 1874 4946
rect 1643 4756 1734 4852
rect 1920 4943 1936 4946
rect 2058 4946 2149 5257
rect 2282 5351 2328 5357
rect 2282 5246 2328 5257
rect 2461 5351 2552 5490
rect 2894 5363 2940 5490
rect 3079 5425 3161 5432
rect 3079 5369 3092 5425
rect 3148 5369 3161 5425
rect 2461 5257 2486 5351
rect 2532 5257 2552 5351
rect 2260 5169 2345 5177
rect 2260 5113 2273 5169
rect 2329 5113 2345 5169
rect 2260 5105 2345 5113
rect 1874 4841 1920 4852
rect 2058 4852 2078 4946
rect 2124 4852 2149 4946
rect 2058 4756 2149 4852
rect 2282 4946 2328 5105
rect 2282 4841 2328 4852
rect 2461 4946 2552 5257
rect 2690 5351 2736 5362
rect 2690 5256 2736 5257
rect 2891 5351 2941 5363
rect 3079 5357 3161 5369
rect 3302 5364 3348 5490
rect 4178 5470 4193 5560
rect 4293 5470 4308 5560
rect 4178 5457 4308 5470
rect 4220 5377 4266 5457
rect 2891 5257 2894 5351
rect 2940 5257 2941 5351
rect 2674 5244 2754 5256
rect 2891 5245 2941 5257
rect 3098 5351 3144 5357
rect 3098 5246 3144 5257
rect 3300 5351 3349 5364
rect 3300 5257 3302 5351
rect 3348 5257 3349 5351
rect 3300 5245 3349 5257
rect 3506 5351 3552 5362
rect 4178 5360 4308 5377
rect 4178 5270 4193 5360
rect 4293 5270 4308 5360
rect 4178 5257 4308 5270
rect 2674 5188 2683 5244
rect 2739 5197 2754 5244
rect 3506 5198 3552 5257
rect 3822 5200 3904 5213
rect 3822 5198 3836 5200
rect 3495 5197 3836 5198
rect 2739 5188 3836 5197
rect 2674 5180 3836 5188
rect 2678 5152 3836 5180
rect 2678 5151 3552 5152
rect 2461 4852 2486 4946
rect 2532 4852 2552 4946
rect 2672 5005 2754 5015
rect 2672 4949 2685 5005
rect 2741 4949 2754 5005
rect 2672 4946 2754 4949
rect 2672 4938 2690 4946
rect 2461 4756 2552 4852
rect 2736 4938 2754 4946
rect 2891 4946 2942 4958
rect 2690 4841 2736 4852
rect 2891 4852 2894 4946
rect 2940 4852 2942 4946
rect 2891 4840 2942 4852
rect 3098 4946 3144 5151
rect 3822 5144 3836 5152
rect 3892 5144 3904 5200
rect 4220 5177 4266 5257
rect 3822 5137 3904 5144
rect 4178 5160 4308 5177
rect 4178 5070 4193 5160
rect 4293 5070 4308 5160
rect 4178 5057 4308 5070
rect 3488 5006 3571 5015
rect 3098 4841 3144 4852
rect 3299 4946 3350 4958
rect 3299 4852 3302 4946
rect 3348 4852 3350 4946
rect 3488 4952 3502 5006
rect 3556 4952 3571 5006
rect 4220 4977 4266 5057
rect 3488 4946 3571 4952
rect 3488 4941 3506 4946
rect 3299 4840 3350 4852
rect 3552 4941 3571 4946
rect 4178 4960 4308 4977
rect 4178 4870 4193 4960
rect 4293 4870 4308 4960
rect 4178 4857 4308 4870
rect 3506 4841 3552 4852
rect 2894 4756 2940 4840
rect 3302 4756 3348 4840
rect 4220 4777 4266 4857
rect 4178 4760 4308 4777
rect 72 4711 156 4721
rect 256 4711 335 4716
rect -3024 4592 -3012 4657
rect -2947 4647 -673 4657
rect -2947 4599 -2796 4647
rect -2327 4599 -2033 4647
rect -1564 4599 -1222 4647
rect -753 4599 -673 4647
rect -2947 4598 -673 4599
rect -2947 4592 -2247 4598
rect -3024 4591 -2247 4592
rect -3024 4587 -2943 4591
rect -2863 4576 -2247 4591
rect -2100 4576 -1484 4598
rect -1289 4576 -673 4598
rect -393 4577 -347 4657
rect 72 4655 92 4711
rect 148 4703 335 4711
rect 148 4655 271 4703
rect 72 4652 156 4655
rect 78 4647 156 4652
rect 256 4652 271 4655
rect 322 4652 335 4703
rect 256 4637 335 4652
rect 446 4710 3357 4756
rect 446 4693 3355 4710
rect -422 4560 -292 4577
rect 446 4566 492 4693
rect 641 4635 699 4637
rect 629 4628 711 4635
rect 629 4572 642 4628
rect 698 4572 711 4628
rect -2839 4484 -2275 4516
rect -2076 4484 -1512 4515
rect -1265 4484 -701 4515
rect -3213 4470 -701 4484
rect -3213 4444 -2724 4470
rect -3213 4376 -3203 4444
rect -3136 4414 -2724 4444
rect -2412 4469 -701 4470
rect -2412 4414 -1961 4469
rect -3136 4413 -1961 4414
rect -1649 4413 -1150 4469
rect -838 4413 -701 4469
rect -422 4470 -407 4560
rect -307 4470 -292 4560
rect -422 4457 -292 4470
rect 242 4554 288 4565
rect 443 4554 494 4566
rect 629 4560 711 4572
rect 854 4566 900 4693
rect 443 4460 446 4554
rect 492 4460 494 4554
rect -3136 4376 -701 4413
rect -393 4377 -347 4457
rect 228 4450 310 4460
rect 228 4394 240 4450
rect 296 4394 310 4450
rect 443 4448 494 4460
rect 650 4554 696 4560
rect 650 4449 696 4460
rect 851 4554 902 4566
rect 851 4460 854 4554
rect 900 4460 902 4554
rect 851 4448 902 4460
rect 1058 4554 1104 4565
rect 1058 4457 1104 4460
rect 1234 4554 1325 4693
rect 1450 4628 1532 4635
rect 1450 4572 1462 4628
rect 1518 4572 1532 4628
rect 1450 4560 1532 4572
rect 1234 4460 1262 4554
rect 1308 4460 1325 4554
rect 228 4385 310 4394
rect 1038 4447 1119 4457
rect 1038 4391 1051 4447
rect 1107 4391 1119 4447
rect 1038 4383 1119 4391
rect -3213 4369 -701 4376
rect -3213 4368 -3122 4369
rect -3213 4364 -3124 4368
rect -2839 4366 -2275 4369
rect -2743 4223 -2692 4366
rect -2743 4149 -2740 4223
rect -2694 4149 -2692 4223
rect -2743 4147 -2692 4149
rect -2580 4223 -2534 4234
rect -2740 4138 -2694 4147
rect -2580 4096 -2534 4149
rect -2420 4223 -2374 4366
rect -2076 4365 -1512 4369
rect -1265 4365 -701 4369
rect -2420 4138 -2374 4149
rect -1980 4222 -1929 4365
rect -1980 4148 -1977 4222
rect -1931 4148 -1929 4222
rect -1980 4146 -1929 4148
rect -1817 4222 -1771 4233
rect -1977 4137 -1931 4146
rect -2165 4115 -2090 4127
rect -2580 4092 -2471 4096
rect -2739 4078 -2650 4092
rect -2739 4050 -2725 4078
rect -2840 4019 -2725 4050
rect -2662 4019 -2650 4078
rect -2580 4050 -2275 4092
rect -2504 4046 -2275 4050
rect -2165 4061 -2156 4115
rect -2102 4061 -2090 4115
rect -1817 4095 -1771 4148
rect -1657 4222 -1611 4365
rect -1657 4137 -1611 4148
rect -1169 4222 -1118 4365
rect -1169 4148 -1166 4222
rect -1120 4148 -1118 4222
rect -1169 4146 -1118 4148
rect -1006 4222 -960 4233
rect -1166 4137 -1120 4146
rect -1006 4095 -960 4148
rect -846 4222 -800 4365
rect -422 4360 -292 4377
rect -422 4270 -407 4360
rect -307 4270 -292 4360
rect 1038 4355 1096 4383
rect 650 4309 1096 4355
rect -422 4257 -292 4270
rect -92 4293 -10 4300
rect 131 4295 210 4309
rect 131 4293 145 4295
rect -393 4177 -347 4257
rect -92 4237 -79 4293
rect -23 4244 145 4293
rect 196 4244 210 4295
rect 523 4270 597 4282
rect 523 4265 533 4270
rect -23 4237 210 4244
rect -92 4228 -10 4237
rect 131 4230 210 4237
rect 326 4219 533 4265
rect -846 4137 -800 4148
rect -422 4160 -292 4177
rect 326 4161 372 4219
rect 523 4214 533 4219
rect 589 4214 597 4270
rect 523 4202 597 4214
rect -1817 4091 -1708 4095
rect -1006 4091 -897 4095
rect -2165 4049 -2090 4061
rect -1976 4077 -1887 4091
rect -1976 4049 -1962 4077
rect -3573 4004 -2650 4019
rect -3573 3956 -2794 4004
rect -2559 3978 -2474 3989
rect -2559 3956 -2548 3978
rect -3573 3941 -2548 3956
rect -2840 3919 -2548 3941
rect -2485 3919 -2474 3978
rect -2840 3910 -2474 3919
rect -2740 3853 -2694 3864
rect -2580 3863 -2534 3864
rect -2740 3699 -2694 3779
rect -2593 3853 -2526 3863
rect -2593 3779 -2580 3853
rect -2534 3779 -2526 3853
rect -2593 3765 -2526 3779
rect -2420 3853 -2374 4046
rect -2321 3955 -2275 4046
rect -2152 4018 -1962 4049
rect -1899 4018 -1887 4077
rect -1817 4064 -1512 4091
rect -1817 4049 -1594 4064
rect -1741 4045 -1594 4049
rect -2152 4003 -1887 4018
rect -1657 4010 -1594 4045
rect -1540 4045 -1512 4064
rect -1165 4077 -1076 4091
rect -1165 4049 -1151 4077
rect -1540 4010 -1528 4045
rect -1657 3997 -1528 4010
rect -1266 4018 -1151 4049
rect -1088 4018 -1076 4077
rect -1006 4056 -701 4091
rect -422 4070 -407 4160
rect -307 4070 -292 4160
rect -422 4057 -292 4070
rect 239 4149 372 4161
rect -1006 4049 -789 4056
rect -930 4045 -789 4049
rect -1266 4003 -1076 4018
rect -1796 3977 -1711 3988
rect -1796 3955 -1785 3977
rect -2321 3918 -1785 3955
rect -1722 3918 -1711 3977
rect -2321 3909 -1711 3918
rect -2420 3768 -2374 3779
rect -1977 3852 -1931 3863
rect -1817 3862 -1771 3863
rect -3025 3687 -2932 3697
rect -2863 3687 -2247 3699
rect -1977 3698 -1931 3778
rect -1830 3852 -1763 3862
rect -1830 3778 -1817 3852
rect -1771 3778 -1763 3852
rect -1830 3764 -1763 3778
rect -1657 3852 -1611 3997
rect -1266 3981 -1220 4003
rect -846 4002 -789 4045
rect -735 4045 -701 4056
rect -735 4002 -725 4045
rect -846 3990 -725 4002
rect -1328 3974 -1220 3981
rect -1328 3920 -1315 3974
rect -1261 3955 -1220 3974
rect -985 3977 -900 3988
rect -985 3955 -974 3977
rect -1261 3920 -974 3955
rect -1328 3918 -974 3920
rect -911 3918 -900 3977
rect -1328 3909 -900 3918
rect -1328 3906 -1259 3909
rect -1657 3767 -1611 3778
rect -1166 3852 -1120 3863
rect -1006 3862 -960 3863
rect -1166 3698 -1120 3778
rect -1019 3852 -952 3862
rect -1019 3778 -1006 3852
rect -960 3778 -952 3852
rect -1019 3764 -952 3778
rect -846 3852 -800 3990
rect -393 3977 -347 4057
rect 239 4055 242 4149
rect 288 4090 372 4149
rect 443 4149 494 4161
rect 288 4055 290 4090
rect 239 4043 290 4055
rect 443 4055 446 4149
rect 492 4055 494 4149
rect 443 4043 494 4055
rect 650 4149 696 4309
rect 1042 4212 1124 4220
rect 650 4044 696 4055
rect 851 4149 902 4161
rect 851 4055 854 4149
rect 900 4055 902 4149
rect 1042 4156 1057 4212
rect 1113 4156 1124 4212
rect 1042 4149 1124 4156
rect 1042 4148 1058 4149
rect 851 4043 902 4055
rect 1104 4148 1124 4149
rect 1234 4149 1325 4460
rect 1466 4554 1512 4560
rect 1466 4449 1512 4460
rect 1643 4554 1734 4693
rect 1643 4460 1670 4554
rect 1716 4460 1734 4554
rect 1445 4377 1530 4392
rect 1445 4321 1458 4377
rect 1514 4321 1530 4377
rect 1445 4311 1530 4321
rect 1058 4044 1104 4055
rect 1234 4055 1262 4149
rect 1308 4055 1325 4149
rect 446 3982 492 4043
rect 854 3982 900 4043
rect 1234 3982 1325 4055
rect 1466 4149 1512 4311
rect 1466 4044 1512 4055
rect 1643 4149 1734 4460
rect 1874 4554 1920 4565
rect 1874 4457 1920 4460
rect 2058 4554 2149 4693
rect 2266 4628 2348 4635
rect 2266 4572 2278 4628
rect 2334 4572 2348 4628
rect 2266 4560 2348 4572
rect 2058 4460 2078 4554
rect 2124 4460 2149 4554
rect 1852 4447 1933 4457
rect 1852 4391 1863 4447
rect 1919 4391 1933 4447
rect 1852 4383 1933 4391
rect 1643 4055 1670 4149
rect 1716 4055 1734 4149
rect 1852 4210 1936 4223
rect 1852 4154 1866 4210
rect 1922 4154 1936 4210
rect 1852 4149 1936 4154
rect 1852 4146 1874 4149
rect 1643 3982 1734 4055
rect 1920 4146 1936 4149
rect 2058 4149 2149 4460
rect 2282 4554 2328 4560
rect 2282 4449 2328 4460
rect 2461 4554 2552 4693
rect 2894 4566 2940 4693
rect 3079 4628 3161 4635
rect 3079 4572 3092 4628
rect 3148 4572 3161 4628
rect 2461 4460 2486 4554
rect 2532 4460 2552 4554
rect 2260 4372 2345 4380
rect 2260 4316 2273 4372
rect 2329 4316 2345 4372
rect 2260 4308 2345 4316
rect 1874 4044 1920 4055
rect 2058 4055 2078 4149
rect 2124 4055 2149 4149
rect 2058 3982 2149 4055
rect 2282 4149 2328 4308
rect 2282 4044 2328 4055
rect 2461 4149 2552 4460
rect 2690 4554 2736 4565
rect 2690 4459 2736 4460
rect 2891 4554 2941 4566
rect 3079 4560 3161 4572
rect 3302 4567 3348 4693
rect 4178 4670 4193 4760
rect 4293 4670 4308 4760
rect 4178 4657 4308 4670
rect 4220 4577 4266 4657
rect 2891 4460 2894 4554
rect 2940 4460 2941 4554
rect 2674 4447 2754 4459
rect 2891 4448 2941 4460
rect 3098 4554 3144 4560
rect 3098 4449 3144 4460
rect 3300 4554 3349 4567
rect 3300 4460 3302 4554
rect 3348 4460 3349 4554
rect 3300 4448 3349 4460
rect 3506 4554 3552 4565
rect 2674 4391 2683 4447
rect 2739 4400 2754 4447
rect 3506 4401 3552 4460
rect 4178 4560 4308 4577
rect 4178 4470 4193 4560
rect 4293 4470 4308 4560
rect 4178 4457 4308 4470
rect 3826 4402 3908 4413
rect 3826 4401 3836 4402
rect 3506 4400 3836 4401
rect 2739 4391 3836 4400
rect 2674 4383 3836 4391
rect 2678 4355 3836 4383
rect 2678 4354 3552 4355
rect 2461 4055 2486 4149
rect 2532 4055 2552 4149
rect 2672 4208 2754 4218
rect 2672 4152 2685 4208
rect 2741 4152 2754 4208
rect 2672 4149 2754 4152
rect 2672 4141 2690 4149
rect 2461 3982 2552 4055
rect 2736 4141 2754 4149
rect 2891 4149 2942 4161
rect 2690 4044 2736 4055
rect 2891 4055 2894 4149
rect 2940 4055 2942 4149
rect 2891 4043 2942 4055
rect 3098 4149 3144 4354
rect 3826 4346 3836 4355
rect 3892 4346 3908 4402
rect 4220 4377 4266 4457
rect 3826 4337 3908 4346
rect 4178 4360 4308 4377
rect 4178 4270 4193 4360
rect 4293 4270 4308 4360
rect 4178 4257 4308 4270
rect 3488 4209 3571 4218
rect 3098 4044 3144 4055
rect 3299 4149 3350 4161
rect 3299 4055 3302 4149
rect 3348 4055 3350 4149
rect 3488 4155 3502 4209
rect 3556 4155 3571 4209
rect 4220 4177 4266 4257
rect 3488 4149 3571 4155
rect 3488 4144 3506 4149
rect 3299 4043 3350 4055
rect 3552 4144 3571 4149
rect 4178 4160 4308 4177
rect 4178 4070 4193 4160
rect 4293 4070 4308 4160
rect 4178 4057 4308 4070
rect 3506 4044 3552 4055
rect 2894 3982 2940 4043
rect 3302 3982 3348 4043
rect 3618 4020 4015 4037
rect 3618 3982 3790 4020
rect -422 3960 -292 3977
rect -422 3870 -407 3960
rect -307 3870 -292 3960
rect 75 3963 167 3981
rect 75 3907 92 3963
rect 148 3907 167 3963
rect 446 3966 3790 3982
rect 3844 3966 4015 4020
rect 4220 3977 4266 4057
rect 446 3952 4015 3966
rect 446 3913 3657 3952
rect 75 3889 167 3907
rect 451 3898 3657 3913
rect 3711 3943 4015 3952
rect 3711 3898 3917 3943
rect 451 3891 3917 3898
rect 3618 3889 3917 3891
rect 3971 3889 4015 3943
rect 3618 3870 4015 3889
rect 4178 3960 4308 3977
rect 4178 3870 4193 3960
rect 4293 3870 4308 3960
rect -422 3857 -292 3870
rect 4178 3857 4308 3870
rect -846 3767 -800 3778
rect -393 3777 -347 3857
rect 4220 3777 4266 3857
rect -422 3760 -292 3777
rect -422 3698 -407 3760
rect -2100 3687 -1484 3698
rect -1289 3687 -407 3698
rect -3538 3620 -3013 3687
rect -2946 3672 -407 3687
rect -2946 3624 -2796 3672
rect -2327 3671 -407 3672
rect -2327 3624 -2033 3671
rect -2946 3623 -2033 3624
rect -1564 3623 -1222 3671
rect -753 3670 -407 3671
rect -307 3743 -292 3760
rect -222 3760 -92 3777
rect -222 3743 -207 3760
rect -307 3670 -207 3743
rect -107 3743 -92 3760
rect -22 3760 108 3777
rect -22 3743 -7 3760
rect -107 3670 -7 3743
rect 93 3743 108 3760
rect 178 3760 308 3777
rect 178 3743 193 3760
rect 93 3670 193 3743
rect 293 3743 308 3760
rect 378 3760 508 3777
rect 378 3743 393 3760
rect 293 3670 393 3743
rect 493 3743 508 3760
rect 578 3760 708 3777
rect 578 3743 593 3760
rect 493 3670 593 3743
rect 693 3743 708 3760
rect 778 3760 908 3777
rect 778 3743 793 3760
rect 693 3670 793 3743
rect 893 3743 908 3760
rect 978 3760 1108 3777
rect 978 3743 993 3760
rect 893 3670 993 3743
rect 1093 3743 1108 3760
rect 1178 3760 1308 3777
rect 1178 3743 1193 3760
rect 1093 3670 1193 3743
rect 1293 3743 1308 3760
rect 1378 3760 1508 3777
rect 1378 3743 1393 3760
rect 1293 3670 1393 3743
rect 1493 3743 1508 3760
rect 1578 3760 1708 3777
rect 1578 3743 1593 3760
rect 1493 3670 1593 3743
rect 1693 3743 1708 3760
rect 1778 3760 1908 3777
rect 1778 3743 1793 3760
rect 1693 3670 1793 3743
rect 1893 3743 1908 3760
rect 1978 3760 2108 3777
rect 1978 3743 1993 3760
rect 1893 3670 1993 3743
rect 2093 3743 2108 3760
rect 2178 3760 2308 3777
rect 2178 3743 2193 3760
rect 2093 3670 2193 3743
rect 2293 3743 2308 3760
rect 2378 3760 2508 3777
rect 2378 3743 2393 3760
rect 2293 3670 2393 3743
rect 2493 3743 2508 3760
rect 2578 3760 2708 3777
rect 2578 3743 2593 3760
rect 2493 3670 2593 3743
rect 2693 3743 2708 3760
rect 2778 3760 2908 3777
rect 2778 3743 2793 3760
rect 2693 3670 2793 3743
rect 2893 3743 2908 3760
rect 2978 3760 3108 3777
rect 2978 3743 2993 3760
rect 2893 3670 2993 3743
rect 3093 3743 3108 3760
rect 3178 3760 3308 3777
rect 3178 3743 3193 3760
rect 3093 3670 3193 3743
rect 3293 3743 3308 3760
rect 3378 3760 3508 3777
rect 3378 3743 3393 3760
rect 3293 3670 3393 3743
rect 3493 3743 3508 3760
rect 3578 3760 3708 3777
rect 3578 3743 3593 3760
rect 3493 3670 3593 3743
rect 3693 3743 3708 3760
rect 3778 3760 3908 3777
rect 3778 3743 3793 3760
rect 3693 3670 3793 3743
rect 3893 3743 3908 3760
rect 3978 3760 4108 3777
rect 3978 3743 3993 3760
rect 3893 3697 3993 3743
rect 3893 3670 3908 3697
rect -753 3657 3908 3670
rect 3978 3670 3993 3697
rect 4093 3743 4108 3760
rect 4178 3760 4308 3777
rect 4178 3743 4193 3760
rect 4093 3697 4193 3743
rect 4093 3670 4108 3697
rect 3978 3657 4108 3670
rect 4178 3670 4193 3697
rect 4293 3670 4308 3760
rect 4178 3657 4308 3670
rect -753 3623 3879 3657
rect -2946 3620 3879 3623
rect -3538 3570 3879 3620
rect -2784 3463 3879 3570
rect -2839 3450 3879 3463
rect 4031 3524 4129 3540
rect 4031 3454 4046 3524
rect 4116 3454 4129 3524
rect -2839 3437 3876 3450
rect 4031 3444 4129 3454
rect -2839 3306 -2791 3437
rect -2646 3306 -2491 3437
rect -2346 3306 -2191 3437
rect -2046 3306 -1891 3437
rect -1746 3306 -1591 3437
rect -1446 3306 -1291 3437
rect -1146 3306 -991 3437
rect -846 3306 -691 3437
rect -546 3306 -391 3437
rect -246 3306 -91 3437
rect 54 3306 209 3437
rect 354 3306 509 3437
rect 654 3306 809 3437
rect 954 3306 1109 3437
rect 1254 3306 1409 3437
rect 1554 3306 1709 3437
rect 1854 3306 2009 3437
rect 2154 3306 2309 3437
rect 2454 3306 2609 3437
rect 2754 3306 2909 3437
rect 3054 3306 3209 3437
rect 3354 3306 3509 3437
rect 3654 3408 3876 3437
rect 3654 3336 3728 3408
rect 3817 3336 3876 3408
rect 3654 3306 3876 3336
rect -2839 3276 3876 3306
rect -3007 3264 -2921 3269
rect -3538 3254 -2921 3264
rect -3538 3198 -2994 3254
rect -2938 3198 -2921 3254
rect -3538 3196 -2921 3198
rect -3007 3186 -2921 3196
rect -2802 3057 -2756 3068
rect -2598 3057 -2552 3068
rect -2620 3004 -2598 3021
rect -2394 3057 -2348 3276
rect -2552 3004 -2535 3021
rect -2620 2944 -2606 3004
rect -2549 2944 -2535 3004
rect -2620 2930 -2598 2944
rect -2802 2769 -2756 2843
rect -2552 2930 -2535 2944
rect -2598 2832 -2552 2843
rect -2190 3057 -2144 3068
rect -2207 3008 -2190 3022
rect -1986 3057 -1940 3068
rect -2144 3008 -2122 3022
rect -2207 2949 -2192 3008
rect -2137 2949 -2122 3008
rect -2207 2931 -2190 2949
rect -2394 2832 -2348 2843
rect -2144 2931 -2122 2949
rect -2190 2832 -2144 2843
rect -1782 3057 -1736 3068
rect -1795 2926 -1782 3016
rect -1578 3057 -1532 3276
rect -1736 3002 -1710 3016
rect -1725 2943 -1710 3002
rect -1986 2769 -1940 2843
rect -1736 2926 -1710 2943
rect -1782 2832 -1736 2843
rect -1374 3057 -1328 3068
rect -1395 3008 -1374 3022
rect -1170 3057 -1124 3068
rect -1328 3008 -1310 3022
rect -1395 2949 -1380 3008
rect -1325 2949 -1310 3008
rect -1395 2931 -1374 2949
rect -1578 2832 -1532 2843
rect -1328 2931 -1310 2949
rect -1374 2832 -1328 2843
rect -966 3057 -920 3068
rect -982 2990 -966 3004
rect -762 3057 -716 3276
rect -920 2990 -897 3004
rect -982 2931 -967 2990
rect -912 2931 -897 2990
rect -982 2913 -966 2931
rect -1170 2769 -1124 2843
rect -920 2913 -897 2931
rect -966 2832 -920 2843
rect -558 3057 -512 3068
rect -572 2924 -558 3015
rect -354 3057 -308 3068
rect -512 3001 -487 3015
rect -502 2942 -487 3001
rect -762 2832 -716 2843
rect -512 2924 -487 2942
rect -558 2832 -512 2843
rect -150 3057 -104 3068
rect -175 2990 -150 3004
rect 54 3057 100 3276
rect -175 2931 -160 2990
rect -175 2913 -150 2931
rect -354 2769 -308 2843
rect -104 2913 -90 3004
rect -150 2832 -104 2843
rect 258 3057 304 3068
rect 240 2995 258 3009
rect 462 3057 508 3068
rect 304 2995 325 3009
rect 240 2936 255 2995
rect 310 2936 325 2995
rect 240 2918 258 2936
rect 54 2832 100 2843
rect 304 2918 325 2936
rect 258 2832 304 2843
rect 666 3057 712 3068
rect 651 2921 666 3012
rect 870 3057 916 3276
rect 712 2998 736 3012
rect 721 2939 736 2998
rect 462 2769 508 2843
rect 712 2921 736 2939
rect 666 2832 712 2843
rect 1074 3057 1120 3068
rect 1061 2931 1074 3022
rect 1278 3057 1324 3068
rect 1120 3008 1146 3022
rect 1131 2949 1146 3008
rect 870 2832 916 2843
rect 1120 2931 1146 2949
rect 1074 2832 1120 2843
rect 1482 3057 1528 3068
rect 1466 2990 1482 3004
rect 1686 3057 1732 3276
rect 1528 2990 1551 3004
rect 1466 2931 1481 2990
rect 1536 2931 1551 2990
rect 1466 2913 1482 2931
rect 1278 2769 1324 2843
rect 1528 2913 1551 2931
rect 1482 2832 1528 2843
rect 1890 3057 1936 3068
rect 1868 2990 1890 3004
rect 2094 3057 2140 3068
rect 1936 2990 1953 3004
rect 1868 2931 1883 2990
rect 1938 2931 1953 2990
rect 1868 2913 1890 2931
rect 1686 2832 1732 2843
rect 1936 2913 1953 2931
rect 1890 2832 1936 2843
rect 2298 3057 2344 3068
rect 2284 2926 2298 3017
rect 2502 3057 2548 3276
rect 2344 3003 2369 3017
rect 2354 2944 2369 3003
rect 2094 2769 2140 2843
rect 2344 2926 2369 2944
rect 2298 2832 2344 2843
rect 2706 3057 2752 3068
rect 2684 2995 2706 3009
rect 2910 3057 2956 3068
rect 2752 2995 2769 3009
rect 2684 2936 2699 2995
rect 2754 2936 2769 2995
rect 2684 2918 2706 2936
rect 2502 2832 2548 2843
rect 2752 2918 2769 2936
rect 2706 2832 2752 2843
rect 3114 3057 3160 3068
rect 3101 2915 3114 3006
rect 3318 3057 3364 3276
rect 3160 2992 3186 3006
rect 3171 2933 3186 2992
rect 2910 2769 2956 2843
rect 3160 2915 3186 2933
rect 3114 2832 3160 2843
rect 3522 3057 3568 3068
rect 3489 2998 3522 3012
rect 3726 3057 3772 3068
rect 3489 2939 3504 2998
rect 3489 2921 3522 2939
rect 3318 2832 3364 2843
rect 3568 2921 3574 3012
rect 3522 2832 3568 2843
rect 3726 2769 3772 2843
rect 4045 2769 4117 3444
rect -3010 2737 -2923 2744
rect -3513 2730 -2923 2737
rect -3513 2677 -2997 2730
rect -2941 2677 -2923 2730
rect -2802 2697 4117 2769
rect -3513 2663 -2923 2677
rect -3513 2660 -2931 2663
rect -2802 2566 -2756 2577
rect -2598 2566 -2552 2577
rect -2618 2499 -2598 2516
rect -2394 2566 -2348 2697
rect -2552 2499 -2533 2516
rect -2618 2440 -2604 2499
rect -2549 2440 -2533 2499
rect -2618 2425 -2598 2440
rect -3005 2236 -2913 2252
rect -3005 2179 -2990 2236
rect -2933 2179 -2913 2236
rect -3005 2164 -2913 2179
rect -2802 2157 -2756 2352
rect -2552 2425 -2533 2440
rect -2598 2341 -2552 2352
rect -2190 2566 -2144 2577
rect -2197 2427 -2190 2518
rect -1986 2566 -1940 2577
rect -2144 2504 -2112 2518
rect -2127 2445 -2112 2504
rect -2394 2341 -2348 2352
rect -2144 2427 -2112 2445
rect -2190 2341 -2144 2352
rect -1782 2566 -1736 2577
rect -1801 2520 -1782 2534
rect -1578 2566 -1532 2697
rect -1736 2520 -1716 2534
rect -1801 2461 -1786 2520
rect -1731 2461 -1716 2520
rect -1801 2443 -1782 2461
rect -1986 2157 -1940 2352
rect -1736 2443 -1716 2461
rect -1782 2341 -1736 2352
rect -1374 2566 -1328 2577
rect -1388 2448 -1374 2539
rect -1170 2566 -1124 2577
rect -1328 2525 -1303 2539
rect -1318 2466 -1303 2525
rect -1578 2341 -1532 2352
rect -1328 2448 -1303 2466
rect -1374 2341 -1328 2352
rect -966 2566 -920 2577
rect -988 2523 -966 2537
rect -762 2566 -716 2697
rect -920 2523 -903 2537
rect -988 2464 -973 2523
rect -918 2464 -903 2523
rect -988 2446 -966 2464
rect -1170 2157 -1124 2352
rect -920 2446 -903 2464
rect -966 2341 -920 2352
rect -558 2566 -512 2577
rect -585 2513 -558 2527
rect -354 2566 -308 2577
rect -585 2454 -570 2513
rect -585 2436 -558 2454
rect -762 2341 -716 2352
rect -512 2436 -500 2527
rect -558 2341 -512 2352
rect -150 2566 -104 2577
rect -162 2438 -150 2529
rect 54 2566 100 2697
rect -104 2515 -77 2529
rect -92 2456 -77 2515
rect -354 2157 -308 2352
rect -104 2438 -77 2456
rect -150 2341 -104 2352
rect 258 2566 304 2577
rect 238 2499 258 2513
rect 462 2566 508 2577
rect 304 2499 323 2513
rect 238 2440 253 2499
rect 308 2440 323 2499
rect 238 2422 258 2440
rect 54 2341 100 2352
rect 304 2422 323 2440
rect 258 2341 304 2352
rect 666 2566 712 2577
rect 647 2514 666 2516
rect 640 2500 666 2514
rect 870 2566 916 2697
rect 712 2514 723 2516
rect 640 2441 655 2500
rect 640 2423 666 2441
rect 462 2157 508 2352
rect 712 2423 725 2514
rect 666 2341 712 2352
rect 1074 2566 1120 2577
rect 1053 2515 1074 2529
rect 1278 2566 1324 2577
rect 1120 2515 1138 2529
rect 1053 2456 1068 2515
rect 1123 2456 1138 2515
rect 1053 2438 1074 2456
rect 870 2341 916 2352
rect 1120 2438 1138 2456
rect 1074 2341 1120 2352
rect 1482 2566 1528 2577
rect 1456 2484 1482 2498
rect 1686 2566 1732 2697
rect 1456 2425 1471 2484
rect 1456 2407 1482 2425
rect 1278 2157 1324 2352
rect 1528 2407 1541 2498
rect 1482 2341 1528 2352
rect 1890 2566 1936 2577
rect 1873 2494 1890 2508
rect 2094 2566 2140 2577
rect 1936 2494 1958 2508
rect 1873 2435 1888 2494
rect 1943 2435 1958 2494
rect 1873 2417 1890 2435
rect 1686 2341 1732 2352
rect 1936 2417 1958 2435
rect 1890 2341 1936 2352
rect 2298 2566 2344 2577
rect 2281 2507 2298 2521
rect 2502 2566 2548 2697
rect 2344 2507 2366 2521
rect 2281 2448 2296 2507
rect 2351 2448 2366 2507
rect 2281 2430 2298 2448
rect 2094 2157 2140 2352
rect 2344 2430 2366 2448
rect 2298 2341 2344 2352
rect 2706 2566 2752 2577
rect 2681 2509 2706 2523
rect 2910 2566 2956 2577
rect 2681 2450 2696 2509
rect 2681 2432 2706 2450
rect 2502 2341 2548 2352
rect 2752 2432 2766 2523
rect 2706 2341 2752 2352
rect 3114 2566 3160 2577
rect 3096 2510 3114 2524
rect 3318 2566 3364 2697
rect 3160 2510 3181 2524
rect 3096 2451 3111 2510
rect 3166 2451 3181 2510
rect 3096 2433 3114 2451
rect 2910 2157 2956 2352
rect 3160 2433 3181 2451
rect 3114 2341 3160 2352
rect 3522 2566 3568 2577
rect 3504 2497 3522 2511
rect 3726 2566 3772 2577
rect 3568 2497 3589 2511
rect 3504 2438 3519 2497
rect 3574 2438 3589 2497
rect 3504 2420 3522 2438
rect 3318 2341 3364 2352
rect 3568 2420 3589 2438
rect 3522 2341 3568 2352
rect 3726 2157 3772 2352
rect -2839 2128 3876 2157
rect -2839 1997 -2795 2128
rect -2650 1997 -2495 2128
rect -2350 1997 -2195 2128
rect -2050 1997 -1895 2128
rect -1750 1997 -1595 2128
rect -1450 1997 -1295 2128
rect -1150 1997 -995 2128
rect -850 1997 -695 2128
rect -550 1997 -395 2128
rect -250 1997 -95 2128
rect 50 1997 205 2128
rect 350 1997 505 2128
rect 650 1997 805 2128
rect 950 1997 1105 2128
rect 1250 1997 1405 2128
rect 1550 1997 1705 2128
rect 1850 1997 2005 2128
rect 2150 1997 2305 2128
rect 2450 1997 2605 2128
rect 2750 1997 2905 2128
rect 3050 1997 3205 2128
rect 3350 1997 3505 2128
rect 3650 2092 3876 2128
rect 3650 2025 3742 2092
rect 3809 2025 3876 2092
rect 3650 1997 3876 2025
rect -2839 1970 3876 1997
<< via1 >>
rect 3661 7621 3716 7677
rect 3862 7618 3917 7674
rect 3659 7487 3714 7543
rect 3867 7482 3922 7538
rect 93 7047 147 7101
rect 642 6963 698 7019
rect 240 6785 296 6841
rect 1462 6963 1518 7019
rect 1051 6782 1107 6838
rect -78 6638 -24 6692
rect 533 6605 589 6661
rect -3203 6336 -3136 6403
rect 1057 6547 1113 6603
rect 1458 6712 1514 6768
rect 2278 6963 2334 7019
rect 1863 6782 1919 6838
rect 1866 6545 1922 6601
rect 3092 6963 3148 7019
rect 2273 6707 2329 6763
rect 2683 6782 2739 6838
rect 2685 6543 2741 6599
rect 3837 6742 3891 6796
rect 3502 6546 3556 6600
rect 92 6246 148 6302
rect 642 6166 698 6222
rect -1600 5946 -1544 6002
rect -1165 5966 -1151 6022
rect -1151 5966 -1109 6022
rect -1299 5809 -1243 5865
rect -621 5980 -565 6036
rect 240 5988 296 6044
rect 1462 6166 1518 6222
rect 1051 5985 1107 6041
rect -79 5831 -23 5887
rect 533 5808 589 5864
rect -3013 5563 -2948 5628
rect 1057 5750 1113 5806
rect 1458 5915 1514 5971
rect 2278 6166 2334 6222
rect 1863 5985 1919 6041
rect 1866 5748 1922 5804
rect 3092 6166 3148 6222
rect 2273 5910 2329 5966
rect 2683 5985 2739 6041
rect 2685 5746 2741 5802
rect 3836 5942 3892 5998
rect 3502 5749 3556 5803
rect -3203 5385 -3136 5452
rect 92 5450 148 5506
rect 642 5369 698 5425
rect -2215 5172 -2161 5226
rect -1009 5216 -955 5270
rect -1340 5120 -1286 5174
rect -1593 4984 -1539 5038
rect 240 5191 296 5247
rect 1462 5369 1518 5425
rect 1051 5188 1107 5244
rect -2088 4864 -2032 4920
rect -2284 4751 -2230 4805
rect -617 4961 -563 5015
rect -79 5039 -23 5095
rect 533 5011 589 5067
rect 1057 4953 1113 5009
rect 1458 5118 1514 5174
rect -238 4782 -182 4838
rect 2278 5369 2334 5425
rect 1863 5188 1919 5244
rect 1866 4951 1922 5007
rect 3092 5369 3148 5425
rect 2273 5113 2329 5169
rect 2683 5188 2739 5244
rect 2685 4949 2741 5005
rect 3836 5144 3892 5200
rect 3502 4952 3556 5006
rect -3012 4592 -2947 4657
rect 92 4655 148 4711
rect 642 4572 698 4628
rect -3203 4376 -3136 4444
rect 240 4394 296 4450
rect 1462 4572 1518 4628
rect 1051 4391 1107 4447
rect -2156 4061 -2102 4115
rect -79 4237 -23 4293
rect 533 4214 589 4270
rect -1594 4010 -1540 4064
rect -789 4002 -735 4056
rect -1315 3920 -1261 3974
rect 1057 4156 1113 4212
rect 1458 4321 1514 4377
rect 2278 4572 2334 4628
rect 1863 4391 1919 4447
rect 1866 4154 1922 4210
rect 3092 4572 3148 4628
rect 2273 4316 2329 4372
rect 2683 4391 2739 4447
rect 2685 4152 2741 4208
rect 3836 4346 3892 4402
rect 3502 4155 3556 4209
rect 92 3960 148 3963
rect 92 3909 95 3960
rect 95 3909 146 3960
rect 146 3909 148 3960
rect 92 3907 148 3909
rect 3790 3966 3844 4020
rect 3657 3898 3711 3952
rect 3917 3889 3971 3943
rect -3013 3620 -2946 3687
rect 4046 3454 4116 3524
rect 3728 3336 3817 3408
rect -2994 3251 -2938 3254
rect -2994 3202 -2989 3251
rect -2989 3202 -2941 3251
rect -2941 3202 -2938 3251
rect -2994 3198 -2938 3202
rect -2606 2944 -2598 3004
rect -2598 2944 -2552 3004
rect -2552 2944 -2549 3004
rect -2192 2949 -2190 3008
rect -2190 2949 -2144 3008
rect -2144 2949 -2137 3008
rect -1780 2943 -1736 3002
rect -1736 2943 -1725 3002
rect -1380 2949 -1374 3008
rect -1374 2949 -1328 3008
rect -1328 2949 -1325 3008
rect -967 2931 -966 2990
rect -966 2931 -920 2990
rect -920 2931 -912 2990
rect -557 2942 -512 3001
rect -512 2942 -502 3001
rect -160 2931 -150 2990
rect -150 2931 -105 2990
rect 255 2936 258 2995
rect 258 2936 304 2995
rect 304 2936 310 2995
rect 666 2939 712 2998
rect 712 2939 721 2998
rect 1076 2949 1120 3008
rect 1120 2949 1131 3008
rect 1481 2931 1482 2990
rect 1482 2931 1528 2990
rect 1528 2931 1536 2990
rect 1883 2931 1890 2990
rect 1890 2931 1936 2990
rect 1936 2931 1938 2990
rect 2299 2944 2344 3003
rect 2344 2944 2354 3003
rect 2699 2936 2706 2995
rect 2706 2936 2752 2995
rect 2752 2936 2754 2995
rect 3116 2933 3160 2992
rect 3160 2933 3171 2992
rect 3504 2939 3522 2998
rect 3522 2939 3559 2998
rect -2604 2440 -2598 2499
rect -2598 2440 -2552 2499
rect -2552 2440 -2549 2499
rect -2990 2231 -2933 2236
rect -2990 2180 -2989 2231
rect -2989 2180 -2941 2231
rect -2941 2180 -2933 2231
rect -2990 2179 -2933 2180
rect -2182 2445 -2144 2504
rect -2144 2445 -2127 2504
rect -1786 2461 -1782 2520
rect -1782 2461 -1736 2520
rect -1736 2461 -1731 2520
rect -1373 2466 -1328 2525
rect -1328 2466 -1318 2525
rect -973 2464 -966 2523
rect -966 2464 -920 2523
rect -920 2464 -918 2523
rect -570 2454 -558 2513
rect -558 2454 -515 2513
rect -147 2456 -104 2515
rect -104 2456 -92 2515
rect 253 2440 258 2499
rect 258 2440 304 2499
rect 304 2440 308 2499
rect 655 2441 666 2500
rect 666 2441 710 2500
rect 1068 2456 1074 2515
rect 1074 2456 1120 2515
rect 1120 2456 1123 2515
rect 1471 2425 1482 2484
rect 1482 2425 1526 2484
rect 1888 2435 1890 2494
rect 1890 2435 1936 2494
rect 1936 2435 1943 2494
rect 2296 2448 2298 2507
rect 2298 2448 2344 2507
rect 2344 2448 2351 2507
rect 2696 2450 2706 2509
rect 2706 2450 2751 2509
rect 3111 2451 3114 2510
rect 3114 2451 3160 2510
rect 3160 2451 3166 2510
rect 3519 2438 3522 2497
rect 3522 2438 3568 2497
rect 3568 2438 3574 2497
rect 3742 2025 3809 2092
<< metal2 >>
rect 3633 7677 3738 7695
rect 3633 7621 3661 7677
rect 3716 7621 3738 7677
rect 3633 7543 3738 7621
rect 3633 7487 3659 7543
rect 3714 7487 3738 7543
rect 81 7101 159 7113
rect 81 7047 93 7101
rect 147 7047 159 7101
rect 81 7039 159 7047
rect -90 6692 -12 6704
rect -90 6638 -78 6692
rect -24 6638 -12 6692
rect -90 6632 -12 6638
rect -3218 6403 -3122 6418
rect -3218 6336 -3203 6403
rect -3136 6336 -3122 6403
rect -3218 6330 -3122 6336
rect -3203 5473 -3136 6330
rect -1165 6031 -734 6057
rect -1176 6022 -734 6031
rect -1610 6002 -1534 6011
rect -2217 5946 -1600 6002
rect -1544 5946 -1534 6002
rect -1176 5966 -1165 6022
rect -1109 6001 -734 6022
rect -1109 5966 -1095 6001
rect -1176 5950 -1095 5966
rect -3025 5628 -2939 5643
rect -3025 5563 -3013 5628
rect -2948 5563 -2939 5628
rect -3025 5556 -2939 5563
rect -3218 5452 -3108 5473
rect -3218 5385 -3203 5452
rect -3136 5385 -3108 5452
rect -3218 5357 -3108 5385
rect -3203 4484 -3136 5357
rect -3013 4665 -2946 5556
rect -2217 5260 -2161 5946
rect -1610 5934 -1534 5946
rect -1315 5894 -1233 5903
rect -1315 5865 -954 5894
rect -1315 5809 -1299 5865
rect -1243 5838 -954 5865
rect -1243 5809 -1233 5838
rect -1315 5798 -1233 5809
rect -1010 5282 -954 5838
rect -1021 5270 -943 5282
rect -2217 5236 -2160 5260
rect -2227 5226 -2149 5236
rect -2227 5172 -2215 5226
rect -2161 5172 -2149 5226
rect -1021 5216 -1009 5270
rect -955 5216 -943 5270
rect -1021 5204 -943 5216
rect -2227 5160 -2149 5172
rect -1354 5175 -1271 5189
rect -1354 5119 -1341 5175
rect -1285 5119 -1271 5175
rect -1354 5105 -1271 5119
rect -1611 5038 -1527 5050
rect -1611 4984 -1593 5038
rect -1539 4984 -1527 5038
rect -1611 4978 -1527 4984
rect -1594 4947 -1537 4978
rect -2098 4920 -2028 4933
rect -2098 4864 -2088 4920
rect -2032 4864 -1912 4920
rect -2098 4852 -2028 4864
rect -2298 4805 -2215 4815
rect -2298 4792 -2284 4805
rect -2366 4751 -2284 4792
rect -2230 4751 -2215 4805
rect -2366 4741 -2215 4751
rect -2366 4736 -2254 4741
rect -3024 4657 -2943 4665
rect -3024 4592 -3012 4657
rect -2947 4592 -2943 4657
rect -3024 4587 -2943 4592
rect -3213 4444 -3124 4484
rect -3213 4376 -3203 4444
rect -3136 4376 -3124 4444
rect -3213 4364 -3124 4376
rect -3013 3697 -2946 4587
rect -2366 4241 -2310 4736
rect -2366 4185 -2101 4241
rect -2157 4127 -2101 4185
rect -2165 4115 -2090 4127
rect -2165 4061 -2156 4115
rect -2102 4061 -2090 4115
rect -2165 4049 -2090 4061
rect -1968 4065 -1912 4864
rect -1593 4728 -1537 4947
rect -1593 4672 -1260 4728
rect -1611 4065 -1528 4067
rect -1968 4064 -1528 4065
rect -1968 4010 -1594 4064
rect -1540 4010 -1528 4064
rect -1968 4009 -1528 4010
rect -1611 3997 -1528 4009
rect -1316 3981 -1260 4672
rect -790 4061 -734 6001
rect -634 6038 -553 6052
rect -79 6038 -23 6632
rect 92 6311 148 7039
rect 629 7019 711 7026
rect 1450 7019 1532 7026
rect 2266 7019 2348 7026
rect 3079 7019 3161 7026
rect 629 6963 642 7019
rect 698 6963 1462 7019
rect 1518 6963 2278 7019
rect 2334 6963 3092 7019
rect 3148 6963 3161 7019
rect 629 6951 711 6963
rect 1450 6951 1532 6963
rect 2266 6951 2348 6963
rect 3079 6951 3161 6963
rect 228 6841 310 6851
rect 228 6785 240 6841
rect 296 6838 310 6841
rect 1038 6838 1119 6848
rect 1852 6838 1933 6848
rect 2674 6838 2754 6850
rect 296 6785 1051 6838
rect 228 6782 1051 6785
rect 1107 6782 1863 6838
rect 1919 6782 2683 6838
rect 2739 6782 2754 6838
rect 228 6776 310 6782
rect 1038 6774 1119 6782
rect 1445 6768 1530 6782
rect 1852 6774 1933 6782
rect 1445 6712 1458 6768
rect 1514 6712 1530 6768
rect 1445 6702 1530 6712
rect 2260 6771 2347 6782
rect 2674 6774 2754 6782
rect 2260 6763 2345 6771
rect 2260 6707 2273 6763
rect 2329 6707 2345 6763
rect 2260 6699 2345 6707
rect 2273 6698 2329 6699
rect 523 6661 597 6673
rect 523 6605 533 6661
rect 589 6609 597 6661
rect 1042 6609 1124 6611
rect 1852 6609 1936 6614
rect 3092 6609 3148 6951
rect 3487 6610 3572 6612
rect 3633 6610 3738 7487
rect 3836 7674 3944 7693
rect 3836 7618 3862 7674
rect 3917 7618 3944 7674
rect 3836 7538 3944 7618
rect 3836 7482 3867 7538
rect 3922 7482 3944 7538
rect 3836 6812 3944 7482
rect 3824 6796 3944 6812
rect 3824 6742 3837 6796
rect 3891 6742 3944 6796
rect 3824 6736 3944 6742
rect 3487 6609 3738 6610
rect 589 6605 3738 6609
rect 523 6603 3738 6605
rect 523 6593 1057 6603
rect 524 6553 1057 6593
rect 1042 6547 1057 6553
rect 1113 6601 3738 6603
rect 1113 6553 1866 6601
rect 1113 6547 1124 6553
rect 1042 6539 1124 6547
rect 1852 6545 1866 6553
rect 1922 6600 3738 6601
rect 1922 6599 3502 6600
rect 1922 6553 2685 6599
rect 1922 6545 1936 6553
rect 1852 6537 1936 6545
rect 2672 6543 2685 6553
rect 2741 6553 3502 6599
rect 2741 6543 2754 6553
rect 2672 6532 2754 6543
rect 3487 6546 3502 6553
rect 3556 6554 3738 6600
rect 3556 6546 3572 6554
rect 3487 6532 3572 6546
rect 80 6302 158 6311
rect 80 6246 92 6302
rect 148 6246 158 6302
rect 80 6237 158 6246
rect -634 6036 -23 6038
rect -634 5980 -621 6036
rect -565 5982 -23 6036
rect -565 5980 -553 5982
rect -634 5970 -553 5980
rect -621 5184 -565 5970
rect -79 5894 -23 5982
rect -93 5887 -15 5894
rect -93 5831 -79 5887
rect -23 5831 -15 5887
rect -93 5822 -15 5831
rect -630 5175 -554 5184
rect -630 5119 -621 5175
rect -565 5119 -554 5175
rect -630 5107 -554 5119
rect -79 5101 -23 5822
rect 92 5517 148 6237
rect 629 6222 711 6229
rect 1450 6222 1532 6229
rect 2266 6222 2348 6229
rect 3079 6222 3161 6229
rect 629 6166 642 6222
rect 698 6166 1462 6222
rect 1518 6166 2278 6222
rect 2334 6166 3092 6222
rect 3148 6166 3161 6222
rect 629 6154 711 6166
rect 1450 6154 1532 6166
rect 2266 6154 2348 6166
rect 3079 6154 3161 6166
rect 228 6044 310 6054
rect 228 5988 240 6044
rect 296 6041 310 6044
rect 1038 6041 1119 6051
rect 1852 6041 1933 6051
rect 2674 6041 2754 6053
rect 296 5988 1051 6041
rect 228 5985 1051 5988
rect 1107 5985 1863 6041
rect 1919 5985 2683 6041
rect 2739 5985 2754 6041
rect 228 5979 310 5985
rect 1038 5977 1119 5985
rect 1445 5971 1530 5985
rect 1852 5977 1933 5985
rect 1445 5915 1458 5971
rect 1514 5915 1530 5971
rect 1445 5905 1530 5915
rect 2260 5974 2347 5985
rect 2674 5977 2754 5985
rect 2260 5966 2345 5974
rect 2260 5910 2273 5966
rect 2329 5910 2345 5966
rect 2260 5902 2345 5910
rect 2273 5901 2329 5902
rect 523 5864 597 5876
rect 523 5808 533 5864
rect 589 5812 597 5864
rect 1042 5812 1124 5814
rect 1852 5812 1936 5817
rect 3092 5812 3148 6154
rect 3487 5812 3572 5815
rect 589 5808 3572 5812
rect 3633 5808 3738 6554
rect 3836 6009 3944 6736
rect 3824 5998 3944 6009
rect 3824 5942 3836 5998
rect 3892 5942 3944 5998
rect 3824 5933 3944 5942
rect 523 5806 3738 5808
rect 523 5796 1057 5806
rect 524 5756 1057 5796
rect 1042 5750 1057 5756
rect 1113 5804 3738 5806
rect 1113 5756 1866 5804
rect 1113 5750 1124 5756
rect 1042 5742 1124 5750
rect 1852 5748 1866 5756
rect 1922 5803 3738 5804
rect 1922 5802 3502 5803
rect 1922 5756 2685 5802
rect 1922 5748 1936 5756
rect 1852 5740 1936 5748
rect 2672 5746 2685 5756
rect 2741 5756 3502 5802
rect 2741 5746 2754 5756
rect 2672 5735 2754 5746
rect 3487 5749 3502 5756
rect 3556 5752 3738 5803
rect 3556 5749 3572 5752
rect 3487 5735 3572 5749
rect 80 5506 158 5517
rect 80 5450 92 5506
rect 148 5450 158 5506
rect 80 5443 158 5450
rect -94 5095 -11 5101
rect -94 5039 -79 5095
rect -23 5039 -11 5095
rect -94 5029 -11 5039
rect -630 5015 -551 5027
rect -630 4961 -617 5015
rect -563 4961 -551 5015
rect -630 4954 -551 4961
rect -618 4838 -562 4954
rect -245 4838 -173 4852
rect -618 4782 -238 4838
rect -182 4782 -173 4838
rect -245 4774 -173 4782
rect -245 4770 -175 4774
rect -79 4300 -23 5029
rect 92 4721 148 5443
rect 629 5425 711 5432
rect 1450 5425 1532 5432
rect 2266 5425 2348 5432
rect 3079 5425 3161 5432
rect 629 5369 642 5425
rect 698 5369 1462 5425
rect 1518 5369 2278 5425
rect 2334 5369 3092 5425
rect 3148 5369 3161 5425
rect 629 5357 711 5369
rect 1450 5357 1532 5369
rect 2266 5357 2348 5369
rect 3079 5357 3161 5369
rect 228 5247 310 5257
rect 228 5191 240 5247
rect 296 5244 310 5247
rect 1038 5244 1119 5254
rect 1852 5244 1933 5254
rect 2674 5244 2754 5256
rect 296 5191 1051 5244
rect 228 5188 1051 5191
rect 1107 5188 1863 5244
rect 1919 5188 2683 5244
rect 2739 5188 2754 5244
rect 228 5182 310 5188
rect 1038 5180 1119 5188
rect 1445 5174 1530 5188
rect 1852 5180 1933 5188
rect 1445 5118 1458 5174
rect 1514 5118 1530 5174
rect 1445 5108 1530 5118
rect 2260 5177 2347 5188
rect 2674 5180 2754 5188
rect 2260 5169 2345 5177
rect 2260 5113 2273 5169
rect 2329 5113 2345 5169
rect 2260 5105 2345 5113
rect 2273 5104 2329 5105
rect 523 5067 597 5079
rect 523 5011 533 5067
rect 589 5015 597 5067
rect 1042 5015 1124 5017
rect 1852 5015 1936 5020
rect 3092 5015 3148 5357
rect 3487 5015 3572 5018
rect 589 5011 3572 5015
rect 523 5009 3572 5011
rect 523 4999 1057 5009
rect 524 4959 1057 4999
rect 1042 4953 1057 4959
rect 1113 5008 3572 5009
rect 3633 5008 3738 5752
rect 3836 5213 3944 5933
rect 3822 5200 3944 5213
rect 3822 5144 3836 5200
rect 3892 5144 3944 5200
rect 3822 5137 3944 5144
rect 1113 5007 3738 5008
rect 1113 4959 1866 5007
rect 1113 4953 1124 4959
rect 1042 4945 1124 4953
rect 1852 4951 1866 4959
rect 1922 5006 3738 5007
rect 1922 5005 3502 5006
rect 1922 4959 2685 5005
rect 1922 4951 1936 4959
rect 1852 4943 1936 4951
rect 2672 4949 2685 4959
rect 2741 4959 3502 5005
rect 2741 4949 2754 4959
rect 2672 4938 2754 4949
rect 3487 4952 3502 4959
rect 3556 4952 3738 5006
rect 3487 4938 3572 4952
rect 78 4711 156 4721
rect 78 4655 92 4711
rect 148 4655 156 4711
rect 78 4647 156 4655
rect -92 4293 -10 4300
rect -92 4237 -79 4293
rect -23 4237 -10 4293
rect -92 4228 -10 4237
rect -802 4056 -725 4061
rect -802 4002 -789 4056
rect -735 4002 -725 4056
rect -802 3990 -725 4002
rect 92 3981 148 4647
rect 629 4628 711 4635
rect 1450 4628 1532 4635
rect 2266 4628 2348 4635
rect 3079 4628 3161 4635
rect 629 4572 642 4628
rect 698 4572 1462 4628
rect 1518 4572 2278 4628
rect 2334 4572 3092 4628
rect 3148 4572 3161 4628
rect 629 4560 711 4572
rect 1450 4560 1532 4572
rect 2266 4560 2348 4572
rect 3079 4560 3161 4572
rect 228 4450 310 4460
rect 228 4394 240 4450
rect 296 4447 310 4450
rect 1038 4447 1119 4457
rect 1852 4447 1933 4457
rect 2674 4447 2754 4459
rect 296 4394 1051 4447
rect 228 4391 1051 4394
rect 1107 4391 1863 4447
rect 1919 4391 2683 4447
rect 2739 4391 2754 4447
rect 228 4385 310 4391
rect 1038 4383 1119 4391
rect 1445 4377 1530 4391
rect 1852 4383 1933 4391
rect 1445 4321 1458 4377
rect 1514 4321 1530 4377
rect 1445 4311 1530 4321
rect 2260 4380 2347 4391
rect 2674 4383 2754 4391
rect 2260 4372 2345 4380
rect 2260 4316 2273 4372
rect 2329 4316 2345 4372
rect 2260 4308 2345 4316
rect 2273 4307 2329 4308
rect 523 4270 597 4282
rect 523 4214 533 4270
rect 589 4218 597 4270
rect 1042 4218 1124 4220
rect 1852 4218 1936 4223
rect 3092 4218 3148 4560
rect 3487 4218 3572 4221
rect 589 4214 3572 4218
rect 523 4212 3572 4214
rect 523 4202 1057 4212
rect 524 4162 1057 4202
rect 1042 4156 1057 4162
rect 1113 4210 3572 4212
rect 1113 4162 1866 4210
rect 1113 4156 1124 4162
rect 1042 4148 1124 4156
rect 1852 4154 1866 4162
rect 1922 4209 3572 4210
rect 1922 4208 3502 4209
rect 1922 4162 2685 4208
rect 1922 4154 1936 4162
rect 1852 4146 1936 4154
rect 2672 4152 2685 4162
rect 2741 4162 3502 4208
rect 2741 4152 2754 4162
rect 2672 4141 2754 4152
rect 3487 4155 3502 4162
rect 3556 4208 3572 4209
rect 3633 4208 3738 4952
rect 3836 4413 3944 5137
rect 3826 4402 3944 4413
rect 3826 4346 3836 4402
rect 3892 4357 3944 4402
rect 3892 4346 3908 4357
rect 3826 4337 3908 4346
rect 3556 4155 3738 4208
rect 3487 4152 3738 4155
rect 3487 4141 3572 4152
rect 3605 4020 4117 4043
rect -1328 3974 -1259 3981
rect -1328 3920 -1315 3974
rect -1261 3920 -1259 3974
rect -1328 3906 -1259 3920
rect 75 3963 167 3981
rect 75 3907 92 3963
rect 148 3907 167 3963
rect 75 3889 167 3907
rect 3605 3966 3790 4020
rect 3844 3966 4117 4020
rect 3605 3952 4117 3966
rect 3605 3898 3657 3952
rect 3711 3943 4117 3952
rect 3711 3898 3917 3943
rect 3605 3889 3917 3898
rect 3971 3889 4117 3943
rect 3605 3870 4117 3889
rect -3025 3687 -2932 3697
rect -3025 3620 -3013 3687
rect -2946 3620 -2932 3687
rect -3025 3608 -2932 3620
rect 4045 3540 4117 3870
rect 4031 3524 4129 3540
rect 4031 3454 4046 3524
rect 4116 3454 4129 3524
rect 4031 3444 4129 3454
rect 3708 3408 3847 3435
rect 3708 3336 3728 3408
rect 3817 3336 3847 3408
rect 3708 3311 3847 3336
rect -3007 3254 -2921 3269
rect -3007 3198 -2994 3254
rect -2938 3198 -2921 3254
rect -3007 3186 -2921 3198
rect -2995 2252 -2937 3186
rect -2620 3004 -2535 3021
rect -2620 2944 -2606 3004
rect -2549 2944 -2535 3004
rect -2620 2930 -2535 2944
rect -2207 3008 -2122 3022
rect -2207 2949 -2192 3008
rect -2137 2949 -2122 3008
rect -2207 2931 -2122 2949
rect -1795 3002 -1710 3016
rect -1795 2943 -1780 3002
rect -1725 2943 -1710 3002
rect -2606 2516 -2549 2930
rect -2189 2518 -2132 2931
rect -1795 2926 -1710 2943
rect -1395 3008 -1310 3022
rect -1395 2949 -1380 3008
rect -1325 2949 -1310 3008
rect -1395 2931 -1310 2949
rect -982 2990 -897 3004
rect -982 2931 -967 2990
rect -912 2931 -897 2990
rect -1781 2534 -1724 2926
rect -1380 2539 -1323 2931
rect -982 2913 -897 2931
rect -572 3001 -487 3015
rect -572 2942 -557 3001
rect -502 2942 -487 3001
rect -572 2924 -487 2942
rect -175 2990 -90 3004
rect -175 2931 -160 2990
rect -105 2931 -90 2990
rect -1801 2520 -1716 2534
rect -2618 2514 -2533 2516
rect -2197 2514 -2112 2518
rect -1801 2514 -1786 2520
rect -2618 2504 -1786 2514
rect -2618 2499 -2182 2504
rect -2618 2440 -2604 2499
rect -2549 2457 -2182 2499
rect -2549 2440 -2533 2457
rect -2618 2425 -2533 2440
rect -2197 2445 -2182 2457
rect -2127 2461 -1786 2504
rect -1731 2514 -1716 2520
rect -1388 2525 -1303 2539
rect -972 2537 -915 2913
rect -1388 2514 -1373 2525
rect -1731 2466 -1373 2514
rect -1318 2514 -1303 2525
rect -988 2523 -903 2537
rect -569 2527 -512 2924
rect -175 2913 -90 2931
rect 240 2995 325 3009
rect 240 2936 255 2995
rect 310 2936 325 2995
rect 240 2918 325 2936
rect 651 2998 736 3012
rect 651 2939 666 2998
rect 721 2939 736 2998
rect 651 2921 736 2939
rect 1061 3008 1146 3022
rect 1061 2949 1076 3008
rect 1131 2949 1146 3008
rect 1061 2931 1146 2949
rect 1466 2990 1551 3004
rect 1466 2931 1481 2990
rect 1536 2931 1551 2990
rect -155 2529 -98 2913
rect -988 2514 -973 2523
rect -1318 2466 -973 2514
rect -1731 2464 -973 2466
rect -918 2514 -903 2523
rect -585 2514 -500 2527
rect -162 2515 -77 2529
rect -162 2514 -147 2515
rect -918 2513 -147 2514
rect -918 2464 -570 2513
rect -1731 2461 -570 2464
rect -2127 2457 -570 2461
rect -2127 2445 -2112 2457
rect -2197 2427 -2112 2445
rect -1801 2443 -1716 2457
rect -1388 2448 -1303 2457
rect -988 2446 -903 2457
rect -585 2454 -570 2457
rect -515 2457 -147 2513
rect -515 2454 -500 2457
rect -585 2436 -500 2454
rect -162 2456 -147 2457
rect -92 2514 -77 2515
rect 254 2514 311 2918
rect 656 2514 713 2921
rect 1070 2529 1127 2931
rect 1466 2913 1551 2931
rect 1868 2990 1953 3004
rect 1868 2931 1883 2990
rect 1938 2931 1953 2990
rect 1868 2913 1953 2931
rect 2284 3003 2369 3017
rect 2284 2944 2299 3003
rect 2354 2944 2369 3003
rect 2284 2926 2369 2944
rect 2684 2995 2769 3009
rect 2684 2936 2699 2995
rect 2754 2936 2769 2995
rect 1053 2515 1138 2529
rect 1053 2514 1068 2515
rect -92 2500 1068 2514
rect -92 2499 655 2500
rect -92 2457 253 2499
rect -92 2456 -77 2457
rect -162 2438 -77 2456
rect 238 2440 253 2457
rect 308 2457 655 2499
rect 308 2440 323 2457
rect 238 2422 323 2440
rect 640 2441 655 2457
rect 710 2457 1068 2500
rect 710 2441 725 2457
rect 640 2423 725 2441
rect 1053 2456 1068 2457
rect 1123 2514 1138 2515
rect 1472 2514 1529 2913
rect 1880 2514 1937 2913
rect 2289 2521 2346 2926
rect 2684 2918 2769 2936
rect 3101 2992 3186 3006
rect 3101 2933 3116 2992
rect 3171 2933 3186 2992
rect 2687 2523 2744 2918
rect 3101 2915 3186 2933
rect 3489 2998 3574 3012
rect 3489 2939 3504 2998
rect 3559 2939 3574 2998
rect 3489 2921 3574 2939
rect 3103 2524 3160 2915
rect 2281 2514 2366 2521
rect 2681 2514 2766 2523
rect 3096 2514 3181 2524
rect 3506 2514 3563 2921
rect 1123 2511 3563 2514
rect 1123 2510 3589 2511
rect 1123 2509 3111 2510
rect 1123 2507 2696 2509
rect 1123 2494 2296 2507
rect 1123 2484 1888 2494
rect 1123 2457 1471 2484
rect 1123 2456 1138 2457
rect 1053 2438 1138 2456
rect 1456 2425 1471 2457
rect 1526 2457 1888 2484
rect 1526 2425 1541 2457
rect 1456 2407 1541 2425
rect 1873 2435 1888 2457
rect 1943 2457 2296 2494
rect 1943 2435 1958 2457
rect 1873 2417 1958 2435
rect 2281 2448 2296 2457
rect 2351 2457 2696 2507
rect 2351 2448 2366 2457
rect 2281 2430 2366 2448
rect 2681 2450 2696 2457
rect 2751 2457 3111 2509
rect 2751 2450 2766 2457
rect 2681 2432 2766 2450
rect 3096 2451 3111 2457
rect 3166 2497 3589 2510
rect 3166 2457 3519 2497
rect 3166 2451 3181 2457
rect 3096 2433 3181 2451
rect 3504 2438 3519 2457
rect 3574 2438 3589 2497
rect 3504 2420 3589 2438
rect -3005 2236 -2913 2252
rect -3005 2179 -2990 2236
rect -2933 2179 -2913 2236
rect -3005 2164 -2913 2179
rect 3742 2103 3809 3311
rect 3725 2092 3828 2103
rect 3725 2025 3742 2092
rect 3809 2025 3828 2092
rect 3725 2010 3828 2025
<< via2 >>
rect -1341 5174 -1285 5175
rect -1341 5120 -1340 5174
rect -1340 5120 -1286 5174
rect -1286 5120 -1285 5174
rect -1341 5119 -1285 5120
rect -621 5119 -565 5175
<< metal3 >>
rect -1354 5175 -1271 5189
rect -630 5175 -554 5184
rect -1354 5119 -1341 5175
rect -1285 5119 -621 5175
rect -565 5119 -554 5175
rect -1354 5105 -1271 5119
rect -630 5107 -554 5119
<< labels >>
flabel metal1 -3384 3241 -3384 3241 0 FreeSans 1600 0 0 0 IM_T
port 0 nsew
flabel metal1 -3340 2694 -3340 2694 0 FreeSans 1600 0 0 0 IM
port 1 nsew
flabel metal1 -3423 3612 -3423 3612 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
flabel metal1 -3204 3981 -3204 3981 0 FreeSans 1600 0 0 0 Ri
port 3 nsew
flabel metal1 -3431 4954 -3431 4954 0 FreeSans 1600 0 0 0 Ci
port 4 nsew
flabel metal1 -3540 5919 -3540 5919 0 FreeSans 1600 0 0 0 Ri-1
port 5 nsew
flabel metal1 -3483 6325 -3483 6325 0 FreeSans 1600 0 0 0 VDD
port 6 nsew
flabel metal2 -517 6019 -517 6019 0 FreeSans 1600 0 0 0 QB
port 7 nsew
flabel via1 -589 4973 -589 4973 0 FreeSans 1600 0 0 0 Q
port 8 nsew
flabel metal1 4074 2797 4074 2797 0 FreeSans 1600 0 0 0 OUT
port 9 nsew
flabel via1 3898 7510 3898 7510 0 FreeSans 1600 0 0 0 OUT+
port 10 nsew
flabel via1 3681 7653 3681 7653 0 FreeSans 1600 0 0 0 OUT-
port 11 nsew
flabel metal2 -540 2480 -540 2480 0 FreeSans 1600 0 0 0 SD
port 12 nsew
flabel metal1 -2821 5929 -2821 5929 0 FreeSans 480 0 0 0 Local_Enc_0.Ri-1
flabel metal1 -1816 6393 -1816 6393 0 FreeSans 480 0 0 0 Local_Enc_0.VDD
flabel metal1 -1812 5606 -1812 5606 0 FreeSans 480 0 0 0 Local_Enc_0.VSS
flabel metal1 -592 4986 -592 4986 0 FreeSans 480 0 0 0 Local_Enc_0.Q
flabel metal1 -518 6013 -518 6013 0 FreeSans 480 0 0 0 Local_Enc_0.QB
flabel metal1 -2821 4951 -2821 4951 0 FreeSans 480 0 0 0 Local_Enc_0.Ci
flabel metal1 -2822 3978 -2822 3978 0 FreeSans 480 0 0 0 Local_Enc_0.Ri
flabel nsubdiffcont -996 5417 -996 5417 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_8.VDD
flabel psubdiffcont -987 4625 -987 4625 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_8.VSS
flabel metal1 -1236 5003 -1236 5003 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_8.B
flabel metal1 -1233 4905 -1233 4905 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_8.A
flabel metal1 -734 5049 -734 5049 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_8.OUT
flabel metal1 -985 4782 -985 4782 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_8.SD
flabel nsubdiffcont -996 4441 -996 4441 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_7.VDD
flabel psubdiffcont -987 3649 -987 3649 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_7.VSS
flabel metal1 -1236 4027 -1236 4027 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_7.B
flabel metal1 -1233 3929 -1233 3929 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_7.A
flabel metal1 -734 4073 -734 4073 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_7.OUT
flabel metal1 -985 3806 -985 3806 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_7.SD
flabel nsubdiffcont -1807 4441 -1807 4441 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_6.VDD
flabel psubdiffcont -1798 3649 -1798 3649 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_6.VSS
flabel metal1 -2047 4027 -2047 4027 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_6.B
flabel metal1 -2044 3929 -2044 3929 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_6.A
flabel metal1 -1545 4073 -1545 4073 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_6.OUT
flabel metal1 -1796 3806 -1796 3806 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_6.SD
flabel nsubdiffcont -1807 5417 -1807 5417 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_5.VDD
flabel psubdiffcont -1798 4625 -1798 4625 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_5.VSS
flabel metal1 -2047 5003 -2047 5003 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_5.B
flabel metal1 -2044 4905 -2044 4905 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_5.A
flabel metal1 -1545 5049 -1545 5049 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_5.OUT
flabel metal1 -1796 4782 -1796 4782 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_5.SD
flabel nsubdiffcont -996 6388 -996 6388 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_4.VDD
flabel psubdiffcont -987 5596 -987 5596 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_4.VSS
flabel metal1 -1236 5974 -1236 5974 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_4.B
flabel metal1 -1233 5876 -1233 5876 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_4.A
flabel metal1 -734 6020 -734 6020 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_4.OUT
flabel metal1 -985 5753 -985 5753 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_4.SD
flabel nsubdiffcont -2570 4442 -2570 4442 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_3.VDD
flabel psubdiffcont -2561 3650 -2561 3650 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_3.VSS
flabel metal1 -2810 4028 -2810 4028 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_3.B
flabel metal1 -2807 3930 -2807 3930 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_3.A
flabel metal1 -2308 4074 -2308 4074 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_3.OUT
flabel metal1 -2559 3807 -2559 3807 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_3.SD
flabel nsubdiffcont -2570 5417 -2570 5417 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_2.VDD
flabel psubdiffcont -2561 4625 -2561 4625 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_2.VSS
flabel metal1 -2810 5003 -2810 5003 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_2.B
flabel metal1 -2807 4905 -2807 4905 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_2.A
flabel metal1 -2308 5049 -2308 5049 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_2.OUT
flabel metal1 -2559 4782 -2559 4782 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_2.SD
flabel nsubdiffcont -1807 6388 -1807 6388 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_1.VDD
flabel psubdiffcont -1798 5596 -1798 5596 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_1.VSS
flabel metal1 -2047 5974 -2047 5974 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_1.B
flabel metal1 -2044 5876 -2044 5876 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_1.A
flabel metal1 -1545 6020 -1545 6020 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_1.OUT
flabel metal1 -1796 5753 -1796 5753 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_1.SD
flabel nsubdiffcont -2570 6388 -2570 6388 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_0.VDD
flabel psubdiffcont -2561 5596 -2561 5596 0 FreeSans 320 0 0 0 Local_Enc_0.NAND_0.VSS
flabel metal1 -2810 5974 -2810 5974 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_0.B
flabel metal1 -2807 5876 -2807 5876 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_0.A
flabel metal1 -2308 6020 -2308 6020 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_0.OUT
flabel metal1 -2559 5753 -2559 5753 0 FreeSans 480 0 0 0 Local_Enc_0.NAND_0.SD
flabel via1 -2972 3227 -2972 3227 0 FreeSans 1600 0 0 0 CM_MSB_V2_0.IM_T
flabel metal1 -1359 3370 -1359 3370 0 FreeSans 1600 0 0 0 CM_MSB_V2_0.VSS
flabel metal1 4018 2734 4018 2734 0 FreeSans 1600 0 0 0 CM_MSB_V2_0.OUT
flabel metal1 -3003 2698 -3003 2698 0 FreeSans 1600 0 0 0 CM_MSB_V2_0.IM
flabel via1 -549 2488 -549 2488 0 FreeSans 1600 0 0 0 CM_MSB_V2_0.SD
<< end >>
