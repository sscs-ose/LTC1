magic
tech gf180mcuD
magscale 1 10
timestamp 1713338890
<< checkpaint >>
rect -6181 -2045 6181 2045
<< psubdiff >>
rect -4181 23 4181 45
rect -4181 -23 -4159 23
rect 4159 -23 4181 23
rect -4181 -45 4181 -23
<< psubdiffcont >>
rect -4159 -23 4159 23
<< metal1 >>
rect -4170 23 4170 34
rect -4170 -23 -4159 23
rect 4159 -23 4170 23
rect -4170 -34 4170 -23
<< end >>
